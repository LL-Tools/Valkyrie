

module b17_C_gen_AntiSAT_k_256_1 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput_f0, keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, 
        keyinput_f5, keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, 
        keyinput_f10, keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, 
        keyinput_f15, keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, 
        keyinput_f20, keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, 
        keyinput_f25, keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, 
        keyinput_f30, keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, 
        keyinput_f35, keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, 
        keyinput_f40, keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, 
        keyinput_f45, keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, 
        keyinput_f50, keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, 
        keyinput_f55, keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, 
        keyinput_f60, keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, 
        keyinput_f65, keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, 
        keyinput_f70, keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, 
        keyinput_f75, keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, 
        keyinput_f80, keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, 
        keyinput_f85, keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, 
        keyinput_f90, keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, 
        keyinput_f95, keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, 
        keyinput_f100, keyinput_f101, keyinput_f102, keyinput_f103, 
        keyinput_f104, keyinput_f105, keyinput_f106, keyinput_f107, 
        keyinput_f108, keyinput_f109, keyinput_f110, keyinput_f111, 
        keyinput_f112, keyinput_f113, keyinput_f114, keyinput_f115, 
        keyinput_f116, keyinput_f117, keyinput_f118, keyinput_f119, 
        keyinput_f120, keyinput_f121, keyinput_f122, keyinput_f123, 
        keyinput_f124, keyinput_f125, keyinput_f126, keyinput_f127, 
        keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3, keyinput_g4, 
        keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8, keyinput_g9, 
        keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13, keyinput_g14, 
        keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18, keyinput_g19, 
        keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23, keyinput_g24, 
        keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28, keyinput_g29, 
        keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33, keyinput_g34, 
        keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38, keyinput_g39, 
        keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43, keyinput_g44, 
        keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48, keyinput_g49, 
        keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53, keyinput_g54, 
        keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58, keyinput_g59, 
        keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63, keyinput_g64, 
        keyinput_g65, keyinput_g66, keyinput_g67, keyinput_g68, keyinput_g69, 
        keyinput_g70, keyinput_g71, keyinput_g72, keyinput_g73, keyinput_g74, 
        keyinput_g75, keyinput_g76, keyinput_g77, keyinput_g78, keyinput_g79, 
        keyinput_g80, keyinput_g81, keyinput_g82, keyinput_g83, keyinput_g84, 
        keyinput_g85, keyinput_g86, keyinput_g87, keyinput_g88, keyinput_g89, 
        keyinput_g90, keyinput_g91, keyinput_g92, keyinput_g93, keyinput_g94, 
        keyinput_g95, keyinput_g96, keyinput_g97, keyinput_g98, keyinput_g99, 
        keyinput_g100, keyinput_g101, keyinput_g102, keyinput_g103, 
        keyinput_g104, keyinput_g105, keyinput_g106, keyinput_g107, 
        keyinput_g108, keyinput_g109, keyinput_g110, keyinput_g111, 
        keyinput_g112, keyinput_g113, keyinput_g114, keyinput_g115, 
        keyinput_g116, keyinput_g117, keyinput_g118, keyinput_g119, 
        keyinput_g120, keyinput_g121, keyinput_g122, keyinput_g123, 
        keyinput_g124, keyinput_g125, keyinput_g126, keyinput_g127, U355, U356, 
        U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, U369, 
        U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, U352, 
        U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, U240, 
        U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, U228, 
        U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, U216, 
        U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, U262, 
        U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, U274, 
        U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, 
        P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, 
        P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, 
        P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, 
        P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, 
        P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, 
        P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, 
        P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, 
        P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, 
        P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, 
        P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, 
        P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, 
        P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, 
        P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, 
        P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, 
        P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, 
        P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, 
        P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, 
        P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, 
        P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, 
        P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, 
        P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, 
        P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, 
        P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, 
        P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, 
        P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, 
        P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, 
        P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, 
        P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, 
        P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, 
        P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, 
        P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, 
        P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, 
        P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, 
        P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, 
        P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, 
        P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, 
        P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, 
        P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, 
        P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, 
        P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, 
        P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, 
        P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, 
        P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, 
        P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, 
        P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, 
        P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, 
        P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, 
        P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, 
        P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, 
        P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, 
        P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, 
        P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, 
        P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, 
        P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, 
        P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, 
        P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, 
        P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, 
        P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, 
        P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, 
        P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, 
        P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, 
        P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, 
        P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, 
        P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, 
        P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, 
        P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, 
        P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, 
        P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, 
        P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, 
        P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, 
        P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, 
        P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, 
        P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, 
        P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, 
        P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, 
        P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, 
        P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, 
        P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, 
        P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, 
        P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, 
        P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, 
        P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, 
        P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, 
        P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, 
        P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, 
        P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, 
        P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, 
        P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, 
        P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, 
        P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, 
        P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, 
        P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, 
        P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, 
        P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, 
        P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, 
        P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, 
        P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, 
        P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, 
        P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, 
        P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, 
        P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, 
        P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, 
        P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, 
        P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, 
        P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, 
        P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, 
        P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, 
        P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, 
        P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, 
        P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, 
        P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, 
        P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, 
        P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, 
        P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, 
        P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, 
        P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, 
        P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, 
        P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, 
        P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, 
        P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, 
        P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, 
        P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, 
        P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, 
        P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, 
        P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, 
        P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, 
        P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, 
        P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, 
        P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, 
        P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, 
        P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, 
        P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, 
        P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, 
        P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, 
        P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, 
        P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, 
        P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, 
        P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, 
        P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, 
        P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, 
        P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, 
        P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, 
        P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, 
        P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, 
        P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, 
        P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, 
        P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, 
        P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, 
        P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, 
        P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, 
        P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, 
        P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, 
        P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, 
        P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, 
        P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, 
        P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, 
        P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, 
        P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, 
        P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, 
        P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, 
        P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, 
        P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, 
        P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, 
        P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, 
        P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, 
        P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, 
        P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, 
        P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, 
        P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, 
        P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, 
        P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, 
        P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, 
        P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, 
        P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, 
        P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, 
        P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, 
        P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, 
        P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, 
        P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, 
        P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, 
        P1_U2802, P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,
         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
         n16611, n16612, n16614, n16615, n16616, n16617, n16618, n16619,
         n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627,
         n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635,
         n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643,
         n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651,
         n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659,
         n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
         n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675,
         n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683,
         n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691,
         n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699,
         n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707,
         n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715,
         n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723,
         n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731,
         n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739,
         n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747,
         n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755,
         n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763,
         n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771,
         n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779,
         n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787,
         n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795,
         n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803,
         n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811,
         n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819,
         n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827,
         n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835,
         n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843,
         n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851,
         n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859,
         n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
         n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875,
         n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883,
         n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891,
         n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899,
         n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
         n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915,
         n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
         n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931,
         n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
         n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947,
         n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
         n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
         n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971,
         n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
         n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987,
         n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995,
         n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
         n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011,
         n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019,
         n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
         n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
         n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043,
         n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051,
         n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059,
         n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067,
         n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075,
         n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083,
         n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091,
         n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
         n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
         n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115,
         n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123,
         n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131,
         n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139,
         n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
         n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
         n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163,
         n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
         n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
         n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187,
         n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195,
         n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203,
         n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211,
         n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
         n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227,
         n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235,
         n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
         n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
         n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
         n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
         n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323,
         n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331,
         n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339,
         n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
         n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355,
         n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
         n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
         n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379,
         n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
         n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395,
         n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403,
         n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
         n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
         n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
         n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435,
         n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
         n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451,
         n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
         n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467,
         n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475,
         n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483,
         n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
         n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499,
         n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507,
         n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515,
         n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523,
         n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
         n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539,
         n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
         n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
         n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
         n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579,
         n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
         n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595,
         n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
         n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611,
         n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619,
         n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627,
         n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635,
         n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643,
         n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651,
         n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659,
         n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667,
         n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
         n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683,
         n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691,
         n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699,
         n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
         n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715,
         n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723,
         n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731,
         n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739,
         n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747,
         n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755,
         n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763,
         n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771,
         n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779,
         n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787,
         n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795,
         n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
         n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811,
         n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
         n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827,
         n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835,
         n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843,
         n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851,
         n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859,
         n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867,
         n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875,
         n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883,
         n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891,
         n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899,
         n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907,
         n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915,
         n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923,
         n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931,
         n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939,
         n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947,
         n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955,
         n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963,
         n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971,
         n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979,
         n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987,
         n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995,
         n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003,
         n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011,
         n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019,
         n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027,
         n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035,
         n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043,
         n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051,
         n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059,
         n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067,
         n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075,
         n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083,
         n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091,
         n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099,
         n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107,
         n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115,
         n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123,
         n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131,
         n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139,
         n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147,
         n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155,
         n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163,
         n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171,
         n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179,
         n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187,
         n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195,
         n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203,
         n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211,
         n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219,
         n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227,
         n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
         n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243,
         n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
         n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259,
         n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267,
         n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275,
         n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283,
         n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291,
         n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299,
         n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
         n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315,
         n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323,
         n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331,
         n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339,
         n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347,
         n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355,
         n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363,
         n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371,
         n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
         n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387,
         n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395,
         n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403,
         n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411,
         n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419,
         n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427,
         n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435,
         n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443,
         n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
         n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459,
         n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467,
         n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475,
         n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483,
         n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491,
         n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499,
         n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507,
         n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515,
         n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523,
         n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531,
         n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539,
         n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547,
         n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555,
         n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563,
         n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
         n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579,
         n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
         n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
         n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603,
         n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611,
         n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619,
         n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627,
         n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635,
         n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643,
         n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
         n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659,
         n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
         n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675,
         n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683,
         n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
         n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699,
         n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707,
         n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
         n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723,
         n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731,
         n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
         n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747,
         n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755,
         n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763,
         n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771,
         n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779,
         n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787,
         n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795,
         n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803,
         n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
         n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
         n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
         n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835,
         n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843,
         n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
         n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
         n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867,
         n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875,
         n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
         n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891,
         n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899,
         n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907,
         n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
         n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923,
         n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
         n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
         n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947,
         n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
         n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963,
         n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
         n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979,
         n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987,
         n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995,
         n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003,
         n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011,
         n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019,
         n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027,
         n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035,
         n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043,
         n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051,
         n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059,
         n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067,
         n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
         n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083,
         n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091,
         n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099,
         n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107,
         n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
         n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123,
         n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131,
         n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139,
         n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
         n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155,
         n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163,
         n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171,
         n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
         n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187,
         n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195,
         n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203,
         n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211,
         n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219,
         n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227,
         n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235,
         n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
         n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251,
         n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
         n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267,
         n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275,
         n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283,
         n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291,
         n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299,
         n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307,
         n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
         n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323,
         n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331,
         n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339,
         n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347,
         n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355,
         n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363,
         n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371,
         n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
         n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
         n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395,
         n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403,
         n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411,
         n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419,
         n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427,
         n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
         n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443,
         n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451,
         n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459,
         n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467,
         n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475,
         n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483,
         n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491,
         n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499,
         n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507,
         n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515,
         n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523,
         n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531,
         n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539,
         n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547,
         n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555,
         n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563,
         n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571,
         n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579,
         n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587,
         n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595,
         n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603,
         n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611,
         n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619,
         n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627,
         n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635,
         n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643,
         n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651,
         n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659,
         n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667,
         n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675,
         n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683,
         n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691,
         n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699,
         n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707,
         n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715,
         n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
         n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731,
         n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739,
         n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747,
         n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755,
         n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763,
         n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771,
         n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779,
         n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787,
         n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
         n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803,
         n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811,
         n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819,
         n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827,
         n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835,
         n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843,
         n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851,
         n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859,
         n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867,
         n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875,
         n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883,
         n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891,
         n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899,
         n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907,
         n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915,
         n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923,
         n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931,
         n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939,
         n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947,
         n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955,
         n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963,
         n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971,
         n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979,
         n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987,
         n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995,
         n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003,
         n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011,
         n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019,
         n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027,
         n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035,
         n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043,
         n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051,
         n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059,
         n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067,
         n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075,
         n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083,
         n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091,
         n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099,
         n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107,
         n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115,
         n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123,
         n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131,
         n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139,
         n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147,
         n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155,
         n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163,
         n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171,
         n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179,
         n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187,
         n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195,
         n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203,
         n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211,
         n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219,
         n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227,
         n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235,
         n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243,
         n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251,
         n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259,
         n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267,
         n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275,
         n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283,
         n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291,
         n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299,
         n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307,
         n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315,
         n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323,
         n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331,
         n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339,
         n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347,
         n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355,
         n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363,
         n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371,
         n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379,
         n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387,
         n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395,
         n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403,
         n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411,
         n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419,
         n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427,
         n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435,
         n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443,
         n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451,
         n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459,
         n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467,
         n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475,
         n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483,
         n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491,
         n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499,
         n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507,
         n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515,
         n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523,
         n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531,
         n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539,
         n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547,
         n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555,
         n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563,
         n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571,
         n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579,
         n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587,
         n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595,
         n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603,
         n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611,
         n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619,
         n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627,
         n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635,
         n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643,
         n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651,
         n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659,
         n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667,
         n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675,
         n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683,
         n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691,
         n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699,
         n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707,
         n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715,
         n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723,
         n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731,
         n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739,
         n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747,
         n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755,
         n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763,
         n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771,
         n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779,
         n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787,
         n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795,
         n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803,
         n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811,
         n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819,
         n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827,
         n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835,
         n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843,
         n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851,
         n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859,
         n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867,
         n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875,
         n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883,
         n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891,
         n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899,
         n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907,
         n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915,
         n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923,
         n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931,
         n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939,
         n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947,
         n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955,
         n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963,
         n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971,
         n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979,
         n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987,
         n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995,
         n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003,
         n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011,
         n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019,
         n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027,
         n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035,
         n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043,
         n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051,
         n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059,
         n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067,
         n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075,
         n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083,
         n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091,
         n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099,
         n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107,
         n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115,
         n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123,
         n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131,
         n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139,
         n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147,
         n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155,
         n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163,
         n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171,
         n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179,
         n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187,
         n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195,
         n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203,
         n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211,
         n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219,
         n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227,
         n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235,
         n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243,
         n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251,
         n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259,
         n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267,
         n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275,
         n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283,
         n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291,
         n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299,
         n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307,
         n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315,
         n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323,
         n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331,
         n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339,
         n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347,
         n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355,
         n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363,
         n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371,
         n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379,
         n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387,
         n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395,
         n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403,
         n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411,
         n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419,
         n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427,
         n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435,
         n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443,
         n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451,
         n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459,
         n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467,
         n21468, n21469, n21470;

  NOR2_X1 U11246 ( .A1(n17817), .A2(n18099), .ZN(n18140) );
  AOI21_X1 U11247 ( .B1(n10094), .B2(n10722), .A(n9924), .ZN(n10093) );
  INV_X1 U11248 ( .A(n18993), .ZN(n18339) );
  AND2_X1 U11249 ( .A1(n10617), .A2(n10610), .ZN(n10716) );
  AND2_X1 U11250 ( .A1(n10617), .A2(n10616), .ZN(n19863) );
  INV_X2 U11251 ( .A(n17312), .ZN(n17292) );
  BUF_X1 U11252 ( .A(n11265), .Z(n11416) );
  INV_X1 U11253 ( .A(n17170), .ZN(n17304) );
  AND2_X1 U11254 ( .A1(n15638), .A2(n9820), .ZN(n15661) );
  CLKBUF_X2 U11255 ( .A(n11522), .Z(n17284) );
  NAND2_X1 U11256 ( .A1(n10639), .A2(n10999), .ZN(n13178) );
  OR2_X1 U11257 ( .A1(n10541), .A2(n10536), .ZN(n10589) );
  NOR2_X1 U11258 ( .A1(n11433), .A2(n11432), .ZN(n11487) );
  OR2_X1 U11259 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n17021) );
  AND2_X1 U11260 ( .A1(n13773), .A2(n11929), .ZN(n11886) );
  BUF_X1 U11261 ( .A(n11967), .Z(n12847) );
  CLKBUF_X2 U11262 ( .A(n11798), .Z(n12806) );
  CLKBUF_X2 U11263 ( .A(n11868), .Z(n12830) );
  INV_X1 U11264 ( .A(n12823), .ZN(n12849) );
  CLKBUF_X2 U11265 ( .A(n9852), .Z(n9821) );
  AND4_X1 U11266 ( .A1(n11784), .A2(n11783), .A3(n11782), .A4(n11781), .ZN(
        n11796) );
  AND2_X2 U11267 ( .A1(n11758), .A2(n11769), .ZN(n12860) );
  AND2_X1 U11268 ( .A1(n11759), .A2(n13941), .ZN(n11798) );
  AND2_X1 U11269 ( .A1(n13924), .A2(n11764), .ZN(n11966) );
  AND2_X1 U11270 ( .A1(n10639), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9808) );
  CLKBUF_X1 U11271 ( .A(n11747), .Z(n9802) );
  AOI21_X1 U11272 ( .B1(n15769), .B2(n11714), .A(n18828), .ZN(n11747) );
  INV_X1 U11273 ( .A(n9848), .ZN(n9803) );
  INV_X2 U11274 ( .A(n9803), .ZN(n9804) );
  OR2_X1 U11275 ( .A1(n10541), .A2(n11225), .ZN(n10512) );
  INV_X1 U11277 ( .A(n10410), .ZN(n9815) );
  OR2_X1 U11278 ( .A1(n10095), .A2(n10093), .ZN(n10092) );
  AND2_X2 U11279 ( .A1(n11757), .A2(n13925), .ZN(n11972) );
  OR2_X1 U11280 ( .A1(n14608), .A2(n14714), .ZN(n14571) );
  AND2_X2 U11281 ( .A1(n10421), .A2(n10444), .ZN(n10665) );
  AND2_X1 U11282 ( .A1(n9833), .A2(n10596), .ZN(n10620) );
  INV_X1 U11283 ( .A(n11939), .ZN(n12983) );
  AND3_X1 U11284 ( .A1(n11848), .A2(n10386), .A3(n11849), .ZN(n13763) );
  AND2_X1 U11285 ( .A1(n10617), .A2(n10611), .ZN(n10708) );
  INV_X2 U11286 ( .A(n11479), .ZN(n17269) );
  INV_X1 U11287 ( .A(n11638), .ZN(n9811) );
  INV_X2 U11288 ( .A(n17237), .ZN(n11444) );
  INV_X2 U11289 ( .A(n11467), .ZN(n17268) );
  INV_X1 U11290 ( .A(n20254), .ZN(n20289) );
  AND2_X2 U11291 ( .A1(n11882), .A2(n11881), .ZN(n11918) );
  AND2_X1 U11292 ( .A1(n15507), .A2(n15508), .ZN(n14902) );
  INV_X1 U11293 ( .A(n11225), .ZN(n10536) );
  INV_X1 U11294 ( .A(n11225), .ZN(n10527) );
  INV_X2 U11295 ( .A(n11219), .ZN(n19470) );
  NOR2_X1 U11297 ( .A1(n11555), .A2(n17809), .ZN(n18135) );
  NAND2_X1 U11298 ( .A1(n17920), .A2(n11548), .ZN(n11551) );
  NOR2_X1 U11299 ( .A1(n17490), .A2(n11518), .ZN(n11546) );
  AND2_X1 U11300 ( .A1(n12780), .A2(n12779), .ZN(n13751) );
  CLKBUF_X3 U11301 ( .A(n10491), .Z(n11217) );
  NAND2_X2 U11302 ( .A1(n19437), .A2(n11225), .ZN(n14159) );
  OR2_X1 U11303 ( .A1(n15570), .A2(n15546), .ZN(n15556) );
  NOR2_X1 U11304 ( .A1(n19764), .A2(n19668), .ZN(n19544) );
  NAND3_X1 U11305 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(P3_EBX_REG_17__SCAN_IN), 
        .A3(n17185), .ZN(n17167) );
  INV_X1 U11306 ( .A(n9890), .ZN(n17245) );
  NOR2_X1 U11307 ( .A1(n17626), .A2(n17627), .ZN(n16526) );
  INV_X1 U11308 ( .A(n17841), .ZN(n17827) );
  NAND2_X1 U11309 ( .A1(n18190), .A2(n18202), .ZN(n18268) );
  NAND2_X1 U11310 ( .A1(n17900), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17899) );
  NAND2_X1 U11311 ( .A1(n15767), .A2(n16648), .ZN(n18791) );
  OR2_X1 U11312 ( .A1(n11559), .A2(n10249), .ZN(n9805) );
  INV_X2 U11313 ( .A(n9888), .ZN(n17291) );
  INV_X1 U11314 ( .A(n17797), .ZN(n17886) );
  AND2_X1 U11315 ( .A1(n11770), .A2(n13910), .ZN(n9806) );
  AND2_X2 U11316 ( .A1(n11770), .A2(n13910), .ZN(n11807) );
  AND2_X1 U11317 ( .A1(n10639), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9807) );
  AND2_X1 U11319 ( .A1(n11759), .A2(n11758), .ZN(n12517) );
  AND2_X1 U11320 ( .A1(n11758), .A2(n13925), .ZN(n11868) );
  AND2_X4 U11321 ( .A1(n11947), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11758) );
  AND2_X1 U11322 ( .A1(n11770), .A2(n11757), .ZN(n11973) );
  NOR2_X2 U11323 ( .A1(n17686), .A2(n17685), .ZN(n17663) );
  NOR2_X4 U11324 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13925) );
  NAND2_X2 U11326 ( .A1(n12700), .A2(n10297), .ZN(n14683) );
  NOR2_X2 U11327 ( .A1(n10907), .A2(n10906), .ZN(n10890) );
  AND2_X1 U11328 ( .A1(n11770), .A2(n11757), .ZN(n9810) );
  AND4_X2 U11329 ( .A1(n11780), .A2(n11779), .A3(n11778), .A4(n11777), .ZN(
        n11797) );
  OR2_X1 U11330 ( .A1(n10050), .A2(n12680), .ZN(n10049) );
  NAND2_X2 U11331 ( .A1(n15650), .A2(n16432), .ZN(n13379) );
  NOR2_X1 U11332 ( .A1(n11433), .A2(n11432), .ZN(n9812) );
  INV_X1 U11333 ( .A(n11487), .ZN(n17170) );
  NOR2_X1 U11334 ( .A1(n18807), .A2(n11434), .ZN(n9813) );
  OAI22_X2 U11335 ( .A1(n14103), .A2(n14102), .B1(n15622), .B2(n19205), .ZN(
        n15311) );
  NAND2_X2 U11336 ( .A1(n15650), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10436) );
  INV_X1 U11337 ( .A(n10410), .ZN(n9814) );
  INV_X1 U11338 ( .A(n10410), .ZN(n16444) );
  NAND2_X2 U11339 ( .A1(n15659), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10410) );
  INV_X1 U11340 ( .A(n13249), .ZN(n9816) );
  INV_X1 U11341 ( .A(n13249), .ZN(n9817) );
  INV_X1 U11342 ( .A(n13249), .ZN(n10634) );
  NAND2_X2 U11343 ( .A1(n15659), .A2(n16432), .ZN(n13249) );
  NAND2_X1 U11344 ( .A1(n17651), .A2(n18015), .ZN(n17650) );
  INV_X4 U11345 ( .A(n16018), .ZN(n14680) );
  AND4_X1 U11346 ( .A1(n10712), .A2(n10711), .A3(n10710), .A4(n10709), .ZN(
        n10722) );
  AND2_X1 U11348 ( .A1(n16401), .A2(n9947), .ZN(n15584) );
  NAND2_X1 U11349 ( .A1(n20306), .A2(n20443), .ZN(n15974) );
  NAND2_X1 U11350 ( .A1(n18783), .A2(n18991), .ZN(n16632) );
  XNOR2_X1 U11351 ( .A(n11551), .B(n11550), .ZN(n17900) );
  NAND2_X1 U11352 ( .A1(n10573), .A2(n10572), .ZN(n10593) );
  NOR2_X1 U11354 ( .A1(n10864), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10871) );
  CLKBUF_X1 U11355 ( .A(n10557), .Z(n11092) );
  NAND2_X1 U11356 ( .A1(n16629), .A2(n19007), .ZN(n16646) );
  NAND2_X1 U11357 ( .A1(n10495), .A2(n10443), .ZN(n10525) );
  BUF_X2 U11358 ( .A(n11264), .Z(n11409) );
  NOR4_X1 U11359 ( .A1(n11669), .A2(n11663), .A3(n11660), .A4(n11661), .ZN(
        n11674) );
  CLKBUF_X1 U11360 ( .A(n10531), .Z(n19464) );
  NOR2_X1 U11361 ( .A1(n11701), .A2(n18355), .ZN(n11703) );
  NOR2_X1 U11362 ( .A1(n18355), .A2(n11671), .ZN(n18796) );
  NAND2_X1 U11363 ( .A1(n12983), .A2(n13630), .ZN(n13779) );
  CLKBUF_X2 U11364 ( .A(n11939), .Z(n12975) );
  NAND2_X1 U11365 ( .A1(n10757), .A2(n10520), .ZN(n10357) );
  CLKBUF_X2 U11366 ( .A(n10757), .Z(n11219) );
  NAND2_X1 U11367 ( .A1(n17370), .A2(n11671), .ZN(n11661) );
  INV_X2 U11369 ( .A(n12074), .ZN(n11928) );
  NOR2_X1 U11370 ( .A1(n11225), .A2(n19437), .ZN(n10499) );
  INV_X1 U11371 ( .A(n13767), .ZN(n13773) );
  INV_X16 U11372 ( .A(n10858), .ZN(n14246) );
  OR3_X1 U11373 ( .A1(n11583), .A2(n11584), .A3(n10016), .ZN(n17516) );
  INV_X1 U11374 ( .A(n20413), .ZN(n9818) );
  NAND2_X1 U11375 ( .A1(n10456), .A2(n10455), .ZN(n10520) );
  BUF_X2 U11376 ( .A(n11909), .Z(n9849) );
  CLKBUF_X2 U11377 ( .A(n10649), .Z(n13217) );
  INV_X1 U11378 ( .A(n11785), .ZN(n9852) );
  CLKBUF_X2 U11379 ( .A(n11807), .Z(n12862) );
  CLKBUF_X2 U11380 ( .A(n11522), .Z(n17273) );
  INV_X2 U11381 ( .A(n13312), .ZN(n13242) );
  INV_X2 U11383 ( .A(n12502), .ZN(n11967) );
  NAND2_X2 U11384 ( .A1(n13941), .A2(n11769), .ZN(n12441) );
  NAND2_X2 U11385 ( .A1(n13925), .A2(n13941), .ZN(n12502) );
  AND2_X4 U11386 ( .A1(n10392), .A2(n15651), .ZN(n13312) );
  INV_X2 U11387 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10256) );
  OAI21_X1 U11388 ( .B1(n15110), .B2(n15111), .A(n14242), .ZN(n14249) );
  XNOR2_X1 U11389 ( .A(n10192), .B(n9930), .ZN(n15435) );
  AND2_X1 U11390 ( .A1(n10280), .A2(n10283), .ZN(n14955) );
  AOI21_X1 U11391 ( .B1(n16260), .B2(n16406), .A(n9907), .ZN(n14273) );
  OR2_X1 U11392 ( .A1(n13336), .A2(n13335), .ZN(n13337) );
  NAND2_X1 U11393 ( .A1(n14977), .A2(n10377), .ZN(n13336) );
  NOR2_X1 U11394 ( .A1(n12788), .A2(n10052), .ZN(n10051) );
  AOI21_X1 U11395 ( .B1(n15498), .B2(n15216), .A(n15215), .ZN(n15260) );
  NAND2_X1 U11396 ( .A1(n14976), .A2(n14978), .ZN(n14977) );
  NAND2_X1 U11397 ( .A1(n9915), .A2(n10112), .ZN(n14555) );
  OR2_X1 U11398 ( .A1(n13309), .A2(n13308), .ZN(n10377) );
  NAND2_X1 U11399 ( .A1(n11081), .A2(n11080), .ZN(n15161) );
  NOR2_X1 U11400 ( .A1(n12721), .A2(n14714), .ZN(n14539) );
  NAND2_X1 U11401 ( .A1(n9892), .A2(n10336), .ZN(n13051) );
  NAND2_X1 U11402 ( .A1(n14985), .A2(n13289), .ZN(n13307) );
  OR2_X1 U11403 ( .A1(n13288), .A2(n13287), .ZN(n13289) );
  AOI21_X1 U11404 ( .B1(n9903), .B2(n17882), .A(n16503), .ZN(n16504) );
  NAND2_X1 U11405 ( .A1(n10273), .A2(n10272), .ZN(n10275) );
  NAND2_X1 U11406 ( .A1(n15606), .A2(n11073), .ZN(n16354) );
  AND2_X1 U11407 ( .A1(n10363), .A2(n10360), .ZN(n9831) );
  AND2_X1 U11408 ( .A1(n13240), .A2(n13264), .ZN(n13241) );
  OAI211_X1 U11409 ( .C1(n11070), .C2(n11071), .A(n11069), .B(n11068), .ZN(
        n15607) );
  NAND2_X1 U11410 ( .A1(n16346), .A2(n10862), .ZN(n10363) );
  NAND2_X1 U11411 ( .A1(n14180), .A2(n12698), .ZN(n12700) );
  NAND2_X1 U11412 ( .A1(n17650), .A2(n10242), .ZN(n11563) );
  OR2_X1 U11413 ( .A1(n15040), .A2(n15039), .ZN(n16211) );
  AND2_X1 U11414 ( .A1(n17670), .A2(n9940), .ZN(n10242) );
  NAND2_X1 U11415 ( .A1(n10021), .A2(n12673), .ZN(n14048) );
  NAND2_X1 U11416 ( .A1(n10093), .A2(n10095), .ZN(n10847) );
  NAND2_X1 U11417 ( .A1(n19283), .A2(n13107), .ZN(n13974) );
  OR2_X1 U11418 ( .A1(n15998), .A2(n12713), .ZN(n14656) );
  NAND2_X1 U11419 ( .A1(n10844), .A2(n10843), .ZN(n11066) );
  AND2_X1 U11420 ( .A1(n9911), .A2(n12699), .ZN(n10297) );
  AND2_X1 U11421 ( .A1(n19209), .A2(n19210), .ZN(n19283) );
  AND2_X1 U11422 ( .A1(n15988), .A2(n14664), .ZN(n12712) );
  NOR2_X1 U11423 ( .A1(n10058), .A2(n10054), .ZN(n10094) );
  OR2_X1 U11424 ( .A1(n10829), .A2(n10828), .ZN(n10844) );
  OAI211_X1 U11425 ( .C1(n16502), .C2(n17993), .A(n16501), .B(n16500), .ZN(
        n16503) );
  NAND2_X1 U11426 ( .A1(n10687), .A2(n9891), .ZN(n10791) );
  NAND2_X1 U11427 ( .A1(n10719), .A2(n10055), .ZN(n10054) );
  AND4_X1 U11428 ( .A1(n10686), .A2(n10685), .A3(n10684), .A4(n10683), .ZN(
        n10687) );
  AOI211_X1 U11429 ( .C1(n10707), .C2(n20136), .A(n19692), .B(n20126), .ZN(
        n19672) );
  NOR2_X1 U11430 ( .A1(n10912), .A2(n10369), .ZN(n10368) );
  NOR2_X1 U11431 ( .A1(n10717), .A2(n10718), .ZN(n10056) );
  NOR2_X1 U11432 ( .A1(n19926), .A2(n19953), .ZN(n10057) );
  OAI21_X1 U11433 ( .B1(n10678), .B2(n13127), .A(n19447), .ZN(n10628) );
  BUF_X1 U11434 ( .A(n10714), .Z(n19798) );
  BUF_X1 U11435 ( .A(n10715), .Z(n19702) );
  NOR2_X1 U11436 ( .A1(n17708), .A2(n17681), .ZN(n11558) );
  OR2_X1 U11437 ( .A1(n10627), .A2(n10606), .ZN(n10678) );
  AOI22_X1 U11438 ( .A1(n18184), .A2(n17917), .B1(n17895), .B2(n18186), .ZN(
        n17885) );
  AND2_X1 U11439 ( .A1(n13592), .A2(n19245), .ZN(n10616) );
  AND2_X1 U11440 ( .A1(n19227), .A2(n19245), .ZN(n10626) );
  CLKBUF_X2 U11441 ( .A(n13081), .Z(n14942) );
  CLKBUF_X1 U11442 ( .A(n14456), .Z(n14508) );
  CLKBUF_X1 U11443 ( .A(n13062), .Z(n14506) );
  NAND2_X1 U11444 ( .A1(n13091), .A2(n13090), .ZN(n13095) );
  NAND2_X1 U11445 ( .A1(n10607), .A2(n10601), .ZN(n19227) );
  NOR2_X1 U11446 ( .A1(n20542), .A2(n20398), .ZN(n20939) );
  INV_X1 U11447 ( .A(n17917), .ZN(n17993) );
  NOR2_X1 U11448 ( .A1(n20542), .A2(n20407), .ZN(n20945) );
  INV_X1 U11449 ( .A(n17988), .ZN(n17975) );
  NOR2_X1 U11450 ( .A1(n20542), .A2(n20415), .ZN(n20951) );
  NAND2_X1 U11451 ( .A1(n10140), .A2(n12107), .ZN(n12108) );
  NOR2_X1 U11452 ( .A1(n20542), .A2(n20422), .ZN(n20957) );
  NOR2_X1 U11453 ( .A1(n20542), .A2(n20429), .ZN(n20963) );
  NOR2_X1 U11454 ( .A1(n20542), .A2(n20436), .ZN(n20971) );
  NOR2_X1 U11455 ( .A1(n20542), .A2(n20447), .ZN(n20978) );
  NOR2_X1 U11456 ( .A1(n20542), .A2(n20387), .ZN(n20923) );
  INV_X1 U11457 ( .A(n13089), .ZN(n19245) );
  NAND2_X2 U11458 ( .A1(n14527), .A2(n13806), .ZN(n14536) );
  NAND2_X1 U11459 ( .A1(n15623), .A2(n11259), .ZN(n15613) );
  NAND2_X1 U11460 ( .A1(n10091), .A2(n10598), .ZN(n10597) );
  AND2_X1 U11461 ( .A1(n10608), .A2(n10605), .ZN(n13089) );
  NAND3_X1 U11462 ( .A1(n18993), .A2(n18783), .A3(n18991), .ZN(n17992) );
  OR2_X1 U11463 ( .A1(n16776), .A2(n16991), .ZN(n10077) );
  CLKBUF_X1 U11464 ( .A(n10599), .Z(n10600) );
  NAND2_X1 U11465 ( .A1(n10046), .A2(n10045), .ZN(n20479) );
  NAND2_X1 U11466 ( .A1(n11216), .A2(n11045), .ZN(n16425) );
  NAND2_X1 U11467 ( .A1(n12090), .A2(n12089), .ZN(n20537) );
  INV_X2 U11468 ( .A(n19293), .ZN(n14945) );
  NOR2_X1 U11469 ( .A1(n16784), .A2(n16949), .ZN(n16777) );
  NAND2_X1 U11470 ( .A1(n10587), .A2(n10586), .ZN(n11117) );
  NAND2_X1 U11471 ( .A1(n10883), .A2(n10952), .ZN(n10882) );
  NOR2_X1 U11472 ( .A1(n13728), .A2(n11244), .ZN(n14084) );
  NOR2_X1 U11473 ( .A1(n17328), .A2(n10262), .ZN(n17306) );
  OAI21_X1 U11474 ( .B1(n12075), .B2(n10299), .A(n9904), .ZN(n12029) );
  NOR2_X1 U11475 ( .A1(n13520), .A2(n19435), .ZN(n19481) );
  AND2_X1 U11476 ( .A1(n10296), .A2(n10295), .ZN(n10545) );
  NAND2_X1 U11477 ( .A1(n10263), .A2(P3_EBX_REG_6__SCAN_IN), .ZN(n17328) );
  AND3_X1 U11478 ( .A1(n10592), .A2(n10591), .A3(n10590), .ZN(n11116) );
  OAI211_X1 U11479 ( .C1(n14253), .C2(n10580), .A(n10579), .B(n10578), .ZN(
        n10582) );
  AND2_X1 U11480 ( .A1(n10871), .A2(n19281), .ZN(n10872) );
  XOR2_X1 U11481 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n16506), .Z(
        n16949) );
  NAND2_X1 U11482 ( .A1(n17943), .A2(n11541), .ZN(n11544) );
  AND3_X1 U11483 ( .A1(n10513), .A2(n10514), .A3(n10515), .ZN(n10544) );
  INV_X1 U11484 ( .A(n10313), .ZN(n11243) );
  AOI21_X1 U11485 ( .B1(n11653), .B2(n11652), .A(n11651), .ZN(n15767) );
  OR2_X1 U11487 ( .A1(n10867), .A2(n10856), .ZN(n10864) );
  AND2_X1 U11488 ( .A1(n10557), .A2(n10561), .ZN(n10539) );
  OAI21_X1 U11489 ( .B1(n11113), .B2(n10576), .A(n10575), .ZN(n10577) );
  OAI211_X1 U11490 ( .C1(n10564), .C2(n13558), .A(n16478), .B(n10563), .ZN(
        n10565) );
  INV_X2 U11492 ( .A(n10589), .ZN(n14255) );
  NAND3_X2 U11493 ( .A1(n18339), .A2(n17554), .A3(n17553), .ZN(n17619) );
  NOR2_X1 U11494 ( .A1(n11935), .A2(n11922), .ZN(n12882) );
  AND2_X2 U11495 ( .A1(n13604), .A2(n20380), .ZN(n12881) );
  OAI22_X1 U11496 ( .A1(n18782), .A2(n15770), .B1(n14219), .B2(n14218), .ZN(
        n15868) );
  AND2_X1 U11497 ( .A1(n13680), .A2(n13679), .ZN(n11235) );
  NAND2_X1 U11498 ( .A1(n11685), .A2(n18775), .ZN(n16629) );
  NOR2_X1 U11499 ( .A1(n10552), .A2(n10551), .ZN(n15638) );
  XNOR2_X1 U11500 ( .A(n11722), .B(n10088), .ZN(n11540) );
  NOR2_X1 U11501 ( .A1(n10803), .A2(n10802), .ZN(n10801) );
  NOR2_X1 U11502 ( .A1(n10224), .A2(n10788), .ZN(n10223) );
  INV_X1 U11503 ( .A(n12772), .ZN(n12764) );
  OR2_X1 U11504 ( .A1(n13638), .A2(n13760), .ZN(n13775) );
  INV_X1 U11505 ( .A(n10813), .ZN(n10224) );
  OR2_X1 U11506 ( .A1(n11884), .A2(n11941), .ZN(n13612) );
  AND2_X1 U11507 ( .A1(n11982), .A2(n20380), .ZN(n12772) );
  AND2_X1 U11508 ( .A1(n11217), .A2(n11022), .ZN(n10550) );
  NOR2_X1 U11509 ( .A1(n10493), .A2(n11022), .ZN(n10517) );
  NOR2_X1 U11510 ( .A1(n17498), .A2(n11537), .ZN(n11538) );
  AND2_X1 U11511 ( .A1(n10531), .A2(n10491), .ZN(n10495) );
  NOR2_X1 U11512 ( .A1(n17987), .A2(n18300), .ZN(n17986) );
  AND2_X2 U11513 ( .A1(n11220), .A2(n11219), .ZN(n11374) );
  CLKBUF_X1 U11514 ( .A(n12898), .Z(n13686) );
  OR2_X1 U11515 ( .A1(n17503), .A2(n11716), .ZN(n11537) );
  XNOR2_X1 U11516 ( .A(n11535), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n17968) );
  INV_X1 U11517 ( .A(n21069), .ZN(n12695) );
  NAND2_X1 U11518 ( .A1(n13075), .A2(n11218), .ZN(n11031) );
  OR2_X1 U11519 ( .A1(n12019), .A2(n12018), .ZN(n12641) );
  NAND2_X1 U11520 ( .A1(n17409), .A2(n18336), .ZN(n11660) );
  AND2_X1 U11521 ( .A1(n11918), .A2(n13753), .ZN(n14026) );
  AND2_X1 U11522 ( .A1(n10757), .A2(n13070), .ZN(n11030) );
  NAND2_X1 U11523 ( .A1(n13763), .A2(n9818), .ZN(n13923) );
  INV_X1 U11524 ( .A(n11916), .ZN(n10115) );
  INV_X1 U11525 ( .A(n10972), .ZN(n14846) );
  NAND3_X1 U11526 ( .A1(n17746), .A2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17737) );
  INV_X1 U11528 ( .A(n10530), .ZN(n19458) );
  XOR2_X1 U11529 ( .A(n17516), .B(n18993), .Z(n19007) );
  NAND2_X1 U11530 ( .A1(n12092), .A2(n12091), .ZN(n12741) );
  INV_X1 U11531 ( .A(n17370), .ZN(n18355) );
  AND2_X1 U11532 ( .A1(n10530), .A2(n11018), .ZN(n10496) );
  CLKBUF_X1 U11533 ( .A(n13075), .Z(n13076) );
  INV_X1 U11534 ( .A(n14159), .ZN(n20169) );
  OAI211_X1 U11535 ( .C1(n9890), .C2(n17124), .A(n11606), .B(n11605), .ZN(
        n17370) );
  NAND2_X1 U11536 ( .A1(n19437), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10972) );
  OR2_X1 U11537 ( .A1(n11917), .A2(n11918), .ZN(n21069) );
  INV_X1 U11538 ( .A(n10520), .ZN(n13070) );
  NOR2_X1 U11539 ( .A1(n17770), .A2(n17769), .ZN(n17746) );
  INV_X1 U11540 ( .A(n17516), .ZN(n18336) );
  OR2_X1 U11541 ( .A1(n12004), .A2(n12003), .ZN(n12694) );
  NAND3_X1 U11542 ( .A1(n11494), .A2(n11495), .A3(n9916), .ZN(n11533) );
  INV_X2 U11543 ( .A(n11917), .ZN(n13753) );
  OAI211_X2 U11544 ( .C1(n17237), .C2(n17287), .A(n11595), .B(n11594), .ZN(
        n18993) );
  INV_X1 U11545 ( .A(n11218), .ZN(n10757) );
  OAI211_X1 U11546 ( .C1(n11638), .C2(n17354), .A(n11576), .B(n11575), .ZN(
        n11701) );
  BUF_X1 U11547 ( .A(n10520), .Z(n13075) );
  AND2_X1 U11548 ( .A1(n10492), .A2(n10502), .ZN(n10443) );
  NAND4_X1 U11549 ( .A1(n11833), .A2(n11832), .A3(n11831), .A4(n11830), .ZN(
        n11929) );
  OAI211_X1 U11550 ( .C1(n9890), .C2(n17110), .A(n11616), .B(n11615), .ZN(
        n11671) );
  INV_X1 U11551 ( .A(n11918), .ZN(n20380) );
  OAI211_X1 U11552 ( .C1(n11523), .C2(n17236), .A(n11627), .B(n11626), .ZN(
        n11663) );
  AOI211_X1 U11553 ( .C1(n17293), .C2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A(
        n11593), .B(n11592), .ZN(n11594) );
  MUX2_X1 U11554 ( .A(n10429), .B(n10428), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10492) );
  NOR2_X1 U11555 ( .A1(n11484), .A2(n11483), .ZN(n17503) );
  NAND2_X1 U11556 ( .A1(n10467), .A2(n10468), .ZN(n11218) );
  AND4_X1 U11557 ( .A1(n11821), .A2(n11820), .A3(n11819), .A4(n11818), .ZN(
        n11832) );
  AND2_X2 U11558 ( .A1(n11776), .A2(n11775), .ZN(n12074) );
  INV_X1 U11559 ( .A(n11910), .ZN(n11911) );
  OR2_X2 U11560 ( .A1(n16582), .A2(n16536), .ZN(n16584) );
  AND4_X1 U11561 ( .A1(n11864), .A2(n11863), .A3(n11862), .A4(n11861), .ZN(
        n11865) );
  AND4_X1 U11562 ( .A1(n11853), .A2(n11852), .A3(n11851), .A4(n11850), .ZN(
        n11866) );
  AND4_X1 U11563 ( .A1(n11802), .A2(n11801), .A3(n11800), .A4(n11799), .ZN(
        n11813) );
  AND4_X1 U11564 ( .A1(n11829), .A2(n11828), .A3(n11827), .A4(n11826), .ZN(
        n11830) );
  NOR2_X1 U11565 ( .A1(n11880), .A2(n11879), .ZN(n11881) );
  AND4_X1 U11566 ( .A1(n11872), .A2(n11871), .A3(n11870), .A4(n11869), .ZN(
        n11882) );
  AND4_X1 U11567 ( .A1(n11897), .A2(n11896), .A3(n11895), .A4(n11894), .ZN(
        n11914) );
  AND4_X1 U11568 ( .A1(n11825), .A2(n11824), .A3(n11823), .A4(n11822), .ZN(
        n11831) );
  AND4_X1 U11569 ( .A1(n11859), .A2(n11858), .A3(n11857), .A4(n11856), .ZN(
        n11863) );
  AND4_X1 U11570 ( .A1(n11789), .A2(n11788), .A3(n11787), .A4(n11786), .ZN(
        n11795) );
  NOR2_X1 U11571 ( .A1(n10435), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10440) );
  CLKBUF_X1 U11572 ( .A(n10694), .Z(n13141) );
  AND2_X1 U11573 ( .A1(n10423), .A2(n10422), .ZN(n10427) );
  NAND2_X1 U11574 ( .A1(n17889), .A2(n16667), .ZN(n17833) );
  NOR2_X1 U11575 ( .A1(n16925), .A2(n17903), .ZN(n17889) );
  INV_X1 U11576 ( .A(n11523), .ZN(n17313) );
  AND2_X2 U11577 ( .A1(n10483), .A2(n10444), .ZN(n13220) );
  INV_X1 U11578 ( .A(n17288), .ZN(n17219) );
  AND4_X1 U11579 ( .A1(n11901), .A2(n11900), .A3(n11899), .A4(n11898), .ZN(
        n11913) );
  AND4_X1 U11580 ( .A1(n11905), .A2(n11904), .A3(n11903), .A4(n11902), .ZN(
        n11912) );
  NAND2_X2 U11581 ( .A1(n18933), .A2(n18864), .ZN(n18926) );
  BUF_X2 U11582 ( .A(n11893), .Z(n9837) );
  INV_X1 U11583 ( .A(n13381), .ZN(n10632) );
  INV_X1 U11584 ( .A(n13381), .ZN(n13392) );
  CLKBUF_X1 U11585 ( .A(n12477), .Z(n12829) );
  NAND2_X2 U11586 ( .A1(n20178), .A2(n20055), .ZN(n20109) );
  NAND2_X2 U11587 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20178), .ZN(n20106) );
  INV_X1 U11588 ( .A(n9888), .ZN(n17154) );
  CLKBUF_X1 U11589 ( .A(n11893), .Z(n9836) );
  INV_X2 U11590 ( .A(n13381), .ZN(n9838) );
  NOR2_X1 U11591 ( .A1(n10195), .A2(n9905), .ZN(n10194) );
  OR2_X1 U11592 ( .A1(n17021), .A2(n11433), .ZN(n9890) );
  INV_X2 U11593 ( .A(n16621), .ZN(n16623) );
  NAND2_X1 U11594 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11429), .ZN(
        n17237) );
  NOR2_X2 U11595 ( .A1(n17931), .A2(n17930), .ZN(n17919) );
  INV_X4 U11596 ( .A(n9856), .ZN(n17309) );
  INV_X2 U11597 ( .A(n18312), .ZN(n9822) );
  NAND2_X2 U11598 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18789), .ZN(
        n17312) );
  INV_X1 U11599 ( .A(n11835), .ZN(n11892) );
  INV_X2 U11600 ( .A(n10469), .ZN(n9834) );
  INV_X2 U11601 ( .A(n10469), .ZN(n10482) );
  NAND2_X1 U11602 ( .A1(n10639), .A2(n16432), .ZN(n13381) );
  AND2_X4 U11603 ( .A1(n10639), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10421) );
  INV_X2 U11604 ( .A(n21081), .ZN(n21038) );
  AND2_X2 U11605 ( .A1(n13312), .A2(n10444), .ZN(n10728) );
  NAND2_X1 U11606 ( .A1(n17949), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17931) );
  NAND2_X1 U11607 ( .A1(n10391), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10469) );
  AND2_X1 U11608 ( .A1(n13644), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11757) );
  NAND4_X1 U11609 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18996), .A3(n19005), 
        .A4(n16655), .ZN(n18842) );
  OR2_X1 U11610 ( .A1(n10255), .A2(n17021), .ZN(n11638) );
  INV_X1 U11611 ( .A(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12608) );
  INV_X1 U11612 ( .A(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12516) );
  AND2_X1 U11613 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11769) );
  AND2_X2 U11614 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13910) );
  NAND2_X1 U11615 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18807) );
  CLKBUF_X1 U11616 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n15662) );
  NOR2_X1 U11617 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10391) );
  NOR2_X1 U11618 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10392) );
  INV_X1 U11619 ( .A(n13773), .ZN(n9823) );
  AND2_X2 U11620 ( .A1(n11813), .A2(n11812), .ZN(n13767) );
  NAND2_X2 U11621 ( .A1(n13040), .A2(n13043), .ZN(n13769) );
  AND2_X1 U11622 ( .A1(n12898), .A2(n11916), .ZN(n13628) );
  INV_X1 U11623 ( .A(n17834), .ZN(n17785) );
  AND2_X2 U11624 ( .A1(n9824), .A2(n10116), .ZN(n13604) );
  NOR2_X1 U11625 ( .A1(n11887), .A2(n11916), .ZN(n9824) );
  INV_X1 U11626 ( .A(n10502), .ZN(n11018) );
  NAND2_X1 U11627 ( .A1(n10059), .A2(n10502), .ZN(n11025) );
  NOR2_X2 U11628 ( .A1(n13974), .A2(n10286), .ZN(n14096) );
  NAND2_X1 U11629 ( .A1(n10116), .A2(n10115), .ZN(n12723) );
  NOR2_X1 U11630 ( .A1(n13628), .A2(n11938), .ZN(n11919) );
  NOR2_X2 U11631 ( .A1(n16700), .A2(n16991), .ZN(n16690) );
  NOR2_X2 U11632 ( .A1(n16747), .A2(n16991), .ZN(n16734) );
  CLKBUF_X1 U11633 ( .A(n12700), .Z(n9825) );
  OR2_X2 U11634 ( .A1(n11935), .A2(n9826), .ZN(n13043) );
  OR2_X1 U11635 ( .A1(n11922), .A2(n11917), .ZN(n9826) );
  NAND2_X1 U11636 ( .A1(n11887), .A2(n9818), .ZN(n9827) );
  NAND2_X1 U11637 ( .A1(n9827), .A2(n11888), .ZN(n11891) );
  NOR2_X2 U11638 ( .A1(n16743), .A2(n16652), .ZN(n16712) );
  NOR3_X2 U11639 ( .A1(n17088), .A2(n16704), .A3(n16718), .ZN(n10260) );
  AND2_X2 U11640 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17213), .ZN(n17185) );
  NAND2_X1 U11641 ( .A1(n10122), .A2(n12108), .ZN(n9828) );
  AND2_X1 U11642 ( .A1(n12074), .A2(n11926), .ZN(n9829) );
  NAND2_X1 U11643 ( .A1(n10122), .A2(n12108), .ZN(n12147) );
  AND2_X1 U11644 ( .A1(n12074), .A2(n11926), .ZN(n11885) );
  CLKBUF_X1 U11645 ( .A(n15187), .Z(n9830) );
  CLKBUF_X1 U11646 ( .A(n15310), .Z(n9832) );
  XNOR2_X1 U11648 ( .A(n10186), .B(n11119), .ZN(n13820) );
  NAND2_X2 U11649 ( .A1(n10125), .A2(n10584), .ZN(n10186) );
  AND2_X1 U11650 ( .A1(n11770), .A2(n13941), .ZN(n11893) );
  INV_X1 U11651 ( .A(n9834), .ZN(n9835) );
  AND2_X2 U11652 ( .A1(n10389), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10639) );
  OR2_X1 U11653 ( .A1(n10603), .A2(n10602), .ZN(n10608) );
  NAND2_X1 U11654 ( .A1(n10603), .A2(n10602), .ZN(n10598) );
  INV_X1 U11655 ( .A(n13392), .ZN(n9839) );
  INV_X2 U11656 ( .A(n10436), .ZN(n9840) );
  INV_X2 U11657 ( .A(n10436), .ZN(n10483) );
  INV_X1 U11658 ( .A(n11785), .ZN(n12854) );
  NAND2_X1 U11659 ( .A1(n10022), .A2(n12664), .ZN(n14016) );
  OR2_X2 U11660 ( .A1(n12689), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14135) );
  NOR2_X4 U11661 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13941) );
  INV_X2 U11662 ( .A(n13379), .ZN(n9841) );
  INV_X1 U11663 ( .A(n13379), .ZN(n9842) );
  NAND2_X2 U11664 ( .A1(n14450), .A2(n14449), .ZN(n14522) );
  NOR2_X2 U11665 ( .A1(n17737), .A2(n17736), .ZN(n17713) );
  NAND2_X2 U11666 ( .A1(n14622), .A2(n12719), .ZN(n10144) );
  OR2_X1 U11667 ( .A1(n14648), .A2(n16018), .ZN(n10043) );
  OR3_X2 U11668 ( .A1(n14648), .A2(n12718), .A3(n9989), .ZN(n10039) );
  NAND2_X1 U11669 ( .A1(n12166), .A2(n12165), .ZN(n12199) );
  OAI21_X1 U11670 ( .B1(n13953), .B2(n12172), .A(n12118), .ZN(n13973) );
  AND2_X1 U11671 ( .A1(n11758), .A2(n11769), .ZN(n9843) );
  AND2_X1 U11672 ( .A1(n11758), .A2(n11769), .ZN(n9844) );
  INV_X1 U11673 ( .A(n9843), .ZN(n9845) );
  NAND2_X1 U11674 ( .A1(n10141), .A2(n10143), .ZN(n20565) );
  INV_X1 U11675 ( .A(n10143), .ZN(n10120) );
  NOR2_X1 U11676 ( .A1(n11811), .A2(n11810), .ZN(n11812) );
  INV_X1 U11677 ( .A(n13141), .ZN(n9846) );
  NOR2_X2 U11678 ( .A1(n14039), .A2(n14068), .ZN(n14069) );
  NAND2_X2 U11679 ( .A1(n12147), .A2(n12110), .ZN(n13953) );
  XOR2_X1 U11680 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n16506), .Z(n9847) );
  AND2_X4 U11681 ( .A1(n14384), .A2(n14386), .ZN(n14359) );
  NOR2_X4 U11682 ( .A1(n14429), .A2(n14487), .ZN(n14384) );
  NAND2_X2 U11683 ( .A1(n11886), .A2(n9829), .ZN(n11888) );
  AND2_X1 U11684 ( .A1(n11770), .A2(n11757), .ZN(n9848) );
  NOR2_X2 U11685 ( .A1(n13972), .A2(n13999), .ZN(n13997) );
  NAND2_X1 U11686 ( .A1(n13921), .A2(n13928), .ZN(n11909) );
  NAND2_X2 U11687 ( .A1(n12627), .A2(n12629), .ZN(n12817) );
  AOI21_X4 U11688 ( .B1(n13024), .B2(n14290), .A(n13023), .ZN(n14563) );
  OR2_X2 U11689 ( .A1(n12817), .A2(n10341), .ZN(n14290) );
  NAND2_X1 U11690 ( .A1(n13921), .A2(n13928), .ZN(n9850) );
  NAND2_X1 U11691 ( .A1(n13921), .A2(n13928), .ZN(n9851) );
  NAND2_X1 U11692 ( .A1(n11758), .A2(n11770), .ZN(n11785) );
  XNOR2_X2 U11693 ( .A(n12085), .B(n12084), .ZN(n12640) );
  NAND2_X1 U11694 ( .A1(n11538), .A2(n11722), .ZN(n11518) );
  NAND2_X1 U11695 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n10256), .ZN(
        n11433) );
  INV_X1 U11696 ( .A(n11471), .ZN(n11523) );
  NAND2_X1 U11697 ( .A1(n17773), .A2(n17886), .ZN(n10248) );
  AOI21_X1 U11698 ( .B1(n10508), .B2(n10507), .A(n19458), .ZN(n10509) );
  CLKBUF_X1 U11699 ( .A(n11961), .Z(n12291) );
  NAND2_X1 U11700 ( .A1(n12164), .A2(n12163), .ZN(n12165) );
  NAND2_X1 U11701 ( .A1(n10043), .A2(n10041), .ZN(n12719) );
  AND2_X1 U11702 ( .A1(n10042), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10041) );
  OR2_X1 U11703 ( .A1(n9860), .A2(n16018), .ZN(n10042) );
  NAND2_X1 U11704 ( .A1(n9886), .A2(n10952), .ZN(n10957) );
  NOR2_X1 U11705 ( .A1(n11225), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11220) );
  NOR2_X1 U11706 ( .A1(n11018), .A2(n10527), .ZN(n10528) );
  AOI21_X1 U11707 ( .B1(n11006), .B2(n10975), .A(n10761), .ZN(n10781) );
  INV_X1 U11708 ( .A(n17495), .ZN(n11722) );
  NOR2_X1 U11709 ( .A1(n15856), .A2(n14425), .ZN(n10149) );
  NOR2_X1 U11710 ( .A1(n12970), .A2(n10160), .ZN(n10159) );
  INV_X1 U11711 ( .A(n14349), .ZN(n10160) );
  NAND2_X1 U11712 ( .A1(n14594), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12721) );
  AND2_X1 U11713 ( .A1(n13485), .A2(n12975), .ZN(n12974) );
  AND2_X1 U11714 ( .A1(n15916), .A2(n14444), .ZN(n10151) );
  INV_X1 U11715 ( .A(n11888), .ZN(n13750) );
  NAND2_X1 U11716 ( .A1(n13767), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12092) );
  NAND2_X1 U11717 ( .A1(n12029), .A2(n12691), .ZN(n12052) );
  NAND2_X1 U11718 ( .A1(n12072), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10298) );
  NAND2_X1 U11719 ( .A1(n11918), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12091) );
  AND2_X1 U11720 ( .A1(n12733), .A2(n12732), .ZN(n12887) );
  NOR2_X1 U11721 ( .A1(n10228), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10227) );
  INV_X1 U11722 ( .A(n10229), .ZN(n10228) );
  NAND2_X1 U11723 ( .A1(n10932), .A2(n10952), .ZN(n10929) );
  AND2_X1 U11724 ( .A1(n19470), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10906) );
  OR2_X1 U11725 ( .A1(n10867), .A2(n19470), .ZN(n10952) );
  INV_X1 U11726 ( .A(n13874), .ZN(n11131) );
  INV_X1 U11727 ( .A(n16266), .ZN(n10292) );
  NAND2_X1 U11728 ( .A1(n10203), .A2(n15235), .ZN(n10202) );
  INV_X1 U11729 ( .A(n10204), .ZN(n10203) );
  INV_X1 U11730 ( .A(n14006), .ZN(n10210) );
  AND4_X1 U11731 ( .A1(n10752), .A2(n10751), .A3(n10750), .A4(n10749), .ZN(
        n10753) );
  AND3_X1 U11732 ( .A1(n10745), .A2(n10744), .A3(n10743), .ZN(n10754) );
  AND4_X1 U11733 ( .A1(n10742), .A2(n10741), .A3(n10740), .A4(n10739), .ZN(
        n10755) );
  AND2_X1 U11734 ( .A1(n13406), .A2(n11220), .ZN(n11264) );
  OR2_X1 U11735 ( .A1(n20167), .A2(n11046), .ZN(n11012) );
  AND2_X1 U11736 ( .A1(n16491), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13537) );
  AND2_X1 U11737 ( .A1(n15641), .A2(n19447), .ZN(n13665) );
  NAND2_X1 U11738 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n11435), .ZN(
        n11434) );
  NAND2_X1 U11739 ( .A1(n18972), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11432) );
  INV_X1 U11740 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17290) );
  NAND2_X1 U11741 ( .A1(n11546), .A2(n11718), .ZN(n11549) );
  OR2_X1 U11742 ( .A1(n11547), .A2(n18251), .ZN(n11548) );
  AOI22_X1 U11743 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18328), .B1(
        n11697), .B2(n11696), .ZN(n11709) );
  AND2_X1 U11744 ( .A1(n14376), .A2(n14364), .ZN(n14362) );
  NOR2_X1 U11745 ( .A1(n13753), .A2(n11918), .ZN(n13485) );
  NOR2_X2 U11746 ( .A1(n13751), .A2(n20180), .ZN(n13764) );
  AOI21_X1 U11747 ( .B1(n14543), .B2(n14542), .A(n14680), .ZN(n10311) );
  NAND2_X1 U11748 ( .A1(n10039), .A2(n16018), .ZN(n14622) );
  INV_X1 U11749 ( .A(n13439), .ZN(n16426) );
  OR2_X1 U11750 ( .A1(n13441), .A2(n16488), .ZN(n13444) );
  AND2_X1 U11751 ( .A1(n15121), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15122) );
  NAND2_X1 U11752 ( .A1(n14947), .A2(n14946), .ZN(n14949) );
  NOR2_X1 U11753 ( .A1(n15140), .A2(n11420), .ZN(n15116) );
  AOI21_X1 U11754 ( .B1(n10367), .B2(n9854), .A(n10365), .ZN(n10364) );
  NAND2_X1 U11755 ( .A1(n15290), .A2(n9898), .ZN(n10366) );
  INV_X1 U11756 ( .A(n15200), .ZN(n10365) );
  NAND2_X1 U11757 ( .A1(n15244), .A2(n15245), .ZN(n15234) );
  NOR2_X1 U11758 ( .A1(n15260), .A2(n15257), .ZN(n15244) );
  NAND2_X1 U11759 ( .A1(n10063), .A2(n10444), .ZN(n10062) );
  NAND2_X1 U11760 ( .A1(n10061), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10060) );
  OR2_X1 U11761 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10255) );
  INV_X1 U11762 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17222) );
  NOR3_X1 U11763 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n18972), .ZN(n11429) );
  INV_X1 U11764 ( .A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17287) );
  OAI211_X1 U11765 ( .C1(n9890), .C2(n15744), .A(n11456), .B(n11455), .ZN(
        n11719) );
  INV_X2 U11766 ( .A(n11447), .ZN(n17274) );
  INV_X1 U11767 ( .A(n13010), .ZN(n17641) );
  NOR2_X1 U11768 ( .A1(n9805), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10247) );
  INV_X1 U11769 ( .A(n18231), .ZN(n18776) );
  NAND2_X1 U11770 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18839), .ZN(n18828) );
  NOR2_X1 U11771 ( .A1(n13444), .A2(n16426), .ZN(n19014) );
  AND2_X1 U11772 ( .A1(n14258), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10172) );
  INV_X1 U11773 ( .A(n16495), .ZN(n17484) );
  OR2_X1 U11774 ( .A1(n12162), .A2(n12161), .ZN(n12669) );
  INV_X1 U11775 ( .A(n11983), .ZN(n12644) );
  AOI21_X1 U11776 ( .B1(n12735), .B2(n12734), .A(n12730), .ZN(n12768) );
  OR2_X1 U11777 ( .A1(n12106), .A2(n12105), .ZN(n12654) );
  NAND2_X1 U11778 ( .A1(n11022), .A2(n10357), .ZN(n11021) );
  NAND2_X1 U11779 ( .A1(n10766), .A2(n10765), .ZN(n10802) );
  NAND2_X1 U11780 ( .A1(n19470), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10765) );
  NAND2_X1 U11781 ( .A1(n10517), .A2(n13426), .ZN(n10537) );
  NAND3_X1 U11782 ( .A1(n10542), .A2(n10512), .A3(n10511), .ZN(n10567) );
  NAND2_X1 U11783 ( .A1(n9838), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10098) );
  AOI22_X1 U11784 ( .A1(n9842), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_7__4__SCAN_IN), .B2(n9815), .ZN(n10097) );
  OR2_X2 U11785 ( .A1(n13820), .A2(n14942), .ZN(n10627) );
  AOI21_X1 U11786 ( .B1(n10781), .B2(n10780), .A(n10779), .ZN(n10783) );
  XNOR2_X1 U11787 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10782) );
  NAND3_X1 U11788 ( .A1(n18964), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11436) );
  NAND2_X1 U11789 ( .A1(n20413), .A2(n11917), .ZN(n11939) );
  INV_X1 U11790 ( .A(n14387), .ZN(n10148) );
  NAND2_X1 U11791 ( .A1(n10023), .A2(n10025), .ZN(n10024) );
  NAND2_X1 U11792 ( .A1(n10023), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n10031) );
  NAND2_X1 U11793 ( .A1(n14291), .A2(n10342), .ZN(n10341) );
  INV_X1 U11794 ( .A(n14300), .ZN(n10342) );
  INV_X1 U11795 ( .A(n14495), .ZN(n10334) );
  INV_X1 U11796 ( .A(n12875), .ZN(n12840) );
  NOR2_X1 U11797 ( .A1(n10351), .A2(n14441), .ZN(n10350) );
  OR2_X1 U11798 ( .A1(n10355), .A2(n10353), .ZN(n10352) );
  INV_X1 U11799 ( .A(n14188), .ZN(n10353) );
  XNOR2_X1 U11800 ( .A(n12674), .B(n12205), .ZN(n12682) );
  NOR2_X1 U11801 ( .A1(n12263), .A2(n12206), .ZN(n12210) );
  AND2_X1 U11802 ( .A1(n20991), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12878) );
  NOR2_X2 U11803 ( .A1(n11928), .A2(n20991), .ZN(n12352) );
  NAND2_X1 U11804 ( .A1(n12719), .A2(n14680), .ZN(n14594) );
  NOR2_X1 U11805 ( .A1(n14189), .A2(n10157), .ZN(n10156) );
  INV_X1 U11806 ( .A(n14194), .ZN(n10157) );
  NOR2_X1 U11807 ( .A1(n10153), .A2(n10155), .ZN(n10152) );
  INV_X1 U11808 ( .A(n10154), .ZN(n10153) );
  INV_X1 U11809 ( .A(n14017), .ZN(n10155) );
  OR2_X1 U11810 ( .A1(n12764), .A2(n12046), .ZN(n12047) );
  AND2_X1 U11811 ( .A1(n13750), .A2(n13025), .ZN(n13914) );
  NOR2_X1 U11812 ( .A1(n13628), .A2(n10030), .ZN(n13637) );
  OAI21_X1 U11813 ( .B1(n21077), .B2(n20989), .A(n15835), .ZN(n20379) );
  NOR2_X1 U11814 ( .A1(n10230), .A2(n9955), .ZN(n10229) );
  INV_X1 U11815 ( .A(n10891), .ZN(n10230) );
  NOR2_X1 U11816 ( .A1(n10220), .A2(n9956), .ZN(n10219) );
  INV_X1 U11817 ( .A(n10221), .ZN(n10220) );
  NAND2_X1 U11818 ( .A1(n10872), .A2(n19129), .ZN(n10883) );
  INV_X1 U11819 ( .A(n13904), .ZN(n10207) );
  INV_X1 U11820 ( .A(n10492), .ZN(n10059) );
  AOI21_X1 U11821 ( .B1(n13241), .B2(n10274), .A(n9954), .ZN(n10273) );
  NAND2_X1 U11822 ( .A1(n15073), .A2(n10274), .ZN(n10272) );
  AND2_X1 U11823 ( .A1(n13186), .A2(n16273), .ZN(n10293) );
  NAND2_X1 U11824 ( .A1(n10180), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10178) );
  NOR2_X1 U11825 ( .A1(n19424), .A2(n10181), .ZN(n10180) );
  INV_X1 U11826 ( .A(n14867), .ZN(n10179) );
  NAND2_X1 U11827 ( .A1(n10597), .A2(n10571), .ZN(n10595) );
  INV_X1 U11828 ( .A(n10582), .ZN(n10594) );
  OR2_X1 U11829 ( .A1(n16223), .A2(n10858), .ZN(n10963) );
  NOR2_X1 U11830 ( .A1(n9857), .A2(n15202), .ZN(n15189) );
  AND2_X1 U11831 ( .A1(n10332), .A2(n10331), .ZN(n10330) );
  INV_X1 U11832 ( .A(n15064), .ZN(n10331) );
  NAND2_X1 U11833 ( .A1(n11176), .A2(n10205), .ZN(n10204) );
  INV_X1 U11834 ( .A(n15264), .ZN(n10205) );
  AND2_X1 U11835 ( .A1(n14901), .A2(n15100), .ZN(n10327) );
  INV_X1 U11836 ( .A(n15291), .ZN(n10110) );
  INV_X1 U11837 ( .A(n13977), .ZN(n11147) );
  INV_X1 U11838 ( .A(n13857), .ZN(n11132) );
  OR2_X1 U11839 ( .A1(n11074), .A2(n10858), .ZN(n11078) );
  NOR2_X1 U11840 ( .A1(n11217), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11228) );
  NOR2_X1 U11841 ( .A1(n10660), .A2(n10659), .ZN(n11231) );
  NAND2_X1 U11842 ( .A1(n13304), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13096) );
  NAND2_X1 U11843 ( .A1(n10497), .A2(n11089), .ZN(n11020) );
  INV_X1 U11844 ( .A(n10523), .ZN(n10497) );
  OR2_X2 U11845 ( .A1(n13820), .A2(n10596), .ZN(n10625) );
  AOI22_X1 U11846 ( .A1(n9838), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(n9807), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10432) );
  AOI22_X1 U11847 ( .A1(n9838), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(n9808), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10437) );
  INV_X1 U11848 ( .A(n10434), .ZN(n10435) );
  NAND2_X1 U11849 ( .A1(n10506), .A2(n10444), .ZN(n10416) );
  AOI21_X1 U11850 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n20140), .A(
        n10786), .ZN(n10971) );
  NOR2_X1 U11851 ( .A1(n18972), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11693) );
  OR2_X1 U11852 ( .A1(n15709), .A2(n9963), .ZN(n10005) );
  NOR2_X1 U11853 ( .A1(n11433), .A2(n18807), .ZN(n11471) );
  NOR3_X1 U11854 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n11432), .ZN(n11522) );
  INV_X1 U11855 ( .A(n18347), .ZN(n11669) );
  INV_X1 U11856 ( .A(n11538), .ZN(n10088) );
  XNOR2_X1 U11857 ( .A(n11534), .B(n11533), .ZN(n11535) );
  NOR2_X1 U11858 ( .A1(n10270), .A2(n10266), .ZN(n10265) );
  INV_X1 U11859 ( .A(n11642), .ZN(n10270) );
  INV_X1 U11860 ( .A(n11643), .ZN(n10271) );
  NAND2_X1 U11861 ( .A1(n13701), .A2(n13463), .ZN(n13501) );
  AND2_X1 U11862 ( .A1(n14408), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14029) );
  NAND2_X1 U11863 ( .A1(n10038), .A2(n10037), .ZN(n12957) );
  NAND2_X1 U11864 ( .A1(n12974), .A2(n14422), .ZN(n10038) );
  NAND2_X1 U11865 ( .A1(n15938), .A2(n9878), .ZN(n14801) );
  NAND2_X1 U11866 ( .A1(n12974), .A2(n10036), .ZN(n10035) );
  OR2_X1 U11867 ( .A1(n14131), .A2(n14130), .ZN(n14185) );
  OR2_X1 U11868 ( .A1(n13043), .A2(n13044), .ZN(n13618) );
  INV_X1 U11869 ( .A(n20180), .ZN(n13757) );
  XNOR2_X1 U11870 ( .A(n12896), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14549) );
  NAND2_X1 U11871 ( .A1(n10340), .A2(n10339), .ZN(n10338) );
  INV_X1 U11872 ( .A(n10341), .ZN(n10340) );
  INV_X1 U11873 ( .A(n13024), .ZN(n10339) );
  AND2_X1 U11874 ( .A1(n9928), .A2(n10344), .ZN(n10343) );
  INV_X1 U11875 ( .A(n14324), .ZN(n10344) );
  NAND2_X1 U11876 ( .A1(n12494), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12536) );
  AND2_X1 U11877 ( .A1(n12321), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12338) );
  CLKBUF_X1 U11878 ( .A(n14435), .Z(n14436) );
  AND2_X1 U11879 ( .A1(n14292), .A2(n12983), .ZN(n13033) );
  INV_X1 U11880 ( .A(n14739), .ZN(n10112) );
  AND2_X1 U11881 ( .A1(n14540), .A2(n14556), .ZN(n14548) );
  INV_X1 U11882 ( .A(n14314), .ZN(n10158) );
  NOR2_X1 U11883 ( .A1(n10162), .A2(n10161), .ZN(n14303) );
  INV_X1 U11884 ( .A(n14301), .ZN(n10161) );
  NAND2_X1 U11885 ( .A1(n10144), .A2(n16018), .ZN(n14612) );
  NAND2_X1 U11886 ( .A1(n10029), .A2(n10027), .ZN(n12948) );
  NAND2_X1 U11887 ( .A1(n12953), .A2(P1_EBX_REG_19__SCAN_IN), .ZN(n10029) );
  NAND2_X1 U11888 ( .A1(n12709), .A2(n10119), .ZN(n10118) );
  NOR2_X1 U11889 ( .A1(n15936), .A2(n15935), .ZN(n15938) );
  AND2_X1 U11890 ( .A1(n13782), .A2(n13781), .ZN(n16101) );
  INV_X1 U11891 ( .A(n13485), .ZN(n13771) );
  NAND2_X1 U11892 ( .A1(n12075), .A2(n21075), .ZN(n10048) );
  NAND2_X1 U11893 ( .A1(n12026), .A2(n12025), .ZN(n12073) );
  OR2_X1 U11894 ( .A1(n12764), .A2(n12023), .ZN(n12026) );
  XNOR2_X1 U11895 ( .A(n12052), .B(n12053), .ZN(n12065) );
  INV_X1 U11896 ( .A(n12109), .ZN(n10122) );
  INV_X1 U11897 ( .A(n20507), .ZN(n10141) );
  NAND2_X1 U11898 ( .A1(n12640), .A2(n13952), .ZN(n20629) );
  NOR2_X1 U11899 ( .A1(n20790), .A2(n20542), .ZN(n20721) );
  OR2_X1 U11900 ( .A1(n20763), .A2(n20762), .ZN(n20785) );
  NOR2_X1 U11901 ( .A1(n20714), .A2(n20542), .ZN(n20888) );
  NAND2_X1 U11902 ( .A1(n13948), .A2(n20377), .ZN(n20762) );
  NAND2_X1 U11903 ( .A1(n12640), .A2(n12108), .ZN(n20925) );
  AOI221_X1 U11904 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n10971), 
        .C1(n13676), .C2(n10971), .A(n10970), .ZN(n11011) );
  NOR2_X1 U11905 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n16463), .ZN(
        n10970) );
  NAND2_X1 U11906 ( .A1(n10526), .A2(n11030), .ZN(n11014) );
  AND2_X1 U11907 ( .A1(n10966), .A2(n10960), .ZN(n16202) );
  NAND2_X1 U11908 ( .A1(n10890), .A2(n10227), .ZN(n10888) );
  AND2_X1 U11909 ( .A1(n14860), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14888) );
  INV_X1 U11910 ( .A(n10897), .ZN(n10899) );
  NAND2_X1 U11911 ( .A1(n9941), .A2(n13976), .ZN(n10288) );
  AND2_X1 U11912 ( .A1(n13106), .A2(n19282), .ZN(n13107) );
  XNOR2_X1 U11913 ( .A(n10275), .B(n13287), .ZN(n14984) );
  INV_X1 U11914 ( .A(n16376), .ZN(n10323) );
  AND2_X1 U11915 ( .A1(n14888), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14890) );
  NAND2_X1 U11916 ( .A1(n16352), .A2(n11076), .ZN(n10306) );
  NAND2_X1 U11917 ( .A1(n10321), .A2(n14264), .ZN(n10315) );
  OR2_X1 U11918 ( .A1(n15040), .A2(n10318), .ZN(n10317) );
  NAND2_X1 U11919 ( .A1(n10358), .A2(n9897), .ZN(n14235) );
  NAND2_X1 U11920 ( .A1(n10962), .A2(n10216), .ZN(n10215) );
  OAI21_X1 U11921 ( .B1(n10969), .B2(n10858), .A(n11426), .ZN(n14234) );
  NAND2_X1 U11922 ( .A1(n15154), .A2(n10956), .ZN(n10064) );
  AND2_X1 U11923 ( .A1(n10309), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10308) );
  NOR2_X1 U11924 ( .A1(n16235), .A2(n10858), .ZN(n15178) );
  AND2_X1 U11925 ( .A1(n15481), .A2(n15482), .ZN(n10137) );
  OR3_X1 U11926 ( .A1(n10914), .A2(n10858), .A3(n15482), .ZN(n15503) );
  OR2_X1 U11927 ( .A1(n15214), .A2(n15534), .ZN(n10107) );
  NAND2_X1 U11928 ( .A1(n15514), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15513) );
  AND3_X1 U11929 ( .A1(n11377), .A2(n11376), .A3(n11375), .ZN(n15521) );
  OR3_X1 U11930 ( .A1(n10915), .A2(n10858), .A3(n15518), .ZN(n15533) );
  AOI21_X1 U11931 ( .B1(n15571), .B2(n9864), .A(n9906), .ZN(n10065) );
  NAND2_X1 U11932 ( .A1(n10191), .A2(n10190), .ZN(n10066) );
  AND3_X1 U11933 ( .A1(n11150), .A2(n11149), .A3(n11148), .ZN(n14006) );
  NAND2_X1 U11934 ( .A1(n11147), .A2(n9929), .ZN(n15303) );
  NOR2_X1 U11935 ( .A1(n16328), .A2(n16329), .ZN(n16327) );
  NAND2_X1 U11936 ( .A1(n11147), .A2(n11146), .ZN(n16324) );
  AND2_X1 U11937 ( .A1(n14087), .A2(n11109), .ZN(n15579) );
  AND2_X1 U11938 ( .A1(n11062), .A2(n14115), .ZN(n15316) );
  AND2_X1 U11939 ( .A1(n11044), .A2(n20027), .ZN(n11216) );
  NAND2_X1 U11940 ( .A1(n13089), .A2(n13537), .ZN(n13091) );
  XNOR2_X1 U11941 ( .A(n13095), .B(n13096), .ZN(n13589) );
  AOI21_X1 U11942 ( .B1(n19227), .B2(n13537), .A(n13094), .ZN(n13590) );
  NAND2_X1 U11943 ( .A1(n20122), .A2(n20160), .ZN(n19668) );
  NOR2_X2 U11944 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20126) );
  OR2_X1 U11945 ( .A1(n19611), .A2(n20130), .ZN(n20127) );
  NAND2_X1 U11946 ( .A1(n20132), .A2(n20160), .ZN(n19921) );
  INV_X1 U11947 ( .A(n10527), .ZN(n19447) );
  OR2_X1 U11948 ( .A1(n20122), .A2(n20160), .ZN(n19899) );
  INV_X1 U11949 ( .A(n19974), .ZN(n19673) );
  CLKBUF_X1 U11950 ( .A(n11016), .Z(n11017) );
  OR2_X1 U11951 ( .A1(n16733), .A2(n16991), .ZN(n10075) );
  NOR2_X1 U11952 ( .A1(n16734), .A2(n16735), .ZN(n16733) );
  INV_X1 U11953 ( .A(n17704), .ZN(n10076) );
  NOR2_X1 U11954 ( .A1(n16777), .A2(n17718), .ZN(n16776) );
  INV_X1 U11955 ( .A(n17336), .ZN(n10263) );
  OR2_X1 U11956 ( .A1(n11503), .A2(n9910), .ZN(n10004) );
  NAND2_X1 U11957 ( .A1(n11470), .A2(n11469), .ZN(n11478) );
  AOI21_X1 U11958 ( .B1(n17268), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n11468), .ZN(n11469) );
  NOR2_X1 U11959 ( .A1(n9888), .A2(n15712), .ZN(n11468) );
  NAND2_X1 U11960 ( .A1(n10017), .A2(n11585), .ZN(n10016) );
  NOR2_X1 U11961 ( .A1(n17714), .A2(n16665), .ZN(n17664) );
  NOR2_X1 U11962 ( .A1(n17833), .A2(n16668), .ZN(n17786) );
  AOI21_X1 U11963 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17734), .A(
        n18719), .ZN(n17834) );
  NOR2_X1 U11964 ( .A1(n15838), .A2(n17886), .ZN(n11565) );
  NOR2_X1 U11965 ( .A1(n17797), .A2(n18113), .ZN(n10249) );
  OR2_X1 U11966 ( .A1(n17782), .A2(n18127), .ZN(n10090) );
  NAND2_X1 U11967 ( .A1(n17928), .A2(n11545), .ZN(n17921) );
  NAND2_X1 U11968 ( .A1(n17967), .A2(n17968), .ZN(n17966) );
  AOI22_X1 U11969 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11595) );
  NAND2_X1 U11970 ( .A1(n15828), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20180) );
  INV_X1 U11971 ( .A(n20660), .ZN(n20881) );
  INV_X1 U11972 ( .A(n14527), .ZN(n14532) );
  AOI21_X1 U11973 ( .B1(n16033), .B2(n14316), .A(n12786), .ZN(n12787) );
  INV_X1 U11974 ( .A(n16031), .ZN(n16033) );
  OR3_X1 U11975 ( .A1(n15816), .A2(n13751), .A3(n20180), .ZN(n20187) );
  OR2_X1 U11976 ( .A1(n21068), .A2(n13960), .ZN(n14689) );
  XNOR2_X1 U11977 ( .A(n12722), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14755) );
  NAND2_X1 U11978 ( .A1(n20565), .A2(n12049), .ZN(n20660) );
  OR2_X1 U11979 ( .A1(n19014), .A2(n14156), .ZN(n19222) );
  AND2_X1 U11980 ( .A1(n19014), .A2(n14147), .ZN(n19226) );
  OAI211_X1 U11981 ( .C1(n15161), .C2(n9993), .A(n10302), .B(n10301), .ZN(
        n14277) );
  NAND2_X1 U11982 ( .A1(n10303), .A2(n14258), .ZN(n10302) );
  XNOR2_X1 U11983 ( .A(n14144), .B(n14143), .ZN(n14276) );
  NAND2_X1 U11984 ( .A1(n15122), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14144) );
  NOR2_X1 U11985 ( .A1(n15513), .A2(n15501), .ZN(n15479) );
  AND2_X1 U11986 ( .A1(n19425), .A2(n20148), .ZN(n16363) );
  INV_X1 U11987 ( .A(n19421), .ZN(n16371) );
  AND2_X1 U11988 ( .A1(n19425), .A2(n13544), .ZN(n19413) );
  INV_X1 U11989 ( .A(n19413), .ZN(n16355) );
  OR2_X1 U11990 ( .A1(n13536), .A2(n14159), .ZN(n19417) );
  XNOR2_X1 U11991 ( .A(n14949), .B(n14260), .ZN(n16260) );
  NAND2_X1 U11992 ( .A1(n10300), .A2(n10304), .ZN(n15115) );
  AOI21_X1 U11993 ( .B1(n15323), .B2(n15325), .A(n15322), .ZN(n15324) );
  NAND2_X1 U11994 ( .A1(n14949), .A2(n14948), .ZN(n15330) );
  OR2_X1 U11995 ( .A1(n14947), .A2(n14946), .ZN(n14948) );
  NAND2_X1 U11996 ( .A1(n15234), .A2(n15233), .ZN(n10192) );
  INV_X1 U11997 ( .A(n20130), .ZN(n20152) );
  INV_X1 U11998 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20147) );
  INV_X1 U11999 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20140) );
  INV_X1 U12000 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20136) );
  NOR2_X1 U12001 ( .A1(n19921), .A2(n19920), .ZN(n19964) );
  NOR2_X1 U12002 ( .A1(n16690), .A2(n16691), .ZN(n16689) );
  AOI21_X1 U12003 ( .B1(n16690), .B2(n16691), .A(n18842), .ZN(n10071) );
  AOI211_X1 U12004 ( .C1(P3_REIP_REG_29__SCAN_IN), .C2(n16694), .A(n16693), 
        .B(n10069), .ZN(n10068) );
  NOR2_X1 U12005 ( .A1(n16698), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n10069) );
  NAND2_X1 U12006 ( .A1(n17135), .A2(P3_EBX_REG_21__SCAN_IN), .ZN(n17120) );
  AOI22_X1 U12007 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11637) );
  AOI211_X1 U12008 ( .C1(n17293), .C2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n11635), .B(n11634), .ZN(n11636) );
  NOR2_X1 U12009 ( .A1(n17167), .A2(n16802), .ZN(n17166) );
  NOR2_X2 U12010 ( .A1(n17250), .A2(n17249), .ZN(n17247) );
  NAND2_X1 U12011 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(P3_EBX_REG_7__SCAN_IN), 
        .ZN(n10262) );
  INV_X1 U12012 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17354) );
  NAND4_X1 U12013 ( .A1(n18991), .A2(n18993), .A3(n17516), .A4(n15868), .ZN(
        n17360) );
  NOR2_X2 U12014 ( .A1(n18366), .A2(n17360), .ZN(n17361) );
  NAND2_X1 U12015 ( .A1(n18796), .A2(n17514), .ZN(n17504) );
  OAI211_X1 U12016 ( .C1(n11565), .C2(n15840), .A(n10235), .B(n10234), .ZN(
        n10233) );
  INV_X1 U12017 ( .A(n11566), .ZN(n10234) );
  OR2_X1 U12018 ( .A1(n15839), .A2(n18951), .ZN(n10235) );
  NOR2_X1 U12019 ( .A1(n17834), .A2(n10015), .ZN(n10014) );
  INV_X1 U12020 ( .A(n17746), .ZN(n10015) );
  NAND3_X1 U12021 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n16655), .A3(n17988), 
        .ZN(n17841) );
  NAND2_X1 U12022 ( .A1(n10236), .A2(n11566), .ZN(n10082) );
  OAI21_X1 U12023 ( .B1(n10238), .B2(n11565), .A(n10237), .ZN(n10236) );
  INV_X1 U12024 ( .A(n11678), .ZN(n10237) );
  OR2_X1 U12025 ( .A1(n15839), .A2(n11675), .ZN(n10238) );
  AND2_X1 U12026 ( .A1(n10233), .A2(n10080), .ZN(n10079) );
  NOR2_X1 U12027 ( .A1(n13017), .A2(n10081), .ZN(n10080) );
  AND2_X1 U12028 ( .A1(n10083), .A2(n9802), .ZN(n10078) );
  INV_X1 U12029 ( .A(n11715), .ZN(n10084) );
  NOR2_X1 U12030 ( .A1(n16530), .A2(n18776), .ZN(n10254) );
  NAND2_X1 U12031 ( .A1(n13018), .A2(n15781), .ZN(n10250) );
  AND2_X1 U12032 ( .A1(n13022), .A2(n17628), .ZN(n10251) );
  NOR2_X2 U12033 ( .A1(n10081), .A2(n13017), .ZN(n18219) );
  INV_X1 U12034 ( .A(n11909), .ZN(n11961) );
  NAND2_X1 U12035 ( .A1(n11883), .A2(n10117), .ZN(n13627) );
  AND2_X1 U12036 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10370) );
  NOR2_X1 U12037 ( .A1(n10057), .A2(n10056), .ZN(n10055) );
  NAND2_X1 U12038 ( .A1(n10721), .A2(n10720), .ZN(n10058) );
  AOI21_X1 U12039 ( .B1(n10703), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n10704), .ZN(n10712) );
  NAND2_X1 U12040 ( .A1(n9807), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10199) );
  NAND2_X1 U12041 ( .A1(n9842), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10197) );
  NOR2_X1 U12042 ( .A1(n10410), .A2(n10196), .ZN(n10195) );
  AND2_X1 U12043 ( .A1(n16432), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10198) );
  NAND2_X1 U12044 ( .A1(n9838), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n10422) );
  NAND2_X1 U12045 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n10423) );
  AOI22_X1 U12046 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9816), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10425) );
  AOI22_X1 U12047 ( .A1(n9838), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10421), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10420) );
  AOI22_X1 U12048 ( .A1(n9840), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10634), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10418) );
  AOI21_X1 U12049 ( .B1(n9814), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A(
        n10444), .ZN(n10451) );
  NAND2_X1 U12050 ( .A1(n13391), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n10450) );
  OAI21_X1 U12051 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n10256), .A(
        n11687), .ZN(n11688) );
  AND2_X1 U12052 ( .A1(n11867), .A2(n11929), .ZN(n11887) );
  AND2_X2 U12053 ( .A1(n10020), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11770) );
  OR2_X1 U12054 ( .A1(n12133), .A2(n12132), .ZN(n12666) );
  OR2_X1 U12055 ( .A1(n12044), .A2(n12043), .ZN(n12642) );
  NAND2_X1 U12056 ( .A1(n12881), .A2(n12992), .ZN(n11930) );
  OR3_X1 U12057 ( .A1(n12761), .A2(n12760), .A3(n12885), .ZN(n12762) );
  AND2_X1 U12058 ( .A1(n13627), .A2(n10023), .ZN(n10030) );
  AOI22_X1 U12059 ( .A1(n9810), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12517), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11760) );
  NAND2_X1 U12060 ( .A1(n11023), .A2(n11217), .ZN(n11024) );
  NAND2_X1 U12061 ( .A1(n14999), .A2(n16222), .ZN(n10232) );
  INV_X1 U12062 ( .A(n14993), .ZN(n10274) );
  INV_X1 U12063 ( .A(n10457), .ZN(n10458) );
  NOR2_X1 U12064 ( .A1(n10129), .A2(n14159), .ZN(n10128) );
  NAND2_X1 U12065 ( .A1(n9820), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10129) );
  AOI22_X1 U12066 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10703), .B1(
        n10817), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10682) );
  AOI22_X1 U12067 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n10823), .B1(
        n10818), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10679) );
  AOI22_X1 U12068 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n10716), .B1(
        n19863), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10683) );
  OR2_X1 U12069 ( .A1(n10675), .A2(n10674), .ZN(n11237) );
  AND2_X1 U12070 ( .A1(n11021), .A2(n11217), .ZN(n10533) );
  INV_X1 U12071 ( .A(n19437), .ZN(n11089) );
  NAND2_X1 U12072 ( .A1(n10609), .A2(n10608), .ZN(n10619) );
  INV_X1 U12073 ( .A(n10616), .ZN(n10618) );
  AOI22_X1 U12074 ( .A1(n9838), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(n9808), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10477) );
  AOI21_X1 U12075 ( .B1(n9816), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A(n9869), 
        .ZN(n10406) );
  AND2_X1 U12076 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n9998) );
  AOI21_X1 U12077 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18801), .A(
        n11686), .ZN(n11692) );
  AND2_X1 U12078 ( .A1(n11706), .A2(n11693), .ZN(n11686) );
  AOI21_X1 U12079 ( .B1(n17291), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n10269), .ZN(n10268) );
  OAI22_X1 U12080 ( .A1(n17312), .A2(n17253), .B1(n17197), .B2(n17252), .ZN(
        n10269) );
  NAND2_X1 U12081 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10267) );
  INV_X1 U12082 ( .A(n11883), .ZN(n11941) );
  NAND2_X1 U12083 ( .A1(n10023), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n10037) );
  AND2_X1 U12084 ( .A1(n10151), .A2(n9974), .ZN(n10150) );
  NAND2_X1 U12085 ( .A1(n10023), .A2(P1_EBX_REG_8__SCAN_IN), .ZN(n10034) );
  AND2_X1 U12086 ( .A1(n10376), .A2(n10346), .ZN(n10345) );
  INV_X1 U12087 ( .A(n14348), .ZN(n10346) );
  NOR2_X1 U12088 ( .A1(n14503), .A2(n14437), .ZN(n10335) );
  NOR2_X1 U12089 ( .A1(n10349), .A2(n10348), .ZN(n10347) );
  INV_X1 U12090 ( .A(n10350), .ZN(n10349) );
  NAND2_X1 U12091 ( .A1(n10356), .A2(n10379), .ZN(n10355) );
  INV_X1 U12092 ( .A(n14191), .ZN(n10356) );
  INV_X1 U12093 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12111) );
  NAND2_X1 U12094 ( .A1(n10023), .A2(n10028), .ZN(n10027) );
  OAI21_X1 U12095 ( .B1(n12665), .B2(n12690), .A(n12671), .ZN(n12672) );
  NOR2_X1 U12096 ( .A1(n13989), .A2(n13887), .ZN(n10154) );
  INV_X1 U12097 ( .A(n12642), .ZN(n12050) );
  OR2_X1 U12098 ( .A1(n12644), .A2(n12092), .ZN(n11981) );
  OR2_X1 U12099 ( .A1(n11980), .A2(n11979), .ZN(n11983) );
  AND2_X1 U12100 ( .A1(n12772), .A2(n13610), .ZN(n12766) );
  NAND2_X1 U12101 ( .A1(n11989), .A2(n11987), .ZN(n10143) );
  AND4_X1 U12102 ( .A1(n11843), .A2(n11842), .A3(n11841), .A4(n11840), .ZN(
        n11849) );
  OR2_X1 U12103 ( .A1(n9850), .A2(n11860), .ZN(n11861) );
  AOI22_X1 U12104 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        P1_INSTQUEUE_REG_10__3__SCAN_IN), .B2(n11973), .ZN(n11850) );
  NAND2_X1 U12105 ( .A1(n20659), .A2(n21075), .ZN(n10140) );
  NAND2_X1 U12106 ( .A1(n9875), .A2(n11217), .ZN(n11032) );
  OR3_X1 U12107 ( .A1(n10934), .A2(n10232), .A3(P2_EBX_REG_26__SCAN_IN), .ZN(
        n10231) );
  NAND2_X1 U12108 ( .A1(n10957), .A2(n10958), .ZN(n10966) );
  NOR3_X1 U12109 ( .A1(n10935), .A2(n10934), .A3(P2_EBX_REG_24__SCAN_IN), .ZN(
        n10949) );
  NOR2_X1 U12110 ( .A1(n10935), .A2(n10934), .ZN(n10945) );
  AND2_X1 U12111 ( .A1(n14142), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14860) );
  NOR2_X1 U12112 ( .A1(n10885), .A2(n10222), .ZN(n10221) );
  INV_X1 U12113 ( .A(n10881), .ZN(n10222) );
  AND2_X1 U12114 ( .A1(n10285), .A2(n14964), .ZN(n10284) );
  INV_X1 U12115 ( .A(n14972), .ZN(n10285) );
  NAND4_X2 U12116 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n15662), .A4(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13177) );
  CLKBUF_X1 U12117 ( .A(n13312), .Z(n13320) );
  INV_X1 U12118 ( .A(n10284), .ZN(n10279) );
  NOR2_X1 U12119 ( .A1(n14954), .A2(n10282), .ZN(n10281) );
  INV_X1 U12120 ( .A(n14964), .ZN(n10282) );
  AND2_X1 U12121 ( .A1(n19447), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13077) );
  NOR2_X1 U12122 ( .A1(n19141), .A2(n10175), .ZN(n10174) );
  INV_X1 U12123 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10175) );
  AOI21_X1 U12124 ( .B1(n10694), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n10643), .ZN(n10644) );
  NAND2_X1 U12125 ( .A1(n10642), .A2(n10641), .ZN(n10643) );
  INV_X1 U12126 ( .A(n14264), .ZN(n10318) );
  NAND2_X1 U12127 ( .A1(n15028), .A2(n13422), .ZN(n10322) );
  INV_X1 U12128 ( .A(n10957), .ZN(n14245) );
  NAND2_X1 U12129 ( .A1(n10218), .A2(n10961), .ZN(n10962) );
  INV_X1 U12130 ( .A(n15137), .ZN(n10218) );
  AND2_X1 U12131 ( .A1(n15137), .A2(n10217), .ZN(n10216) );
  NAND2_X1 U12132 ( .A1(n15148), .A2(n10961), .ZN(n10217) );
  NOR2_X1 U12133 ( .A1(n10955), .A2(n10954), .ZN(n10956) );
  AND2_X1 U12134 ( .A1(n14987), .A2(n14980), .ZN(n10213) );
  AND2_X1 U12135 ( .A1(n15413), .A2(n15075), .ZN(n10332) );
  AND2_X1 U12136 ( .A1(n9883), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10309) );
  AND2_X1 U12137 ( .A1(n19053), .A2(n14246), .ZN(n10919) );
  INV_X1 U12138 ( .A(n15503), .ZN(n10105) );
  AND2_X1 U12139 ( .A1(n9929), .A2(n10209), .ZN(n10208) );
  INV_X1 U12140 ( .A(n15302), .ZN(n10209) );
  NOR2_X1 U12141 ( .A1(n10189), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10190) );
  AOI21_X1 U12142 ( .B1(n15575), .B2(n10880), .A(n15546), .ZN(n10188) );
  AND2_X1 U12143 ( .A1(n15592), .A2(n9927), .ZN(n10362) );
  NOR2_X1 U12144 ( .A1(n14924), .A2(n10325), .ZN(n10324) );
  INV_X1 U12145 ( .A(n16400), .ZN(n10325) );
  AND2_X1 U12146 ( .A1(n11071), .A2(n15314), .ZN(n11065) );
  OR2_X1 U12147 ( .A1(n10841), .A2(n10840), .ZN(n11258) );
  OAI21_X1 U12148 ( .B1(n11064), .B2(n14246), .A(n19178), .ZN(n10852) );
  AND3_X1 U12149 ( .A1(n11130), .A2(n11129), .A3(n11128), .ZN(n13874) );
  INV_X1 U12150 ( .A(n11237), .ZN(n11051) );
  NAND2_X1 U12151 ( .A1(n10760), .A2(n10759), .ZN(n10803) );
  NAND2_X1 U12152 ( .A1(n11231), .A2(n11219), .ZN(n10760) );
  NAND2_X1 U12153 ( .A1(n10294), .A2(n10126), .ZN(n10546) );
  INV_X1 U12154 ( .A(n10545), .ZN(n10294) );
  INV_X1 U12155 ( .A(n10544), .ZN(n10126) );
  NAND2_X1 U12156 ( .A1(n13426), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n10314) );
  OR2_X1 U12157 ( .A1(n10778), .A2(n10777), .ZN(n11245) );
  NAND2_X1 U12158 ( .A1(n11088), .A2(n10378), .ZN(n11207) );
  NAND2_X1 U12159 ( .A1(n13071), .A2(n20136), .ZN(n13092) );
  NOR2_X1 U12160 ( .A1(n13332), .A2(n19457), .ZN(n13087) );
  AND2_X2 U12161 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15659) );
  NAND2_X1 U12162 ( .A1(n13088), .A2(n13087), .ZN(n13100) );
  NAND2_X1 U12163 ( .A1(n10405), .A2(n10404), .ZN(n10531) );
  INV_X1 U12164 ( .A(n10492), .ZN(n10530) );
  OR2_X1 U12165 ( .A1(n10786), .A2(n10784), .ZN(n10994) );
  AND2_X1 U12166 ( .A1(n17268), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n9999) );
  NAND2_X1 U12167 ( .A1(n10011), .A2(n10010), .ZN(n10009) );
  INV_X1 U12168 ( .A(n15718), .ZN(n10011) );
  AND2_X1 U12169 ( .A1(n17268), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n10001) );
  AND2_X1 U12170 ( .A1(n11474), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n10000) );
  AND2_X1 U12171 ( .A1(n17268), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n10003) );
  AND2_X1 U12172 ( .A1(n17268), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n10002) );
  AOI22_X1 U12173 ( .A1(n9812), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11474), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11585) );
  AOI21_X1 U12174 ( .B1(n17292), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n10018), .ZN(n10017) );
  NOR2_X1 U12175 ( .A1(n11638), .A2(n17317), .ZN(n10018) );
  NAND2_X1 U12176 ( .A1(n11444), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11579) );
  AND4_X1 U12177 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16667) );
  NAND2_X1 U12178 ( .A1(n17899), .A2(n11553), .ZN(n11556) );
  AOI211_X1 U12179 ( .C1(n17293), .C2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n11574), .B(n11573), .ZN(n11575) );
  AOI211_X1 U12180 ( .C1(n17293), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n11614), .B(n11613), .ZN(n11615) );
  INV_X1 U12181 ( .A(n11654), .ZN(n11672) );
  NOR3_X1 U12182 ( .A1(n11671), .A2(n11701), .A3(n11663), .ZN(n11659) );
  AND2_X1 U12183 ( .A1(n12889), .A2(n12888), .ZN(n13480) );
  NAND2_X1 U12184 ( .A1(n10023), .A2(n21097), .ZN(n12943) );
  NOR2_X1 U12185 ( .A1(n21382), .A2(n15934), .ZN(n15920) );
  NOR2_X1 U12186 ( .A1(n21302), .A2(n15955), .ZN(n15939) );
  INV_X1 U12187 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n20219) );
  NAND2_X1 U12188 ( .A1(n20276), .A2(n14408), .ZN(n20250) );
  NAND2_X1 U12189 ( .A1(n10023), .A2(n21313), .ZN(n12972) );
  NAND2_X1 U12190 ( .A1(n14362), .A2(n10159), .ZN(n14327) );
  AND2_X1 U12191 ( .A1(n12963), .A2(n12962), .ZN(n14349) );
  NAND2_X1 U12192 ( .A1(n14362), .A2(n14349), .ZN(n14351) );
  AND2_X1 U12193 ( .A1(n14424), .A2(n9977), .ZN(n14376) );
  NAND2_X1 U12194 ( .A1(n14424), .A2(n10149), .ZN(n15853) );
  NAND2_X1 U12195 ( .A1(n10026), .A2(n10024), .ZN(n12920) );
  NAND2_X1 U12196 ( .A1(n12953), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n10026) );
  NAND2_X1 U12197 ( .A1(n10032), .A2(n10031), .ZN(n12906) );
  NAND2_X1 U12198 ( .A1(n12974), .A2(n10033), .ZN(n10032) );
  AOI21_X1 U12199 ( .B1(n12675), .B2(n12352), .A(n12198), .ZN(n14068) );
  OR2_X1 U12200 ( .A1(n12846), .A2(n14565), .ZN(n12895) );
  AOI22_X1 U12201 ( .A1(n12845), .A2(n12844), .B1(n12843), .B2(n14567), .ZN(
        n14291) );
  NAND2_X1 U12202 ( .A1(n12582), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12789) );
  AND2_X1 U12203 ( .A1(n14599), .A2(n12843), .ZN(n12577) );
  NOR2_X1 U12204 ( .A1(n12536), .A2(n14615), .ZN(n12537) );
  NAND2_X1 U12205 ( .A1(n12537), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12580) );
  AND2_X1 U12206 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n12493), .ZN(
        n12494) );
  AND2_X1 U12207 ( .A1(n12499), .A2(n12498), .ZN(n14372) );
  NOR2_X1 U12208 ( .A1(n12434), .A2(n14642), .ZN(n12435) );
  NAND2_X1 U12209 ( .A1(n12415), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12434) );
  CLKBUF_X1 U12210 ( .A(n14427), .Z(n14428) );
  NOR2_X1 U12211 ( .A1(n12379), .A2(n12339), .ZN(n12380) );
  NAND2_X1 U12212 ( .A1(n12338), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12379) );
  INV_X1 U12213 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12302) );
  AND2_X1 U12214 ( .A1(n12267), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12268) );
  NAND2_X1 U12215 ( .A1(n12285), .A2(n12284), .ZN(n14449) );
  NOR2_X1 U12216 ( .A1(n12248), .A2(n12247), .ZN(n12267) );
  INV_X1 U12217 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12247) );
  OR2_X1 U12218 ( .A1(n12229), .A2(n20219), .ZN(n12248) );
  NAND2_X1 U12219 ( .A1(n12207), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12229) );
  NOR2_X1 U12220 ( .A1(n12210), .A2(n12209), .ZN(n12211) );
  AND2_X1 U12221 ( .A1(n12191), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12207) );
  AND2_X1 U12222 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n12138), .ZN(
        n12167) );
  INV_X1 U12223 ( .A(n13897), .ZN(n12081) );
  NAND2_X1 U12224 ( .A1(n10023), .A2(n21410), .ZN(n12981) );
  NOR2_X1 U12225 ( .A1(n10144), .A2(n10114), .ZN(n10113) );
  INV_X1 U12226 ( .A(n14585), .ZN(n10114) );
  OR2_X1 U12227 ( .A1(n14648), .A2(n9989), .ZN(n14629) );
  NAND2_X1 U12228 ( .A1(n14424), .A2(n12949), .ZN(n15855) );
  NAND2_X1 U12229 ( .A1(n14648), .A2(n14647), .ZN(n14646) );
  NOR2_X1 U12230 ( .A1(n16097), .A2(n14696), .ZN(n14813) );
  NAND2_X1 U12231 ( .A1(n15938), .A2(n10151), .ZN(n15919) );
  NAND2_X1 U12232 ( .A1(n10023), .A2(n21299), .ZN(n12933) );
  AND2_X1 U12233 ( .A1(n15938), .A2(n14444), .ZN(n15917) );
  NAND2_X1 U12234 ( .A1(n14195), .A2(n9877), .ZN(n15936) );
  NOR2_X1 U12235 ( .A1(n14185), .A2(n14184), .ZN(n14195) );
  NAND2_X1 U12236 ( .A1(n10023), .A2(n21142), .ZN(n12924) );
  NAND2_X1 U12237 ( .A1(n14195), .A2(n14194), .ZN(n14197) );
  NAND2_X1 U12238 ( .A1(n10023), .A2(n21376), .ZN(n12915) );
  AND2_X1 U12239 ( .A1(n12910), .A2(n10152), .ZN(n14050) );
  NAND2_X1 U12240 ( .A1(n12910), .A2(n12909), .ZN(n13988) );
  XNOR2_X1 U12241 ( .A(n13694), .B(n12636), .ZN(n13749) );
  NAND2_X1 U12242 ( .A1(n14825), .A2(n21075), .ZN(n12784) );
  NAND2_X1 U12243 ( .A1(n12983), .A2(n12903), .ZN(n12902) );
  AND2_X1 U12244 ( .A1(n13783), .A2(n13780), .ZN(n20360) );
  NAND2_X1 U12245 ( .A1(n13783), .A2(n13914), .ZN(n20361) );
  NAND2_X1 U12246 ( .A1(n12056), .A2(n12055), .ZN(n12084) );
  OR2_X1 U12247 ( .A1(n12052), .A2(n12054), .ZN(n12055) );
  INV_X1 U12248 ( .A(n12108), .ZN(n13952) );
  INV_X1 U12249 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13928) );
  NAND2_X1 U12250 ( .A1(n10333), .A2(n11960), .ZN(n13622) );
  AND3_X1 U12251 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21075), .A3(n20379), 
        .ZN(n20444) );
  INV_X1 U12252 ( .A(n20590), .ZN(n20880) );
  NAND2_X1 U12253 ( .A1(n20374), .A2(n20373), .ZN(n20440) );
  NAND2_X1 U12254 ( .A1(n20374), .A2(n20372), .ZN(n20441) );
  AOI21_X1 U12255 ( .B1(n20843), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n20542), 
        .ZN(n20932) );
  AND2_X1 U12256 ( .A1(n16145), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15828) );
  INV_X1 U12257 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n10226) );
  NAND2_X1 U12258 ( .A1(n10929), .A2(n10930), .ZN(n10935) );
  AND2_X1 U12259 ( .A1(n10890), .A2(n10229), .ZN(n10896) );
  NAND2_X1 U12260 ( .A1(n19182), .A2(n9934), .ZN(n19037) );
  NAND2_X1 U12261 ( .A1(n10882), .A2(n10219), .ZN(n10903) );
  AND2_X1 U12262 ( .A1(n19470), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10885) );
  NAND2_X1 U12263 ( .A1(n10882), .A2(n10881), .ZN(n10886) );
  AND2_X1 U12264 ( .A1(n19470), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10856) );
  AND3_X1 U12265 ( .A1(n11186), .A2(n11185), .A3(n11184), .ZN(n15202) );
  OR2_X1 U12266 ( .A1(n11279), .A2(n11278), .ZN(n13106) );
  AND3_X1 U12267 ( .A1(n11135), .A2(n11134), .A3(n11133), .ZN(n13904) );
  NAND2_X1 U12268 ( .A1(n11132), .A2(n11131), .ZN(n13905) );
  NOR2_X1 U12269 ( .A1(n14159), .A2(n11025), .ZN(n10127) );
  INV_X1 U12270 ( .A(n15028), .ZN(n10319) );
  AND2_X1 U12271 ( .A1(n13331), .A2(n13338), .ZN(n14962) );
  AND2_X1 U12272 ( .A1(n10330), .A2(n10329), .ZN(n10328) );
  INV_X1 U12273 ( .A(n15054), .ZN(n10329) );
  AND2_X1 U12274 ( .A1(n15412), .A2(n15413), .ZN(n15415) );
  OR2_X1 U12275 ( .A1(n13264), .A2(n9957), .ZN(n10291) );
  AND2_X1 U12276 ( .A1(n13562), .A2(n20041), .ZN(n19372) );
  NAND2_X1 U12277 ( .A1(n10184), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10183) );
  NOR2_X1 U12278 ( .A1(n16198), .A2(n10185), .ZN(n10184) );
  INV_X1 U12279 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10185) );
  INV_X1 U12280 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16198) );
  NOR3_X1 U12281 ( .A1(n15168), .A2(n15158), .A3(n16198), .ZN(n15149) );
  OR2_X1 U12282 ( .A1(n15182), .A2(n15171), .ZN(n15168) );
  AND2_X1 U12283 ( .A1(n14890), .A2(n9978), .ZN(n15193) );
  AND3_X1 U12284 ( .A1(n11189), .A2(n11188), .A3(n11187), .ZN(n15190) );
  NAND2_X1 U12285 ( .A1(n14890), .A2(n9881), .ZN(n15205) );
  AND2_X1 U12286 ( .A1(n14890), .A2(n9961), .ZN(n15206) );
  AND2_X1 U12287 ( .A1(n14890), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14858) );
  NOR2_X1 U12288 ( .A1(n14881), .A2(n19091), .ZN(n14880) );
  AND3_X1 U12289 ( .A1(n11160), .A2(n11159), .A3(n11158), .ZN(n15523) );
  NAND2_X1 U12290 ( .A1(n14878), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14881) );
  AND2_X1 U12291 ( .A1(n14874), .A2(n10173), .ZN(n14878) );
  AND2_X1 U12292 ( .A1(n9876), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10173) );
  NAND2_X1 U12293 ( .A1(n14874), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14876) );
  AND2_X1 U12294 ( .A1(n14873), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14874) );
  NOR2_X1 U12295 ( .A1(n14872), .A2(n16351), .ZN(n14873) );
  INV_X1 U12296 ( .A(n16354), .ZN(n10134) );
  NAND2_X1 U12297 ( .A1(n10179), .A2(n10177), .ZN(n14872) );
  NOR2_X1 U12298 ( .A1(n10178), .A2(n10182), .ZN(n10177) );
  INV_X1 U12299 ( .A(n10178), .ZN(n10176) );
  NAND2_X1 U12300 ( .A1(n10179), .A2(n10180), .ZN(n14870) );
  NOR2_X1 U12301 ( .A1(n14867), .A2(n19424), .ZN(n14871) );
  NAND2_X1 U12302 ( .A1(n14078), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14867) );
  XNOR2_X1 U12303 ( .A(n10594), .B(n10593), .ZN(n10124) );
  AND2_X1 U12304 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14078) );
  AND2_X1 U12305 ( .A1(n13443), .A2(n13442), .ZN(n13535) );
  NOR2_X1 U12306 ( .A1(n9862), .A2(n14241), .ZN(n14242) );
  NAND2_X1 U12307 ( .A1(n14262), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10305) );
  NOR2_X1 U12308 ( .A1(n14961), .A2(n11206), .ZN(n14947) );
  NAND2_X1 U12309 ( .A1(n14997), .A2(n10211), .ZN(n14961) );
  AND2_X1 U12310 ( .A1(n9959), .A2(n10212), .ZN(n10211) );
  INV_X1 U12311 ( .A(n14959), .ZN(n10212) );
  NOR2_X1 U12312 ( .A1(n16189), .A2(n10858), .ZN(n15137) );
  INV_X1 U12313 ( .A(n15135), .ZN(n15133) );
  AND2_X1 U12314 ( .A1(n10964), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15166) );
  NAND2_X1 U12315 ( .A1(n15189), .A2(n11190), .ZN(n15192) );
  INV_X1 U12316 ( .A(n15190), .ZN(n11190) );
  AND3_X1 U12317 ( .A1(n11193), .A2(n11192), .A3(n11191), .ZN(n14996) );
  NOR2_X1 U12318 ( .A1(n15192), .A2(n14996), .ZN(n14997) );
  NAND2_X1 U12319 ( .A1(n15412), .A2(n10330), .ZN(n15066) );
  INV_X1 U12320 ( .A(n15292), .ZN(n10369) );
  NAND2_X1 U12321 ( .A1(n10201), .A2(n14894), .ZN(n10200) );
  INV_X1 U12322 ( .A(n10202), .ZN(n10201) );
  NOR2_X1 U12323 ( .A1(n15265), .A2(n10202), .ZN(n15238) );
  AND3_X1 U12324 ( .A1(n11175), .A2(n11174), .A3(n11173), .ZN(n15009) );
  NOR2_X1 U12325 ( .A1(n15265), .A2(n10204), .ZN(n15236) );
  NAND2_X1 U12326 ( .A1(n14902), .A2(n9879), .ZN(n15465) );
  INV_X1 U12327 ( .A(n15462), .ZN(n10326) );
  AND3_X1 U12328 ( .A1(n11172), .A2(n11171), .A3(n11170), .ZN(n15264) );
  NAND2_X1 U12329 ( .A1(n14904), .A2(n15017), .ZN(n15265) );
  NAND2_X1 U12330 ( .A1(n14902), .A2(n10327), .ZN(n15463) );
  AND2_X1 U12331 ( .A1(n14902), .A2(n14901), .ZN(n15101) );
  NOR2_X1 U12332 ( .A1(n9855), .A2(n14172), .ZN(n14906) );
  AND2_X1 U12333 ( .A1(n10111), .A2(n15504), .ZN(n15287) );
  OAI21_X1 U12334 ( .B1(n15213), .B2(n10106), .A(n10104), .ZN(n10111) );
  AOI21_X1 U12335 ( .B1(n10109), .B2(n10107), .A(n10105), .ZN(n10104) );
  INV_X1 U12336 ( .A(n10107), .ZN(n10106) );
  AND2_X1 U12337 ( .A1(n15273), .A2(n10902), .ZN(n15286) );
  INV_X1 U12338 ( .A(n15559), .ZN(n11345) );
  AND2_X1 U12339 ( .A1(n11147), .A2(n10208), .ZN(n15305) );
  NAND2_X1 U12340 ( .A1(n9831), .A2(n10875), .ZN(n10191) );
  NAND2_X1 U12341 ( .A1(n10363), .A2(n10360), .ZN(n15571) );
  NOR2_X1 U12342 ( .A1(n16321), .A2(n10361), .ZN(n10360) );
  INV_X1 U12343 ( .A(n10362), .ZN(n10361) );
  AND3_X1 U12344 ( .A1(n11145), .A2(n11144), .A3(n11143), .ZN(n16326) );
  AND2_X1 U12345 ( .A1(n9870), .A2(n13978), .ZN(n10206) );
  NAND2_X1 U12346 ( .A1(n16354), .A2(n9853), .ZN(n10130) );
  AND2_X1 U12347 ( .A1(n14246), .A2(n11374), .ZN(n11262) );
  OR2_X1 U12348 ( .A1(n11063), .A2(n15629), .ZN(n15314) );
  OAI21_X1 U12349 ( .B1(n14072), .B2(n10811), .A(n10810), .ZN(n14103) );
  AND2_X1 U12350 ( .A1(n10214), .A2(n9942), .ZN(n14107) );
  AND2_X1 U12351 ( .A1(n14107), .A2(n14106), .ZN(n14109) );
  AND3_X1 U12352 ( .A1(n11253), .A2(n11252), .A3(n11251), .ZN(n14105) );
  INV_X1 U12353 ( .A(n11059), .ZN(n11060) );
  INV_X1 U12354 ( .A(n11058), .ZN(n11061) );
  OAI21_X1 U12355 ( .B1(n14076), .B2(n14246), .A(n14161), .ZN(n14072) );
  INV_X1 U12356 ( .A(n10598), .ZN(n10604) );
  NAND2_X1 U12357 ( .A1(n11224), .A2(n11223), .ZN(n13680) );
  AND2_X1 U12358 ( .A1(n11238), .A2(n11222), .ZN(n11223) );
  XNOR2_X1 U12359 ( .A(n11235), .B(n11236), .ZN(n13714) );
  NAND2_X1 U12360 ( .A1(n11217), .A2(n10357), .ZN(n11232) );
  XNOR2_X1 U12361 ( .A(n11243), .B(n11242), .ZN(n13727) );
  INV_X1 U12362 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15651) );
  OAI21_X1 U12363 ( .B1(n13088), .B2(n13087), .A(n13100), .ZN(n13746) );
  NAND2_X1 U12364 ( .A1(n11038), .A2(n10988), .ZN(n15641) );
  CLKBUF_X1 U12365 ( .A(n11020), .Z(n13674) );
  OR2_X1 U12367 ( .A1(n20021), .A2(n19426), .ZN(n19427) );
  INV_X1 U12368 ( .A(n19481), .ZN(n19484) );
  NAND2_X2 U12369 ( .A1(n10442), .A2(n10441), .ZN(n10502) );
  NAND4_X1 U12370 ( .A1(n9893), .A2(n10433), .A3(n10432), .A4(n10431), .ZN(
        n10442) );
  NOR2_X1 U12371 ( .A1(n19436), .A2(n19435), .ZN(n19480) );
  AND2_X1 U12372 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19965), .ZN(
        n13082) );
  NAND2_X1 U12373 ( .A1(n19611), .A2(n20152), .ZN(n19920) );
  INV_X1 U12374 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n16479) );
  NAND2_X1 U12375 ( .A1(n11674), .A2(n11701), .ZN(n11685) );
  OAI21_X1 U12376 ( .B1(n11698), .B2(n11708), .A(n11709), .ZN(n18777) );
  NOR2_X1 U12377 ( .A1(n16723), .A2(n16991), .ZN(n16714) );
  OR2_X1 U12378 ( .A1(n17023), .A2(n16670), .ZN(n16852) );
  NAND2_X1 U12379 ( .A1(n19008), .A2(n17516), .ZN(n16654) );
  NOR2_X1 U12380 ( .A1(n15708), .A2(n10005), .ZN(n15710) );
  INV_X1 U12381 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17153) );
  NOR2_X1 U12382 ( .A1(n17297), .A2(n10006), .ZN(n17299) );
  NAND2_X1 U12383 ( .A1(n10008), .A2(n10007), .ZN(n10006) );
  INV_X1 U12384 ( .A(n17298), .ZN(n10008) );
  INV_X1 U12385 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17317) );
  NOR2_X1 U12386 ( .A1(n18854), .A2(n16646), .ZN(n17515) );
  INV_X1 U12387 ( .A(n18775), .ZN(n17554) );
  NOR2_X1 U12388 ( .A1(n16692), .A2(n16657), .ZN(n16520) );
  NAND2_X1 U12389 ( .A1(n16526), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16657) );
  NAND2_X1 U12390 ( .A1(n17663), .A2(n10072), .ZN(n17626) );
  NOR2_X1 U12391 ( .A1(n10074), .A2(n10073), .ZN(n10072) );
  INV_X1 U12392 ( .A(n17662), .ZN(n10074) );
  NOR2_X1 U12393 ( .A1(n17684), .A2(n18031), .ZN(n17669) );
  INV_X1 U12394 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17685) );
  AND2_X1 U12395 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17949) );
  NAND2_X1 U12396 ( .A1(n17797), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10089) );
  OR2_X1 U12397 ( .A1(n17706), .A2(n18060), .ZN(n18018) );
  NOR2_X1 U12398 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17727), .ZN(
        n17705) );
  NOR2_X1 U12399 ( .A1(n18148), .A2(n11554), .ZN(n18122) );
  NAND2_X1 U12400 ( .A1(n10243), .A2(n17886), .ZN(n17781) );
  NAND2_X1 U12401 ( .A1(n17828), .A2(n10244), .ZN(n10243) );
  AND2_X1 U12402 ( .A1(n10245), .A2(n9984), .ZN(n10244) );
  NAND2_X1 U12403 ( .A1(n18122), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18099) );
  NOR2_X1 U12404 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10245) );
  NOR2_X1 U12405 ( .A1(n11742), .A2(n17893), .ZN(n17817) );
  NOR2_X1 U12406 ( .A1(n11701), .A2(n11669), .ZN(n18786) );
  NAND2_X1 U12407 ( .A1(n16646), .A2(n10019), .ZN(n11670) );
  AND2_X1 U12408 ( .A1(n11654), .A2(n18993), .ZN(n10019) );
  INV_X1 U12409 ( .A(n17817), .ZN(n18184) );
  AND2_X1 U12410 ( .A1(n11553), .A2(n10240), .ZN(n10239) );
  NOR2_X1 U12411 ( .A1(n17797), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10240) );
  NAND2_X1 U12412 ( .A1(n17921), .A2(n17922), .ZN(n17920) );
  XNOR2_X1 U12413 ( .A(n11544), .B(n11543), .ZN(n17929) );
  XNOR2_X1 U12414 ( .A(n11540), .B(n11539), .ZN(n17945) );
  NAND2_X1 U12415 ( .A1(n10086), .A2(n10085), .ZN(n17944) );
  NAND2_X1 U12416 ( .A1(n17954), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10085) );
  NAND2_X1 U12417 ( .A1(n17955), .A2(n10087), .ZN(n10086) );
  OR2_X1 U12418 ( .A1(n17954), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10087) );
  NAND2_X1 U12419 ( .A1(n17944), .A2(n17945), .ZN(n17943) );
  XNOR2_X1 U12420 ( .A(n11533), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17981) );
  NOR2_X2 U12421 ( .A1(n19007), .A2(n15770), .ZN(n18811) );
  NOR2_X1 U12422 ( .A1(n18972), .A2(n18809), .ZN(n18789) );
  NAND2_X1 U12423 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18809) );
  INV_X1 U12424 ( .A(n18811), .ZN(n18792) );
  NAND3_X1 U12425 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15775) );
  NAND2_X1 U12426 ( .A1(n10271), .A2(n10265), .ZN(n10264) );
  INV_X1 U12427 ( .A(n11663), .ZN(n18351) );
  INV_X1 U12428 ( .A(n11671), .ZN(n18360) );
  NAND2_X1 U12429 ( .A1(n18996), .A2(n18334), .ZN(n18486) );
  MUX2_X1 U12430 ( .A(n12989), .B(n12988), .S(n12987), .Z(n14418) );
  INV_X1 U12431 ( .A(n20292), .ZN(n20218) );
  INV_X1 U12432 ( .A(n20255), .ZN(n20288) );
  AND2_X1 U12433 ( .A1(n14549), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12897) );
  AND2_X1 U12434 ( .A1(n14408), .A2(n14031), .ZN(n20254) );
  INV_X1 U12435 ( .A(n15960), .ZN(n20245) );
  NOR2_X2 U12436 ( .A1(n12991), .A2(n12990), .ZN(n20272) );
  INV_X1 U12437 ( .A(n14029), .ZN(n12991) );
  INV_X1 U12438 ( .A(n20276), .ZN(n20285) );
  INV_X1 U12439 ( .A(n20272), .ZN(n20295) );
  AND2_X1 U12440 ( .A1(n14029), .A2(n13000), .ZN(n20292) );
  INV_X1 U12441 ( .A(n15974), .ZN(n20303) );
  AND2_X2 U12442 ( .A1(n13029), .A2(n13757), .ZN(n20306) );
  INV_X1 U12443 ( .A(n12880), .ZN(n10337) );
  INV_X1 U12444 ( .A(n14454), .ZN(n14505) );
  NAND2_X1 U12445 ( .A1(n13049), .A2(n13048), .ZN(n14527) );
  OR2_X1 U12446 ( .A1(n14532), .A2(n13806), .ZN(n14530) );
  AND2_X1 U12447 ( .A1(n13647), .A2(n13764), .ZN(n20310) );
  INV_X1 U12448 ( .A(n20308), .ZN(n20319) );
  INV_X1 U12449 ( .A(n13824), .ZN(n20351) );
  AND2_X1 U12450 ( .A1(n21069), .A2(n16146), .ZN(n13700) );
  OR2_X1 U12451 ( .A1(n20348), .A2(n11917), .ZN(n13824) );
  AOI21_X1 U12452 ( .B1(n10348), .B2(n14515), .A(n14514), .ZN(n16004) );
  INV_X1 U12453 ( .A(n14521), .ZN(n15932) );
  INV_X1 U12454 ( .A(n16038), .ZN(n16027) );
  OAI21_X1 U12455 ( .B1(n14548), .B2(n14547), .A(n14546), .ZN(n14690) );
  NAND2_X1 U12456 ( .A1(n10312), .A2(n10310), .ZN(n14546) );
  NAND2_X1 U12457 ( .A1(n14545), .A2(n14680), .ZN(n10312) );
  OAI21_X1 U12458 ( .B1(n14702), .B2(n20355), .A(n14701), .ZN(n14703) );
  AOI21_X1 U12459 ( .B1(n14734), .B2(n14700), .A(n14699), .ZN(n14701) );
  OR2_X1 U12460 ( .A1(n13033), .A2(n13032), .ZN(n13036) );
  XNOR2_X1 U12461 ( .A(n14597), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16047) );
  NAND2_X1 U12462 ( .A1(n10040), .A2(n14680), .ZN(n14621) );
  NAND2_X1 U12463 ( .A1(n14648), .A2(n9860), .ZN(n10040) );
  OAI21_X1 U12464 ( .B1(n13886), .B2(n16105), .A(n20361), .ZN(n16114) );
  NAND2_X1 U12465 ( .A1(n9825), .A2(n12699), .ZN(n14200) );
  NAND2_X1 U12466 ( .A1(n12681), .A2(n12680), .ZN(n14137) );
  AND2_X1 U12467 ( .A1(n13783), .A2(n15803), .ZN(n20366) );
  AND2_X1 U12468 ( .A1(n13783), .A2(n13770), .ZN(n20357) );
  NAND2_X1 U12469 ( .A1(n10299), .A2(n12073), .ZN(n10045) );
  NAND2_X1 U12470 ( .A1(n10047), .A2(n12072), .ZN(n10046) );
  NAND2_X1 U12471 ( .A1(n10048), .A2(n12073), .ZN(n10047) );
  INV_X1 U12472 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20791) );
  INV_X1 U12473 ( .A(n9885), .ZN(n12066) );
  INV_X1 U12474 ( .A(n12065), .ZN(n12067) );
  NAND2_X1 U12475 ( .A1(n13954), .A2(n20376), .ZN(n20763) );
  INV_X1 U12476 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20371) );
  OAI21_X1 U12477 ( .B1(n13947), .B2(n16151), .A(n20542), .ZN(n20370) );
  INV_X2 U12478 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13644) );
  AND2_X1 U12479 ( .A1(n12882), .A2(n11917), .ZN(n15803) );
  NOR2_X1 U12480 ( .A1(n13751), .A2(n20799), .ZN(n14834) );
  NOR2_X1 U12481 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14825) );
  OAI21_X1 U12482 ( .B1(n20559), .B2(n20543), .A(n20888), .ZN(n20561) );
  OR2_X1 U12483 ( .A1(n20629), .A2(n20880), .ZN(n20624) );
  OR2_X1 U12484 ( .A1(n20629), .A2(n20851), .ZN(n20622) );
  OAI211_X1 U12485 ( .C1(n20684), .C2(n20799), .A(n20721), .B(n20668), .ZN(
        n20686) );
  OR2_X1 U12486 ( .A1(n20763), .A2(n20851), .ZN(n20739) );
  INV_X1 U12487 ( .A(n20739), .ZN(n20746) );
  AOI22_X1 U12488 ( .A1(n20797), .A2(n20794), .B1(n20790), .B2(n20789), .ZN(
        n20842) );
  OAI211_X1 U12489 ( .C1(n20913), .C2(n20889), .A(n20888), .B(n20887), .ZN(
        n20915) );
  INV_X1 U12490 ( .A(n20792), .ZN(n20924) );
  INV_X1 U12491 ( .A(n20804), .ZN(n20940) );
  INV_X1 U12492 ( .A(n20809), .ZN(n20946) );
  INV_X1 U12493 ( .A(n20814), .ZN(n20952) );
  INV_X1 U12494 ( .A(n20819), .ZN(n20958) );
  OR2_X1 U12495 ( .A1(n20925), .A2(n20880), .ZN(n20969) );
  INV_X1 U12496 ( .A(n20986), .ZN(n20966) );
  INV_X1 U12497 ( .A(n20824), .ZN(n20964) );
  INV_X1 U12498 ( .A(n20829), .ZN(n20972) );
  OR2_X1 U12499 ( .A1(n20925), .A2(n20762), .ZN(n20986) );
  INV_X1 U12500 ( .A(n20835), .ZN(n20980) );
  INV_X1 U12501 ( .A(n14834), .ZN(n15835) );
  INV_X2 U12502 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20991) );
  INV_X1 U12503 ( .A(n13648), .ZN(n20989) );
  INV_X1 U12504 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20799) );
  NAND2_X1 U12505 ( .A1(n13438), .A2(n13437), .ZN(n14150) );
  CLKBUF_X1 U12506 ( .A(n11014), .Z(n11015) );
  NOR2_X1 U12507 ( .A1(n10167), .A2(n9964), .ZN(n10164) );
  INV_X1 U12508 ( .A(n10169), .ZN(n10167) );
  AND2_X1 U12509 ( .A1(n16152), .A2(n10171), .ZN(n10165) );
  INV_X1 U12510 ( .A(n10170), .ZN(n10166) );
  NAND2_X1 U12511 ( .A1(n16180), .A2(n16181), .ZN(n16179) );
  NAND2_X1 U12512 ( .A1(n16206), .A2(n19182), .ZN(n16193) );
  NAND2_X1 U12513 ( .A1(n16215), .A2(n19182), .ZN(n16207) );
  NAND2_X1 U12514 ( .A1(n16207), .A2(n16208), .ZN(n16206) );
  NAND2_X1 U12515 ( .A1(n16228), .A2(n19182), .ZN(n16216) );
  NAND2_X1 U12516 ( .A1(n16216), .A2(n16217), .ZN(n16215) );
  NAND2_X1 U12517 ( .A1(n16155), .A2(n19182), .ZN(n16255) );
  NAND2_X1 U12518 ( .A1(n15795), .A2(n15796), .ZN(n16155) );
  INV_X1 U12519 ( .A(n19239), .ZN(n19207) );
  NAND2_X1 U12520 ( .A1(n19014), .A2(n14160), .ZN(n19204) );
  CLKBUF_X1 U12521 ( .A(n14153), .Z(n19198) );
  INV_X1 U12522 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n19233) );
  NAND2_X1 U12523 ( .A1(n9902), .A2(n13337), .ZN(n10283) );
  NAND2_X1 U12524 ( .A1(n14963), .A2(n14964), .ZN(n10280) );
  OR2_X1 U12525 ( .A1(n11373), .A2(n11372), .ZN(n19263) );
  OR2_X1 U12526 ( .A1(n11358), .A2(n11357), .ZN(n19264) );
  NAND2_X1 U12527 ( .A1(n10287), .A2(n19269), .ZN(n10286) );
  INV_X1 U12528 ( .A(n10288), .ZN(n10287) );
  OR2_X1 U12529 ( .A1(n11327), .A2(n11326), .ZN(n14004) );
  OR2_X1 U12530 ( .A1(n11312), .A2(n11311), .ZN(n19276) );
  INV_X1 U12531 ( .A(n19289), .ZN(n19278) );
  NAND2_X1 U12532 ( .A1(n19293), .A2(n11217), .ZN(n19289) );
  NOR2_X1 U12533 ( .A1(n14973), .A2(n14972), .ZN(n14971) );
  NAND2_X1 U12534 ( .A1(n13337), .A2(n13339), .ZN(n14973) );
  AND2_X1 U12535 ( .A1(n13678), .A2(n13520), .ZN(n19300) );
  AND2_X1 U12536 ( .A1(n13678), .A2(n19436), .ZN(n19299) );
  AND2_X1 U12537 ( .A1(n19347), .A2(n13406), .ZN(n19298) );
  AND2_X1 U12538 ( .A1(n19361), .A2(n19348), .ZN(n19338) );
  INV_X1 U12539 ( .A(n19361), .ZN(n19342) );
  INV_X1 U12540 ( .A(n19348), .ZN(n19357) );
  INV_X1 U12541 ( .A(n19325), .ZN(n19365) );
  OR2_X1 U12542 ( .A1(n19298), .A2(n13678), .ZN(n19325) );
  OR2_X1 U12543 ( .A1(n14150), .A2(n19447), .ZN(n14152) );
  INV_X1 U12544 ( .A(n15330), .ZN(n16169) );
  INV_X1 U12545 ( .A(n19425), .ZN(n16316) );
  INV_X1 U12546 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16351) );
  INV_X1 U12547 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19424) );
  INV_X1 U12548 ( .A(n16363), .ZN(n19416) );
  XNOR2_X1 U12549 ( .A(n14235), .B(n10375), .ZN(n15131) );
  INV_X1 U12550 ( .A(n15157), .ZN(n16214) );
  CLKBUF_X1 U12551 ( .A(n15176), .Z(n15177) );
  INV_X1 U12552 ( .A(n15386), .ZN(n16262) );
  NAND2_X1 U12553 ( .A1(n15220), .A2(n9883), .ZN(n15419) );
  XNOR2_X1 U12554 ( .A(n10101), .B(n15219), .ZN(n15434) );
  NAND2_X1 U12555 ( .A1(n10102), .A2(n15232), .ZN(n10101) );
  NAND2_X1 U12556 ( .A1(n15234), .A2(n15218), .ZN(n10102) );
  INV_X1 U12557 ( .A(n10135), .ZN(n15502) );
  OAI21_X1 U12558 ( .B1(n15479), .B2(n9960), .A(n10136), .ZN(n10135) );
  NOR2_X1 U12559 ( .A1(n15509), .A2(n10137), .ZN(n10136) );
  NAND2_X1 U12560 ( .A1(n15287), .A2(n15286), .ZN(n15498) );
  NAND2_X1 U12561 ( .A1(n10103), .A2(n10107), .ZN(n15506) );
  NAND2_X1 U12562 ( .A1(n15213), .A2(n10108), .ZN(n10103) );
  NAND2_X1 U12563 ( .A1(n15213), .A2(n15291), .ZN(n15536) );
  AND2_X1 U12564 ( .A1(n15303), .A2(n14007), .ZN(n19135) );
  INV_X1 U12565 ( .A(n15406), .ZN(n15597) );
  INV_X1 U12566 ( .A(n16425), .ZN(n16407) );
  INV_X1 U12567 ( .A(n16412), .ZN(n16387) );
  CLKBUF_X1 U12568 ( .A(n9833), .Z(n13821) );
  INV_X1 U12569 ( .A(n16416), .ZN(n16390) );
  INV_X1 U12570 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20165) );
  NAND2_X1 U12571 ( .A1(n15643), .A2(n13556), .ZN(n20160) );
  INV_X1 U12572 ( .A(n20122), .ZN(n20132) );
  INV_X1 U12573 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16463) );
  XNOR2_X1 U12574 ( .A(n13589), .B(n13591), .ZN(n20130) );
  OAI21_X1 U12575 ( .B1(n13817), .B2(n13818), .A(n13819), .ZN(n20122) );
  INV_X1 U12576 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13676) );
  AOI21_X1 U12577 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16490), .A(n13670), .ZN(
        n20123) );
  INV_X1 U12578 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19462) );
  INV_X1 U12579 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n19468) );
  INV_X1 U12580 ( .A(n19544), .ZN(n19528) );
  OR2_X1 U12581 ( .A1(n19554), .A2(n19673), .ZN(n19573) );
  INV_X1 U12582 ( .A(n19563), .ZN(n19572) );
  NOR2_X1 U12583 ( .A1(n19709), .A2(n20127), .ZN(n19628) );
  NOR2_X1 U12584 ( .A1(n19613), .A2(n19610), .ZN(n19634) );
  INV_X1 U12585 ( .A(n19676), .ZN(n19694) );
  OR2_X1 U12586 ( .A1(n19704), .A2(n19703), .ZN(n19729) );
  INV_X1 U12587 ( .A(n19758), .ZN(n19750) );
  NOR2_X1 U12588 ( .A1(n19899), .A2(n19764), .ZN(n19823) );
  NOR2_X1 U12589 ( .A1(n19899), .A2(n20127), .ZN(n19865) );
  OAI22_X1 U12590 ( .A1(n19463), .A2(n19482), .B1(n20420), .B2(n19484), .ZN(
        n19947) );
  OAI22_X1 U12591 ( .A1(n19469), .A2(n19482), .B1(n20427), .B2(n19484), .ZN(
        n19950) );
  OAI21_X1 U12592 ( .B1(n19933), .B2(n19932), .A(n19931), .ZN(n19960) );
  OAI22_X1 U12593 ( .A1(n13065), .A2(n19484), .B1(n19483), .B2(n19482), .ZN(
        n19958) );
  AND2_X1 U12594 ( .A1(n19447), .A2(n19485), .ZN(n19980) );
  INV_X1 U12595 ( .A(n19782), .ZN(n19994) );
  AND2_X1 U12596 ( .A1(n19458), .A2(n19485), .ZN(n19992) );
  INV_X1 U12597 ( .A(n19523), .ZN(n19998) );
  INV_X1 U12598 ( .A(n19817), .ZN(n20006) );
  INV_X1 U12599 ( .A(n19950), .ZN(n20009) );
  INV_X1 U12600 ( .A(n19820), .ZN(n20012) );
  INV_X1 U12601 ( .A(n19954), .ZN(n20015) );
  AND2_X1 U12602 ( .A1(n13082), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20017) );
  NOR2_X2 U12603 ( .A1(n19899), .A2(n19920), .ZN(n20021) );
  AND2_X1 U12604 ( .A1(n19485), .A2(n11217), .ZN(n20016) );
  INV_X1 U12605 ( .A(n19964), .ZN(n20025) );
  OR2_X1 U12606 ( .A1(n15864), .A2(n20158), .ZN(n16488) );
  INV_X1 U12607 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20158) );
  INV_X1 U12608 ( .A(n16650), .ZN(n19008) );
  INV_X1 U12609 ( .A(n10075), .ZN(n16724) );
  NOR2_X1 U12610 ( .A1(n16769), .A2(n16669), .ZN(n16750) );
  INV_X1 U12611 ( .A(n10077), .ZN(n16768) );
  NOR2_X1 U12612 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16801), .ZN(n16786) );
  NOR2_X1 U12613 ( .A1(n18898), .A2(n16816), .ZN(n16800) );
  NOR2_X1 U12614 ( .A1(n18891), .A2(n16852), .ZN(n16845) );
  INV_X1 U12615 ( .A(n16949), .ZN(n16959) );
  NOR2_X1 U12616 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16893), .ZN(n16876) );
  NOR2_X1 U12617 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16965), .ZN(n16946) );
  NOR2_X1 U12618 ( .A1(n18774), .A2(n16654), .ZN(n17009) );
  INV_X1 U12619 ( .A(n16969), .ZN(n17018) );
  INV_X1 U12620 ( .A(n17026), .ZN(n17030) );
  INV_X1 U12621 ( .A(n16766), .ZN(n17032) );
  NOR2_X1 U12622 ( .A1(n10260), .A2(n17361), .ZN(n17083) );
  NAND2_X1 U12623 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17096), .ZN(n17088) );
  AND2_X1 U12624 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n17100), .ZN(n17096) );
  NOR2_X1 U12625 ( .A1(n17040), .A2(n17097), .ZN(n17100) );
  NOR2_X1 U12626 ( .A1(n17038), .A2(n17120), .ZN(n17101) );
  NOR2_X1 U12627 ( .A1(n17167), .A2(n9965), .ZN(n17135) );
  INV_X1 U12628 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n10261) );
  INV_X1 U12629 ( .A(n17229), .ZN(n17213) );
  NAND2_X1 U12630 ( .A1(n17247), .A2(P3_EBX_REG_12__SCAN_IN), .ZN(n15757) );
  NAND2_X1 U12631 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17267), .ZN(n17249) );
  AND2_X1 U12632 ( .A1(n17306), .A2(P3_EBX_REG_9__SCAN_IN), .ZN(n17267) );
  NOR2_X1 U12633 ( .A1(n17360), .A2(n17342), .ZN(n17337) );
  INV_X1 U12634 ( .A(n17376), .ZN(n17372) );
  NOR2_X1 U12635 ( .A1(n17581), .A2(n17385), .ZN(n17381) );
  INV_X1 U12636 ( .A(n17399), .ZN(n17395) );
  NAND2_X1 U12637 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17395), .ZN(n17394) );
  NOR2_X1 U12638 ( .A1(n17409), .A2(n17404), .ZN(n17400) );
  NOR2_X1 U12639 ( .A1(n17560), .A2(n17437), .ZN(n17431) );
  NOR2_X1 U12640 ( .A1(n17620), .A2(n17455), .ZN(n17448) );
  INV_X1 U12641 ( .A(n17473), .ZN(n17477) );
  AOI211_X1 U12642 ( .C1(n11497), .C2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n11517), .B(n11516), .ZN(n17487) );
  AND2_X1 U12643 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17492), .ZN(n17489) );
  INV_X1 U12644 ( .A(n11719), .ZN(n17490) );
  NOR2_X1 U12645 ( .A1(n17453), .A2(n17493), .ZN(n17492) );
  AOI211_X1 U12646 ( .C1(n17200), .C2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n11506), .B(n11505), .ZN(n17495) );
  OR2_X1 U12647 ( .A1(n11482), .A2(n11481), .ZN(n11483) );
  OR3_X1 U12648 ( .A1(n11478), .A2(n11477), .A3(n11476), .ZN(n11484) );
  AND2_X1 U12649 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11481) );
  NOR3_X1 U12650 ( .A1(n17591), .A2(n17510), .A3(n17501), .ZN(n17506) );
  INV_X1 U12651 ( .A(n17509), .ZN(n17507) );
  AOI21_X2 U12652 ( .B1(n15870), .B2(n15869), .A(n18828), .ZN(n17514) );
  NOR2_X1 U12653 ( .A1(n18796), .A2(n17494), .ZN(n17509) );
  INV_X1 U12654 ( .A(n17504), .ZN(n17508) );
  CLKBUF_X1 U12655 ( .A(n17617), .Z(n17604) );
  OAI211_X1 U12656 ( .C1(n18339), .C2(n18988), .A(n17554), .B(n17553), .ZN(
        n17617) );
  INV_X1 U12657 ( .A(n16499), .ZN(n16501) );
  AND2_X1 U12658 ( .A1(n18308), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n10012) );
  INV_X1 U12659 ( .A(n10014), .ZN(n17760) );
  NAND2_X1 U12660 ( .A1(n17786), .A2(n9935), .ZN(n17770) );
  INV_X1 U12661 ( .A(n17895), .ZN(n17860) );
  INV_X1 U12662 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17903) );
  INV_X1 U12663 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17930) );
  INV_X1 U12664 ( .A(n18463), .ZN(n18719) );
  INV_X1 U12665 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18015) );
  NOR2_X1 U12666 ( .A1(n10246), .A2(n9805), .ZN(n17680) );
  INV_X1 U12667 ( .A(n10248), .ZN(n10246) );
  NAND2_X1 U12668 ( .A1(n17828), .A2(n18152), .ZN(n17818) );
  NAND2_X1 U12669 ( .A1(n17955), .A2(n17954), .ZN(n17953) );
  INV_X1 U12670 ( .A(n18310), .ZN(n18294) );
  INV_X1 U12671 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18801) );
  INV_X1 U12672 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18330) );
  INV_X1 U12673 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18328) );
  INV_X1 U12674 ( .A(n18828), .ZN(n18991) );
  NOR2_X1 U12675 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18996), .ZN(n18839) );
  INV_X1 U12676 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18996) );
  INV_X1 U12677 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18862) );
  NAND2_X1 U12678 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18862), .ZN(n19003) );
  AND2_X2 U12679 ( .A1(n13061), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20373)
         );
  INV_X1 U12680 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21375) );
  CLKBUF_X1 U12681 ( .A(n16618), .Z(n16617) );
  OAI21_X1 U12682 ( .B1(n14755), .B2(n20187), .A(n10051), .ZN(P1_U2972) );
  INV_X1 U12683 ( .A(n12787), .ZN(n10052) );
  OAI21_X1 U12684 ( .B1(n16047), .B2(n20187), .A(n10145), .ZN(P1_U2974) );
  INV_X1 U12685 ( .A(n10146), .ZN(n10145) );
  OAI21_X1 U12686 ( .B1(n14600), .B2(n14689), .A(n10147), .ZN(n10146) );
  AOI21_X1 U12687 ( .B1(n16033), .B2(n14599), .A(n14598), .ZN(n10147) );
  NAND2_X1 U12688 ( .A1(n10168), .A2(n10170), .ZN(n16170) );
  AOI211_X1 U12689 ( .C1(n16363), .C2(n16260), .A(n14279), .B(n14278), .ZN(
        n14280) );
  NAND2_X1 U12690 ( .A1(n15435), .A2(n16366), .ZN(n15243) );
  OAI211_X1 U12691 ( .C1(n16413), .C2(n15330), .A(n15329), .B(n10372), .ZN(
        n15331) );
  OAI21_X1 U12692 ( .B1(n16689), .B2(n10070), .A(n10067), .ZN(P3_U2642) );
  AND2_X1 U12693 ( .A1(n16697), .A2(n10068), .ZN(n10067) );
  INV_X1 U12694 ( .A(n10071), .ZN(n10070) );
  OAI21_X1 U12695 ( .B1(n10259), .B2(n17082), .A(n10257), .ZN(P3_U2674) );
  AOI21_X1 U12696 ( .B1(n10260), .B2(n17082), .A(n10258), .ZN(n10257) );
  INV_X1 U12697 ( .A(n17083), .ZN(n10259) );
  NOR2_X1 U12698 ( .A1(n17358), .A2(n17379), .ZN(n10258) );
  NOR3_X1 U12699 ( .A1(n17167), .A2(n17409), .A3(n16802), .ZN(n17149) );
  INV_X1 U12700 ( .A(n17306), .ZN(n17326) );
  AOI211_X1 U12701 ( .C1(n10014), .C2(n10013), .A(n17750), .B(n10012), .ZN(
        n17755) );
  AOI22_X1 U12702 ( .A1(n17749), .A2(n17759), .B1(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10013) );
  AOI21_X1 U12703 ( .B1(n10079), .B2(n10082), .A(n10078), .ZN(n11754) );
  OAI21_X1 U12704 ( .B1(n16502), .B2(n18304), .A(n11751), .ZN(n11752) );
  OAI21_X1 U12705 ( .B1(n10253), .B2(n10252), .A(n9865), .ZN(P3_U2834) );
  OR2_X1 U12706 ( .A1(n9822), .A2(n15781), .ZN(n10252) );
  AOI211_X1 U12707 ( .C1(n13015), .C2(n13014), .A(n10254), .B(n13013), .ZN(
        n10253) );
  NAND4_X2 U12708 ( .A1(n18964), .A2(n10256), .A3(n11435), .A4(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11467) );
  OR3_X2 U12709 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n18807), .ZN(n9856) );
  OR3_X1 U12710 ( .A1(n17021), .A2(n10256), .A3(n11435), .ZN(n11479) );
  AND2_X1 U12711 ( .A1(n11077), .A2(n10306), .ZN(n9853) );
  NAND2_X1 U12712 ( .A1(n10354), .A2(n10379), .ZN(n14170) );
  NAND2_X1 U12713 ( .A1(n10373), .A2(n10928), .ZN(n9854) );
  OR2_X1 U12714 ( .A1(n14097), .A2(n15523), .ZN(n9855) );
  OR2_X1 U12715 ( .A1(n15265), .A2(n10200), .ZN(n9857) );
  AND2_X1 U12716 ( .A1(n14359), .A2(n10345), .ZN(n14337) );
  NAND2_X1 U12717 ( .A1(n12360), .A2(n9953), .ZN(n14395) );
  AND2_X1 U12718 ( .A1(n11131), .A2(n10207), .ZN(n9858) );
  AND2_X1 U12719 ( .A1(n14522), .A2(n10350), .ZN(n14442) );
  AND2_X1 U12720 ( .A1(n10540), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9859) );
  AND2_X1 U12721 ( .A1(n14647), .A2(n9992), .ZN(n9860) );
  AND2_X1 U12722 ( .A1(n10359), .A2(n9927), .ZN(n9861) );
  INV_X1 U12723 ( .A(n12072), .ZN(n10299) );
  NAND2_X1 U12724 ( .A1(n14522), .A2(n14523), .ZN(n14440) );
  NOR3_X1 U12725 ( .A1(n14240), .A2(n10858), .A3(n15325), .ZN(n9862) );
  NAND2_X1 U12726 ( .A1(n14359), .A2(n9928), .ZN(n14323) );
  NOR2_X1 U12727 ( .A1(n14992), .A2(n14993), .ZN(n9863) );
  INV_X1 U12728 ( .A(n10880), .ZN(n10189) );
  NOR2_X1 U12729 ( .A1(n10189), .A2(n10187), .ZN(n9864) );
  AND3_X1 U12730 ( .A1(n9919), .A2(n10251), .A3(n10250), .ZN(n9865) );
  NAND2_X1 U12731 ( .A1(n10444), .A2(n10371), .ZN(n9866) );
  AND2_X1 U12732 ( .A1(n10099), .A2(n10098), .ZN(n9867) );
  AND2_X1 U12733 ( .A1(n11079), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9868) );
  AND2_X1 U12734 ( .A1(n15650), .A2(n9918), .ZN(n9869) );
  AND2_X1 U12735 ( .A1(n9858), .A2(n14920), .ZN(n9870) );
  OR2_X1 U12736 ( .A1(n10398), .A2(n10096), .ZN(n9871) );
  NAND2_X1 U12737 ( .A1(n14997), .A2(n9959), .ZN(n14958) );
  AND3_X1 U12738 ( .A1(n10962), .A2(n10956), .A3(n9948), .ZN(n9872) );
  NOR3_X1 U12739 ( .A1(n11442), .A2(n11441), .A3(n9932), .ZN(n9873) );
  AND2_X1 U12740 ( .A1(n10219), .A2(n9962), .ZN(n9874) );
  INV_X2 U12741 ( .A(n12127), .ZN(n12038) );
  OR2_X1 U12742 ( .A1(n13974), .A2(n13108), .ZN(n13975) );
  NAND2_X1 U12743 ( .A1(n16401), .A2(n16400), .ZN(n14923) );
  NAND2_X1 U12744 ( .A1(n15013), .A2(n10293), .ZN(n15001) );
  NAND2_X1 U12745 ( .A1(n11031), .A2(n10516), .ZN(n9875) );
  INV_X1 U12746 ( .A(n19182), .ZN(n19192) );
  INV_X1 U12747 ( .A(n15199), .ZN(n10367) );
  AND2_X1 U12748 ( .A1(n10174), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9876) );
  AND2_X1 U12749 ( .A1(n10156), .A2(n9981), .ZN(n9877) );
  AND2_X1 U12750 ( .A1(n10150), .A2(n14403), .ZN(n9878) );
  AND2_X1 U12751 ( .A1(n10326), .A2(n10327), .ZN(n9879) );
  INV_X1 U12752 ( .A(n16171), .ZN(n10171) );
  AND2_X1 U12753 ( .A1(n11132), .A2(n9858), .ZN(n9880) );
  AND2_X1 U12754 ( .A1(n9961), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9881) );
  AND2_X1 U12755 ( .A1(n10149), .A2(n10148), .ZN(n9882) );
  AND2_X1 U12756 ( .A1(n15397), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9883) );
  AND3_X1 U12757 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .A3(P3_EBX_REG_12__SCAN_IN), .ZN(n9884) );
  OR2_X1 U12758 ( .A1(n10648), .A2(n10647), .ZN(n11221) );
  AND2_X2 U12759 ( .A1(n13312), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10748) );
  AND2_X1 U12760 ( .A1(n9840), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10694) );
  AND2_X1 U12761 ( .A1(n10142), .A2(n12051), .ZN(n9885) );
  NOR2_X2 U12762 ( .A1(n11434), .A2(n11432), .ZN(n11519) );
  OR2_X1 U12763 ( .A1(n10935), .A2(n10231), .ZN(n9886) );
  OR2_X1 U12764 ( .A1(n11435), .A2(n11436), .ZN(n9887) );
  INV_X2 U12765 ( .A(n11448), .ZN(n17293) );
  OR2_X1 U12766 ( .A1(n17021), .A2(n11434), .ZN(n9888) );
  NAND2_X1 U12767 ( .A1(n14359), .A2(n10376), .ZN(n14347) );
  NAND2_X1 U12768 ( .A1(n10092), .A2(n10847), .ZN(n11063) );
  AND2_X1 U12769 ( .A1(n10882), .A2(n10221), .ZN(n9889) );
  AND4_X1 U12770 ( .A1(n10682), .A2(n10681), .A3(n10680), .A4(n10679), .ZN(
        n9891) );
  NAND2_X1 U12771 ( .A1(n10277), .A2(n10276), .ZN(n14953) );
  AND2_X1 U12772 ( .A1(n12360), .A2(n10335), .ZN(n14394) );
  NAND2_X1 U12773 ( .A1(n12360), .A2(n12359), .ZN(n14438) );
  INV_X2 U12774 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10444) );
  OR3_X1 U12775 ( .A1(n12817), .A2(n10337), .A3(n10338), .ZN(n9892) );
  AND2_X1 U12776 ( .A1(n10430), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9893) );
  NAND2_X2 U12777 ( .A1(n10131), .A2(n10130), .ZN(n15220) );
  NAND2_X1 U12778 ( .A1(n13101), .A2(n13100), .ZN(n13818) );
  XNOR2_X1 U12779 ( .A(n13307), .B(n13308), .ZN(n14976) );
  OR3_X1 U12780 ( .A1(n10935), .A2(n10934), .A3(n10232), .ZN(n9894) );
  AND2_X1 U12781 ( .A1(n10705), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n9895) );
  OAI21_X1 U12782 ( .B1(n11063), .B2(n14246), .A(n19189), .ZN(n10814) );
  AND3_X1 U12783 ( .A1(n11226), .A2(n20136), .A3(n10314), .ZN(n9896) );
  INV_X1 U12784 ( .A(n10144), .ZN(n14608) );
  AND2_X1 U12785 ( .A1(n10215), .A2(n15132), .ZN(n9897) );
  INV_X1 U12786 ( .A(n16019), .ZN(n10119) );
  NAND2_X1 U12787 ( .A1(n10359), .A2(n10362), .ZN(n16317) );
  AND2_X1 U12788 ( .A1(n10368), .A2(n10367), .ZN(n9898) );
  OAI22_X1 U12789 ( .A1(n9835), .A2(n10397), .B1(n13242), .B2(n19468), .ZN(
        n10398) );
  AND3_X1 U12790 ( .A1(n10452), .A2(n10451), .A3(n10450), .ZN(n9899) );
  AND2_X1 U12791 ( .A1(n10882), .A2(n9874), .ZN(n10897) );
  AND2_X1 U12792 ( .A1(n10132), .A2(n9853), .ZN(n9900) );
  AND2_X1 U12793 ( .A1(n10402), .A2(n10444), .ZN(n9901) );
  AND2_X1 U12794 ( .A1(n13339), .A2(n10284), .ZN(n9902) );
  AND2_X1 U12795 ( .A1(n10082), .A2(n10233), .ZN(n9903) );
  AND2_X1 U12796 ( .A1(n12073), .A2(n10298), .ZN(n9904) );
  AND2_X1 U12797 ( .A1(n10639), .A2(n10198), .ZN(n9905) );
  NOR2_X1 U12798 ( .A1(n10188), .A2(n10187), .ZN(n9906) );
  NOR2_X1 U12799 ( .A1(n10396), .A2(n10395), .ZN(n10503) );
  AND2_X1 U12800 ( .A1(n15053), .A2(n15048), .ZN(n15037) );
  NAND2_X1 U12801 ( .A1(n14272), .A2(n14271), .ZN(n9907) );
  NAND2_X1 U12802 ( .A1(n15220), .A2(n10308), .ZN(n15172) );
  INV_X1 U12803 ( .A(n15172), .ZN(n11081) );
  AND2_X1 U12804 ( .A1(n15220), .A2(n10309), .ZN(n9908) );
  AND2_X1 U12805 ( .A1(n14359), .A2(n10343), .ZN(n12627) );
  AND2_X1 U12806 ( .A1(n15220), .A2(n15397), .ZN(n9909) );
  AND2_X1 U12808 ( .A1(n11444), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n9910) );
  OR2_X1 U12809 ( .A1(n14680), .A2(n16126), .ZN(n9911) );
  OR2_X1 U12810 ( .A1(n11235), .A2(n11236), .ZN(n9912) );
  AND3_X1 U12811 ( .A1(n10510), .A2(n10502), .A3(n10509), .ZN(n9913) );
  AND2_X1 U12812 ( .A1(n10097), .A2(n10402), .ZN(n9914) );
  AND2_X1 U12813 ( .A1(n10113), .A2(n12721), .ZN(n9915) );
  OR2_X1 U12814 ( .A1(n17312), .A2(n17359), .ZN(n9916) );
  NOR2_X1 U12815 ( .A1(n11502), .A2(n10004), .ZN(n9917) );
  AND2_X1 U12816 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n9918) );
  NAND3_X1 U12817 ( .A1(n17624), .A2(n17640), .A3(n18219), .ZN(n9919) );
  OAI21_X1 U12818 ( .B1(n16505), .B2(n18185), .A(n10084), .ZN(n10083) );
  INV_X1 U12819 ( .A(n10307), .ZN(n10133) );
  NOR2_X1 U12820 ( .A1(n16352), .A2(n11076), .ZN(n10307) );
  AND2_X1 U12821 ( .A1(n10849), .A2(n10855), .ZN(n9920) );
  INV_X1 U12822 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11435) );
  INV_X1 U12823 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18964) );
  INV_X1 U12824 ( .A(n10588), .ZN(n14259) );
  INV_X2 U12825 ( .A(n14259), .ZN(n14250) );
  INV_X1 U12826 ( .A(n10574), .ZN(n11113) );
  INV_X1 U12827 ( .A(n12190), .ZN(n12263) );
  INV_X1 U12828 ( .A(n12263), .ZN(n12879) );
  NOR2_X1 U12829 ( .A1(n15557), .A2(n11345), .ZN(n15539) );
  AND2_X1 U12830 ( .A1(n14997), .A2(n14987), .ZN(n14979) );
  AND2_X1 U12831 ( .A1(n17853), .A2(n18193), .ZN(n17828) );
  NAND2_X1 U12832 ( .A1(n17828), .A2(n10245), .ZN(n17796) );
  AND2_X1 U12833 ( .A1(n14424), .A2(n9882), .ZN(n9921) );
  NOR2_X1 U12834 ( .A1(n15540), .A2(n15521), .ZN(n15507) );
  NOR2_X1 U12835 ( .A1(n14119), .A2(n10355), .ZN(n14187) );
  NAND2_X1 U12836 ( .A1(n14874), .A2(n9876), .ZN(n14865) );
  NAND2_X1 U12837 ( .A1(n15412), .A2(n10332), .ZN(n15063) );
  INV_X1 U12838 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n16491) );
  AND2_X1 U12839 ( .A1(n10179), .A2(n10176), .ZN(n9922) );
  AND2_X1 U12840 ( .A1(n10324), .A2(n15598), .ZN(n9923) );
  INV_X1 U12841 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10020) );
  NOR2_X1 U12842 ( .A1(n14174), .A2(n19257), .ZN(n15014) );
  AND2_X1 U12843 ( .A1(n11254), .A2(n10527), .ZN(n9924) );
  AND2_X1 U12844 ( .A1(n14874), .A2(n10174), .ZN(n9925) );
  NAND2_X1 U12845 ( .A1(n13763), .A2(n20413), .ZN(n11916) );
  OR2_X1 U12846 ( .A1(n15265), .A2(n15264), .ZN(n9926) );
  AND2_X1 U12847 ( .A1(n16343), .A2(n16358), .ZN(n9927) );
  AND2_X1 U12848 ( .A1(n10345), .A2(n14338), .ZN(n9928) );
  AND2_X1 U12849 ( .A1(n11146), .A2(n10210), .ZN(n9929) );
  NAND2_X1 U12850 ( .A1(n10191), .A2(n10880), .ZN(n15299) );
  AND2_X1 U12851 ( .A1(n14906), .A2(n14905), .ZN(n14904) );
  AND2_X1 U12852 ( .A1(n15232), .A2(n15231), .ZN(n9930) );
  NOR2_X1 U12853 ( .A1(n15465), .A2(n15091), .ZN(n15090) );
  AND3_X1 U12854 ( .A1(n10223), .A2(n10795), .A3(n10849), .ZN(n9931) );
  AND2_X1 U12855 ( .A1(n10801), .A2(n10797), .ZN(n10795) );
  INV_X1 U12856 ( .A(n10531), .ZN(n11022) );
  OR2_X1 U12857 ( .A1(n12285), .A2(n12284), .ZN(n14448) );
  INV_X1 U12858 ( .A(n10100), .ZN(n11096) );
  NOR2_X1 U12859 ( .A1(n15073), .A2(n13241), .ZN(n14992) );
  AND2_X1 U12860 ( .A1(n11444), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n9932) );
  NOR2_X1 U12861 ( .A1(n14801), .A2(n14802), .ZN(n14424) );
  INV_X1 U12862 ( .A(n14119), .ZN(n10354) );
  AND2_X1 U12863 ( .A1(n10208), .A2(n14098), .ZN(n9933) );
  INV_X1 U12864 ( .A(n13887), .ZN(n12909) );
  OAI21_X1 U12865 ( .B1(n12665), .B2(n12172), .A(n12171), .ZN(n14040) );
  OR2_X1 U12866 ( .A1(n19038), .A2(n19042), .ZN(n9934) );
  AND2_X1 U12867 ( .A1(n15090), .A2(n15445), .ZN(n14854) );
  AND2_X1 U12868 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n9935) );
  XOR2_X1 U12869 ( .A(n14680), .B(n14737), .Z(n9936) );
  AND2_X1 U12870 ( .A1(n10925), .A2(n10924), .ZN(n15230) );
  INV_X1 U12871 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n19177) );
  NAND2_X1 U12872 ( .A1(n15013), .A2(n16273), .ZN(n9937) );
  NAND2_X1 U12873 ( .A1(n14362), .A2(n9968), .ZN(n10162) );
  AND2_X1 U12874 ( .A1(n10035), .A2(n10034), .ZN(n9938) );
  OR2_X1 U12875 ( .A1(n16494), .A2(n18780), .ZN(n9939) );
  NAND2_X1 U12876 ( .A1(n10223), .A2(n10795), .ZN(n10225) );
  OR2_X1 U12877 ( .A1(n17886), .A2(n17995), .ZN(n9940) );
  AND2_X1 U12878 ( .A1(n19276), .A2(n14004), .ZN(n9941) );
  INV_X1 U12879 ( .A(n10109), .ZN(n10108) );
  OR2_X1 U12880 ( .A1(n15214), .A2(n10110), .ZN(n10109) );
  AND2_X1 U12881 ( .A1(n14997), .A2(n10213), .ZN(n14968) );
  OR2_X1 U12882 ( .A1(n11118), .A2(n11117), .ZN(n9942) );
  INV_X1 U12883 ( .A(n11030), .ZN(n10516) );
  AND2_X1 U12884 ( .A1(n10227), .A2(n10226), .ZN(n9943) );
  AND2_X1 U12885 ( .A1(n10152), .A2(n14049), .ZN(n9944) );
  AND2_X1 U12886 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n15662), .ZN(n9945) );
  NAND2_X1 U12887 ( .A1(n19470), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n9946) );
  AND2_X1 U12888 ( .A1(n9923), .A2(n10323), .ZN(n9947) );
  NAND2_X1 U12889 ( .A1(n15135), .A2(n15148), .ZN(n9948) );
  INV_X1 U12890 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n19107) );
  NAND2_X1 U12891 ( .A1(n12135), .A2(n12134), .ZN(n12146) );
  INV_X1 U12892 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10053) );
  INV_X1 U12893 ( .A(n9802), .ZN(n10081) );
  INV_X1 U12894 ( .A(n11228), .ZN(n13420) );
  INV_X1 U12895 ( .A(n12058), .ZN(n12891) );
  INV_X1 U12896 ( .A(n12891), .ZN(n12843) );
  NOR2_X1 U12897 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12058) );
  INV_X1 U12898 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n16450) );
  NAND2_X1 U12899 ( .A1(n16401), .A2(n9923), .ZN(n15599) );
  NOR2_X1 U12900 ( .A1(n14085), .A2(n14105), .ZN(n14104) );
  AND2_X1 U12901 ( .A1(n14096), .A2(n13109), .ZN(n9949) );
  NAND2_X1 U12902 ( .A1(n17899), .A2(n10239), .ZN(n17869) );
  AND2_X1 U12903 ( .A1(n12910), .A2(n10154), .ZN(n9950) );
  NAND2_X1 U12904 ( .A1(n11147), .A2(n9933), .ZN(n14097) );
  AND2_X1 U12905 ( .A1(n17247), .A2(n9884), .ZN(n9951) );
  AND2_X1 U12906 ( .A1(n14195), .A2(n10156), .ZN(n9952) );
  AND2_X1 U12907 ( .A1(n14396), .A2(n10335), .ZN(n9953) );
  AND2_X1 U12908 ( .A1(n13264), .A2(n13263), .ZN(n9954) );
  NOR2_X1 U12909 ( .A1(n15168), .A2(n10183), .ZN(n15121) );
  AND2_X1 U12910 ( .A1(n19470), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n9955) );
  AND2_X1 U12911 ( .A1(n19470), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n9956) );
  AND2_X1 U12912 ( .A1(n10293), .A2(n10292), .ZN(n9957) );
  AND2_X1 U12913 ( .A1(n15938), .A2(n10150), .ZN(n9958) );
  AND2_X1 U12914 ( .A1(n10213), .A2(n14969), .ZN(n9959) );
  AND2_X1 U12915 ( .A1(n16416), .A2(n15480), .ZN(n9960) );
  AND2_X1 U12916 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n9961) );
  NAND2_X1 U12917 ( .A1(n19470), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n9962) );
  INV_X1 U12918 ( .A(n17409), .ZN(n18366) );
  OAI211_X2 U12919 ( .C1(n11638), .C2(n17222), .A(n11637), .B(n11636), .ZN(
        n17409) );
  AND2_X1 U12920 ( .A1(n11444), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n9963) );
  AND2_X1 U12921 ( .A1(n19182), .A2(n10165), .ZN(n9964) );
  OR3_X1 U12922 ( .A1(n17409), .A2(n16802), .A3(n10261), .ZN(n9965) );
  OR2_X1 U12923 ( .A1(n15168), .A2(n15158), .ZN(n9966) );
  AND2_X1 U12924 ( .A1(n11553), .A2(n10241), .ZN(n9967) );
  AND2_X1 U12925 ( .A1(n10159), .A2(n10158), .ZN(n9968) );
  NAND2_X1 U12926 ( .A1(n19283), .A2(n19282), .ZN(n9969) );
  OR2_X1 U12927 ( .A1(n13974), .A2(n10288), .ZN(n10289) );
  INV_X1 U12928 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10196) );
  INV_X1 U12929 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16249) );
  AND2_X1 U12930 ( .A1(n19182), .A2(n10171), .ZN(n9970) );
  AND2_X1 U12931 ( .A1(n11132), .A2(n9870), .ZN(n9971) );
  AND2_X1 U12932 ( .A1(n16401), .A2(n10324), .ZN(n9972) );
  INV_X1 U12933 ( .A(n10321), .ZN(n10320) );
  OR2_X1 U12934 ( .A1(n11419), .A2(n10322), .ZN(n10321) );
  AND2_X1 U12935 ( .A1(n9957), .A2(n13264), .ZN(n9973) );
  AND2_X1 U12936 ( .A1(n15896), .A2(n15897), .ZN(n9974) );
  AND2_X1 U12937 ( .A1(n17899), .A2(n9967), .ZN(n9975) );
  AND2_X1 U12938 ( .A1(n9953), .A2(n10334), .ZN(n9976) );
  AND2_X1 U12939 ( .A1(n9882), .A2(n14374), .ZN(n9977) );
  AND2_X1 U12940 ( .A1(n9881), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9978) );
  AND2_X1 U12941 ( .A1(n10320), .A2(n10318), .ZN(n9979) );
  OR2_X1 U12942 ( .A1(n10702), .A2(n10701), .ZN(n11250) );
  NOR2_X1 U12943 ( .A1(n11419), .A2(n10319), .ZN(n9980) );
  AOI21_X1 U12944 ( .B1(n19182), .B2(n16152), .A(n10171), .ZN(n10170) );
  INV_X1 U12945 ( .A(n13520), .ZN(n19436) );
  INV_X1 U12946 ( .A(n11474), .ZN(n11447) );
  INV_X1 U12947 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10241) );
  INV_X1 U12948 ( .A(n14523), .ZN(n10351) );
  INV_X1 U12949 ( .A(n14513), .ZN(n10348) );
  OR2_X1 U12950 ( .A1(n12929), .A2(n12928), .ZN(n9981) );
  OR2_X1 U12951 ( .A1(n18990), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n9982) );
  NAND2_X1 U12952 ( .A1(n12881), .A2(n11917), .ZN(n13040) );
  AND2_X2 U12953 ( .A1(n10053), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15650) );
  AND2_X1 U12954 ( .A1(n11444), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n9983) );
  INV_X1 U12955 ( .A(n10138), .ZN(n13921) );
  NAND2_X1 U12956 ( .A1(n13910), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10138) );
  AND2_X1 U12957 ( .A1(n17851), .A2(n11555), .ZN(n9984) );
  NOR3_X1 U12958 ( .A1(n15687), .A2(n15688), .A3(n9983), .ZN(n9985) );
  AND2_X1 U12959 ( .A1(n17310), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n9986) );
  NOR2_X1 U12960 ( .A1(n15717), .A2(n10009), .ZN(n9987) );
  AND2_X1 U12961 ( .A1(n9884), .A2(P3_EBX_REG_15__SCAN_IN), .ZN(n9988) );
  INV_X1 U12962 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n10036) );
  INV_X1 U12963 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n10033) );
  INV_X1 U12964 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n10025) );
  INV_X1 U12965 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n10028) );
  NAND2_X1 U12966 ( .A1(n15857), .A2(n14691), .ZN(n9989) );
  INV_X1 U12967 ( .A(n14153), .ZN(n20032) );
  AND2_X1 U12968 ( .A1(n11444), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n9990) );
  AND2_X1 U12969 ( .A1(n11444), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n9991) );
  NOR2_X1 U12970 ( .A1(n10305), .A2(n15148), .ZN(n10304) );
  AND2_X1 U12971 ( .A1(n14767), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9992) );
  OR2_X1 U12972 ( .A1(n10303), .A2(n14258), .ZN(n9993) );
  NOR3_X1 U12973 ( .A1(n17223), .A2(n17224), .A3(n9990), .ZN(n9994) );
  NOR3_X1 U12974 ( .A1(n17280), .A2(n17279), .A3(n9991), .ZN(n9995) );
  AND2_X1 U12975 ( .A1(n17310), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n9996) );
  NOR2_X1 U12976 ( .A1(n14542), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9997) );
  INV_X1 U12977 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10073) );
  INV_X1 U12978 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10181) );
  INV_X1 U12979 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10182) );
  INV_X1 U12980 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14936) );
  NOR2_X1 U12981 ( .A1(n19463), .A2(n18463), .ZN(n18743) );
  OR2_X1 U12982 ( .A1(n18486), .A2(n18627), .ZN(n18463) );
  NAND2_X1 U12983 ( .A1(n11444), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10007) );
  NAND2_X1 U12984 ( .A1(n11444), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n14225) );
  NAND2_X1 U12985 ( .A1(n11444), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n17189) );
  AOI21_X1 U12986 ( .B1(n11444), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A(
        n10002), .ZN(n17256) );
  AOI22_X1 U12987 ( .A1(n11444), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__5__SCAN_IN), .B2(n17293), .ZN(n17131) );
  AOI21_X1 U12988 ( .B1(n11444), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A(
        n10003), .ZN(n17201) );
  AOI21_X1 U12989 ( .B1(n11444), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n10001), .ZN(n17155) );
  AOI21_X1 U12990 ( .B1(n11444), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n10000), .ZN(n17171) );
  AOI21_X1 U12991 ( .B1(n11444), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n9996), .ZN(n17311) );
  AOI21_X1 U12992 ( .B1(n11444), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n9986), .ZN(n15737) );
  AOI21_X1 U12993 ( .B1(n11444), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n9999), .ZN(n17109) );
  AOI21_X1 U12994 ( .B1(n11444), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n9998), .ZN(n15725) );
  NAND2_X1 U12995 ( .A1(n11444), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n10010) );
  INV_X1 U12996 ( .A(n10304), .ZN(n10303) );
  NOR2_X2 U12997 ( .A1(n18347), .A2(n18365), .ZN(n18738) );
  NOR2_X1 U12998 ( .A1(n10264), .A2(n11645), .ZN(n18347) );
  NAND2_X2 U12999 ( .A1(n16632), .A2(n9982), .ZN(n17988) );
  OAI21_X2 U13000 ( .B1(n18776), .B2(n18782), .A(n9939), .ZN(n18783) );
  INV_X2 U13001 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18972) );
  NAND2_X1 U13002 ( .A1(n14016), .A2(n14015), .ZN(n10021) );
  NAND2_X1 U13003 ( .A1(n13984), .A2(n13983), .ZN(n10022) );
  CLKBUF_X1 U13004 ( .A(n12983), .Z(n10023) );
  OR2_X1 U13005 ( .A1(n13030), .A2(n10023), .ZN(n12982) );
  NAND2_X1 U13006 ( .A1(n12638), .A2(n10044), .ZN(n12650) );
  NAND2_X1 U13007 ( .A1(n13749), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10044) );
  NAND2_X1 U13008 ( .A1(n13692), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13694) );
  XNOR2_X2 U13009 ( .A(n11989), .B(n11988), .ZN(n12075) );
  OAI211_X2 U13010 ( .C1(n12681), .C2(n10050), .A(n14134), .B(n10049), .ZN(
        n14180) );
  INV_X2 U13011 ( .A(n14135), .ZN(n10050) );
  NAND2_X1 U13012 ( .A1(n13070), .A2(n11218), .ZN(n10493) );
  AND2_X1 U13013 ( .A1(n9820), .A2(n10499), .ZN(n11088) );
  NAND2_X2 U13014 ( .A1(n10062), .A2(n10060), .ZN(n19437) );
  NAND4_X1 U13015 ( .A1(n10474), .A2(n10477), .A3(n10475), .A4(n10476), .ZN(
        n10061) );
  NAND4_X1 U13016 ( .A1(n10473), .A2(n10470), .A3(n10472), .A4(n10471), .ZN(
        n10063) );
  XNOR2_X2 U13017 ( .A(n15134), .B(n15133), .ZN(n15146) );
  NAND2_X2 U13018 ( .A1(n10064), .A2(n15132), .ZN(n15134) );
  NOR2_X2 U13019 ( .A1(n10944), .A2(n10943), .ZN(n15154) );
  AND2_X2 U13020 ( .A1(n10066), .A2(n10065), .ZN(n15290) );
  AND2_X2 U13021 ( .A1(n10075), .A2(n17654), .ZN(n16723) );
  AND2_X2 U13022 ( .A1(n10077), .A2(n10076), .ZN(n16767) );
  NOR2_X2 U13023 ( .A1(n15777), .A2(n16519), .ZN(n15838) );
  OR2_X2 U13024 ( .A1(n13010), .A2(n10089), .ZN(n15777) );
  OR2_X2 U13025 ( .A1(n11563), .A2(n18008), .ZN(n13010) );
  NOR2_X2 U13026 ( .A1(n17773), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17772) );
  NAND3_X1 U13027 ( .A1(n10090), .A2(n17781), .A3(n10382), .ZN(n17773) );
  NAND2_X1 U13028 ( .A1(n10595), .A2(n10581), .ZN(n10125) );
  INV_X1 U13029 ( .A(n10599), .ZN(n10091) );
  AND3_X2 U13030 ( .A1(n10790), .A2(n10791), .A3(n11250), .ZN(n10095) );
  AND2_X2 U13031 ( .A1(n10677), .A2(n10676), .ZN(n10790) );
  NAND4_X1 U13032 ( .A1(n9867), .A2(n10403), .A3(n10097), .A4(n9901), .ZN(
        n10404) );
  NAND2_X1 U13033 ( .A1(n9867), .A2(n9914), .ZN(n10096) );
  NAND2_X1 U13034 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10099) );
  INV_X2 U13035 ( .A(n10537), .ZN(n11085) );
  NAND2_X1 U13036 ( .A1(n10127), .A2(n11085), .ZN(n10100) );
  AND2_X1 U13037 ( .A1(n10128), .A2(n11085), .ZN(n10574) );
  INV_X1 U13038 ( .A(n13627), .ZN(n10116) );
  NAND2_X1 U13039 ( .A1(n11885), .A2(n13767), .ZN(n10117) );
  INV_X1 U13040 ( .A(n11834), .ZN(n11883) );
  NAND2_X2 U13041 ( .A1(n10118), .A2(n12716), .ZN(n14648) );
  XNOR2_X2 U13042 ( .A(n10333), .B(n11960), .ZN(n13909) );
  NAND2_X2 U13043 ( .A1(n12049), .A2(n11951), .ZN(n10333) );
  NAND2_X2 U13044 ( .A1(n20507), .A2(n10120), .ZN(n12049) );
  XNOR2_X2 U13045 ( .A(n11933), .B(n11946), .ZN(n20507) );
  NAND2_X1 U13046 ( .A1(n10121), .A2(n10311), .ZN(n10310) );
  NAND3_X1 U13047 ( .A1(n14540), .A2(n9997), .A3(n14556), .ZN(n10121) );
  XNOR2_X1 U13048 ( .A(n14548), .B(n9936), .ZN(n14730) );
  NAND2_X1 U13049 ( .A1(n12108), .A2(n12146), .ZN(n10123) );
  NAND2_X2 U13050 ( .A1(n12085), .A2(n10139), .ZN(n12109) );
  NOR2_X2 U13051 ( .A1(n10123), .A2(n12109), .ZN(n12166) );
  NAND2_X2 U13052 ( .A1(n12674), .A2(n12692), .ZN(n14639) );
  INV_X1 U13053 ( .A(n13081), .ZN(n10596) );
  XNOR2_X1 U13054 ( .A(n10595), .B(n10124), .ZN(n13081) );
  NAND2_X1 U13055 ( .A1(n10790), .A2(n10791), .ZN(n11057) );
  AOI21_X1 U13056 ( .B1(n9853), .B2(n10307), .A(n9868), .ZN(n10131) );
  NAND2_X1 U13057 ( .A1(n10134), .A2(n10133), .ZN(n10132) );
  NAND2_X1 U13058 ( .A1(n10132), .A2(n10306), .ZN(n16341) );
  NAND3_X1 U13059 ( .A1(n13910), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11835) );
  NAND2_X1 U13060 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11779) );
  NAND2_X2 U13061 ( .A1(n14683), .A2(n12701), .ZN(n16019) );
  INV_X1 U13062 ( .A(n12084), .ZN(n10139) );
  OAI21_X1 U13063 ( .B1(n12166), .B2(n12165), .A(n12199), .ZN(n12665) );
  NAND3_X1 U13064 ( .A1(n20565), .A2(n21075), .A3(n12049), .ZN(n10142) );
  NAND2_X1 U13065 ( .A1(n12910), .A2(n9944), .ZN(n14131) );
  INV_X1 U13066 ( .A(n10162), .ZN(n14313) );
  NAND2_X1 U13067 ( .A1(n16192), .A2(n9970), .ZN(n10163) );
  OAI211_X1 U13068 ( .C1(n16192), .C2(n10166), .A(n10163), .B(n10164), .ZN(
        n16172) );
  NAND2_X1 U13069 ( .A1(n16192), .A2(n19182), .ZN(n16180) );
  NAND2_X1 U13070 ( .A1(n16192), .A2(n19182), .ZN(n10168) );
  AOI21_X1 U13071 ( .B1(n10170), .B2(n19192), .A(n20032), .ZN(n10169) );
  AOI21_X4 U13072 ( .B1(n14276), .B2(n16491), .A(n10172), .ZN(n19182) );
  NAND2_X1 U13073 ( .A1(n10186), .A2(n11119), .ZN(n10214) );
  INV_X1 U13074 ( .A(n15300), .ZN(n10187) );
  NAND3_X1 U13075 ( .A1(n10193), .A2(n10194), .A3(n10390), .ZN(n10396) );
  AND2_X1 U13076 ( .A1(n10197), .A2(n10199), .ZN(n10193) );
  INV_X2 U13077 ( .A(n13379), .ZN(n13391) );
  NAND2_X1 U13078 ( .A1(n11132), .A2(n10206), .ZN(n13977) );
  INV_X1 U13079 ( .A(n13379), .ZN(n10633) );
  INV_X2 U13080 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16432) );
  NAND3_X1 U13081 ( .A1(n10223), .A2(n9920), .A3(n10795), .ZN(n10867) );
  NAND2_X1 U13082 ( .A1(n10795), .A2(n10813), .ZN(n10812) );
  INV_X1 U13083 ( .A(n10225), .ZN(n10850) );
  NAND2_X1 U13084 ( .A1(n10890), .A2(n9943), .ZN(n10932) );
  AND2_X1 U13085 ( .A1(n10890), .A2(n10891), .ZN(n10893) );
  NAND2_X1 U13086 ( .A1(n10248), .A2(n10247), .ZN(n11560) );
  NOR2_X2 U13087 ( .A1(n17772), .A2(n17797), .ZN(n17741) );
  NAND3_X1 U13088 ( .A1(n11644), .A2(n10268), .A3(n10267), .ZN(n10266) );
  NAND2_X1 U13089 ( .A1(n17247), .A2(n9988), .ZN(n17229) );
  INV_X1 U13090 ( .A(n10275), .ZN(n13288) );
  NAND3_X1 U13091 ( .A1(n13337), .A2(n10278), .A3(n13339), .ZN(n10276) );
  NAND2_X1 U13092 ( .A1(n14963), .A2(n10281), .ZN(n10277) );
  NOR2_X1 U13093 ( .A1(n14954), .A2(n10279), .ZN(n10278) );
  INV_X1 U13094 ( .A(n10289), .ZN(n14003) );
  NAND2_X1 U13095 ( .A1(n15013), .A2(n9973), .ZN(n10290) );
  AND2_X1 U13096 ( .A1(n15013), .A2(n9957), .ZN(n13240) );
  OAI211_X1 U13097 ( .C1(n15013), .C2(n13264), .A(n10291), .B(n10290), .ZN(
        n15072) );
  NAND2_X1 U13098 ( .A1(n10505), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10415) );
  NAND4_X1 U13099 ( .A1(n10414), .A2(n10412), .A3(n10411), .A4(n10413), .ZN(
        n10505) );
  INV_X1 U13100 ( .A(n10543), .ZN(n10295) );
  NAND2_X1 U13101 ( .A1(n10540), .A2(n9945), .ZN(n10296) );
  OAI21_X2 U13102 ( .B1(n13953), .B2(n12690), .A(n12655), .ZN(n12656) );
  INV_X1 U13103 ( .A(n15161), .ZN(n10300) );
  NAND2_X1 U13104 ( .A1(n15161), .A2(n14258), .ZN(n10301) );
  OR2_X1 U13105 ( .A1(n15161), .A2(n15148), .ZN(n15140) );
  OAI21_X1 U13106 ( .B1(n13714), .B2(n13713), .A(n9912), .ZN(n10313) );
  AND2_X1 U13107 ( .A1(n15040), .A2(n9980), .ZN(n13421) );
  NAND2_X1 U13108 ( .A1(n15040), .A2(n10320), .ZN(n14265) );
  NAND2_X1 U13109 ( .A1(n15040), .A2(n9979), .ZN(n10316) );
  NAND2_X1 U13110 ( .A1(n15040), .A2(n15028), .ZN(n15030) );
  NAND3_X1 U13111 ( .A1(n10317), .A2(n10316), .A3(n10315), .ZN(n16164) );
  AND2_X2 U13112 ( .A1(n15412), .A2(n10328), .ZN(n15053) );
  NAND2_X1 U13113 ( .A1(n13971), .A2(n13973), .ZN(n13972) );
  AND2_X2 U13114 ( .A1(n12360), .A2(n9976), .ZN(n14427) );
  NOR2_X1 U13115 ( .A1(n12817), .A2(n10338), .ZN(n13023) );
  OAI21_X1 U13116 ( .B1(n12817), .B2(n10338), .A(n10337), .ZN(n10336) );
  NOR2_X1 U13117 ( .A1(n12817), .A2(n14300), .ZN(n14289) );
  NAND2_X1 U13118 ( .A1(n14522), .A2(n10347), .ZN(n14435) );
  NOR2_X2 U13119 ( .A1(n14119), .A2(n10352), .ZN(n12285) );
  INV_X1 U13120 ( .A(n10357), .ZN(n13405) );
  AND2_X1 U13121 ( .A1(n10536), .A2(n10357), .ZN(n11086) );
  AOI21_X1 U13122 ( .B1(n19458), .B2(n10357), .A(n11018), .ZN(n10521) );
  MUX2_X1 U13123 ( .A(n10549), .B(n10357), .S(n19458), .Z(n10552) );
  NAND2_X1 U13124 ( .A1(n15154), .A2(n9872), .ZN(n10358) );
  CLKBUF_X1 U13125 ( .A(n10363), .Z(n10359) );
  NAND2_X1 U13126 ( .A1(n15290), .A2(n15292), .ZN(n15213) );
  AOI21_X1 U13127 ( .B1(n15290), .B2(n10368), .A(n9854), .ZN(n15198) );
  NAND2_X1 U13128 ( .A1(n10366), .A2(n10364), .ZN(n15187) );
  NAND2_X1 U13129 ( .A1(n15659), .A2(n10370), .ZN(n10371) );
  NAND2_X1 U13130 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n11556), .ZN(
        n13019) );
  NAND2_X1 U13131 ( .A1(n17986), .A2(n17981), .ZN(n17980) );
  NAND2_X1 U13132 ( .A1(n13817), .A2(n13818), .ZN(n13819) );
  INV_X1 U13133 ( .A(n13080), .ZN(n13817) );
  NAND2_X1 U13134 ( .A1(n14984), .A2(n14986), .ZN(n14985) );
  OR2_X1 U13135 ( .A1(n13769), .A2(n11931), .ZN(n11932) );
  AOI22_X1 U13136 ( .A1(n11798), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11972), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11755) );
  AND4_X1 U13137 ( .A1(n10615), .A2(n10614), .A3(n10613), .A4(n10612), .ZN(
        n10631) );
  NAND2_X1 U13138 ( .A1(n10532), .A2(n10516), .ZN(n11034) );
  AND2_X1 U13139 ( .A1(n10620), .A2(n10626), .ZN(n10714) );
  AND2_X2 U13140 ( .A1(n10620), .A2(n10616), .ZN(n19739) );
  NAND2_X1 U13141 ( .A1(n13895), .A2(n12083), .ZN(n13971) );
  NOR2_X1 U13142 ( .A1(n9823), .A2(n21075), .ZN(n11982) );
  NAND2_X1 U13143 ( .A1(n20306), .A2(n14455), .ZN(n15973) );
  INV_X1 U13144 ( .A(n15973), .ZN(n13038) );
  INV_X1 U13145 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12729) );
  NAND2_X1 U13146 ( .A1(n11216), .A2(n11211), .ZN(n16413) );
  INV_X1 U13147 ( .A(n16413), .ZN(n16406) );
  OR2_X1 U13148 ( .A1(n15328), .A2(n16416), .ZN(n10372) );
  NOR2_X1 U13149 ( .A1(n10926), .A2(n15230), .ZN(n10373) );
  INV_X1 U13150 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10961) );
  AND2_X1 U13151 ( .A1(n11004), .A2(n11219), .ZN(n10374) );
  AND2_X1 U13152 ( .A1(n14234), .A2(n15109), .ZN(n10375) );
  AND2_X1 U13153 ( .A1(n14372), .A2(n14360), .ZN(n10376) );
  AND2_X1 U13154 ( .A1(n10494), .A2(n11217), .ZN(n10378) );
  NAND3_X1 U13155 ( .A1(n12228), .A2(n12227), .A3(n12226), .ZN(n10379) );
  AND3_X1 U13156 ( .A1(n17705), .A2(n18060), .A3(n18048), .ZN(n10380) );
  INV_X1 U13157 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12753) );
  INV_X2 U13158 ( .A(n19003), .ZN(n18933) );
  AND2_X1 U13159 ( .A1(n9841), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10381) );
  INV_X1 U13160 ( .A(n17882), .ZN(n17898) );
  NOR2_X2 U13161 ( .A1(n17992), .A2(n17484), .ZN(n17882) );
  NAND2_X1 U13162 ( .A1(n14265), .A2(n13423), .ZN(n15321) );
  INV_X1 U13163 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11554) );
  OR2_X1 U13164 ( .A1(n17886), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10382) );
  INV_X2 U13165 ( .A(n17361), .ZN(n17358) );
  OR2_X1 U13166 ( .A1(n19372), .A2(n19402), .ZN(n19370) );
  INV_X1 U13167 ( .A(n11519), .ZN(n11498) );
  NOR2_X2 U13168 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20933) );
  NOR2_X1 U13169 ( .A1(n20719), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10383) );
  NOR2_X1 U13170 ( .A1(n17734), .A2(n17827), .ZN(n17973) );
  NOR2_X1 U13171 ( .A1(n17975), .A2(n17989), .ZN(n17734) );
  INV_X1 U13172 ( .A(n17494), .ZN(n17449) );
  AND2_X1 U13173 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10384) );
  AND2_X1 U13174 ( .A1(n13098), .A2(n13097), .ZN(n10385) );
  NAND2_X1 U13175 ( .A1(n13819), .A2(n13104), .ZN(n19209) );
  AND4_X1 U13176 ( .A1(n11839), .A2(n11838), .A3(n11837), .A4(n11836), .ZN(
        n10386) );
  INV_X1 U13177 ( .A(n11798), .ZN(n12611) );
  OAI21_X1 U13178 ( .B1(n12074), .B2(n11926), .A(n11929), .ZN(n11834) );
  OR2_X1 U13179 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n12753), .ZN(
        n12726) );
  INV_X1 U13180 ( .A(n12742), .ZN(n12737) );
  OR2_X1 U13181 ( .A1(n12750), .A2(n13753), .ZN(n12769) );
  AND4_X1 U13182 ( .A1(n12033), .A2(n12032), .A3(n12031), .A4(n12030), .ZN(
        n12037) );
  AND2_X1 U13183 ( .A1(n16432), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10779) );
  OR2_X1 U13184 ( .A1(n12764), .A2(n12148), .ZN(n12164) );
  INV_X1 U13185 ( .A(n12769), .ZN(n12770) );
  NAND2_X1 U13186 ( .A1(n12728), .A2(n12727), .ZN(n12735) );
  INV_X1 U13187 ( .A(n12200), .ZN(n12201) );
  AND2_X1 U13188 ( .A1(n12048), .A2(n12047), .ZN(n12053) );
  NAND2_X1 U13189 ( .A1(n14848), .A2(n9913), .ZN(n10511) );
  AND3_X1 U13190 ( .A1(n10623), .A2(n10622), .A3(n10621), .ZN(n10630) );
  NOR2_X1 U13191 ( .A1(n11228), .A2(n10384), .ZN(n11222) );
  OR2_X1 U13192 ( .A1(n12764), .A2(n12173), .ZN(n12189) );
  INV_X1 U13193 ( .A(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11908) );
  INV_X1 U13194 ( .A(n12208), .ZN(n12209) );
  OR2_X1 U13195 ( .A1(n12764), .A2(n12119), .ZN(n12135) );
  OAI211_X1 U13196 ( .C1(n9851), .C2(n12608), .A(n11809), .B(n11808), .ZN(
        n11810) );
  NAND2_X1 U13197 ( .A1(n12028), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12691) );
  OR2_X1 U13198 ( .A1(n12187), .A2(n12186), .ZN(n12683) );
  AND2_X1 U13199 ( .A1(n10783), .A2(n10782), .ZN(n10786) );
  OR2_X1 U13200 ( .A1(n13284), .A2(n13286), .ZN(n13311) );
  OR2_X1 U13201 ( .A1(n13238), .A2(n13237), .ZN(n13258) );
  AOI22_X1 U13202 ( .A1(n9838), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10421), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10447) );
  NAND2_X1 U13203 ( .A1(n19470), .A2(n10758), .ZN(n10759) );
  AND2_X1 U13204 ( .A1(n19470), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n10934) );
  AND4_X1 U13205 ( .A1(n10738), .A2(n10737), .A3(n10736), .A4(n10735), .ZN(
        n10756) );
  INV_X1 U13206 ( .A(n11066), .ZN(n10845) );
  INV_X1 U13207 ( .A(n14437), .ZN(n12359) );
  AND2_X1 U13208 ( .A1(n12189), .A2(n12188), .ZN(n12200) );
  AND2_X1 U13209 ( .A1(n12581), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12582) );
  INV_X1 U13210 ( .A(n12492), .ZN(n12493) );
  OR2_X1 U13211 ( .A1(n11888), .A2(n21075), .ZN(n12875) );
  NOR2_X1 U13212 ( .A1(n12112), .A2(n12111), .ZN(n12138) );
  INV_X1 U13213 ( .A(n11847), .ZN(n11848) );
  INV_X1 U13214 ( .A(n14173), .ZN(n13110) );
  AND2_X1 U13215 ( .A1(n11411), .A2(n11410), .ZN(n15054) );
  AND2_X1 U13216 ( .A1(n16248), .A2(n10938), .ZN(n10939) );
  AND2_X1 U13217 ( .A1(n11399), .A2(n11398), .ZN(n15462) );
  INV_X1 U13218 ( .A(n16326), .ZN(n11146) );
  INV_X1 U13219 ( .A(n16342), .ZN(n11077) );
  AND2_X1 U13220 ( .A1(n20165), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10975) );
  NAND2_X1 U13221 ( .A1(n13077), .A2(n13076), .ZN(n13332) );
  NOR2_X1 U13222 ( .A1(n10627), .A2(n10618), .ZN(n10706) );
  INV_X1 U13223 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17272) );
  INV_X1 U13224 ( .A(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17252) );
  OR2_X1 U13225 ( .A1(n12895), .A2(n12894), .ZN(n12896) );
  OAI211_X1 U13226 ( .C1(n11953), .C2(n10020), .A(n11959), .B(n11958), .ZN(
        n11960) );
  AND2_X1 U13227 ( .A1(n12790), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12791) );
  NOR2_X1 U13228 ( .A1(n12414), .A2(n14402), .ZN(n12415) );
  NOR2_X1 U13229 ( .A1(n12303), .A2(n12302), .ZN(n12321) );
  INV_X1 U13230 ( .A(n13997), .ZN(n14042) );
  INV_X1 U13231 ( .A(n12974), .ZN(n12952) );
  AND2_X1 U13232 ( .A1(n11926), .A2(n11917), .ZN(n13610) );
  NAND2_X1 U13233 ( .A1(n13620), .A2(n13619), .ZN(n15805) );
  OR2_X1 U13234 ( .A1(n19414), .A2(n14155), .ZN(n14156) );
  AND2_X1 U13235 ( .A1(n19263), .A2(n19264), .ZN(n13109) );
  OR2_X1 U13236 ( .A1(n11341), .A2(n11340), .ZN(n19269) );
  INV_X1 U13237 ( .A(n13332), .ZN(n13304) );
  AND2_X1 U13238 ( .A1(n11401), .A2(n11400), .ZN(n15091) );
  AND3_X1 U13239 ( .A1(n11153), .A2(n11152), .A3(n11151), .ZN(n15302) );
  INV_X1 U13240 ( .A(n15109), .ZN(n14241) );
  OR2_X1 U13241 ( .A1(n10920), .A2(n15251), .ZN(n15245) );
  OR2_X1 U13242 ( .A1(n10879), .A2(n10878), .ZN(n16319) );
  NAND2_X1 U13243 ( .A1(n11061), .A2(n11060), .ZN(n14115) );
  BUF_X1 U13244 ( .A(n10713), .Z(n19582) );
  INV_X1 U13245 ( .A(n10823), .ZN(n19926) );
  AND2_X1 U13246 ( .A1(n11213), .A2(n15638), .ZN(n15658) );
  INV_X1 U13247 ( .A(n13012), .ZN(n13013) );
  NOR2_X1 U13248 ( .A1(n11558), .A2(n10380), .ZN(n11559) );
  INV_X1 U13249 ( .A(n18185), .ZN(n18229) );
  INV_X1 U13250 ( .A(n17487), .ZN(n11718) );
  NOR2_X1 U13251 ( .A1(n11662), .A2(n11647), .ZN(n11681) );
  INV_X1 U13252 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14402) );
  INV_X1 U13253 ( .A(n20250), .ZN(n15951) );
  AND2_X1 U13254 ( .A1(n15832), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12893) );
  NAND2_X1 U13255 ( .A1(n14029), .A2(n12994), .ZN(n20276) );
  AND2_X1 U13256 ( .A1(n12973), .A2(n12972), .ZN(n14314) );
  INV_X1 U13257 ( .A(n14424), .ZN(n14800) );
  NAND2_X1 U13258 ( .A1(n12791), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12846) );
  INV_X1 U13259 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14615) );
  AND2_X1 U13260 ( .A1(n12167), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12191) );
  NAND2_X1 U13261 ( .A1(n12766), .A2(n12887), .ZN(n12780) );
  AND2_X1 U13262 ( .A1(n10119), .A2(n14674), .ZN(n16009) );
  NOR2_X1 U13263 ( .A1(n13793), .A2(n20366), .ZN(n16105) );
  INV_X1 U13264 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14826) );
  INV_X1 U13265 ( .A(n12640), .ZN(n20376) );
  OR2_X1 U13266 ( .A1(n13948), .A2(n20479), .ZN(n20851) );
  AND2_X1 U13267 ( .A1(n13948), .A2(n20479), .ZN(n20590) );
  INV_X1 U13268 ( .A(n20933), .ZN(n20926) );
  AND2_X1 U13269 ( .A1(n13946), .A2(n13945), .ZN(n15822) );
  AND2_X1 U13270 ( .A1(n11102), .A2(n11101), .ZN(n16430) );
  OR3_X1 U13271 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n14150), .A3(n14149), .ZN(
        n14151) );
  AND3_X1 U13272 ( .A1(n11205), .A2(n11204), .A3(n11203), .ZN(n14959) );
  AND2_X1 U13273 ( .A1(n19347), .A2(n13427), .ZN(n13678) );
  AND3_X1 U13274 ( .A1(n11163), .A2(n11162), .A3(n11161), .ZN(n14172) );
  INV_X1 U13275 ( .A(n14873), .ZN(n14875) );
  INV_X1 U13276 ( .A(n19414), .ZN(n19176) );
  OR2_X1 U13277 ( .A1(n19501), .A2(n19496), .ZN(n19542) );
  OR2_X1 U13278 ( .A1(n19702), .A2(n19701), .ZN(n19708) );
  OR2_X1 U13279 ( .A1(n19611), .A2(n20152), .ZN(n19764) );
  NAND2_X1 U13280 ( .A1(n19611), .A2(n20130), .ZN(n19898) );
  NAND3_X1 U13281 ( .A1(n20126), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19974), 
        .ZN(n19435) );
  INV_X1 U13282 ( .A(n19480), .ZN(n19482) );
  NAND2_X1 U13283 ( .A1(n16491), .A2(n16479), .ZN(n16478) );
  NOR2_X1 U13284 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16846), .ZN(n16829) );
  NOR2_X1 U13285 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16943), .ZN(n16915) );
  INV_X1 U13286 ( .A(n17009), .ZN(n17023) );
  INV_X1 U13287 ( .A(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17236) );
  NOR2_X1 U13288 ( .A1(n18015), .A2(n17660), .ZN(n17997) );
  INV_X1 U13289 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17736) );
  INV_X1 U13290 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17769) );
  INV_X1 U13291 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16868) );
  INV_X1 U13292 ( .A(n11542), .ZN(n11543) );
  INV_X1 U13293 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18060) );
  NOR2_X1 U13294 ( .A1(n18797), .A2(n18791), .ZN(n18285) );
  NOR2_X1 U13295 ( .A1(n18163), .A2(n17851), .ZN(n18176) );
  OAI221_X1 U13296 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(n19005), .C1(n18965), 
        .C2(P3_STATE2_REG_2__SCAN_IN), .A(n18954), .ZN(n18334) );
  INV_X1 U13297 ( .A(n17989), .ZN(n17824) );
  NOR2_X1 U13298 ( .A1(n15893), .A2(n13005), .ZN(n14357) );
  NOR2_X1 U13299 ( .A1(n15915), .A2(n15894), .ZN(n14398) );
  NOR2_X1 U13300 ( .A1(n21381), .A2(n20210), .ZN(n15963) );
  OR3_X1 U13301 ( .A1(n13501), .A2(n12893), .A3(n12892), .ZN(n14408) );
  INV_X1 U13302 ( .A(n14530), .ZN(n14534) );
  NAND2_X1 U13303 ( .A1(n13047), .A2(n13757), .ZN(n13048) );
  INV_X1 U13304 ( .A(n13745), .ZN(n13845) );
  AOI21_X1 U13305 ( .B1(n12579), .B2(n12578), .A(n12577), .ZN(n14338) );
  NAND2_X1 U13306 ( .A1(n12435), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12492) );
  NAND2_X1 U13307 ( .A1(n12380), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12414) );
  NAND2_X1 U13308 ( .A1(n12268), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12303) );
  INV_X1 U13309 ( .A(n14689), .ZN(n20374) );
  INV_X1 U13310 ( .A(n20187), .ZN(n16034) );
  NAND2_X1 U13311 ( .A1(n13766), .A2(n13765), .ZN(n13783) );
  NOR2_X1 U13312 ( .A1(n14706), .A2(n14813), .ZN(n15859) );
  OR2_X1 U13313 ( .A1(n16104), .A2(n13802), .ZN(n14796) );
  INV_X1 U13314 ( .A(n20369), .ZN(n16106) );
  OR2_X1 U13315 ( .A1(n20366), .A2(n20360), .ZN(n16104) );
  NAND2_X1 U13316 ( .A1(n12658), .A2(n12657), .ZN(n13984) );
  INV_X1 U13317 ( .A(n20355), .ZN(n16135) );
  NAND2_X1 U13318 ( .A1(n21075), .A2(n20379), .ZN(n20542) );
  OAI22_X1 U13319 ( .A1(n20391), .A2(n20390), .B1(n20663), .B2(n20538), .ZN(
        n20448) );
  AND2_X1 U13320 ( .A1(n20376), .A2(n13953), .ZN(n20480) );
  AND2_X1 U13321 ( .A1(n20480), .A2(n20457), .ZN(n20502) );
  AND2_X1 U13322 ( .A1(n20480), .A2(n20590), .ZN(n20532) );
  NOR2_X2 U13323 ( .A1(n20512), .A2(n20762), .ZN(n20560) );
  INV_X1 U13324 ( .A(n20622), .ZN(n20618) );
  INV_X1 U13325 ( .A(n20624), .ZN(n20653) );
  INV_X1 U13326 ( .A(n20664), .ZN(n20685) );
  INV_X1 U13327 ( .A(n20784), .ZN(n20657) );
  INV_X1 U13328 ( .A(n20783), .ZN(n20741) );
  OAI21_X1 U13329 ( .B1(n20761), .B2(n20760), .A(n20759), .ZN(n20780) );
  INV_X1 U13330 ( .A(n20785), .ZN(n20837) );
  OR2_X1 U13331 ( .A1(n13948), .A2(n20377), .ZN(n20784) );
  NOR2_X2 U13332 ( .A1(n20925), .A2(n20851), .ZN(n20914) );
  INV_X1 U13333 ( .A(n20969), .ZN(n20982) );
  INV_X1 U13334 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n16145) );
  INV_X1 U13335 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n21007) );
  AND2_X1 U13336 ( .A1(n21038), .A2(n21007), .ZN(n21043) );
  NAND2_X1 U13337 ( .A1(n16255), .A2(n16256), .ZN(n16254) );
  INV_X1 U13338 ( .A(n19204), .ZN(n19241) );
  AND2_X1 U13339 ( .A1(n19014), .A2(n16482), .ZN(n19239) );
  INV_X1 U13340 ( .A(n19222), .ZN(n19242) );
  NOR2_X1 U13341 ( .A1(n19182), .A2(n20032), .ZN(n19251) );
  INV_X1 U13342 ( .A(n15189), .ZN(n15204) );
  INV_X1 U13343 ( .A(n11217), .ZN(n13426) );
  INV_X1 U13344 ( .A(n19347), .ZN(n19356) );
  INV_X1 U13345 ( .A(n13504), .ZN(n19405) );
  INV_X1 U13346 ( .A(n13469), .ZN(n19407) );
  INV_X1 U13347 ( .A(n19417), .ZN(n16366) );
  AND2_X1 U13348 ( .A1(n13535), .A2(n20168), .ZN(n19421) );
  INV_X1 U13349 ( .A(n13095), .ZN(n15643) );
  XNOR2_X1 U13350 ( .A(n13746), .B(n10385), .ZN(n19611) );
  OAI21_X2 U13351 ( .B1(n20121), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n15867), 
        .ZN(n19974) );
  NOR2_X1 U13352 ( .A1(n20132), .A2(n20160), .ZN(n19576) );
  INV_X1 U13353 ( .A(n19606), .ZN(n19592) );
  OAI21_X1 U13354 ( .B1(n19617), .B2(n19616), .A(n19615), .ZN(n19635) );
  NOR2_X1 U13355 ( .A1(n19668), .A2(n19898), .ZN(n19663) );
  NOR2_X1 U13356 ( .A1(n19709), .A2(n19898), .ZN(n19685) );
  NOR2_X1 U13357 ( .A1(n19709), .A2(n19920), .ZN(n19758) );
  NOR2_X1 U13358 ( .A1(n19921), .A2(n19764), .ZN(n19790) );
  NOR2_X1 U13359 ( .A1(n19921), .A2(n20127), .ZN(n19840) );
  NOR2_X1 U13360 ( .A1(n19921), .A2(n19898), .ZN(n19890) );
  NOR2_X2 U13361 ( .A1(n19899), .A2(n19898), .ZN(n19959) );
  OAI22_X1 U13362 ( .A1(n19474), .A2(n19482), .B1(n20434), .B2(n19484), .ZN(
        n19954) );
  AND4_X1 U13363 ( .A1(n13669), .A2(n13668), .A3(n13667), .A4(n13666), .ZN(
        n16474) );
  INV_X1 U13364 ( .A(n14851), .ZN(n20047) );
  INV_X1 U13365 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20055) );
  NAND4_X1 U13366 ( .A1(n18355), .A2(n11659), .A3(n11672), .A4(n17516), .ZN(
        n18775) );
  NOR2_X1 U13367 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16740), .ZN(n16726) );
  NOR2_X1 U13368 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16759), .ZN(n16744) );
  NOR2_X1 U13369 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16780), .ZN(n16763) );
  NOR2_X1 U13370 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16818), .ZN(n16811) );
  NOR2_X1 U13371 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16865), .ZN(n16853) );
  NOR2_X1 U13372 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16906), .ZN(n16905) );
  INV_X1 U13373 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16920) );
  INV_X1 U13374 ( .A(n17034), .ZN(n16973) );
  NAND2_X1 U13375 ( .A1(n16649), .A2(n16650), .ZN(n17034) );
  NOR2_X1 U13376 ( .A1(n17576), .A2(n17394), .ZN(n17389) );
  NOR4_X1 U13377 ( .A1(n17568), .A2(n17558), .A3(n17444), .A4(n17410), .ZN(
        n17405) );
  NAND2_X1 U13378 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17448), .ZN(n17444) );
  INV_X1 U13379 ( .A(n17552), .ZN(n17517) );
  NOR2_X1 U13380 ( .A1(n17684), .A2(n18030), .ZN(n17661) );
  INV_X1 U13381 ( .A(n13019), .ZN(n18186) );
  INV_X1 U13382 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18127) );
  NOR2_X1 U13383 ( .A1(n18993), .A2(n18268), .ZN(n18231) );
  INV_X1 U13384 ( .A(n18312), .ZN(n18308) );
  INV_X1 U13385 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18965) );
  INV_X1 U13386 ( .A(n18816), .ZN(n18815) );
  INV_X1 U13387 ( .A(n18437), .ZN(n18426) );
  INV_X1 U13388 ( .A(n18484), .ZN(n18473) );
  INV_X1 U13389 ( .A(n18533), .ZN(n18526) );
  INV_X1 U13390 ( .A(n18549), .ZN(n18553) );
  INV_X1 U13391 ( .A(n18600), .ZN(n18602) );
  INV_X1 U13392 ( .A(n18626), .ZN(n18619) );
  INV_X1 U13393 ( .A(n18652), .ZN(n18643) );
  INV_X1 U13394 ( .A(n18331), .ZN(n18582) );
  INV_X1 U13395 ( .A(n18711), .ZN(n18701) );
  AND2_X1 U13396 ( .A1(n18536), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18724) );
  NAND2_X1 U13397 ( .A1(n13764), .A2(n12881), .ZN(n13701) );
  INV_X1 U13398 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20848) );
  AND2_X1 U13399 ( .A1(n13007), .A2(n13006), .ZN(n13008) );
  NAND2_X1 U13400 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n14398), .ZN(n15893) );
  NAND2_X1 U13401 ( .A1(n14408), .A2(n12897), .ZN(n15960) );
  INV_X1 U13402 ( .A(n14418), .ZN(n14702) );
  NAND2_X1 U13403 ( .A1(n20310), .A2(n20380), .ZN(n13816) );
  INV_X1 U13404 ( .A(n20310), .ZN(n20338) );
  OR2_X1 U13405 ( .A1(n20348), .A2(n13753), .ZN(n13745) );
  NAND2_X1 U13406 ( .A1(n16038), .A2(n13695), .ZN(n16031) );
  NAND2_X1 U13407 ( .A1(n20187), .A2(n12781), .ZN(n16038) );
  NAND2_X1 U13408 ( .A1(n13783), .A2(n13776), .ZN(n20355) );
  INV_X1 U13409 ( .A(n20357), .ZN(n16112) );
  INV_X1 U13410 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20843) );
  NAND2_X1 U13411 ( .A1(n20480), .A2(n20657), .ZN(n20477) );
  AOI22_X1 U13412 ( .A1(n20482), .A2(n20485), .B1(n10383), .B2(n20714), .ZN(
        n20506) );
  AOI22_X1 U13413 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20511), .B1(n20515), 
        .B2(n20510), .ZN(n20536) );
  OR2_X1 U13414 ( .A1(n20629), .A2(n20784), .ZN(n20589) );
  AOI22_X1 U13415 ( .A1(n20597), .A2(n20594), .B1(n20790), .B2(n10383), .ZN(
        n20628) );
  OR2_X1 U13416 ( .A1(n20629), .A2(n20762), .ZN(n20664) );
  NAND2_X1 U13417 ( .A1(n20658), .A2(n20657), .ZN(n20712) );
  AOI22_X1 U13418 ( .A1(n20718), .A2(n20716), .B1(n20714), .B2(n20882), .ZN(
        n20750) );
  OR2_X1 U13419 ( .A1(n20763), .A2(n20880), .ZN(n20783) );
  INV_X1 U13420 ( .A(n20923), .ZN(n20803) );
  INV_X1 U13421 ( .A(n20963), .ZN(n20828) );
  OR2_X1 U13422 ( .A1(n20925), .A2(n20784), .ZN(n20878) );
  INV_X1 U13423 ( .A(n20965), .ZN(n20909) );
  INV_X1 U13424 ( .A(n20852), .ZN(n20938) );
  INV_X1 U13425 ( .A(n20860), .ZN(n20956) );
  INV_X1 U13426 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n21075) );
  INV_X1 U13427 ( .A(n21058), .ZN(n20993) );
  INV_X1 U13428 ( .A(n21054), .ZN(n21058) );
  INV_X1 U13429 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21332) );
  INV_X1 U13430 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n21381) );
  INV_X1 U13431 ( .A(n14848), .ZN(n13447) );
  INV_X1 U13432 ( .A(n19252), .ZN(n19223) );
  INV_X1 U13433 ( .A(n19226), .ZN(n19246) );
  AND2_X2 U13434 ( .A1(n13557), .A2(n20027), .ZN(n19293) );
  NAND2_X1 U13435 ( .A1(n19347), .A2(n13426), .ZN(n19348) );
  AND2_X1 U13436 ( .A1(n13404), .A2(n20027), .ZN(n19347) );
  NAND2_X1 U13437 ( .A1(n19347), .A2(n13405), .ZN(n19361) );
  NAND2_X1 U13438 ( .A1(n19372), .A2(n14846), .ZN(n19367) );
  INV_X1 U13439 ( .A(n19372), .ZN(n19404) );
  OR2_X1 U13440 ( .A1(n14150), .A2(n13449), .ZN(n13469) );
  INV_X1 U13441 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n19091) );
  INV_X1 U13442 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n19141) );
  INV_X1 U13443 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19153) );
  NAND2_X1 U13444 ( .A1(n13533), .A2(n13532), .ZN(n19425) );
  NAND2_X1 U13445 ( .A1(n11216), .A2(n11047), .ZN(n16416) );
  NAND2_X1 U13446 ( .A1(n11216), .A2(n11215), .ZN(n16412) );
  INV_X1 U13447 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n19457) );
  AND2_X1 U13448 ( .A1(n19434), .A2(n19974), .ZN(n19487) );
  NAND2_X1 U13449 ( .A1(n19500), .A2(n19576), .ZN(n19563) );
  OR2_X1 U13450 ( .A1(n19668), .A2(n20127), .ZN(n19606) );
  INV_X1 U13451 ( .A(n19628), .ZN(n19638) );
  INV_X1 U13452 ( .A(n19663), .ZN(n19661) );
  INV_X1 U13453 ( .A(n19685), .ZN(n19697) );
  INV_X1 U13454 ( .A(n19723), .ZN(n19732) );
  INV_X1 U13455 ( .A(n19790), .ZN(n19789) );
  INV_X1 U13456 ( .A(n19823), .ZN(n19811) );
  INV_X1 U13457 ( .A(n19976), .ZN(n19839) );
  INV_X1 U13458 ( .A(n19840), .ZN(n19859) );
  INV_X1 U13459 ( .A(n19865), .ZN(n19889) );
  INV_X1 U13460 ( .A(n19890), .ZN(n19918) );
  AOI21_X1 U13461 ( .B1(n19930), .B2(n19932), .A(n19928), .ZN(n19963) );
  INV_X1 U13462 ( .A(n19947), .ZN(n20003) );
  INV_X1 U13463 ( .A(n19958), .ZN(n20026) );
  INV_X1 U13464 ( .A(n20119), .ZN(n20035) );
  OR2_X1 U13465 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19017), .ZN(n20175) );
  NOR2_X1 U13466 ( .A1(n18828), .A2(n18777), .ZN(n17553) );
  INV_X1 U13467 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17676) );
  NAND2_X1 U13468 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n17034), .ZN(n16969) );
  INV_X1 U13469 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16875) );
  INV_X1 U13470 ( .A(n17007), .ZN(n17031) );
  INV_X1 U13471 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17331) );
  AND2_X1 U13472 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17463), .ZN(n17466) );
  NOR2_X1 U13473 ( .A1(n17603), .A2(n17479), .ZN(n17482) );
  NAND2_X1 U13474 ( .A1(n17517), .A2(n17516), .ZN(n17534) );
  NAND2_X1 U13475 ( .A1(n17553), .A2(n17515), .ZN(n17552) );
  INV_X1 U13476 ( .A(n17794), .ZN(n17774) );
  INV_X1 U13477 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18113) );
  INV_X1 U13478 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17851) );
  INV_X1 U13479 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18214) );
  OR2_X1 U13480 ( .A1(n18068), .A2(n17637), .ZN(n13022) );
  INV_X1 U13481 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18048) );
  INV_X1 U13482 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18096) );
  INV_X1 U13483 ( .A(n18219), .ZN(n18237) );
  NAND2_X1 U13484 ( .A1(n18312), .A2(n10081), .ZN(n18310) );
  INV_X1 U13485 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18820) );
  AOI211_X1 U13486 ( .C1(n18991), .C2(n18815), .A(n18335), .B(n15773), .ZN(
        n18973) );
  INV_X1 U13487 ( .A(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n18373) );
  INV_X1 U13488 ( .A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18387) );
  INV_X1 U13489 ( .A(n18507), .ZN(n18505) );
  INV_X1 U13490 ( .A(n18720), .ZN(n18684) );
  INV_X1 U13491 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18942) );
  INV_X1 U13492 ( .A(n18939), .ZN(n18936) );
  NOR2_X1 U13493 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13435), .ZN(n16618)
         );
  INV_X1 U13494 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20059) );
  OAI21_X1 U13495 ( .B1(n14459), .B2(n15974), .A(n13039), .ZN(P1_U2842) );
  OAI21_X1 U13496 ( .B1(n15131), .B2(n16425), .A(n11428), .ZN(P2_U3017) );
  INV_X1 U13497 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10695) );
  INV_X1 U13498 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10387) );
  OAI22_X1 U13499 ( .A1(n10436), .A2(n10695), .B1(n13249), .B2(n10387), .ZN(
        n10388) );
  INV_X1 U13500 ( .A(n10388), .ZN(n10390) );
  INV_X1 U13501 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10389) );
  INV_X1 U13502 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10394) );
  INV_X1 U13503 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10393) );
  OAI22_X1 U13504 ( .A1(n9835), .A2(n10394), .B1(n13242), .B2(n10393), .ZN(
        n10395) );
  NAND2_X1 U13505 ( .A1(n10503), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10405) );
  INV_X1 U13506 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10397) );
  INV_X1 U13507 ( .A(n10398), .ZN(n10403) );
  INV_X1 U13508 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10400) );
  INV_X1 U13509 ( .A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10399) );
  OAI22_X1 U13510 ( .A1(n10436), .A2(n10400), .B1(n13249), .B2(n10399), .ZN(
        n10401) );
  INV_X1 U13511 ( .A(n10401), .ZN(n10402) );
  AOI22_X1 U13512 ( .A1(n9838), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10421), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10409) );
  AOI22_X1 U13513 ( .A1(n10482), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13312), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10408) );
  AOI22_X1 U13514 ( .A1(n9841), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(n9814), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10407) );
  NAND4_X1 U13515 ( .A1(n10409), .A2(n10408), .A3(n10407), .A4(n10406), .ZN(
        n10506) );
  AOI22_X1 U13516 ( .A1(n9838), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(n9808), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10414) );
  AOI22_X1 U13517 ( .A1(n10482), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13312), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10413) );
  AOI22_X1 U13518 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9816), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10412) );
  AOI22_X1 U13519 ( .A1(n9841), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9815), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10411) );
  NAND2_X1 U13520 ( .A1(n10416), .A2(n10415), .ZN(n10491) );
  AOI22_X1 U13521 ( .A1(n10482), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13312), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10419) );
  AOI22_X1 U13522 ( .A1(n13391), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9815), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10417) );
  NAND4_X1 U13523 ( .A1(n10420), .A2(n10419), .A3(n10418), .A4(n10417), .ZN(
        n10429) );
  AOI22_X1 U13524 ( .A1(n9834), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13312), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10426) );
  AOI22_X1 U13525 ( .A1(n13391), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9814), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10424) );
  NAND4_X1 U13526 ( .A1(n10427), .A2(n10426), .A3(n10425), .A4(n10424), .ZN(
        n10428) );
  AOI22_X1 U13527 ( .A1(n9842), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9815), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10430) );
  AOI22_X1 U13528 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10634), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10433) );
  AOI22_X1 U13529 ( .A1(n10482), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13312), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10431) );
  AOI22_X1 U13530 ( .A1(n9834), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13312), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10434) );
  AOI22_X1 U13531 ( .A1(n9840), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10634), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10439) );
  AOI22_X1 U13532 ( .A1(n13391), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9814), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10438) );
  NAND4_X1 U13533 ( .A1(n10440), .A2(n10439), .A3(n10438), .A4(n10437), .ZN(
        n10441) );
  AOI22_X1 U13534 ( .A1(n9841), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(n9814), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10445) );
  AND2_X1 U13535 ( .A1(n10445), .A2(n10444), .ZN(n10449) );
  AOI22_X1 U13536 ( .A1(n9840), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(n9817), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10448) );
  AOI22_X1 U13537 ( .A1(n9834), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13312), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10446) );
  NAND4_X1 U13538 ( .A1(n10449), .A2(n10448), .A3(n10447), .A4(n10446), .ZN(
        n10456) );
  AOI22_X1 U13539 ( .A1(n9834), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13312), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10452) );
  AOI22_X1 U13540 ( .A1(n9840), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9817), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10454) );
  AOI22_X1 U13541 ( .A1(n13392), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9807), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10453) );
  NAND3_X1 U13542 ( .A1(n9899), .A2(n10454), .A3(n10453), .ZN(n10455) );
  AOI22_X1 U13543 ( .A1(n10482), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13312), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10457) );
  NOR2_X1 U13544 ( .A1(n10458), .A2(n10444), .ZN(n10462) );
  AOI22_X1 U13545 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10634), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10461) );
  AOI22_X1 U13546 ( .A1(n13392), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10421), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10460) );
  AOI22_X1 U13547 ( .A1(n9841), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9815), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10459) );
  NAND4_X1 U13548 ( .A1(n10462), .A2(n10461), .A3(n10460), .A4(n10459), .ZN(
        n10468) );
  NOR2_X1 U13549 ( .A1(n10381), .A2(n9866), .ZN(n10466) );
  AOI22_X1 U13550 ( .A1(n9840), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10634), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10465) );
  AOI22_X1 U13551 ( .A1(n9838), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10421), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10464) );
  AOI22_X1 U13552 ( .A1(n9834), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13312), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10463) );
  NAND4_X1 U13553 ( .A1(n10466), .A2(n10465), .A3(n10464), .A4(n10463), .ZN(
        n10467) );
  NOR2_X2 U13554 ( .A1(n10525), .A2(n11031), .ZN(n11016) );
  AOI22_X1 U13555 ( .A1(n13392), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10421), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10473) );
  AOI22_X1 U13556 ( .A1(n9834), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13312), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10472) );
  AOI22_X1 U13557 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10634), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10471) );
  AOI22_X1 U13558 ( .A1(n13391), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9815), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10470) );
  AOI22_X1 U13559 ( .A1(n9834), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13312), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10476) );
  AOI22_X1 U13560 ( .A1(n9840), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9816), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10475) );
  AOI22_X1 U13561 ( .A1(n9841), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9814), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10474) );
  NAND2_X1 U13562 ( .A1(n11016), .A2(n14846), .ZN(n10541) );
  AOI22_X1 U13563 ( .A1(n13392), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9808), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10481) );
  AOI22_X1 U13564 ( .A1(n9834), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13312), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10480) );
  AOI22_X1 U13565 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9816), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10479) );
  AOI22_X1 U13566 ( .A1(n13391), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9815), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10478) );
  NAND4_X1 U13567 ( .A1(n10481), .A2(n10480), .A3(n10479), .A4(n10478), .ZN(
        n10489) );
  AOI22_X1 U13568 ( .A1(n13392), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9808), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10487) );
  AOI22_X1 U13569 ( .A1(n10482), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13312), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U13570 ( .A1(n9840), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9817), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10485) );
  AOI22_X1 U13571 ( .A1(n13391), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9814), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10484) );
  NAND4_X1 U13572 ( .A1(n10487), .A2(n10486), .A3(n10485), .A4(n10484), .ZN(
        n10488) );
  MUX2_X2 U13573 ( .A(n10489), .B(n10488), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n11225) );
  INV_X1 U13574 ( .A(n10589), .ZN(n10490) );
  NAND2_X1 U13575 ( .A1(n10490), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10515) );
  AOI22_X1 U13576 ( .A1(n10574), .A2(P2_EBX_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10514) );
  INV_X1 U13577 ( .A(n10493), .ZN(n10494) );
  NAND3_X1 U13578 ( .A1(n10496), .A2(n11030), .A3(n10495), .ZN(n10523) );
  NAND2_X1 U13579 ( .A1(n11207), .A2(n11020), .ZN(n10498) );
  NAND2_X1 U13580 ( .A1(n10498), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10542) );
  INV_X1 U13581 ( .A(n10499), .ZN(n10500) );
  NAND2_X2 U13582 ( .A1(n10500), .A2(n14159), .ZN(n14848) );
  INV_X1 U13583 ( .A(n11031), .ZN(n10501) );
  NAND2_X1 U13584 ( .A1(n10501), .A2(n10536), .ZN(n10549) );
  INV_X1 U13585 ( .A(n10549), .ZN(n10510) );
  INV_X1 U13586 ( .A(n10503), .ZN(n10504) );
  NAND4_X1 U13587 ( .A1(n10505), .A2(n10504), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10508) );
  NAND4_X1 U13588 ( .A1(n10506), .A2(n9871), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n10444), .ZN(n10507) );
  NAND2_X1 U13589 ( .A1(n10567), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10513) );
  NAND2_X1 U13590 ( .A1(n10516), .A2(n10550), .ZN(n10519) );
  INV_X1 U13591 ( .A(n10517), .ZN(n10518) );
  NAND2_X1 U13592 ( .A1(n10519), .A2(n10518), .ZN(n10522) );
  NAND2_X1 U13593 ( .A1(n10522), .A2(n10521), .ZN(n10524) );
  NAND3_X1 U13594 ( .A1(n10524), .A2(n11089), .A3(n10523), .ZN(n10557) );
  INV_X1 U13595 ( .A(n10525), .ZN(n10526) );
  NAND2_X1 U13596 ( .A1(n11014), .A2(n10528), .ZN(n11212) );
  NOR2_X1 U13597 ( .A1(n11016), .A2(n10972), .ZN(n10529) );
  NAND2_X1 U13598 ( .A1(n11212), .A2(n10529), .ZN(n10561) );
  NAND2_X1 U13599 ( .A1(n10537), .A2(n10530), .ZN(n10535) );
  AND2_X1 U13600 ( .A1(n11031), .A2(n19464), .ZN(n10532) );
  NAND2_X1 U13601 ( .A1(n11034), .A2(n10533), .ZN(n11083) );
  NAND2_X1 U13602 ( .A1(n11083), .A2(n19458), .ZN(n10534) );
  NAND2_X1 U13603 ( .A1(n10535), .A2(n10534), .ZN(n10556) );
  NAND2_X1 U13604 ( .A1(n10556), .A2(n20169), .ZN(n10538) );
  NAND2_X1 U13605 ( .A1(n10537), .A2(n11086), .ZN(n10560) );
  NAND2_X1 U13606 ( .A1(n10560), .A2(n11089), .ZN(n10558) );
  NAND3_X1 U13607 ( .A1(n10539), .A2(n10538), .A3(n10558), .ZN(n10540) );
  OAI211_X1 U13608 ( .C1(n16478), .C2(n16450), .A(n10542), .B(n10541), .ZN(
        n10543) );
  NAND2_X1 U13609 ( .A1(n10545), .A2(n10544), .ZN(n10571) );
  NAND2_X1 U13610 ( .A1(n10546), .A2(n10571), .ZN(n10599) );
  NAND2_X1 U13611 ( .A1(n20169), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10547) );
  NOR2_X1 U13612 ( .A1(n10547), .A2(n11025), .ZN(n10548) );
  OAI22_X1 U13613 ( .A1(n9859), .A2(n10548), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n10574), .ZN(n10555) );
  NAND2_X1 U13614 ( .A1(n14848), .A2(n10550), .ZN(n10551) );
  NOR2_X1 U13615 ( .A1(n16478), .A2(n20165), .ZN(n10553) );
  AOI21_X1 U13616 ( .B1(n15661), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10553), 
        .ZN(n10554) );
  NAND2_X1 U13617 ( .A1(n10555), .A2(n10554), .ZN(n10603) );
  NAND2_X1 U13618 ( .A1(n10558), .A2(n11092), .ZN(n10559) );
  AOI21_X1 U13619 ( .B1(n10556), .B2(n10560), .A(n10559), .ZN(n10570) );
  INV_X1 U13620 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n10562) );
  OAI21_X1 U13621 ( .B1(n10589), .B2(n10562), .A(n10561), .ZN(n10566) );
  INV_X1 U13622 ( .A(n10574), .ZN(n10564) );
  INV_X1 U13623 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13558) );
  NAND2_X1 U13624 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10563) );
  NOR2_X1 U13625 ( .A1(n10566), .A2(n10565), .ZN(n10569) );
  NAND2_X1 U13626 ( .A1(n10588), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10568) );
  OAI211_X1 U13627 ( .C1(n10570), .C2(n16491), .A(n10569), .B(n10568), .ZN(
        n10602) );
  BUF_X1 U13628 ( .A(n9859), .Z(n10585) );
  NAND2_X1 U13629 ( .A1(n10585), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10573) );
  AOI21_X1 U13630 ( .B1(n16491), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10572) );
  INV_X1 U13631 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n10580) );
  NAND2_X1 U13632 ( .A1(n10588), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10579) );
  INV_X1 U13633 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n10576) );
  NAND2_X1 U13634 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10575) );
  INV_X1 U13635 ( .A(n10577), .ZN(n10578) );
  NAND2_X1 U13636 ( .A1(n10593), .A2(n10582), .ZN(n10581) );
  INV_X1 U13637 ( .A(n10593), .ZN(n10583) );
  NAND2_X1 U13638 ( .A1(n10583), .A2(n10594), .ZN(n10584) );
  NAND2_X1 U13639 ( .A1(n10585), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10587) );
  OR2_X1 U13640 ( .A1(n16478), .A2(n20140), .ZN(n10586) );
  AOI22_X1 U13641 ( .A1(n14254), .A2(P2_EBX_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10592) );
  NAND2_X1 U13642 ( .A1(n10588), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10591) );
  NAND2_X1 U13643 ( .A1(n14255), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n10590) );
  XNOR2_X2 U13644 ( .A(n11117), .B(n11116), .ZN(n11119) );
  NAND2_X1 U13646 ( .A1(n10604), .A2(n10600), .ZN(n10601) );
  INV_X1 U13647 ( .A(n10604), .ZN(n10605) );
  INV_X1 U13648 ( .A(n10626), .ZN(n10606) );
  NOR2_X2 U13649 ( .A1(n10625), .A2(n10606), .ZN(n10707) );
  AND2_X2 U13650 ( .A1(n9833), .A2(n14942), .ZN(n10617) );
  INV_X1 U13651 ( .A(n10607), .ZN(n10609) );
  INV_X1 U13652 ( .A(n10619), .ZN(n10610) );
  AOI22_X1 U13653 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10707), .B1(
        n10716), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10615) );
  NOR2_X1 U13654 ( .A1(n10625), .A2(n10619), .ZN(n10715) );
  AND2_X2 U13655 ( .A1(n10620), .A2(n10610), .ZN(n10817) );
  AOI22_X1 U13656 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10715), .B1(
        n10817), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10614) );
  INV_X1 U13657 ( .A(n19227), .ZN(n13592) );
  NAND2_X1 U13658 ( .A1(n13089), .A2(n10600), .ZN(n10624) );
  INV_X1 U13659 ( .A(n10624), .ZN(n10611) );
  AND2_X2 U13660 ( .A1(n10620), .A2(n10611), .ZN(n10818) );
  AOI22_X1 U13661 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19739), .B1(
        n10818), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10613) );
  AOI22_X1 U13662 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n10708), .B1(
        n10823), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10612) );
  NOR2_X2 U13663 ( .A1(n10625), .A2(n10618), .ZN(n19607) );
  AOI22_X1 U13664 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19607), .B1(
        n19863), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10623) );
  NOR2_X1 U13665 ( .A1(n10627), .A2(n10619), .ZN(n10713) );
  AOI22_X1 U13666 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10706), .B1(
        n10713), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10622) );
  NOR2_X2 U13667 ( .A1(n10627), .A2(n10624), .ZN(n19494) );
  AOI22_X1 U13668 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19494), .B1(
        n10714), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10621) );
  NOR2_X2 U13669 ( .A1(n10625), .A2(n10624), .ZN(n10705) );
  INV_X1 U13670 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13127) );
  NOR2_X1 U13671 ( .A1(n9895), .A2(n10628), .ZN(n10629) );
  NAND3_X1 U13672 ( .A1(n10631), .A2(n10630), .A3(n10629), .ZN(n10677) );
  AND2_X2 U13673 ( .A1(n9838), .A2(n10444), .ZN(n10688) );
  AND2_X2 U13674 ( .A1(n9838), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10689) );
  AOI22_X1 U13675 ( .A1(n10688), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10689), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10638) );
  AND2_X2 U13676 ( .A1(n9841), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10650) );
  AND2_X2 U13677 ( .A1(n10634), .A2(n10444), .ZN(n13187) );
  AOI22_X1 U13678 ( .A1(n10650), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13187), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10637) );
  AND2_X2 U13679 ( .A1(n13391), .A2(n10444), .ZN(n13218) );
  AND2_X2 U13680 ( .A1(n9815), .A2(n10444), .ZN(n13219) );
  AOI22_X1 U13681 ( .A1(n13218), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13219), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10636) );
  AND2_X1 U13682 ( .A1(n10634), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10649) );
  AOI22_X1 U13683 ( .A1(n13220), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10649), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10635) );
  NAND4_X1 U13684 ( .A1(n10638), .A2(n10637), .A3(n10636), .A4(n10635), .ZN(
        n10648) );
  NAND2_X1 U13685 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13201) );
  INV_X1 U13686 ( .A(n13201), .ZN(n10999) );
  INV_X1 U13687 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n19936) );
  INV_X1 U13688 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n19446) );
  OAI22_X1 U13689 ( .A1(n13178), .A2(n19936), .B1(n13177), .B2(n19446), .ZN(
        n10640) );
  INV_X1 U13690 ( .A(n10640), .ZN(n10646) );
  AND2_X2 U13691 ( .A1(n9834), .A2(n10444), .ZN(n13225) );
  AND2_X2 U13692 ( .A1(n9834), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13226) );
  AOI22_X1 U13693 ( .A1(n13225), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13226), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10645) );
  AOI22_X1 U13694 ( .A1(n10728), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10748), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10642) );
  NAND2_X1 U13695 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n10641) );
  NAND3_X1 U13696 ( .A1(n10646), .A2(n10645), .A3(n10644), .ZN(n10647) );
  INV_X1 U13697 ( .A(n11221), .ZN(n10661) );
  INV_X1 U13698 ( .A(n13177), .ZN(n13228) );
  AOI22_X1 U13699 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n13228), .ZN(n10654) );
  AOI22_X1 U13700 ( .A1(n13220), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13217), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10653) );
  AOI22_X1 U13701 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n13218), .B1(
        n10650), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10652) );
  AOI22_X1 U13702 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n13219), .B1(
        n13226), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10651) );
  NAND4_X1 U13703 ( .A1(n10654), .A2(n10653), .A3(n10652), .A4(n10651), .ZN(
        n10660) );
  AOI22_X1 U13704 ( .A1(n10688), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n10728), .ZN(n10658) );
  INV_X1 U13705 ( .A(n13178), .ZN(n13227) );
  AOI22_X1 U13706 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n13187), .B1(
        n13227), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10657) );
  AOI22_X1 U13707 ( .A1(n10689), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n10748), .ZN(n10656) );
  AOI22_X1 U13708 ( .A1(n10694), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n13225), .ZN(n10655) );
  NAND4_X1 U13709 ( .A1(n10658), .A2(n10657), .A3(n10656), .A4(n10655), .ZN(
        n10659) );
  NOR2_X1 U13710 ( .A1(n10661), .A2(n11231), .ZN(n10662) );
  NAND2_X1 U13711 ( .A1(n10536), .A2(n10662), .ZN(n11052) );
  INV_X1 U13712 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10663) );
  OAI22_X1 U13713 ( .A1(n13178), .A2(n10663), .B1(n13177), .B2(n19457), .ZN(
        n10664) );
  AOI21_X1 U13714 ( .B1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B2(n10694), .A(
        n10664), .ZN(n10669) );
  AOI22_X1 U13715 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10728), .B1(
        n10748), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10668) );
  AOI22_X1 U13716 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n13225), .B1(
        n13226), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10667) );
  NAND2_X1 U13717 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n10666) );
  NAND4_X1 U13718 ( .A1(n10669), .A2(n10668), .A3(n10667), .A4(n10666), .ZN(
        n10675) );
  AOI22_X1 U13719 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10688), .B1(
        n10689), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10673) );
  AOI22_X1 U13720 ( .A1(n10650), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13187), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10672) );
  AOI22_X1 U13721 ( .A1(n13218), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13219), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10671) );
  AOI22_X1 U13722 ( .A1(n13220), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13217), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10670) );
  NAND4_X1 U13723 ( .A1(n10673), .A2(n10672), .A3(n10671), .A4(n10670), .ZN(
        n10674) );
  NAND2_X1 U13724 ( .A1(n11052), .A2(n11051), .ZN(n10676) );
  INV_X1 U13725 ( .A(n10678), .ZN(n10703) );
  AOI22_X1 U13726 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10713), .B1(
        n19739), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10681) );
  AOI22_X1 U13727 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10706), .B1(
        n19494), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10680) );
  AOI22_X1 U13728 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10715), .B1(
        n10707), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10686) );
  AOI22_X1 U13729 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19607), .B1(
        n10714), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10685) );
  AOI22_X1 U13730 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10705), .B1(
        n10708), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10684) );
  AOI22_X1 U13731 ( .A1(n10688), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10689), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10693) );
  AOI22_X1 U13732 ( .A1(n10650), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13187), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10692) );
  AOI22_X1 U13733 ( .A1(n13218), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13219), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10691) );
  AOI22_X1 U13734 ( .A1(n13220), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13217), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10690) );
  NAND4_X1 U13735 ( .A1(n10693), .A2(n10692), .A3(n10691), .A4(n10690), .ZN(
        n10702) );
  OAI22_X1 U13736 ( .A1(n13178), .A2(n10695), .B1(n13177), .B2(n19468), .ZN(
        n10696) );
  AOI21_X1 U13737 ( .B1(n10694), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A(
        n10696), .ZN(n10700) );
  AOI22_X1 U13738 ( .A1(n10728), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10748), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10699) );
  AOI22_X1 U13739 ( .A1(n13225), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13226), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10698) );
  NAND2_X1 U13740 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10697) );
  NAND4_X1 U13741 ( .A1(n10700), .A2(n10699), .A3(n10698), .A4(n10697), .ZN(
        n10701) );
  AND2_X1 U13742 ( .A1(n10818), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10704) );
  AOI22_X1 U13743 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n10705), .B1(
        n19607), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10711) );
  AOI22_X1 U13744 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19440), .B1(
        n19494), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10710) );
  AOI22_X1 U13745 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n10707), .B1(
        n10708), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10709) );
  AOI22_X1 U13746 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19582), .B1(
        n19739), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10721) );
  AOI22_X1 U13747 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19798), .B1(
        n19863), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10720) );
  AOI22_X1 U13748 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19702), .B1(
        n10716), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10719) );
  INV_X1 U13749 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10718) );
  INV_X1 U13750 ( .A(n10817), .ZN(n10717) );
  AOI22_X1 U13751 ( .A1(n10650), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13220), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10726) );
  AOI22_X1 U13752 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10688), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10725) );
  AOI22_X1 U13753 ( .A1(n13218), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10694), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10724) );
  AOI22_X1 U13754 ( .A1(n13217), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13219), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10723) );
  NAND4_X1 U13755 ( .A1(n10726), .A2(n10725), .A3(n10724), .A4(n10723), .ZN(
        n10734) );
  INV_X1 U13756 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13871) );
  OAI22_X1 U13757 ( .A1(n13178), .A2(n19953), .B1(n13177), .B2(n13871), .ZN(
        n10727) );
  AOI21_X1 U13758 ( .B1(n13187), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A(
        n10727), .ZN(n10732) );
  AOI22_X1 U13759 ( .A1(n10728), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13226), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10731) );
  AOI22_X1 U13760 ( .A1(n13225), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10748), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10730) );
  NAND2_X1 U13761 ( .A1(n10689), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10729) );
  NAND4_X1 U13762 ( .A1(n10732), .A2(n10731), .A3(n10730), .A4(n10729), .ZN(
        n10733) );
  NOR2_X1 U13763 ( .A1(n10734), .A2(n10733), .ZN(n11254) );
  NAND2_X1 U13764 ( .A1(n10650), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10738) );
  NAND2_X1 U13765 ( .A1(n10694), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10737) );
  NAND2_X1 U13766 ( .A1(n13218), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10736) );
  NAND2_X1 U13767 ( .A1(n13217), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10735) );
  NAND2_X1 U13768 ( .A1(n10688), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10742) );
  NAND2_X1 U13769 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10741) );
  NAND2_X1 U13770 ( .A1(n13220), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10740) );
  NAND2_X1 U13771 ( .A1(n13219), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10739) );
  NAND2_X1 U13772 ( .A1(n10689), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10745) );
  NAND2_X1 U13773 ( .A1(n10728), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10744) );
  NAND2_X1 U13774 ( .A1(n13225), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10743) );
  INV_X1 U13775 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10746) );
  INV_X1 U13776 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13105) );
  OAI22_X1 U13777 ( .A1(n13178), .A2(n10746), .B1(n13177), .B2(n13105), .ZN(
        n10747) );
  INV_X1 U13778 ( .A(n10747), .ZN(n10752) );
  NAND2_X1 U13779 ( .A1(n10748), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10751) );
  NAND2_X1 U13780 ( .A1(n13226), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10750) );
  NAND2_X1 U13781 ( .A1(n13187), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10749) );
  AND4_X2 U13782 ( .A1(n10756), .A2(n10755), .A3(n10754), .A4(n10753), .ZN(
        n10858) );
  OR2_X1 U13783 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(
        n10758) );
  MUX2_X1 U13784 ( .A(n16450), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        n15662), .Z(n11006) );
  NOR2_X1 U13785 ( .A1(n15651), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10761) );
  INV_X1 U13786 ( .A(n10781), .ZN(n10763) );
  XNOR2_X1 U13787 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n10762) );
  XNOR2_X1 U13788 ( .A(n10763), .B(n10762), .ZN(n10993) );
  INV_X1 U13789 ( .A(n10993), .ZN(n10764) );
  NAND2_X1 U13790 ( .A1(n14159), .A2(n10764), .ZN(n11004) );
  OAI21_X1 U13791 ( .B1(n11051), .B2(n14159), .A(n10374), .ZN(n10766) );
  AOI22_X1 U13792 ( .A1(n10688), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10689), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10770) );
  AOI22_X1 U13793 ( .A1(n10650), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13187), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10769) );
  AOI22_X1 U13794 ( .A1(n13218), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13219), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10768) );
  AOI22_X1 U13795 ( .A1(n13220), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13217), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10767) );
  NAND4_X1 U13796 ( .A1(n10770), .A2(n10769), .A3(n10768), .A4(n10767), .ZN(
        n10778) );
  INV_X1 U13797 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10771) );
  OAI22_X1 U13798 ( .A1(n13178), .A2(n10771), .B1(n13177), .B2(n19462), .ZN(
        n10772) );
  AOI21_X1 U13799 ( .B1(n10694), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A(
        n10772), .ZN(n10776) );
  AOI22_X1 U13800 ( .A1(n10728), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10748), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10775) );
  AOI22_X1 U13801 ( .A1(n13225), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13226), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10774) );
  NAND2_X1 U13802 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n10773) );
  NAND4_X1 U13803 ( .A1(n10776), .A2(n10775), .A3(n10774), .A4(n10773), .ZN(
        n10777) );
  NAND2_X1 U13804 ( .A1(n20147), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10780) );
  NOR2_X1 U13805 ( .A1(n10783), .A2(n10782), .ZN(n10784) );
  INV_X1 U13806 ( .A(n10994), .ZN(n10785) );
  MUX2_X1 U13807 ( .A(n11245), .B(n10785), .S(n14159), .Z(n10982) );
  INV_X1 U13808 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n14164) );
  MUX2_X1 U13809 ( .A(n10982), .B(n14164), .S(n19470), .Z(n10797) );
  NAND3_X1 U13810 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n10971), .A3(
        n13676), .ZN(n10996) );
  MUX2_X1 U13811 ( .A(n10996), .B(n11250), .S(n20169), .Z(n10787) );
  INV_X1 U13812 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n19292) );
  MUX2_X1 U13813 ( .A(n10787), .B(n19292), .S(n19470), .Z(n10813) );
  MUX2_X1 U13814 ( .A(n11254), .B(P2_EBX_REG_5__SCAN_IN), .S(n19470), .Z(
        n10788) );
  NAND2_X1 U13815 ( .A1(n10812), .A2(n10788), .ZN(n10789) );
  NAND2_X1 U13816 ( .A1(n10225), .A2(n10789), .ZN(n19189) );
  INV_X1 U13817 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15629) );
  XNOR2_X1 U13818 ( .A(n10814), .B(n15629), .ZN(n15310) );
  INV_X1 U13819 ( .A(n10790), .ZN(n10793) );
  INV_X1 U13820 ( .A(n10791), .ZN(n10792) );
  NAND2_X1 U13821 ( .A1(n10793), .A2(n10792), .ZN(n10794) );
  NAND2_X1 U13822 ( .A1(n11057), .A2(n10794), .ZN(n14076) );
  INV_X1 U13823 ( .A(n10795), .ZN(n10796) );
  OAI21_X1 U13824 ( .B1(n10797), .B2(n10801), .A(n10796), .ZN(n14161) );
  AND2_X1 U13825 ( .A1(n10053), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10798) );
  NOR2_X1 U13826 ( .A1(n10975), .A2(n10798), .ZN(n10976) );
  MUX2_X1 U13827 ( .A(n11221), .B(n10976), .S(n14159), .Z(n11007) );
  MUX2_X1 U13828 ( .A(n11007), .B(P2_EBX_REG_0__SCAN_IN), .S(n19470), .Z(
        n19240) );
  NAND2_X1 U13829 ( .A1(n19240), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13546) );
  INV_X1 U13830 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n13593) );
  NAND3_X1 U13831 ( .A1(n19470), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n10799) );
  NAND2_X1 U13832 ( .A1(n10803), .A2(n10799), .ZN(n19221) );
  NOR2_X1 U13833 ( .A1(n13546), .A2(n19221), .ZN(n10800) );
  NAND2_X1 U13834 ( .A1(n13546), .A2(n19221), .ZN(n13545) );
  OAI21_X1 U13835 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n10800), .A(
        n13545), .ZN(n13596) );
  INV_X1 U13836 ( .A(n10801), .ZN(n10805) );
  NAND2_X1 U13837 ( .A1(n10803), .A2(n10802), .ZN(n10804) );
  NAND2_X1 U13838 ( .A1(n10805), .A2(n10804), .ZN(n10807) );
  INV_X1 U13839 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10806) );
  XNOR2_X1 U13840 ( .A(n10807), .B(n10806), .ZN(n13595) );
  OR2_X1 U13841 ( .A1(n13596), .A2(n13595), .ZN(n13735) );
  INV_X1 U13842 ( .A(n10807), .ZN(n14939) );
  NAND2_X1 U13843 ( .A1(n14939), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10808) );
  NAND2_X1 U13844 ( .A1(n13735), .A2(n10808), .ZN(n10809) );
  AND2_X1 U13845 ( .A1(n10809), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10811) );
  INV_X1 U13846 ( .A(n10809), .ZN(n14074) );
  INV_X1 U13847 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14073) );
  NAND2_X1 U13848 ( .A1(n14074), .A2(n14073), .ZN(n10810) );
  OAI21_X1 U13849 ( .B1(n10795), .B2(n10813), .A(n10812), .ZN(n19205) );
  INV_X1 U13850 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15622) );
  XNOR2_X1 U13851 ( .A(n19205), .B(n15622), .ZN(n14102) );
  NAND2_X1 U13852 ( .A1(n15310), .A2(n15311), .ZN(n10816) );
  NAND2_X1 U13853 ( .A1(n10814), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10815) );
  NAND2_X1 U13854 ( .A1(n10816), .A2(n10815), .ZN(n15616) );
  INV_X1 U13855 ( .A(n10847), .ZN(n10846) );
  AOI22_X1 U13856 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10703), .B1(
        n10817), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10822) );
  AOI22_X1 U13857 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19440), .B1(
        n10818), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10821) );
  AOI22_X1 U13858 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n10716), .B1(
        n19863), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10820) );
  AOI22_X1 U13859 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19702), .B1(
        n10708), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10819) );
  NAND4_X1 U13860 ( .A1(n10822), .A2(n10821), .A3(n10820), .A4(n10819), .ZN(
        n10829) );
  AOI22_X1 U13861 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10707), .B1(
        n10705), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10827) );
  AOI22_X1 U13862 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19582), .B1(
        n19739), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10826) );
  AOI22_X1 U13863 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19494), .B1(
        n10823), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10825) );
  AOI22_X1 U13864 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19607), .B1(
        n19798), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10824) );
  NAND4_X1 U13865 ( .A1(n10827), .A2(n10826), .A3(n10825), .A4(n10824), .ZN(
        n10828) );
  AOI22_X1 U13866 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10688), .B1(
        n10689), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10833) );
  AOI22_X1 U13867 ( .A1(n10650), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13187), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10832) );
  AOI22_X1 U13868 ( .A1(n13218), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13219), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10831) );
  AOI22_X1 U13869 ( .A1(n13220), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13217), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10830) );
  NAND4_X1 U13870 ( .A1(n10833), .A2(n10832), .A3(n10831), .A4(n10830), .ZN(
        n10841) );
  INV_X1 U13871 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10834) );
  INV_X1 U13872 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19479) );
  OAI22_X1 U13873 ( .A1(n13178), .A2(n10834), .B1(n13177), .B2(n19479), .ZN(
        n10835) );
  AOI21_X1 U13874 ( .B1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B2(n10694), .A(
        n10835), .ZN(n10839) );
  AOI22_X1 U13875 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10728), .B1(
        n10748), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10838) );
  AOI22_X1 U13876 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n13225), .B1(
        n13226), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10837) );
  NAND2_X1 U13877 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n10836) );
  NAND4_X1 U13878 ( .A1(n10839), .A2(n10838), .A3(n10837), .A4(n10836), .ZN(
        n10840) );
  INV_X1 U13879 ( .A(n11258), .ZN(n10842) );
  NAND2_X1 U13880 ( .A1(n10842), .A2(n10527), .ZN(n10843) );
  NAND2_X1 U13881 ( .A1(n10846), .A2(n10845), .ZN(n11074) );
  NAND2_X1 U13882 ( .A1(n10847), .A2(n11066), .ZN(n10848) );
  NAND2_X1 U13883 ( .A1(n11074), .A2(n10848), .ZN(n11064) );
  INV_X1 U13884 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n13878) );
  MUX2_X1 U13885 ( .A(n11258), .B(n13878), .S(n19470), .Z(n10849) );
  NOR2_X1 U13886 ( .A1(n10850), .A2(n10849), .ZN(n10851) );
  OR2_X1 U13887 ( .A1(n9931), .A2(n10851), .ZN(n19178) );
  INV_X1 U13888 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16392) );
  XNOR2_X1 U13889 ( .A(n10852), .B(n16392), .ZN(n15617) );
  NAND2_X1 U13890 ( .A1(n15616), .A2(n15617), .ZN(n16346) );
  NAND2_X1 U13891 ( .A1(n10852), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16345) );
  INV_X1 U13892 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n10853) );
  MUX2_X1 U13893 ( .A(n14246), .B(n10853), .S(n19470), .Z(n10855) );
  INV_X1 U13894 ( .A(n10855), .ZN(n10854) );
  XNOR2_X1 U13895 ( .A(n9931), .B(n10854), .ZN(n19169) );
  NAND2_X1 U13896 ( .A1(n19169), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16357) );
  NAND2_X1 U13897 ( .A1(n10867), .A2(n10856), .ZN(n10857) );
  NAND2_X1 U13898 ( .A1(n10864), .A2(n10857), .ZN(n14926) );
  NOR2_X1 U13899 ( .A1(n14926), .A2(n10858), .ZN(n10859) );
  NAND2_X1 U13900 ( .A1(n10859), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16344) );
  AND3_X1 U13901 ( .A1(n16345), .A2(n16357), .A3(n16344), .ZN(n10862) );
  INV_X1 U13902 ( .A(n10859), .ZN(n10860) );
  INV_X1 U13903 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16395) );
  NAND2_X1 U13904 ( .A1(n10860), .A2(n16395), .ZN(n16343) );
  INV_X1 U13905 ( .A(n19169), .ZN(n10861) );
  INV_X1 U13906 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11076) );
  NAND2_X1 U13907 ( .A1(n10861), .A2(n11076), .ZN(n16358) );
  AND2_X1 U13908 ( .A1(n19470), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10863) );
  MUX2_X1 U13909 ( .A(n11219), .B(n10863), .S(n10864), .Z(n10865) );
  NOR2_X1 U13910 ( .A1(n10865), .A2(n10871), .ZN(n19152) );
  NAND2_X1 U13911 ( .A1(n19152), .A2(n14246), .ZN(n10866) );
  NAND2_X1 U13912 ( .A1(n10866), .A2(n15596), .ZN(n15592) );
  INV_X1 U13913 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n19281) );
  NOR2_X1 U13914 ( .A1(n10871), .A2(n19281), .ZN(n10868) );
  NAND2_X1 U13915 ( .A1(n19470), .A2(n10868), .ZN(n10869) );
  NAND2_X1 U13916 ( .A1(n10952), .A2(n10869), .ZN(n10870) );
  AOI21_X1 U13917 ( .B1(n10871), .B2(n19281), .A(n10870), .ZN(n19145) );
  AOI21_X1 U13918 ( .B1(n19145), .B2(n14246), .A(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16321) );
  INV_X1 U13919 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n19129) );
  INV_X1 U13920 ( .A(n10872), .ZN(n10873) );
  AND3_X1 U13921 ( .A1(n19470), .A2(P2_EBX_REG_11__SCAN_IN), .A3(n10873), .ZN(
        n10874) );
  NOR2_X1 U13922 ( .A1(n10882), .A2(n10874), .ZN(n19128) );
  AOI21_X1 U13923 ( .B1(n19128), .B2(n14246), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15575) );
  INV_X1 U13924 ( .A(n15575), .ZN(n10875) );
  AND2_X1 U13925 ( .A1(n14246), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10876) );
  NAND2_X1 U13926 ( .A1(n19152), .A2(n10876), .ZN(n16318) );
  AND2_X1 U13927 ( .A1(n14246), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10877) );
  NAND2_X1 U13928 ( .A1(n19128), .A2(n10877), .ZN(n15573) );
  INV_X1 U13929 ( .A(n19145), .ZN(n10879) );
  NAND2_X1 U13930 ( .A1(n14246), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10878) );
  AND3_X1 U13931 ( .A1(n16318), .A2(n15573), .A3(n16319), .ZN(n10880) );
  NAND2_X1 U13932 ( .A1(n19470), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10881) );
  NAND3_X1 U13933 ( .A1(n19470), .A2(n10883), .A3(P2_EBX_REG_12__SCAN_IN), 
        .ZN(n10884) );
  AND2_X1 U13934 ( .A1(n10886), .A2(n10884), .ZN(n19122) );
  NAND2_X1 U13935 ( .A1(n19122), .A2(n14246), .ZN(n15300) );
  INV_X1 U13936 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15546) );
  AND2_X1 U13937 ( .A1(n10886), .A2(n10885), .ZN(n10887) );
  OR2_X1 U13938 ( .A1(n10887), .A2(n9889), .ZN(n19108) );
  INV_X1 U13939 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15545) );
  OAI21_X1 U13940 ( .B1(n19108), .B2(n10858), .A(n15545), .ZN(n15292) );
  NAND2_X1 U13941 ( .A1(n10897), .A2(n9946), .ZN(n10907) );
  NAND2_X1 U13942 ( .A1(n19470), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10891) );
  AND3_X1 U13943 ( .A1(n10888), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n19470), .ZN(
        n10889) );
  NOR2_X1 U13944 ( .A1(n10929), .A2(n10889), .ZN(n14896) );
  AOI21_X1 U13945 ( .B1(n14896), .B2(n14246), .A(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15212) );
  INV_X1 U13946 ( .A(n15212), .ZN(n10911) );
  XNOR2_X1 U13947 ( .A(n10893), .B(n9955), .ZN(n19053) );
  NOR2_X1 U13948 ( .A1(n10919), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15247) );
  NOR2_X1 U13949 ( .A1(n10890), .A2(n10891), .ZN(n10892) );
  OR2_X1 U13950 ( .A1(n10893), .A2(n10892), .ZN(n19065) );
  INV_X1 U13951 ( .A(n19065), .ZN(n10894) );
  AOI21_X1 U13952 ( .B1(n10894), .B2(n14246), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15258) );
  NOR2_X1 U13953 ( .A1(n15247), .A2(n15258), .ZN(n15233) );
  NAND2_X1 U13954 ( .A1(n19470), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10895) );
  XNOR2_X1 U13955 ( .A(n10896), .B(n10895), .ZN(n19039) );
  INV_X1 U13956 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15436) );
  OAI21_X1 U13957 ( .B1(n19039), .B2(n10858), .A(n15436), .ZN(n15231) );
  NAND2_X1 U13958 ( .A1(n15233), .A2(n15231), .ZN(n15217) );
  NAND3_X1 U13959 ( .A1(n10899), .A2(P2_EBX_REG_16__SCAN_IN), .A3(n19470), 
        .ZN(n10898) );
  OAI211_X1 U13960 ( .C1(n10899), .C2(P2_EBX_REG_16__SCAN_IN), .A(n10898), .B(
        n10952), .ZN(n14908) );
  OR2_X1 U13961 ( .A1(n14908), .A2(n10858), .ZN(n10901) );
  INV_X1 U13962 ( .A(n10901), .ZN(n10900) );
  NAND2_X1 U13963 ( .A1(n10900), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15273) );
  INV_X1 U13964 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15501) );
  NAND2_X1 U13965 ( .A1(n10901), .A2(n15501), .ZN(n10902) );
  XNOR2_X1 U13966 ( .A(n10903), .B(n9962), .ZN(n19089) );
  NAND2_X1 U13967 ( .A1(n19089), .A2(n14246), .ZN(n10904) );
  INV_X1 U13968 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15482) );
  NAND2_X1 U13969 ( .A1(n10904), .A2(n15482), .ZN(n15504) );
  XNOR2_X1 U13970 ( .A(n9889), .B(n9956), .ZN(n19100) );
  NAND2_X1 U13971 ( .A1(n19100), .A2(n14246), .ZN(n10905) );
  INV_X1 U13972 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15518) );
  NAND2_X1 U13973 ( .A1(n10905), .A2(n15518), .ZN(n15534) );
  AND2_X1 U13974 ( .A1(n10907), .A2(n10906), .ZN(n10908) );
  OR2_X1 U13975 ( .A1(n10908), .A2(n10890), .ZN(n19078) );
  INV_X1 U13976 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15483) );
  OAI21_X1 U13977 ( .B1(n19078), .B2(n10858), .A(n15483), .ZN(n15272) );
  NAND4_X1 U13978 ( .A1(n15286), .A2(n15504), .A3(n15534), .A4(n15272), .ZN(
        n10909) );
  NOR2_X1 U13979 ( .A1(n15217), .A2(n10909), .ZN(n10910) );
  NAND2_X1 U13980 ( .A1(n10911), .A2(n10910), .ZN(n10912) );
  NAND2_X1 U13981 ( .A1(n14246), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10913) );
  NOR2_X1 U13982 ( .A1(n19065), .A2(n10913), .ZN(n15257) );
  INV_X1 U13983 ( .A(n19089), .ZN(n10914) );
  INV_X1 U13984 ( .A(n19100), .ZN(n10915) );
  INV_X1 U13985 ( .A(n19108), .ZN(n10917) );
  AND2_X1 U13986 ( .A1(n14246), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10916) );
  NAND2_X1 U13987 ( .A1(n10917), .A2(n10916), .ZN(n15291) );
  NAND3_X1 U13988 ( .A1(n15503), .A2(n15533), .A3(n15291), .ZN(n10918) );
  NOR2_X1 U13989 ( .A1(n15257), .A2(n10918), .ZN(n10923) );
  INV_X1 U13990 ( .A(n10919), .ZN(n10920) );
  INV_X1 U13991 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15251) );
  INV_X1 U13992 ( .A(n19078), .ZN(n10922) );
  AND2_X1 U13993 ( .A1(n14246), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10921) );
  NAND2_X1 U13994 ( .A1(n10922), .A2(n10921), .ZN(n15271) );
  AND2_X1 U13995 ( .A1(n15271), .A2(n15273), .ZN(n15216) );
  NAND3_X1 U13996 ( .A1(n10923), .A2(n15245), .A3(n15216), .ZN(n10926) );
  INV_X1 U13997 ( .A(n19039), .ZN(n10925) );
  AND2_X1 U13998 ( .A1(n14246), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10924) );
  AND2_X1 U13999 ( .A1(n14246), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10927) );
  AND2_X1 U14000 ( .A1(n14896), .A2(n10927), .ZN(n15211) );
  INV_X1 U14001 ( .A(n15211), .ZN(n10928) );
  NAND2_X1 U14002 ( .A1(n19470), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10930) );
  INV_X1 U14003 ( .A(n10930), .ZN(n10931) );
  NAND2_X1 U14004 ( .A1(n10932), .A2(n10931), .ZN(n10933) );
  AND2_X1 U14005 ( .A1(n10935), .A2(n10933), .ZN(n15791) );
  AOI21_X1 U14006 ( .B1(n15791), .B2(n14246), .A(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15199) );
  NAND3_X1 U14007 ( .A1(n15791), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n14246), .ZN(n15200) );
  AND2_X1 U14008 ( .A1(n10935), .A2(n10934), .ZN(n10936) );
  NOR2_X1 U14009 ( .A1(n10945), .A2(n10936), .ZN(n16248) );
  NAND2_X1 U14010 ( .A1(n16248), .A2(n14246), .ZN(n10937) );
  XNOR2_X1 U14011 ( .A(n10937), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15188) );
  INV_X1 U14012 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15395) );
  NOR2_X1 U14013 ( .A1(n10858), .A2(n15395), .ZN(n10938) );
  AOI21_X1 U14014 ( .B1(n15187), .B2(n15188), .A(n10939), .ZN(n15176) );
  NAND2_X1 U14015 ( .A1(n19470), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10940) );
  MUX2_X1 U14016 ( .A(n10940), .B(P2_EBX_REG_24__SCAN_IN), .S(n10945), .Z(
        n10941) );
  NAND2_X1 U14017 ( .A1(n10941), .A2(n10952), .ZN(n16235) );
  AOI21_X1 U14018 ( .B1(n10942), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15178), .ZN(n10944) );
  INV_X1 U14019 ( .A(n15176), .ZN(n10942) );
  NOR2_X1 U14020 ( .A1(n10942), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10943) );
  INV_X1 U14021 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n14999) );
  INV_X1 U14022 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n16222) );
  NAND3_X1 U14023 ( .A1(n19470), .A2(P2_EBX_REG_26__SCAN_IN), .A3(n9894), .ZN(
        n10946) );
  NAND2_X1 U14024 ( .A1(n14245), .A2(n10946), .ZN(n10947) );
  INV_X1 U14025 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15359) );
  NOR3_X1 U14026 ( .A1(n10947), .A2(n10858), .A3(n15359), .ZN(n10965) );
  INV_X1 U14027 ( .A(n10947), .ZN(n16212) );
  AOI21_X1 U14028 ( .B1(n16212), .B2(n14246), .A(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10948) );
  NOR2_X1 U14029 ( .A1(n10965), .A2(n10948), .ZN(n15156) );
  INV_X1 U14030 ( .A(n15156), .ZN(n10955) );
  NOR2_X1 U14031 ( .A1(n10949), .A2(n16222), .ZN(n10950) );
  NAND2_X1 U14032 ( .A1(n19470), .A2(n10950), .ZN(n10951) );
  AND2_X1 U14033 ( .A1(n10952), .A2(n10951), .ZN(n10953) );
  NAND2_X1 U14034 ( .A1(n9894), .A2(n10953), .ZN(n16223) );
  INV_X1 U14035 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15369) );
  NAND2_X1 U14036 ( .A1(n10963), .A2(n15369), .ZN(n15165) );
  INV_X1 U14037 ( .A(n15165), .ZN(n10954) );
  NAND2_X1 U14038 ( .A1(n19470), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10958) );
  INV_X1 U14039 ( .A(n10958), .ZN(n10959) );
  NAND2_X1 U14040 ( .A1(n10959), .A2(n9886), .ZN(n10960) );
  NAND2_X1 U14041 ( .A1(n16202), .A2(n14246), .ZN(n15135) );
  INV_X1 U14042 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15148) );
  NAND2_X1 U14043 ( .A1(n19470), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n10967) );
  XOR2_X1 U14044 ( .A(n10967), .B(n10966), .Z(n16189) );
  INV_X1 U14045 ( .A(n10963), .ZN(n10964) );
  NOR2_X1 U14046 ( .A1(n15166), .A2(n10965), .ZN(n15132) );
  NAND2_X1 U14047 ( .A1(n19470), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14237) );
  INV_X1 U14048 ( .A(n10966), .ZN(n10968) );
  NAND2_X1 U14049 ( .A1(n10968), .A2(n10967), .ZN(n14236) );
  XOR2_X1 U14050 ( .A(n14237), .B(n14236), .Z(n10969) );
  INV_X1 U14051 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11426) );
  INV_X1 U14052 ( .A(n10969), .ZN(n16176) );
  NAND3_X1 U14053 ( .A1(n16176), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14246), .ZN(n15109) );
  NAND2_X1 U14054 ( .A1(n10972), .A2(n19447), .ZN(n10973) );
  NAND2_X1 U14055 ( .A1(n10973), .A2(n10993), .ZN(n10981) );
  NAND2_X1 U14056 ( .A1(n10976), .A2(n11006), .ZN(n10974) );
  NAND2_X1 U14057 ( .A1(n20169), .A2(n10974), .ZN(n10980) );
  XNOR2_X1 U14058 ( .A(n11006), .B(n10975), .ZN(n10989) );
  NAND2_X1 U14059 ( .A1(n19447), .A2(n10989), .ZN(n10978) );
  INV_X1 U14060 ( .A(n10976), .ZN(n10992) );
  OAI21_X1 U14061 ( .B1(n10989), .B2(n10992), .A(n10993), .ZN(n10977) );
  NAND3_X1 U14062 ( .A1(n10978), .A2(n11089), .A3(n10977), .ZN(n10979) );
  AOI22_X1 U14063 ( .A1(n11004), .A2(n10981), .B1(n10980), .B2(n10979), .ZN(
        n10984) );
  NAND2_X1 U14064 ( .A1(n10982), .A2(n10996), .ZN(n11008) );
  NAND2_X1 U14065 ( .A1(n11008), .A2(n14159), .ZN(n10983) );
  OAI21_X1 U14066 ( .B1(n10984), .B2(n10994), .A(n10983), .ZN(n10985) );
  OAI21_X1 U14067 ( .B1(n10996), .B2(n14159), .A(n10985), .ZN(n10986) );
  OR2_X1 U14068 ( .A1(n11011), .A2(n10986), .ZN(n10987) );
  MUX2_X1 U14069 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n10987), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n11038) );
  NAND2_X1 U14070 ( .A1(n11011), .A2(n14846), .ZN(n10988) );
  NAND2_X1 U14071 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n14851) );
  INV_X1 U14072 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19017) );
  NOR2_X1 U14073 ( .A1(n19017), .A2(n20055), .ZN(n20048) );
  NAND2_X1 U14074 ( .A1(n19017), .A2(n20055), .ZN(n20050) );
  INV_X1 U14075 ( .A(n20050), .ZN(n20036) );
  NOR3_X1 U14076 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20048), .A3(n20036), 
        .ZN(n20041) );
  INV_X1 U14077 ( .A(n20041), .ZN(n14845) );
  NOR2_X1 U14078 ( .A1(n20047), .A2(n14845), .ZN(n13663) );
  NAND3_X1 U14079 ( .A1(n13665), .A2(n13663), .A3(n11018), .ZN(n11043) );
  NOR3_X1 U14080 ( .A1(n10994), .A2(n10989), .A3(n10993), .ZN(n10990) );
  AND2_X1 U14081 ( .A1(n10996), .A2(n10990), .ZN(n10991) );
  OR2_X1 U14082 ( .A1(n11011), .A2(n10991), .ZN(n13441) );
  NOR3_X1 U14083 ( .A1(n10994), .A2(n10993), .A3(n10992), .ZN(n10995) );
  NAND2_X1 U14084 ( .A1(n10996), .A2(n10995), .ZN(n10997) );
  NAND2_X1 U14085 ( .A1(n10997), .A2(n16479), .ZN(n10998) );
  OR2_X1 U14086 ( .A1(n13441), .A2(n10998), .ZN(n11003) );
  AOI21_X1 U14087 ( .B1(n15662), .B2(n10999), .A(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13671) );
  NAND2_X1 U14088 ( .A1(n13178), .A2(n13671), .ZN(n11001) );
  INV_X1 U14089 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n11000) );
  NAND2_X1 U14090 ( .A1(n11001), .A2(n11000), .ZN(n11002) );
  NAND2_X1 U14091 ( .A1(n11002), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n20157) );
  NAND2_X1 U14092 ( .A1(n11003), .A2(n20157), .ZN(n16477) );
  NAND2_X1 U14093 ( .A1(n16477), .A2(n19447), .ZN(n11013) );
  INV_X1 U14094 ( .A(n11004), .ZN(n11005) );
  AOI21_X1 U14095 ( .B1(n11007), .B2(n11006), .A(n11005), .ZN(n11009) );
  NOR2_X1 U14096 ( .A1(n11009), .A2(n11008), .ZN(n11010) );
  OR2_X1 U14097 ( .A1(n11011), .A2(n11010), .ZN(n20167) );
  AND2_X1 U14098 ( .A1(n10536), .A2(n19437), .ZN(n20168) );
  INV_X1 U14099 ( .A(n20168), .ZN(n11046) );
  NAND2_X1 U14100 ( .A1(n11013), .A2(n11012), .ZN(n13443) );
  INV_X1 U14101 ( .A(n11015), .ZN(n16464) );
  MUX2_X1 U14102 ( .A(n11017), .B(n11018), .S(n10527), .Z(n11019) );
  NAND2_X1 U14103 ( .A1(n11019), .A2(n14851), .ZN(n11036) );
  NAND2_X1 U14104 ( .A1(n11021), .A2(n10502), .ZN(n11028) );
  NAND2_X1 U14105 ( .A1(n10536), .A2(n11022), .ZN(n11098) );
  NAND2_X1 U14106 ( .A1(n11098), .A2(n11089), .ZN(n11023) );
  NAND2_X1 U14107 ( .A1(n11024), .A2(n10502), .ZN(n11026) );
  NAND2_X1 U14108 ( .A1(n11026), .A2(n11025), .ZN(n11027) );
  AOI21_X1 U14109 ( .B1(n13674), .B2(n11028), .A(n11027), .ZN(n11102) );
  INV_X1 U14110 ( .A(n13441), .ZN(n16427) );
  AND2_X1 U14111 ( .A1(n16427), .A2(n13663), .ZN(n11029) );
  NAND2_X1 U14112 ( .A1(n11017), .A2(n11029), .ZN(n11033) );
  NAND2_X1 U14113 ( .A1(n11032), .A2(n20168), .ZN(n11100) );
  AND3_X1 U14114 ( .A1(n11034), .A2(n11033), .A3(n11100), .ZN(n11035) );
  AND2_X1 U14115 ( .A1(n11102), .A2(n11035), .ZN(n13667) );
  OAI21_X1 U14116 ( .B1(n13441), .B2(n11036), .A(n13667), .ZN(n11037) );
  AOI21_X1 U14117 ( .B1(n13443), .B2(n16464), .A(n11037), .ZN(n11042) );
  INV_X1 U14118 ( .A(n13665), .ZN(n11040) );
  AOI21_X1 U14119 ( .B1(n11038), .B2(n11089), .A(n19464), .ZN(n11039) );
  NAND2_X1 U14120 ( .A1(n11040), .A2(n11039), .ZN(n11041) );
  NAND3_X1 U14121 ( .A1(n11043), .A2(n11042), .A3(n11041), .ZN(n11044) );
  NAND2_X1 U14122 ( .A1(n16479), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15864) );
  INV_X1 U14123 ( .A(n16488), .ZN(n20027) );
  NOR2_X1 U14124 ( .A1(n11015), .A2(n14159), .ZN(n11045) );
  NOR2_X1 U14125 ( .A1(n11015), .A2(n11046), .ZN(n11047) );
  INV_X1 U14126 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n16421) );
  NOR2_X1 U14127 ( .A1(n11221), .A2(n16421), .ZN(n13534) );
  INV_X1 U14128 ( .A(n11231), .ZN(n11048) );
  NAND2_X1 U14129 ( .A1(n13534), .A2(n11048), .ZN(n11050) );
  NOR2_X1 U14130 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n11221), .ZN(
        n11049) );
  XOR2_X1 U14131 ( .A(n11231), .B(n11049), .Z(n13549) );
  NAND2_X1 U14132 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13549), .ZN(
        n13548) );
  NAND2_X1 U14133 ( .A1(n11050), .A2(n13548), .ZN(n11053) );
  XOR2_X1 U14134 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n11053), .Z(
        n13600) );
  XNOR2_X1 U14135 ( .A(n11052), .B(n11051), .ZN(n13599) );
  NAND2_X1 U14136 ( .A1(n13600), .A2(n13599), .ZN(n13598) );
  NAND2_X1 U14137 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11053), .ZN(
        n11054) );
  NAND2_X1 U14138 ( .A1(n13598), .A2(n11054), .ZN(n11055) );
  XNOR2_X1 U14139 ( .A(n11055), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14077) );
  NAND2_X1 U14140 ( .A1(n11055), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11056) );
  OAI21_X1 U14141 ( .B1(n14076), .B2(n14077), .A(n11056), .ZN(n11058) );
  XNOR2_X1 U14142 ( .A(n11057), .B(n11250), .ZN(n11059) );
  NAND2_X1 U14143 ( .A1(n11058), .A2(n11059), .ZN(n14114) );
  NAND2_X1 U14144 ( .A1(n14114), .A2(n15622), .ZN(n11062) );
  NAND2_X1 U14145 ( .A1(n11063), .A2(n15629), .ZN(n15313) );
  NAND2_X1 U14146 ( .A1(n15316), .A2(n15313), .ZN(n11070) );
  INV_X1 U14147 ( .A(n11064), .ZN(n11071) );
  NAND2_X1 U14148 ( .A1(n11065), .A2(n11070), .ZN(n11069) );
  INV_X1 U14149 ( .A(n15314), .ZN(n11067) );
  NAND2_X1 U14150 ( .A1(n11067), .A2(n11066), .ZN(n11068) );
  NAND2_X1 U14151 ( .A1(n15607), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15606) );
  NAND2_X1 U14152 ( .A1(n11070), .A2(n15314), .ZN(n11072) );
  NAND2_X1 U14153 ( .A1(n11072), .A2(n11071), .ZN(n11073) );
  NAND2_X1 U14154 ( .A1(n11074), .A2(n10858), .ZN(n11075) );
  NAND2_X1 U14155 ( .A1(n11078), .A2(n11075), .ZN(n16352) );
  XNOR2_X1 U14156 ( .A(n11078), .B(n16395), .ZN(n16342) );
  INV_X1 U14157 ( .A(n11078), .ZN(n11079) );
  AND3_X1 U14158 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15467) );
  NAND2_X1 U14159 ( .A1(n15467), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15438) );
  NOR2_X1 U14160 ( .A1(n15438), .A2(n15251), .ZN(n15437) );
  AND2_X1 U14161 ( .A1(n15437), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15389) );
  AND2_X1 U14162 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15544) );
  NAND2_X1 U14163 ( .A1(n15544), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15388) );
  AND2_X1 U14164 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15580) );
  NAND2_X1 U14165 ( .A1(n15580), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15525) );
  NOR2_X1 U14166 ( .A1(n15388), .A2(n15525), .ZN(n15478) );
  AND2_X1 U14167 ( .A1(n15389), .A2(n15478), .ZN(n15391) );
  NAND2_X1 U14168 ( .A1(n15391), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15407) );
  INV_X1 U14169 ( .A(n15407), .ZN(n15397) );
  NAND2_X1 U14170 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15356) );
  INV_X1 U14171 ( .A(n15356), .ZN(n11080) );
  INV_X1 U14172 ( .A(n15140), .ZN(n15147) );
  AOI21_X1 U14173 ( .B1(n15147), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11082) );
  NAND2_X1 U14174 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11420) );
  NOR2_X1 U14175 ( .A1(n11082), .A2(n15116), .ZN(n15129) );
  NAND2_X1 U14176 ( .A1(n11083), .A2(n19447), .ZN(n15636) );
  NAND2_X1 U14177 ( .A1(n15636), .A2(n11100), .ZN(n11084) );
  NAND2_X1 U14178 ( .A1(n11084), .A2(n19458), .ZN(n11095) );
  OAI21_X1 U14179 ( .B1(n11085), .B2(n11086), .A(n14848), .ZN(n11087) );
  NAND2_X1 U14180 ( .A1(n11087), .A2(n9820), .ZN(n11094) );
  NAND2_X1 U14181 ( .A1(n11085), .A2(n11088), .ZN(n13403) );
  OAI22_X1 U14182 ( .A1(n14848), .A2(n19464), .B1(n11089), .B2(n10502), .ZN(
        n11090) );
  INV_X1 U14183 ( .A(n11090), .ZN(n11091) );
  AND2_X1 U14184 ( .A1(n13403), .A2(n11091), .ZN(n11093) );
  NAND4_X1 U14185 ( .A1(n11095), .A2(n11094), .A3(n11093), .A4(n11092), .ZN(
        n16449) );
  OR2_X1 U14186 ( .A1(n16449), .A2(n11096), .ZN(n11097) );
  NAND2_X1 U14187 ( .A1(n11216), .A2(n11097), .ZN(n11106) );
  INV_X1 U14188 ( .A(n11106), .ZN(n15481) );
  INV_X1 U14189 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15649) );
  NOR2_X1 U14190 ( .A1(n15649), .A2(n16421), .ZN(n13724) );
  AND2_X1 U14191 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13724), .ZN(
        n13732) );
  INV_X1 U14192 ( .A(n11098), .ZN(n11099) );
  AND2_X1 U14193 ( .A1(n11100), .A2(n11099), .ZN(n11101) );
  NAND2_X1 U14194 ( .A1(n11216), .A2(n16430), .ZN(n15480) );
  INV_X1 U14195 ( .A(n15480), .ZN(n13731) );
  NOR2_X1 U14196 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13724), .ZN(
        n13733) );
  INV_X1 U14197 ( .A(n13733), .ZN(n14088) );
  AOI22_X1 U14198 ( .A1(n15481), .A2(n13732), .B1(n13731), .B2(n14088), .ZN(
        n16394) );
  INV_X1 U14199 ( .A(n16394), .ZN(n14110) );
  NAND3_X1 U14200 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16393) );
  NOR4_X1 U14201 ( .A1(n16392), .A2(n11076), .A3(n16395), .A4(n16393), .ZN(
        n11107) );
  NAND2_X1 U14202 ( .A1(n14110), .A2(n11107), .ZN(n15406) );
  NAND2_X1 U14203 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11103) );
  NOR2_X1 U14204 ( .A1(n15407), .A2(n11103), .ZN(n11110) );
  NAND2_X1 U14205 ( .A1(n15597), .A2(n11110), .ZN(n15378) );
  INV_X1 U14206 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15377) );
  NOR3_X1 U14207 ( .A1(n15378), .A2(n15356), .A3(n15377), .ZN(n15336) );
  INV_X1 U14208 ( .A(n15336), .ZN(n11422) );
  NOR2_X1 U14209 ( .A1(n11422), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15346) );
  NOR2_X1 U14210 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11106), .ZN(
        n13725) );
  INV_X1 U14211 ( .A(n11216), .ZN(n11105) );
  INV_X1 U14212 ( .A(n16478), .ZN(n11104) );
  AND2_X2 U14213 ( .A1(n11104), .A2(n20126), .ZN(n19414) );
  NAND2_X1 U14214 ( .A1(n11105), .A2(n19176), .ZN(n16417) );
  OAI21_X1 U14215 ( .B1(n11106), .B2(n13724), .A(n16417), .ZN(n15439) );
  NOR2_X1 U14216 ( .A1(n13725), .A2(n15439), .ZN(n14087) );
  NAND2_X1 U14217 ( .A1(n15480), .A2(n11106), .ZN(n16420) );
  NAND2_X1 U14218 ( .A1(n14088), .A2(n11107), .ZN(n11108) );
  NAND2_X1 U14219 ( .A1(n16420), .A2(n11108), .ZN(n11109) );
  INV_X1 U14220 ( .A(n15579), .ZN(n15595) );
  INV_X1 U14221 ( .A(n16420), .ZN(n16386) );
  OAI22_X1 U14222 ( .A1(n16386), .A2(n11110), .B1(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15378), .ZN(n11111) );
  NOR2_X1 U14223 ( .A1(n15595), .A2(n11111), .ZN(n15376) );
  NAND2_X1 U14224 ( .A1(n16420), .A2(n15356), .ZN(n11112) );
  NAND2_X1 U14225 ( .A1(n15376), .A2(n11112), .ZN(n15348) );
  NOR2_X1 U14226 ( .A1(n15346), .A2(n15348), .ZN(n15339) );
  INV_X1 U14227 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20104) );
  INV_X4 U14228 ( .A(n11113), .ZN(n14254) );
  AOI22_X1 U14229 ( .A1(n14254), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n11114) );
  OAI21_X1 U14230 ( .B1(n14253), .B2(n20104), .A(n11114), .ZN(n11115) );
  AOI21_X1 U14231 ( .B1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n14250), .A(
        n11115), .ZN(n11206) );
  INV_X1 U14232 ( .A(n11116), .ZN(n11118) );
  INV_X1 U14233 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n11123) );
  AND2_X1 U14234 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11120) );
  AOI21_X1 U14235 ( .B1(n14254), .B2(P2_EBX_REG_4__SCAN_IN), .A(n11120), .ZN(
        n11122) );
  NAND2_X1 U14236 ( .A1(n14250), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11121) );
  OAI211_X1 U14237 ( .C1(n14253), .C2(n11123), .A(n11122), .B(n11121), .ZN(
        n14106) );
  INV_X1 U14238 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n11127) );
  AND2_X1 U14239 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11124) );
  AOI21_X1 U14240 ( .B1(n14254), .B2(P2_EBX_REG_5__SCAN_IN), .A(n11124), .ZN(
        n11126) );
  NAND2_X1 U14241 ( .A1(n14250), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11125) );
  OAI211_X1 U14242 ( .C1(n14253), .C2(n11127), .A(n11126), .B(n11125), .ZN(
        n13858) );
  NAND2_X1 U14243 ( .A1(n14109), .A2(n13858), .ZN(n13857) );
  AOI22_X1 U14244 ( .A1(n14254), .A2(P2_EBX_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11130) );
  NAND2_X1 U14245 ( .A1(n14250), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11129) );
  NAND2_X1 U14246 ( .A1(n14255), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11128) );
  AOI22_X1 U14247 ( .A1(n14254), .A2(P2_EBX_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11135) );
  NAND2_X1 U14248 ( .A1(n14250), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11134) );
  NAND2_X1 U14249 ( .A1(n14255), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n11133) );
  INV_X1 U14250 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n14928) );
  AND2_X1 U14251 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11136) );
  AOI21_X1 U14252 ( .B1(n14254), .B2(P2_EBX_REG_8__SCAN_IN), .A(n11136), .ZN(
        n11138) );
  NAND2_X1 U14253 ( .A1(n14250), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11137) );
  OAI211_X1 U14254 ( .C1(n14253), .C2(n14928), .A(n11138), .B(n11137), .ZN(
        n14920) );
  INV_X1 U14255 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n11142) );
  AND2_X1 U14256 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11139) );
  AOI21_X1 U14257 ( .B1(n14254), .B2(P2_EBX_REG_9__SCAN_IN), .A(n11139), .ZN(
        n11141) );
  NAND2_X1 U14258 ( .A1(n14250), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11140) );
  OAI211_X1 U14259 ( .C1(n14253), .C2(n11142), .A(n11141), .B(n11140), .ZN(
        n13978) );
  AOI22_X1 U14260 ( .A1(n14254), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n11145) );
  NAND2_X1 U14261 ( .A1(n14250), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11144) );
  NAND2_X1 U14262 ( .A1(n14255), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11143) );
  AOI22_X1 U14263 ( .A1(n14254), .A2(P2_EBX_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11150) );
  NAND2_X1 U14264 ( .A1(n14250), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11149) );
  NAND2_X1 U14265 ( .A1(n14255), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n11148) );
  AOI22_X1 U14266 ( .A1(n14254), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n11153) );
  NAND2_X1 U14267 ( .A1(n14250), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11152) );
  NAND2_X1 U14268 ( .A1(n14255), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11151) );
  INV_X1 U14269 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n11157) );
  AND2_X1 U14270 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11154) );
  AOI21_X1 U14271 ( .B1(n14254), .B2(P2_EBX_REG_13__SCAN_IN), .A(n11154), .ZN(
        n11156) );
  NAND2_X1 U14272 ( .A1(n14250), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11155) );
  OAI211_X1 U14273 ( .C1(n14253), .C2(n11157), .A(n11156), .B(n11155), .ZN(
        n14098) );
  AOI22_X1 U14274 ( .A1(n14254), .A2(P2_EBX_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n11160) );
  NAND2_X1 U14275 ( .A1(n14250), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11159) );
  NAND2_X1 U14276 ( .A1(n14255), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11158) );
  AOI22_X1 U14277 ( .A1(n14254), .A2(P2_EBX_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n11163) );
  NAND2_X1 U14278 ( .A1(n14250), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11162) );
  NAND2_X1 U14279 ( .A1(n14255), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11161) );
  INV_X1 U14280 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n14910) );
  AND2_X1 U14281 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11164) );
  AOI21_X1 U14282 ( .B1(n14254), .B2(P2_EBX_REG_16__SCAN_IN), .A(n11164), .ZN(
        n11166) );
  NAND2_X1 U14283 ( .A1(n14250), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11165) );
  OAI211_X1 U14284 ( .C1(n14253), .C2(n14910), .A(n11166), .B(n11165), .ZN(
        n14905) );
  INV_X1 U14285 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20081) );
  AND2_X1 U14286 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11167) );
  AOI21_X1 U14287 ( .B1(n14254), .B2(P2_EBX_REG_17__SCAN_IN), .A(n11167), .ZN(
        n11169) );
  NAND2_X1 U14288 ( .A1(n14250), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11168) );
  OAI211_X1 U14289 ( .C1(n14253), .C2(n20081), .A(n11169), .B(n11168), .ZN(
        n15017) );
  AOI22_X1 U14290 ( .A1(n14254), .A2(P2_EBX_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11172) );
  NAND2_X1 U14291 ( .A1(n14250), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11171) );
  NAND2_X1 U14292 ( .A1(n14255), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11170) );
  AOI22_X1 U14293 ( .A1(n14254), .A2(P2_EBX_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n11175) );
  NAND2_X1 U14294 ( .A1(n14250), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11174) );
  NAND2_X1 U14295 ( .A1(n14255), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11173) );
  INV_X1 U14296 ( .A(n15009), .ZN(n11176) );
  INV_X1 U14297 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n11180) );
  AND2_X1 U14298 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11177) );
  AOI21_X1 U14299 ( .B1(n14254), .B2(P2_EBX_REG_20__SCAN_IN), .A(n11177), .ZN(
        n11179) );
  NAND2_X1 U14300 ( .A1(n14250), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11178) );
  OAI211_X1 U14301 ( .C1(n14253), .C2(n11180), .A(n11179), .B(n11178), .ZN(
        n15235) );
  INV_X1 U14302 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20088) );
  AND2_X1 U14303 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11181) );
  AOI21_X1 U14304 ( .B1(n14254), .B2(P2_EBX_REG_21__SCAN_IN), .A(n11181), .ZN(
        n11183) );
  NAND2_X1 U14305 ( .A1(n14250), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11182) );
  OAI211_X1 U14306 ( .C1(n14253), .C2(n20088), .A(n11183), .B(n11182), .ZN(
        n14894) );
  AOI22_X1 U14307 ( .A1(n14254), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11186) );
  NAND2_X1 U14308 ( .A1(n14250), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11185) );
  NAND2_X1 U14309 ( .A1(n14255), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11184) );
  AOI22_X1 U14310 ( .A1(n14254), .A2(P2_EBX_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n11189) );
  NAND2_X1 U14311 ( .A1(n14250), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11188) );
  NAND2_X1 U14312 ( .A1(n14255), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11187) );
  AOI22_X1 U14313 ( .A1(n14254), .A2(P2_EBX_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n11193) );
  NAND2_X1 U14314 ( .A1(n14250), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11192) );
  NAND2_X1 U14315 ( .A1(n14255), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11191) );
  INV_X1 U14316 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20096) );
  AND2_X1 U14317 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11194) );
  AOI21_X1 U14318 ( .B1(n14254), .B2(P2_EBX_REG_25__SCAN_IN), .A(n11194), .ZN(
        n11196) );
  NAND2_X1 U14319 ( .A1(n14250), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11195) );
  OAI211_X1 U14320 ( .C1(n14253), .C2(n20096), .A(n11196), .B(n11195), .ZN(
        n14987) );
  INV_X1 U14321 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20098) );
  AND2_X1 U14322 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11197) );
  AOI21_X1 U14323 ( .B1(n14254), .B2(P2_EBX_REG_26__SCAN_IN), .A(n11197), .ZN(
        n11199) );
  NAND2_X1 U14324 ( .A1(n14250), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11198) );
  OAI211_X1 U14325 ( .C1(n14253), .C2(n20098), .A(n11199), .B(n11198), .ZN(
        n14980) );
  INV_X1 U14326 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20101) );
  AND2_X1 U14327 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11200) );
  AOI21_X1 U14328 ( .B1(n14254), .B2(P2_EBX_REG_27__SCAN_IN), .A(n11200), .ZN(
        n11202) );
  NAND2_X1 U14329 ( .A1(n14250), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11201) );
  OAI211_X1 U14330 ( .C1(n14253), .C2(n20101), .A(n11202), .B(n11201), .ZN(
        n14969) );
  AOI22_X1 U14331 ( .A1(n14254), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n11205) );
  NAND2_X1 U14332 ( .A1(n14250), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11204) );
  NAND2_X1 U14333 ( .A1(n14255), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11203) );
  AOI21_X1 U14334 ( .B1(n11206), .B2(n14961), .A(n14947), .ZN(n16178) );
  INV_X1 U14335 ( .A(n15661), .ZN(n11210) );
  AND2_X1 U14336 ( .A1(n11207), .A2(n13674), .ZN(n11208) );
  NAND2_X1 U14337 ( .A1(n11017), .A2(n19437), .ZN(n13436) );
  NAND2_X1 U14338 ( .A1(n11208), .A2(n13436), .ZN(n16437) );
  NAND2_X1 U14339 ( .A1(n16437), .A2(n10527), .ZN(n11209) );
  NAND2_X1 U14340 ( .A1(n11210), .A2(n11209), .ZN(n11211) );
  NAND2_X1 U14341 ( .A1(n16178), .A2(n16406), .ZN(n11425) );
  INV_X1 U14342 ( .A(n11212), .ZN(n11213) );
  INV_X1 U14343 ( .A(n15658), .ZN(n16428) );
  NAND2_X1 U14344 ( .A1(n13436), .A2(n13674), .ZN(n13439) );
  NAND2_X1 U14345 ( .A1(n13439), .A2(n19447), .ZN(n11214) );
  NAND2_X1 U14346 ( .A1(n16428), .A2(n11214), .ZN(n11215) );
  AND2_X1 U14347 ( .A1(n11218), .A2(n11217), .ZN(n13406) );
  AND2_X1 U14348 ( .A1(n11225), .A2(n20136), .ZN(n11265) );
  AOI222_X1 U14349 ( .A1(P2_REIP_REG_29__SCAN_IN), .A2(n11409), .B1(n11406), 
        .B2(P2_EAX_REG_29__SCAN_IN), .C1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), 
        .C2(n11416), .ZN(n11419) );
  NAND2_X1 U14350 ( .A1(n11374), .A2(n11221), .ZN(n11224) );
  NAND2_X1 U14351 ( .A1(n13405), .A2(n11265), .ZN(n11238) );
  NAND2_X1 U14352 ( .A1(n11264), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11227) );
  INV_X1 U14353 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n13682) );
  NAND2_X1 U14354 ( .A1(n11225), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11226) );
  NAND2_X1 U14355 ( .A1(n11227), .A2(n9896), .ZN(n13679) );
  AOI22_X1 U14356 ( .A1(n11228), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n11265), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11230) );
  NAND2_X1 U14357 ( .A1(n11264), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11229) );
  NAND2_X1 U14358 ( .A1(n11230), .A2(n11229), .ZN(n11236) );
  INV_X1 U14359 ( .A(n11374), .ZN(n11393) );
  OR2_X1 U14360 ( .A1(n11231), .A2(n11393), .ZN(n11234) );
  MUX2_X1 U14361 ( .A(n11232), .B(n16450), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n11233) );
  NAND2_X1 U14362 ( .A1(n11234), .A2(n11233), .ZN(n13713) );
  NAND2_X1 U14363 ( .A1(n11374), .A2(n11237), .ZN(n11239) );
  OAI211_X1 U14364 ( .C1(n20136), .C2(n20147), .A(n11239), .B(n11238), .ZN(
        n11242) );
  INV_X2 U14365 ( .A(n13420), .ZN(n11406) );
  AOI22_X1 U14366 ( .A1(n11406), .A2(P2_EAX_REG_2__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n11416), .ZN(n11241) );
  NAND2_X1 U14367 ( .A1(n11409), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11240) );
  NAND2_X1 U14368 ( .A1(n11241), .A2(n11240), .ZN(n13726) );
  NOR2_X1 U14369 ( .A1(n13727), .A2(n13726), .ZN(n13728) );
  NOR2_X1 U14370 ( .A1(n11243), .A2(n11242), .ZN(n11244) );
  NAND2_X1 U14371 ( .A1(n11409), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11249) );
  AOI22_X1 U14372 ( .A1(n11416), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11248) );
  NAND2_X1 U14373 ( .A1(n11374), .A2(n11245), .ZN(n11247) );
  NAND2_X1 U14374 ( .A1(n11406), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11246) );
  NAND4_X1 U14375 ( .A1(n11249), .A2(n11248), .A3(n11247), .A4(n11246), .ZN(
        n14083) );
  NAND2_X1 U14376 ( .A1(n14084), .A2(n14083), .ZN(n14085) );
  AOI22_X1 U14377 ( .A1(n11406), .A2(P2_EAX_REG_4__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n11416), .ZN(n11253) );
  NAND2_X1 U14378 ( .A1(n11409), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11252) );
  NAND2_X1 U14379 ( .A1(n11374), .A2(n11250), .ZN(n11251) );
  INV_X1 U14380 ( .A(n11254), .ZN(n11255) );
  AOI22_X1 U14381 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n11409), .B1(n11374), 
        .B2(n11255), .ZN(n11257) );
  AOI22_X1 U14382 ( .A1(n11406), .A2(P2_EAX_REG_5__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n11416), .ZN(n11256) );
  NAND2_X1 U14383 ( .A1(n11257), .A2(n11256), .ZN(n15624) );
  NAND2_X1 U14384 ( .A1(n14104), .A2(n15624), .ZN(n15623) );
  NAND2_X1 U14385 ( .A1(n11374), .A2(n11258), .ZN(n11259) );
  AOI22_X1 U14386 ( .A1(n11406), .A2(P2_EAX_REG_6__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n11416), .ZN(n11261) );
  NAND2_X1 U14387 ( .A1(n11409), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11260) );
  NAND2_X1 U14388 ( .A1(n11261), .A2(n11260), .ZN(n15612) );
  AOI21_X1 U14389 ( .B1(n15613), .B2(n15612), .A(n11262), .ZN(n11263) );
  INV_X2 U14390 ( .A(n11263), .ZN(n16401) );
  INV_X1 U14391 ( .A(n11264), .ZN(n13418) );
  INV_X1 U14392 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n20065) );
  INV_X1 U14393 ( .A(n11265), .ZN(n13419) );
  INV_X1 U14394 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19388) );
  OAI222_X1 U14395 ( .A1(n13418), .A2(n20065), .B1(n13419), .B2(n11076), .C1(
        n13420), .C2(n19388), .ZN(n16400) );
  NOR2_X1 U14396 ( .A1(n13419), .A2(n16395), .ZN(n11281) );
  AOI22_X1 U14397 ( .A1(n10688), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10689), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11269) );
  AOI22_X1 U14398 ( .A1(n13218), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13141), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11268) );
  AOI22_X1 U14399 ( .A1(n10650), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13219), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11267) );
  AOI22_X1 U14400 ( .A1(n13220), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13217), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11266) );
  NAND4_X1 U14401 ( .A1(n11269), .A2(n11268), .A3(n11267), .A4(n11266), .ZN(
        n11279) );
  AOI22_X1 U14402 ( .A1(n10728), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13226), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11277) );
  AOI22_X1 U14403 ( .A1(n13225), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10748), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11276) );
  INV_X1 U14404 ( .A(n13187), .ZN(n13231) );
  INV_X1 U14405 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11272) );
  NAND2_X1 U14406 ( .A1(n13227), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11271) );
  NAND2_X1 U14407 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n13228), .ZN(
        n11270) );
  OAI211_X1 U14408 ( .C1(n13231), .C2(n11272), .A(n11271), .B(n11270), .ZN(
        n11273) );
  INV_X1 U14409 ( .A(n11273), .ZN(n11275) );
  NAND2_X1 U14410 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11274) );
  NAND4_X1 U14411 ( .A1(n11277), .A2(n11276), .A3(n11275), .A4(n11274), .ZN(
        n11278) );
  INV_X1 U14412 ( .A(n13106), .ZN(n19285) );
  OAI22_X1 U14413 ( .A1(n13418), .A2(n14928), .B1(n11393), .B2(n19285), .ZN(
        n11280) );
  AOI211_X1 U14414 ( .C1(n11406), .C2(P2_EAX_REG_8__SCAN_IN), .A(n11281), .B(
        n11280), .ZN(n14924) );
  AOI22_X1 U14415 ( .A1(n11406), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n11416), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11297) );
  NAND2_X1 U14416 ( .A1(n11409), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11296) );
  AOI22_X1 U14417 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10688), .B1(
        n10689), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11285) );
  AOI22_X1 U14418 ( .A1(n10650), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13187), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11284) );
  AOI22_X1 U14419 ( .A1(n13218), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13219), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11283) );
  AOI22_X1 U14420 ( .A1(n13220), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13217), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11282) );
  NAND4_X1 U14421 ( .A1(n11285), .A2(n11284), .A3(n11283), .A4(n11282), .ZN(
        n11294) );
  INV_X1 U14422 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11287) );
  INV_X1 U14423 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11286) );
  OAI22_X1 U14424 ( .A1(n13178), .A2(n11287), .B1(n13177), .B2(n11286), .ZN(
        n11288) );
  AOI21_X1 U14425 ( .B1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n13141), .A(
        n11288), .ZN(n11292) );
  AOI22_X1 U14426 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10728), .B1(
        n10748), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11291) );
  AOI22_X1 U14427 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n13225), .B1(
        n13226), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11290) );
  NAND2_X1 U14428 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11289) );
  NAND4_X1 U14429 ( .A1(n11292), .A2(n11291), .A3(n11290), .A4(n11289), .ZN(
        n11293) );
  NOR2_X1 U14430 ( .A1(n11294), .A2(n11293), .ZN(n13108) );
  INV_X1 U14431 ( .A(n13108), .ZN(n13976) );
  NAND2_X1 U14432 ( .A1(n11374), .A2(n13976), .ZN(n11295) );
  NAND3_X1 U14433 ( .A1(n11297), .A2(n11296), .A3(n11295), .ZN(n15598) );
  INV_X1 U14434 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n11298) );
  INV_X1 U14435 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16329) );
  OAI22_X1 U14436 ( .A1(n13420), .A2(n11298), .B1(n16329), .B2(n13419), .ZN(
        n11314) );
  AOI22_X1 U14437 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10688), .B1(
        n10689), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11302) );
  AOI22_X1 U14438 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n13141), .B1(
        n13220), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11301) );
  AOI22_X1 U14439 ( .A1(n13218), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13217), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11300) );
  AOI22_X1 U14440 ( .A1(n10650), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13219), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11299) );
  NAND4_X1 U14441 ( .A1(n11302), .A2(n11301), .A3(n11300), .A4(n11299), .ZN(
        n11312) );
  AOI22_X1 U14442 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10728), .B1(
        n13226), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11310) );
  AOI22_X1 U14443 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n13225), .B1(
        n10748), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11309) );
  INV_X1 U14444 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11305) );
  NAND2_X1 U14445 ( .A1(n13227), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11304) );
  NAND2_X1 U14446 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n13228), .ZN(
        n11303) );
  OAI211_X1 U14447 ( .C1(n13231), .C2(n11305), .A(n11304), .B(n11303), .ZN(
        n11306) );
  INV_X1 U14448 ( .A(n11306), .ZN(n11308) );
  NAND2_X1 U14449 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n11307) );
  NAND4_X1 U14450 ( .A1(n11310), .A2(n11309), .A3(n11308), .A4(n11307), .ZN(
        n11311) );
  INV_X1 U14451 ( .A(n19276), .ZN(n14002) );
  NOR2_X1 U14452 ( .A1(n11393), .A2(n14002), .ZN(n11313) );
  AOI211_X1 U14453 ( .C1(n11409), .C2(P2_REIP_REG_10__SCAN_IN), .A(n11314), 
        .B(n11313), .ZN(n16376) );
  AOI22_X1 U14454 ( .A1(n11406), .A2(P2_EAX_REG_11__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n11416), .ZN(n11330) );
  NAND2_X1 U14455 ( .A1(n11409), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n11329) );
  AOI22_X1 U14456 ( .A1(n10688), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10689), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11318) );
  AOI22_X1 U14457 ( .A1(n10650), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13187), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11317) );
  AOI22_X1 U14458 ( .A1(n13218), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13219), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11316) );
  AOI22_X1 U14459 ( .A1(n13220), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13217), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11315) );
  NAND4_X1 U14460 ( .A1(n11318), .A2(n11317), .A3(n11316), .A4(n11315), .ZN(
        n11327) );
  INV_X1 U14461 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11320) );
  INV_X1 U14462 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11319) );
  OAI22_X1 U14463 ( .A1(n13178), .A2(n11320), .B1(n13177), .B2(n11319), .ZN(
        n11321) );
  AOI21_X1 U14464 ( .B1(n13141), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A(
        n11321), .ZN(n11325) );
  AOI22_X1 U14465 ( .A1(n10728), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10748), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11324) );
  AOI22_X1 U14466 ( .A1(n13225), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13226), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11323) );
  NAND2_X1 U14467 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n11322) );
  NAND4_X1 U14468 ( .A1(n11325), .A2(n11324), .A3(n11323), .A4(n11322), .ZN(
        n11326) );
  NAND2_X1 U14469 ( .A1(n11374), .A2(n14004), .ZN(n11328) );
  NAND3_X1 U14470 ( .A1(n11330), .A2(n11329), .A3(n11328), .ZN(n15585) );
  NAND2_X1 U14471 ( .A1(n15584), .A2(n15585), .ZN(n15557) );
  AOI22_X1 U14472 ( .A1(n11406), .A2(P2_EAX_REG_12__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n11416), .ZN(n11344) );
  NAND2_X1 U14473 ( .A1(n11409), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11343) );
  AOI22_X1 U14474 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10688), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11334) );
  AOI22_X1 U14475 ( .A1(n13218), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13141), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11333) );
  AOI22_X1 U14476 ( .A1(n13220), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13187), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11332) );
  AOI22_X1 U14477 ( .A1(n13217), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13219), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11331) );
  NAND4_X1 U14478 ( .A1(n11334), .A2(n11333), .A3(n11332), .A4(n11331), .ZN(
        n11341) );
  INV_X1 U14479 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13314) );
  OAI22_X1 U14480 ( .A1(n13178), .A2(n10196), .B1(n13177), .B2(n13314), .ZN(
        n11335) );
  AOI21_X1 U14481 ( .B1(n10650), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n11335), .ZN(n11339) );
  AOI22_X1 U14482 ( .A1(n10728), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10748), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11338) );
  AOI22_X1 U14483 ( .A1(n13225), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13226), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11337) );
  NAND2_X1 U14484 ( .A1(n10689), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11336) );
  NAND4_X1 U14485 ( .A1(n11339), .A2(n11338), .A3(n11337), .A4(n11336), .ZN(
        n11340) );
  NAND2_X1 U14486 ( .A1(n11374), .A2(n19269), .ZN(n11342) );
  NAND3_X1 U14487 ( .A1(n11344), .A2(n11343), .A3(n11342), .ZN(n15559) );
  AOI22_X1 U14488 ( .A1(n10688), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10689), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11349) );
  AOI22_X1 U14489 ( .A1(n10650), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13187), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11348) );
  AOI22_X1 U14490 ( .A1(n13218), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13219), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11347) );
  AOI22_X1 U14491 ( .A1(n13220), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13217), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11346) );
  NAND4_X1 U14492 ( .A1(n11349), .A2(n11348), .A3(n11347), .A4(n11346), .ZN(
        n11358) );
  INV_X1 U14493 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11351) );
  INV_X1 U14494 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11350) );
  OAI22_X1 U14495 ( .A1(n13178), .A2(n11351), .B1(n13177), .B2(n11350), .ZN(
        n11352) );
  AOI21_X1 U14496 ( .B1(n13141), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A(
        n11352), .ZN(n11356) );
  AOI22_X1 U14497 ( .A1(n10728), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10748), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11355) );
  AOI22_X1 U14498 ( .A1(n13225), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13226), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11354) );
  NAND2_X1 U14499 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11353) );
  NAND4_X1 U14500 ( .A1(n11356), .A2(n11355), .A3(n11354), .A4(n11353), .ZN(
        n11357) );
  AOI22_X1 U14501 ( .A1(n11409), .A2(P2_REIP_REG_13__SCAN_IN), .B1(n11374), 
        .B2(n19264), .ZN(n11360) );
  AOI22_X1 U14502 ( .A1(n11406), .A2(P2_EAX_REG_13__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n11416), .ZN(n11359) );
  NAND2_X1 U14503 ( .A1(n11360), .A2(n11359), .ZN(n15541) );
  NAND2_X1 U14504 ( .A1(n15539), .A2(n15541), .ZN(n15540) );
  AOI22_X1 U14505 ( .A1(n11406), .A2(P2_EAX_REG_14__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n11416), .ZN(n11377) );
  NAND2_X1 U14506 ( .A1(n11409), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11376) );
  AOI22_X1 U14507 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n10689), .B1(
        n10688), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11364) );
  AOI22_X1 U14508 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n13141), .B1(
        n13220), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11363) );
  AOI22_X1 U14509 ( .A1(n10650), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13217), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11362) );
  AOI22_X1 U14510 ( .A1(n13218), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13219), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11361) );
  NAND4_X1 U14511 ( .A1(n11364), .A2(n11363), .A3(n11362), .A4(n11361), .ZN(
        n11373) );
  AOI22_X1 U14512 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10728), .B1(
        n13225), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11371) );
  AOI22_X1 U14513 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n10748), .B1(
        n13226), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11370) );
  INV_X1 U14514 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13359) );
  NAND2_X1 U14515 ( .A1(n13227), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11366) );
  NAND2_X1 U14516 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n13228), .ZN(
        n11365) );
  OAI211_X1 U14517 ( .C1(n13231), .C2(n13359), .A(n11366), .B(n11365), .ZN(
        n11367) );
  INV_X1 U14518 ( .A(n11367), .ZN(n11369) );
  NAND2_X1 U14519 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n11368) );
  NAND4_X1 U14520 ( .A1(n11371), .A2(n11370), .A3(n11369), .A4(n11368), .ZN(
        n11372) );
  NAND2_X1 U14521 ( .A1(n11374), .A2(n19263), .ZN(n11375) );
  AOI22_X1 U14522 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10688), .B1(
        n10689), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11381) );
  AOI22_X1 U14523 ( .A1(n10650), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13187), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11380) );
  AOI22_X1 U14524 ( .A1(n13218), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13219), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11379) );
  AOI22_X1 U14525 ( .A1(n13220), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13217), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11378) );
  NAND4_X1 U14526 ( .A1(n11381), .A2(n11380), .A3(n11379), .A4(n11378), .ZN(
        n11390) );
  INV_X1 U14527 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11383) );
  INV_X1 U14528 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11382) );
  OAI22_X1 U14529 ( .A1(n13178), .A2(n11383), .B1(n13177), .B2(n11382), .ZN(
        n11384) );
  AOI21_X1 U14530 ( .B1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n13141), .A(
        n11384), .ZN(n11388) );
  AOI22_X1 U14531 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10728), .B1(
        n10748), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11387) );
  AOI22_X1 U14532 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n13225), .B1(
        n13226), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11386) );
  NAND2_X1 U14533 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11385) );
  NAND4_X1 U14534 ( .A1(n11388), .A2(n11387), .A3(n11386), .A4(n11385), .ZN(
        n11389) );
  NOR2_X1 U14535 ( .A1(n11390), .A2(n11389), .ZN(n14173) );
  AOI22_X1 U14536 ( .A1(n11406), .A2(P2_EAX_REG_15__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n11416), .ZN(n11392) );
  NAND2_X1 U14537 ( .A1(n11409), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11391) );
  OAI211_X1 U14538 ( .C1(n14173), .C2(n11393), .A(n11392), .B(n11391), .ZN(
        n15508) );
  AOI22_X1 U14539 ( .A1(n11406), .A2(P2_EAX_REG_16__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n11416), .ZN(n11395) );
  NAND2_X1 U14540 ( .A1(n11409), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11394) );
  NAND2_X1 U14541 ( .A1(n11395), .A2(n11394), .ZN(n14901) );
  AOI22_X1 U14542 ( .A1(n11406), .A2(P2_EAX_REG_17__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n11416), .ZN(n11397) );
  NAND2_X1 U14543 ( .A1(n11409), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11396) );
  NAND2_X1 U14544 ( .A1(n11397), .A2(n11396), .ZN(n15100) );
  AOI22_X1 U14545 ( .A1(n11406), .A2(P2_EAX_REG_18__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n11416), .ZN(n11399) );
  NAND2_X1 U14546 ( .A1(n11409), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11398) );
  AOI22_X1 U14547 ( .A1(n11406), .A2(P2_EAX_REG_19__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n11416), .ZN(n11401) );
  NAND2_X1 U14548 ( .A1(n11409), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11400) );
  AOI22_X1 U14549 ( .A1(n11406), .A2(P2_EAX_REG_20__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n11416), .ZN(n11403) );
  NAND2_X1 U14550 ( .A1(n11409), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11402) );
  NAND2_X1 U14551 ( .A1(n11403), .A2(n11402), .ZN(n15445) );
  INV_X1 U14552 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n15082) );
  INV_X1 U14553 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15221) );
  OAI222_X1 U14554 ( .A1(n13418), .A2(n20088), .B1(n13420), .B2(n15082), .C1(
        n15221), .C2(n13419), .ZN(n14856) );
  AND2_X2 U14555 ( .A1(n14854), .A2(n14856), .ZN(n15412) );
  AOI22_X1 U14556 ( .A1(n11406), .A2(P2_EAX_REG_22__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n11416), .ZN(n11405) );
  NAND2_X1 U14557 ( .A1(n11409), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11404) );
  NAND2_X1 U14558 ( .A1(n11405), .A2(n11404), .ZN(n15413) );
  INV_X1 U14559 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20092) );
  INV_X1 U14560 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n13575) );
  OAI222_X1 U14561 ( .A1(n13418), .A2(n20092), .B1(n13420), .B2(n13575), .C1(
        n15395), .C2(n13419), .ZN(n15075) );
  AOI22_X1 U14562 ( .A1(n11406), .A2(P2_EAX_REG_24__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n11416), .ZN(n11408) );
  NAND2_X1 U14563 ( .A1(n11409), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11407) );
  AND2_X1 U14564 ( .A1(n11408), .A2(n11407), .ZN(n15064) );
  AOI22_X1 U14565 ( .A1(n11406), .A2(P2_EAX_REG_25__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n11416), .ZN(n11411) );
  NAND2_X1 U14566 ( .A1(n11409), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11410) );
  AOI22_X1 U14567 ( .A1(n11406), .A2(P2_EAX_REG_26__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n11416), .ZN(n11413) );
  NAND2_X1 U14568 ( .A1(n11409), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11412) );
  NAND2_X1 U14569 ( .A1(n11413), .A2(n11412), .ZN(n15048) );
  AOI22_X1 U14570 ( .A1(n11406), .A2(P2_EAX_REG_27__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n11416), .ZN(n11415) );
  NAND2_X1 U14571 ( .A1(n11409), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11414) );
  NAND2_X1 U14572 ( .A1(n11415), .A2(n11414), .ZN(n15038) );
  AND2_X2 U14573 ( .A1(n15037), .A2(n15038), .ZN(n15040) );
  AOI22_X1 U14574 ( .A1(n11406), .A2(P2_EAX_REG_28__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n11416), .ZN(n11418) );
  NAND2_X1 U14575 ( .A1(n11409), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11417) );
  NAND2_X1 U14576 ( .A1(n11418), .A2(n11417), .ZN(n15028) );
  AOI21_X1 U14577 ( .B1(n11419), .B2(n15030), .A(n13421), .ZN(n16177) );
  NOR2_X1 U14578 ( .A1(n19176), .A2(n20104), .ZN(n15120) );
  INV_X1 U14579 ( .A(n11420), .ZN(n14262) );
  AOI21_X1 U14580 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11421) );
  NOR3_X1 U14581 ( .A1(n11422), .A2(n14262), .A3(n11421), .ZN(n11423) );
  AOI211_X1 U14582 ( .C1(n16387), .C2(n16177), .A(n15120), .B(n11423), .ZN(
        n11424) );
  OAI211_X1 U14583 ( .C1(n15339), .C2(n11426), .A(n11425), .B(n11424), .ZN(
        n11427) );
  AOI21_X1 U14584 ( .B1(n16390), .B2(n15129), .A(n11427), .ZN(n11428) );
  INV_X1 U14585 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18951) );
  NOR2_X1 U14586 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18951), .ZN(
        n11675) );
  INV_X1 U14587 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16519) );
  NOR2_X2 U14588 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11436), .ZN(
        n11474) );
  AOI22_X1 U14589 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11443) );
  OR2_X2 U14590 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n15775), .ZN(
        n11448) );
  INV_X1 U14591 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17063) );
  AOI22_X1 U14592 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11431) );
  AOI22_X1 U14593 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11430) );
  OAI211_X1 U14594 ( .C1(n11448), .C2(n17063), .A(n11431), .B(n11430), .ZN(
        n11442) );
  INV_X2 U14595 ( .A(n11479), .ZN(n17211) );
  AOI22_X1 U14596 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11440) );
  AOI22_X1 U14597 ( .A1(n17313), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11439) );
  NOR2_X2 U14598 ( .A1(n18807), .A2(n11434), .ZN(n11497) );
  AOI22_X1 U14599 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17309), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11438) );
  INV_X2 U14600 ( .A(n9887), .ZN(n17310) );
  NAND2_X1 U14601 ( .A1(n17310), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11437) );
  NAND4_X1 U14602 ( .A1(n11440), .A2(n11439), .A3(n11438), .A4(n11437), .ZN(
        n11441) );
  OAI211_X1 U14603 ( .C1(n17312), .C2(n17222), .A(n11443), .B(n9873), .ZN(
        n16495) );
  INV_X1 U14604 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15744) );
  AOI22_X1 U14605 ( .A1(n17313), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17310), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11456) );
  INV_X1 U14606 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17339) );
  AOI22_X1 U14607 ( .A1(n11497), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11446) );
  AOI22_X1 U14608 ( .A1(n17304), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11445) );
  OAI211_X1 U14609 ( .C1(n17312), .C2(n17339), .A(n11446), .B(n11445), .ZN(
        n11454) );
  INV_X2 U14610 ( .A(n11638), .ZN(n17285) );
  AOI22_X1 U14611 ( .A1(n9811), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17309), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11452) );
  AOI22_X1 U14612 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11451) );
  AOI22_X1 U14613 ( .A1(n11474), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11450) );
  NAND2_X1 U14614 ( .A1(n17268), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11449) );
  NAND4_X1 U14615 ( .A1(n11452), .A2(n11451), .A3(n11450), .A4(n11449), .ZN(
        n11453) );
  AOI211_X1 U14616 ( .C1(n11444), .C2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A(
        n11454), .B(n11453), .ZN(n11455) );
  AOI22_X1 U14617 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11466) );
  INV_X1 U14618 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17347) );
  AOI22_X1 U14619 ( .A1(n11497), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17291), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11458) );
  AOI22_X1 U14620 ( .A1(n17313), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17285), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11457) );
  OAI211_X1 U14621 ( .C1(n17312), .C2(n17347), .A(n11458), .B(n11457), .ZN(
        n11464) );
  INV_X1 U14622 ( .A(n9890), .ZN(n17314) );
  AOI22_X1 U14623 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17309), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11462) );
  AOI22_X1 U14624 ( .A1(n9812), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11461) );
  AOI22_X1 U14625 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11519), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11460) );
  NAND2_X1 U14626 ( .A1(n17310), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11459) );
  NAND4_X1 U14627 ( .A1(n11462), .A2(n11461), .A3(n11460), .A4(n11459), .ZN(
        n11463) );
  AOI211_X1 U14628 ( .C1(n17293), .C2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A(
        n11464), .B(n11463), .ZN(n11465) );
  OAI211_X1 U14629 ( .C1(n17237), .C2(n17153), .A(n11466), .B(n11465), .ZN(
        n11725) );
  INV_X1 U14630 ( .A(n11725), .ZN(n17498) );
  AOI22_X1 U14631 ( .A1(n9812), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17310), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11470) );
  INV_X1 U14632 ( .A(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15712) );
  AOI22_X1 U14633 ( .A1(n11522), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11519), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11473) );
  AOI22_X1 U14634 ( .A1(n11471), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11472) );
  OAI211_X1 U14635 ( .C1(n17312), .C2(n17354), .A(n11473), .B(n11472), .ZN(
        n11477) );
  INV_X1 U14636 ( .A(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17179) );
  AOI22_X1 U14637 ( .A1(n11474), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11475) );
  OAI21_X1 U14638 ( .B1(n17237), .B2(n17179), .A(n11475), .ZN(n11476) );
  INV_X1 U14639 ( .A(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17169) );
  AOI22_X1 U14640 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17309), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11480) );
  OAI21_X1 U14641 ( .B1(n11479), .B2(n17169), .A(n11480), .ZN(n11482) );
  INV_X1 U14642 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17359) );
  AOI22_X1 U14643 ( .A1(n17310), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11495) );
  AOI22_X1 U14644 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11486) );
  AOI22_X1 U14645 ( .A1(n17313), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11519), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11485) );
  OAI211_X1 U14646 ( .C1(n11448), .C2(n17290), .A(n11486), .B(n11485), .ZN(
        n11493) );
  AOI22_X1 U14647 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17291), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11491) );
  AOI22_X1 U14648 ( .A1(n17285), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17309), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11490) );
  AOI22_X1 U14649 ( .A1(n11487), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11522), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11489) );
  NAND2_X1 U14650 ( .A1(n11474), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11488) );
  NAND4_X1 U14651 ( .A1(n11491), .A2(n11490), .A3(n11489), .A4(n11488), .ZN(
        n11492) );
  AOI211_X1 U14652 ( .C1(n11444), .C2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A(
        n11493), .B(n11492), .ZN(n11494) );
  INV_X1 U14653 ( .A(n11533), .ZN(n11716) );
  INV_X2 U14654 ( .A(n11523), .ZN(n17200) );
  INV_X1 U14655 ( .A(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17138) );
  AOI22_X1 U14656 ( .A1(n17304), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11496) );
  OAI21_X1 U14657 ( .B1(n9856), .B2(n17138), .A(n11496), .ZN(n11506) );
  INV_X1 U14658 ( .A(n11497), .ZN(n17288) );
  INV_X1 U14659 ( .A(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17232) );
  INV_X2 U14660 ( .A(n11498), .ZN(n17325) );
  AOI22_X1 U14661 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11504) );
  INV_X1 U14662 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15732) );
  INV_X1 U14663 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17343) );
  OAI22_X1 U14664 ( .A1(n17197), .A2(n15732), .B1(n17312), .B2(n17343), .ZN(
        n11503) );
  AOI22_X1 U14665 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11501) );
  AOI22_X1 U14666 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17285), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11500) );
  AOI22_X1 U14667 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11499) );
  NAND3_X1 U14668 ( .A1(n11501), .A2(n11500), .A3(n11499), .ZN(n11502) );
  OAI211_X1 U14669 ( .C1(n17288), .C2(n17232), .A(n11504), .B(n9917), .ZN(
        n11505) );
  INV_X1 U14670 ( .A(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17053) );
  AOI22_X1 U14671 ( .A1(n17285), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11507) );
  OAI21_X1 U14672 ( .B1(n9888), .B2(n17053), .A(n11507), .ZN(n11517) );
  INV_X1 U14673 ( .A(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11515) );
  AOI22_X1 U14674 ( .A1(n17309), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11514) );
  INV_X1 U14675 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17108) );
  AOI22_X1 U14676 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11508) );
  OAI21_X1 U14677 ( .B1(n17237), .B2(n17108), .A(n11508), .ZN(n11512) );
  INV_X1 U14678 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17333) );
  AOI22_X1 U14679 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11510) );
  AOI22_X1 U14680 ( .A1(n17313), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9812), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11509) );
  OAI211_X1 U14681 ( .C1(n17312), .C2(n17333), .A(n11510), .B(n11509), .ZN(
        n11511) );
  AOI211_X1 U14682 ( .C1(n17293), .C2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A(
        n11512), .B(n11511), .ZN(n11513) );
  OAI211_X1 U14683 ( .C1(n17197), .C2(n11515), .A(n11514), .B(n11513), .ZN(
        n11516) );
  NOR2_X4 U14684 ( .A1(n17484), .A2(n11549), .ZN(n17797) );
  INV_X1 U14685 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n18008) );
  INV_X1 U14686 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18029) );
  NOR2_X1 U14687 ( .A1(n18029), .A2(n18015), .ZN(n17995) );
  XNOR2_X1 U14688 ( .A(n11719), .B(n11518), .ZN(n11542) );
  NAND2_X1 U14689 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n11716), .ZN(
        n11532) );
  AOI22_X1 U14690 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17293), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11531) );
  INV_X1 U14691 ( .A(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18396) );
  AOI22_X1 U14692 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__0__SCAN_IN), .B2(n17309), .ZN(n11521) );
  AOI22_X1 U14693 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n11519), .B1(
        n17291), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11520) );
  OAI211_X1 U14694 ( .C1(n11467), .C2(n18396), .A(n11521), .B(n11520), .ZN(
        n11529) );
  AOI22_X1 U14695 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n11487), .B1(
        P3_INSTQUEUE_REG_3__0__SCAN_IN), .B2(n17273), .ZN(n11527) );
  AOI22_X1 U14696 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n11497), .B1(
        P3_INSTQUEUE_REG_13__0__SCAN_IN), .B2(n17211), .ZN(n11526) );
  AOI22_X1 U14697 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17285), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11525) );
  NAND2_X1 U14698 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n17310), .ZN(
        n11524) );
  NAND4_X1 U14699 ( .A1(n11527), .A2(n11526), .A3(n11525), .A4(n11524), .ZN(
        n11528) );
  AOI211_X1 U14700 ( .C1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .C2(n11444), .A(
        n11529), .B(n11528), .ZN(n11530) );
  OAI211_X1 U14701 ( .C1(n17317), .C2(n17312), .A(n11531), .B(n11530), .ZN(
        n17978) );
  INV_X1 U14702 ( .A(n17978), .ZN(n17987) );
  INV_X1 U14703 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18300) );
  NAND2_X1 U14704 ( .A1(n11532), .A2(n17980), .ZN(n17967) );
  INV_X1 U14705 ( .A(n17503), .ZN(n11534) );
  INV_X1 U14706 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18284) );
  OR2_X1 U14707 ( .A1(n18284), .A2(n11535), .ZN(n11536) );
  NAND2_X1 U14708 ( .A1(n17966), .A2(n11536), .ZN(n17955) );
  XNOR2_X1 U14709 ( .A(n11537), .B(n11725), .ZN(n17954) );
  INV_X1 U14710 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n17956) );
  INV_X1 U14711 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11539) );
  NAND2_X1 U14712 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n11540), .ZN(
        n11541) );
  NAND2_X1 U14713 ( .A1(n11542), .A2(n11544), .ZN(n11545) );
  NAND2_X1 U14714 ( .A1(n17929), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17928) );
  XOR2_X1 U14715 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n11718), .Z(
        n17916) );
  XOR2_X1 U14716 ( .A(n11546), .B(n17916), .Z(n17922) );
  XOR2_X1 U14717 ( .A(n17487), .B(n11546), .Z(n11547) );
  INV_X1 U14718 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18251) );
  AOI21_X1 U14719 ( .B1(n17484), .B2(n11549), .A(n17797), .ZN(n11552) );
  INV_X1 U14720 ( .A(n11552), .ZN(n11550) );
  NAND2_X1 U14721 ( .A1(n11552), .A2(n11551), .ZN(n11553) );
  NOR3_X2 U14722 ( .A1(n17869), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17853) );
  INV_X1 U14723 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18193) );
  INV_X1 U14724 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18152) );
  INV_X1 U14725 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11555) );
  INV_X1 U14726 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18205) );
  NOR2_X1 U14727 ( .A1(n18214), .A2(n18205), .ZN(n18189) );
  NAND2_X1 U14728 ( .A1(n18189), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18163) );
  NAND2_X1 U14729 ( .A1(n18176), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18148) );
  NOR2_X2 U14730 ( .A1(n18099), .A2(n13019), .ZN(n17782) );
  NOR2_X1 U14731 ( .A1(n18127), .A2(n18113), .ZN(n18104) );
  INV_X1 U14732 ( .A(n18104), .ZN(n17757) );
  INV_X1 U14733 ( .A(n17782), .ZN(n17708) );
  NOR2_X1 U14734 ( .A1(n17757), .A2(n17708), .ZN(n17725) );
  NOR2_X1 U14735 ( .A1(n17741), .A2(n17725), .ZN(n17726) );
  INV_X1 U14736 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18084) );
  NOR2_X1 U14737 ( .A1(n18096), .A2(n18084), .ZN(n18074) );
  NAND3_X1 U14738 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n18074), .ZN(n17706) );
  NOR2_X1 U14739 ( .A1(n17726), .A2(n18018), .ZN(n17691) );
  NOR2_X1 U14740 ( .A1(n17757), .A2(n18018), .ZN(n18043) );
  INV_X1 U14741 ( .A(n18043), .ZN(n17996) );
  NOR2_X1 U14742 ( .A1(n17996), .A2(n18048), .ZN(n11743) );
  INV_X1 U14743 ( .A(n11743), .ZN(n17681) );
  INV_X1 U14744 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18107) );
  NAND2_X1 U14745 ( .A1(n18107), .A2(n17886), .ZN(n17761) );
  NOR2_X1 U14746 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17761), .ZN(
        n11557) );
  NAND2_X1 U14747 ( .A1(n11557), .A2(n18084), .ZN(n17727) );
  INV_X1 U14748 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17684) );
  NAND3_X1 U14749 ( .A1(n17691), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n11560), .ZN(n11562) );
  INV_X1 U14750 ( .A(n11560), .ZN(n17671) );
  NOR2_X1 U14751 ( .A1(n17797), .A2(n17671), .ZN(n11561) );
  AOI221_X1 U14752 ( .B1(n17797), .B2(n18029), .C1(n11562), .C2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n11561), .ZN(n17651) );
  NAND2_X1 U14753 ( .A1(n17797), .A2(n11562), .ZN(n17670) );
  AND2_X2 U14754 ( .A1(n18008), .A2(n11563), .ZN(n17640) );
  NOR2_X1 U14755 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17797), .ZN(
        n11564) );
  NAND2_X1 U14756 ( .A1(n17640), .A2(n11564), .ZN(n15778) );
  NOR2_X2 U14757 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15778), .ZN(
        n15839) );
  INV_X1 U14758 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15840) );
  NOR2_X1 U14759 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n15840), .ZN(
        n11678) );
  AOI22_X1 U14760 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17886), .B1(
        n17797), .B2(n18951), .ZN(n11566) );
  AOI22_X1 U14761 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11576) );
  AOI22_X1 U14762 ( .A1(n17309), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11568) );
  AOI22_X1 U14763 ( .A1(n11497), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17200), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11567) );
  OAI211_X1 U14764 ( .C1(n11467), .C2(n17272), .A(n11568), .B(n11567), .ZN(
        n11574) );
  AOI22_X1 U14765 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9812), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11572) );
  AOI22_X1 U14766 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11519), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11571) );
  AOI22_X1 U14767 ( .A1(n17310), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17292), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11570) );
  NAND2_X1 U14768 ( .A1(n11444), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11569) );
  NAND4_X1 U14769 ( .A1(n11572), .A2(n11571), .A3(n11570), .A4(n11569), .ZN(
        n11573) );
  INV_X1 U14770 ( .A(n11701), .ZN(n18343) );
  AOI22_X1 U14771 ( .A1(n17309), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17273), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11578) );
  AOI22_X1 U14772 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11519), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11577) );
  OAI211_X1 U14773 ( .C1(n11467), .C2(n18373), .A(n11578), .B(n11577), .ZN(
        n11584) );
  AOI22_X1 U14774 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11497), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11582) );
  AOI22_X1 U14775 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17200), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11581) );
  AOI22_X1 U14776 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17310), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11580) );
  NAND4_X1 U14777 ( .A1(n11582), .A2(n11581), .A3(n11580), .A4(n11579), .ZN(
        n11583) );
  AOI22_X1 U14778 ( .A1(n17285), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17309), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11587) );
  AOI22_X1 U14779 ( .A1(n11497), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11586) );
  OAI211_X1 U14780 ( .C1(n17312), .C2(n17290), .A(n11587), .B(n11586), .ZN(
        n11593) );
  AOI22_X1 U14781 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17200), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11591) );
  AOI22_X1 U14782 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9812), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11590) );
  AOI22_X1 U14783 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11589) );
  NAND2_X1 U14784 ( .A1(n17310), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11588) );
  NAND4_X1 U14785 ( .A1(n11591), .A2(n11590), .A3(n11589), .A4(n11588), .ZN(
        n11592) );
  NAND2_X1 U14786 ( .A1(n18336), .A2(n18993), .ZN(n11596) );
  NAND2_X1 U14787 ( .A1(n18343), .A2(n11596), .ZN(n11662) );
  INV_X1 U14788 ( .A(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17124) );
  AOI22_X1 U14789 ( .A1(n17310), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17273), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11606) );
  INV_X1 U14790 ( .A(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17122) );
  AOI22_X1 U14791 ( .A1(n11497), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9812), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11598) );
  AOI22_X1 U14792 ( .A1(n17313), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11597) );
  OAI211_X1 U14793 ( .C1(n17312), .C2(n17122), .A(n11598), .B(n11597), .ZN(
        n11604) );
  AOI22_X1 U14794 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11602) );
  AOI22_X1 U14795 ( .A1(n17285), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17309), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11601) );
  AOI22_X1 U14796 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11600) );
  NAND2_X1 U14797 ( .A1(n11444), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11599) );
  NAND4_X1 U14798 ( .A1(n11602), .A2(n11601), .A3(n11600), .A4(n11599), .ZN(
        n11603) );
  AOI211_X1 U14799 ( .C1(n17293), .C2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n11604), .B(n11603), .ZN(n11605) );
  INV_X1 U14800 ( .A(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17110) );
  AOI22_X1 U14801 ( .A1(n17310), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11616) );
  AOI22_X1 U14802 ( .A1(n11497), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11487), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11608) );
  AOI22_X1 U14803 ( .A1(n9811), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17309), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11607) );
  OAI211_X1 U14804 ( .C1(n11467), .C2(n18387), .A(n11608), .B(n11607), .ZN(
        n11614) );
  AOI22_X1 U14805 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17273), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11612) );
  AOI22_X1 U14806 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11519), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11611) );
  AOI22_X1 U14807 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17292), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11610) );
  NAND2_X1 U14808 ( .A1(n11444), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11609) );
  NAND4_X1 U14809 ( .A1(n11612), .A2(n11611), .A3(n11610), .A4(n11609), .ZN(
        n11613) );
  INV_X1 U14810 ( .A(n18796), .ZN(n11656) );
  AOI22_X1 U14811 ( .A1(n17310), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17309), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11627) );
  INV_X1 U14812 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11619) );
  AOI22_X1 U14813 ( .A1(n17304), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11618) );
  AOI22_X1 U14814 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11497), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11617) );
  OAI211_X1 U14815 ( .C1(n17312), .C2(n11619), .A(n11618), .B(n11617), .ZN(
        n11625) );
  AOI22_X1 U14816 ( .A1(n17285), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17273), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11623) );
  AOI22_X1 U14817 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11519), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11622) );
  AOI22_X1 U14818 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11621) );
  NAND2_X1 U14819 ( .A1(n11444), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11620) );
  NAND4_X1 U14820 ( .A1(n11623), .A2(n11622), .A3(n11621), .A4(n11620), .ZN(
        n11624) );
  AOI211_X1 U14821 ( .C1(n17293), .C2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n11625), .B(n11624), .ZN(n11626) );
  NOR2_X1 U14822 ( .A1(n18360), .A2(n17370), .ZN(n11650) );
  INV_X1 U14823 ( .A(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17071) );
  AOI22_X1 U14824 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9813), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11629) );
  AOI22_X1 U14825 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11628) );
  OAI211_X1 U14826 ( .C1(n17237), .C2(n17071), .A(n11629), .B(n11628), .ZN(
        n11635) );
  AOI22_X1 U14827 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11487), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11633) );
  AOI22_X1 U14828 ( .A1(n17309), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11632) );
  AOI22_X1 U14829 ( .A1(n17310), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11631) );
  NAND2_X1 U14830 ( .A1(n17292), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11630) );
  NAND4_X1 U14831 ( .A1(n11633), .A2(n11632), .A3(n11631), .A4(n11630), .ZN(
        n11634) );
  INV_X1 U14832 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17254) );
  AOI22_X1 U14833 ( .A1(n9811), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11640) );
  AOI22_X1 U14834 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11519), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11639) );
  OAI211_X1 U14835 ( .C1(n17237), .C2(n17254), .A(n11640), .B(n11639), .ZN(
        n11645) );
  AOI22_X1 U14836 ( .A1(n11497), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17273), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11644) );
  AOI22_X1 U14837 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17309), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11641) );
  OAI21_X1 U14838 ( .B1(n17170), .B2(n17153), .A(n11641), .ZN(n11643) );
  INV_X1 U14839 ( .A(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17253) );
  AOI22_X1 U14840 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11642) );
  NAND2_X1 U14841 ( .A1(n17409), .A2(n11669), .ZN(n11654) );
  AOI211_X1 U14842 ( .C1(n11656), .C2(n11663), .A(n11650), .B(n11654), .ZN(
        n11646) );
  INV_X1 U14843 ( .A(n11646), .ZN(n11647) );
  NAND2_X1 U14844 ( .A1(n18343), .A2(n18993), .ZN(n11648) );
  NOR2_X1 U14845 ( .A1(n18360), .A2(n11648), .ZN(n11713) );
  NAND2_X1 U14846 ( .A1(n11681), .A2(n11713), .ZN(n16494) );
  INV_X1 U14847 ( .A(n16494), .ZN(n18779) );
  NAND2_X1 U14848 ( .A1(n18779), .A2(n16495), .ZN(n13017) );
  INV_X1 U14849 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15781) );
  NOR2_X1 U14850 ( .A1(n18008), .A2(n15781), .ZN(n15788) );
  NAND2_X1 U14851 ( .A1(n15788), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16510) );
  INV_X1 U14852 ( .A(n16510), .ZN(n11750) );
  NOR2_X1 U14853 ( .A1(n18148), .A2(n13019), .ZN(n17810) );
  NAND2_X1 U14854 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17810), .ZN(
        n17809) );
  NAND2_X1 U14855 ( .A1(n11743), .A2(n18135), .ZN(n18030) );
  NAND2_X1 U14856 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17661), .ZN(
        n17660) );
  NAND3_X1 U14857 ( .A1(n11750), .A2(n17997), .A3(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11649) );
  XOR2_X1 U14858 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n11649), .Z(
        n16505) );
  NAND2_X1 U14859 ( .A1(n17484), .A2(n18779), .ZN(n18185) );
  NAND2_X1 U14860 ( .A1(n11650), .A2(n18786), .ZN(n14219) );
  NOR2_X1 U14861 ( .A1(n14219), .A2(n18993), .ZN(n11653) );
  INV_X1 U14862 ( .A(n11660), .ZN(n11652) );
  NAND2_X1 U14863 ( .A1(n17554), .A2(n18993), .ZN(n16647) );
  NAND2_X1 U14864 ( .A1(n16646), .A2(n16647), .ZN(n11651) );
  NAND2_X1 U14865 ( .A1(n18339), .A2(n17516), .ZN(n11655) );
  AOI21_X1 U14866 ( .B1(n17409), .B2(n11656), .A(n11655), .ZN(n11682) );
  INV_X1 U14867 ( .A(n11682), .ZN(n11657) );
  OAI21_X1 U14868 ( .B1(n11659), .B2(n11703), .A(n11657), .ZN(n11668) );
  NAND2_X1 U14869 ( .A1(n11671), .A2(n11703), .ZN(n11710) );
  INV_X1 U14870 ( .A(n11710), .ZN(n11658) );
  NOR2_X1 U14871 ( .A1(n11659), .A2(n11658), .ZN(n11667) );
  AOI22_X1 U14872 ( .A1(n18796), .A2(n18351), .B1(n18347), .B2(n11660), .ZN(
        n11666) );
  NAND2_X1 U14873 ( .A1(n17409), .A2(n11661), .ZN(n11664) );
  AOI22_X1 U14874 ( .A1(n11664), .A2(n11663), .B1(n11662), .B2(n11661), .ZN(
        n11665) );
  OAI211_X1 U14875 ( .C1(n11667), .C2(n17516), .A(n11666), .B(n11665), .ZN(
        n11683) );
  AOI21_X1 U14876 ( .B1(n11669), .B2(n11668), .A(n11683), .ZN(n11673) );
  NAND2_X1 U14877 ( .A1(n11670), .A2(n11673), .ZN(n18785) );
  AOI21_X2 U14878 ( .B1(n18786), .B2(n15767), .A(n18785), .ZN(n18190) );
  NOR2_X1 U14879 ( .A1(n18351), .A2(n11671), .ZN(n18787) );
  NAND3_X1 U14880 ( .A1(n11703), .A2(n11672), .A3(n18787), .ZN(n15770) );
  NAND2_X1 U14881 ( .A1(n11674), .A2(n11673), .ZN(n16648) );
  NOR2_X4 U14882 ( .A1(n18811), .A2(n18791), .ZN(n18202) );
  INV_X1 U14883 ( .A(n18268), .ZN(n18126) );
  INV_X1 U14884 ( .A(n11675), .ZN(n11680) );
  AOI21_X1 U14885 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18264) );
  NAND3_X1 U14886 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11676) );
  NOR2_X1 U14887 ( .A1(n18264), .A2(n11676), .ZN(n18226) );
  NAND4_X1 U14888 ( .A1(n18226), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18121) );
  NOR2_X1 U14889 ( .A1(n18121), .A2(n18099), .ZN(n18053) );
  NAND3_X1 U14890 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11677) );
  INV_X1 U14891 ( .A(n11676), .ZN(n18252) );
  NAND3_X1 U14892 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n18252), .ZN(n18224) );
  OR2_X1 U14893 ( .A1(n11677), .A2(n18224), .ZN(n18149) );
  NOR2_X1 U14894 ( .A1(n18099), .A2(n18149), .ZN(n18050) );
  NOR2_X1 U14895 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18791), .ZN(
        n18302) );
  INV_X1 U14896 ( .A(n18190), .ZN(n18797) );
  NOR2_X1 U14897 ( .A1(n18302), .A2(n18285), .ZN(n18097) );
  AOI22_X1 U14898 ( .A1(n18811), .A2(n18053), .B1(n18050), .B2(n18097), .ZN(
        n13020) );
  NOR2_X1 U14899 ( .A1(n18048), .A2(n17684), .ZN(n18019) );
  NAND2_X1 U14900 ( .A1(n18043), .A2(n18019), .ZN(n11745) );
  NOR2_X1 U14901 ( .A1(n13020), .A2(n11745), .ZN(n18016) );
  NAND2_X1 U14902 ( .A1(n17995), .A2(n18016), .ZN(n15786) );
  NAND2_X1 U14903 ( .A1(n11750), .A2(n11678), .ZN(n11679) );
  OAI22_X1 U14904 ( .A1(n18126), .A2(n11680), .B1(n15786), .B2(n11679), .ZN(
        n11715) );
  INV_X1 U14905 ( .A(n11681), .ZN(n11684) );
  AOI211_X1 U14906 ( .C1(n11685), .C2(n11684), .A(n11683), .B(n11682), .ZN(
        n15769) );
  OAI22_X1 U14907 ( .A1(n18964), .A2(n18801), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11706) );
  AOI22_X1 U14908 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(n18330), .B2(n10256), .ZN(
        n11691) );
  OR2_X1 U14909 ( .A1(n11691), .A2(n11692), .ZN(n11687) );
  OAI22_X1 U14910 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18328), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n11688), .ZN(n11694) );
  NOR2_X1 U14911 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18328), .ZN(
        n11689) );
  NAND2_X1 U14912 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11688), .ZN(
        n11695) );
  AOI22_X1 U14913 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n11694), .B1(
        n11689), .B2(n11695), .ZN(n11705) );
  OAI21_X1 U14914 ( .B1(n11692), .B2(n11691), .A(n11705), .ZN(n11690) );
  AOI21_X1 U14915 ( .B1(n11692), .B2(n11691), .A(n11690), .ZN(n11699) );
  AOI21_X1 U14916 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n18972), .A(
        n11693), .ZN(n11704) );
  XNOR2_X1 U14917 ( .A(n11706), .B(n11693), .ZN(n11698) );
  INV_X1 U14918 ( .A(n11699), .ZN(n11708) );
  INV_X1 U14919 ( .A(n11694), .ZN(n11697) );
  NAND2_X1 U14920 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n11695), .ZN(
        n11696) );
  AOI21_X1 U14921 ( .B1(n11699), .B2(n11704), .A(n18777), .ZN(n16493) );
  NAND2_X2 U14922 ( .A1(n18933), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18922) );
  NOR2_X1 U14923 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18849) );
  INV_X1 U14924 ( .A(n18849), .ZN(n11700) );
  NAND3_X1 U14925 ( .A1(n18862), .A2(n18922), .A3(n11700), .ZN(n18854) );
  INV_X1 U14926 ( .A(n18854), .ZN(n18992) );
  XOR2_X1 U14927 ( .A(n18993), .B(n11701), .Z(n11702) );
  NAND2_X1 U14928 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n18988) );
  OAI21_X1 U14929 ( .B1(n18992), .B2(n11702), .A(n18988), .ZN(n16630) );
  NOR3_X1 U14930 ( .A1(n11703), .A2(n18777), .A3(n16630), .ZN(n11712) );
  NAND3_X1 U14931 ( .A1(n11706), .A2(n11705), .A3(n11704), .ZN(n11707) );
  NAND3_X1 U14932 ( .A1(n11709), .A2(n11708), .A3(n11707), .ZN(n18782) );
  AOI21_X1 U14933 ( .B1(n18351), .B2(n11710), .A(n18782), .ZN(n11711) );
  AOI211_X1 U14934 ( .C1(n16493), .C2(n11713), .A(n11712), .B(n11711), .ZN(
        n11714) );
  NAND2_X1 U14935 ( .A1(n17978), .A2(n11533), .ZN(n11728) );
  NAND2_X1 U14936 ( .A1(n17503), .A2(n11728), .ZN(n11726) );
  NAND2_X1 U14937 ( .A1(n11726), .A2(n11725), .ZN(n11723) );
  NOR2_X1 U14938 ( .A1(n17495), .A2(n11723), .ZN(n11720) );
  NAND2_X1 U14939 ( .A1(n11720), .A2(n11719), .ZN(n17912) );
  INV_X1 U14940 ( .A(n17912), .ZN(n17914) );
  NAND2_X1 U14941 ( .A1(n11718), .A2(n17914), .ZN(n11717) );
  NOR2_X1 U14942 ( .A1(n11717), .A2(n17484), .ZN(n11741) );
  INV_X1 U14943 ( .A(n11741), .ZN(n11737) );
  XOR2_X1 U14944 ( .A(n16495), .B(n11717), .Z(n17906) );
  XNOR2_X1 U14945 ( .A(n17912), .B(n11718), .ZN(n11736) );
  XOR2_X1 U14946 ( .A(n11720), .B(n11719), .Z(n11721) );
  NAND2_X1 U14947 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n11721), .ZN(
        n11735) );
  INV_X1 U14948 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18257) );
  XNOR2_X1 U14949 ( .A(n18257), .B(n11721), .ZN(n17934) );
  XNOR2_X1 U14950 ( .A(n11723), .B(n11722), .ZN(n11724) );
  NAND2_X1 U14951 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n11724), .ZN(
        n11734) );
  XOR2_X1 U14952 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n11724), .Z(
        n17942) );
  XOR2_X1 U14953 ( .A(n11726), .B(n11725), .Z(n11727) );
  NAND2_X1 U14954 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n11727), .ZN(
        n11733) );
  XNOR2_X1 U14955 ( .A(n17956), .B(n11727), .ZN(n17960) );
  XOR2_X1 U14956 ( .A(n17503), .B(n11728), .Z(n11731) );
  OR2_X1 U14957 ( .A1(n18284), .A2(n11731), .ZN(n11732) );
  AOI21_X1 U14958 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n11533), .A(
        n17978), .ZN(n11730) );
  NOR2_X1 U14959 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n11533), .ZN(
        n11729) );
  AOI221_X1 U14960 ( .B1(n17978), .B2(n11533), .C1(n11730), .C2(n18300), .A(
        n11729), .ZN(n17971) );
  XNOR2_X1 U14961 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n11731), .ZN(
        n17970) );
  NAND2_X1 U14962 ( .A1(n17971), .A2(n17970), .ZN(n17969) );
  NAND2_X1 U14963 ( .A1(n11732), .A2(n17969), .ZN(n17959) );
  NAND2_X1 U14964 ( .A1(n17960), .A2(n17959), .ZN(n17958) );
  NAND2_X1 U14965 ( .A1(n11733), .A2(n17958), .ZN(n17941) );
  NAND2_X1 U14966 ( .A1(n17942), .A2(n17941), .ZN(n17940) );
  NAND2_X1 U14967 ( .A1(n11734), .A2(n17940), .ZN(n17933) );
  NAND2_X1 U14968 ( .A1(n17934), .A2(n17933), .ZN(n17932) );
  NAND2_X1 U14969 ( .A1(n11735), .A2(n17932), .ZN(n17913) );
  AOI222_X1 U14970 ( .A1(n11736), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B1(
        n11736), .B2(n17913), .C1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(
        n17913), .ZN(n17907) );
  NAND2_X1 U14971 ( .A1(n17906), .A2(n17907), .ZN(n17905) );
  NAND2_X1 U14972 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17905), .ZN(
        n11740) );
  NOR2_X1 U14973 ( .A1(n11737), .A2(n11740), .ZN(n11742) );
  NOR2_X1 U14974 ( .A1(n17906), .A2(n17907), .ZN(n11739) );
  NOR2_X1 U14975 ( .A1(n11741), .A2(n11740), .ZN(n11738) );
  AOI211_X1 U14976 ( .C1(n11741), .C2(n11740), .A(n11739), .B(n11738), .ZN(
        n17894) );
  NOR2_X1 U14977 ( .A1(n17894), .A2(n10241), .ZN(n17893) );
  NAND2_X1 U14978 ( .A1(n18140), .A2(n11743), .ZN(n18031) );
  NAND2_X1 U14979 ( .A1(n17995), .A2(n17669), .ZN(n17633) );
  NOR2_X1 U14980 ( .A1(n16510), .A2(n17633), .ZN(n16528) );
  NAND2_X1 U14981 ( .A1(n16528), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11744) );
  XOR2_X1 U14982 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n11744), .Z(
        n16502) );
  NAND2_X1 U14983 ( .A1(n9802), .A2(n18231), .ZN(n18304) );
  NOR2_X1 U14984 ( .A1(n18300), .A2(n18149), .ZN(n18147) );
  INV_X1 U14985 ( .A(n18147), .ZN(n18211) );
  NOR2_X1 U14986 ( .A1(n18099), .A2(n18211), .ZN(n18072) );
  INV_X1 U14987 ( .A(n11745), .ZN(n17994) );
  NAND2_X1 U14988 ( .A1(n17994), .A2(n17995), .ZN(n16511) );
  NOR2_X1 U14989 ( .A1(n16511), .A2(n18008), .ZN(n13021) );
  AOI21_X1 U14990 ( .B1(n18072), .B2(n13021), .A(n18190), .ZN(n11749) );
  INV_X1 U14991 ( .A(n16511), .ZN(n11746) );
  AOI21_X1 U14992 ( .B1(n18053), .B2(n11746), .A(n18792), .ZN(n18001) );
  INV_X1 U14993 ( .A(n18791), .ZN(n18799) );
  AOI21_X1 U14994 ( .B1(n11746), .B2(n18050), .A(n18799), .ZN(n11748) );
  NOR4_X1 U14995 ( .A1(n11749), .A2(n18001), .A3(n11748), .A4(n10081), .ZN(
        n13011) );
  NAND2_X1 U14996 ( .A1(n18965), .A2(n18942), .ZN(n18944) );
  OR3_X2 U14997 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), 
        .A3(n18944), .ZN(n18312) );
  AOI221_X1 U14998 ( .B1(n18126), .B2(n13011), .C1(n11750), .C2(n13011), .A(
        n9822), .ZN(n15844) );
  AOI22_X1 U14999 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n15844), .B1(
        n18308), .B2(P3_REIP_REG_31__SCAN_IN), .ZN(n11751) );
  INV_X1 U15000 ( .A(n11752), .ZN(n11753) );
  NAND2_X1 U15001 ( .A1(n11754), .A2(n11753), .ZN(P3_U2831) );
  INV_X2 U15002 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11947) );
  AND2_X2 U15003 ( .A1(n13925), .A2(n13910), .ZN(n11974) );
  AOI22_X1 U15004 ( .A1(n9844), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11974), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11756) );
  NOR2_X1 U15005 ( .A1(n10020), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11759) );
  NAND2_X1 U15006 ( .A1(n11756), .A2(n11755), .ZN(n11763) );
  AOI22_X1 U15007 ( .A1(n12854), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11868), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11761) );
  NAND2_X1 U15008 ( .A1(n11761), .A2(n11760), .ZN(n11762) );
  NOR2_X1 U15009 ( .A1(n11763), .A2(n11762), .ZN(n11776) );
  NAND2_X1 U15010 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11768) );
  NAND3_X2 U15011 ( .A1(n13924), .A2(n13644), .A3(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11855) );
  INV_X2 U15012 ( .A(n11855), .ZN(n12476) );
  NOR2_X1 U15013 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11764) );
  AOI22_X1 U15014 ( .A1(n12476), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11966), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11767) );
  NAND2_X1 U15015 ( .A1(n11967), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11766) );
  NAND2_X1 U15016 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11765) );
  NAND4_X1 U15017 ( .A1(n11768), .A2(n11767), .A3(n11766), .A4(n11765), .ZN(
        n11774) );
  INV_X1 U15018 ( .A(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12822) );
  INV_X4 U15019 ( .A(n12441), .ZN(n12344) );
  NAND2_X1 U15020 ( .A1(n12344), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11772) );
  NAND2_X1 U15021 ( .A1(n9806), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11771) );
  OAI211_X1 U15022 ( .C1(n9851), .C2(n12822), .A(n11772), .B(n11771), .ZN(
        n11773) );
  NOR2_X1 U15023 ( .A1(n11774), .A2(n11773), .ZN(n11775) );
  AOI22_X1 U15024 ( .A1(n12476), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11966), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11780) );
  NAND2_X1 U15025 ( .A1(n11967), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11778) );
  NAND2_X1 U15026 ( .A1(n9837), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11777) );
  NAND2_X1 U15027 ( .A1(n11798), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11784) );
  NAND2_X1 U15028 ( .A1(n11972), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11783) );
  NAND2_X1 U15029 ( .A1(n9844), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11782) );
  NAND2_X1 U15030 ( .A1(n11974), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11781) );
  NAND2_X1 U15031 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11789) );
  NAND2_X1 U15032 ( .A1(n12854), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11788) );
  NAND2_X1 U15033 ( .A1(n12517), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11787) );
  NAND2_X1 U15034 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11786) );
  INV_X1 U15035 ( .A(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11792) );
  NAND2_X1 U15036 ( .A1(n12344), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11791) );
  NAND2_X1 U15037 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11790) );
  OAI211_X1 U15038 ( .C1(n9850), .C2(n11792), .A(n11791), .B(n11790), .ZN(
        n11793) );
  INV_X1 U15039 ( .A(n11793), .ZN(n11794) );
  NAND4_X4 U15040 ( .A1(n11794), .A2(n11796), .A3(n11795), .A4(n11797), .ZN(
        n11926) );
  AOI22_X1 U15041 ( .A1(n11798), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11972), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11802) );
  AOI22_X1 U15042 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12517), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11801) );
  AOI22_X1 U15043 ( .A1(n9852), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11868), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11800) );
  AOI22_X1 U15044 ( .A1(n9844), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11974), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11799) );
  NAND2_X1 U15045 ( .A1(n11967), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11806) );
  NAND2_X1 U15046 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11805) );
  AOI22_X1 U15047 ( .A1(n12476), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11966), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11804) );
  NAND2_X1 U15048 ( .A1(n9836), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11803) );
  NAND4_X1 U15049 ( .A1(n11806), .A2(n11805), .A3(n11804), .A4(n11803), .ZN(
        n11811) );
  NAND2_X1 U15050 ( .A1(n12344), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11809) );
  NAND2_X1 U15051 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11808) );
  INV_X1 U15052 ( .A(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11816) );
  NAND2_X1 U15053 ( .A1(n9806), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11815) );
  NAND2_X1 U15054 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11814) );
  OAI211_X1 U15055 ( .C1(n11835), .C2(n11816), .A(n11815), .B(n11814), .ZN(
        n11817) );
  INV_X1 U15056 ( .A(n11817), .ZN(n11833) );
  AOI22_X1 U15057 ( .A1(n12476), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11966), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11821) );
  NAND2_X1 U15058 ( .A1(n11961), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11820) );
  NAND2_X1 U15059 ( .A1(n11974), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11819) );
  NAND2_X1 U15060 ( .A1(n11967), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11818) );
  NAND2_X1 U15061 ( .A1(n9852), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11825) );
  NAND2_X1 U15062 ( .A1(n9837), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11824) );
  NAND2_X1 U15063 ( .A1(n12517), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11823) );
  NAND2_X1 U15064 ( .A1(n12344), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11822) );
  NAND2_X1 U15065 ( .A1(n11972), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11829) );
  NAND2_X1 U15066 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11828) );
  NAND2_X1 U15067 ( .A1(n11798), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11827) );
  NAND2_X1 U15068 ( .A1(n12860), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11826) );
  AOI22_X1 U15069 ( .A1(n12476), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11966), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11839) );
  INV_X1 U15070 ( .A(n11835), .ZN(n12477) );
  NAND2_X1 U15071 ( .A1(n12477), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11838) );
  NAND2_X1 U15072 ( .A1(n11967), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11837) );
  INV_X1 U15073 ( .A(n9837), .ZN(n12503) );
  NAND2_X1 U15074 ( .A1(n9837), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11836) );
  AOI22_X1 U15075 ( .A1(n11798), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11972), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11843) );
  AOI22_X1 U15076 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12517), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11842) );
  AOI22_X1 U15077 ( .A1(n9852), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11868), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11841) );
  AOI22_X1 U15078 ( .A1(n12860), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11974), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11840) );
  INV_X1 U15079 ( .A(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11846) );
  NAND2_X1 U15080 ( .A1(n12344), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n11845) );
  NAND2_X1 U15081 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n11844) );
  OAI211_X1 U15082 ( .C1(n9851), .C2(n11846), .A(n11845), .B(n11844), .ZN(
        n11847) );
  AOI22_X1 U15083 ( .A1(n12517), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11798), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11853) );
  AOI22_X1 U15084 ( .A1(n11972), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12344), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11852) );
  AOI22_X1 U15085 ( .A1(n9843), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11974), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11851) );
  AOI22_X1 U15086 ( .A1(n12854), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11807), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11864) );
  NAND2_X1 U15087 ( .A1(n9837), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n11859) );
  NAND2_X1 U15088 ( .A1(n11966), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11858) );
  INV_X1 U15089 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11854) );
  OR2_X1 U15090 ( .A1(n12502), .A2(n11854), .ZN(n11857) );
  INV_X2 U15091 ( .A(n11855), .ZN(n12848) );
  NAND2_X1 U15092 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11856) );
  NAND2_X1 U15093 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11862) );
  INV_X1 U15094 ( .A(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11860) );
  NAND2_X4 U15095 ( .A1(n11866), .A2(n11865), .ZN(n20413) );
  NAND2_X1 U15096 ( .A1(n12074), .A2(n13767), .ZN(n11867) );
  AOI22_X1 U15097 ( .A1(n11798), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11972), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11872) );
  AOI22_X1 U15098 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12517), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11871) );
  AOI22_X1 U15099 ( .A1(n9852), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11868), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11870) );
  AOI22_X1 U15100 ( .A1(n9843), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11974), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11869) );
  AOI22_X1 U15101 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11966), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11876) );
  NAND2_X1 U15102 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11875) );
  NAND2_X1 U15103 ( .A1(n11967), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11874) );
  NAND2_X1 U15104 ( .A1(n9837), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11873) );
  NAND4_X1 U15105 ( .A1(n11876), .A2(n11875), .A3(n11874), .A4(n11873), .ZN(
        n11880) );
  NAND2_X1 U15106 ( .A1(n12344), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11878) );
  NAND2_X1 U15107 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11877) );
  OAI211_X1 U15108 ( .C1(n9851), .C2(n12516), .A(n11878), .B(n11877), .ZN(
        n11879) );
  XNOR2_X1 U15109 ( .A(n21007), .B(P1_STATE_REG_1__SCAN_IN), .ZN(n12992) );
  INV_X1 U15110 ( .A(n9829), .ZN(n11940) );
  NAND2_X1 U15111 ( .A1(n11940), .A2(n9823), .ZN(n11884) );
  NAND2_X1 U15112 ( .A1(n13612), .A2(n11888), .ZN(n11921) );
  AND2_X2 U15113 ( .A1(n13767), .A2(n11926), .ZN(n13630) );
  NAND2_X1 U15114 ( .A1(n11926), .A2(n11928), .ZN(n11889) );
  MUX2_X1 U15115 ( .A(n13630), .B(n11889), .S(n13763), .Z(n11890) );
  NAND2_X2 U15116 ( .A1(n11891), .A2(n11890), .ZN(n11935) );
  NAND2_X1 U15117 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11897) );
  AOI22_X1 U15118 ( .A1(n12476), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11966), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11896) );
  NAND2_X1 U15119 ( .A1(n11967), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11895) );
  NAND2_X1 U15120 ( .A1(n9837), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11894) );
  NAND2_X1 U15121 ( .A1(n9843), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11901) );
  NAND2_X1 U15122 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11900) );
  NAND2_X1 U15123 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11899) );
  NAND2_X1 U15124 ( .A1(n11974), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11898) );
  NAND2_X1 U15125 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11905) );
  NAND2_X1 U15126 ( .A1(n11798), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11904) );
  NAND2_X1 U15127 ( .A1(n11972), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11903) );
  NAND2_X1 U15128 ( .A1(n12344), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11902) );
  NAND2_X1 U15129 ( .A1(n9852), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11907) );
  NAND2_X1 U15130 ( .A1(n12517), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11906) );
  OAI211_X1 U15131 ( .C1(n9851), .C2(n11908), .A(n11907), .B(n11906), .ZN(
        n11910) );
  NAND4_X4 U15132 ( .A1(n11914), .A2(n11913), .A3(n11912), .A4(n11911), .ZN(
        n11917) );
  NAND2_X1 U15133 ( .A1(n13923), .A2(n13753), .ZN(n11915) );
  OAI21_X1 U15134 ( .B1(n11935), .B2(n11915), .A(n11918), .ZN(n11920) );
  OR2_X4 U15135 ( .A1(n11918), .A2(n20413), .ZN(n12976) );
  NAND2_X1 U15136 ( .A1(n11939), .A2(n12976), .ZN(n12898) );
  OR2_X1 U15137 ( .A1(n11918), .A2(n13763), .ZN(n13633) );
  OAI211_X1 U15138 ( .C1(n21069), .C2(n9823), .A(n13779), .B(n13633), .ZN(
        n11938) );
  NAND4_X1 U15139 ( .A1(n11930), .A2(n11921), .A3(n11920), .A4(n11919), .ZN(
        n11923) );
  NAND2_X1 U15140 ( .A1(n13630), .A2(n11918), .ZN(n11922) );
  OAI21_X2 U15141 ( .B1(n11923), .B2(n13769), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11952) );
  INV_X1 U15142 ( .A(n15828), .ZN(n15824) );
  NAND2_X1 U15143 ( .A1(n15824), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11948) );
  NAND2_X1 U15144 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11955) );
  OAI21_X1 U15145 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n11955), .ZN(n20719) );
  OR2_X1 U15146 ( .A1(n12784), .A2(n20719), .ZN(n11924) );
  AND2_X1 U15147 ( .A1(n11948), .A2(n11924), .ZN(n11925) );
  OAI21_X2 U15148 ( .B1(n11952), .B2(n11947), .A(n11925), .ZN(n11933) );
  INV_X1 U15149 ( .A(n13923), .ZN(n11927) );
  INV_X1 U15150 ( .A(n11926), .ZN(n13026) );
  NAND3_X1 U15151 ( .A1(n11927), .A2(n14026), .A3(n13026), .ZN(n13638) );
  NAND2_X1 U15152 ( .A1(n11928), .A2(n20443), .ZN(n13760) );
  NAND2_X1 U15153 ( .A1(n11930), .A2(n13775), .ZN(n11931) );
  NAND2_X2 U15154 ( .A1(n11932), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11946) );
  MUX2_X1 U15155 ( .A(n12784), .B(n15828), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n11934) );
  OAI21_X2 U15156 ( .B1(n11952), .B2(n13644), .A(n11934), .ZN(n11989) );
  NAND2_X1 U15157 ( .A1(n11935), .A2(n14026), .ZN(n13635) );
  OR2_X1 U15158 ( .A1(n13923), .A2(n11928), .ZN(n13777) );
  NAND2_X1 U15159 ( .A1(n14825), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20183) );
  INV_X1 U15160 ( .A(n20183), .ZN(n11936) );
  NAND2_X1 U15161 ( .A1(n11918), .A2(n11917), .ZN(n14028) );
  NAND3_X1 U15162 ( .A1(n13777), .A2(n11936), .A3(n14028), .ZN(n11937) );
  NOR2_X1 U15163 ( .A1(n11938), .A2(n11937), .ZN(n11945) );
  INV_X1 U15164 ( .A(n14026), .ZN(n13482) );
  AND2_X1 U15165 ( .A1(n13482), .A2(n12975), .ZN(n13503) );
  NAND2_X1 U15166 ( .A1(n11940), .A2(n20413), .ZN(n11942) );
  AOI22_X1 U15167 ( .A1(n13503), .A2(n11942), .B1(n12695), .B2(n11941), .ZN(
        n11944) );
  NAND3_X1 U15168 ( .A1(n13612), .A2(n11888), .A3(n11917), .ZN(n11943) );
  NAND4_X1 U15169 ( .A1(n13635), .A2(n11945), .A3(n11944), .A4(n11943), .ZN(
        n11987) );
  INV_X1 U15170 ( .A(n11946), .ZN(n11950) );
  NAND2_X1 U15171 ( .A1(n11948), .A2(n11947), .ZN(n11949) );
  NAND2_X1 U15172 ( .A1(n11950), .A2(n11949), .ZN(n11951) );
  INV_X1 U15174 ( .A(n12784), .ZN(n11957) );
  INV_X1 U15175 ( .A(n11955), .ZN(n11954) );
  NAND2_X1 U15176 ( .A1(n11954), .A2(n12753), .ZN(n20752) );
  NAND2_X1 U15177 ( .A1(n11955), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11956) );
  NAND2_X1 U15178 ( .A1(n20752), .A2(n11956), .ZN(n20389) );
  NAND2_X1 U15179 ( .A1(n11957), .A2(n20389), .ZN(n11959) );
  NAND2_X1 U15180 ( .A1(n15824), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11958) );
  INV_X1 U15181 ( .A(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11964) );
  NAND2_X1 U15182 ( .A1(n12344), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n11963) );
  NAND2_X1 U15183 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n11962) );
  OAI211_X1 U15184 ( .C1(n9849), .C2(n11964), .A(n11963), .B(n11962), .ZN(
        n11965) );
  INV_X1 U15185 ( .A(n11965), .ZN(n11971) );
  INV_X1 U15186 ( .A(n11966), .ZN(n11994) );
  INV_X2 U15187 ( .A(n11994), .ZN(n12801) );
  AOI22_X1 U15188 ( .A1(n12476), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12801), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11970) );
  INV_X2 U15189 ( .A(n12503), .ZN(n12858) );
  AOI22_X1 U15190 ( .A1(n12858), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12847), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11969) );
  NAND2_X1 U15191 ( .A1(n12477), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11968) );
  NAND4_X1 U15192 ( .A1(n11971), .A2(n11970), .A3(n11969), .A4(n11968), .ZN(
        n11980) );
  INV_X1 U15193 ( .A(n11972), .ZN(n12127) );
  AOI22_X1 U15194 ( .A1(n12806), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11978) );
  INV_X2 U15195 ( .A(n12826), .ZN(n12859) );
  AOI22_X1 U15196 ( .A1(n9804), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12859), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11977) );
  AOI22_X1 U15197 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12830), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11976) );
  INV_X1 U15198 ( .A(n11974), .ZN(n12823) );
  AOI22_X1 U15199 ( .A1(n9843), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12849), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11975) );
  NAND4_X1 U15200 ( .A1(n11978), .A2(n11977), .A3(n11976), .A4(n11975), .ZN(
        n11979) );
  OAI21_X2 U15201 ( .B1(n13909), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11981), 
        .ZN(n11986) );
  INV_X1 U15202 ( .A(n12091), .ZN(n11984) );
  AOI22_X1 U15203 ( .A1(n12772), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11984), .B2(n11983), .ZN(n11985) );
  XNOR2_X2 U15204 ( .A(n11986), .B(n11985), .ZN(n12085) );
  INV_X1 U15205 ( .A(n11987), .ZN(n11988) );
  INV_X1 U15206 ( .A(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11992) );
  NAND2_X1 U15207 ( .A1(n12344), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11991) );
  NAND2_X1 U15208 ( .A1(n9806), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11990) );
  OAI211_X1 U15209 ( .C1(n9849), .C2(n11992), .A(n11991), .B(n11990), .ZN(
        n11993) );
  INV_X1 U15210 ( .A(n11993), .ZN(n11998) );
  AOI22_X1 U15211 ( .A1(n12476), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12801), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11997) );
  AOI22_X1 U15212 ( .A1(n12858), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12847), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11996) );
  NAND2_X1 U15213 ( .A1(n12477), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11995) );
  NAND4_X1 U15214 ( .A1(n11998), .A2(n11997), .A3(n11996), .A4(n11995), .ZN(
        n12004) );
  AOI22_X1 U15215 ( .A1(n12806), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12002) );
  AOI22_X1 U15216 ( .A1(n9810), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12859), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12001) );
  AOI22_X1 U15217 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12830), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12000) );
  AOI22_X1 U15218 ( .A1(n9843), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12849), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11999) );
  NAND4_X1 U15219 ( .A1(n12002), .A2(n12001), .A3(n12000), .A4(n11999), .ZN(
        n12003) );
  NAND2_X1 U15220 ( .A1(n9823), .A2(n12694), .ZN(n12027) );
  INV_X1 U15221 ( .A(n12694), .ZN(n12005) );
  NAND2_X1 U15222 ( .A1(n9823), .A2(n12005), .ZN(n12020) );
  NAND2_X1 U15223 ( .A1(n12847), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12009) );
  NAND2_X1 U15224 ( .A1(n12849), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12008) );
  NAND2_X1 U15225 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12007) );
  NAND2_X1 U15226 ( .A1(n12801), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12006) );
  AND4_X1 U15227 ( .A1(n12009), .A2(n12008), .A3(n12007), .A4(n12006), .ZN(
        n12013) );
  AOI22_X1 U15228 ( .A1(n12830), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12012) );
  NAND2_X1 U15229 ( .A1(n12477), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12011) );
  NAND2_X1 U15230 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12010) );
  NAND4_X1 U15231 ( .A1(n12013), .A2(n12012), .A3(n12011), .A4(n12010), .ZN(
        n12019) );
  AOI22_X1 U15232 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11807), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12017) );
  AOI22_X1 U15233 ( .A1(n11973), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12858), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12016) );
  AOI22_X1 U15234 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12806), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12015) );
  AOI22_X1 U15235 ( .A1(n12038), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12860), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12014) );
  NAND4_X1 U15236 ( .A1(n12017), .A2(n12016), .A3(n12015), .A4(n12014), .ZN(
        n12018) );
  MUX2_X1 U15237 ( .A(n12027), .B(n12020), .S(n12641), .Z(n12021) );
  INV_X1 U15238 ( .A(n12021), .ZN(n12022) );
  NAND2_X1 U15239 ( .A1(n12022), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12072) );
  INV_X1 U15240 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12023) );
  AOI21_X1 U15241 ( .B1(n11918), .B2(n12641), .A(n21075), .ZN(n12024) );
  AND2_X1 U15242 ( .A1(n12024), .A2(n12027), .ZN(n12025) );
  INV_X1 U15243 ( .A(n12027), .ZN(n12028) );
  NAND2_X1 U15244 ( .A1(n12858), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12033) );
  NAND2_X1 U15245 ( .A1(n12801), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12032) );
  NAND2_X1 U15246 ( .A1(n12849), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12031) );
  NAND2_X1 U15247 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12030) );
  AOI22_X1 U15248 ( .A1(n9810), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12036) );
  NAND2_X1 U15249 ( .A1(n12477), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12035) );
  NAND2_X1 U15250 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12034) );
  NAND4_X1 U15251 ( .A1(n12037), .A2(n12036), .A3(n12035), .A4(n12034), .ZN(
        n12044) );
  AOI22_X1 U15252 ( .A1(n12806), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12830), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12042) );
  AOI22_X1 U15253 ( .A1(n9806), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12859), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12041) );
  AOI22_X1 U15254 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12860), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12040) );
  AOI22_X1 U15255 ( .A1(n12038), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12847), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12039) );
  NAND4_X1 U15256 ( .A1(n12042), .A2(n12041), .A3(n12040), .A4(n12039), .ZN(
        n12043) );
  OAI22_X1 U15257 ( .A1(n12092), .A2(n12694), .B1(n12091), .B2(n12050), .ZN(
        n12045) );
  INV_X1 U15258 ( .A(n12045), .ZN(n12048) );
  INV_X1 U15259 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12046) );
  OR2_X1 U15260 ( .A1(n12050), .A2(n12092), .ZN(n12051) );
  NAND2_X1 U15261 ( .A1(n12065), .A2(n9885), .ZN(n12056) );
  INV_X1 U15262 ( .A(n12053), .ZN(n12054) );
  NAND2_X1 U15263 ( .A1(n12640), .A2(n12352), .ZN(n12063) );
  INV_X1 U15264 ( .A(n13760), .ZN(n12057) );
  NAND2_X1 U15265 ( .A1(n12057), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12116) );
  XNOR2_X1 U15266 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20290) );
  AOI21_X1 U15267 ( .B1(n12843), .B2(n20290), .A(n12878), .ZN(n12060) );
  NOR2_X2 U15268 ( .A1(n20443), .A2(n20991), .ZN(n12190) );
  NAND2_X1 U15269 ( .A1(n12879), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n12059) );
  OAI211_X1 U15270 ( .C1(n12116), .C2(n10020), .A(n12060), .B(n12059), .ZN(
        n12061) );
  INV_X1 U15271 ( .A(n12061), .ZN(n12062) );
  NAND2_X1 U15272 ( .A1(n12063), .A2(n12062), .ZN(n12064) );
  NAND2_X1 U15273 ( .A1(n12878), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12083) );
  NAND2_X1 U15274 ( .A1(n12064), .A2(n12083), .ZN(n13894) );
  INV_X1 U15275 ( .A(n13894), .ZN(n12082) );
  XNOR2_X2 U15276 ( .A(n12067), .B(n12066), .ZN(n13948) );
  NAND2_X1 U15277 ( .A1(n13948), .A2(n12352), .ZN(n12071) );
  AOI22_X1 U15278 ( .A1(n12879), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20991), .ZN(n12069) );
  INV_X1 U15279 ( .A(n12116), .ZN(n12136) );
  NAND2_X1 U15280 ( .A1(n12136), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12068) );
  AND2_X1 U15281 ( .A1(n12069), .A2(n12068), .ZN(n12070) );
  NAND2_X1 U15282 ( .A1(n12071), .A2(n12070), .ZN(n13790) );
  AOI21_X1 U15283 ( .B1(n20479), .B2(n12074), .A(n20991), .ZN(n13691) );
  NAND2_X1 U15284 ( .A1(n12075), .A2(n12352), .ZN(n12079) );
  AOI22_X1 U15285 ( .A1(n12879), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20991), .ZN(n12077) );
  NAND2_X1 U15286 ( .A1(n12136), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12076) );
  AND2_X1 U15287 ( .A1(n12077), .A2(n12076), .ZN(n12078) );
  NAND2_X1 U15288 ( .A1(n12079), .A2(n12078), .ZN(n13690) );
  NAND2_X1 U15289 ( .A1(n13691), .A2(n13690), .ZN(n13689) );
  OR2_X1 U15290 ( .A1(n13690), .A2(n12891), .ZN(n12080) );
  NAND2_X1 U15291 ( .A1(n13689), .A2(n12080), .ZN(n13789) );
  NAND2_X1 U15292 ( .A1(n13790), .A2(n13789), .ZN(n13897) );
  NAND2_X1 U15293 ( .A1(n12082), .A2(n12081), .ZN(n13895) );
  INV_X1 U15294 ( .A(n11953), .ZN(n12086) );
  NAND2_X1 U15295 ( .A1(n12086), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12090) );
  NOR3_X1 U15296 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12753), .A3(
        n20791), .ZN(n20635) );
  NAND2_X1 U15297 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20635), .ZN(
        n20631) );
  NAND2_X1 U15298 ( .A1(n12729), .A2(n20631), .ZN(n12087) );
  NAND3_X1 U15299 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20922) );
  INV_X1 U15300 ( .A(n20922), .ZN(n20934) );
  NAND2_X1 U15301 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20934), .ZN(
        n20918) );
  NAND2_X1 U15302 ( .A1(n12087), .A2(n20918), .ZN(n20661) );
  OAI22_X1 U15303 ( .A1(n12784), .A2(n20661), .B1(n15828), .B2(n12729), .ZN(
        n12088) );
  INV_X1 U15304 ( .A(n12088), .ZN(n12089) );
  XNOR2_X2 U15305 ( .A(n13622), .B(n20537), .ZN(n20659) );
  INV_X1 U15306 ( .A(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12095) );
  NAND2_X1 U15307 ( .A1(n12344), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n12094) );
  NAND2_X1 U15308 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n12093) );
  OAI211_X1 U15309 ( .C1(n9849), .C2(n12095), .A(n12094), .B(n12093), .ZN(
        n12096) );
  INV_X1 U15310 ( .A(n12096), .ZN(n12100) );
  AOI22_X1 U15311 ( .A1(n12476), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12801), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12099) );
  AOI22_X1 U15312 ( .A1(n12858), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12847), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12098) );
  NAND2_X1 U15313 ( .A1(n12477), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12097) );
  NAND4_X1 U15314 ( .A1(n12100), .A2(n12099), .A3(n12098), .A4(n12097), .ZN(
        n12106) );
  AOI22_X1 U15315 ( .A1(n12806), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12104) );
  AOI22_X1 U15316 ( .A1(n9804), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12859), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12103) );
  AOI22_X1 U15317 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12830), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12102) );
  AOI22_X1 U15318 ( .A1(n9844), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12849), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12101) );
  NAND4_X1 U15319 ( .A1(n12104), .A2(n12103), .A3(n12102), .A4(n12101), .ZN(
        n12105) );
  AOI22_X1 U15320 ( .A1(n12772), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12741), .B2(n12654), .ZN(n12107) );
  NAND2_X1 U15321 ( .A1(n12109), .A2(n13952), .ZN(n12110) );
  INV_X1 U15322 ( .A(n12352), .ZN(n12172) );
  NAND2_X1 U15323 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12112) );
  INV_X1 U15324 ( .A(n12112), .ZN(n12113) );
  INV_X1 U15325 ( .A(n12138), .ZN(n12139) );
  OAI21_X1 U15326 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n12113), .A(
        n12139), .ZN(n14056) );
  AOI22_X1 U15327 ( .A1(n12843), .A2(n14056), .B1(n12878), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12115) );
  NAND2_X1 U15328 ( .A1(n12190), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n12114) );
  OAI211_X1 U15329 ( .C1(n12116), .C2(n13928), .A(n12115), .B(n12114), .ZN(
        n12117) );
  INV_X1 U15330 ( .A(n12117), .ZN(n12118) );
  INV_X1 U15331 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12119) );
  INV_X1 U15332 ( .A(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12610) );
  NAND2_X1 U15333 ( .A1(n12344), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n12121) );
  NAND2_X1 U15334 ( .A1(n11807), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n12120) );
  OAI211_X1 U15335 ( .C1(n9849), .C2(n12610), .A(n12121), .B(n12120), .ZN(
        n12122) );
  INV_X1 U15336 ( .A(n12122), .ZN(n12126) );
  AOI22_X1 U15337 ( .A1(n12476), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12801), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12125) );
  AOI22_X1 U15338 ( .A1(n12858), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12847), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12124) );
  NAND2_X1 U15339 ( .A1(n12477), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12123) );
  NAND4_X1 U15340 ( .A1(n12126), .A2(n12125), .A3(n12124), .A4(n12123), .ZN(
        n12133) );
  AOI22_X1 U15341 ( .A1(n12806), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12131) );
  AOI22_X1 U15342 ( .A1(n9804), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12859), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12130) );
  AOI22_X1 U15343 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12830), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12129) );
  AOI22_X1 U15344 ( .A1(n12860), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12849), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12128) );
  NAND4_X1 U15345 ( .A1(n12131), .A2(n12130), .A3(n12129), .A4(n12128), .ZN(
        n12132) );
  NAND2_X1 U15346 ( .A1(n12741), .A2(n12666), .ZN(n12134) );
  XNOR2_X1 U15347 ( .A(n9828), .B(n12146), .ZN(n12659) );
  NAND2_X1 U15348 ( .A1(n12136), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12144) );
  INV_X1 U15349 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20268) );
  AOI21_X1 U15350 ( .B1(n20268), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12137) );
  AOI21_X1 U15351 ( .B1(n12190), .B2(P1_EAX_REG_4__SCAN_IN), .A(n12137), .ZN(
        n12143) );
  INV_X1 U15352 ( .A(n12167), .ZN(n12141) );
  NAND2_X1 U15353 ( .A1(n20268), .A2(n12139), .ZN(n12140) );
  NAND2_X1 U15354 ( .A1(n12141), .A2(n12140), .ZN(n20267) );
  NOR2_X1 U15355 ( .A1(n20267), .A2(n12891), .ZN(n12142) );
  AOI21_X1 U15356 ( .B1(n12144), .B2(n12143), .A(n12142), .ZN(n12145) );
  AOI21_X1 U15357 ( .B1(n12659), .B2(n12352), .A(n12145), .ZN(n13999) );
  INV_X1 U15358 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12148) );
  NAND2_X1 U15359 ( .A1(n9843), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n12152) );
  NAND2_X1 U15360 ( .A1(n12849), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n12151) );
  NAND2_X1 U15361 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n12150) );
  NAND2_X1 U15362 ( .A1(n12801), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n12149) );
  AND4_X1 U15363 ( .A1(n12152), .A2(n12151), .A3(n12150), .A4(n12149), .ZN(
        n12156) );
  AOI22_X1 U15364 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n12830), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12155) );
  NAND2_X1 U15365 ( .A1(n12829), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12154) );
  NAND2_X1 U15366 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n12153) );
  NAND4_X1 U15367 ( .A1(n12156), .A2(n12155), .A3(n12154), .A4(n12153), .ZN(
        n12162) );
  AOI22_X1 U15368 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12806), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12160) );
  AOI22_X1 U15369 ( .A1(n9804), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12862), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12159) );
  AOI22_X1 U15370 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n12858), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12158) );
  AOI22_X1 U15371 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n9821), .B1(
        n12847), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12157) );
  NAND4_X1 U15372 ( .A1(n12160), .A2(n12159), .A3(n12158), .A4(n12157), .ZN(
        n12161) );
  NAND2_X1 U15373 ( .A1(n12741), .A2(n12669), .ZN(n12163) );
  NOR2_X1 U15374 ( .A1(n12167), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12168) );
  NOR2_X1 U15375 ( .A1(n12191), .A2(n12168), .ZN(n20253) );
  INV_X1 U15376 ( .A(n12878), .ZN(n12169) );
  INV_X1 U15377 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16039) );
  OAI22_X1 U15378 ( .A1(n20253), .A2(n12891), .B1(n12169), .B2(n16039), .ZN(
        n12170) );
  AOI21_X1 U15379 ( .B1(n12190), .B2(P1_EAX_REG_5__SCAN_IN), .A(n12170), .ZN(
        n12171) );
  NAND2_X1 U15380 ( .A1(n13997), .A2(n14040), .ZN(n14039) );
  INV_X1 U15381 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12173) );
  INV_X1 U15382 ( .A(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12176) );
  NAND2_X1 U15383 ( .A1(n12344), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n12175) );
  NAND2_X1 U15384 ( .A1(n12862), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n12174) );
  OAI211_X1 U15385 ( .C1(n9849), .C2(n12176), .A(n12175), .B(n12174), .ZN(
        n12177) );
  INV_X1 U15386 ( .A(n12177), .ZN(n12181) );
  AOI22_X1 U15387 ( .A1(n12476), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12801), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12180) );
  AOI22_X1 U15388 ( .A1(n12858), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12847), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12179) );
  NAND2_X1 U15389 ( .A1(n12829), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12178) );
  NAND4_X1 U15390 ( .A1(n12181), .A2(n12180), .A3(n12179), .A4(n12178), .ZN(
        n12187) );
  AOI22_X1 U15391 ( .A1(n12806), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12185) );
  AOI22_X1 U15392 ( .A1(n9804), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12859), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12184) );
  AOI22_X1 U15393 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12830), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12183) );
  AOI22_X1 U15394 ( .A1(n12860), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12849), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12182) );
  NAND4_X1 U15395 ( .A1(n12185), .A2(n12184), .A3(n12183), .A4(n12182), .ZN(
        n12186) );
  NAND2_X1 U15396 ( .A1(n12741), .A2(n12683), .ZN(n12188) );
  NAND2_X1 U15397 ( .A1(n12199), .A2(n12200), .ZN(n12675) );
  INV_X1 U15398 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n12197) );
  INV_X1 U15399 ( .A(n12207), .ZN(n12195) );
  INV_X1 U15400 ( .A(n12191), .ZN(n12193) );
  INV_X1 U15401 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12192) );
  NAND2_X1 U15402 ( .A1(n12193), .A2(n12192), .ZN(n12194) );
  NAND2_X1 U15403 ( .A1(n12195), .A2(n12194), .ZN(n20240) );
  AOI22_X1 U15404 ( .A1(n20240), .A2(n12843), .B1(n12878), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12196) );
  OAI21_X1 U15405 ( .B1(n12263), .B2(n12197), .A(n12196), .ZN(n12198) );
  INV_X1 U15406 ( .A(n12199), .ZN(n12202) );
  NAND2_X1 U15407 ( .A1(n12202), .A2(n12201), .ZN(n12674) );
  INV_X1 U15408 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12204) );
  NAND2_X1 U15409 ( .A1(n12741), .A2(n12694), .ZN(n12203) );
  OAI21_X1 U15410 ( .B1(n12764), .B2(n12204), .A(n12203), .ZN(n12205) );
  NAND2_X1 U15411 ( .A1(n12682), .A2(n12352), .ZN(n12212) );
  INV_X1 U15412 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n12206) );
  OAI21_X1 U15413 ( .B1(n12207), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n12229), .ZN(n20228) );
  AOI22_X1 U15414 ( .A1(n20228), .A2(n12843), .B1(n12878), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12208) );
  NAND2_X1 U15415 ( .A1(n12212), .A2(n12211), .ZN(n14120) );
  NAND2_X1 U15416 ( .A1(n14069), .A2(n14120), .ZN(n14119) );
  AOI22_X1 U15417 ( .A1(n9804), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9821), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12216) );
  AOI22_X1 U15418 ( .A1(n12806), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9844), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12215) );
  AOI22_X1 U15419 ( .A1(n12862), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12214) );
  AOI22_X1 U15420 ( .A1(n12038), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12849), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12213) );
  AND4_X1 U15421 ( .A1(n12216), .A2(n12215), .A3(n12214), .A4(n12213), .ZN(
        n12223) );
  AOI22_X1 U15422 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12830), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12222) );
  AOI22_X1 U15423 ( .A1(n12858), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12847), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12219) );
  INV_X1 U15424 ( .A(n12848), .ZN(n12821) );
  AOI22_X1 U15425 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12801), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12218) );
  NAND2_X1 U15426 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12217) );
  AND3_X1 U15427 ( .A1(n12219), .A2(n12218), .A3(n12217), .ZN(n12221) );
  NAND2_X1 U15428 ( .A1(n12829), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12220) );
  NAND4_X1 U15429 ( .A1(n12223), .A2(n12222), .A3(n12221), .A4(n12220), .ZN(
        n12224) );
  NAND2_X1 U15430 ( .A1(n12352), .A2(n12224), .ZN(n12228) );
  NAND2_X1 U15431 ( .A1(n12190), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n12227) );
  INV_X1 U15432 ( .A(n12229), .ZN(n12225) );
  XNOR2_X1 U15433 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n12225), .ZN(
        n20214) );
  AOI22_X1 U15434 ( .A1(n12843), .A2(n20214), .B1(n12878), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12226) );
  XOR2_X1 U15435 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n12248), .Z(n20206) );
  AOI22_X1 U15436 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12233) );
  AOI22_X1 U15437 ( .A1(n9804), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12859), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12232) );
  AOI22_X1 U15438 ( .A1(n12860), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12830), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12231) );
  AOI22_X1 U15439 ( .A1(n12806), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12849), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12230) );
  NAND4_X1 U15440 ( .A1(n12233), .A2(n12232), .A3(n12231), .A4(n12230), .ZN(
        n12242) );
  INV_X1 U15441 ( .A(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12387) );
  NAND2_X1 U15442 ( .A1(n12344), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12235) );
  NAND2_X1 U15443 ( .A1(n12862), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12234) );
  OAI211_X1 U15444 ( .C1(n9849), .C2(n12387), .A(n12235), .B(n12234), .ZN(
        n12236) );
  INV_X1 U15445 ( .A(n12236), .ZN(n12240) );
  AOI22_X1 U15446 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12801), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12239) );
  AOI22_X1 U15447 ( .A1(n12858), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12847), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12238) );
  NAND2_X1 U15448 ( .A1(n12829), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12237) );
  NAND4_X1 U15449 ( .A1(n12240), .A2(n12239), .A3(n12238), .A4(n12237), .ZN(
        n12241) );
  OAI21_X1 U15450 ( .B1(n12242), .B2(n12241), .A(n12352), .ZN(n12245) );
  NAND2_X1 U15451 ( .A1(n12190), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12244) );
  NAND2_X1 U15452 ( .A1(n12878), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12243) );
  NAND3_X1 U15453 ( .A1(n12245), .A2(n12244), .A3(n12243), .ZN(n12246) );
  AOI21_X1 U15454 ( .B1(n20206), .B2(n12058), .A(n12246), .ZN(n14191) );
  XNOR2_X1 U15455 ( .A(n12267), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15956) );
  NAND2_X1 U15456 ( .A1(n15956), .A2(n12058), .ZN(n12266) );
  INV_X1 U15457 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n14217) );
  AOI22_X1 U15458 ( .A1(n12806), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12830), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12252) );
  AOI22_X1 U15459 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12860), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12251) );
  AOI22_X1 U15460 ( .A1(n12038), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12847), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12250) );
  AOI22_X1 U15461 ( .A1(n9804), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12249) );
  AND4_X1 U15462 ( .A1(n12252), .A2(n12251), .A3(n12250), .A4(n12249), .ZN(
        n12259) );
  AOI22_X1 U15463 ( .A1(n12862), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12859), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12258) );
  AOI22_X1 U15464 ( .A1(n12858), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12849), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12255) );
  NAND2_X1 U15465 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n12254) );
  AOI22_X1 U15466 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12801), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12253) );
  AND3_X1 U15467 ( .A1(n12255), .A2(n12254), .A3(n12253), .ZN(n12257) );
  NAND2_X1 U15468 ( .A1(n12829), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n12256) );
  NAND4_X1 U15469 ( .A1(n12259), .A2(n12258), .A3(n12257), .A4(n12256), .ZN(
        n12260) );
  NAND2_X1 U15470 ( .A1(n12352), .A2(n12260), .ZN(n12262) );
  NAND2_X1 U15471 ( .A1(n12878), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12261) );
  OAI211_X1 U15472 ( .C1(n12263), .C2(n14217), .A(n12262), .B(n12261), .ZN(
        n12264) );
  INV_X1 U15473 ( .A(n12264), .ZN(n12265) );
  NAND2_X1 U15474 ( .A1(n12266), .A2(n12265), .ZN(n14188) );
  NAND2_X1 U15475 ( .A1(n12879), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n12270) );
  OAI21_X1 U15476 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n12268), .A(
        n12303), .ZN(n16026) );
  AOI22_X1 U15477 ( .A1(n12843), .A2(n16026), .B1(n12878), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12269) );
  NAND2_X1 U15478 ( .A1(n12270), .A2(n12269), .ZN(n12284) );
  AOI22_X1 U15479 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12274) );
  AOI22_X1 U15480 ( .A1(n12858), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12806), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12273) );
  AOI22_X1 U15481 ( .A1(n9804), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12272) );
  AOI22_X1 U15482 ( .A1(n12830), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12847), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12271) );
  AND4_X1 U15483 ( .A1(n12274), .A2(n12273), .A3(n12272), .A4(n12271), .ZN(
        n12281) );
  AOI22_X1 U15484 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12862), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12280) );
  AOI22_X1 U15485 ( .A1(n12860), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12849), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12277) );
  NAND2_X1 U15486 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n12276) );
  AOI22_X1 U15487 ( .A1(n12476), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12801), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12275) );
  AND3_X1 U15488 ( .A1(n12277), .A2(n12276), .A3(n12275), .ZN(n12279) );
  NAND2_X1 U15489 ( .A1(n12829), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12278) );
  NAND4_X1 U15490 ( .A1(n12281), .A2(n12280), .A3(n12279), .A4(n12278), .ZN(
        n12282) );
  NAND2_X1 U15491 ( .A1(n12352), .A2(n12282), .ZN(n14453) );
  INV_X1 U15492 ( .A(n14453), .ZN(n12283) );
  NAND2_X1 U15493 ( .A1(n14448), .A2(n12283), .ZN(n14450) );
  INV_X1 U15494 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14528) );
  XNOR2_X1 U15495 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n12303), .ZN(
        n16014) );
  INV_X1 U15496 ( .A(n16014), .ZN(n12286) );
  AOI22_X1 U15497 ( .A1(n12878), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n12843), .B2(n12286), .ZN(n12301) );
  AOI22_X1 U15498 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12806), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12290) );
  AOI22_X1 U15499 ( .A1(n12858), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12289) );
  AOI22_X1 U15500 ( .A1(n12862), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9843), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12288) );
  AOI22_X1 U15501 ( .A1(n9804), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12287) );
  AND4_X1 U15502 ( .A1(n12290), .A2(n12289), .A3(n12288), .A4(n12287), .ZN(
        n12298) );
  AOI22_X1 U15503 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12830), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12297) );
  AOI22_X1 U15504 ( .A1(n12847), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12849), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12294) );
  NAND2_X1 U15505 ( .A1(n12291), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n12293) );
  AOI22_X1 U15506 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12801), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12292) );
  AND3_X1 U15507 ( .A1(n12294), .A2(n12293), .A3(n12292), .ZN(n12296) );
  NAND2_X1 U15508 ( .A1(n12829), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12295) );
  NAND4_X1 U15509 ( .A1(n12298), .A2(n12297), .A3(n12296), .A4(n12295), .ZN(
        n12299) );
  NAND2_X1 U15510 ( .A1(n12352), .A2(n12299), .ZN(n12300) );
  OAI211_X1 U15511 ( .C1(n12263), .C2(n14528), .A(n12301), .B(n12300), .ZN(
        n14523) );
  XNOR2_X1 U15512 ( .A(n12321), .B(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15929) );
  AOI22_X1 U15513 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12307) );
  AOI22_X1 U15514 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n12858), .B1(
        n9844), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12306) );
  AOI22_X1 U15515 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n12862), .B1(
        n12847), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12305) );
  AOI22_X1 U15516 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12304) );
  NAND4_X1 U15517 ( .A1(n12307), .A2(n12306), .A3(n12305), .A4(n12304), .ZN(
        n12316) );
  INV_X1 U15518 ( .A(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12458) );
  NAND2_X1 U15519 ( .A1(n12830), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n12309) );
  NAND2_X1 U15520 ( .A1(n9804), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n12308) );
  OAI211_X1 U15521 ( .C1(n9849), .C2(n12458), .A(n12309), .B(n12308), .ZN(
        n12310) );
  INV_X1 U15522 ( .A(n12310), .ZN(n12314) );
  AOI22_X1 U15523 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12801), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12313) );
  AOI22_X1 U15524 ( .A1(n12806), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12849), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12312) );
  NAND2_X1 U15525 ( .A1(n12829), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12311) );
  NAND4_X1 U15526 ( .A1(n12314), .A2(n12313), .A3(n12312), .A4(n12311), .ZN(
        n12315) );
  OAI21_X1 U15527 ( .B1(n12316), .B2(n12315), .A(n12352), .ZN(n12319) );
  NAND2_X1 U15528 ( .A1(n12879), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n12318) );
  NAND2_X1 U15529 ( .A1(n12878), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12317) );
  NAND3_X1 U15530 ( .A1(n12319), .A2(n12318), .A3(n12317), .ZN(n12320) );
  AOI21_X1 U15531 ( .B1(n15929), .B2(n12058), .A(n12320), .ZN(n14441) );
  XOR2_X1 U15532 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n12338), .Z(
        n16003) );
  INV_X1 U15533 ( .A(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12825) );
  NAND2_X1 U15534 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12323) );
  NAND2_X1 U15535 ( .A1(n12038), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n12322) );
  OAI211_X1 U15536 ( .C1(n9849), .C2(n12825), .A(n12323), .B(n12322), .ZN(
        n12324) );
  INV_X1 U15537 ( .A(n12324), .ZN(n12328) );
  AOI22_X1 U15538 ( .A1(n12476), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12801), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12327) );
  AOI22_X1 U15539 ( .A1(n12847), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12849), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12326) );
  NAND2_X1 U15540 ( .A1(n12829), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n12325) );
  NAND4_X1 U15541 ( .A1(n12328), .A2(n12327), .A3(n12326), .A4(n12325), .ZN(
        n12334) );
  AOI22_X1 U15542 ( .A1(n9804), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12806), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12332) );
  AOI22_X1 U15543 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12830), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12331) );
  AOI22_X1 U15544 ( .A1(n12858), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12860), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12330) );
  AOI22_X1 U15545 ( .A1(n12862), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12329) );
  NAND4_X1 U15546 ( .A1(n12332), .A2(n12331), .A3(n12330), .A4(n12329), .ZN(
        n12333) );
  OR2_X1 U15547 ( .A1(n12334), .A2(n12333), .ZN(n12335) );
  AOI22_X1 U15548 ( .A1(n12352), .A2(n12335), .B1(n12878), .B2(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12337) );
  NAND2_X1 U15549 ( .A1(n12879), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12336) );
  OAI211_X1 U15550 ( .C1(n16003), .C2(n12891), .A(n12337), .B(n12336), .ZN(
        n14513) );
  INV_X1 U15551 ( .A(n14435), .ZN(n12360) );
  INV_X1 U15552 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12339) );
  XNOR2_X1 U15553 ( .A(n12379), .B(n12339), .ZN(n15907) );
  AOI22_X1 U15554 ( .A1(n12862), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12343) );
  AOI22_X1 U15555 ( .A1(n9804), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12806), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12342) );
  AOI22_X1 U15556 ( .A1(n9843), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12830), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12341) );
  AOI22_X1 U15557 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12849), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12340) );
  NAND4_X1 U15558 ( .A1(n12343), .A2(n12342), .A3(n12341), .A4(n12340), .ZN(
        n12354) );
  INV_X1 U15559 ( .A(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12500) );
  NAND2_X1 U15560 ( .A1(n12344), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12346) );
  NAND2_X1 U15561 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n12345) );
  OAI211_X1 U15562 ( .C1(n9849), .C2(n12500), .A(n12346), .B(n12345), .ZN(
        n12347) );
  INV_X1 U15563 ( .A(n12347), .ZN(n12351) );
  AOI22_X1 U15564 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12801), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12350) );
  AOI22_X1 U15565 ( .A1(n12858), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12847), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12349) );
  NAND2_X1 U15566 ( .A1(n12477), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n12348) );
  NAND4_X1 U15567 ( .A1(n12351), .A2(n12350), .A3(n12349), .A4(n12348), .ZN(
        n12353) );
  OAI21_X1 U15568 ( .B1(n12354), .B2(n12353), .A(n12352), .ZN(n12357) );
  NAND2_X1 U15569 ( .A1(n12879), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12356) );
  NAND2_X1 U15570 ( .A1(n12878), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12355) );
  NAND3_X1 U15571 ( .A1(n12357), .A2(n12356), .A3(n12355), .ZN(n12358) );
  AOI21_X1 U15572 ( .B1(n15907), .B2(n12058), .A(n12358), .ZN(n14437) );
  INV_X1 U15573 ( .A(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12363) );
  NAND2_X1 U15574 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12362) );
  NAND2_X1 U15575 ( .A1(n12830), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12361) );
  OAI211_X1 U15576 ( .C1(n9849), .C2(n12363), .A(n12362), .B(n12361), .ZN(
        n12364) );
  INV_X1 U15577 ( .A(n12364), .ZN(n12368) );
  AOI22_X1 U15578 ( .A1(n12476), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12801), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12367) );
  AOI22_X1 U15579 ( .A1(n12858), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12849), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12366) );
  NAND2_X1 U15580 ( .A1(n12477), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12365) );
  NAND4_X1 U15581 ( .A1(n12368), .A2(n12367), .A3(n12366), .A4(n12365), .ZN(
        n12374) );
  AOI22_X1 U15582 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12806), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12372) );
  AOI22_X1 U15583 ( .A1(n9804), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9843), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12371) );
  AOI22_X1 U15584 ( .A1(n12862), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12847), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12370) );
  AOI22_X1 U15585 ( .A1(n12038), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12369) );
  NAND4_X1 U15586 ( .A1(n12372), .A2(n12371), .A3(n12370), .A4(n12369), .ZN(
        n12373) );
  NOR2_X1 U15587 ( .A1(n12374), .A2(n12373), .ZN(n12378) );
  NAND2_X1 U15588 ( .A1(n20991), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12375) );
  NAND2_X1 U15589 ( .A1(n12891), .A2(n12375), .ZN(n12376) );
  AOI21_X1 U15590 ( .B1(n12190), .B2(P1_EAX_REG_16__SCAN_IN), .A(n12376), .ZN(
        n12377) );
  OAI21_X1 U15591 ( .B1(n12875), .B2(n12378), .A(n12377), .ZN(n12382) );
  OAI21_X1 U15592 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12380), .A(
        n12414), .ZN(n15996) );
  OR2_X1 U15593 ( .A1(n12891), .A2(n15996), .ZN(n12381) );
  NAND2_X1 U15594 ( .A1(n12382), .A2(n12381), .ZN(n14503) );
  INV_X1 U15595 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n12399) );
  AOI22_X1 U15596 ( .A1(n9804), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11972), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12386) );
  AOI22_X1 U15597 ( .A1(n12806), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12830), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12385) );
  AOI22_X1 U15598 ( .A1(n12860), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12849), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12384) );
  AOI22_X1 U15599 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12383) );
  NAND4_X1 U15600 ( .A1(n12386), .A2(n12385), .A3(n12384), .A4(n12383), .ZN(
        n12396) );
  INV_X1 U15601 ( .A(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12394) );
  INV_X1 U15602 ( .A(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12388) );
  OAI22_X1 U15603 ( .A1(n12821), .A2(n12388), .B1(n11994), .B2(n12387), .ZN(
        n12391) );
  INV_X1 U15604 ( .A(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12544) );
  INV_X1 U15605 ( .A(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12389) );
  OAI22_X1 U15606 ( .A1(n12503), .A2(n12544), .B1(n12502), .B2(n12389), .ZN(
        n12390) );
  AOI211_X1 U15607 ( .C1(n12829), .C2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A(
        n12391), .B(n12390), .ZN(n12393) );
  AOI22_X1 U15608 ( .A1(n12862), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12859), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12392) );
  OAI211_X1 U15609 ( .C1(n9849), .C2(n12394), .A(n12393), .B(n12392), .ZN(
        n12395) );
  OAI21_X1 U15610 ( .B1(n12396), .B2(n12395), .A(n12840), .ZN(n12398) );
  XOR2_X1 U15611 ( .A(n12414), .B(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .Z(
        n14653) );
  AOI22_X1 U15612 ( .A1(n14653), .A2(n12058), .B1(n12878), .B2(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12397) );
  OAI211_X1 U15613 ( .C1(n12263), .C2(n12399), .A(n12398), .B(n12397), .ZN(
        n14396) );
  AOI22_X1 U15614 ( .A1(n9804), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12806), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12403) );
  AOI22_X1 U15615 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12830), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12402) );
  AOI22_X1 U15616 ( .A1(n12862), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12401) );
  AOI22_X1 U15617 ( .A1(n12858), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12847), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12400) );
  AND4_X1 U15618 ( .A1(n12403), .A2(n12402), .A3(n12401), .A4(n12400), .ZN(
        n12412) );
  INV_X1 U15619 ( .A(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12405) );
  INV_X1 U15620 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12404) );
  OAI22_X1 U15621 ( .A1(n11785), .A2(n12405), .B1(n9845), .B2(n12404), .ZN(
        n12410) );
  INV_X1 U15622 ( .A(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12408) );
  AOI22_X1 U15623 ( .A1(n12038), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12849), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12407) );
  AOI22_X1 U15624 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12801), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12406) );
  OAI211_X1 U15625 ( .C1(n9849), .C2(n12408), .A(n12407), .B(n12406), .ZN(
        n12409) );
  AOI211_X1 U15626 ( .C1(n12829), .C2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n12410), .B(n12409), .ZN(n12411) );
  AOI21_X1 U15627 ( .B1(n12412), .B2(n12411), .A(n12875), .ZN(n12417) );
  INV_X1 U15628 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13660) );
  OAI21_X1 U15629 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n20848), .A(
        n20991), .ZN(n12413) );
  OAI21_X1 U15630 ( .B1(n12263), .B2(n13660), .A(n12413), .ZN(n12416) );
  OAI21_X1 U15631 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n12415), .A(
        n12434), .ZN(n15889) );
  OAI22_X1 U15632 ( .A1(n12417), .A2(n12416), .B1(n12891), .B2(n15889), .ZN(
        n14495) );
  XNOR2_X1 U15633 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n12434), .ZN(
        n15883) );
  INV_X1 U15634 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14642) );
  OAI21_X1 U15635 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n14642), .A(n12891), 
        .ZN(n12432) );
  AOI22_X1 U15636 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12862), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12421) );
  AOI22_X1 U15637 ( .A1(n11972), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9844), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12420) );
  AOI22_X1 U15638 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12830), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12419) );
  AOI22_X1 U15639 ( .A1(n12806), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12849), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12418) );
  AND4_X1 U15640 ( .A1(n12421), .A2(n12420), .A3(n12419), .A4(n12418), .ZN(
        n12430) );
  INV_X1 U15641 ( .A(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12423) );
  INV_X1 U15642 ( .A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12422) );
  OAI22_X1 U15643 ( .A1(n9803), .A2(n12423), .B1(n12441), .B2(n12422), .ZN(
        n12428) );
  INV_X1 U15644 ( .A(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12426) );
  AOI22_X1 U15645 ( .A1(n12858), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12847), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12425) );
  AOI22_X1 U15646 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12801), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12424) );
  OAI211_X1 U15647 ( .C1(n9849), .C2(n12426), .A(n12425), .B(n12424), .ZN(
        n12427) );
  AOI211_X1 U15648 ( .C1(n12829), .C2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n12428), .B(n12427), .ZN(n12429) );
  AOI21_X1 U15649 ( .B1(n12430), .B2(n12429), .A(n12875), .ZN(n12431) );
  AOI211_X1 U15650 ( .C1(n12190), .C2(P1_EAX_REG_19__SCAN_IN), .A(n12432), .B(
        n12431), .ZN(n12433) );
  AOI21_X1 U15651 ( .B1(n12843), .B2(n15883), .A(n12433), .ZN(n14431) );
  NAND2_X1 U15652 ( .A1(n14427), .A2(n14431), .ZN(n14429) );
  OAI21_X1 U15653 ( .B1(n12435), .B2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n12492), .ZN(n15984) );
  AOI22_X1 U15654 ( .A1(n12862), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12859), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12439) );
  AOI22_X1 U15655 ( .A1(n12038), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12830), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12438) );
  AOI22_X1 U15656 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11974), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12437) );
  AOI22_X1 U15657 ( .A1(n12806), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12847), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12436) );
  AND4_X1 U15658 ( .A1(n12439), .A2(n12438), .A3(n12437), .A4(n12436), .ZN(
        n12449) );
  INV_X1 U15659 ( .A(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12442) );
  INV_X1 U15660 ( .A(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12440) );
  OAI22_X1 U15661 ( .A1(n9803), .A2(n12442), .B1(n12441), .B2(n12440), .ZN(
        n12447) );
  INV_X1 U15662 ( .A(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12445) );
  AOI22_X1 U15663 ( .A1(n12858), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12860), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12444) );
  AOI22_X1 U15664 ( .A1(n12476), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12801), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12443) );
  OAI211_X1 U15665 ( .C1(n9849), .C2(n12445), .A(n12444), .B(n12443), .ZN(
        n12446) );
  AOI211_X1 U15666 ( .C1(n12829), .C2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n12447), .B(n12446), .ZN(n12448) );
  AOI21_X1 U15667 ( .B1(n12449), .B2(n12448), .A(n12875), .ZN(n12453) );
  INV_X1 U15668 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n12451) );
  NAND2_X1 U15669 ( .A1(n12879), .A2(P1_EAX_REG_20__SCAN_IN), .ZN(n12450) );
  OAI211_X1 U15670 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n12451), .A(n12450), 
        .B(n12891), .ZN(n12452) );
  OAI22_X1 U15671 ( .A1(n15984), .A2(n12891), .B1(n12453), .B2(n12452), .ZN(
        n14487) );
  AOI22_X1 U15672 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12858), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12457) );
  AOI22_X1 U15673 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n9804), .B1(
        n12859), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12456) );
  AOI22_X1 U15674 ( .A1(n12806), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12860), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12455) );
  AOI22_X1 U15675 ( .A1(n12038), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12454) );
  NAND4_X1 U15676 ( .A1(n12457), .A2(n12456), .A3(n12455), .A4(n12454), .ZN(
        n12468) );
  INV_X1 U15677 ( .A(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12466) );
  INV_X1 U15678 ( .A(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12459) );
  OAI22_X1 U15679 ( .A1(n12821), .A2(n12459), .B1(n11994), .B2(n12458), .ZN(
        n12463) );
  INV_X1 U15680 ( .A(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12461) );
  INV_X1 U15681 ( .A(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12460) );
  OAI22_X1 U15682 ( .A1(n12461), .A2(n12502), .B1(n12823), .B2(n12460), .ZN(
        n12462) );
  AOI211_X1 U15683 ( .C1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .C2(n12829), .A(
        n12463), .B(n12462), .ZN(n12465) );
  AOI22_X1 U15684 ( .A1(n12862), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12830), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12464) );
  OAI211_X1 U15685 ( .C1(n12466), .C2(n9849), .A(n12465), .B(n12464), .ZN(
        n12467) );
  OAI21_X1 U15686 ( .B1(n12468), .B2(n12467), .A(n12840), .ZN(n12471) );
  INV_X1 U15687 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14633) );
  AOI21_X1 U15688 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14633), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12469) );
  AOI21_X1 U15689 ( .B1(n12190), .B2(P1_EAX_REG_21__SCAN_IN), .A(n12469), .ZN(
        n12470) );
  XNOR2_X1 U15690 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n12492), .ZN(
        n14637) );
  AOI22_X1 U15691 ( .A1(n12471), .A2(n12470), .B1(n12843), .B2(n14637), .ZN(
        n14386) );
  INV_X1 U15692 ( .A(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12474) );
  NAND2_X1 U15693 ( .A1(n12862), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12473) );
  NAND2_X1 U15694 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n12472) );
  OAI211_X1 U15695 ( .C1(n9849), .C2(n12474), .A(n12473), .B(n12472), .ZN(
        n12475) );
  INV_X1 U15696 ( .A(n12475), .ZN(n12481) );
  AOI22_X1 U15697 ( .A1(n12476), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12801), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12480) );
  AOI22_X1 U15698 ( .A1(n12858), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12847), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12479) );
  NAND2_X1 U15699 ( .A1(n12477), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n12478) );
  NAND4_X1 U15700 ( .A1(n12481), .A2(n12480), .A3(n12479), .A4(n12478), .ZN(
        n12487) );
  AOI22_X1 U15701 ( .A1(n9804), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12806), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12485) );
  AOI22_X1 U15702 ( .A1(n11972), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12830), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12484) );
  AOI22_X1 U15703 ( .A1(n12860), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11974), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12483) );
  AOI22_X1 U15704 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12482) );
  NAND4_X1 U15705 ( .A1(n12485), .A2(n12484), .A3(n12483), .A4(n12482), .ZN(
        n12486) );
  NOR2_X1 U15706 ( .A1(n12487), .A2(n12486), .ZN(n12491) );
  NAND2_X1 U15707 ( .A1(n20991), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12488) );
  NAND2_X1 U15708 ( .A1(n12891), .A2(n12488), .ZN(n12489) );
  AOI21_X1 U15709 ( .B1(n12190), .B2(P1_EAX_REG_22__SCAN_IN), .A(n12489), .ZN(
        n12490) );
  OAI21_X1 U15710 ( .B1(n12875), .B2(n12491), .A(n12490), .ZN(n12499) );
  INV_X1 U15711 ( .A(n12494), .ZN(n12496) );
  INV_X1 U15712 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12495) );
  NAND2_X1 U15713 ( .A1(n12496), .A2(n12495), .ZN(n12497) );
  NAND2_X1 U15714 ( .A1(n12536), .A2(n12497), .ZN(n14625) );
  OR2_X1 U15715 ( .A1(n14625), .A2(n12891), .ZN(n12498) );
  XNOR2_X1 U15716 ( .A(n12536), .B(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14619) );
  INV_X1 U15717 ( .A(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12508) );
  INV_X1 U15718 ( .A(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12501) );
  OAI22_X1 U15719 ( .A1(n12821), .A2(n12501), .B1(n11994), .B2(n12500), .ZN(
        n12505) );
  INV_X1 U15720 ( .A(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12852) );
  INV_X1 U15721 ( .A(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12857) );
  OAI22_X1 U15722 ( .A1(n12503), .A2(n12852), .B1(n12502), .B2(n12857), .ZN(
        n12504) );
  AOI211_X1 U15723 ( .C1(n12829), .C2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n12505), .B(n12504), .ZN(n12507) );
  AOI22_X1 U15724 ( .A1(n9843), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12849), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12506) );
  OAI211_X1 U15725 ( .C1(n9849), .C2(n12508), .A(n12507), .B(n12506), .ZN(
        n12514) );
  AOI22_X1 U15726 ( .A1(n12806), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12512) );
  AOI22_X1 U15727 ( .A1(n9804), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12859), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12511) );
  AOI22_X1 U15728 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12830), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12510) );
  AOI22_X1 U15729 ( .A1(n12862), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12509) );
  NAND4_X1 U15730 ( .A1(n12512), .A2(n12511), .A3(n12510), .A4(n12509), .ZN(
        n12513) );
  NOR2_X1 U15731 ( .A1(n12514), .A2(n12513), .ZN(n12541) );
  INV_X1 U15732 ( .A(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12524) );
  INV_X1 U15733 ( .A(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12515) );
  OAI22_X1 U15734 ( .A1(n12823), .A2(n12516), .B1(n12821), .B2(n12515), .ZN(
        n12521) );
  INV_X1 U15735 ( .A(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12519) );
  INV_X1 U15736 ( .A(n12517), .ZN(n12826) );
  INV_X1 U15737 ( .A(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12518) );
  OAI22_X1 U15738 ( .A1(n9803), .A2(n12519), .B1(n12826), .B2(n12518), .ZN(
        n12520) );
  AOI211_X1 U15739 ( .C1(n12829), .C2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n12521), .B(n12520), .ZN(n12523) );
  AOI22_X1 U15740 ( .A1(n12862), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12522) );
  OAI211_X1 U15741 ( .C1(n9849), .C2(n12524), .A(n12523), .B(n12522), .ZN(
        n12530) );
  AOI22_X1 U15742 ( .A1(n12858), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12860), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12528) );
  AOI22_X1 U15743 ( .A1(n12806), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12527) );
  AOI22_X1 U15744 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12830), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12526) );
  AOI22_X1 U15745 ( .A1(n11967), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12801), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12525) );
  NAND4_X1 U15746 ( .A1(n12528), .A2(n12527), .A3(n12526), .A4(n12525), .ZN(
        n12529) );
  NOR2_X1 U15747 ( .A1(n12530), .A2(n12529), .ZN(n12540) );
  XOR2_X1 U15748 ( .A(n12541), .B(n12540), .Z(n12534) );
  INV_X1 U15749 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n12532) );
  NOR2_X1 U15750 ( .A1(n20848), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12531) );
  OAI22_X1 U15751 ( .A1(n12263), .A2(n12532), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n12531), .ZN(n12533) );
  AOI21_X1 U15752 ( .B1(n12534), .B2(n12840), .A(n12533), .ZN(n12535) );
  AOI21_X1 U15753 ( .B1(n12843), .B2(n14619), .A(n12535), .ZN(n14360) );
  INV_X1 U15754 ( .A(n12537), .ZN(n12538) );
  INV_X1 U15755 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14352) );
  NAND2_X1 U15756 ( .A1(n12538), .A2(n14352), .ZN(n12539) );
  NAND2_X1 U15757 ( .A1(n12580), .A2(n12539), .ZN(n14604) );
  NOR2_X1 U15758 ( .A1(n12541), .A2(n12540), .ZN(n12561) );
  NAND2_X1 U15759 ( .A1(n12861), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12543) );
  NAND2_X1 U15760 ( .A1(n12862), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12542) );
  OAI211_X1 U15761 ( .C1(n9849), .C2(n12544), .A(n12543), .B(n12542), .ZN(
        n12545) );
  INV_X1 U15762 ( .A(n12545), .ZN(n12549) );
  AOI22_X1 U15763 ( .A1(n12476), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12801), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12548) );
  AOI22_X1 U15764 ( .A1(n12858), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12847), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12547) );
  NAND2_X1 U15765 ( .A1(n12829), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12546) );
  NAND4_X1 U15766 ( .A1(n12549), .A2(n12548), .A3(n12547), .A4(n12546), .ZN(
        n12555) );
  AOI22_X1 U15767 ( .A1(n12806), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12553) );
  AOI22_X1 U15768 ( .A1(n9804), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12859), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12552) );
  AOI22_X1 U15769 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12830), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12551) );
  AOI22_X1 U15770 ( .A1(n12860), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12849), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12550) );
  NAND4_X1 U15771 ( .A1(n12553), .A2(n12552), .A3(n12551), .A4(n12550), .ZN(
        n12554) );
  OR2_X1 U15772 ( .A1(n12555), .A2(n12554), .ZN(n12560) );
  XNOR2_X1 U15773 ( .A(n12561), .B(n12560), .ZN(n12558) );
  AOI21_X1 U15774 ( .B1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n20991), .A(
        n12058), .ZN(n12557) );
  NAND2_X1 U15775 ( .A1(n12879), .A2(P1_EAX_REG_24__SCAN_IN), .ZN(n12556) );
  OAI211_X1 U15776 ( .C1(n12558), .C2(n12875), .A(n12557), .B(n12556), .ZN(
        n12559) );
  OAI21_X1 U15777 ( .B1(n12891), .B2(n14604), .A(n12559), .ZN(n14348) );
  NAND2_X1 U15778 ( .A1(n12561), .A2(n12560), .ZN(n12585) );
  INV_X1 U15779 ( .A(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12568) );
  INV_X1 U15780 ( .A(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12564) );
  AOI22_X1 U15781 ( .A1(n9804), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12806), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12563) );
  AOI22_X1 U15782 ( .A1(n11972), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12848), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12562) );
  OAI211_X1 U15783 ( .C1(n9849), .C2(n12564), .A(n12563), .B(n12562), .ZN(
        n12565) );
  INV_X1 U15784 ( .A(n12565), .ZN(n12567) );
  AOI22_X1 U15785 ( .A1(n12862), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12830), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12566) );
  OAI211_X1 U15786 ( .C1(n11835), .C2(n12568), .A(n12567), .B(n12566), .ZN(
        n12574) );
  AOI22_X1 U15787 ( .A1(n12858), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9844), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12572) );
  AOI22_X1 U15788 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12849), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12571) );
  AOI22_X1 U15789 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12570) );
  AOI22_X1 U15790 ( .A1(n11967), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12801), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12569) );
  NAND4_X1 U15791 ( .A1(n12572), .A2(n12571), .A3(n12570), .A4(n12569), .ZN(
        n12573) );
  NOR2_X1 U15792 ( .A1(n12574), .A2(n12573), .ZN(n12586) );
  XOR2_X1 U15793 ( .A(n12585), .B(n12586), .Z(n12575) );
  NAND2_X1 U15794 ( .A1(n12575), .A2(n12840), .ZN(n12579) );
  INV_X1 U15795 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14593) );
  AOI21_X1 U15796 ( .B1(n14593), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12576) );
  AOI21_X1 U15797 ( .B1(n12190), .B2(P1_EAX_REG_25__SCAN_IN), .A(n12576), .ZN(
        n12578) );
  XNOR2_X1 U15798 ( .A(n12580), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14599) );
  INV_X1 U15799 ( .A(n12580), .ZN(n12581) );
  INV_X1 U15800 ( .A(n12582), .ZN(n12583) );
  INV_X1 U15801 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14330) );
  NAND2_X1 U15802 ( .A1(n12583), .A2(n14330), .ZN(n12584) );
  NAND2_X1 U15803 ( .A1(n12789), .A2(n12584), .ZN(n14588) );
  NOR2_X1 U15804 ( .A1(n12586), .A2(n12585), .ZN(n12606) );
  INV_X1 U15805 ( .A(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12589) );
  NAND2_X1 U15806 ( .A1(n12861), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12588) );
  NAND2_X1 U15807 ( .A1(n12862), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n12587) );
  OAI211_X1 U15808 ( .C1(n9849), .C2(n12589), .A(n12588), .B(n12587), .ZN(
        n12590) );
  INV_X1 U15809 ( .A(n12590), .ZN(n12594) );
  AOI22_X1 U15810 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12801), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12593) );
  AOI22_X1 U15811 ( .A1(n12858), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12847), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12592) );
  NAND2_X1 U15812 ( .A1(n12829), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n12591) );
  NAND4_X1 U15813 ( .A1(n12594), .A2(n12593), .A3(n12592), .A4(n12591), .ZN(
        n12600) );
  AOI22_X1 U15814 ( .A1(n12806), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11972), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12598) );
  AOI22_X1 U15815 ( .A1(n9804), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12859), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12597) );
  AOI22_X1 U15816 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12830), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12596) );
  AOI22_X1 U15817 ( .A1(n9844), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12849), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12595) );
  NAND4_X1 U15818 ( .A1(n12598), .A2(n12597), .A3(n12596), .A4(n12595), .ZN(
        n12599) );
  OR2_X1 U15819 ( .A1(n12600), .A2(n12599), .ZN(n12605) );
  XNOR2_X1 U15820 ( .A(n12606), .B(n12605), .ZN(n12603) );
  AOI21_X1 U15821 ( .B1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n20991), .A(
        n12058), .ZN(n12602) );
  NAND2_X1 U15822 ( .A1(n12879), .A2(P1_EAX_REG_26__SCAN_IN), .ZN(n12601) );
  OAI211_X1 U15823 ( .C1(n12603), .C2(n12875), .A(n12602), .B(n12601), .ZN(
        n12604) );
  OAI21_X1 U15824 ( .B1(n12891), .B2(n14588), .A(n12604), .ZN(n14324) );
  NAND2_X1 U15825 ( .A1(n12606), .A2(n12605), .ZN(n12795) );
  INV_X1 U15826 ( .A(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12616) );
  INV_X1 U15827 ( .A(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12607) );
  OAI22_X1 U15828 ( .A1(n12823), .A2(n12608), .B1(n12821), .B2(n12607), .ZN(
        n12613) );
  INV_X1 U15829 ( .A(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12609) );
  OAI22_X1 U15830 ( .A1(n12611), .A2(n12610), .B1(n12127), .B2(n12609), .ZN(
        n12612) );
  AOI211_X1 U15831 ( .C1(n12829), .C2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n12613), .B(n12612), .ZN(n12615) );
  AOI22_X1 U15832 ( .A1(n12862), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12859), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12614) );
  OAI211_X1 U15833 ( .C1(n9849), .C2(n12616), .A(n12615), .B(n12614), .ZN(
        n12622) );
  AOI22_X1 U15834 ( .A1(n12858), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12860), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12620) );
  AOI22_X1 U15835 ( .A1(n9804), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12830), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12619) );
  AOI22_X1 U15836 ( .A1(n11967), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12801), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12618) );
  AOI22_X1 U15837 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12617) );
  NAND4_X1 U15838 ( .A1(n12620), .A2(n12619), .A3(n12618), .A4(n12617), .ZN(
        n12621) );
  NOR2_X1 U15839 ( .A1(n12622), .A2(n12621), .ZN(n12796) );
  XOR2_X1 U15840 ( .A(n12795), .B(n12796), .Z(n12623) );
  NAND2_X1 U15841 ( .A1(n12623), .A2(n12840), .ZN(n12626) );
  INV_X1 U15842 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12785) );
  AOI21_X1 U15843 ( .B1(n12785), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12624) );
  AOI21_X1 U15844 ( .B1(n12190), .B2(P1_EAX_REG_27__SCAN_IN), .A(n12624), .ZN(
        n12625) );
  XNOR2_X1 U15845 ( .A(n12789), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14316) );
  AOI22_X1 U15846 ( .A1(n12626), .A2(n12625), .B1(n12843), .B2(n14316), .ZN(
        n12629) );
  BUF_X1 U15847 ( .A(n12817), .Z(n12628) );
  OAI21_X1 U15848 ( .B1(n12627), .B2(n12629), .A(n12628), .ZN(n14312) );
  NAND2_X1 U15849 ( .A1(n21075), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n21068) );
  NAND2_X1 U15850 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n20933), .ZN(n13960) );
  NOR2_X1 U15851 ( .A1(n14312), .A2(n14689), .ZN(n12788) );
  INV_X1 U15852 ( .A(n13610), .ZN(n12690) );
  NAND2_X1 U15853 ( .A1(n11918), .A2(n20413), .ZN(n12645) );
  OAI21_X1 U15854 ( .B1(n21069), .B2(n12641), .A(n12645), .ZN(n12630) );
  INV_X1 U15855 ( .A(n12630), .ZN(n12631) );
  OAI21_X1 U15856 ( .B1(n20479), .B2(n12690), .A(n12631), .ZN(n13692) );
  NAND2_X1 U15857 ( .A1(n9885), .A2(n11917), .ZN(n12635) );
  XNOR2_X1 U15858 ( .A(n12642), .B(n12641), .ZN(n12632) );
  OAI211_X1 U15859 ( .C1(n21069), .C2(n12632), .A(n10115), .B(n11926), .ZN(
        n12633) );
  INV_X1 U15860 ( .A(n12633), .ZN(n12634) );
  NAND2_X1 U15861 ( .A1(n12635), .A2(n12634), .ZN(n12636) );
  INV_X1 U15862 ( .A(n12636), .ZN(n12637) );
  OR2_X1 U15863 ( .A1(n13694), .A2(n12637), .ZN(n12638) );
  INV_X1 U15864 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12639) );
  XNOR2_X1 U15865 ( .A(n12650), .B(n12639), .ZN(n13792) );
  NAND2_X1 U15866 ( .A1(n12640), .A2(n13610), .ZN(n12649) );
  NAND2_X1 U15867 ( .A1(n12642), .A2(n12641), .ZN(n12643) );
  NAND2_X1 U15868 ( .A1(n12643), .A2(n12644), .ZN(n12653) );
  OAI21_X1 U15869 ( .B1(n12644), .B2(n12643), .A(n12653), .ZN(n12647) );
  INV_X1 U15870 ( .A(n12645), .ZN(n12646) );
  AOI21_X1 U15871 ( .B1(n12695), .B2(n12647), .A(n12646), .ZN(n12648) );
  NAND2_X1 U15872 ( .A1(n12649), .A2(n12648), .ZN(n13791) );
  NAND2_X1 U15873 ( .A1(n13792), .A2(n13791), .ZN(n12652) );
  NAND2_X1 U15874 ( .A1(n12650), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12651) );
  NAND2_X1 U15875 ( .A1(n12652), .A2(n12651), .ZN(n13884) );
  NAND2_X1 U15876 ( .A1(n12653), .A2(n12654), .ZN(n12668) );
  OAI211_X1 U15877 ( .C1(n12654), .C2(n12653), .A(n12695), .B(n12668), .ZN(
        n12655) );
  INV_X1 U15878 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13985) );
  XNOR2_X1 U15879 ( .A(n12656), .B(n13985), .ZN(n13885) );
  NAND2_X1 U15880 ( .A1(n13884), .A2(n13885), .ZN(n12658) );
  NAND2_X1 U15881 ( .A1(n12656), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12657) );
  NAND2_X1 U15882 ( .A1(n12659), .A2(n13610), .ZN(n12662) );
  XNOR2_X1 U15883 ( .A(n12668), .B(n12666), .ZN(n12660) );
  NAND2_X1 U15884 ( .A1(n12660), .A2(n12695), .ZN(n12661) );
  NAND2_X1 U15885 ( .A1(n12662), .A2(n12661), .ZN(n12663) );
  INV_X1 U15886 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13986) );
  XNOR2_X1 U15887 ( .A(n12663), .B(n13986), .ZN(n13983) );
  NAND2_X1 U15888 ( .A1(n12663), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12664) );
  INV_X1 U15889 ( .A(n12666), .ZN(n12667) );
  NOR2_X1 U15890 ( .A1(n12668), .A2(n12667), .ZN(n12670) );
  NAND2_X1 U15891 ( .A1(n12670), .A2(n12669), .ZN(n12685) );
  OAI211_X1 U15892 ( .C1(n12670), .C2(n12669), .A(n12685), .B(n12695), .ZN(
        n12671) );
  INV_X1 U15893 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12913) );
  XNOR2_X1 U15894 ( .A(n12672), .B(n12913), .ZN(n14015) );
  NAND2_X1 U15895 ( .A1(n12672), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12673) );
  NAND3_X1 U15896 ( .A1(n12674), .A2(n12675), .A3(n13610), .ZN(n12678) );
  XNOR2_X1 U15897 ( .A(n12685), .B(n12683), .ZN(n12676) );
  NAND2_X1 U15898 ( .A1(n12676), .A2(n12695), .ZN(n12677) );
  NAND2_X1 U15899 ( .A1(n12678), .A2(n12677), .ZN(n12679) );
  INV_X1 U15900 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14202) );
  XNOR2_X1 U15901 ( .A(n12679), .B(n14202), .ZN(n14047) );
  NAND2_X1 U15902 ( .A1(n14048), .A2(n14047), .ZN(n12681) );
  NAND2_X1 U15903 ( .A1(n12679), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12680) );
  NAND2_X1 U15904 ( .A1(n12682), .A2(n13610), .ZN(n12688) );
  INV_X1 U15905 ( .A(n12683), .ZN(n12684) );
  OR2_X1 U15906 ( .A1(n12685), .A2(n12684), .ZN(n12693) );
  XNOR2_X1 U15907 ( .A(n12693), .B(n12694), .ZN(n12686) );
  NAND2_X1 U15908 ( .A1(n12686), .A2(n12695), .ZN(n12687) );
  NAND2_X1 U15909 ( .A1(n12688), .A2(n12687), .ZN(n12689) );
  NAND2_X1 U15910 ( .A1(n12689), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14134) );
  NOR2_X1 U15911 ( .A1(n12691), .A2(n12690), .ZN(n12692) );
  INV_X1 U15912 ( .A(n12693), .ZN(n12696) );
  NAND3_X1 U15913 ( .A1(n12696), .A2(n12695), .A3(n12694), .ZN(n12697) );
  NAND2_X1 U15914 ( .A1(n14639), .A2(n12697), .ZN(n14178) );
  OR2_X1 U15915 ( .A1(n14178), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12698) );
  NAND2_X1 U15916 ( .A1(n14178), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12699) );
  INV_X1 U15917 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16126) );
  NAND2_X1 U15918 ( .A1(n14680), .A2(n16126), .ZN(n12701) );
  NAND2_X1 U15919 ( .A1(n16018), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15999) );
  INV_X1 U15920 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14812) );
  NAND2_X1 U15921 ( .A1(n14639), .A2(n14812), .ZN(n12702) );
  NAND2_X1 U15922 ( .A1(n15999), .A2(n12702), .ZN(n14675) );
  INV_X1 U15923 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12703) );
  NAND2_X1 U15924 ( .A1(n14639), .A2(n12703), .ZN(n16010) );
  NAND2_X1 U15925 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12704) );
  NAND2_X1 U15926 ( .A1(n14639), .A2(n12704), .ZN(n14674) );
  NAND2_X1 U15927 ( .A1(n16010), .A2(n14674), .ZN(n12705) );
  NOR2_X1 U15928 ( .A1(n14675), .A2(n12705), .ZN(n15997) );
  INV_X1 U15929 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16087) );
  NAND2_X1 U15930 ( .A1(n14639), .A2(n16087), .ZN(n12706) );
  NAND2_X1 U15931 ( .A1(n15997), .A2(n12706), .ZN(n14663) );
  NAND2_X1 U15932 ( .A1(n16018), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15988) );
  OAI21_X1 U15933 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A(n16018), .ZN(n14664) );
  XNOR2_X1 U15934 ( .A(n14639), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15990) );
  INV_X1 U15935 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16084) );
  NAND2_X1 U15936 ( .A1(n14639), .A2(n16084), .ZN(n15986) );
  NAND2_X1 U15937 ( .A1(n15990), .A2(n15986), .ZN(n12707) );
  AOI21_X1 U15938 ( .B1(n14663), .B2(n12712), .A(n12707), .ZN(n14655) );
  OAI21_X1 U15939 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n16018), .A(
        n14655), .ZN(n12708) );
  INV_X1 U15940 ( .A(n12708), .ZN(n12709) );
  INV_X1 U15941 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12710) );
  NAND2_X1 U15942 ( .A1(n12710), .A2(n16132), .ZN(n12711) );
  NAND2_X1 U15943 ( .A1(n16018), .A2(n12711), .ZN(n16007) );
  NAND2_X1 U15944 ( .A1(n16018), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16011) );
  NAND2_X1 U15945 ( .A1(n16007), .A2(n16011), .ZN(n15998) );
  INV_X1 U15946 ( .A(n12712), .ZN(n12713) );
  NOR2_X1 U15947 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12714) );
  NOR2_X1 U15948 ( .A1(n14680), .A2(n12714), .ZN(n12715) );
  NOR2_X1 U15949 ( .A1(n14656), .A2(n12715), .ZN(n12716) );
  XNOR2_X1 U15950 ( .A(n14680), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14647) );
  AND2_X1 U15951 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14767) );
  NAND3_X1 U15952 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14714) );
  INV_X1 U15953 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15857) );
  INV_X1 U15954 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14691) );
  INV_X1 U15955 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12717) );
  NAND2_X1 U15956 ( .A1(n16061), .A2(n12717), .ZN(n12718) );
  NOR2_X1 U15957 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12720) );
  INV_X1 U15958 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16040) );
  AND2_X1 U15959 ( .A1(n12720), .A2(n16040), .ZN(n14585) );
  MUX2_X1 U15960 ( .A(n14539), .B(n9915), .S(n16018), .Z(n12722) );
  AND2_X1 U15961 ( .A1(n11888), .A2(n11918), .ZN(n12724) );
  NOR2_X1 U15962 ( .A1(n12723), .A2(n12724), .ZN(n13613) );
  NAND2_X1 U15963 ( .A1(n13613), .A2(n13630), .ZN(n15816) );
  MUX2_X1 U15964 ( .A(n20791), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n12738) );
  NAND2_X1 U15965 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20843), .ZN(
        n12742) );
  NAND2_X1 U15966 ( .A1(n12738), .A2(n12737), .ZN(n12736) );
  NAND2_X1 U15967 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n20791), .ZN(
        n12725) );
  NAND2_X1 U15968 ( .A1(n12736), .A2(n12725), .ZN(n12755) );
  NAND2_X1 U15969 ( .A1(n12755), .A2(n12726), .ZN(n12728) );
  NAND2_X1 U15970 ( .A1(n12753), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12727) );
  MUX2_X1 U15971 ( .A(n12729), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12734) );
  NOR2_X1 U15972 ( .A1(n13928), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12730) );
  NAND2_X1 U15973 ( .A1(n20371), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12731) );
  NAND2_X1 U15974 ( .A1(n12768), .A2(n12731), .ZN(n12733) );
  INV_X1 U15975 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13626) );
  NAND2_X1 U15976 ( .A1(n13626), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n12732) );
  NAND2_X1 U15977 ( .A1(n12887), .A2(n12741), .ZN(n12778) );
  XNOR2_X1 U15978 ( .A(n12735), .B(n12734), .ZN(n12884) );
  OAI21_X1 U15979 ( .B1(n12738), .B2(n12737), .A(n12736), .ZN(n12883) );
  NAND2_X1 U15980 ( .A1(n12741), .A2(n11917), .ZN(n12740) );
  NAND2_X1 U15981 ( .A1(n13026), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12739) );
  NAND2_X1 U15982 ( .A1(n12740), .A2(n12739), .ZN(n12750) );
  NOR2_X1 U15983 ( .A1(n12883), .A2(n12750), .ZN(n12749) );
  INV_X1 U15984 ( .A(n12741), .ZN(n12761) );
  OAI21_X1 U15985 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20843), .A(
        n12742), .ZN(n12744) );
  NOR2_X1 U15986 ( .A1(n12761), .A2(n12744), .ZN(n12748) );
  INV_X1 U15987 ( .A(n13630), .ZN(n12746) );
  OR2_X1 U15988 ( .A1(n11926), .A2(n11918), .ZN(n12743) );
  NAND2_X1 U15989 ( .A1(n12743), .A2(n13753), .ZN(n12760) );
  INV_X1 U15990 ( .A(n12744), .ZN(n12745) );
  OAI211_X1 U15991 ( .C1(n11918), .C2(n12746), .A(n12760), .B(n12745), .ZN(
        n12747) );
  OAI21_X1 U15992 ( .B1(n12766), .B2(n12748), .A(n12747), .ZN(n12751) );
  NAND2_X1 U15993 ( .A1(n12749), .A2(n12751), .ZN(n12759) );
  INV_X1 U15994 ( .A(n12750), .ZN(n12752) );
  OAI211_X1 U15995 ( .C1(n12752), .C2(n12751), .A(n12883), .B(n12769), .ZN(
        n12758) );
  MUX2_X1 U15996 ( .A(n12753), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n12754) );
  XNOR2_X1 U15997 ( .A(n12755), .B(n12754), .ZN(n12885) );
  NAND2_X1 U15998 ( .A1(n12772), .A2(n12885), .ZN(n12756) );
  OAI211_X1 U15999 ( .C1(n12761), .C2(n12885), .A(n12756), .B(n12760), .ZN(
        n12757) );
  NAND3_X1 U16000 ( .A1(n12759), .A2(n12758), .A3(n12757), .ZN(n12763) );
  AOI22_X1 U16001 ( .A1(n12764), .A2(n12884), .B1(n12763), .B2(n12762), .ZN(
        n12765) );
  AOI21_X1 U16002 ( .B1(n12766), .B2(n12884), .A(n12765), .ZN(n12775) );
  NOR2_X1 U16003 ( .A1(n20371), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12767) );
  NAND2_X1 U16004 ( .A1(n12768), .A2(n12767), .ZN(n12888) );
  NOR2_X1 U16005 ( .A1(n12772), .A2(n12888), .ZN(n12774) );
  INV_X1 U16006 ( .A(n12888), .ZN(n12771) );
  NAND3_X1 U16007 ( .A1(n12772), .A2(n12771), .A3(n12770), .ZN(n12773) );
  OAI21_X1 U16008 ( .B1(n12775), .B2(n12774), .A(n12773), .ZN(n12776) );
  AOI21_X1 U16009 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n21075), .A(
        n12776), .ZN(n12777) );
  NAND2_X1 U16010 ( .A1(n12778), .A2(n12777), .ZN(n12779) );
  NAND2_X1 U16011 ( .A1(n12784), .A2(n20926), .ZN(n21065) );
  NAND2_X1 U16012 ( .A1(n21065), .A2(n21075), .ZN(n12781) );
  NAND2_X1 U16013 ( .A1(n21075), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12783) );
  NAND2_X1 U16014 ( .A1(n20848), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12782) );
  NAND2_X1 U16015 ( .A1(n12783), .A2(n12782), .ZN(n13695) );
  OR2_X2 U16016 ( .A1(n12784), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20369) );
  INV_X1 U16017 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21412) );
  OAI22_X1 U16018 ( .A1(n16038), .A2(n12785), .B1(n20369), .B2(n21412), .ZN(
        n12786) );
  INV_X1 U16019 ( .A(n12789), .ZN(n12790) );
  INV_X1 U16020 ( .A(n12791), .ZN(n12793) );
  INV_X1 U16021 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12792) );
  NAND2_X1 U16022 ( .A1(n12793), .A2(n12792), .ZN(n12794) );
  NAND2_X1 U16023 ( .A1(n12846), .A2(n12794), .ZN(n14580) );
  NOR2_X1 U16024 ( .A1(n12796), .A2(n12795), .ZN(n12819) );
  INV_X1 U16025 ( .A(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12799) );
  NAND2_X1 U16026 ( .A1(n12861), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12798) );
  NAND2_X1 U16027 ( .A1(n12862), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n12797) );
  OAI211_X1 U16028 ( .C1(n9849), .C2(n12799), .A(n12798), .B(n12797), .ZN(
        n12800) );
  INV_X1 U16029 ( .A(n12800), .ZN(n12805) );
  AOI22_X1 U16030 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12801), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12804) );
  AOI22_X1 U16031 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n12858), .B1(
        n12847), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12803) );
  NAND2_X1 U16032 ( .A1(n12829), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n12802) );
  NAND4_X1 U16033 ( .A1(n12805), .A2(n12804), .A3(n12803), .A4(n12802), .ZN(
        n12812) );
  AOI22_X1 U16034 ( .A1(n12806), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11972), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12810) );
  AOI22_X1 U16035 ( .A1(n9804), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12859), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12809) );
  AOI22_X1 U16036 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n9821), .B1(
        n12830), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12808) );
  AOI22_X1 U16037 ( .A1(n9844), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11974), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12807) );
  NAND4_X1 U16038 ( .A1(n12810), .A2(n12809), .A3(n12808), .A4(n12807), .ZN(
        n12811) );
  OR2_X1 U16039 ( .A1(n12812), .A2(n12811), .ZN(n12818) );
  XNOR2_X1 U16040 ( .A(n12819), .B(n12818), .ZN(n12815) );
  AOI21_X1 U16041 ( .B1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20991), .A(
        n12058), .ZN(n12814) );
  NAND2_X1 U16042 ( .A1(n12879), .A2(P1_EAX_REG_28__SCAN_IN), .ZN(n12813) );
  OAI211_X1 U16043 ( .C1(n12815), .C2(n12875), .A(n12814), .B(n12813), .ZN(
        n12816) );
  OAI21_X1 U16044 ( .B1(n12891), .B2(n14580), .A(n12816), .ZN(n14300) );
  NAND2_X1 U16045 ( .A1(n12819), .A2(n12818), .ZN(n12869) );
  INV_X1 U16046 ( .A(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12833) );
  INV_X1 U16047 ( .A(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12820) );
  OAI22_X1 U16048 ( .A1(n12823), .A2(n12822), .B1(n12821), .B2(n12820), .ZN(
        n12828) );
  INV_X1 U16049 ( .A(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12824) );
  OAI22_X1 U16050 ( .A1(n12826), .A2(n12825), .B1(n12127), .B2(n12824), .ZN(
        n12827) );
  AOI211_X1 U16051 ( .C1(n12829), .C2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n12828), .B(n12827), .ZN(n12832) );
  AOI22_X1 U16052 ( .A1(n12830), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12831) );
  OAI211_X1 U16053 ( .C1(n9849), .C2(n12833), .A(n12832), .B(n12831), .ZN(
        n12839) );
  AOI22_X1 U16054 ( .A1(n9804), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12806), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12837) );
  AOI22_X1 U16055 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12862), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12836) );
  AOI22_X1 U16056 ( .A1(n12858), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12860), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12835) );
  AOI22_X1 U16057 ( .A1(n11967), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12801), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12834) );
  NAND4_X1 U16058 ( .A1(n12837), .A2(n12836), .A3(n12835), .A4(n12834), .ZN(
        n12838) );
  NOR2_X1 U16059 ( .A1(n12839), .A2(n12838), .ZN(n12870) );
  XOR2_X1 U16060 ( .A(n12869), .B(n12870), .Z(n12841) );
  NAND2_X1 U16061 ( .A1(n12841), .A2(n12840), .ZN(n12845) );
  INV_X1 U16062 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14565) );
  NOR2_X1 U16063 ( .A1(n14565), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12842) );
  AOI211_X1 U16064 ( .C1(n12190), .C2(P1_EAX_REG_29__SCAN_IN), .A(n12058), .B(
        n12842), .ZN(n12844) );
  XNOR2_X1 U16065 ( .A(n12846), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14567) );
  INV_X1 U16066 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12894) );
  XNOR2_X1 U16067 ( .A(n12895), .B(n12894), .ZN(n14561) );
  AOI22_X1 U16068 ( .A1(n9804), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12847), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12851) );
  AOI22_X1 U16069 ( .A1(n12849), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12848), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12850) );
  OAI211_X1 U16070 ( .C1(n9849), .C2(n12852), .A(n12851), .B(n12850), .ZN(
        n12853) );
  INV_X1 U16071 ( .A(n12853), .ZN(n12856) );
  AOI22_X1 U16072 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12830), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12855) );
  OAI211_X1 U16073 ( .C1(n11835), .C2(n12857), .A(n12856), .B(n12855), .ZN(
        n12868) );
  AOI22_X1 U16074 ( .A1(n12858), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12038), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12866) );
  AOI22_X1 U16075 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12806), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12865) );
  AOI22_X1 U16076 ( .A1(n9844), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12801), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12864) );
  AOI22_X1 U16077 ( .A1(n12862), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12861), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12863) );
  NAND4_X1 U16078 ( .A1(n12866), .A2(n12865), .A3(n12864), .A4(n12863), .ZN(
        n12867) );
  NOR2_X1 U16079 ( .A1(n12868), .A2(n12867), .ZN(n12872) );
  NOR2_X1 U16080 ( .A1(n12870), .A2(n12869), .ZN(n12871) );
  XOR2_X1 U16081 ( .A(n12872), .B(n12871), .Z(n12876) );
  AOI21_X1 U16082 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20991), .A(
        n12058), .ZN(n12874) );
  NAND2_X1 U16083 ( .A1(n12879), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n12873) );
  OAI211_X1 U16084 ( .C1(n12876), .C2(n12875), .A(n12874), .B(n12873), .ZN(
        n12877) );
  OAI21_X1 U16085 ( .B1(n12891), .B2(n14561), .A(n12877), .ZN(n13024) );
  AOI22_X1 U16086 ( .A1(n12879), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n12878), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12880) );
  INV_X1 U16087 ( .A(n13051), .ZN(n14554) );
  NOR3_X1 U16088 ( .A1(n12885), .A2(n12884), .A3(n12883), .ZN(n12886) );
  OR2_X1 U16089 ( .A1(n12887), .A2(n12886), .ZN(n12889) );
  NOR2_X1 U16090 ( .A1(n13480), .A2(n20180), .ZN(n12890) );
  NAND2_X1 U16091 ( .A1(n12882), .A2(n12890), .ZN(n13463) );
  NAND2_X1 U16092 ( .A1(n20991), .A2(n16145), .ZN(n15834) );
  NOR2_X1 U16093 ( .A1(n20799), .A2(n15834), .ZN(n15832) );
  OAI21_X1 U16094 ( .B1(n12891), .B2(n21068), .A(n20369), .ZN(n12892) );
  AOI22_X1 U16095 ( .A1(P1_EBX_REG_31__SCAN_IN), .A2(n13686), .B1(n13771), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12989) );
  MUX2_X1 U16096 ( .A(n12974), .B(n12983), .S(P1_EBX_REG_1__SCAN_IN), .Z(
        n12899) );
  INV_X1 U16097 ( .A(n12899), .ZN(n12901) );
  INV_X1 U16098 ( .A(n13686), .ZN(n12921) );
  NAND2_X1 U16099 ( .A1(n12921), .A2(n14826), .ZN(n12900) );
  NAND2_X1 U16100 ( .A1(n12901), .A2(n12900), .ZN(n12904) );
  INV_X1 U16101 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n12903) );
  OAI21_X1 U16102 ( .B1(n12976), .B2(n12903), .A(n12902), .ZN(n13687) );
  XNOR2_X1 U16103 ( .A(n12904), .B(n13687), .ZN(n13772) );
  AOI21_X1 U16104 ( .B1(n13772), .B2(n13485), .A(n12904), .ZN(n13798) );
  NOR2_X1 U16105 ( .A1(n13686), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12905) );
  NOR2_X1 U16106 ( .A1(n12906), .A2(n12905), .ZN(n13797) );
  NAND2_X1 U16107 ( .A1(n13798), .A2(n13797), .ZN(n13796) );
  INV_X1 U16108 ( .A(n13796), .ZN(n12910) );
  INV_X1 U16109 ( .A(n12976), .ZN(n12953) );
  MUX2_X1 U16110 ( .A(n12983), .B(n12953), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n12908) );
  AND2_X1 U16111 ( .A1(n13771), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12907) );
  NOR2_X1 U16112 ( .A1(n12908), .A2(n12907), .ZN(n13887) );
  NAND2_X1 U16113 ( .A1(n12975), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12911) );
  OAI211_X1 U16114 ( .C1(n13771), .C2(P1_EBX_REG_4__SCAN_IN), .A(n12911), .B(
        n12976), .ZN(n12912) );
  OAI21_X1 U16115 ( .B1(n12952), .B2(P1_EBX_REG_4__SCAN_IN), .A(n12912), .ZN(
        n13989) );
  NAND2_X1 U16116 ( .A1(n12976), .A2(n12913), .ZN(n12914) );
  OAI211_X1 U16117 ( .C1(n13771), .C2(P1_EBX_REG_5__SCAN_IN), .A(n12975), .B(
        n12914), .ZN(n12916) );
  INV_X1 U16118 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n21376) );
  NAND2_X1 U16119 ( .A1(n12916), .A2(n12915), .ZN(n14017) );
  MUX2_X1 U16120 ( .A(n12974), .B(n12983), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n12918) );
  NOR2_X1 U16121 ( .A1(n13686), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12917) );
  NOR2_X1 U16122 ( .A1(n12918), .A2(n12917), .ZN(n14049) );
  AND2_X1 U16123 ( .A1(n13771), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12919) );
  NOR2_X1 U16124 ( .A1(n12920), .A2(n12919), .ZN(n14130) );
  INV_X1 U16125 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16141) );
  NAND2_X1 U16126 ( .A1(n12921), .A2(n16141), .ZN(n12922) );
  NAND2_X1 U16127 ( .A1(n9938), .A2(n12922), .ZN(n14184) );
  NAND2_X1 U16128 ( .A1(n12976), .A2(n16126), .ZN(n12923) );
  OAI211_X1 U16129 ( .C1(n13771), .C2(P1_EBX_REG_9__SCAN_IN), .A(n12975), .B(
        n12923), .ZN(n12925) );
  INV_X1 U16130 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n21142) );
  NAND2_X1 U16131 ( .A1(n12925), .A2(n12924), .ZN(n14194) );
  NAND2_X1 U16132 ( .A1(n12975), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12926) );
  OAI211_X1 U16133 ( .C1(n13771), .C2(P1_EBX_REG_10__SCAN_IN), .A(n12926), .B(
        n12976), .ZN(n12927) );
  OAI21_X1 U16134 ( .B1(n12952), .B2(P1_EBX_REG_10__SCAN_IN), .A(n12927), .ZN(
        n14189) );
  MUX2_X1 U16135 ( .A(n12983), .B(n12953), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n12929) );
  AND2_X1 U16136 ( .A1(n13771), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12928) );
  NAND2_X1 U16137 ( .A1(n12975), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12930) );
  OAI211_X1 U16138 ( .C1(n13771), .C2(P1_EBX_REG_12__SCAN_IN), .A(n12930), .B(
        n12976), .ZN(n12931) );
  OAI21_X1 U16139 ( .B1(n12952), .B2(P1_EBX_REG_12__SCAN_IN), .A(n12931), .ZN(
        n15935) );
  NAND2_X1 U16140 ( .A1(n12976), .A2(n14812), .ZN(n12932) );
  OAI211_X1 U16141 ( .C1(n13771), .C2(P1_EBX_REG_13__SCAN_IN), .A(n12975), .B(
        n12932), .ZN(n12934) );
  INV_X1 U16142 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n21299) );
  NAND2_X1 U16143 ( .A1(n12934), .A2(n12933), .ZN(n14444) );
  MUX2_X1 U16144 ( .A(n12974), .B(n12983), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n12936) );
  NOR2_X1 U16145 ( .A1(n13686), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12935) );
  NOR2_X1 U16146 ( .A1(n12936), .A2(n12935), .ZN(n15916) );
  INV_X1 U16147 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n21197) );
  NAND2_X1 U16148 ( .A1(n12974), .A2(n21197), .ZN(n12939) );
  NAND2_X1 U16149 ( .A1(n12975), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12937) );
  OAI211_X1 U16150 ( .C1(n13771), .C2(P1_EBX_REG_16__SCAN_IN), .A(n12937), .B(
        n12976), .ZN(n12938) );
  AND2_X1 U16151 ( .A1(n12939), .A2(n12938), .ZN(n15896) );
  MUX2_X1 U16152 ( .A(n12975), .B(n12976), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n12941) );
  NAND2_X1 U16153 ( .A1(n13771), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12940) );
  NAND2_X1 U16154 ( .A1(n12941), .A2(n12940), .ZN(n15897) );
  INV_X1 U16155 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14798) );
  NAND2_X1 U16156 ( .A1(n12976), .A2(n14798), .ZN(n12942) );
  OAI211_X1 U16157 ( .C1(n13771), .C2(P1_EBX_REG_17__SCAN_IN), .A(n12975), .B(
        n12942), .ZN(n12944) );
  INV_X1 U16158 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n21097) );
  NAND2_X1 U16159 ( .A1(n12944), .A2(n12943), .ZN(n14403) );
  NAND2_X1 U16160 ( .A1(n12975), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12945) );
  OAI211_X1 U16161 ( .C1(n13771), .C2(P1_EBX_REG_18__SCAN_IN), .A(n12945), .B(
        n12976), .ZN(n12946) );
  OAI21_X1 U16162 ( .B1(n12952), .B2(P1_EBX_REG_18__SCAN_IN), .A(n12946), .ZN(
        n14802) );
  AND2_X1 U16163 ( .A1(n13771), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12947) );
  NOR2_X1 U16164 ( .A1(n12948), .A2(n12947), .ZN(n14425) );
  INV_X1 U16165 ( .A(n14425), .ZN(n12949) );
  NAND2_X1 U16166 ( .A1(n12975), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12950) );
  OAI211_X1 U16167 ( .C1(n13771), .C2(P1_EBX_REG_20__SCAN_IN), .A(n12950), .B(
        n12976), .ZN(n12951) );
  OAI21_X1 U16168 ( .B1(n12952), .B2(P1_EBX_REG_20__SCAN_IN), .A(n12951), .ZN(
        n15856) );
  MUX2_X1 U16169 ( .A(n12983), .B(n12953), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n12955) );
  AND2_X1 U16170 ( .A1(n13771), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12954) );
  NOR2_X1 U16171 ( .A1(n12955), .A2(n12954), .ZN(n14387) );
  NOR2_X1 U16172 ( .A1(n13686), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12956) );
  NOR2_X1 U16173 ( .A1(n12957), .A2(n12956), .ZN(n14374) );
  INV_X1 U16174 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14611) );
  NAND2_X1 U16175 ( .A1(n12976), .A2(n14611), .ZN(n12958) );
  OAI211_X1 U16176 ( .C1(n13771), .C2(P1_EBX_REG_23__SCAN_IN), .A(n12975), .B(
        n12958), .ZN(n12960) );
  INV_X1 U16177 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n21195) );
  NAND2_X1 U16178 ( .A1(n12983), .A2(n21195), .ZN(n12959) );
  NAND2_X1 U16179 ( .A1(n12960), .A2(n12959), .ZN(n14364) );
  INV_X1 U16180 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n21363) );
  NAND2_X1 U16181 ( .A1(n12974), .A2(n21363), .ZN(n12963) );
  NAND2_X1 U16182 ( .A1(n12975), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12961) );
  OAI211_X1 U16183 ( .C1(n13771), .C2(P1_EBX_REG_24__SCAN_IN), .A(n12961), .B(
        n12976), .ZN(n12962) );
  INV_X1 U16184 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n12964) );
  NAND2_X1 U16185 ( .A1(n12974), .A2(n12964), .ZN(n12967) );
  NAND2_X1 U16186 ( .A1(n12975), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12965) );
  OAI211_X1 U16187 ( .C1(n13771), .C2(P1_EBX_REG_26__SCAN_IN), .A(n12965), .B(
        n12976), .ZN(n12966) );
  AND2_X1 U16188 ( .A1(n12967), .A2(n12966), .ZN(n14326) );
  MUX2_X1 U16189 ( .A(n12975), .B(n12976), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n12969) );
  NAND2_X1 U16190 ( .A1(n13771), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12968) );
  NAND2_X1 U16191 ( .A1(n12969), .A2(n12968), .ZN(n14339) );
  NAND2_X1 U16192 ( .A1(n14326), .A2(n14339), .ZN(n12970) );
  INV_X1 U16193 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14573) );
  NAND2_X1 U16194 ( .A1(n12976), .A2(n14573), .ZN(n12971) );
  OAI211_X1 U16195 ( .C1(n13771), .C2(P1_EBX_REG_27__SCAN_IN), .A(n12975), .B(
        n12971), .ZN(n12973) );
  INV_X1 U16196 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n21313) );
  INV_X1 U16197 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n21315) );
  NAND2_X1 U16198 ( .A1(n12974), .A2(n21315), .ZN(n12979) );
  NAND2_X1 U16199 ( .A1(n12975), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12977) );
  OAI211_X1 U16200 ( .C1(n13771), .C2(P1_EBX_REG_28__SCAN_IN), .A(n12977), .B(
        n12976), .ZN(n12978) );
  AND2_X1 U16201 ( .A1(n12979), .A2(n12978), .ZN(n14301) );
  OR2_X1 U16202 ( .A1(n13771), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n12980) );
  OAI21_X1 U16203 ( .B1(n13686), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n12980), .ZN(n13030) );
  INV_X1 U16204 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n21410) );
  NAND2_X1 U16205 ( .A1(n12982), .A2(n12981), .ZN(n14293) );
  NAND2_X1 U16206 ( .A1(n14303), .A2(n14293), .ZN(n14292) );
  NOR2_X1 U16207 ( .A1(n13033), .A2(n12989), .ZN(n12988) );
  INV_X1 U16208 ( .A(n14292), .ZN(n12986) );
  NAND2_X1 U16209 ( .A1(n13686), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n12985) );
  NAND2_X1 U16210 ( .A1(n13771), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12984) );
  NAND2_X1 U16211 ( .A1(n12985), .A2(n12984), .ZN(n13034) );
  NAND2_X1 U16212 ( .A1(n12986), .A2(n13034), .ZN(n12987) );
  NAND2_X1 U16213 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21064) );
  NAND2_X1 U16214 ( .A1(n21064), .A2(n20848), .ZN(n15825) );
  NAND3_X1 U16215 ( .A1(n13485), .A2(P1_EBX_REG_31__SCAN_IN), .A3(n15825), 
        .ZN(n12990) );
  NAND2_X1 U16216 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n12997) );
  INV_X1 U16217 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20999) );
  NAND2_X1 U16218 ( .A1(n12992), .A2(n20999), .ZN(n21073) );
  NAND2_X1 U16219 ( .A1(n13753), .A2(n21073), .ZN(n13759) );
  INV_X1 U16220 ( .A(n15825), .ZN(n12993) );
  NAND2_X1 U16221 ( .A1(n13759), .A2(n12993), .ZN(n12998) );
  NOR2_X1 U16222 ( .A1(n12998), .A2(n11918), .ZN(n12994) );
  INV_X1 U16223 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n21310) );
  NOR2_X1 U16224 ( .A1(n21310), .A2(n21412), .ZN(n12996) );
  NAND3_X1 U16225 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .A3(P1_REIP_REG_24__SCAN_IN), .ZN(n12995) );
  AND3_X1 U16226 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(P1_REIP_REG_21__SCAN_IN), 
        .A3(P1_REIP_REG_23__SCAN_IN), .ZN(n13004) );
  NAND3_X1 U16227 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(P1_REIP_REG_19__SCAN_IN), 
        .A3(P1_REIP_REG_18__SCAN_IN), .ZN(n14373) );
  INV_X1 U16228 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n21341) );
  INV_X1 U16229 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21382) );
  INV_X1 U16230 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n21384) );
  INV_X1 U16231 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n21019) );
  INV_X1 U16232 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21379) );
  NAND3_X1 U16233 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .ZN(n20274) );
  NOR2_X1 U16234 ( .A1(n21332), .A2(n20274), .ZN(n20275) );
  NAND3_X1 U16235 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(n20275), .ZN(n20227) );
  NOR3_X1 U16236 ( .A1(n21019), .A2(n21379), .A3(n20227), .ZN(n13003) );
  NAND2_X1 U16237 ( .A1(n13003), .A2(n14408), .ZN(n20202) );
  NOR3_X1 U16238 ( .A1(n21384), .A2(n21381), .A3(n20202), .ZN(n15952) );
  NAND3_X1 U16239 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .A3(n15952), .ZN(n15926) );
  NOR3_X1 U16240 ( .A1(n21341), .A2(n21382), .A3(n15926), .ZN(n15895) );
  NAND4_X1 U16241 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .A3(P1_REIP_REG_16__SCAN_IN), .A4(n15895), .ZN(n14397) );
  OAI21_X1 U16242 ( .B1(n14373), .B2(n14397), .A(n20250), .ZN(n15875) );
  OAI21_X1 U16243 ( .B1(n15951), .B2(n13004), .A(n15875), .ZN(n14368) );
  AOI21_X1 U16244 ( .B1(n12995), .B2(n20250), .A(n14368), .ZN(n14333) );
  OAI21_X1 U16245 ( .B1(n15951), .B2(n12996), .A(n14333), .ZN(n14304) );
  AOI21_X1 U16246 ( .B1(n12997), .B2(n20250), .A(n14304), .ZN(n14288) );
  INV_X1 U16247 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n21048) );
  INV_X1 U16248 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n21300) );
  OAI211_X1 U16249 ( .C1(n13753), .C2(n21300), .A(n12998), .B(n20380), .ZN(
        n12999) );
  INV_X1 U16250 ( .A(n12999), .ZN(n13000) );
  AND2_X2 U16251 ( .A1(n14408), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20255) );
  AOI22_X1 U16252 ( .A1(n20292), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n20255), .ZN(n13001) );
  OAI21_X1 U16253 ( .B1(n14288), .B2(n21048), .A(n13001), .ZN(n13002) );
  AOI21_X1 U16254 ( .B1(n14418), .B2(n20272), .A(n13002), .ZN(n13007) );
  INV_X1 U16255 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n21302) );
  NAND2_X1 U16256 ( .A1(n20285), .A2(n13003), .ZN(n20210) );
  NAND2_X1 U16257 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n15963), .ZN(n15955) );
  NAND2_X1 U16258 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(n15939), .ZN(n15934) );
  NAND2_X1 U16259 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n15920), .ZN(n15915) );
  NAND2_X1 U16260 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n15894) );
  INV_X1 U16261 ( .A(n14373), .ZN(n14367) );
  NAND2_X1 U16262 ( .A1(n14367), .A2(n13004), .ZN(n13005) );
  NAND4_X1 U16263 ( .A1(n14357), .A2(P1_REIP_REG_25__SCAN_IN), .A3(
        P1_REIP_REG_24__SCAN_IN), .A4(P1_REIP_REG_26__SCAN_IN), .ZN(n14319) );
  NOR3_X1 U16264 ( .A1(n14319), .A2(n21412), .A3(n21310), .ZN(n14298) );
  NAND4_X1 U16265 ( .A1(n14298), .A2(P1_REIP_REG_29__SCAN_IN), .A3(
        P1_REIP_REG_30__SCAN_IN), .A4(n21048), .ZN(n13006) );
  OAI21_X1 U16266 ( .B1(n14554), .B2(n15960), .A(n13008), .ZN(P1_U2809) );
  INV_X1 U16267 ( .A(n15788), .ZN(n13009) );
  NOR2_X1 U16268 ( .A1(n13009), .A2(n17633), .ZN(n16530) );
  AOI21_X1 U16269 ( .B1(n13010), .B2(n17797), .A(n17640), .ZN(n17625) );
  AOI22_X1 U16270 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17886), .B1(
        n17797), .B2(n15781), .ZN(n17624) );
  NOR2_X1 U16271 ( .A1(n17625), .A2(n17624), .ZN(n17623) );
  INV_X1 U16272 ( .A(n17623), .ZN(n13015) );
  AOI21_X1 U16273 ( .B1(n17641), .B2(n17797), .A(n13017), .ZN(n13014) );
  NAND2_X1 U16274 ( .A1(n15788), .A2(n17997), .ZN(n16518) );
  OAI21_X1 U16275 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18202), .A(
        n13011), .ZN(n15780) );
  AOI21_X1 U16276 ( .B1(n16518), .B2(n18229), .A(n15780), .ZN(n13012) );
  NAND2_X1 U16277 ( .A1(n17797), .A2(n17641), .ZN(n13016) );
  NAND2_X1 U16278 ( .A1(n9802), .A2(n18779), .ZN(n18311) );
  NOR2_X1 U16279 ( .A1(n13016), .A2(n18311), .ZN(n13018) );
  NAND2_X1 U16280 ( .A1(n18308), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17628) );
  AOI22_X1 U16281 ( .A1(n18231), .A2(n18184), .B1(n18229), .B2(n18186), .ZN(
        n18098) );
  OAI21_X1 U16282 ( .B1(n18098), .B2(n18099), .A(n13020), .ZN(n18042) );
  NAND2_X1 U16283 ( .A1(n9802), .A2(n18042), .ZN(n18068) );
  NAND2_X1 U16284 ( .A1(n13021), .A2(n15781), .ZN(n17637) );
  INV_X1 U16285 ( .A(n14563), .ZN(n14459) );
  AND2_X1 U16286 ( .A1(n13485), .A2(n10115), .ZN(n13025) );
  NAND2_X1 U16287 ( .A1(n13751), .A2(n13914), .ZN(n13617) );
  INV_X1 U16288 ( .A(n20443), .ZN(n14455) );
  NAND4_X1 U16289 ( .A1(n13026), .A2(n9823), .A3(n14455), .A4(n11928), .ZN(
        n13027) );
  NOR2_X1 U16290 ( .A1(n13027), .A2(n13923), .ZN(n13045) );
  NAND2_X1 U16291 ( .A1(n13045), .A2(n13485), .ZN(n13028) );
  NAND2_X1 U16292 ( .A1(n13617), .A2(n13028), .ZN(n13029) );
  INV_X1 U16293 ( .A(n13030), .ZN(n13031) );
  AND2_X1 U16294 ( .A1(n14303), .A2(n13031), .ZN(n13032) );
  INV_X1 U16295 ( .A(n13034), .ZN(n13035) );
  XNOR2_X1 U16296 ( .A(n13036), .B(n13035), .ZN(n14727) );
  INV_X1 U16297 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n21385) );
  NOR2_X1 U16298 ( .A1(n20306), .A2(n21385), .ZN(n13037) );
  AOI21_X1 U16299 ( .B1(n14727), .B2(n13038), .A(n13037), .ZN(n13039) );
  INV_X1 U16300 ( .A(n21064), .ZN(n16146) );
  NOR2_X1 U16301 ( .A1(n13482), .A2(n11916), .ZN(n13041) );
  NAND2_X1 U16302 ( .A1(n13750), .A2(n13041), .ZN(n13912) );
  OAI21_X1 U16303 ( .B1(n13040), .B2(n16146), .A(n13912), .ZN(n13042) );
  NAND2_X1 U16304 ( .A1(n13042), .A2(n13764), .ZN(n13049) );
  NOR2_X1 U16305 ( .A1(n16146), .A2(n13480), .ZN(n13752) );
  INV_X1 U16306 ( .A(n13752), .ZN(n13044) );
  NAND2_X1 U16307 ( .A1(n13045), .A2(n14026), .ZN(n13046) );
  NAND2_X1 U16308 ( .A1(n13618), .A2(n13046), .ZN(n13047) );
  AND2_X1 U16309 ( .A1(n14527), .A2(n14455), .ZN(n13050) );
  NAND2_X1 U16310 ( .A1(n13051), .A2(n13050), .ZN(n13069) );
  NOR4_X1 U16311 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n13055) );
  NOR4_X1 U16312 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n13054) );
  NOR4_X1 U16313 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13053) );
  NOR4_X1 U16314 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n13052) );
  AND4_X1 U16315 ( .A1(n13055), .A2(n13054), .A3(n13053), .A4(n13052), .ZN(
        n13060) );
  NOR4_X1 U16316 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n13058) );
  NOR4_X1 U16317 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n13057) );
  NOR4_X1 U16318 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n13056) );
  INV_X1 U16319 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n21011) );
  AND4_X1 U16320 ( .A1(n13058), .A2(n13057), .A3(n13056), .A4(n21011), .ZN(
        n13059) );
  NAND2_X1 U16321 ( .A1(n13060), .A2(n13059), .ZN(n13061) );
  NOR3_X1 U16322 ( .A1(n14532), .A2(n20373), .A3(n13760), .ZN(n13062) );
  AOI22_X1 U16323 ( .A1(n14506), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14532), .ZN(n13063) );
  INV_X1 U16324 ( .A(n13063), .ZN(n13067) );
  INV_X1 U16325 ( .A(n20373), .ZN(n20372) );
  NOR2_X1 U16326 ( .A1(n13760), .A2(n20372), .ZN(n13064) );
  NAND2_X1 U16327 ( .A1(n14527), .A2(n13064), .ZN(n14454) );
  INV_X1 U16328 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n13065) );
  NOR2_X1 U16329 ( .A1(n14454), .A2(n13065), .ZN(n13066) );
  NOR2_X1 U16330 ( .A1(n13067), .A2(n13066), .ZN(n13068) );
  NAND2_X1 U16331 ( .A1(n13069), .A2(n13068), .ZN(P1_U2873) );
  NAND2_X1 U16332 ( .A1(n9833), .A2(n13537), .ZN(n13074) );
  NAND2_X1 U16333 ( .A1(n13070), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13071) );
  NAND2_X1 U16334 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19924) );
  INV_X1 U16335 ( .A(n19924), .ZN(n19965) );
  OAI21_X1 U16336 ( .B1(n13082), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n20126), .ZN(n13072) );
  NOR2_X1 U16337 ( .A1(n13072), .A2(n20017), .ZN(n19860) );
  AOI21_X1 U16338 ( .B1(n13092), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19860), .ZN(n13073) );
  NAND2_X1 U16339 ( .A1(n13074), .A2(n13073), .ZN(n13079) );
  NOR2_X1 U16340 ( .A1(n13332), .A2(n19462), .ZN(n13078) );
  NAND2_X1 U16341 ( .A1(n13079), .A2(n13078), .ZN(n13103) );
  OAI21_X1 U16342 ( .B1(n13079), .B2(n13078), .A(n13103), .ZN(n13080) );
  NAND2_X1 U16343 ( .A1(n13081), .A2(n13537), .ZN(n13086) );
  NAND2_X1 U16344 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19829) );
  NAND2_X1 U16345 ( .A1(n19829), .A2(n20147), .ZN(n13084) );
  INV_X1 U16346 ( .A(n13082), .ZN(n13083) );
  AND2_X1 U16347 ( .A1(n13084), .A2(n13083), .ZN(n19609) );
  AOI22_X1 U16348 ( .A1(n13092), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n20126), .B2(n19609), .ZN(n13085) );
  NAND2_X1 U16349 ( .A1(n13086), .A2(n13085), .ZN(n13088) );
  INV_X1 U16350 ( .A(n13746), .ZN(n13099) );
  AOI22_X1 U16351 ( .A1(n13092), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20126), .B2(n20165), .ZN(n13090) );
  NAND2_X1 U16352 ( .A1(n13092), .A2(n15662), .ZN(n13093) );
  NAND2_X1 U16353 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20165), .ZN(
        n19795) );
  NAND2_X1 U16354 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n16450), .ZN(
        n19763) );
  NAND2_X1 U16355 ( .A1(n19795), .A2(n19763), .ZN(n19671) );
  NAND2_X1 U16356 ( .A1(n20126), .A2(n19671), .ZN(n19797) );
  NAND2_X1 U16357 ( .A1(n13093), .A2(n19797), .ZN(n13094) );
  NAND2_X1 U16358 ( .A1(n13589), .A2(n13590), .ZN(n13098) );
  NAND2_X1 U16359 ( .A1(n15643), .A2(n13096), .ZN(n13097) );
  NAND2_X1 U16360 ( .A1(n13099), .A2(n10385), .ZN(n13101) );
  NAND2_X1 U16361 ( .A1(n13070), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13102) );
  AND2_X1 U16362 ( .A1(n13103), .A2(n13102), .ZN(n13104) );
  NOR2_X1 U16363 ( .A1(n13332), .A2(n19468), .ZN(n19210) );
  NAND2_X1 U16364 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13872) );
  NOR2_X1 U16365 ( .A1(n13105), .A2(n13872), .ZN(n19282) );
  NAND2_X1 U16366 ( .A1(n9949), .A2(n13110), .ZN(n14174) );
  AOI22_X1 U16367 ( .A1(n10688), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10689), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13114) );
  AOI22_X1 U16368 ( .A1(n10650), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13187), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13113) );
  AOI22_X1 U16369 ( .A1(n13218), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13219), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13112) );
  AOI22_X1 U16370 ( .A1(n13220), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13217), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13111) );
  NAND4_X1 U16371 ( .A1(n13114), .A2(n13113), .A3(n13112), .A4(n13111), .ZN(
        n13122) );
  INV_X1 U16372 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13115) );
  OAI22_X1 U16373 ( .A1(n13178), .A2(n19446), .B1(n13177), .B2(n13115), .ZN(
        n13116) );
  AOI21_X1 U16374 ( .B1(n13141), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n13116), .ZN(n13120) );
  AOI22_X1 U16375 ( .A1(n10728), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10748), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13119) );
  AOI22_X1 U16376 ( .A1(n13225), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13226), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13118) );
  NAND2_X1 U16377 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n13117) );
  NAND4_X1 U16378 ( .A1(n13120), .A2(n13119), .A3(n13118), .A4(n13117), .ZN(
        n13121) );
  NOR2_X1 U16379 ( .A1(n13122), .A2(n13121), .ZN(n19257) );
  AOI22_X1 U16380 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10688), .B1(
        n10689), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13126) );
  AOI22_X1 U16381 ( .A1(n10650), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13187), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13125) );
  AOI22_X1 U16382 ( .A1(n13218), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13219), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13124) );
  AOI22_X1 U16383 ( .A1(n13220), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13217), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13123) );
  NAND4_X1 U16384 ( .A1(n13126), .A2(n13125), .A3(n13124), .A4(n13123), .ZN(
        n13134) );
  INV_X1 U16385 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19452) );
  OAI22_X1 U16386 ( .A1(n13178), .A2(n19452), .B1(n13177), .B2(n13127), .ZN(
        n13128) );
  AOI21_X1 U16387 ( .B1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n13141), .A(
        n13128), .ZN(n13132) );
  AOI22_X1 U16388 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10728), .B1(
        n10748), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13131) );
  AOI22_X1 U16389 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n13225), .B1(
        n13226), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13130) );
  NAND2_X1 U16390 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n13129) );
  NAND4_X1 U16391 ( .A1(n13132), .A2(n13131), .A3(n13130), .A4(n13129), .ZN(
        n13133) );
  OR2_X1 U16392 ( .A1(n13134), .A2(n13133), .ZN(n15015) );
  AND2_X2 U16393 ( .A1(n15014), .A2(n15015), .ZN(n15013) );
  AOI22_X1 U16394 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10688), .B1(
        n10689), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13138) );
  AOI22_X1 U16395 ( .A1(n10650), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13187), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13137) );
  AOI22_X1 U16396 ( .A1(n13218), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13219), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13136) );
  AOI22_X1 U16397 ( .A1(n13220), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13217), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13135) );
  NAND4_X1 U16398 ( .A1(n13138), .A2(n13137), .A3(n13136), .A4(n13135), .ZN(
        n13147) );
  INV_X1 U16399 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13139) );
  OAI22_X1 U16400 ( .A1(n13178), .A2(n19457), .B1(n13177), .B2(n13139), .ZN(
        n13140) );
  AOI21_X1 U16401 ( .B1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n13141), .A(
        n13140), .ZN(n13145) );
  AOI22_X1 U16402 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10728), .B1(
        n10748), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13144) );
  AOI22_X1 U16403 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n13225), .B1(
        n13226), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13143) );
  NAND2_X1 U16404 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n13142) );
  NAND4_X1 U16405 ( .A1(n13145), .A2(n13144), .A3(n13143), .A4(n13142), .ZN(
        n13146) );
  OR2_X1 U16406 ( .A1(n13147), .A2(n13146), .ZN(n16273) );
  AOI22_X1 U16407 ( .A1(n10688), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10689), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13151) );
  AOI22_X1 U16408 ( .A1(n10650), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13187), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13150) );
  AOI22_X1 U16409 ( .A1(n13218), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13219), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13149) );
  AOI22_X1 U16410 ( .A1(n13220), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13217), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13148) );
  NAND4_X1 U16411 ( .A1(n13151), .A2(n13150), .A3(n13149), .A4(n13148), .ZN(
        n13159) );
  INV_X1 U16412 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13152) );
  OAI22_X1 U16413 ( .A1(n13178), .A2(n13871), .B1(n13177), .B2(n13152), .ZN(
        n13153) );
  AOI21_X1 U16414 ( .B1(n13141), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n13153), .ZN(n13157) );
  AOI22_X1 U16415 ( .A1(n10728), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10748), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13156) );
  AOI22_X1 U16416 ( .A1(n13225), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13226), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13155) );
  NAND2_X1 U16417 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n13154) );
  NAND4_X1 U16418 ( .A1(n13157), .A2(n13156), .A3(n13155), .A4(n13154), .ZN(
        n13158) );
  OR2_X1 U16419 ( .A1(n13159), .A2(n13158), .ZN(n15003) );
  AOI22_X1 U16420 ( .A1(n10688), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10689), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13163) );
  AOI22_X1 U16421 ( .A1(n10650), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13187), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13162) );
  AOI22_X1 U16422 ( .A1(n13218), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13219), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13161) );
  AOI22_X1 U16423 ( .A1(n13220), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13217), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13160) );
  NAND4_X1 U16424 ( .A1(n13163), .A2(n13162), .A3(n13161), .A4(n13160), .ZN(
        n13171) );
  INV_X1 U16425 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13164) );
  OAI22_X1 U16426 ( .A1(n13178), .A2(n19468), .B1(n13177), .B2(n13164), .ZN(
        n13165) );
  AOI21_X1 U16427 ( .B1(n13141), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A(
        n13165), .ZN(n13169) );
  AOI22_X1 U16428 ( .A1(n10728), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10748), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13168) );
  AOI22_X1 U16429 ( .A1(n13225), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13226), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13167) );
  NAND2_X1 U16430 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n13166) );
  NAND4_X1 U16431 ( .A1(n13169), .A2(n13168), .A3(n13167), .A4(n13166), .ZN(
        n13170) );
  NOR2_X1 U16432 ( .A1(n13171), .A2(n13170), .ZN(n16271) );
  AOI22_X1 U16433 ( .A1(n10688), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10689), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13175) );
  AOI22_X1 U16434 ( .A1(n10650), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13187), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13174) );
  AOI22_X1 U16435 ( .A1(n13218), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13219), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13173) );
  AOI22_X1 U16436 ( .A1(n13220), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13217), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13172) );
  NAND4_X1 U16437 ( .A1(n13175), .A2(n13174), .A3(n13173), .A4(n13172), .ZN(
        n13185) );
  INV_X1 U16438 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13176) );
  OAI22_X1 U16439 ( .A1(n13178), .A2(n19462), .B1(n13177), .B2(n13176), .ZN(
        n13179) );
  AOI21_X1 U16440 ( .B1(n13141), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n13179), .ZN(n13183) );
  AOI22_X1 U16441 ( .A1(n10728), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10748), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13182) );
  AOI22_X1 U16442 ( .A1(n13225), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13226), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13181) );
  NAND2_X1 U16443 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n13180) );
  NAND4_X1 U16444 ( .A1(n13183), .A2(n13182), .A3(n13181), .A4(n13180), .ZN(
        n13184) );
  NOR2_X1 U16445 ( .A1(n13185), .A2(n13184), .ZN(n15007) );
  NOR2_X1 U16446 ( .A1(n16271), .A2(n15007), .ZN(n15002) );
  AND2_X1 U16447 ( .A1(n15003), .A2(n15002), .ZN(n13186) );
  AOI22_X1 U16448 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10688), .B1(
        n10689), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13191) );
  AOI22_X1 U16449 ( .A1(n10650), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13187), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13190) );
  AOI22_X1 U16450 ( .A1(n13218), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13219), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13189) );
  AOI22_X1 U16451 ( .A1(n13220), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10649), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13188) );
  NAND4_X1 U16452 ( .A1(n13191), .A2(n13190), .A3(n13189), .A4(n13188), .ZN(
        n13200) );
  INV_X1 U16453 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13194) );
  AOI22_X1 U16454 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n13225), .B1(
        n13226), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13193) );
  AOI22_X1 U16455 ( .A1(n13227), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n13228), .ZN(n13192) );
  OAI211_X1 U16456 ( .C1(n13194), .C2(n9846), .A(n13193), .B(n13192), .ZN(
        n13199) );
  INV_X1 U16457 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13197) );
  INV_X1 U16458 ( .A(n10665), .ZN(n13196) );
  AOI22_X1 U16459 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n10748), .B1(
        n10728), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13195) );
  OAI21_X1 U16460 ( .B1(n13197), .B2(n13196), .A(n13195), .ZN(n13198) );
  NOR3_X1 U16461 ( .A1(n13200), .A2(n13199), .A3(n13198), .ZN(n16266) );
  AOI22_X1 U16462 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13391), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13208) );
  AOI22_X1 U16463 ( .A1(n9815), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(n9834), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13207) );
  AOI22_X1 U16464 ( .A1(n10632), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9817), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13206) );
  INV_X1 U16465 ( .A(n10421), .ZN(n13388) );
  INV_X1 U16466 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13203) );
  OAI21_X2 U16467 ( .B1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n13201), .ZN(n13390) );
  NAND2_X1 U16468 ( .A1(n13320), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n13202) );
  OAI211_X1 U16469 ( .C1(n13388), .C2(n13203), .A(n13390), .B(n13202), .ZN(
        n13204) );
  INV_X1 U16470 ( .A(n13204), .ZN(n13205) );
  NAND4_X1 U16471 ( .A1(n13208), .A2(n13207), .A3(n13206), .A4(n13205), .ZN(
        n13216) );
  AOI22_X1 U16472 ( .A1(n9840), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9842), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13214) );
  AOI22_X1 U16473 ( .A1(n10634), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13320), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13213) );
  AOI22_X1 U16474 ( .A1(n10632), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9815), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13212) );
  NAND2_X1 U16475 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n13210) );
  AOI21_X1 U16476 ( .B1(n10482), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A(
        n13390), .ZN(n13209) );
  AND2_X1 U16477 ( .A1(n13210), .A2(n13209), .ZN(n13211) );
  NAND4_X1 U16478 ( .A1(n13214), .A2(n13213), .A3(n13212), .A4(n13211), .ZN(
        n13215) );
  AND2_X1 U16479 ( .A1(n13216), .A2(n13215), .ZN(n13261) );
  NAND2_X1 U16480 ( .A1(n19447), .A2(n13261), .ZN(n13239) );
  AOI22_X1 U16481 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10688), .B1(
        n10689), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13224) );
  AOI22_X1 U16482 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n13141), .B1(
        n10650), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13223) );
  AOI22_X1 U16483 ( .A1(n13218), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13217), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13222) );
  AOI22_X1 U16484 ( .A1(n13220), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13219), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13221) );
  NAND4_X1 U16485 ( .A1(n13224), .A2(n13223), .A3(n13222), .A4(n13221), .ZN(
        n13238) );
  AOI22_X1 U16486 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n13225), .B1(
        n10728), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13236) );
  AOI22_X1 U16487 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n10748), .B1(
        n13226), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13235) );
  INV_X1 U16488 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13378) );
  NAND2_X1 U16489 ( .A1(n13227), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n13230) );
  NAND2_X1 U16490 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n13228), .ZN(
        n13229) );
  OAI211_X1 U16491 ( .C1(n13231), .C2(n13378), .A(n13230), .B(n13229), .ZN(
        n13232) );
  INV_X1 U16492 ( .A(n13232), .ZN(n13234) );
  NAND2_X1 U16493 ( .A1(n10665), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n13233) );
  NAND4_X1 U16494 ( .A1(n13236), .A2(n13235), .A3(n13234), .A4(n13233), .ZN(
        n13237) );
  XNOR2_X1 U16495 ( .A(n13239), .B(n13258), .ZN(n13264) );
  NAND2_X1 U16496 ( .A1(n10527), .A2(n13261), .ZN(n15074) );
  NOR2_X2 U16497 ( .A1(n15072), .A2(n15074), .ZN(n15073) );
  AOI22_X1 U16498 ( .A1(n10632), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10633), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13248) );
  INV_X1 U16499 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13243) );
  OAI21_X1 U16500 ( .B1(n13242), .B2(n13243), .A(n13390), .ZN(n13244) );
  AOI21_X1 U16501 ( .B1(n9807), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A(n13244), .ZN(n13247) );
  AOI22_X1 U16502 ( .A1(n9817), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13246) );
  AOI22_X1 U16503 ( .A1(n9840), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n16444), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13245) );
  NAND4_X1 U16504 ( .A1(n13248), .A2(n13247), .A3(n13246), .A4(n13245), .ZN(
        n13257) );
  AOI22_X1 U16505 ( .A1(n10632), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10633), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13255) );
  AOI22_X1 U16506 ( .A1(n9816), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13254) );
  AOI22_X1 U16507 ( .A1(n9840), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n16444), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13253) );
  NAND2_X1 U16508 ( .A1(n9808), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n13251) );
  AOI21_X1 U16509 ( .B1(n13320), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A(
        n13390), .ZN(n13250) );
  AND2_X1 U16510 ( .A1(n13251), .A2(n13250), .ZN(n13252) );
  NAND4_X1 U16511 ( .A1(n13255), .A2(n13254), .A3(n13253), .A4(n13252), .ZN(
        n13256) );
  NAND2_X1 U16512 ( .A1(n13257), .A2(n13256), .ZN(n13260) );
  NAND2_X1 U16513 ( .A1(n13258), .A2(n13261), .ZN(n13265) );
  XOR2_X1 U16514 ( .A(n13260), .B(n13265), .Z(n13259) );
  NAND2_X1 U16515 ( .A1(n13259), .A2(n13304), .ZN(n14993) );
  INV_X1 U16516 ( .A(n13260), .ZN(n13266) );
  NAND2_X1 U16517 ( .A1(n10536), .A2(n13266), .ZN(n14995) );
  INV_X1 U16518 ( .A(n13261), .ZN(n13262) );
  NOR2_X1 U16519 ( .A1(n14995), .A2(n13262), .ZN(n13263) );
  INV_X1 U16520 ( .A(n13265), .ZN(n13267) );
  NAND2_X1 U16521 ( .A1(n13267), .A2(n13266), .ZN(n13284) );
  AOI22_X1 U16522 ( .A1(n10632), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10633), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13274) );
  AOI22_X1 U16523 ( .A1(n10634), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13273) );
  AOI22_X1 U16524 ( .A1(n9840), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n16444), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13272) );
  INV_X1 U16525 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13269) );
  NAND2_X1 U16526 ( .A1(n13312), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n13268) );
  OAI211_X1 U16527 ( .C1(n13388), .C2(n13269), .A(n13390), .B(n13268), .ZN(
        n13270) );
  INV_X1 U16528 ( .A(n13270), .ZN(n13271) );
  NAND4_X1 U16529 ( .A1(n13274), .A2(n13273), .A3(n13272), .A4(n13271), .ZN(
        n13283) );
  AOI22_X1 U16530 ( .A1(n10632), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10633), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13281) );
  AOI22_X1 U16531 ( .A1(n9817), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9834), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13280) );
  AOI22_X1 U16532 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n16444), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13279) );
  INV_X1 U16533 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13276) );
  INV_X1 U16534 ( .A(n13390), .ZN(n13322) );
  NAND2_X1 U16535 ( .A1(n13320), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n13275) );
  OAI211_X1 U16536 ( .C1(n13388), .C2(n13276), .A(n13322), .B(n13275), .ZN(
        n13277) );
  INV_X1 U16537 ( .A(n13277), .ZN(n13278) );
  NAND4_X1 U16538 ( .A1(n13281), .A2(n13280), .A3(n13279), .A4(n13278), .ZN(
        n13282) );
  NAND2_X1 U16539 ( .A1(n13283), .A2(n13282), .ZN(n13286) );
  NAND2_X1 U16540 ( .A1(n13284), .A2(n13286), .ZN(n13285) );
  NAND3_X1 U16541 ( .A1(n13311), .A2(n13304), .A3(n13285), .ZN(n13287) );
  NOR2_X1 U16542 ( .A1(n19447), .A2(n13286), .ZN(n14986) );
  AOI22_X1 U16543 ( .A1(n10632), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10633), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13295) );
  INV_X1 U16544 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13290) );
  OAI21_X1 U16545 ( .B1(n13242), .B2(n13290), .A(n13390), .ZN(n13291) );
  AOI21_X1 U16546 ( .B1(n9808), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A(n13291), .ZN(n13294) );
  AOI22_X1 U16547 ( .A1(n9816), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13293) );
  AOI22_X1 U16548 ( .A1(n9840), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n16444), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13292) );
  NAND4_X1 U16549 ( .A1(n13295), .A2(n13294), .A3(n13293), .A4(n13292), .ZN(
        n13303) );
  AOI22_X1 U16550 ( .A1(n10632), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10633), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13301) );
  AOI22_X1 U16551 ( .A1(n9816), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9834), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13300) );
  AOI22_X1 U16552 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n16444), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13299) );
  NAND2_X1 U16553 ( .A1(n10421), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n13297) );
  AOI21_X1 U16554 ( .B1(n13320), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n13390), .ZN(n13296) );
  AND2_X1 U16555 ( .A1(n13297), .A2(n13296), .ZN(n13298) );
  NAND4_X1 U16556 ( .A1(n13301), .A2(n13300), .A3(n13299), .A4(n13298), .ZN(
        n13302) );
  AND2_X1 U16557 ( .A1(n13303), .A2(n13302), .ZN(n13306) );
  XNOR2_X1 U16558 ( .A(n13311), .B(n13306), .ZN(n13305) );
  NAND2_X1 U16559 ( .A1(n13305), .A2(n13304), .ZN(n13308) );
  INV_X1 U16560 ( .A(n13306), .ZN(n13310) );
  NOR2_X1 U16561 ( .A1(n19447), .A2(n13310), .ZN(n14978) );
  INV_X1 U16562 ( .A(n13307), .ZN(n13309) );
  NOR2_X1 U16563 ( .A1(n13311), .A2(n13310), .ZN(n13331) );
  INV_X1 U16564 ( .A(n13331), .ZN(n13334) );
  AOI22_X1 U16565 ( .A1(n10632), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10633), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13319) );
  AOI22_X1 U16566 ( .A1(n9817), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13318) );
  AOI22_X1 U16567 ( .A1(n9840), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n16444), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13317) );
  NAND2_X1 U16568 ( .A1(n13312), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n13313) );
  OAI211_X1 U16569 ( .C1(n13388), .C2(n13314), .A(n13390), .B(n13313), .ZN(
        n13315) );
  INV_X1 U16570 ( .A(n13315), .ZN(n13316) );
  NAND4_X1 U16571 ( .A1(n13319), .A2(n13318), .A3(n13317), .A4(n13316), .ZN(
        n13330) );
  AOI22_X1 U16572 ( .A1(n10632), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10633), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13328) );
  AOI22_X1 U16573 ( .A1(n9817), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9834), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13327) );
  AOI22_X1 U16574 ( .A1(n9840), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16444), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13326) );
  INV_X1 U16575 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13323) );
  NAND2_X1 U16576 ( .A1(n13320), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n13321) );
  OAI211_X1 U16577 ( .C1(n13388), .C2(n13323), .A(n13322), .B(n13321), .ZN(
        n13324) );
  INV_X1 U16578 ( .A(n13324), .ZN(n13325) );
  NAND4_X1 U16579 ( .A1(n13328), .A2(n13327), .A3(n13326), .A4(n13325), .ZN(
        n13329) );
  AND2_X1 U16580 ( .A1(n13330), .A2(n13329), .ZN(n13338) );
  INV_X1 U16581 ( .A(n13338), .ZN(n13333) );
  AOI211_X1 U16582 ( .C1(n13334), .C2(n13333), .A(n13332), .B(n14962), .ZN(
        n13335) );
  NAND2_X1 U16583 ( .A1(n13336), .A2(n13335), .ZN(n13339) );
  NAND2_X1 U16584 ( .A1(n10527), .A2(n13338), .ZN(n14972) );
  INV_X1 U16585 ( .A(n13339), .ZN(n14963) );
  AOI22_X1 U16586 ( .A1(n10632), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10633), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13345) );
  INV_X1 U16587 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13340) );
  OAI21_X1 U16588 ( .B1(n13242), .B2(n13340), .A(n13390), .ZN(n13341) );
  AOI21_X1 U16589 ( .B1(n10421), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n13341), .ZN(n13344) );
  AOI22_X1 U16590 ( .A1(n9816), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(n9834), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13343) );
  AOI22_X1 U16591 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n16444), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13342) );
  NAND4_X1 U16592 ( .A1(n13345), .A2(n13344), .A3(n13343), .A4(n13342), .ZN(
        n13353) );
  AOI22_X1 U16593 ( .A1(n10632), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10633), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13351) );
  AOI22_X1 U16594 ( .A1(n10634), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13350) );
  AOI22_X1 U16595 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n16444), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13349) );
  NAND2_X1 U16596 ( .A1(n9807), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n13347) );
  AOI21_X1 U16597 ( .B1(n13320), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n13390), .ZN(n13346) );
  AND2_X1 U16598 ( .A1(n13347), .A2(n13346), .ZN(n13348) );
  NAND4_X1 U16599 ( .A1(n13351), .A2(n13350), .A3(n13349), .A4(n13348), .ZN(
        n13352) );
  AND2_X1 U16600 ( .A1(n13353), .A2(n13352), .ZN(n14964) );
  INV_X1 U16601 ( .A(n14962), .ZN(n13355) );
  NAND2_X1 U16602 ( .A1(n19447), .A2(n14964), .ZN(n13354) );
  NOR2_X1 U16603 ( .A1(n13355), .A2(n13354), .ZN(n13374) );
  AOI22_X1 U16604 ( .A1(n9840), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10633), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13364) );
  INV_X1 U16605 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13356) );
  OAI21_X1 U16606 ( .B1(n13242), .B2(n13356), .A(n13390), .ZN(n13357) );
  AOI21_X1 U16607 ( .B1(n9807), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A(n13357), .ZN(n13363) );
  AOI22_X1 U16608 ( .A1(n9817), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13362) );
  INV_X1 U16609 ( .A(n16444), .ZN(n16440) );
  INV_X1 U16610 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13358) );
  OAI22_X1 U16611 ( .A1(n13381), .A2(n13359), .B1(n16440), .B2(n13358), .ZN(
        n13360) );
  INV_X1 U16612 ( .A(n13360), .ZN(n13361) );
  NAND4_X1 U16613 ( .A1(n13364), .A2(n13363), .A3(n13362), .A4(n13361), .ZN(
        n13372) );
  AOI22_X1 U16614 ( .A1(n10632), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10633), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13370) );
  AOI22_X1 U16615 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9834), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13369) );
  AOI22_X1 U16616 ( .A1(n9817), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n16444), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13368) );
  NAND2_X1 U16617 ( .A1(n9808), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n13366) );
  AOI21_X1 U16618 ( .B1(n13320), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n13390), .ZN(n13365) );
  AND2_X1 U16619 ( .A1(n13366), .A2(n13365), .ZN(n13367) );
  NAND4_X1 U16620 ( .A1(n13370), .A2(n13369), .A3(n13368), .A4(n13367), .ZN(
        n13371) );
  AND2_X1 U16621 ( .A1(n13372), .A2(n13371), .ZN(n13373) );
  NAND2_X1 U16622 ( .A1(n13374), .A2(n13373), .ZN(n13375) );
  OAI21_X1 U16623 ( .B1(n13374), .B2(n13373), .A(n13375), .ZN(n14954) );
  INV_X1 U16624 ( .A(n13375), .ZN(n13376) );
  NOR2_X1 U16625 ( .A1(n14953), .A2(n13376), .ZN(n13400) );
  INV_X1 U16626 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13377) );
  OAI21_X1 U16627 ( .B1(n13242), .B2(n13377), .A(n13390), .ZN(n13383) );
  INV_X1 U16628 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13380) );
  OAI22_X1 U16629 ( .A1(n9839), .A2(n13380), .B1(n13379), .B2(n13378), .ZN(
        n13382) );
  AOI211_X1 U16630 ( .C1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .C2(n9808), .A(
        n13383), .B(n13382), .ZN(n13386) );
  AOI22_X1 U16631 ( .A1(n9840), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13385) );
  AOI22_X1 U16632 ( .A1(n10634), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n16444), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13384) );
  NAND3_X1 U16633 ( .A1(n13386), .A2(n13385), .A3(n13384), .ZN(n13398) );
  INV_X1 U16634 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13387) );
  NOR2_X1 U16635 ( .A1(n13388), .A2(n13387), .ZN(n13389) );
  AOI211_X1 U16636 ( .C1(n9834), .C2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n13390), .B(n13389), .ZN(n13396) );
  AOI22_X1 U16637 ( .A1(n16444), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13320), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13395) );
  AOI22_X1 U16638 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9817), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13394) );
  AOI22_X1 U16639 ( .A1(n10632), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10633), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13393) );
  NAND4_X1 U16640 ( .A1(n13396), .A2(n13395), .A3(n13394), .A4(n13393), .ZN(
        n13397) );
  NAND2_X1 U16641 ( .A1(n13398), .A2(n13397), .ZN(n13399) );
  XNOR2_X1 U16642 ( .A(n13400), .B(n13399), .ZN(n14952) );
  AND2_X1 U16643 ( .A1(n14848), .A2(n14851), .ZN(n13440) );
  NAND2_X1 U16644 ( .A1(n13439), .A2(n13440), .ZN(n13401) );
  NOR2_X1 U16645 ( .A1(n13441), .A2(n13401), .ZN(n13402) );
  AOI21_X1 U16646 ( .B1(n15641), .B2(n16430), .A(n13402), .ZN(n13668) );
  NAND2_X1 U16647 ( .A1(n13668), .A2(n13403), .ZN(n13404) );
  NOR4_X1 U16648 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n13410) );
  NOR4_X1 U16649 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n13409) );
  NOR4_X1 U16650 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n13408) );
  NOR4_X1 U16651 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n13407) );
  NAND4_X1 U16652 ( .A1(n13410), .A2(n13409), .A3(n13408), .A4(n13407), .ZN(
        n13415) );
  NOR4_X1 U16653 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n13413) );
  NOR4_X1 U16654 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n13412) );
  NOR4_X1 U16655 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n13411) );
  NAND4_X1 U16656 ( .A1(n13413), .A2(n13412), .A3(n13411), .A4(n20059), .ZN(
        n13414) );
  OAI21_X4 U16657 ( .B1(n13415), .B2(n13414), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13520) );
  NAND2_X1 U16658 ( .A1(n13520), .A2(BUF2_REG_14__SCAN_IN), .ZN(n13417) );
  INV_X1 U16659 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n16554) );
  OR2_X1 U16660 ( .A1(n13520), .A2(n16554), .ZN(n13416) );
  NAND2_X1 U16661 ( .A1(n13417), .A2(n13416), .ZN(n19406) );
  INV_X1 U16662 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13424) );
  INV_X1 U16663 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15325) );
  INV_X1 U16664 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n20107) );
  OAI222_X1 U16665 ( .A1(n13420), .A2(n13424), .B1(n13419), .B2(n15325), .C1(
        n20107), .C2(n13418), .ZN(n13422) );
  OR2_X1 U16666 ( .A1(n13421), .A2(n13422), .ZN(n13423) );
  OAI22_X1 U16667 ( .A1(n19348), .A2(n15321), .B1(n19347), .B2(n13424), .ZN(
        n13425) );
  AOI21_X1 U16668 ( .B1(n19298), .B2(n19406), .A(n13425), .ZN(n13429) );
  NOR2_X1 U16669 ( .A1(n13426), .A2(n13076), .ZN(n13427) );
  AOI22_X1 U16670 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19299), .B1(n19300), .B2(
        BUF2_REG_30__SCAN_IN), .ZN(n13428) );
  AND2_X1 U16671 ( .A1(n13429), .A2(n13428), .ZN(n13430) );
  OAI21_X1 U16672 ( .B1(n14952), .B2(n19361), .A(n13430), .ZN(P2_U2889) );
  NOR2_X1 U16673 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13432) );
  NOR4_X1 U16674 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13431) );
  NAND4_X1 U16675 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13432), .A4(n13431), .ZN(n13435) );
  NOR3_X1 U16676 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(P1_D_C_N_REG_SCAN_IN), .A3(
        n21375), .ZN(n13434) );
  NOR4_X1 U16677 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(P1_BE_N_REG_2__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n13433)
         );
  NAND4_X1 U16678 ( .A1(n20373), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13434), .A4(
        n13433), .ZN(U214) );
  NOR2_X1 U16679 ( .A1(n13520), .A2(n13435), .ZN(n16536) );
  NAND2_X1 U16680 ( .A1(n16536), .A2(U214), .ZN(U212) );
  NOR2_X1 U16681 ( .A1(n13444), .A2(n13674), .ZN(n19232) );
  INV_X1 U16682 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n20177) );
  INV_X1 U16683 ( .A(n13444), .ZN(n13438) );
  INV_X1 U16684 ( .A(n13436), .ZN(n13437) );
  NAND2_X1 U16685 ( .A1(n20126), .A2(n16479), .ZN(n13445) );
  OAI211_X1 U16686 ( .C1(n19232), .C2(n20177), .A(n14150), .B(n13445), .ZN(
        P2_U2814) );
  NOR4_X1 U16687 ( .A1(n13441), .A2(n13440), .A3(n16426), .A4(n13663), .ZN(
        n16466) );
  NOR2_X1 U16688 ( .A1(n16466), .A2(n16488), .ZN(n20173) );
  NOR2_X1 U16689 ( .A1(n11015), .A2(n16488), .ZN(n13442) );
  NAND2_X1 U16690 ( .A1(n13535), .A2(n19437), .ZN(n13533) );
  OAI21_X1 U16691 ( .B1(n20173), .B2(n11000), .A(n13533), .ZN(P2_U2819) );
  NOR2_X1 U16692 ( .A1(n19014), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n13446)
         );
  AOI22_X1 U16693 ( .A1(n19014), .A2(n13447), .B1(n13446), .B2(n13445), .ZN(
        P2_U3612) );
  INV_X1 U16694 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13451) );
  INV_X1 U16695 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13450) );
  INV_X1 U16696 ( .A(n14150), .ZN(n13448) );
  OAI21_X1 U16697 ( .B1(n10527), .B2(n14851), .A(n13448), .ZN(n13459) );
  INV_X1 U16698 ( .A(n13459), .ZN(n13504) );
  NAND2_X1 U16699 ( .A1(n19447), .A2(n14851), .ZN(n13449) );
  AOI22_X1 U16700 ( .A1(n19436), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n13520), .ZN(n19308) );
  OAI222_X1 U16701 ( .A1(n14152), .A2(n13451), .B1(n13450), .B2(n13504), .C1(
        n13469), .C2(n19308), .ZN(P2_U2982) );
  INV_X2 U16702 ( .A(n14152), .ZN(n19409) );
  AOI22_X1 U16703 ( .A1(P2_LWORD_REG_6__SCAN_IN), .A2(n13459), .B1(n19409), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n13452) );
  OAI22_X1 U16704 ( .A1(n13520), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n19436), .ZN(n19476) );
  INV_X1 U16705 ( .A(n19476), .ZN(n16278) );
  NAND2_X1 U16706 ( .A1(n19407), .A2(n16278), .ZN(n13472) );
  NAND2_X1 U16707 ( .A1(n13452), .A2(n13472), .ZN(P2_U2973) );
  AOI22_X1 U16708 ( .A1(P2_LWORD_REG_5__SCAN_IN), .A2(n13459), .B1(n19409), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n13454) );
  AOI22_X1 U16709 ( .A1(n19436), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n13520), .ZN(n19471) );
  INV_X1 U16710 ( .A(n19471), .ZN(n13453) );
  NAND2_X1 U16711 ( .A1(n19407), .A2(n13453), .ZN(n13474) );
  NAND2_X1 U16712 ( .A1(n13454), .A2(n13474), .ZN(P2_U2972) );
  AOI22_X1 U16713 ( .A1(P2_LWORD_REG_7__SCAN_IN), .A2(n13459), .B1(n19409), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n13455) );
  AOI22_X1 U16714 ( .A1(n19436), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n13520), .ZN(n19488) );
  INV_X1 U16715 ( .A(n19488), .ZN(n15077) );
  NAND2_X1 U16716 ( .A1(n19407), .A2(n15077), .ZN(n13507) );
  NAND2_X1 U16717 ( .A1(n13455), .A2(n13507), .ZN(P2_U2974) );
  AOI22_X1 U16718 ( .A1(P2_LWORD_REG_9__SCAN_IN), .A2(n13459), .B1(n19409), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n13458) );
  INV_X1 U16719 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16564) );
  OR2_X1 U16720 ( .A1(n13520), .A2(n16564), .ZN(n13457) );
  NAND2_X1 U16721 ( .A1(n13520), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13456) );
  AND2_X1 U16722 ( .A1(n13457), .A2(n13456), .ZN(n19322) );
  INV_X1 U16723 ( .A(n19322), .ZN(n15057) );
  NAND2_X1 U16724 ( .A1(n19407), .A2(n15057), .ZN(n13505) );
  NAND2_X1 U16725 ( .A1(n13458), .A2(n13505), .ZN(P2_U2976) );
  AOI22_X1 U16726 ( .A1(P2_LWORD_REG_11__SCAN_IN), .A2(n13459), .B1(n19409), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n13462) );
  INV_X1 U16727 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n16560) );
  OR2_X1 U16728 ( .A1(n13520), .A2(n16560), .ZN(n13461) );
  NAND2_X1 U16729 ( .A1(n13520), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13460) );
  AND2_X1 U16730 ( .A1(n13461), .A2(n13460), .ZN(n19317) );
  INV_X1 U16731 ( .A(n19317), .ZN(n15041) );
  NAND2_X1 U16732 ( .A1(n19407), .A2(n15041), .ZN(n13516) );
  NAND2_X1 U16733 ( .A1(n13462), .A2(n13516), .ZN(P2_U2978) );
  INV_X1 U16734 ( .A(n13463), .ZN(n13465) );
  INV_X1 U16735 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n21392) );
  NOR2_X1 U16736 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20926), .ZN(n14400) );
  INV_X1 U16737 ( .A(n14400), .ZN(n13464) );
  OAI211_X1 U16738 ( .C1(n13465), .C2(n21392), .A(n13701), .B(n13464), .ZN(
        P1_U2801) );
  AOI22_X1 U16739 ( .A1(P2_UWORD_REG_2__SCAN_IN), .A2(n13459), .B1(n19409), 
        .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n13466) );
  INV_X1 U16740 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16578) );
  INV_X1 U16741 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18342) );
  AOI22_X1 U16742 ( .A1(n19436), .A2(n16578), .B1(n18342), .B2(n13520), .ZN(
        n16291) );
  INV_X1 U16743 ( .A(n16291), .ZN(n19453) );
  OR2_X1 U16744 ( .A1(n13469), .A2(n19453), .ZN(n13528) );
  NAND2_X1 U16745 ( .A1(n13466), .A2(n13528), .ZN(P2_U2954) );
  AOI22_X1 U16746 ( .A1(P2_UWORD_REG_1__SCAN_IN), .A2(n13459), .B1(n19409), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n13468) );
  AOI22_X1 U16747 ( .A1(n19436), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13520), .ZN(n19448) );
  INV_X1 U16748 ( .A(n19448), .ZN(n13467) );
  NAND2_X1 U16749 ( .A1(n19407), .A2(n13467), .ZN(n13511) );
  NAND2_X1 U16750 ( .A1(n13468), .A2(n13511), .ZN(P2_U2953) );
  AOI22_X1 U16751 ( .A1(P2_UWORD_REG_0__SCAN_IN), .A2(n13459), .B1(n19409), 
        .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n13470) );
  INV_X1 U16752 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16585) );
  INV_X1 U16753 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18329) );
  AOI22_X1 U16754 ( .A1(n19436), .A2(n16585), .B1(n18329), .B2(n13520), .ZN(
        n19297) );
  INV_X1 U16755 ( .A(n19297), .ZN(n19438) );
  OR2_X1 U16756 ( .A1(n13469), .A2(n19438), .ZN(n13530) );
  NAND2_X1 U16757 ( .A1(n13470), .A2(n13530), .ZN(P2_U2952) );
  AOI22_X1 U16758 ( .A1(P2_UWORD_REG_3__SCAN_IN), .A2(n13459), .B1(n19409), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n13471) );
  AOI22_X1 U16759 ( .A1(n19436), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13520), .ZN(n19459) );
  INV_X1 U16760 ( .A(n19459), .ZN(n15093) );
  NAND2_X1 U16761 ( .A1(n19407), .A2(n15093), .ZN(n13518) );
  NAND2_X1 U16762 ( .A1(n13471), .A2(n13518), .ZN(P2_U2955) );
  AOI22_X1 U16763 ( .A1(P2_UWORD_REG_6__SCAN_IN), .A2(n13459), .B1(n19409), 
        .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n13473) );
  NAND2_X1 U16764 ( .A1(n13473), .A2(n13472), .ZN(P2_U2958) );
  AOI22_X1 U16765 ( .A1(P2_UWORD_REG_5__SCAN_IN), .A2(n19405), .B1(n19409), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n13475) );
  NAND2_X1 U16766 ( .A1(n13475), .A2(n13474), .ZN(P2_U2957) );
  AOI22_X1 U16767 ( .A1(P2_UWORD_REG_4__SCAN_IN), .A2(n19405), .B1(n19409), 
        .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n13476) );
  OAI22_X1 U16768 ( .A1(n13520), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n19436), .ZN(n19465) );
  INV_X1 U16769 ( .A(n19465), .ZN(n16285) );
  NAND2_X1 U16770 ( .A1(n19407), .A2(n16285), .ZN(n13509) );
  NAND2_X1 U16771 ( .A1(n13476), .A2(n13509), .ZN(P2_U2956) );
  INV_X1 U16772 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13567) );
  NAND2_X1 U16773 ( .A1(n13520), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13478) );
  INV_X1 U16774 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16562) );
  OR2_X1 U16775 ( .A1(n13520), .A2(n16562), .ZN(n13477) );
  NAND2_X1 U16776 ( .A1(n13478), .A2(n13477), .ZN(n19319) );
  NAND2_X1 U16777 ( .A1(n19407), .A2(n19319), .ZN(n13497) );
  NAND2_X1 U16778 ( .A1(n19405), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13479) );
  OAI211_X1 U16779 ( .C1(n13567), .C2(n14152), .A(n13497), .B(n13479), .ZN(
        P2_U2962) );
  INV_X1 U16780 ( .A(n13480), .ZN(n13492) );
  AND2_X1 U16781 ( .A1(n12882), .A2(n13492), .ZN(n13481) );
  OR2_X1 U16782 ( .A1(n13481), .A2(n12881), .ZN(n13484) );
  NAND2_X1 U16783 ( .A1(n13751), .A2(n13482), .ZN(n13483) );
  NAND2_X1 U16784 ( .A1(n13484), .A2(n13483), .ZN(n20181) );
  INV_X1 U16785 ( .A(n21073), .ZN(n21070) );
  OR2_X1 U16786 ( .A1(n13485), .A2(n21070), .ZN(n13486) );
  AND2_X1 U16787 ( .A1(n13486), .A2(n21064), .ZN(n13605) );
  INV_X1 U16788 ( .A(n13605), .ZN(n13488) );
  NAND2_X1 U16789 ( .A1(n14026), .A2(n21064), .ZN(n13487) );
  NAND2_X1 U16790 ( .A1(n13488), .A2(n13487), .ZN(n13489) );
  NOR2_X1 U16791 ( .A1(n20181), .A2(n13489), .ZN(n15815) );
  OR2_X1 U16792 ( .A1(n15815), .A2(n20180), .ZN(n20186) );
  INV_X1 U16793 ( .A(n12881), .ZN(n13490) );
  NAND3_X1 U16794 ( .A1(n13490), .A2(n13912), .A3(n15816), .ZN(n13494) );
  INV_X1 U16795 ( .A(n12882), .ZN(n13615) );
  INV_X1 U16796 ( .A(n13914), .ZN(n13491) );
  OAI22_X1 U16797 ( .A1(n13615), .A2(n13492), .B1(n13751), .B2(n13491), .ZN(
        n13493) );
  AOI21_X1 U16798 ( .B1(n13494), .B2(n13751), .A(n13493), .ZN(n15817) );
  NAND2_X1 U16799 ( .A1(n20186), .A2(P1_MORE_REG_SCAN_IN), .ZN(n13495) );
  OAI21_X1 U16800 ( .B1(n20186), .B2(n15817), .A(n13495), .ZN(P1_U3484) );
  NAND2_X1 U16801 ( .A1(n19405), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13496) );
  OAI211_X1 U16802 ( .C1(n11298), .C2(n14152), .A(n13497), .B(n13496), .ZN(
        P2_U2977) );
  INV_X1 U16803 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19386) );
  MUX2_X1 U16804 ( .A(BUF1_REG_8__SCAN_IN), .B(BUF2_REG_8__SCAN_IN), .S(n13520), .Z(n19326) );
  NAND2_X1 U16805 ( .A1(n19407), .A2(n19326), .ZN(n13500) );
  NAND2_X1 U16806 ( .A1(n19405), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13498) );
  OAI211_X1 U16807 ( .C1(n19386), .C2(n14152), .A(n13500), .B(n13498), .ZN(
        P2_U2975) );
  INV_X1 U16808 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13581) );
  NAND2_X1 U16809 ( .A1(n19405), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13499) );
  OAI211_X1 U16810 ( .C1(n13581), .C2(n14152), .A(n13500), .B(n13499), .ZN(
        P2_U2960) );
  INV_X1 U16811 ( .A(n13501), .ZN(n21067) );
  OAI21_X1 U16812 ( .B1(n14400), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n21067), 
        .ZN(n13502) );
  OAI21_X1 U16813 ( .B1(n13503), .B2(n21067), .A(n13502), .ZN(P1_U3487) );
  AOI22_X1 U16814 ( .A1(P2_UWORD_REG_9__SCAN_IN), .A2(n19405), .B1(n19409), 
        .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n13506) );
  NAND2_X1 U16815 ( .A1(n13506), .A2(n13505), .ZN(P2_U2961) );
  AOI22_X1 U16816 ( .A1(P2_UWORD_REG_7__SCAN_IN), .A2(n19405), .B1(n19409), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n13508) );
  NAND2_X1 U16817 ( .A1(n13508), .A2(n13507), .ZN(P2_U2959) );
  AOI22_X1 U16818 ( .A1(P2_LWORD_REG_4__SCAN_IN), .A2(n19405), .B1(n19409), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n13510) );
  NAND2_X1 U16819 ( .A1(n13510), .A2(n13509), .ZN(P2_U2971) );
  AOI22_X1 U16820 ( .A1(P2_LWORD_REG_1__SCAN_IN), .A2(n19405), .B1(n19409), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n13512) );
  NAND2_X1 U16821 ( .A1(n13512), .A2(n13511), .ZN(P2_U2968) );
  AOI22_X1 U16822 ( .A1(P2_LWORD_REG_12__SCAN_IN), .A2(n19405), .B1(n19409), 
        .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n13515) );
  INV_X1 U16823 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16558) );
  OR2_X1 U16824 ( .A1(n13520), .A2(n16558), .ZN(n13514) );
  NAND2_X1 U16825 ( .A1(n13520), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13513) );
  AND2_X1 U16826 ( .A1(n13514), .A2(n13513), .ZN(n19315) );
  INV_X1 U16827 ( .A(n19315), .ZN(n15031) );
  NAND2_X1 U16828 ( .A1(n19407), .A2(n15031), .ZN(n13526) );
  NAND2_X1 U16829 ( .A1(n13515), .A2(n13526), .ZN(P2_U2979) );
  AOI22_X1 U16830 ( .A1(P2_UWORD_REG_11__SCAN_IN), .A2(n19405), .B1(n19409), 
        .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n13517) );
  NAND2_X1 U16831 ( .A1(n13517), .A2(n13516), .ZN(P2_U2963) );
  AOI22_X1 U16832 ( .A1(P2_LWORD_REG_3__SCAN_IN), .A2(n19405), .B1(n19409), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n13519) );
  NAND2_X1 U16833 ( .A1(n13519), .A2(n13518), .ZN(P2_U2970) );
  AOI22_X1 U16834 ( .A1(P2_LWORD_REG_13__SCAN_IN), .A2(n19405), .B1(n19409), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n13523) );
  INV_X1 U16835 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16556) );
  OR2_X1 U16836 ( .A1(n13520), .A2(n16556), .ZN(n13522) );
  NAND2_X1 U16837 ( .A1(n13520), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13521) );
  AND2_X1 U16838 ( .A1(n13522), .A2(n13521), .ZN(n19312) );
  INV_X1 U16839 ( .A(n19312), .ZN(n15023) );
  NAND2_X1 U16840 ( .A1(n19407), .A2(n15023), .ZN(n13524) );
  NAND2_X1 U16841 ( .A1(n13523), .A2(n13524), .ZN(P2_U2980) );
  AOI22_X1 U16842 ( .A1(P2_UWORD_REG_13__SCAN_IN), .A2(n19405), .B1(n19409), 
        .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n13525) );
  NAND2_X1 U16843 ( .A1(n13525), .A2(n13524), .ZN(P2_U2965) );
  AOI22_X1 U16844 ( .A1(P2_UWORD_REG_12__SCAN_IN), .A2(n19405), .B1(n19409), 
        .B2(P2_EAX_REG_28__SCAN_IN), .ZN(n13527) );
  NAND2_X1 U16845 ( .A1(n13527), .A2(n13526), .ZN(P2_U2964) );
  AOI22_X1 U16846 ( .A1(P2_LWORD_REG_2__SCAN_IN), .A2(n19405), .B1(n19409), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n13529) );
  NAND2_X1 U16847 ( .A1(n13529), .A2(n13528), .ZN(P2_U2969) );
  AOI22_X1 U16848 ( .A1(P2_LWORD_REG_0__SCAN_IN), .A2(n19405), .B1(n19409), 
        .B2(P2_EAX_REG_0__SCAN_IN), .ZN(n13531) );
  NAND2_X1 U16849 ( .A1(n13531), .A2(n13530), .ZN(P2_U2967) );
  NOR2_X1 U16850 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20029) );
  OR2_X1 U16851 ( .A1(n20126), .A2(n20029), .ZN(n20156) );
  NAND2_X1 U16852 ( .A1(n20156), .A2(n16491), .ZN(n13532) );
  AND2_X1 U16853 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20148) );
  AOI21_X1 U16854 ( .B1(n11221), .B2(n16421), .A(n13534), .ZN(n16414) );
  INV_X1 U16855 ( .A(n13535), .ZN(n13536) );
  OAI21_X1 U16856 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n19240), .A(
        n13546), .ZN(n16424) );
  NAND2_X1 U16857 ( .A1(n19414), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n16422) );
  OAI21_X1 U16858 ( .B1(n19417), .B2(n16424), .A(n16422), .ZN(n13542) );
  INV_X1 U16859 ( .A(n13537), .ZN(n13539) );
  INV_X1 U16860 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19612) );
  NAND2_X1 U16861 ( .A1(n19612), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13538) );
  NAND2_X1 U16862 ( .A1(n13539), .A2(n13538), .ZN(n13544) );
  OAI21_X1 U16863 ( .B1(n16316), .B2(n13544), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13540) );
  INV_X1 U16864 ( .A(n13540), .ZN(n13541) );
  AOI211_X1 U16865 ( .C1(n16414), .C2(n19421), .A(n13542), .B(n13541), .ZN(
        n13543) );
  OAI21_X1 U16866 ( .B1(n19245), .B2(n19416), .A(n13543), .ZN(P2_U3014) );
  OAI22_X1 U16867 ( .A1(n13592), .A2(n19416), .B1(n16355), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13554) );
  OAI21_X1 U16868 ( .B1(n13546), .B2(n19221), .A(n13545), .ZN(n13547) );
  XNOR2_X1 U16869 ( .A(n13547), .B(n15649), .ZN(n13716) );
  OAI21_X1 U16870 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13549), .A(
        n13548), .ZN(n13550) );
  INV_X1 U16871 ( .A(n13550), .ZN(n13715) );
  AND2_X1 U16872 ( .A1(n19414), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n13719) );
  AOI21_X1 U16873 ( .B1(n19421), .B2(n13715), .A(n13719), .ZN(n13552) );
  OR2_X1 U16874 ( .A1(n19425), .A2(n19233), .ZN(n13551) );
  OAI211_X1 U16875 ( .C1(n13716), .C2(n19417), .A(n13552), .B(n13551), .ZN(
        n13553) );
  OR2_X1 U16876 ( .A1(n13554), .A2(n13553), .ZN(P2_U3013) );
  NAND2_X1 U16877 ( .A1(n19447), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13555) );
  NAND4_X1 U16878 ( .A1(n13555), .A2(n13076), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n20136), .ZN(n13556) );
  INV_X1 U16879 ( .A(n15641), .ZN(n16431) );
  NAND2_X1 U16880 ( .A1(n16431), .A2(n15658), .ZN(n13666) );
  NAND2_X1 U16881 ( .A1(n13666), .A2(n10100), .ZN(n13557) );
  MUX2_X1 U16882 ( .A(n13558), .B(n19245), .S(n19293), .Z(n13559) );
  OAI21_X1 U16883 ( .B1(n20160), .B2(n19289), .A(n13559), .ZN(P2_U2887) );
  INV_X1 U16884 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13564) );
  NOR2_X1 U16885 ( .A1(n13674), .A2(n16488), .ZN(n13560) );
  NAND2_X1 U16886 ( .A1(n13665), .A2(n13560), .ZN(n13561) );
  NAND2_X1 U16887 ( .A1(n13561), .A2(n14152), .ZN(n13562) );
  NAND2_X1 U16888 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n15866) );
  NOR2_X1 U16889 ( .A1(n15866), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19397) );
  CLKBUF_X1 U16890 ( .A(n19397), .Z(n19402) );
  INV_X2 U16891 ( .A(n19370), .ZN(n19396) );
  AOI22_X1 U16892 ( .A1(n19402), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19396), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13563) );
  OAI21_X1 U16893 ( .B1(n13564), .B2(n19367), .A(n13563), .ZN(P2_U2935) );
  INV_X1 U16894 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n15102) );
  AOI22_X1 U16895 ( .A1(n19402), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19396), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13565) );
  OAI21_X1 U16896 ( .B1(n15102), .B2(n19367), .A(n13565), .ZN(P2_U2934) );
  AOI22_X1 U16897 ( .A1(n19402), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19396), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13566) );
  OAI21_X1 U16898 ( .B1(n13567), .B2(n19367), .A(n13566), .ZN(P2_U2925) );
  INV_X1 U16899 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n13569) );
  AOI22_X1 U16900 ( .A1(n19402), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19396), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13568) );
  OAI21_X1 U16901 ( .B1(n13569), .B2(n19367), .A(n13568), .ZN(P2_U2926) );
  INV_X1 U16902 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n13571) );
  AOI22_X1 U16903 ( .A1(n19402), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19396), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13570) );
  OAI21_X1 U16904 ( .B1(n13571), .B2(n19367), .A(n13570), .ZN(P2_U2922) );
  INV_X1 U16905 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n13573) );
  AOI22_X1 U16906 ( .A1(n19402), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19396), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13572) );
  OAI21_X1 U16907 ( .B1(n13573), .B2(n19367), .A(n13572), .ZN(P2_U2932) );
  AOI22_X1 U16908 ( .A1(n19402), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19396), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13574) );
  OAI21_X1 U16909 ( .B1(n13575), .B2(n19367), .A(n13574), .ZN(P2_U2928) );
  INV_X1 U16910 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13577) );
  AOI22_X1 U16911 ( .A1(n19402), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19396), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13576) );
  OAI21_X1 U16912 ( .B1(n13577), .B2(n19367), .A(n13576), .ZN(P2_U2923) );
  INV_X1 U16913 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13579) );
  AOI22_X1 U16914 ( .A1(n19402), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19396), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13578) );
  OAI21_X1 U16915 ( .B1(n13579), .B2(n19367), .A(n13578), .ZN(P2_U2929) );
  AOI22_X1 U16916 ( .A1(n19402), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19396), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13580) );
  OAI21_X1 U16917 ( .B1(n13581), .B2(n19367), .A(n13580), .ZN(P2_U2927) );
  INV_X1 U16918 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13583) );
  AOI22_X1 U16919 ( .A1(n19402), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19396), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13582) );
  OAI21_X1 U16920 ( .B1(n13583), .B2(n19367), .A(n13582), .ZN(P2_U2933) );
  AOI22_X1 U16921 ( .A1(n19402), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19396), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13584) );
  OAI21_X1 U16922 ( .B1(n15082), .B2(n19367), .A(n13584), .ZN(P2_U2930) );
  INV_X1 U16923 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13586) );
  AOI22_X1 U16924 ( .A1(n19402), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19396), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13585) );
  OAI21_X1 U16925 ( .B1(n13586), .B2(n19367), .A(n13585), .ZN(P2_U2931) );
  INV_X1 U16926 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n13588) );
  AOI22_X1 U16927 ( .A1(n19402), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19396), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13587) );
  OAI21_X1 U16928 ( .B1(n13588), .B2(n19367), .A(n13587), .ZN(P2_U2924) );
  INV_X1 U16929 ( .A(n13590), .ZN(n13591) );
  MUX2_X1 U16930 ( .A(n13593), .B(n13592), .S(n19293), .Z(n13594) );
  OAI21_X1 U16931 ( .B1(n20130), .B2(n19289), .A(n13594), .ZN(P2_U2886) );
  AOI21_X1 U16932 ( .B1(n19233), .B2(n14936), .A(n14078), .ZN(n14934) );
  NAND2_X1 U16933 ( .A1(n13596), .A2(n13595), .ZN(n13734) );
  NAND3_X1 U16934 ( .A1(n13735), .A2(n16366), .A3(n13734), .ZN(n13597) );
  OAI21_X1 U16935 ( .B1(n19425), .B2(n14936), .A(n13597), .ZN(n13602) );
  OAI21_X1 U16936 ( .B1(n13600), .B2(n13599), .A(n13598), .ZN(n13722) );
  OAI22_X1 U16937 ( .A1(n10580), .A2(n19176), .B1(n16371), .B2(n13722), .ZN(
        n13601) );
  AOI211_X1 U16938 ( .C1(n19413), .C2(n14934), .A(n13602), .B(n13601), .ZN(
        n13603) );
  OAI21_X1 U16939 ( .B1(n10596), .B2(n19416), .A(n13603), .ZN(P2_U3012) );
  NAND2_X1 U16940 ( .A1(n15803), .A2(n21070), .ZN(n13646) );
  INV_X1 U16941 ( .A(n13604), .ZN(n13639) );
  NAND2_X1 U16942 ( .A1(n13646), .A2(n13639), .ZN(n13606) );
  NAND2_X1 U16943 ( .A1(n13606), .A2(n13605), .ZN(n13607) );
  NAND2_X1 U16944 ( .A1(n13607), .A2(n13912), .ZN(n13609) );
  INV_X1 U16945 ( .A(n13751), .ZN(n13608) );
  NAND2_X1 U16946 ( .A1(n13609), .A2(n13608), .ZN(n13620) );
  AOI21_X1 U16947 ( .B1(n13610), .B2(n12074), .A(n11918), .ZN(n13611) );
  NAND2_X1 U16948 ( .A1(n13612), .A2(n13611), .ZN(n13634) );
  NAND2_X1 U16949 ( .A1(n13613), .A2(n13634), .ZN(n13614) );
  NAND2_X1 U16950 ( .A1(n13615), .A2(n13614), .ZN(n13756) );
  INV_X1 U16951 ( .A(n13763), .ZN(n20405) );
  OR2_X1 U16952 ( .A1(n14028), .A2(n20405), .ZN(n13616) );
  AND4_X1 U16953 ( .A1(n13618), .A2(n13756), .A3(n13617), .A4(n13616), .ZN(
        n13619) );
  INV_X1 U16954 ( .A(n15805), .ZN(n13621) );
  NAND2_X1 U16955 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n13648) );
  NAND2_X1 U16956 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20989), .ZN(n16151) );
  INV_X1 U16957 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n21319) );
  OAI22_X1 U16958 ( .A1(n13621), .A2(n20180), .B1(n16151), .B2(n21319), .ZN(
        n13624) );
  AOI21_X1 U16959 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21075), .A(n13624), 
        .ZN(n14843) );
  INV_X1 U16960 ( .A(n14843), .ZN(n14831) );
  INV_X1 U16961 ( .A(n20537), .ZN(n20788) );
  OR2_X1 U16962 ( .A1(n13622), .A2(n20788), .ZN(n13623) );
  XNOR2_X1 U16963 ( .A(n13623), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20271) );
  INV_X1 U16964 ( .A(n13043), .ZN(n13942) );
  NAND4_X1 U16965 ( .A1(n20271), .A2(n14825), .A3(n13942), .A4(n13624), .ZN(
        n13625) );
  OAI21_X1 U16966 ( .B1(n14831), .B2(n13626), .A(n13625), .ZN(P1_U3468) );
  AOI21_X1 U16967 ( .B1(n15803), .B2(n14825), .A(n14843), .ZN(n13645) );
  INV_X1 U16968 ( .A(n12075), .ZN(n13968) );
  OAI211_X1 U16969 ( .C1(n11928), .C2(n13763), .A(n20443), .B(n13923), .ZN(
        n13629) );
  NAND2_X1 U16970 ( .A1(n13629), .A2(n11917), .ZN(n13632) );
  OR2_X1 U16971 ( .A1(n13630), .A2(n14028), .ZN(n13631) );
  AND4_X1 U16972 ( .A1(n13634), .A2(n13633), .A3(n13632), .A4(n13631), .ZN(
        n13636) );
  AND3_X1 U16973 ( .A1(n13637), .A2(n13636), .A3(n13635), .ZN(n13778) );
  AND2_X1 U16974 ( .A1(n13638), .A2(n13779), .ZN(n13640) );
  NAND4_X1 U16975 ( .A1(n13043), .A2(n13778), .A3(n13640), .A4(n13639), .ZN(
        n14824) );
  INV_X1 U16976 ( .A(n14824), .ZN(n13641) );
  OAI22_X1 U16977 ( .A1(n13968), .A2(n13641), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n11888), .ZN(n15802) );
  OAI22_X1 U16978 ( .A1(n16145), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15835), .ZN(n13642) );
  AOI21_X1 U16979 ( .B1(n15802), .B2(n14825), .A(n13642), .ZN(n13643) );
  OAI22_X1 U16980 ( .A1(n13645), .A2(n13644), .B1(n13643), .B2(n14843), .ZN(
        P1_U3474) );
  INV_X1 U16981 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n21206) );
  NAND2_X1 U16982 ( .A1(n12881), .A2(n13753), .ZN(n13774) );
  OR2_X1 U16983 ( .A1(n13774), .A2(n21073), .ZN(n15826) );
  NAND2_X1 U16984 ( .A1(n15826), .A2(n13646), .ZN(n13647) );
  NOR2_X1 U16985 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n13648), .ZN(n20336) );
  INV_X1 U16986 ( .A(n20336), .ZN(n20308) );
  NOR2_X4 U16987 ( .A1(n20310), .A2(n20319), .ZN(n15849) );
  AOI22_X1 U16988 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20319), .B1(n15849), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13649) );
  OAI21_X1 U16989 ( .B1(n21206), .B2(n13816), .A(n13649), .ZN(P1_U2908) );
  INV_X1 U16990 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13651) );
  AOI22_X1 U16991 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20336), .B1(n15849), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13650) );
  OAI21_X1 U16992 ( .B1(n13651), .B2(n13816), .A(n13650), .ZN(P1_U2917) );
  INV_X1 U16993 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13653) );
  AOI22_X1 U16994 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20319), .B1(n15849), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13652) );
  OAI21_X1 U16995 ( .B1(n13653), .B2(n13816), .A(n13652), .ZN(P1_U2916) );
  INV_X1 U16996 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13706) );
  AOI22_X1 U16997 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20319), .B1(n15849), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13654) );
  OAI21_X1 U16998 ( .B1(n13706), .B2(n13816), .A(n13654), .ZN(P1_U2912) );
  INV_X1 U16999 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13656) );
  AOI22_X1 U17000 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20319), .B1(n15849), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13655) );
  OAI21_X1 U17001 ( .B1(n13656), .B2(n13816), .A(n13655), .ZN(P1_U2915) );
  INV_X1 U17002 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n21326) );
  AOI22_X1 U17003 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20319), .B1(n15849), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13657) );
  OAI21_X1 U17004 ( .B1(n21326), .B2(n13816), .A(n13657), .ZN(P1_U2914) );
  AOI22_X1 U17005 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20319), .B1(n15849), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13658) );
  OAI21_X1 U17006 ( .B1(n12532), .B2(n13816), .A(n13658), .ZN(P1_U2913) );
  AOI22_X1 U17007 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20319), .B1(n15849), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13659) );
  OAI21_X1 U17008 ( .B1(n13660), .B2(n13816), .A(n13659), .ZN(P1_U2918) );
  INV_X1 U17009 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13712) );
  AOI22_X1 U17010 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20319), .B1(n15849), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13661) );
  OAI21_X1 U17011 ( .B1(n13712), .B2(n13816), .A(n13661), .ZN(P1_U2911) );
  INV_X1 U17012 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n21350) );
  AOI22_X1 U17013 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20319), .B1(n15849), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13662) );
  OAI21_X1 U17014 ( .B1(n21350), .B2(n13816), .A(n13662), .ZN(P1_U2909) );
  NOR2_X1 U17015 ( .A1(n16491), .A2(n15866), .ZN(n16490) );
  INV_X1 U17016 ( .A(n13663), .ZN(n14148) );
  NOR2_X1 U17017 ( .A1(n13674), .A2(n14148), .ZN(n13664) );
  NAND2_X1 U17018 ( .A1(n13665), .A2(n13664), .ZN(n13669) );
  OAI22_X1 U17019 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20136), .B1(n16474), 
        .B2(n16488), .ZN(n13670) );
  INV_X1 U17020 ( .A(n20123), .ZN(n13677) );
  INV_X1 U17021 ( .A(n13671), .ZN(n13672) );
  NAND2_X1 U17022 ( .A1(n10527), .A2(n13672), .ZN(n13673) );
  NOR2_X1 U17023 ( .A1(n13674), .A2(n13673), .ZN(n16465) );
  NAND3_X1 U17024 ( .A1(n13677), .A2(n16465), .A3(n20029), .ZN(n13675) );
  OAI21_X1 U17025 ( .B1(n13677), .B2(n13676), .A(n13675), .ZN(P2_U3595) );
  NOR2_X1 U17026 ( .A1(n13680), .A2(n13679), .ZN(n13681) );
  OR2_X1 U17027 ( .A1(n11235), .A2(n13681), .ZN(n19237) );
  OAI22_X1 U17028 ( .A1(n19348), .A2(n19237), .B1(n19347), .B2(n13682), .ZN(
        n13684) );
  NOR2_X1 U17029 ( .A1(n20160), .A2(n19237), .ZN(n19360) );
  AOI211_X1 U17030 ( .C1(n20160), .C2(n19237), .A(n19361), .B(n19360), .ZN(
        n13683) );
  AOI211_X1 U17031 ( .C1(n19297), .C2(n19325), .A(n13684), .B(n13683), .ZN(
        n13685) );
  INV_X1 U17032 ( .A(n13685), .ZN(P2_U2919) );
  NOR2_X1 U17033 ( .A1(n13686), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13688) );
  OR2_X1 U17034 ( .A1(n13688), .A2(n13687), .ZN(n20354) );
  OAI21_X1 U17035 ( .B1(n13691), .B2(n13690), .A(n13689), .ZN(n14038) );
  OAI222_X1 U17036 ( .A1(n20354), .A2(n15973), .B1(n12903), .B2(n20306), .C1(
        n14038), .C2(n15974), .ZN(P1_U2872) );
  OR2_X1 U17037 ( .A1(n13692), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13693) );
  AND2_X1 U17038 ( .A1(n13694), .A2(n13693), .ZN(n20358) );
  INV_X1 U17039 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13697) );
  OAI21_X1 U17040 ( .B1(n16027), .B2(n13695), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13696) );
  OAI21_X1 U17041 ( .B1(n13697), .B2(n20369), .A(n13696), .ZN(n13698) );
  AOI21_X1 U17042 ( .B1(n20358), .B2(n16034), .A(n13698), .ZN(n13699) );
  OAI21_X1 U17043 ( .B1(n14689), .B2(n14038), .A(n13699), .ZN(P1_U2999) );
  INV_X1 U17044 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n21316) );
  OR2_X2 U17045 ( .A1(n13701), .A2(n13700), .ZN(n20348) );
  MUX2_X1 U17046 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n20373), .Z(
        n14467) );
  NAND2_X1 U17047 ( .A1(n13845), .A2(n14467), .ZN(n20342) );
  NAND2_X1 U17048 ( .A1(n20348), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n13702) );
  OAI211_X1 U17049 ( .C1(n21316), .C2(n13824), .A(n20342), .B(n13702), .ZN(
        P1_U2947) );
  INV_X1 U17050 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n21179) );
  MUX2_X1 U17051 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n20373), .Z(
        n14516) );
  NAND2_X1 U17052 ( .A1(n13845), .A2(n14516), .ZN(n20352) );
  NAND2_X1 U17053 ( .A1(n20348), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n13703) );
  OAI211_X1 U17054 ( .C1(n21179), .C2(n13824), .A(n20352), .B(n13703), .ZN(
        P1_U2951) );
  MUX2_X1 U17055 ( .A(DATAI_11_), .B(BUF1_REG_11__SCAN_IN), .S(n20373), .Z(
        n14533) );
  NAND2_X1 U17056 ( .A1(n13845), .A2(n14533), .ZN(n20344) );
  NAND2_X1 U17057 ( .A1(n20348), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n13704) );
  OAI211_X1 U17058 ( .C1(n21350), .C2(n13824), .A(n20344), .B(n13704), .ZN(
        P1_U2948) );
  MUX2_X1 U17059 ( .A(DATAI_8_), .B(BUF1_REG_8__SCAN_IN), .S(n20373), .Z(
        n14473) );
  NAND2_X1 U17060 ( .A1(n13845), .A2(n14473), .ZN(n13709) );
  NAND2_X1 U17061 ( .A1(n20348), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n13705) );
  OAI211_X1 U17062 ( .C1(n13706), .C2(n13824), .A(n13709), .B(n13705), .ZN(
        P1_U2945) );
  INV_X1 U17063 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13814) );
  MUX2_X1 U17064 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n20373), .Z(
        n14519) );
  NAND2_X1 U17065 ( .A1(n13845), .A2(n14519), .ZN(n20349) );
  NAND2_X1 U17066 ( .A1(n20348), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n13707) );
  OAI211_X1 U17067 ( .C1(n13814), .C2(n13824), .A(n20349), .B(n13707), .ZN(
        P1_U2950) );
  INV_X1 U17068 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20323) );
  NAND2_X1 U17069 ( .A1(n20348), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n13708) );
  OAI211_X1 U17070 ( .C1(n20323), .C2(n13824), .A(n13709), .B(n13708), .ZN(
        P1_U2960) );
  MUX2_X1 U17071 ( .A(DATAI_12_), .B(BUF1_REG_12__SCAN_IN), .S(n20373), .Z(
        n14526) );
  NAND2_X1 U17072 ( .A1(n13845), .A2(n14526), .ZN(n20346) );
  NAND2_X1 U17073 ( .A1(n20348), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n13710) );
  OAI211_X1 U17074 ( .C1(n21206), .C2(n13824), .A(n20346), .B(n13710), .ZN(
        P1_U2949) );
  MUX2_X1 U17075 ( .A(DATAI_9_), .B(BUF1_REG_9__SCAN_IN), .S(n20373), .Z(
        n14470) );
  NAND2_X1 U17076 ( .A1(n13845), .A2(n14470), .ZN(n20340) );
  NAND2_X1 U17077 ( .A1(n20348), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n13711) );
  OAI211_X1 U17078 ( .C1(n13712), .C2(n13824), .A(n20340), .B(n13711), .ZN(
        P1_U2946) );
  XNOR2_X1 U17079 ( .A(n13714), .B(n13713), .ZN(n20154) );
  INV_X1 U17080 ( .A(n20154), .ZN(n13863) );
  AOI22_X1 U17081 ( .A1(n16390), .A2(n13715), .B1(n16406), .B2(n19227), .ZN(
        n13721) );
  AOI211_X1 U17082 ( .C1(n15649), .C2(n16421), .A(n16386), .B(n13724), .ZN(
        n13718) );
  OAI22_X1 U17083 ( .A1(n15649), .A2(n16417), .B1(n16425), .B2(n13716), .ZN(
        n13717) );
  NOR3_X1 U17084 ( .A1(n13719), .A2(n13718), .A3(n13717), .ZN(n13720) );
  OAI211_X1 U17085 ( .C1(n16412), .C2(n13863), .A(n13721), .B(n13720), .ZN(
        P2_U3045) );
  OAI22_X1 U17086 ( .A1(n10580), .A2(n19176), .B1(n16416), .B2(n13722), .ZN(
        n13723) );
  AOI21_X1 U17087 ( .B1(n13725), .B2(n13724), .A(n13723), .ZN(n13742) );
  NAND2_X1 U17088 ( .A1(n13727), .A2(n13726), .ZN(n13730) );
  INV_X1 U17089 ( .A(n13728), .ZN(n13729) );
  NAND2_X1 U17090 ( .A1(n13730), .A2(n13729), .ZN(n20145) );
  NAND2_X1 U17091 ( .A1(n20145), .A2(n16387), .ZN(n13739) );
  OAI21_X1 U17092 ( .B1(n13733), .B2(n13732), .A(n13731), .ZN(n13738) );
  NAND2_X1 U17093 ( .A1(n16406), .A2(n14942), .ZN(n13737) );
  NAND3_X1 U17094 ( .A1(n16407), .A2(n13735), .A3(n13734), .ZN(n13736) );
  NAND4_X1 U17095 ( .A1(n13739), .A2(n13738), .A3(n13737), .A4(n13736), .ZN(
        n13740) );
  AOI21_X1 U17096 ( .B1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n15439), .A(
        n13740), .ZN(n13741) );
  NAND2_X1 U17097 ( .A1(n13742), .A2(n13741), .ZN(P2_U3044) );
  INV_X1 U17098 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14511) );
  INV_X1 U17099 ( .A(DATAI_15_), .ZN(n13744) );
  INV_X1 U17100 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13743) );
  MUX2_X1 U17101 ( .A(n13744), .B(n13743), .S(n20373), .Z(n14512) );
  INV_X1 U17102 ( .A(n20348), .ZN(n13825) );
  INV_X1 U17103 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20309) );
  OAI222_X1 U17104 ( .A1(n13824), .A2(n14511), .B1(n13745), .B2(n14512), .C1(
        n13825), .C2(n20309), .ZN(P1_U2967) );
  NAND2_X1 U17105 ( .A1(n19611), .A2(n19278), .ZN(n13748) );
  NAND2_X1 U17106 ( .A1(n14942), .A2(n19293), .ZN(n13747) );
  OAI211_X1 U17107 ( .C1(n19293), .C2(n10576), .A(n13748), .B(n13747), .ZN(
        P2_U2885) );
  XNOR2_X1 U17108 ( .A(n13749), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13883) );
  NAND3_X1 U17109 ( .A1(n13751), .A2(n13750), .A3(n11917), .ZN(n13755) );
  OAI211_X1 U17110 ( .C1(n13753), .C2(n21070), .A(n20405), .B(n13752), .ZN(
        n13754) );
  NAND3_X1 U17111 ( .A1(n13756), .A2(n13755), .A3(n13754), .ZN(n13758) );
  NAND2_X1 U17112 ( .A1(n13758), .A2(n13757), .ZN(n13766) );
  NAND3_X1 U17113 ( .A1(n13604), .A2(n21064), .A3(n13759), .ZN(n13761) );
  NAND3_X1 U17114 ( .A1(n13761), .A2(n20380), .A3(n13760), .ZN(n13762) );
  NAND3_X1 U17115 ( .A1(n13764), .A2(n13763), .A3(n13762), .ZN(n13765) );
  OAI211_X1 U17116 ( .C1(n9823), .C2(n13775), .A(n15816), .B(n13912), .ZN(
        n13768) );
  OR2_X1 U17117 ( .A1(n13769), .A2(n13768), .ZN(n13770) );
  XNOR2_X1 U17118 ( .A(n13772), .B(n13771), .ZN(n14413) );
  INV_X1 U17119 ( .A(n14413), .ZN(n13787) );
  OAI21_X1 U17120 ( .B1(n13775), .B2(n13773), .A(n13774), .ZN(n13776) );
  INV_X1 U17121 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n21391) );
  INV_X1 U17122 ( .A(n20361), .ZN(n13802) );
  INV_X1 U17123 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20362) );
  OAI211_X1 U17124 ( .C1(n13779), .C2(n20380), .A(n13778), .B(n13777), .ZN(
        n13780) );
  NAND2_X1 U17125 ( .A1(n20360), .A2(n20362), .ZN(n13782) );
  OR2_X1 U17126 ( .A1(n13783), .A2(n16106), .ZN(n13781) );
  INV_X1 U17127 ( .A(n16101), .ZN(n14709) );
  AOI21_X1 U17128 ( .B1(n13802), .B2(n20362), .A(n14709), .ZN(n20359) );
  OAI22_X1 U17129 ( .A1(n20369), .A2(n21391), .B1(n14826), .B2(n20359), .ZN(
        n13786) );
  INV_X1 U17130 ( .A(n14796), .ZN(n14717) );
  NOR2_X1 U17131 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n20366), .ZN(
        n13784) );
  NOR3_X1 U17132 ( .A1(n14717), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n13784), .ZN(n13785) );
  AOI211_X1 U17133 ( .C1(n13787), .C2(n16135), .A(n13786), .B(n13785), .ZN(
        n13788) );
  OAI21_X1 U17134 ( .B1(n13883), .B2(n16112), .A(n13788), .ZN(P1_U3030) );
  INV_X1 U17135 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n14409) );
  OAI21_X1 U17136 ( .B1(n13790), .B2(n13789), .A(n13897), .ZN(n14417) );
  OAI222_X1 U17137 ( .A1(n14413), .A2(n15973), .B1(n14409), .B2(n20306), .C1(
        n14417), .C2(n15974), .ZN(P1_U2871) );
  XNOR2_X1 U17138 ( .A(n13792), .B(n13791), .ZN(n13902) );
  INV_X1 U17139 ( .A(n16104), .ZN(n14707) );
  OAI21_X1 U17140 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n14707), .A(
        n16101), .ZN(n13795) );
  NAND2_X1 U17141 ( .A1(n20360), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14695) );
  INV_X1 U17142 ( .A(n14695), .ZN(n13793) );
  OAI21_X1 U17143 ( .B1(n14826), .B2(n16105), .A(n12639), .ZN(n13794) );
  OAI21_X1 U17144 ( .B1(n12639), .B2(n13795), .A(n13794), .ZN(n13804) );
  NOR2_X1 U17145 ( .A1(n12639), .A2(n14826), .ZN(n14694) );
  INV_X1 U17146 ( .A(n14694), .ZN(n13886) );
  OAI21_X1 U17147 ( .B1(n20362), .B2(n14826), .A(n12639), .ZN(n14203) );
  OAI21_X1 U17148 ( .B1(n13886), .B2(n20362), .A(n14203), .ZN(n13801) );
  INV_X1 U17149 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n21009) );
  NOR2_X1 U17150 ( .A1(n20369), .A2(n21009), .ZN(n13800) );
  OAI21_X1 U17151 ( .B1(n13798), .B2(n13797), .A(n13796), .ZN(n20301) );
  NOR2_X1 U17152 ( .A1(n20301), .A2(n20355), .ZN(n13799) );
  AOI211_X1 U17153 ( .C1(n13802), .C2(n13801), .A(n13800), .B(n13799), .ZN(
        n13803) );
  OAI211_X1 U17154 ( .C1(n13902), .C2(n16112), .A(n13804), .B(n13803), .ZN(
        P1_U3029) );
  OR2_X1 U17155 ( .A1(n9829), .A2(n14455), .ZN(n13806) );
  INV_X1 U17156 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16580) );
  NAND2_X1 U17157 ( .A1(n20373), .A2(n16580), .ZN(n13805) );
  OAI21_X1 U17158 ( .B1(n20373), .B2(DATAI_1_), .A(n13805), .ZN(n20398) );
  INV_X1 U17159 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20335) );
  OAI222_X1 U17160 ( .A1(n14530), .A2(n20398), .B1(n14527), .B2(n20335), .C1(
        n14536), .C2(n14417), .ZN(P1_U2903) );
  NAND2_X1 U17161 ( .A1(n20372), .A2(DATAI_0_), .ZN(n13808) );
  NAND2_X1 U17162 ( .A1(n20373), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13807) );
  AND2_X1 U17163 ( .A1(n13808), .A2(n13807), .ZN(n20387) );
  INV_X1 U17164 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20339) );
  OAI222_X1 U17165 ( .A1(n14038), .A2(n14536), .B1(n14530), .B2(n20387), .C1(
        n14527), .C2(n20339), .ZN(P1_U2904) );
  AOI22_X1 U17166 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20319), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n15849), .ZN(n13809) );
  OAI21_X1 U17167 ( .B1(n21179), .B2(n13816), .A(n13809), .ZN(P1_U2906) );
  AOI22_X1 U17168 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20319), .B1(n15849), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13810) );
  OAI21_X1 U17169 ( .B1(n21316), .B2(n13816), .A(n13810), .ZN(P1_U2910) );
  INV_X1 U17170 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13812) );
  AOI22_X1 U17171 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20319), .B1(n15849), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13811) );
  OAI21_X1 U17172 ( .B1(n13812), .B2(n13816), .A(n13811), .ZN(P1_U2920) );
  AOI22_X1 U17173 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20319), .B1(n15849), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13813) );
  OAI21_X1 U17174 ( .B1(n13814), .B2(n13816), .A(n13813), .ZN(P1_U2907) );
  AOI22_X1 U17175 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20319), .B1(n15849), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13815) );
  OAI21_X1 U17176 ( .B1(n12399), .B2(n13816), .A(n13815), .ZN(P1_U2919) );
  NAND2_X1 U17177 ( .A1(n14945), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n13823) );
  NAND2_X1 U17178 ( .A1(n13821), .A2(n19293), .ZN(n13822) );
  OAI211_X1 U17179 ( .C1(n20122), .C2(n19289), .A(n13823), .B(n13822), .ZN(
        P2_U2884) );
  AOI22_X1 U17180 ( .A1(n20351), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20348), .ZN(n13826) );
  INV_X1 U17181 ( .A(n20398), .ZN(n14500) );
  NAND2_X1 U17182 ( .A1(n13845), .A2(n14500), .ZN(n13832) );
  NAND2_X1 U17183 ( .A1(n13826), .A2(n13832), .ZN(P1_U2953) );
  AOI22_X1 U17184 ( .A1(n20351), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20348), .ZN(n13827) );
  INV_X1 U17185 ( .A(n20387), .ZN(n14507) );
  NAND2_X1 U17186 ( .A1(n13845), .A2(n14507), .ZN(n13853) );
  NAND2_X1 U17187 ( .A1(n13827), .A2(n13853), .ZN(P1_U2952) );
  AOI22_X1 U17188 ( .A1(n20351), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20348), .ZN(n13829) );
  INV_X1 U17189 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16574) );
  NAND2_X1 U17190 ( .A1(n20373), .A2(n16574), .ZN(n13828) );
  OAI21_X1 U17191 ( .B1(n20373), .B2(DATAI_4_), .A(n13828), .ZN(n20422) );
  INV_X1 U17192 ( .A(n20422), .ZN(n14488) );
  NAND2_X1 U17193 ( .A1(n13845), .A2(n14488), .ZN(n13847) );
  NAND2_X1 U17194 ( .A1(n13829), .A2(n13847), .ZN(P1_U2956) );
  AOI22_X1 U17195 ( .A1(n20351), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20348), .ZN(n13831) );
  NAND2_X1 U17196 ( .A1(n20373), .A2(n16578), .ZN(n13830) );
  OAI21_X1 U17197 ( .B1(n20373), .B2(DATAI_2_), .A(n13830), .ZN(n20407) );
  INV_X1 U17198 ( .A(n20407), .ZN(n14496) );
  NAND2_X1 U17199 ( .A1(n13845), .A2(n14496), .ZN(n13836) );
  NAND2_X1 U17200 ( .A1(n13831), .A2(n13836), .ZN(P1_U2939) );
  AOI22_X1 U17201 ( .A1(n20351), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20348), .ZN(n13833) );
  NAND2_X1 U17202 ( .A1(n13833), .A2(n13832), .ZN(P1_U2938) );
  AOI22_X1 U17203 ( .A1(n20351), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20348), .ZN(n13835) );
  INV_X1 U17204 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16576) );
  NAND2_X1 U17205 ( .A1(n20373), .A2(n16576), .ZN(n13834) );
  OAI21_X1 U17206 ( .B1(n20373), .B2(DATAI_3_), .A(n13834), .ZN(n20415) );
  INV_X1 U17207 ( .A(n20415), .ZN(n14492) );
  NAND2_X1 U17208 ( .A1(n13845), .A2(n14492), .ZN(n13842) );
  NAND2_X1 U17209 ( .A1(n13835), .A2(n13842), .ZN(P1_U2955) );
  AOI22_X1 U17210 ( .A1(n20351), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20348), .ZN(n13837) );
  NAND2_X1 U17211 ( .A1(n13837), .A2(n13836), .ZN(P1_U2954) );
  AOI22_X1 U17212 ( .A1(n20351), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20348), .ZN(n13839) );
  INV_X1 U17213 ( .A(DATAI_7_), .ZN(n21394) );
  NAND2_X1 U17214 ( .A1(n20373), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13838) );
  OAI21_X1 U17215 ( .B1(n20373), .B2(n21394), .A(n13838), .ZN(n14477) );
  NAND2_X1 U17216 ( .A1(n13845), .A2(n14477), .ZN(n13849) );
  NAND2_X1 U17217 ( .A1(n13839), .A2(n13849), .ZN(P1_U2959) );
  AOI22_X1 U17218 ( .A1(n20351), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20348), .ZN(n13841) );
  INV_X1 U17219 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16570) );
  NAND2_X1 U17220 ( .A1(n20373), .A2(n16570), .ZN(n13840) );
  OAI21_X1 U17221 ( .B1(n20373), .B2(DATAI_6_), .A(n13840), .ZN(n20436) );
  INV_X1 U17222 ( .A(n20436), .ZN(n14480) );
  NAND2_X1 U17223 ( .A1(n13845), .A2(n14480), .ZN(n13851) );
  NAND2_X1 U17224 ( .A1(n13841), .A2(n13851), .ZN(P1_U2958) );
  AOI22_X1 U17225 ( .A1(n20351), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20348), .ZN(n13843) );
  NAND2_X1 U17226 ( .A1(n13843), .A2(n13842), .ZN(P1_U2940) );
  AOI22_X1 U17227 ( .A1(n20351), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20348), .ZN(n13846) );
  INV_X1 U17228 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16572) );
  NAND2_X1 U17229 ( .A1(n20373), .A2(n16572), .ZN(n13844) );
  OAI21_X1 U17230 ( .B1(n20373), .B2(DATAI_5_), .A(n13844), .ZN(n20429) );
  INV_X1 U17231 ( .A(n20429), .ZN(n14484) );
  NAND2_X1 U17232 ( .A1(n13845), .A2(n14484), .ZN(n13855) );
  NAND2_X1 U17233 ( .A1(n13846), .A2(n13855), .ZN(P1_U2942) );
  AOI22_X1 U17234 ( .A1(n20351), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20348), .ZN(n13848) );
  NAND2_X1 U17235 ( .A1(n13848), .A2(n13847), .ZN(P1_U2941) );
  AOI22_X1 U17236 ( .A1(n20351), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20348), .ZN(n13850) );
  NAND2_X1 U17237 ( .A1(n13850), .A2(n13849), .ZN(P1_U2944) );
  AOI22_X1 U17238 ( .A1(n20351), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20348), .ZN(n13852) );
  NAND2_X1 U17239 ( .A1(n13852), .A2(n13851), .ZN(P1_U2943) );
  AOI22_X1 U17240 ( .A1(n20351), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20348), .ZN(n13854) );
  NAND2_X1 U17241 ( .A1(n13854), .A2(n13853), .ZN(P1_U2937) );
  AOI22_X1 U17242 ( .A1(n20351), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20348), .ZN(n13856) );
  NAND2_X1 U17243 ( .A1(n13856), .A2(n13855), .ZN(P1_U2957) );
  INV_X1 U17244 ( .A(n19283), .ZN(n19212) );
  XOR2_X1 U17245 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n19212), .Z(n13862)
         );
  OR2_X1 U17246 ( .A1(n14109), .A2(n13858), .ZN(n13859) );
  AND2_X1 U17247 ( .A1(n13857), .A2(n13859), .ZN(n19195) );
  INV_X1 U17248 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n19202) );
  NOR2_X1 U17249 ( .A1(n19293), .A2(n19202), .ZN(n13860) );
  AOI21_X1 U17250 ( .B1(n19195), .B2(n19293), .A(n13860), .ZN(n13861) );
  OAI21_X1 U17251 ( .B1(n13862), .B2(n19289), .A(n13861), .ZN(P2_U2882) );
  XNOR2_X1 U17252 ( .A(n19611), .B(n20145), .ZN(n13867) );
  NAND2_X1 U17253 ( .A1(n20130), .A2(n13863), .ZN(n13864) );
  OAI21_X1 U17254 ( .B1(n20130), .B2(n13863), .A(n13864), .ZN(n19359) );
  NOR2_X1 U17255 ( .A1(n19359), .A2(n19360), .ZN(n19358) );
  INV_X1 U17256 ( .A(n13864), .ZN(n13865) );
  NOR2_X1 U17257 ( .A1(n19358), .A2(n13865), .ZN(n13866) );
  NOR2_X1 U17258 ( .A1(n13866), .A2(n13867), .ZN(n19332) );
  AOI21_X1 U17259 ( .B1(n13867), .B2(n13866), .A(n19332), .ZN(n13870) );
  AOI22_X1 U17260 ( .A1(n20145), .A2(n19357), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19356), .ZN(n13869) );
  NAND2_X1 U17261 ( .A1(n19325), .A2(n16291), .ZN(n13868) );
  OAI211_X1 U17262 ( .C1(n13870), .C2(n19361), .A(n13869), .B(n13868), .ZN(
        P2_U2917) );
  NOR2_X1 U17263 ( .A1(n19212), .A2(n13871), .ZN(n13873) );
  OR2_X1 U17264 ( .A1(n19212), .A2(n13872), .ZN(n13903) );
  OAI211_X1 U17265 ( .C1(n13873), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n19278), .B(n13903), .ZN(n13877) );
  NAND2_X1 U17266 ( .A1(n13857), .A2(n13874), .ZN(n13875) );
  NAND2_X1 U17267 ( .A1(n13905), .A2(n13875), .ZN(n16368) );
  INV_X1 U17268 ( .A(n16368), .ZN(n19185) );
  NAND2_X1 U17269 ( .A1(n19185), .A2(n19293), .ZN(n13876) );
  OAI211_X1 U17270 ( .C1(n19293), .C2(n13878), .A(n13877), .B(n13876), .ZN(
        P2_U2881) );
  INV_X1 U17271 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13881) );
  OAI22_X1 U17272 ( .A1(n16038), .A2(n13881), .B1(n20369), .B2(n21391), .ZN(
        n13880) );
  NOR2_X1 U17273 ( .A1(n14417), .A2(n14689), .ZN(n13879) );
  AOI211_X1 U17274 ( .C1(n16033), .C2(n13881), .A(n13880), .B(n13879), .ZN(
        n13882) );
  OAI21_X1 U17275 ( .B1(n13883), .B2(n20187), .A(n13882), .ZN(P1_U2998) );
  XNOR2_X1 U17276 ( .A(n13885), .B(n13884), .ZN(n13996) );
  NAND2_X1 U17277 ( .A1(n14203), .A2(n16114), .ZN(n14128) );
  INV_X1 U17278 ( .A(n14128), .ZN(n13890) );
  NAND2_X1 U17279 ( .A1(n13796), .A2(n13887), .ZN(n13888) );
  NAND2_X1 U17280 ( .A1(n13988), .A2(n13888), .ZN(n14055) );
  INV_X1 U17281 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n21012) );
  OAI22_X1 U17282 ( .A1(n14055), .A2(n20355), .B1(n21012), .B2(n20369), .ZN(
        n13889) );
  AOI21_X1 U17283 ( .B1(n13890), .B2(n13985), .A(n13889), .ZN(n13893) );
  OAI21_X1 U17284 ( .B1(n14707), .B2(n14694), .A(n16101), .ZN(n14205) );
  INV_X1 U17285 ( .A(n14205), .ZN(n13891) );
  OAI21_X1 U17286 ( .B1(n20361), .B2(n14203), .A(n13891), .ZN(n14020) );
  NAND2_X1 U17287 ( .A1(n14020), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13892) );
  OAI211_X1 U17288 ( .C1(n13996), .C2(n16112), .A(n13893), .B(n13892), .ZN(
        P1_U3028) );
  CLKBUF_X1 U17289 ( .A(n13894), .Z(n13898) );
  INV_X1 U17290 ( .A(n13895), .ZN(n13896) );
  AOI21_X1 U17291 ( .B1(n13898), .B2(n13897), .A(n13896), .ZN(n20304) );
  AOI22_X1 U17292 ( .A1(n16027), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n16106), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13899) );
  OAI21_X1 U17293 ( .B1(n20290), .B2(n16031), .A(n13899), .ZN(n13900) );
  AOI21_X1 U17294 ( .B1(n20304), .B2(n20374), .A(n13900), .ZN(n13901) );
  OAI21_X1 U17295 ( .B1(n20187), .B2(n13902), .A(n13901), .ZN(P1_U2997) );
  XOR2_X1 U17296 ( .A(n13903), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n13908)
         );
  AND2_X1 U17297 ( .A1(n13905), .A2(n13904), .ZN(n13906) );
  OR2_X1 U17298 ( .A1(n13906), .A2(n9880), .ZN(n19171) );
  MUX2_X1 U17299 ( .A(n19171), .B(n10853), .S(n14945), .Z(n13907) );
  OAI21_X1 U17300 ( .B1(n13908), .B2(n19289), .A(n13907), .ZN(P2_U2880) );
  NOR2_X1 U17301 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n16145), .ZN(n13938) );
  INV_X1 U17302 ( .A(n13909), .ZN(n20384) );
  NOR2_X1 U17303 ( .A1(n13910), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13927) );
  INV_X1 U17304 ( .A(n13927), .ZN(n13911) );
  NAND2_X1 U17305 ( .A1(n13911), .A2(n10138), .ZN(n13915) );
  NOR3_X1 U17306 ( .A1(n14824), .A2(n13923), .A3(n13915), .ZN(n13919) );
  INV_X1 U17307 ( .A(n15803), .ZN(n14820) );
  XNOR2_X1 U17308 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13917) );
  INV_X1 U17309 ( .A(n13912), .ZN(n13913) );
  OR2_X1 U17310 ( .A1(n13914), .A2(n13913), .ZN(n13932) );
  INV_X1 U17311 ( .A(n13932), .ZN(n13916) );
  INV_X1 U17312 ( .A(n13915), .ZN(n14833) );
  OAI22_X1 U17313 ( .A1(n14820), .A2(n13917), .B1(n13916), .B2(n14833), .ZN(
        n13918) );
  AOI211_X1 U17314 ( .C1(n20384), .C2(n14824), .A(n13919), .B(n13918), .ZN(
        n14838) );
  INV_X1 U17315 ( .A(n14838), .ZN(n13920) );
  MUX2_X1 U17316 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n13920), .S(
        n15805), .Z(n15811) );
  AOI22_X1 U17317 ( .A1(n13938), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n16145), .B2(n15811), .ZN(n13940) );
  OAI21_X1 U17318 ( .B1(n13921), .B2(n13928), .A(n9849), .ZN(n13922) );
  INV_X1 U17319 ( .A(n13922), .ZN(n14840) );
  OR2_X1 U17320 ( .A1(n13923), .A2(n14840), .ZN(n13935) );
  XNOR2_X1 U17321 ( .A(n13924), .B(n13928), .ZN(n13933) );
  INV_X1 U17322 ( .A(n13925), .ZN(n13926) );
  OAI21_X1 U17323 ( .B1(n13927), .B2(n13928), .A(n13926), .ZN(n13930) );
  NAND2_X1 U17324 ( .A1(n13910), .A2(n13928), .ZN(n13929) );
  NAND2_X1 U17325 ( .A1(n13930), .A2(n13929), .ZN(n13931) );
  AOI22_X1 U17326 ( .A1(n15803), .A2(n13933), .B1(n13932), .B2(n13931), .ZN(
        n13934) );
  OAI21_X1 U17327 ( .B1(n14824), .B2(n13935), .A(n13934), .ZN(n13936) );
  AOI21_X1 U17328 ( .B1(n20659), .B2(n14824), .A(n13936), .ZN(n14842) );
  NOR2_X1 U17329 ( .A1(n15805), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13937) );
  AOI21_X1 U17330 ( .B1(n14842), .B2(n15805), .A(n13937), .ZN(n15801) );
  AOI22_X1 U17331 ( .A1(n13938), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n16145), .B2(n15801), .ZN(n13939) );
  NOR2_X1 U17332 ( .A1(n13940), .A2(n13939), .ZN(n15819) );
  INV_X1 U17333 ( .A(n13941), .ZN(n14821) );
  NAND2_X1 U17334 ( .A1(n15819), .A2(n14821), .ZN(n13965) );
  AND2_X1 U17335 ( .A1(n15805), .A2(n16145), .ZN(n13943) );
  NAND3_X1 U17336 ( .A1(n20271), .A2(n13942), .A3(n13943), .ZN(n13946) );
  INV_X1 U17337 ( .A(n13943), .ZN(n13944) );
  NAND3_X1 U17338 ( .A1(n13944), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(
        n21319), .ZN(n13945) );
  AND3_X1 U17339 ( .A1(n13965), .A2(n15822), .A3(n21319), .ZN(n13947) );
  INV_X1 U17340 ( .A(n15834), .ZN(n21077) );
  AND2_X1 U17341 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20799), .ZN(n13967) );
  AOI21_X1 U17342 ( .B1(n13948), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20926), 
        .ZN(n20929) );
  OAI21_X1 U17343 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n13948), .A(n20929), 
        .ZN(n13949) );
  OAI21_X1 U17344 ( .B1(n20660), .B2(n13967), .A(n13949), .ZN(n13950) );
  NAND2_X1 U17345 ( .A1(n20370), .A2(n13950), .ZN(n13951) );
  OAI21_X1 U17346 ( .B1(n20370), .B2(n20791), .A(n13951), .ZN(P1_U3477) );
  MUX2_X1 U17347 ( .A(n20925), .B(n20629), .S(n13948), .Z(n13955) );
  INV_X1 U17348 ( .A(n13953), .ZN(n13954) );
  AOI21_X1 U17349 ( .B1(n13955), .B2(n20763), .A(n13960), .ZN(n13958) );
  NAND2_X1 U17350 ( .A1(n20933), .A2(n20848), .ZN(n20786) );
  INV_X1 U17351 ( .A(n20659), .ZN(n13956) );
  OAI22_X1 U17352 ( .A1(n13953), .A2(n20786), .B1(n13956), .B2(n13967), .ZN(
        n13957) );
  OAI21_X1 U17353 ( .B1(n13958), .B2(n13957), .A(n20370), .ZN(n13959) );
  OAI21_X1 U17354 ( .B1(n12729), .B2(n20370), .A(n13959), .ZN(P1_U3475) );
  NOR2_X1 U17355 ( .A1(n13909), .A2(n13967), .ZN(n13963) );
  INV_X1 U17356 ( .A(n13948), .ZN(n20633) );
  NOR2_X1 U17357 ( .A1(n20633), .A2(n13960), .ZN(n13961) );
  MUX2_X1 U17358 ( .A(n13961), .B(n20929), .S(n12640), .Z(n13962) );
  OAI21_X1 U17359 ( .B1(n13963), .B2(n13962), .A(n20370), .ZN(n13964) );
  OAI21_X1 U17360 ( .B1(n12753), .B2(n20370), .A(n13964), .ZN(P1_U3476) );
  AND2_X1 U17361 ( .A1(n15822), .A2(n20989), .ZN(n13966) );
  AND2_X1 U17362 ( .A1(n13966), .A2(n13965), .ZN(n15829) );
  OAI22_X1 U17363 ( .A1(n20479), .A2(n20926), .B1(n13968), .B2(n13967), .ZN(
        n13969) );
  OAI21_X1 U17364 ( .B1(n15829), .B2(n13969), .A(n20370), .ZN(n13970) );
  OAI21_X1 U17365 ( .B1(n20370), .B2(n20843), .A(n13970), .ZN(P1_U3478) );
  CLKBUF_X1 U17366 ( .A(n13972), .Z(n13998) );
  OAI21_X1 U17367 ( .B1(n13971), .B2(n13973), .A(n13998), .ZN(n14067) );
  INV_X1 U17368 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n21199) );
  OAI222_X1 U17369 ( .A1(n14067), .A2(n15974), .B1(n20306), .B2(n21199), .C1(
        n14055), .C2(n15973), .ZN(P1_U2869) );
  INV_X1 U17370 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n19165) );
  INV_X1 U17371 ( .A(n13974), .ZN(n19284) );
  OAI211_X1 U17372 ( .C1(n19284), .C2(n13976), .A(n19278), .B(n13975), .ZN(
        n13981) );
  OR2_X1 U17373 ( .A1(n9971), .A2(n13978), .ZN(n13979) );
  AND2_X1 U17374 ( .A1(n13977), .A2(n13979), .ZN(n19159) );
  NAND2_X1 U17375 ( .A1(n19159), .A2(n19293), .ZN(n13980) );
  OAI211_X1 U17376 ( .C1(n19293), .C2(n19165), .A(n13981), .B(n13980), .ZN(
        P2_U2878) );
  INV_X1 U17377 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20333) );
  INV_X1 U17378 ( .A(n20304), .ZN(n13982) );
  OAI222_X1 U17379 ( .A1(n14530), .A2(n20407), .B1(n14527), .B2(n20333), .C1(
        n14536), .C2(n13982), .ZN(P1_U2902) );
  INV_X1 U17380 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20331) );
  OAI222_X1 U17381 ( .A1(n14530), .A2(n20415), .B1(n14527), .B2(n20331), .C1(
        n14536), .C2(n14067), .ZN(P1_U2901) );
  XNOR2_X1 U17382 ( .A(n13984), .B(n13983), .ZN(n14014) );
  AOI21_X1 U17383 ( .B1(n13986), .B2(n13985), .A(n14128), .ZN(n13987) );
  NAND2_X1 U17384 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14019) );
  AOI22_X1 U17385 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n14020), .B1(
        n13987), .B2(n14019), .ZN(n13991) );
  AOI21_X1 U17386 ( .B1(n13989), .B2(n13988), .A(n9950), .ZN(n20273) );
  NOR2_X1 U17387 ( .A1(n20369), .A2(n21332), .ZN(n14010) );
  AOI21_X1 U17388 ( .B1(n20273), .B2(n16135), .A(n14010), .ZN(n13990) );
  OAI211_X1 U17389 ( .C1(n16112), .C2(n14014), .A(n13991), .B(n13990), .ZN(
        P1_U3027) );
  INV_X1 U17390 ( .A(n14067), .ZN(n13994) );
  AOI22_X1 U17391 ( .A1(n16027), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n16106), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n13992) );
  OAI21_X1 U17392 ( .B1(n14056), .B2(n16031), .A(n13992), .ZN(n13993) );
  AOI21_X1 U17393 ( .B1(n13994), .B2(n20374), .A(n13993), .ZN(n13995) );
  OAI21_X1 U17394 ( .B1(n20187), .B2(n13996), .A(n13995), .ZN(P1_U2996) );
  AOI21_X1 U17395 ( .B1(n13999), .B2(n13998), .A(n13997), .ZN(n20282) );
  INV_X1 U17396 ( .A(n20282), .ZN(n14001) );
  INV_X1 U17397 ( .A(n20306), .ZN(n14433) );
  AOI22_X1 U17398 ( .A1(n20273), .A2(n13038), .B1(P1_EBX_REG_4__SCAN_IN), .B2(
        n14433), .ZN(n14000) );
  OAI21_X1 U17399 ( .B1(n14001), .B2(n15974), .A(n14000), .ZN(P1_U2868) );
  INV_X1 U17400 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20329) );
  OAI222_X1 U17401 ( .A1(n14001), .A2(n14536), .B1(n14527), .B2(n20329), .C1(
        n14530), .C2(n20422), .ZN(P1_U2900) );
  NOR2_X1 U17402 ( .A1(n13975), .A2(n14002), .ZN(n14005) );
  OAI211_X1 U17403 ( .C1(n14005), .C2(n14004), .A(n10289), .B(n19278), .ZN(
        n14009) );
  NAND2_X1 U17404 ( .A1(n16324), .A2(n14006), .ZN(n14007) );
  NAND2_X1 U17405 ( .A1(n19135), .A2(n19293), .ZN(n14008) );
  OAI211_X1 U17406 ( .C1(n19293), .C2(n19129), .A(n14009), .B(n14008), .ZN(
        P2_U2876) );
  AOI21_X1 U17407 ( .B1(n16027), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n14010), .ZN(n14011) );
  OAI21_X1 U17408 ( .B1(n20267), .B2(n16031), .A(n14011), .ZN(n14012) );
  AOI21_X1 U17409 ( .B1(n20282), .B2(n20374), .A(n14012), .ZN(n14013) );
  OAI21_X1 U17410 ( .B1(n20187), .B2(n14014), .A(n14013), .ZN(P1_U2995) );
  XNOR2_X1 U17411 ( .A(n14016), .B(n14015), .ZN(n16032) );
  NOR2_X1 U17412 ( .A1(n9950), .A2(n14017), .ZN(n14018) );
  OR2_X1 U17413 ( .A1(n14050), .A2(n14018), .ZN(n20263) );
  INV_X1 U17414 ( .A(n20263), .ZN(n14024) );
  NAND2_X1 U17415 ( .A1(n16106), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n16036) );
  INV_X1 U17416 ( .A(n16036), .ZN(n14023) );
  NOR2_X1 U17417 ( .A1(n14019), .A2(n14128), .ZN(n14021) );
  NAND3_X1 U17418 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14201) );
  AOI21_X1 U17419 ( .B1(n14796), .B2(n14201), .A(n14020), .ZN(n14129) );
  INV_X1 U17420 ( .A(n14129), .ZN(n14051) );
  MUX2_X1 U17421 ( .A(n14021), .B(n14051), .S(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(n14022) );
  AOI211_X1 U17422 ( .C1(n16135), .C2(n14024), .A(n14023), .B(n14022), .ZN(
        n14025) );
  OAI21_X1 U17423 ( .B1(n16112), .B2(n16032), .A(n14025), .ZN(P1_U3026) );
  NAND2_X1 U17424 ( .A1(n14029), .A2(n14026), .ZN(n14027) );
  NAND2_X1 U17425 ( .A1(n14027), .A2(n15960), .ZN(n20297) );
  INV_X1 U17426 ( .A(n20297), .ZN(n14416) );
  INV_X1 U17427 ( .A(n14028), .ZN(n21074) );
  AND2_X1 U17428 ( .A1(n14029), .A2(n21074), .ZN(n20286) );
  NAND2_X1 U17429 ( .A1(n20250), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n14035) );
  INV_X1 U17430 ( .A(n20354), .ZN(n14030) );
  NAND2_X1 U17431 ( .A1(n20272), .A2(n14030), .ZN(n14034) );
  NAND2_X1 U17432 ( .A1(n20292), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n14033) );
  NOR2_X1 U17433 ( .A1(n14549), .A2(n16145), .ZN(n14031) );
  OAI21_X1 U17434 ( .B1(n20255), .B2(n20254), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14032) );
  NAND4_X1 U17435 ( .A1(n14035), .A2(n14034), .A3(n14033), .A4(n14032), .ZN(
        n14036) );
  AOI21_X1 U17436 ( .B1(n12075), .B2(n20286), .A(n14036), .ZN(n14037) );
  OAI21_X1 U17437 ( .B1(n14038), .B2(n14416), .A(n14037), .ZN(P1_U2840) );
  INV_X1 U17438 ( .A(n14040), .ZN(n14041) );
  NAND2_X1 U17439 ( .A1(n14042), .A2(n14041), .ZN(n14043) );
  AND2_X1 U17440 ( .A1(n14039), .A2(n14043), .ZN(n20265) );
  OAI22_X1 U17441 ( .A1(n20263), .A2(n15973), .B1(n21376), .B2(n20306), .ZN(
        n14044) );
  AOI21_X1 U17442 ( .B1(n20265), .B2(n20303), .A(n14044), .ZN(n14045) );
  INV_X1 U17443 ( .A(n14045), .ZN(P1_U2867) );
  INV_X1 U17444 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n20327) );
  INV_X1 U17445 ( .A(n20265), .ZN(n14046) );
  OAI222_X1 U17446 ( .A1(n14530), .A2(n20429), .B1(n14527), .B2(n20327), .C1(
        n14536), .C2(n14046), .ZN(P1_U2899) );
  XNOR2_X1 U17447 ( .A(n14048), .B(n14047), .ZN(n14127) );
  OAI21_X1 U17448 ( .B1(n14050), .B2(n14049), .A(n14131), .ZN(n14071) );
  INV_X1 U17449 ( .A(n14071), .ZN(n20239) );
  INV_X1 U17450 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n21365) );
  NOR2_X1 U17451 ( .A1(n20369), .A2(n21365), .ZN(n14123) );
  NOR2_X1 U17452 ( .A1(n14201), .A2(n14128), .ZN(n14052) );
  MUX2_X1 U17453 ( .A(n14052), .B(n14051), .S(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .Z(n14053) );
  AOI211_X1 U17454 ( .C1(n16135), .C2(n20239), .A(n14123), .B(n14053), .ZN(
        n14054) );
  OAI21_X1 U17455 ( .B1(n16112), .B2(n14127), .A(n14054), .ZN(P1_U3025) );
  INV_X1 U17456 ( .A(n14055), .ZN(n14064) );
  NAND3_X1 U17457 ( .A1(n21012), .A2(P1_REIP_REG_2__SCAN_IN), .A3(
        P1_REIP_REG_1__SCAN_IN), .ZN(n14060) );
  INV_X1 U17458 ( .A(n14056), .ZN(n14057) );
  AOI22_X1 U17459 ( .A1(n14057), .A2(n20254), .B1(n20255), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14059) );
  NAND2_X1 U17460 ( .A1(n20292), .A2(P1_EBX_REG_3__SCAN_IN), .ZN(n14058) );
  OAI211_X1 U17461 ( .C1(n14060), .C2(n20276), .A(n14059), .B(n14058), .ZN(
        n14063) );
  INV_X1 U17462 ( .A(n14408), .ZN(n20252) );
  NAND2_X1 U17463 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .ZN(n14061) );
  OAI21_X1 U17464 ( .B1(n20252), .B2(n14061), .A(n20250), .ZN(n20299) );
  NOR2_X1 U17465 ( .A1(n20299), .A2(n21012), .ZN(n14062) );
  AOI211_X1 U17466 ( .C1(n14064), .C2(n20272), .A(n14063), .B(n14062), .ZN(
        n14066) );
  NAND2_X1 U17467 ( .A1(n20659), .A2(n20286), .ZN(n14065) );
  OAI211_X1 U17468 ( .C1(n14067), .C2(n14416), .A(n14066), .B(n14065), .ZN(
        P1_U2837) );
  AND2_X1 U17469 ( .A1(n14039), .A2(n14068), .ZN(n14070) );
  OR2_X1 U17470 ( .A1(n14070), .A2(n14069), .ZN(n14122) );
  OAI222_X1 U17471 ( .A1(n14122), .A2(n15974), .B1(n21328), .B2(n20306), .C1(
        n14071), .C2(n15973), .ZN(P1_U2866) );
  MUX2_X1 U17472 ( .A(n14073), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .S(
        n14072), .Z(n14075) );
  XNOR2_X1 U17473 ( .A(n14075), .B(n14074), .ZN(n14095) );
  XOR2_X1 U17474 ( .A(n14077), .B(n14076), .Z(n14093) );
  OAI21_X1 U17475 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n14078), .A(
        n14867), .ZN(n14868) );
  AOI22_X1 U17476 ( .A1(n16316), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n19414), .B2(P2_REIP_REG_3__SCAN_IN), .ZN(n14080) );
  NAND2_X1 U17477 ( .A1(n13821), .A2(n16363), .ZN(n14079) );
  OAI211_X1 U17478 ( .C1(n16355), .C2(n14868), .A(n14080), .B(n14079), .ZN(
        n14081) );
  AOI21_X1 U17479 ( .B1(n14093), .B2(n19421), .A(n14081), .ZN(n14082) );
  OAI21_X1 U17480 ( .B1(n14095), .B2(n19417), .A(n14082), .ZN(P2_U3011) );
  OR2_X1 U17481 ( .A1(n14084), .A2(n14083), .ZN(n14086) );
  NAND2_X1 U17482 ( .A1(n14086), .A2(n14085), .ZN(n20137) );
  OAI21_X1 U17483 ( .B1(n15480), .B2(n14088), .A(n14087), .ZN(n15608) );
  INV_X1 U17484 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n20060) );
  NOR2_X1 U17485 ( .A1(n20060), .A2(n19176), .ZN(n14089) );
  AOI221_X1 U17486 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n15608), .C1(
        n14073), .C2(n14110), .A(n14089), .ZN(n14091) );
  NAND2_X1 U17487 ( .A1(n13821), .A2(n16406), .ZN(n14090) );
  OAI211_X1 U17488 ( .C1(n20137), .C2(n16412), .A(n14091), .B(n14090), .ZN(
        n14092) );
  AOI21_X1 U17489 ( .B1(n16390), .B2(n14093), .A(n14092), .ZN(n14094) );
  OAI21_X1 U17490 ( .B1(n14095), .B2(n16425), .A(n14094), .ZN(P2_U3043) );
  OAI222_X1 U17491 ( .A1(n14530), .A2(n20436), .B1(n14527), .B2(n12197), .C1(
        n14536), .C2(n14122), .ZN(P1_U2898) );
  XNOR2_X1 U17492 ( .A(n14096), .B(n19264), .ZN(n14101) );
  OR2_X1 U17493 ( .A1(n15305), .A2(n14098), .ZN(n14099) );
  NAND2_X1 U17494 ( .A1(n14097), .A2(n14099), .ZN(n19113) );
  INV_X1 U17495 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n19118) );
  MUX2_X1 U17496 ( .A(n19113), .B(n19118), .S(n14945), .Z(n14100) );
  OAI21_X1 U17497 ( .B1(n14101), .B2(n19289), .A(n14100), .ZN(P2_U2874) );
  XNOR2_X1 U17498 ( .A(n14103), .B(n14102), .ZN(n19418) );
  AOI21_X1 U17499 ( .B1(n14105), .B2(n14085), .A(n14104), .ZN(n19339) );
  NOR2_X1 U17500 ( .A1(n14107), .A2(n14106), .ZN(n14108) );
  OR2_X1 U17501 ( .A1(n14109), .A2(n14108), .ZN(n19415) );
  NOR2_X1 U17502 ( .A1(n19415), .A2(n16413), .ZN(n14113) );
  NAND2_X1 U17503 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n14110), .ZN(
        n15621) );
  AOI21_X1 U17504 ( .B1(n16420), .B2(n14073), .A(n15608), .ZN(n15630) );
  NAND2_X1 U17505 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19414), .ZN(n14111) );
  OAI221_X1 U17506 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n15621), .C1(
        n15622), .C2(n15630), .A(n14111), .ZN(n14112) );
  AOI211_X1 U17507 ( .C1(n16387), .C2(n19339), .A(n14113), .B(n14112), .ZN(
        n14118) );
  NAND2_X1 U17508 ( .A1(n14115), .A2(n14114), .ZN(n14116) );
  XNOR2_X1 U17509 ( .A(n14116), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19420) );
  NAND2_X1 U17510 ( .A1(n19420), .A2(n16390), .ZN(n14117) );
  OAI211_X1 U17511 ( .C1(n16425), .C2(n19418), .A(n14118), .B(n14117), .ZN(
        P2_U3042) );
  OR2_X1 U17512 ( .A1(n14069), .A2(n14120), .ZN(n14121) );
  AND2_X1 U17513 ( .A1(n14119), .A2(n14121), .ZN(n20237) );
  INV_X1 U17514 ( .A(n20237), .ZN(n14141) );
  INV_X1 U17515 ( .A(n14477), .ZN(n20447) );
  OAI222_X1 U17516 ( .A1(n14141), .A2(n14536), .B1(n14530), .B2(n20447), .C1(
        n14527), .C2(n12206), .ZN(P1_U2897) );
  INV_X1 U17517 ( .A(n14122), .ZN(n20246) );
  AOI21_X1 U17518 ( .B1(n16027), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n14123), .ZN(n14124) );
  OAI21_X1 U17519 ( .B1(n20240), .B2(n16031), .A(n14124), .ZN(n14125) );
  AOI21_X1 U17520 ( .B1(n20246), .B2(n20374), .A(n14125), .ZN(n14126) );
  OAI21_X1 U17521 ( .B1(n14127), .B2(n20187), .A(n14126), .ZN(P1_U2993) );
  NOR3_X1 U17522 ( .A1(n14202), .A2(n14201), .A3(n14128), .ZN(n16139) );
  INV_X1 U17523 ( .A(n16139), .ZN(n14140) );
  OAI21_X1 U17524 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n14717), .A(
        n14129), .ZN(n16137) );
  NAND2_X1 U17525 ( .A1(n14131), .A2(n14130), .ZN(n14132) );
  NAND2_X1 U17526 ( .A1(n14185), .A2(n14132), .ZN(n20235) );
  OAI22_X1 U17527 ( .A1(n20235), .A2(n20355), .B1(n21379), .B2(n20369), .ZN(
        n14133) );
  AOI21_X1 U17528 ( .B1(n16137), .B2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n14133), .ZN(n14139) );
  NAND2_X1 U17529 ( .A1(n14135), .A2(n14134), .ZN(n14136) );
  XNOR2_X1 U17530 ( .A(n14137), .B(n14136), .ZN(n16028) );
  NAND2_X1 U17531 ( .A1(n16028), .A2(n20357), .ZN(n14138) );
  OAI211_X1 U17532 ( .C1(n14140), .C2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n14139), .B(n14138), .ZN(P1_U3024) );
  OAI222_X1 U17533 ( .A1(n20235), .A2(n15973), .B1(n20306), .B2(n10025), .C1(
        n14141), .C2(n15974), .ZN(P1_U2865) );
  INV_X1 U17534 ( .A(n19232), .ZN(n19247) );
  NAND2_X1 U17535 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n14880), .ZN(
        n14883) );
  INV_X1 U17536 ( .A(n14883), .ZN(n14142) );
  NAND2_X1 U17537 ( .A1(n15193), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15182) );
  INV_X1 U17538 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15171) );
  INV_X1 U17539 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15158) );
  INV_X1 U17540 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14143) );
  INV_X1 U17541 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14258) );
  AOI22_X1 U17542 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16491), .ZN(n19256) );
  AOI22_X1 U17543 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n19233), .B2(n16491), .ZN(
        n15648) );
  NAND2_X1 U17544 ( .A1(n19256), .A2(n15648), .ZN(n15647) );
  NOR2_X1 U17545 ( .A1(n14934), .A2(n15647), .ZN(n14869) );
  NOR2_X1 U17546 ( .A1(n19192), .A2(n14869), .ZN(n14145) );
  XNOR2_X1 U17547 ( .A(n14145), .B(n14868), .ZN(n14146) );
  NOR4_X1 U17548 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(P2_STATE2_REG_0__SCAN_IN), .A4(n16479), .ZN(n14153) );
  NAND2_X1 U17549 ( .A1(n14146), .A2(n19198), .ZN(n14169) );
  NAND2_X1 U17550 ( .A1(n19612), .A2(n14851), .ZN(n14157) );
  NOR2_X1 U17551 ( .A1(n14159), .A2(n14157), .ZN(n14147) );
  NOR2_X1 U17552 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n14148), .ZN(n16158) );
  INV_X1 U17553 ( .A(n14157), .ZN(n14149) );
  OAI21_X4 U17554 ( .B1(n14152), .B2(n16158), .A(n14151), .ZN(n19250) );
  INV_X1 U17555 ( .A(n19250), .ZN(n19203) );
  NOR3_X1 U17556 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n15864), .A3(n20136), 
        .ZN(n16475) );
  INV_X1 U17557 ( .A(n16475), .ZN(n14154) );
  NAND2_X1 U17558 ( .A1(n20032), .A2(n14154), .ZN(n14155) );
  NAND2_X1 U17559 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n14157), .ZN(n14158) );
  NOR2_X1 U17560 ( .A1(n14159), .A2(n14158), .ZN(n14160) );
  INV_X1 U17561 ( .A(n14161), .ZN(n14162) );
  AOI22_X1 U17562 ( .A1(n19242), .A2(P2_REIP_REG_3__SCAN_IN), .B1(n19241), 
        .B2(n14162), .ZN(n14163) );
  OAI21_X1 U17563 ( .B1(n19203), .B2(n14164), .A(n14163), .ZN(n14167) );
  INV_X1 U17564 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14165) );
  NOR2_X2 U17565 ( .A1(n19242), .A2(n20136), .ZN(n19252) );
  AND2_X1 U17566 ( .A1(n20168), .A2(n16158), .ZN(n16482) );
  OAI22_X1 U17567 ( .A1(n14165), .A2(n19223), .B1(n19207), .B2(n20137), .ZN(
        n14166) );
  AOI211_X1 U17568 ( .C1(n19226), .C2(n13821), .A(n14167), .B(n14166), .ZN(
        n14168) );
  OAI211_X1 U17569 ( .C1(n19247), .C2(n20122), .A(n14169), .B(n14168), .ZN(
        P2_U2852) );
  OAI21_X1 U17570 ( .B1(n10354), .B2(n10379), .A(n14170), .ZN(n20217) );
  AOI22_X1 U17571 ( .A1(n14534), .A2(n14473), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n14532), .ZN(n14171) );
  OAI21_X1 U17572 ( .B1(n20217), .B2(n14536), .A(n14171), .ZN(P1_U2896) );
  INV_X1 U17573 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n14177) );
  AOI21_X1 U17574 ( .B1(n14172), .B2(n9855), .A(n14906), .ZN(n19093) );
  NAND2_X1 U17575 ( .A1(n19093), .A2(n19293), .ZN(n14176) );
  OAI211_X1 U17576 ( .C1(n9949), .C2(n13110), .A(n19278), .B(n14174), .ZN(
        n14175) );
  OAI211_X1 U17577 ( .C1(n19293), .C2(n14177), .A(n14176), .B(n14175), .ZN(
        P2_U2872) );
  XNOR2_X1 U17578 ( .A(n14178), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14179) );
  XNOR2_X1 U17579 ( .A(n14180), .B(n14179), .ZN(n16138) );
  NAND2_X1 U17580 ( .A1(n16138), .A2(n16034), .ZN(n14183) );
  NOR2_X1 U17581 ( .A1(n20369), .A2(n21019), .ZN(n16134) );
  NOR2_X1 U17582 ( .A1(n16031), .A2(n20214), .ZN(n14181) );
  AOI211_X1 U17583 ( .C1(n16027), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16134), .B(n14181), .ZN(n14182) );
  OAI211_X1 U17584 ( .C1(n14689), .C2(n20217), .A(n14183), .B(n14182), .ZN(
        P1_U2991) );
  AND2_X1 U17585 ( .A1(n14185), .A2(n14184), .ZN(n14186) );
  OR2_X1 U17586 ( .A1(n14195), .A2(n14186), .ZN(n20215) );
  OAI222_X1 U17587 ( .A1(n20215), .A2(n15973), .B1(n20306), .B2(n10036), .C1(
        n20217), .C2(n15974), .ZN(P1_U2864) );
  XNOR2_X1 U17588 ( .A(n14187), .B(n14188), .ZN(n15961) );
  AOI21_X1 U17589 ( .B1(n14189), .B2(n14197), .A(n9952), .ZN(n16123) );
  AOI22_X1 U17590 ( .A1(n16123), .A2(n13038), .B1(P1_EBX_REG_10__SCAN_IN), 
        .B2(n14433), .ZN(n14190) );
  OAI21_X1 U17591 ( .B1(n15961), .B2(n15974), .A(n14190), .ZN(P1_U2862) );
  AND2_X1 U17592 ( .A1(n14170), .A2(n14191), .ZN(n14192) );
  OR2_X1 U17593 ( .A1(n14192), .A2(n14187), .ZN(n20203) );
  AOI22_X1 U17594 ( .A1(n14534), .A2(n14470), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n14532), .ZN(n14193) );
  OAI21_X1 U17595 ( .B1(n20203), .B2(n14536), .A(n14193), .ZN(P1_U2895) );
  OR2_X1 U17596 ( .A1(n14195), .A2(n14194), .ZN(n14196) );
  AND2_X1 U17597 ( .A1(n14197), .A2(n14196), .ZN(n20208) );
  AOI22_X1 U17598 ( .A1(n20208), .A2(n13038), .B1(P1_EBX_REG_9__SCAN_IN), .B2(
        n14433), .ZN(n14198) );
  OAI21_X1 U17599 ( .B1(n20203), .B2(n15974), .A(n14198), .ZN(P1_U2863) );
  XNOR2_X1 U17600 ( .A(n14680), .B(n16126), .ZN(n14199) );
  XNOR2_X1 U17601 ( .A(n14200), .B(n14199), .ZN(n14211) );
  INV_X1 U17602 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16140) );
  NOR4_X1 U17603 ( .A1(n16141), .A2(n16140), .A3(n14202), .A4(n14201), .ZN(
        n14693) );
  NAND2_X1 U17604 ( .A1(n14693), .A2(n14203), .ZN(n16124) );
  AND2_X1 U17605 ( .A1(n14796), .A2(n16124), .ZN(n14204) );
  NOR2_X1 U17606 ( .A1(n14205), .A2(n14204), .ZN(n16133) );
  NOR2_X1 U17607 ( .A1(n20369), .A2(n21381), .ZN(n14213) );
  AOI21_X1 U17608 ( .B1(n20208), .B2(n16135), .A(n14213), .ZN(n14208) );
  INV_X1 U17609 ( .A(n16114), .ZN(n16125) );
  NOR2_X1 U17610 ( .A1(n16125), .A2(n16124), .ZN(n14206) );
  NAND2_X1 U17611 ( .A1(n14206), .A2(n16126), .ZN(n14207) );
  OAI211_X1 U17612 ( .C1(n16133), .C2(n16126), .A(n14208), .B(n14207), .ZN(
        n14209) );
  AOI21_X1 U17613 ( .B1(n14211), .B2(n20357), .A(n14209), .ZN(n14210) );
  INV_X1 U17614 ( .A(n14210), .ZN(P1_U3022) );
  NAND2_X1 U17615 ( .A1(n14211), .A2(n16034), .ZN(n14215) );
  NOR2_X1 U17616 ( .A1(n16031), .A2(n20206), .ZN(n14212) );
  AOI211_X1 U17617 ( .C1(n16027), .C2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n14213), .B(n14212), .ZN(n14214) );
  OAI211_X1 U17618 ( .C1(n14689), .C2(n20203), .A(n14215), .B(n14214), .ZN(
        P1_U2990) );
  INV_X1 U17619 ( .A(n14467), .ZN(n14216) );
  OAI222_X1 U17620 ( .A1(n14527), .A2(n14217), .B1(n14530), .B2(n14216), .C1(
        n14536), .C2(n15961), .ZN(P1_U2894) );
  INV_X1 U17621 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17250) );
  INV_X1 U17622 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n16933) );
  INV_X1 U17623 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17332) );
  NAND2_X1 U17624 ( .A1(n18366), .A2(n18351), .ZN(n14218) );
  INV_X1 U17625 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n14220) );
  NAND2_X1 U17626 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17350) );
  NOR2_X1 U17627 ( .A1(n14220), .A2(n17350), .ZN(n17340) );
  NAND3_X1 U17628 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n17340), .ZN(n17342) );
  NAND2_X1 U17629 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17337), .ZN(n17336) );
  INV_X1 U17630 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n14221) );
  NAND2_X1 U17631 ( .A1(n18366), .A2(n17247), .ZN(n17264) );
  NOR2_X1 U17632 ( .A1(n14221), .A2(n17264), .ZN(n15758) );
  AOI21_X1 U17633 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n15758), .A(
        P3_EBX_REG_14__SCAN_IN), .ZN(n14222) );
  NOR2_X1 U17634 ( .A1(n9951), .A2(n14222), .ZN(n14233) );
  AOI22_X1 U17635 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14232) );
  AOI22_X1 U17636 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14224) );
  AOI22_X1 U17637 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14223) );
  OAI211_X1 U17638 ( .C1(n17312), .C2(n18387), .A(n14224), .B(n14223), .ZN(
        n14230) );
  AOI22_X1 U17639 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9812), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14228) );
  AOI22_X1 U17640 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17309), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14227) );
  AOI22_X1 U17641 ( .A1(n17310), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14226) );
  NAND4_X1 U17642 ( .A1(n14228), .A2(n14227), .A3(n14226), .A4(n14225), .ZN(
        n14229) );
  AOI211_X1 U17643 ( .C1(n17293), .C2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n14230), .B(n14229), .ZN(n14231) );
  OAI211_X1 U17644 ( .C1(n9890), .C2(n17108), .A(n14232), .B(n14231), .ZN(
        n17454) );
  MUX2_X1 U17645 ( .A(n14233), .B(n17454), .S(n17361), .Z(P3_U2689) );
  NAND2_X1 U17646 ( .A1(n14235), .A2(n14234), .ZN(n15110) );
  INV_X1 U17647 ( .A(n14236), .ZN(n14238) );
  NAND2_X1 U17648 ( .A1(n14238), .A2(n14237), .ZN(n14243) );
  NAND2_X1 U17649 ( .A1(n19470), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14239) );
  XNOR2_X1 U17650 ( .A(n14243), .B(n14239), .ZN(n16167) );
  AOI21_X1 U17651 ( .B1(n16167), .B2(n14246), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15111) );
  INV_X1 U17652 ( .A(n16167), .ZN(n14240) );
  NOR2_X1 U17653 ( .A1(n14243), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14244) );
  MUX2_X1 U17654 ( .A(n14245), .B(n14244), .S(n19470), .Z(n16157) );
  NAND2_X1 U17655 ( .A1(n16157), .A2(n14246), .ZN(n14247) );
  XNOR2_X1 U17656 ( .A(n14247), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14248) );
  XNOR2_X1 U17657 ( .A(n14249), .B(n14248), .ZN(n14281) );
  AOI22_X1 U17658 ( .A1(n14254), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n14252) );
  NAND2_X1 U17659 ( .A1(n14250), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14251) );
  OAI211_X1 U17660 ( .C1(n14253), .C2(n20107), .A(n14252), .B(n14251), .ZN(
        n14946) );
  AOI22_X1 U17661 ( .A1(n14254), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n14257) );
  NAND2_X1 U17662 ( .A1(n14255), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14256) );
  OAI211_X1 U17663 ( .C1(n14259), .C2(n14258), .A(n14257), .B(n14256), .ZN(
        n14260) );
  INV_X1 U17664 ( .A(n14277), .ZN(n14261) );
  NAND2_X1 U17665 ( .A1(n14261), .A2(n16390), .ZN(n14272) );
  NAND2_X1 U17666 ( .A1(n14262), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14266) );
  AND2_X1 U17667 ( .A1(n16420), .A2(n14266), .ZN(n14263) );
  NOR2_X1 U17668 ( .A1(n15348), .A2(n14263), .ZN(n15326) );
  OAI21_X1 U17669 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16386), .A(
        n15326), .ZN(n14270) );
  AOI222_X1 U17670 ( .A1(n11409), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n11406), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n11416), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14264) );
  NAND2_X1 U17671 ( .A1(n19414), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14275) );
  OAI21_X1 U17672 ( .B1(n16164), .B2(n16412), .A(n14275), .ZN(n14269) );
  INV_X1 U17673 ( .A(n14266), .ZN(n14267) );
  NAND2_X1 U17674 ( .A1(n15336), .A2(n14267), .ZN(n15319) );
  NOR3_X1 U17675 ( .A1(n15319), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15325), .ZN(n14268) );
  AOI211_X1 U17676 ( .C1(n14270), .C2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n14269), .B(n14268), .ZN(n14271) );
  OAI21_X1 U17677 ( .B1(n14281), .B2(n16425), .A(n14273), .ZN(P2_U3015) );
  NAND2_X1 U17678 ( .A1(n16316), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14274) );
  OAI211_X1 U17679 ( .C1(n16355), .C2(n14276), .A(n14275), .B(n14274), .ZN(
        n14279) );
  NOR2_X1 U17680 ( .A1(n14277), .A2(n16371), .ZN(n14278) );
  OAI21_X1 U17681 ( .B1(n14281), .B2(n19417), .A(n14280), .ZN(P2_U2983) );
  AOI21_X1 U17682 ( .B1(n14298), .B2(P1_REIP_REG_29__SCAN_IN), .A(
        P1_REIP_REG_30__SCAN_IN), .ZN(n14287) );
  NAND2_X1 U17683 ( .A1(n14563), .A2(n20245), .ZN(n14286) );
  NAND2_X1 U17684 ( .A1(n20292), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n14283) );
  NAND2_X1 U17685 ( .A1(n20255), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14282) );
  OAI211_X1 U17686 ( .C1(n14561), .C2(n20289), .A(n14283), .B(n14282), .ZN(
        n14284) );
  AOI21_X1 U17687 ( .B1(n14727), .B2(n20272), .A(n14284), .ZN(n14285) );
  OAI211_X1 U17688 ( .C1(n14288), .C2(n14287), .A(n14286), .B(n14285), .ZN(
        P1_U2810) );
  OAI21_X1 U17689 ( .B1(n14289), .B2(n14291), .A(n14290), .ZN(n14570) );
  INV_X1 U17690 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21408) );
  OAI21_X1 U17691 ( .B1(n14303), .B2(n14293), .A(n14292), .ZN(n14731) );
  AOI22_X1 U17692 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n20255), .B1(
        n20254), .B2(n14567), .ZN(n14294) );
  OAI21_X1 U17693 ( .B1(n20218), .B2(n21410), .A(n14294), .ZN(n14295) );
  AOI21_X1 U17694 ( .B1(n14304), .B2(P1_REIP_REG_29__SCAN_IN), .A(n14295), 
        .ZN(n14296) );
  OAI21_X1 U17695 ( .B1(n14731), .B2(n20295), .A(n14296), .ZN(n14297) );
  AOI21_X1 U17696 ( .B1(n14298), .B2(n21408), .A(n14297), .ZN(n14299) );
  OAI21_X1 U17697 ( .B1(n14570), .B2(n15960), .A(n14299), .ZN(P1_U2811) );
  AOI21_X1 U17698 ( .B1(n14300), .B2(n12628), .A(n14289), .ZN(n14582) );
  INV_X1 U17699 ( .A(n14582), .ZN(n14464) );
  NOR2_X1 U17700 ( .A1(n14313), .A2(n14301), .ZN(n14302) );
  OR2_X1 U17701 ( .A1(n14303), .A2(n14302), .ZN(n14744) );
  INV_X1 U17702 ( .A(n14744), .ZN(n14310) );
  NAND2_X1 U17703 ( .A1(n14304), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14307) );
  INV_X1 U17704 ( .A(n14580), .ZN(n14305) );
  AOI22_X1 U17705 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n20255), .B1(
        n20254), .B2(n14305), .ZN(n14306) );
  OAI211_X1 U17706 ( .C1(n21315), .C2(n20218), .A(n14307), .B(n14306), .ZN(
        n14309) );
  NOR3_X1 U17707 ( .A1(n14319), .A2(P1_REIP_REG_28__SCAN_IN), .A3(n21412), 
        .ZN(n14308) );
  AOI211_X1 U17708 ( .C1(n14310), .C2(n20272), .A(n14309), .B(n14308), .ZN(
        n14311) );
  OAI21_X1 U17709 ( .B1(n14464), .B2(n15960), .A(n14311), .ZN(P1_U2812) );
  NAND2_X1 U17710 ( .A1(n14327), .A2(n14314), .ZN(n14315) );
  NAND2_X1 U17711 ( .A1(n10162), .A2(n14315), .ZN(n14419) );
  INV_X1 U17712 ( .A(n14419), .ZN(n14753) );
  AOI22_X1 U17713 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n20255), .B1(
        n20254), .B2(n14316), .ZN(n14318) );
  NAND2_X1 U17714 ( .A1(n20292), .A2(P1_EBX_REG_27__SCAN_IN), .ZN(n14317) );
  OAI211_X1 U17715 ( .C1(n14333), .C2(n21412), .A(n14318), .B(n14317), .ZN(
        n14321) );
  NOR2_X1 U17716 ( .A1(n14319), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14320) );
  AOI211_X1 U17717 ( .C1(n14753), .C2(n20272), .A(n14321), .B(n14320), .ZN(
        n14322) );
  OAI21_X1 U17718 ( .B1(n14312), .B2(n15960), .A(n14322), .ZN(P1_U2813) );
  AOI21_X1 U17719 ( .B1(n14324), .B2(n14323), .A(n12627), .ZN(n14325) );
  INV_X1 U17720 ( .A(n14325), .ZN(n14591) );
  INV_X1 U17721 ( .A(n14351), .ZN(n14340) );
  AOI21_X1 U17722 ( .B1(n14340), .B2(n14339), .A(n14326), .ZN(n14329) );
  INV_X1 U17723 ( .A(n14327), .ZN(n14328) );
  NOR2_X1 U17724 ( .A1(n14329), .A2(n14328), .ZN(n14757) );
  INV_X1 U17725 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n21037) );
  OAI22_X1 U17726 ( .A1(n14330), .A2(n20288), .B1(n20289), .B2(n14588), .ZN(
        n14331) );
  AOI21_X1 U17727 ( .B1(n20292), .B2(P1_EBX_REG_26__SCAN_IN), .A(n14331), .ZN(
        n14332) );
  OAI21_X1 U17728 ( .B1(n14333), .B2(n21037), .A(n14332), .ZN(n14334) );
  AOI21_X1 U17729 ( .B1(n14757), .B2(n20272), .A(n14334), .ZN(n14336) );
  NAND4_X1 U17730 ( .A1(n14357), .A2(P1_REIP_REG_25__SCAN_IN), .A3(
        P1_REIP_REG_24__SCAN_IN), .A4(n21037), .ZN(n14335) );
  OAI211_X1 U17731 ( .C1(n14591), .C2(n15960), .A(n14336), .B(n14335), .ZN(
        P1_U2814) );
  XNOR2_X1 U17732 ( .A(n14337), .B(n14338), .ZN(n14600) );
  XOR2_X1 U17733 ( .A(P1_REIP_REG_25__SCAN_IN), .B(P1_REIP_REG_24__SCAN_IN), 
        .Z(n14345) );
  XNOR2_X1 U17734 ( .A(n14340), .B(n14339), .ZN(n16042) );
  INV_X1 U17735 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n21325) );
  AOI22_X1 U17736 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n20255), .B1(
        n20254), .B2(n14599), .ZN(n14341) );
  OAI21_X1 U17737 ( .B1(n20218), .B2(n21325), .A(n14341), .ZN(n14342) );
  AOI21_X1 U17738 ( .B1(n14368), .B2(P1_REIP_REG_25__SCAN_IN), .A(n14342), 
        .ZN(n14343) );
  OAI21_X1 U17739 ( .B1(n16042), .B2(n20295), .A(n14343), .ZN(n14344) );
  AOI21_X1 U17740 ( .B1(n14357), .B2(n14345), .A(n14344), .ZN(n14346) );
  OAI21_X1 U17741 ( .B1(n14600), .B2(n15960), .A(n14346), .ZN(P1_U2815) );
  AOI21_X1 U17742 ( .B1(n14348), .B2(n14347), .A(n14337), .ZN(n14606) );
  INV_X1 U17743 ( .A(n14606), .ZN(n14476) );
  INV_X1 U17744 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21413) );
  OR2_X1 U17745 ( .A1(n14362), .A2(n14349), .ZN(n14350) );
  NAND2_X1 U17746 ( .A1(n14351), .A2(n14350), .ZN(n16049) );
  OAI22_X1 U17747 ( .A1(n14352), .A2(n20288), .B1(n20289), .B2(n14604), .ZN(
        n14354) );
  NOR2_X1 U17748 ( .A1(n20218), .A2(n21363), .ZN(n14353) );
  AOI211_X1 U17749 ( .C1(n14368), .C2(P1_REIP_REG_24__SCAN_IN), .A(n14354), 
        .B(n14353), .ZN(n14355) );
  OAI21_X1 U17750 ( .B1(n16049), .B2(n20295), .A(n14355), .ZN(n14356) );
  AOI21_X1 U17751 ( .B1(n14357), .B2(n21413), .A(n14356), .ZN(n14358) );
  OAI21_X1 U17752 ( .B1(n14476), .B2(n15960), .A(n14358), .ZN(P1_U2816) );
  AND2_X1 U17753 ( .A1(n14359), .A2(n14372), .ZN(n14361) );
  OAI21_X1 U17754 ( .B1(n14361), .B2(n14360), .A(n14347), .ZN(n14616) );
  INV_X1 U17755 ( .A(n14362), .ZN(n14363) );
  OAI21_X1 U17756 ( .B1(n14376), .B2(n14364), .A(n14363), .ZN(n14421) );
  INV_X1 U17757 ( .A(n14421), .ZN(n14768) );
  AOI22_X1 U17758 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n20255), .B1(
        n20254), .B2(n14619), .ZN(n14365) );
  OAI21_X1 U17759 ( .B1(n20218), .B2(n21195), .A(n14365), .ZN(n14366) );
  AOI21_X1 U17760 ( .B1(n14768), .B2(n20272), .A(n14366), .ZN(n14371) );
  INV_X1 U17761 ( .A(n15893), .ZN(n15877) );
  NAND3_X1 U17762 ( .A1(n15877), .A2(P1_REIP_REG_21__SCAN_IN), .A3(n14367), 
        .ZN(n14383) );
  INV_X1 U17763 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21309) );
  NOR2_X1 U17764 ( .A1(n14383), .A2(n21309), .ZN(n14369) );
  OAI21_X1 U17765 ( .B1(n14369), .B2(P1_REIP_REG_23__SCAN_IN), .A(n14368), 
        .ZN(n14370) );
  OAI211_X1 U17766 ( .C1(n14616), .C2(n15960), .A(n14371), .B(n14370), .ZN(
        P1_U2817) );
  XOR2_X1 U17767 ( .A(n14372), .B(n14359), .Z(n14624) );
  NAND2_X1 U17768 ( .A1(n14624), .A2(n20245), .ZN(n14382) );
  OR3_X1 U17769 ( .A1(n15893), .A2(n14373), .A3(P1_REIP_REG_21__SCAN_IN), .ZN(
        n14392) );
  AOI21_X1 U17770 ( .B1(n15875), .B2(n14392), .A(n21309), .ZN(n14380) );
  NOR2_X1 U17771 ( .A1(n9921), .A2(n14374), .ZN(n14375) );
  OR2_X1 U17772 ( .A1(n14376), .A2(n14375), .ZN(n16060) );
  INV_X1 U17773 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14422) );
  OAI22_X1 U17774 ( .A1(n16060), .A2(n20295), .B1(n20218), .B2(n14422), .ZN(
        n14377) );
  INV_X1 U17775 ( .A(n14377), .ZN(n14378) );
  OAI21_X1 U17776 ( .B1(n14625), .B2(n20289), .A(n14378), .ZN(n14379) );
  AOI211_X1 U17777 ( .C1(n20255), .C2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n14380), .B(n14379), .ZN(n14381) );
  OAI211_X1 U17778 ( .C1(P1_REIP_REG_22__SCAN_IN), .C2(n14383), .A(n14382), 
        .B(n14381), .ZN(P1_U2818) );
  INV_X1 U17779 ( .A(n14359), .ZN(n14385) );
  OAI21_X1 U17780 ( .B1(n14386), .B2(n14384), .A(n14385), .ZN(n14634) );
  AND2_X1 U17781 ( .A1(n15853), .A2(n14387), .ZN(n14388) );
  NOR2_X1 U17782 ( .A1(n9921), .A2(n14388), .ZN(n14423) );
  INV_X1 U17783 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n21369) );
  NOR2_X1 U17784 ( .A1(n15875), .A2(n21369), .ZN(n14391) );
  INV_X1 U17785 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n21415) );
  AOI22_X1 U17786 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n20255), .B1(
        n20254), .B2(n14637), .ZN(n14389) );
  OAI21_X1 U17787 ( .B1(n20218), .B2(n21415), .A(n14389), .ZN(n14390) );
  AOI211_X1 U17788 ( .C1(n14423), .C2(n20272), .A(n14391), .B(n14390), .ZN(
        n14393) );
  OAI211_X1 U17789 ( .C1(n14634), .C2(n15960), .A(n14393), .B(n14392), .ZN(
        P1_U2819) );
  OAI21_X1 U17790 ( .B1(n14394), .B2(n14396), .A(n14395), .ZN(n14662) );
  AND2_X1 U17791 ( .A1(n20250), .A2(n14397), .ZN(n15887) );
  OAI21_X1 U17792 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n14398), .A(n15887), 
        .ZN(n14407) );
  INV_X1 U17793 ( .A(n14653), .ZN(n14399) );
  NAND2_X1 U17794 ( .A1(n20254), .A2(n14399), .ZN(n14401) );
  NAND2_X1 U17795 ( .A1(n14408), .A2(n14400), .ZN(n20256) );
  OAI211_X1 U17796 ( .C1(n20288), .C2(n14402), .A(n14401), .B(n20256), .ZN(
        n14405) );
  OAI21_X1 U17797 ( .B1(n9958), .B2(n14403), .A(n14801), .ZN(n14432) );
  NOR2_X1 U17798 ( .A1(n14432), .A2(n20295), .ZN(n14404) );
  AOI211_X1 U17799 ( .C1(n20292), .C2(P1_EBX_REG_17__SCAN_IN), .A(n14405), .B(
        n14404), .ZN(n14406) );
  OAI211_X1 U17800 ( .C1(n14662), .C2(n15960), .A(n14407), .B(n14406), .ZN(
        P1_U2823) );
  OAI22_X1 U17801 ( .A1(n20289), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n21391), .B2(n14408), .ZN(n14411) );
  OAI22_X1 U17802 ( .A1(n20218), .A2(n14409), .B1(P1_REIP_REG_1__SCAN_IN), 
        .B2(n20276), .ZN(n14410) );
  AOI211_X1 U17803 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n20255), .A(
        n14411), .B(n14410), .ZN(n14412) );
  OAI21_X1 U17804 ( .B1(n20295), .B2(n14413), .A(n14412), .ZN(n14414) );
  AOI21_X1 U17805 ( .B1(n20881), .B2(n20286), .A(n14414), .ZN(n14415) );
  OAI21_X1 U17806 ( .B1(n14417), .B2(n14416), .A(n14415), .ZN(P1_U2839) );
  OAI22_X1 U17807 ( .A1(n14702), .A2(n15973), .B1(n20306), .B2(n21300), .ZN(
        P1_U2841) );
  OAI222_X1 U17808 ( .A1(n14731), .A2(n15973), .B1(n21410), .B2(n20306), .C1(
        n14570), .C2(n15974), .ZN(P1_U2843) );
  OAI222_X1 U17809 ( .A1(n14464), .A2(n15974), .B1(n21315), .B2(n20306), .C1(
        n14744), .C2(n15973), .ZN(P1_U2844) );
  OAI222_X1 U17810 ( .A1(n14312), .A2(n15974), .B1(n21313), .B2(n20306), .C1(
        n14419), .C2(n15973), .ZN(P1_U2845) );
  AOI22_X1 U17811 ( .A1(n14757), .A2(n13038), .B1(P1_EBX_REG_26__SCAN_IN), 
        .B2(n14433), .ZN(n14420) );
  OAI21_X1 U17812 ( .B1(n14591), .B2(n15974), .A(n14420), .ZN(P1_U2846) );
  OAI222_X1 U17813 ( .A1(n15974), .A2(n14600), .B1(n21325), .B2(n20306), .C1(
        n15973), .C2(n16042), .ZN(P1_U2847) );
  OAI222_X1 U17814 ( .A1(n14476), .A2(n15974), .B1(n21363), .B2(n20306), .C1(
        n16049), .C2(n15973), .ZN(P1_U2848) );
  OAI222_X1 U17815 ( .A1(n14616), .A2(n15974), .B1(n21195), .B2(n20306), .C1(
        n14421), .C2(n15973), .ZN(P1_U2849) );
  INV_X1 U17816 ( .A(n14624), .ZN(n14483) );
  OAI222_X1 U17817 ( .A1(n16060), .A2(n15973), .B1(n14422), .B2(n20306), .C1(
        n14483), .C2(n15974), .ZN(P1_U2850) );
  INV_X1 U17818 ( .A(n14423), .ZN(n14784) );
  OAI222_X1 U17819 ( .A1(n14784), .A2(n15973), .B1(n20306), .B2(n21415), .C1(
        n14634), .C2(n15974), .ZN(P1_U2851) );
  NAND2_X1 U17820 ( .A1(n14800), .A2(n14425), .ZN(n14426) );
  NAND2_X1 U17821 ( .A1(n15855), .A2(n14426), .ZN(n15879) );
  BUF_X1 U17822 ( .A(n14429), .Z(n14430) );
  OAI21_X1 U17823 ( .B1(n14428), .B2(n14431), .A(n14430), .ZN(n15880) );
  OAI222_X1 U17824 ( .A1(n15879), .A2(n15973), .B1(n20306), .B2(n10028), .C1(
        n15880), .C2(n15974), .ZN(P1_U2853) );
  INV_X1 U17825 ( .A(n14432), .ZN(n14816) );
  AOI22_X1 U17826 ( .A1(n14816), .A2(n13038), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n14433), .ZN(n14434) );
  OAI21_X1 U17827 ( .B1(n14662), .B2(n15974), .A(n14434), .ZN(P1_U2855) );
  INV_X1 U17828 ( .A(n14436), .ZN(n14514) );
  OAI21_X1 U17829 ( .B1(n14514), .B2(n12359), .A(n14438), .ZN(n15910) );
  INV_X1 U17830 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14439) );
  INV_X1 U17831 ( .A(n15919), .ZN(n15898) );
  XNOR2_X1 U17832 ( .A(n15898), .B(n15897), .ZN(n15906) );
  OAI222_X1 U17833 ( .A1(n15974), .A2(n15910), .B1(n14439), .B2(n20306), .C1(
        n15973), .C2(n15906), .ZN(P1_U2857) );
  AND2_X1 U17834 ( .A1(n14440), .A2(n14441), .ZN(n14443) );
  OR2_X1 U17835 ( .A1(n14443), .A2(n14442), .ZN(n14521) );
  NOR2_X1 U17836 ( .A1(n15938), .A2(n14444), .ZN(n14445) );
  OR2_X1 U17837 ( .A1(n15917), .A2(n14445), .ZN(n16092) );
  OAI22_X1 U17838 ( .A1(n16092), .A2(n15973), .B1(n21299), .B2(n20306), .ZN(
        n14446) );
  AOI21_X1 U17839 ( .B1(n15932), .B2(n20303), .A(n14446), .ZN(n14447) );
  INV_X1 U17840 ( .A(n14447), .ZN(P1_U2859) );
  OAI21_X1 U17841 ( .B1(n9952), .B2(n9981), .A(n15936), .ZN(n16116) );
  INV_X1 U17842 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n21318) );
  NAND2_X1 U17843 ( .A1(n14449), .A2(n14448), .ZN(n14452) );
  INV_X1 U17844 ( .A(n14450), .ZN(n14451) );
  AOI21_X1 U17845 ( .B1(n14453), .B2(n14452), .A(n14451), .ZN(n16023) );
  INV_X1 U17846 ( .A(n16023), .ZN(n14537) );
  OAI222_X1 U17847 ( .A1(n16116), .A2(n15973), .B1(n20306), .B2(n21318), .C1(
        n14537), .C2(n15974), .ZN(P1_U2861) );
  AOI22_X1 U17848 ( .A1(n14505), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n14532), .ZN(n14458) );
  NOR3_X1 U17849 ( .A1(n14532), .A2(n14455), .A3(n11926), .ZN(n14456) );
  AOI22_X1 U17850 ( .A1(n14508), .A2(n14516), .B1(n14506), .B2(DATAI_30_), 
        .ZN(n14457) );
  OAI211_X1 U17851 ( .C1(n14459), .C2(n14536), .A(n14458), .B(n14457), .ZN(
        P1_U2874) );
  AOI22_X1 U17852 ( .A1(n14505), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n14532), .ZN(n14461) );
  AOI22_X1 U17853 ( .A1(n14508), .A2(n14519), .B1(n14506), .B2(DATAI_29_), 
        .ZN(n14460) );
  OAI211_X1 U17854 ( .C1(n14570), .C2(n14536), .A(n14461), .B(n14460), .ZN(
        P1_U2875) );
  AOI22_X1 U17855 ( .A1(n14505), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n14532), .ZN(n14463) );
  AOI22_X1 U17856 ( .A1(n14508), .A2(n14526), .B1(n14506), .B2(DATAI_28_), 
        .ZN(n14462) );
  OAI211_X1 U17857 ( .C1(n14464), .C2(n14536), .A(n14463), .B(n14462), .ZN(
        P1_U2876) );
  AOI22_X1 U17858 ( .A1(n14505), .A2(BUF1_REG_27__SCAN_IN), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(n14532), .ZN(n14466) );
  AOI22_X1 U17859 ( .A1(n14508), .A2(n14533), .B1(n14506), .B2(DATAI_27_), 
        .ZN(n14465) );
  OAI211_X1 U17860 ( .C1(n14312), .C2(n14536), .A(n14466), .B(n14465), .ZN(
        P1_U2877) );
  AOI22_X1 U17861 ( .A1(n14505), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n14532), .ZN(n14469) );
  AOI22_X1 U17862 ( .A1(n14508), .A2(n14467), .B1(n14506), .B2(DATAI_26_), 
        .ZN(n14468) );
  OAI211_X1 U17863 ( .C1(n14591), .C2(n14536), .A(n14469), .B(n14468), .ZN(
        P1_U2878) );
  AOI22_X1 U17864 ( .A1(n14505), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n14532), .ZN(n14472) );
  AOI22_X1 U17865 ( .A1(n14508), .A2(n14470), .B1(n14506), .B2(DATAI_25_), 
        .ZN(n14471) );
  OAI211_X1 U17866 ( .C1(n14600), .C2(n14536), .A(n14472), .B(n14471), .ZN(
        P1_U2879) );
  AOI22_X1 U17867 ( .A1(n14505), .A2(BUF1_REG_24__SCAN_IN), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(n14532), .ZN(n14475) );
  AOI22_X1 U17868 ( .A1(n14508), .A2(n14473), .B1(n14506), .B2(DATAI_24_), 
        .ZN(n14474) );
  OAI211_X1 U17869 ( .C1(n14476), .C2(n14536), .A(n14475), .B(n14474), .ZN(
        P1_U2880) );
  AOI22_X1 U17870 ( .A1(n14505), .A2(BUF1_REG_23__SCAN_IN), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(n14532), .ZN(n14479) );
  AOI22_X1 U17871 ( .A1(n14508), .A2(n14477), .B1(n14506), .B2(DATAI_23_), 
        .ZN(n14478) );
  OAI211_X1 U17872 ( .C1(n14616), .C2(n14536), .A(n14479), .B(n14478), .ZN(
        P1_U2881) );
  AOI22_X1 U17873 ( .A1(n14505), .A2(BUF1_REG_22__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n14532), .ZN(n14482) );
  AOI22_X1 U17874 ( .A1(n14508), .A2(n14480), .B1(n14506), .B2(DATAI_22_), 
        .ZN(n14481) );
  OAI211_X1 U17875 ( .C1(n14483), .C2(n14536), .A(n14482), .B(n14481), .ZN(
        P1_U2882) );
  AOI22_X1 U17876 ( .A1(n14505), .A2(BUF1_REG_21__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n14532), .ZN(n14486) );
  AOI22_X1 U17877 ( .A1(n14508), .A2(n14484), .B1(n14506), .B2(DATAI_21_), 
        .ZN(n14485) );
  OAI211_X1 U17878 ( .C1(n14634), .C2(n14536), .A(n14486), .B(n14485), .ZN(
        P1_U2883) );
  AOI21_X1 U17879 ( .B1(n14487), .B2(n14430), .A(n14384), .ZN(n15981) );
  INV_X1 U17880 ( .A(n15981), .ZN(n14491) );
  AOI22_X1 U17881 ( .A1(n14505), .A2(BUF1_REG_20__SCAN_IN), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(n14532), .ZN(n14490) );
  AOI22_X1 U17882 ( .A1(n14508), .A2(n14488), .B1(n14506), .B2(DATAI_20_), 
        .ZN(n14489) );
  OAI211_X1 U17883 ( .C1(n14491), .C2(n14536), .A(n14490), .B(n14489), .ZN(
        P1_U2884) );
  AOI22_X1 U17884 ( .A1(n14505), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n14532), .ZN(n14494) );
  AOI22_X1 U17885 ( .A1(n14508), .A2(n14492), .B1(n14506), .B2(DATAI_19_), 
        .ZN(n14493) );
  OAI211_X1 U17886 ( .C1(n15880), .C2(n14536), .A(n14494), .B(n14493), .ZN(
        P1_U2885) );
  AOI21_X1 U17887 ( .B1(n14495), .B2(n14395), .A(n14428), .ZN(n15970) );
  INV_X1 U17888 ( .A(n15970), .ZN(n14499) );
  AOI22_X1 U17889 ( .A1(n14505), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n14532), .ZN(n14498) );
  AOI22_X1 U17890 ( .A1(n14508), .A2(n14496), .B1(n14506), .B2(DATAI_18_), 
        .ZN(n14497) );
  OAI211_X1 U17891 ( .C1(n14499), .C2(n14536), .A(n14498), .B(n14497), .ZN(
        P1_U2886) );
  AOI22_X1 U17892 ( .A1(n14505), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n14532), .ZN(n14502) );
  AOI22_X1 U17893 ( .A1(n14508), .A2(n14500), .B1(n14506), .B2(DATAI_17_), 
        .ZN(n14501) );
  OAI211_X1 U17894 ( .C1(n14662), .C2(n14536), .A(n14502), .B(n14501), .ZN(
        P1_U2887) );
  AND2_X1 U17895 ( .A1(n14438), .A2(n14503), .ZN(n14504) );
  OR2_X1 U17896 ( .A1(n14394), .A2(n14504), .ZN(n15985) );
  AOI22_X1 U17897 ( .A1(n14505), .A2(BUF1_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n14532), .ZN(n14510) );
  AOI22_X1 U17898 ( .A1(n14508), .A2(n14507), .B1(n14506), .B2(DATAI_16_), 
        .ZN(n14509) );
  OAI211_X1 U17899 ( .C1(n15985), .C2(n14536), .A(n14510), .B(n14509), .ZN(
        P1_U2888) );
  OAI222_X1 U17900 ( .A1(n15910), .A2(n14536), .B1(n14530), .B2(n14512), .C1(
        n14527), .C2(n14511), .ZN(P1_U2889) );
  INV_X1 U17901 ( .A(n14442), .ZN(n14515) );
  INV_X1 U17902 ( .A(n16004), .ZN(n14518) );
  AOI22_X1 U17903 ( .A1(n14534), .A2(n14516), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n14532), .ZN(n14517) );
  OAI21_X1 U17904 ( .B1(n14518), .B2(n14536), .A(n14517), .ZN(P1_U2890) );
  AOI22_X1 U17905 ( .A1(n14534), .A2(n14519), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n14532), .ZN(n14520) );
  OAI21_X1 U17906 ( .B1(n14521), .B2(n14536), .A(n14520), .ZN(P1_U2891) );
  INV_X1 U17907 ( .A(n14522), .ZN(n14524) );
  NAND2_X1 U17908 ( .A1(n14524), .A2(n10351), .ZN(n14525) );
  AND2_X1 U17909 ( .A1(n14440), .A2(n14525), .ZN(n16015) );
  INV_X1 U17910 ( .A(n16015), .ZN(n14531) );
  INV_X1 U17911 ( .A(n14526), .ZN(n14529) );
  OAI222_X1 U17912 ( .A1(n14531), .A2(n14536), .B1(n14530), .B2(n14529), .C1(
        n14528), .C2(n14527), .ZN(P1_U2892) );
  AOI22_X1 U17913 ( .A1(n14534), .A2(n14533), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n14532), .ZN(n14535) );
  OAI21_X1 U17914 ( .B1(n14537), .B2(n14536), .A(n14535), .ZN(P1_U2893) );
  INV_X1 U17915 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14538) );
  NAND2_X1 U17916 ( .A1(n14573), .A2(n14538), .ZN(n14739) );
  NAND2_X1 U17917 ( .A1(n14555), .A2(n16018), .ZN(n14540) );
  AND2_X1 U17918 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14698) );
  NAND2_X1 U17919 ( .A1(n14539), .A2(n14698), .ZN(n14556) );
  NAND2_X1 U17920 ( .A1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14544) );
  NOR2_X1 U17921 ( .A1(n14544), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14700) );
  MUX2_X1 U17922 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n14700), .S(
        n14680), .Z(n14543) );
  INV_X1 U17923 ( .A(n14543), .ZN(n14547) );
  INV_X1 U17924 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14737) );
  INV_X1 U17925 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14541) );
  NAND2_X1 U17926 ( .A1(n14737), .A2(n14541), .ZN(n14542) );
  OAI21_X1 U17927 ( .B1(n14556), .B2(n14544), .A(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14545) );
  INV_X1 U17928 ( .A(n14549), .ZN(n14551) );
  NOR2_X1 U17929 ( .A1(n20369), .A2(n21048), .ZN(n14699) );
  AOI21_X1 U17930 ( .B1(n16027), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14699), .ZN(n14550) );
  OAI21_X1 U17931 ( .B1(n14551), .B2(n16031), .A(n14550), .ZN(n14552) );
  AOI21_X1 U17932 ( .B1(n14690), .B2(n16034), .A(n14552), .ZN(n14553) );
  OAI21_X1 U17933 ( .B1(n14554), .B2(n14689), .A(n14553), .ZN(P1_U2968) );
  NOR2_X1 U17934 ( .A1(n14555), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14558) );
  NOR2_X1 U17935 ( .A1(n14556), .A2(n14737), .ZN(n14557) );
  MUX2_X1 U17936 ( .A(n14558), .B(n14557), .S(n14680), .Z(n14559) );
  XNOR2_X1 U17937 ( .A(n14559), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14729) );
  NAND2_X1 U17938 ( .A1(n16106), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14723) );
  NAND2_X1 U17939 ( .A1(n16027), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14560) );
  OAI211_X1 U17940 ( .C1(n16031), .C2(n14561), .A(n14723), .B(n14560), .ZN(
        n14562) );
  AOI21_X1 U17941 ( .B1(n14563), .B2(n20374), .A(n14562), .ZN(n14564) );
  OAI21_X1 U17942 ( .B1(n20187), .B2(n14729), .A(n14564), .ZN(P1_U2969) );
  NOR2_X1 U17943 ( .A1(n20369), .A2(n21408), .ZN(n14733) );
  NOR2_X1 U17944 ( .A1(n16038), .A2(n14565), .ZN(n14566) );
  AOI211_X1 U17945 ( .C1(n16033), .C2(n14567), .A(n14733), .B(n14566), .ZN(
        n14569) );
  NAND2_X1 U17946 ( .A1(n14730), .A2(n16034), .ZN(n14568) );
  OAI211_X1 U17947 ( .C1(n14570), .C2(n14689), .A(n14569), .B(n14568), .ZN(
        P1_U2970) );
  NAND2_X1 U17948 ( .A1(n14612), .A2(n14571), .ZN(n14575) );
  AND3_X1 U17949 ( .A1(n14575), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14577) );
  INV_X1 U17950 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14572) );
  NAND3_X1 U17951 ( .A1(n14585), .A2(n14573), .A3(n14572), .ZN(n14574) );
  NOR2_X1 U17952 ( .A1(n14575), .A2(n14574), .ZN(n14576) );
  MUX2_X1 U17953 ( .A(n14577), .B(n14576), .S(n16018), .Z(n14578) );
  XNOR2_X1 U17954 ( .A(n14578), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14748) );
  OR2_X1 U17955 ( .A1(n20369), .A2(n21310), .ZN(n14743) );
  NAND2_X1 U17956 ( .A1(n16027), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14579) );
  OAI211_X1 U17957 ( .C1(n16031), .C2(n14580), .A(n14743), .B(n14579), .ZN(
        n14581) );
  AOI21_X1 U17958 ( .B1(n14582), .B2(n20374), .A(n14581), .ZN(n14583) );
  OAI21_X1 U17959 ( .B1(n20187), .B2(n14748), .A(n14583), .ZN(P1_U2971) );
  NOR2_X1 U17960 ( .A1(n10144), .A2(n14680), .ZN(n14609) );
  NOR3_X1 U17961 ( .A1(n14608), .A2(n16018), .A3(n14714), .ZN(n14584) );
  AOI21_X1 U17962 ( .B1(n14609), .B2(n14585), .A(n14584), .ZN(n14586) );
  XNOR2_X1 U17963 ( .A(n14586), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14756) );
  NOR2_X1 U17964 ( .A1(n20369), .A2(n21037), .ZN(n14760) );
  AOI21_X1 U17965 ( .B1(n16027), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n14760), .ZN(n14587) );
  OAI21_X1 U17966 ( .B1(n14588), .B2(n16031), .A(n14587), .ZN(n14589) );
  AOI21_X1 U17967 ( .B1(n14756), .B2(n16034), .A(n14589), .ZN(n14590) );
  OAI21_X1 U17968 ( .B1(n14591), .B2(n14689), .A(n14590), .ZN(P1_U2973) );
  INV_X1 U17969 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n14592) );
  OAI22_X1 U17970 ( .A1(n16038), .A2(n14593), .B1(n20369), .B2(n14592), .ZN(
        n14598) );
  NAND2_X1 U17971 ( .A1(n14594), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14601) );
  NAND2_X1 U17972 ( .A1(n16018), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14595) );
  OAI211_X1 U17973 ( .C1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n16018), .A(
        n14612), .B(n14595), .ZN(n14596) );
  AOI21_X1 U17974 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n14601), .A(
        n14596), .ZN(n14597) );
  MUX2_X1 U17975 ( .A(n14680), .B(n14609), .S(n14601), .Z(n14602) );
  XNOR2_X1 U17976 ( .A(n14602), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16048) );
  AOI22_X1 U17977 ( .A1(n16027), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        n16106), .B2(P1_REIP_REG_24__SCAN_IN), .ZN(n14603) );
  OAI21_X1 U17978 ( .B1(n14604), .B2(n16031), .A(n14603), .ZN(n14605) );
  AOI21_X1 U17979 ( .B1(n14606), .B2(n20374), .A(n14605), .ZN(n14607) );
  OAI21_X1 U17980 ( .B1(n16048), .B2(n20187), .A(n14607), .ZN(P1_U2975) );
  XNOR2_X1 U17981 ( .A(n14608), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14614) );
  NAND2_X1 U17982 ( .A1(n14609), .A2(n14611), .ZN(n14610) );
  OAI21_X1 U17983 ( .B1(n14612), .B2(n14611), .A(n14610), .ZN(n14613) );
  AOI21_X1 U17984 ( .B1(n14614), .B2(n14680), .A(n14613), .ZN(n14775) );
  NAND2_X1 U17985 ( .A1(n16106), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n14769) );
  OAI21_X1 U17986 ( .B1(n16038), .B2(n14615), .A(n14769), .ZN(n14618) );
  NOR2_X1 U17987 ( .A1(n14616), .A2(n14689), .ZN(n14617) );
  AOI211_X1 U17988 ( .C1(n16033), .C2(n14619), .A(n14618), .B(n14617), .ZN(
        n14620) );
  OAI21_X1 U17989 ( .B1(n14775), .B2(n20187), .A(n14620), .ZN(P1_U2976) );
  NAND2_X1 U17990 ( .A1(n14622), .A2(n14621), .ZN(n14623) );
  INV_X1 U17991 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14711) );
  XNOR2_X1 U17992 ( .A(n14623), .B(n14711), .ZN(n16070) );
  NAND2_X1 U17993 ( .A1(n14624), .A2(n20374), .ZN(n14628) );
  NOR2_X1 U17994 ( .A1(n20369), .A2(n21309), .ZN(n16063) );
  NOR2_X1 U17995 ( .A1(n16031), .A2(n14625), .ZN(n14626) );
  AOI211_X1 U17996 ( .C1(n16027), .C2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16063), .B(n14626), .ZN(n14627) );
  OAI211_X1 U17997 ( .C1(n20187), .C2(n16070), .A(n14628), .B(n14627), .ZN(
        P1_U2977) );
  OR2_X1 U17998 ( .A1(n20369), .A2(n21369), .ZN(n14780) );
  NOR2_X1 U17999 ( .A1(n14629), .A2(n14680), .ZN(n15851) );
  NAND2_X1 U18000 ( .A1(n14639), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14630) );
  NOR2_X1 U18001 ( .A1(n14646), .A2(n14630), .ZN(n15850) );
  AOI22_X1 U18002 ( .A1(n12717), .A2(n15851), .B1(n15850), .B2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14631) );
  XNOR2_X1 U18003 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n14631), .ZN(
        n14782) );
  NAND2_X1 U18004 ( .A1(n16034), .A2(n14782), .ZN(n14632) );
  OAI211_X1 U18005 ( .C1(n16038), .C2(n14633), .A(n14780), .B(n14632), .ZN(
        n14636) );
  NOR2_X1 U18006 ( .A1(n14634), .A2(n14689), .ZN(n14635) );
  AOI211_X1 U18007 ( .C1(n16033), .C2(n14637), .A(n14636), .B(n14635), .ZN(
        n14638) );
  INV_X1 U18008 ( .A(n14638), .ZN(P1_U2978) );
  OAI21_X1 U18009 ( .B1(n14639), .B2(n14691), .A(n14646), .ZN(n14641) );
  XNOR2_X1 U18010 ( .A(n14680), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14640) );
  XNOR2_X1 U18011 ( .A(n14641), .B(n14640), .ZN(n14792) );
  NAND2_X1 U18012 ( .A1(n16106), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n14788) );
  OAI21_X1 U18013 ( .B1(n16038), .B2(n14642), .A(n14788), .ZN(n14644) );
  NOR2_X1 U18014 ( .A1(n15880), .A2(n14689), .ZN(n14643) );
  AOI211_X1 U18015 ( .C1(n16033), .C2(n15883), .A(n14644), .B(n14643), .ZN(
        n14645) );
  OAI21_X1 U18016 ( .B1(n14792), .B2(n20187), .A(n14645), .ZN(P1_U2980) );
  OAI21_X1 U18017 ( .B1(n14648), .B2(n14647), .A(n14646), .ZN(n14810) );
  NAND2_X1 U18018 ( .A1(n15970), .A2(n20374), .ZN(n14651) );
  INV_X1 U18019 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21378) );
  NOR2_X1 U18020 ( .A1(n20369), .A2(n21378), .ZN(n14804) );
  NOR2_X1 U18021 ( .A1(n16031), .A2(n15889), .ZN(n14649) );
  AOI211_X1 U18022 ( .C1(n16027), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n14804), .B(n14649), .ZN(n14650) );
  OAI211_X1 U18023 ( .C1(n20187), .C2(n14810), .A(n14651), .B(n14650), .ZN(
        P1_U2981) );
  INV_X1 U18024 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n14652) );
  NOR2_X1 U18025 ( .A1(n20369), .A2(n14652), .ZN(n14815) );
  NOR2_X1 U18026 ( .A1(n16031), .A2(n14653), .ZN(n14654) );
  AOI211_X1 U18027 ( .C1(n16027), .C2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n14815), .B(n14654), .ZN(n14661) );
  NOR2_X1 U18028 ( .A1(n14680), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14658) );
  OAI21_X1 U18029 ( .B1(n10119), .B2(n14656), .A(n14655), .ZN(n14657) );
  MUX2_X1 U18030 ( .A(n14680), .B(n14658), .S(n14657), .Z(n14659) );
  XNOR2_X1 U18031 ( .A(n14659), .B(n14798), .ZN(n14811) );
  NAND2_X1 U18032 ( .A1(n14811), .A2(n16034), .ZN(n14660) );
  OAI211_X1 U18033 ( .C1(n14662), .C2(n14689), .A(n14661), .B(n14660), .ZN(
        P1_U2982) );
  OR2_X1 U18034 ( .A1(n16019), .A2(n14663), .ZN(n14667) );
  INV_X1 U18035 ( .A(n14664), .ZN(n14665) );
  NOR2_X1 U18036 ( .A1(n15998), .A2(n14665), .ZN(n14666) );
  NAND2_X1 U18037 ( .A1(n14667), .A2(n14666), .ZN(n15987) );
  NAND2_X1 U18038 ( .A1(n15988), .A2(n15986), .ZN(n14668) );
  XNOR2_X1 U18039 ( .A(n15987), .B(n14668), .ZN(n16081) );
  INV_X1 U18040 ( .A(n16081), .ZN(n14673) );
  INV_X1 U18041 ( .A(n15910), .ZN(n14671) );
  NOR2_X1 U18042 ( .A1(n20369), .A2(n21136), .ZN(n16078) );
  AOI21_X1 U18043 ( .B1(n16027), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16078), .ZN(n14669) );
  OAI21_X1 U18044 ( .B1(n15907), .B2(n16031), .A(n14669), .ZN(n14670) );
  AOI21_X1 U18045 ( .B1(n14671), .B2(n20374), .A(n14670), .ZN(n14672) );
  OAI21_X1 U18046 ( .B1(n14673), .B2(n20187), .A(n14672), .ZN(P1_U2984) );
  OAI21_X1 U18047 ( .B1(n16009), .B2(n15998), .A(n16010), .ZN(n14676) );
  XNOR2_X1 U18048 ( .A(n14676), .B(n14675), .ZN(n16093) );
  AOI22_X1 U18049 ( .A1(n16027), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n16106), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n14677) );
  OAI21_X1 U18050 ( .B1(n15929), .B2(n16031), .A(n14677), .ZN(n14678) );
  AOI21_X1 U18051 ( .B1(n15932), .B2(n20374), .A(n14678), .ZN(n14679) );
  OAI21_X1 U18052 ( .B1(n20187), .B2(n16093), .A(n14679), .ZN(P1_U2986) );
  NAND2_X1 U18053 ( .A1(n14683), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14682) );
  XNOR2_X1 U18054 ( .A(n16019), .B(n16132), .ZN(n14681) );
  MUX2_X1 U18055 ( .A(n14682), .B(n14681), .S(n14680), .Z(n14685) );
  NOR3_X1 U18056 ( .A1(n14683), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n14680), .ZN(n16020) );
  INV_X1 U18057 ( .A(n16020), .ZN(n14684) );
  NAND2_X1 U18058 ( .A1(n14685), .A2(n14684), .ZN(n16129) );
  NAND2_X1 U18059 ( .A1(n16129), .A2(n16034), .ZN(n14688) );
  NOR2_X1 U18060 ( .A1(n20369), .A2(n21384), .ZN(n16122) );
  NOR2_X1 U18061 ( .A1(n16031), .A2(n15956), .ZN(n14686) );
  AOI211_X1 U18062 ( .C1(n16027), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16122), .B(n14686), .ZN(n14687) );
  OAI211_X1 U18063 ( .C1(n15961), .C2(n14689), .A(n14688), .B(n14687), .ZN(
        P1_U2989) );
  INV_X1 U18064 ( .A(n14690), .ZN(n14721) );
  INV_X1 U18065 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16061) );
  INV_X1 U18066 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16077) );
  NOR2_X1 U18067 ( .A1(n16084), .A2(n16077), .ZN(n16072) );
  NAND4_X1 U18068 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A4(n16072), .ZN(n14803) );
  NOR2_X1 U18069 ( .A1(n14691), .A2(n14803), .ZN(n14704) );
  INV_X1 U18070 ( .A(n14704), .ZN(n14706) );
  NAND2_X1 U18071 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16127) );
  NOR2_X1 U18072 ( .A1(n16127), .A2(n16124), .ZN(n16115) );
  AND2_X1 U18073 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16115), .ZN(
        n16109) );
  NAND2_X1 U18074 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n16109), .ZN(
        n14793) );
  INV_X1 U18075 ( .A(n16127), .ZN(n14692) );
  NAND3_X1 U18076 ( .A1(n14694), .A2(n14693), .A3(n14692), .ZN(n16103) );
  NOR3_X1 U18077 ( .A1(n12710), .A2(n12703), .A3(n16103), .ZN(n14705) );
  INV_X1 U18078 ( .A(n14705), .ZN(n14794) );
  OAI22_X1 U18079 ( .A1(n20361), .A2(n14793), .B1(n14794), .B2(n14695), .ZN(
        n16097) );
  NAND2_X1 U18080 ( .A1(n20366), .A2(n14705), .ZN(n16100) );
  INV_X1 U18081 ( .A(n16100), .ZN(n14696) );
  NAND2_X1 U18082 ( .A1(n14767), .A2(n15859), .ZN(n16065) );
  NOR4_X1 U18083 ( .A1(n16061), .A2(n14711), .A3(n14611), .A4(n16065), .ZN(
        n16057) );
  AND2_X1 U18084 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n16057), .ZN(
        n16041) );
  NAND2_X1 U18085 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14716) );
  INV_X1 U18086 ( .A(n14716), .ZN(n14697) );
  NAND2_X1 U18087 ( .A1(n16041), .A2(n14697), .ZN(n14751) );
  INV_X1 U18088 ( .A(n14698), .ZN(n14740) );
  NOR2_X1 U18089 ( .A1(n14751), .A2(n14740), .ZN(n14734) );
  INV_X1 U18090 ( .A(n14703), .ZN(n14720) );
  NAND2_X1 U18091 ( .A1(n14705), .A2(n14704), .ZN(n14785) );
  NOR2_X1 U18092 ( .A1(n14706), .A2(n14793), .ZN(n14787) );
  NAND2_X1 U18093 ( .A1(n14707), .A2(n14787), .ZN(n14710) );
  INV_X1 U18094 ( .A(n14767), .ZN(n14708) );
  AOI211_X1 U18095 ( .C1(n14785), .C2(n14710), .A(n14709), .B(n14708), .ZN(
        n14776) );
  NOR2_X1 U18096 ( .A1(n16061), .A2(n14711), .ZN(n14766) );
  NAND2_X1 U18097 ( .A1(n14776), .A2(n14766), .ZN(n14712) );
  AND2_X1 U18098 ( .A1(n14717), .A2(n16101), .ZN(n14777) );
  INV_X1 U18099 ( .A(n14777), .ZN(n14718) );
  NAND2_X1 U18100 ( .A1(n14712), .A2(n14718), .ZN(n14765) );
  OR2_X1 U18101 ( .A1(n20361), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14713) );
  AND2_X1 U18102 ( .A1(n14765), .A2(n14713), .ZN(n16052) );
  NAND2_X1 U18103 ( .A1(n14796), .A2(n14714), .ZN(n14715) );
  NAND2_X1 U18104 ( .A1(n16052), .A2(n14715), .ZN(n16043) );
  AOI21_X1 U18105 ( .B1(n14796), .B2(n14716), .A(n16043), .ZN(n14750) );
  INV_X1 U18106 ( .A(n14750), .ZN(n14746) );
  AOI21_X1 U18107 ( .B1(n14740), .B2(n14796), .A(n14746), .ZN(n14738) );
  OAI211_X1 U18108 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n14717), .A(
        n14738), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14722) );
  NAND3_X1 U18109 ( .A1(n14722), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14718), .ZN(n14719) );
  OAI211_X1 U18110 ( .C1(n14721), .C2(n16112), .A(n14720), .B(n14719), .ZN(
        P1_U3000) );
  INV_X1 U18111 ( .A(n14722), .ZN(n14725) );
  AOI21_X1 U18112 ( .B1(n14734), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14724) );
  OAI21_X1 U18113 ( .B1(n14725), .B2(n14724), .A(n14723), .ZN(n14726) );
  AOI21_X1 U18114 ( .B1(n14727), .B2(n16135), .A(n14726), .ZN(n14728) );
  OAI21_X1 U18115 ( .B1(n14729), .B2(n16112), .A(n14728), .ZN(P1_U3001) );
  NAND2_X1 U18116 ( .A1(n14730), .A2(n20357), .ZN(n14736) );
  NOR2_X1 U18117 ( .A1(n14731), .A2(n20355), .ZN(n14732) );
  AOI211_X1 U18118 ( .C1(n14734), .C2(n14737), .A(n14733), .B(n14732), .ZN(
        n14735) );
  OAI211_X1 U18119 ( .C1(n14738), .C2(n14737), .A(n14736), .B(n14735), .ZN(
        P1_U3002) );
  INV_X1 U18120 ( .A(n14751), .ZN(n14741) );
  NAND3_X1 U18121 ( .A1(n14741), .A2(n14740), .A3(n14739), .ZN(n14742) );
  OAI211_X1 U18122 ( .C1(n14744), .C2(n20355), .A(n14743), .B(n14742), .ZN(
        n14745) );
  AOI21_X1 U18123 ( .B1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n14746), .A(
        n14745), .ZN(n14747) );
  OAI21_X1 U18124 ( .B1(n14748), .B2(n16112), .A(n14747), .ZN(P1_U3003) );
  NAND2_X1 U18125 ( .A1(n16106), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14749) );
  OAI221_X1 U18126 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14751), 
        .C1(n14573), .C2(n14750), .A(n14749), .ZN(n14752) );
  AOI21_X1 U18127 ( .B1(n14753), .B2(n16135), .A(n14752), .ZN(n14754) );
  OAI21_X1 U18128 ( .B1(n14755), .B2(n16112), .A(n14754), .ZN(P1_U3004) );
  INV_X1 U18129 ( .A(n14756), .ZN(n14764) );
  NOR2_X1 U18130 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n16040), .ZN(
        n14761) );
  INV_X1 U18131 ( .A(n14757), .ZN(n14758) );
  NOR2_X1 U18132 ( .A1(n14758), .A2(n20355), .ZN(n14759) );
  AOI211_X1 U18133 ( .C1(n16041), .C2(n14761), .A(n14760), .B(n14759), .ZN(
        n14763) );
  NAND2_X1 U18134 ( .A1(n16043), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14762) );
  OAI211_X1 U18135 ( .C1(n14764), .C2(n16112), .A(n14763), .B(n14762), .ZN(
        P1_U3005) );
  INV_X1 U18136 ( .A(n14765), .ZN(n14773) );
  NAND3_X1 U18137 ( .A1(n14767), .A2(n14766), .A3(n14611), .ZN(n16053) );
  INV_X1 U18138 ( .A(n15859), .ZN(n14771) );
  NAND2_X1 U18139 ( .A1(n14768), .A2(n16135), .ZN(n14770) );
  OAI211_X1 U18140 ( .C1(n16053), .C2(n14771), .A(n14770), .B(n14769), .ZN(
        n14772) );
  AOI21_X1 U18141 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n14773), .A(
        n14772), .ZN(n14774) );
  OAI21_X1 U18142 ( .B1(n14775), .B2(n16112), .A(n14774), .ZN(P1_U3008) );
  NOR2_X1 U18143 ( .A1(n14777), .A2(n14776), .ZN(n16067) );
  INV_X1 U18144 ( .A(n16065), .ZN(n14778) );
  AOI22_X1 U18145 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n16067), .B1(
        n16061), .B2(n14778), .ZN(n14779) );
  NAND2_X1 U18146 ( .A1(n14780), .A2(n14779), .ZN(n14781) );
  AOI21_X1 U18147 ( .B1(n20357), .B2(n14782), .A(n14781), .ZN(n14783) );
  OAI21_X1 U18148 ( .B1(n14784), .B2(n20355), .A(n14783), .ZN(P1_U3010) );
  AOI22_X1 U18149 ( .A1(n20366), .A2(n15857), .B1(n16104), .B2(n14785), .ZN(
        n14786) );
  OAI211_X1 U18150 ( .C1(n14787), .C2(n20361), .A(n16101), .B(n14786), .ZN(
        n15858) );
  NAND2_X1 U18151 ( .A1(n15858), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14789) );
  OAI211_X1 U18152 ( .C1(n15879), .C2(n20355), .A(n14789), .B(n14788), .ZN(
        n14790) );
  AOI21_X1 U18153 ( .B1(n15859), .B2(n15857), .A(n14790), .ZN(n14791) );
  OAI21_X1 U18154 ( .B1(n14792), .B2(n16112), .A(n14791), .ZN(P1_U3012) );
  NOR2_X1 U18155 ( .A1(n14812), .A2(n14793), .ZN(n16088) );
  OAI21_X1 U18156 ( .B1(n14812), .B2(n14794), .A(n16104), .ZN(n14795) );
  OAI211_X1 U18157 ( .C1(n16088), .C2(n20361), .A(n16101), .B(n14795), .ZN(
        n16096) );
  AOI21_X1 U18158 ( .B1(n16087), .B2(n14796), .A(n16096), .ZN(n16085) );
  INV_X1 U18159 ( .A(n16072), .ZN(n14797) );
  OAI21_X1 U18160 ( .B1(n14798), .B2(n14797), .A(n14796), .ZN(n14799) );
  NAND2_X1 U18161 ( .A1(n16085), .A2(n14799), .ZN(n14814) );
  AOI21_X1 U18162 ( .B1(n14802), .B2(n14801), .A(n14424), .ZN(n15969) );
  INV_X1 U18163 ( .A(n15969), .ZN(n14807) );
  NOR3_X1 U18164 ( .A1(n14813), .A2(n14803), .A3(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14805) );
  NOR2_X1 U18165 ( .A1(n14805), .A2(n14804), .ZN(n14806) );
  OAI21_X1 U18166 ( .B1(n14807), .B2(n20355), .A(n14806), .ZN(n14808) );
  AOI21_X1 U18167 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n14814), .A(
        n14808), .ZN(n14809) );
  OAI21_X1 U18168 ( .B1(n14810), .B2(n16112), .A(n14809), .ZN(P1_U3013) );
  INV_X1 U18169 ( .A(n14811), .ZN(n14819) );
  NOR3_X1 U18170 ( .A1(n14813), .A2(n16087), .A3(n14812), .ZN(n16080) );
  OAI221_X1 U18171 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n16072), 
        .C1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n16080), .A(n14814), .ZN(
        n14818) );
  AOI21_X1 U18172 ( .B1(n14816), .B2(n16135), .A(n14815), .ZN(n14817) );
  OAI211_X1 U18173 ( .C1(n14819), .C2(n16112), .A(n14818), .B(n14817), .ZN(
        P1_U3014) );
  NOR2_X1 U18174 ( .A1(n14820), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14823) );
  NOR3_X1 U18175 ( .A1(n11888), .A2(n13910), .A3(n13941), .ZN(n14822) );
  AOI211_X1 U18176 ( .C1(n20881), .C2(n14824), .A(n14823), .B(n14822), .ZN(
        n15804) );
  INV_X1 U18177 ( .A(n14825), .ZN(n14841) );
  INV_X1 U18178 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14827) );
  AOI22_X1 U18179 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n14827), .B2(n14826), .ZN(
        n14836) );
  INV_X1 U18180 ( .A(n14836), .ZN(n14829) );
  NOR2_X1 U18181 ( .A1(n16145), .A2(n20362), .ZN(n14835) );
  NOR3_X1 U18182 ( .A1(n13941), .A2(n13910), .A3(n15835), .ZN(n14828) );
  AOI21_X1 U18183 ( .B1(n14829), .B2(n14835), .A(n14828), .ZN(n14830) );
  OAI21_X1 U18184 ( .B1(n15804), .B2(n14841), .A(n14830), .ZN(n14832) );
  MUX2_X1 U18185 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14832), .S(
        n14831), .Z(P1_U3473) );
  AOI22_X1 U18186 ( .A1(n14836), .A2(n14835), .B1(n14834), .B2(n14833), .ZN(
        n14837) );
  OAI21_X1 U18187 ( .B1(n14838), .B2(n14841), .A(n14837), .ZN(n14839) );
  MUX2_X1 U18188 ( .A(n14839), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n14843), .Z(P1_U3472) );
  OAI22_X1 U18189 ( .A1(n14842), .A2(n14841), .B1(n14840), .B2(n15835), .ZN(
        n14844) );
  MUX2_X1 U18190 ( .A(n14844), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n14843), .Z(P1_U3469) );
  AOI22_X1 U18191 ( .A1(n14846), .A2(n19612), .B1(P2_STATE2_REG_0__SCAN_IN), 
        .B2(n14845), .ZN(n14849) );
  NOR2_X1 U18192 ( .A1(n20047), .A2(n20158), .ZN(n14847) );
  AOI21_X1 U18193 ( .B1(n16479), .B2(n20158), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n16483) );
  OAI22_X1 U18194 ( .A1(n14849), .A2(n14848), .B1(n14847), .B2(n16483), .ZN(
        n14853) );
  AOI21_X1 U18195 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n16478), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n14850) );
  AOI211_X1 U18196 ( .C1(n19402), .C2(n14851), .A(n14850), .B(n19014), .ZN(
        n14852) );
  MUX2_X1 U18197 ( .A(n14853), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n14852), 
        .Z(P2_U3610) );
  INV_X1 U18198 ( .A(n15412), .ZN(n14855) );
  OAI21_X1 U18199 ( .B1(n14854), .B2(n14856), .A(n14855), .ZN(n15429) );
  NOR2_X1 U18200 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n14858), .ZN(
        n14857) );
  NOR2_X1 U18201 ( .A1(n15206), .A2(n14857), .ZN(n15224) );
  INV_X1 U18202 ( .A(n14858), .ZN(n14859) );
  OAI21_X1 U18203 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n14890), .A(
        n14859), .ZN(n15240) );
  INV_X1 U18204 ( .A(n15240), .ZN(n19042) );
  INV_X1 U18205 ( .A(n14888), .ZN(n14863) );
  INV_X1 U18206 ( .A(n14860), .ZN(n14886) );
  INV_X1 U18207 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n14861) );
  NAND2_X1 U18208 ( .A1(n14886), .A2(n14861), .ZN(n14862) );
  NAND2_X1 U18209 ( .A1(n14863), .A2(n14862), .ZN(n19063) );
  INV_X1 U18210 ( .A(n19063), .ZN(n14887) );
  OR2_X1 U18211 ( .A1(n14880), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14864) );
  NAND2_X1 U18212 ( .A1(n14864), .A2(n14883), .ZN(n15282) );
  INV_X1 U18213 ( .A(n15282), .ZN(n14915) );
  OAI21_X1 U18214 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n14878), .A(
        n14881), .ZN(n19099) );
  INV_X1 U18215 ( .A(n19099), .ZN(n14879) );
  OR2_X1 U18216 ( .A1(n9925), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14866) );
  NAND2_X1 U18217 ( .A1(n14865), .A2(n14866), .ZN(n19121) );
  INV_X1 U18218 ( .A(n19121), .ZN(n14877) );
  OAI21_X1 U18219 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n14874), .A(
        n14876), .ZN(n16333) );
  INV_X1 U18220 ( .A(n16333), .ZN(n19143) );
  AOI21_X1 U18221 ( .B1(n16351), .B2(n14872), .A(n14873), .ZN(n16340) );
  AOI21_X1 U18222 ( .B1(n19177), .B2(n14870), .A(n9922), .ZN(n19184) );
  AOI21_X1 U18223 ( .B1(n19424), .B2(n14867), .A(n14871), .ZN(n19412) );
  NAND2_X1 U18224 ( .A1(n14869), .A2(n14868), .ZN(n19214) );
  NOR2_X1 U18225 ( .A1(n19412), .A2(n19214), .ZN(n19191) );
  OAI21_X1 U18226 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n14871), .A(
        n14870), .ZN(n19194) );
  NAND2_X1 U18227 ( .A1(n19191), .A2(n19194), .ZN(n19181) );
  NOR2_X1 U18228 ( .A1(n19184), .A2(n19181), .ZN(n19166) );
  OAI21_X1 U18229 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n9922), .A(
        n14872), .ZN(n19168) );
  NAND2_X1 U18230 ( .A1(n19166), .A2(n19168), .ZN(n14921) );
  NOR2_X1 U18231 ( .A1(n16340), .A2(n14921), .ZN(n19156) );
  AOI21_X1 U18232 ( .B1(n19153), .B2(n14875), .A(n14874), .ZN(n16334) );
  INV_X1 U18233 ( .A(n16334), .ZN(n19158) );
  NAND2_X1 U18234 ( .A1(n19156), .A2(n19158), .ZN(n19142) );
  NOR2_X1 U18235 ( .A1(n19143), .A2(n19142), .ZN(n19132) );
  AOI21_X1 U18236 ( .B1(n19141), .B2(n14876), .A(n9925), .ZN(n16310) );
  INV_X1 U18237 ( .A(n16310), .ZN(n19134) );
  NAND2_X1 U18238 ( .A1(n19132), .A2(n19134), .ZN(n19119) );
  NOR2_X1 U18239 ( .A1(n14877), .A2(n19119), .ZN(n19110) );
  AOI21_X1 U18240 ( .B1(n19107), .B2(n14865), .A(n14878), .ZN(n15295) );
  INV_X1 U18241 ( .A(n15295), .ZN(n19112) );
  NAND2_X1 U18242 ( .A1(n19110), .A2(n19112), .ZN(n19097) );
  NOR2_X1 U18243 ( .A1(n14879), .A2(n19097), .ZN(n19086) );
  AOI21_X1 U18244 ( .B1(n19091), .B2(n14881), .A(n14880), .ZN(n19088) );
  INV_X1 U18245 ( .A(n19088), .ZN(n14882) );
  NAND2_X1 U18246 ( .A1(n19086), .A2(n14882), .ZN(n14913) );
  NOR2_X1 U18247 ( .A1(n14915), .A2(n14913), .ZN(n19075) );
  INV_X1 U18248 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14884) );
  NAND2_X1 U18249 ( .A1(n14884), .A2(n14883), .ZN(n14885) );
  NAND2_X1 U18250 ( .A1(n14886), .A2(n14885), .ZN(n19085) );
  NAND2_X1 U18251 ( .A1(n19075), .A2(n19085), .ZN(n19062) );
  NOR2_X1 U18252 ( .A1(n14887), .A2(n19062), .ZN(n19050) );
  NOR2_X1 U18253 ( .A1(n14888), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14889) );
  NOR2_X1 U18254 ( .A1(n14890), .A2(n14889), .ZN(n19052) );
  INV_X1 U18255 ( .A(n19052), .ZN(n15252) );
  NAND2_X1 U18256 ( .A1(n19050), .A2(n15252), .ZN(n19038) );
  INV_X1 U18257 ( .A(n19037), .ZN(n14891) );
  INV_X1 U18258 ( .A(n15224), .ZN(n15793) );
  AOI221_X1 U18259 ( .B1(n15224), .B2(n14891), .C1(n15793), .C2(n19037), .A(
        n20032), .ZN(n14893) );
  INV_X1 U18260 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15222) );
  OAI22_X1 U18261 ( .A1(n15222), .A2(n19223), .B1(n20088), .B2(n19222), .ZN(
        n14892) );
  AOI211_X1 U18262 ( .C1(P2_EBX_REG_21__SCAN_IN), .C2(n19250), .A(n14893), .B(
        n14892), .ZN(n14900) );
  OR2_X1 U18263 ( .A1(n15238), .A2(n14894), .ZN(n14895) );
  NAND2_X1 U18264 ( .A1(n9857), .A2(n14895), .ZN(n15428) );
  INV_X1 U18265 ( .A(n14896), .ZN(n14897) );
  OAI22_X1 U18266 ( .A1(n15428), .A2(n19246), .B1(n14897), .B2(n19204), .ZN(
        n14898) );
  INV_X1 U18267 ( .A(n14898), .ZN(n14899) );
  OAI211_X1 U18268 ( .C1(n15429), .C2(n19207), .A(n14900), .B(n14899), .ZN(
        P2_U2834) );
  NOR2_X1 U18269 ( .A1(n14902), .A2(n14901), .ZN(n14903) );
  OR2_X1 U18270 ( .A1(n15101), .A2(n14903), .ZN(n19302) );
  NOR2_X1 U18271 ( .A1(n14906), .A2(n14905), .ZN(n14907) );
  OR2_X1 U18272 ( .A1(n14904), .A2(n14907), .ZN(n19262) );
  INV_X1 U18273 ( .A(n19262), .ZN(n15285) );
  NOR2_X1 U18274 ( .A1(n14908), .A2(n19204), .ZN(n14912) );
  AOI22_X1 U18275 ( .A1(P2_EBX_REG_16__SCAN_IN), .A2(n19250), .B1(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n19252), .ZN(n14909) );
  OAI211_X1 U18276 ( .C1(n19222), .C2(n14910), .A(n14909), .B(n19176), .ZN(
        n14911) );
  AOI211_X1 U18277 ( .C1(n15285), .C2(n19226), .A(n14912), .B(n14911), .ZN(
        n14918) );
  NAND2_X1 U18278 ( .A1(n19182), .A2(n14913), .ZN(n14914) );
  XNOR2_X1 U18279 ( .A(n14915), .B(n14914), .ZN(n14916) );
  NAND2_X1 U18280 ( .A1(n14916), .A2(n19198), .ZN(n14917) );
  OAI211_X1 U18281 ( .C1(n19302), .C2(n19207), .A(n14918), .B(n14917), .ZN(
        P2_U2839) );
  INV_X1 U18282 ( .A(n9971), .ZN(n14919) );
  OAI21_X1 U18283 ( .B1(n9880), .B2(n14920), .A(n14919), .ZN(n19288) );
  NAND2_X1 U18284 ( .A1(n19182), .A2(n14921), .ZN(n14922) );
  XNOR2_X1 U18285 ( .A(n16340), .B(n14922), .ZN(n14925) );
  AOI21_X1 U18286 ( .B1(n14924), .B2(n14923), .A(n9972), .ZN(n19324) );
  AOI22_X1 U18287 ( .A1(n19198), .A2(n14925), .B1(n19239), .B2(n19324), .ZN(
        n14932) );
  INV_X1 U18288 ( .A(n14926), .ZN(n14930) );
  AOI22_X1 U18289 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19252), .B1(
        P2_EBX_REG_8__SCAN_IN), .B2(n19250), .ZN(n14927) );
  OAI211_X1 U18290 ( .C1(n19222), .C2(n14928), .A(n14927), .B(n19176), .ZN(
        n14929) );
  AOI21_X1 U18291 ( .B1(n14930), .B2(n19241), .A(n14929), .ZN(n14931) );
  OAI211_X1 U18292 ( .C1(n19246), .C2(n19288), .A(n14932), .B(n14931), .ZN(
        P2_U2847) );
  INV_X1 U18293 ( .A(n19611), .ZN(n20143) );
  NAND2_X1 U18294 ( .A1(n19182), .A2(n15647), .ZN(n14933) );
  XNOR2_X1 U18295 ( .A(n14934), .B(n14933), .ZN(n14935) );
  NAND2_X1 U18296 ( .A1(n14935), .A2(n19198), .ZN(n14944) );
  INV_X1 U18297 ( .A(n20145), .ZN(n19333) );
  OAI22_X1 U18298 ( .A1(n19203), .A2(n10576), .B1(n10580), .B2(n19222), .ZN(
        n14938) );
  NOR2_X1 U18299 ( .A1(n19223), .A2(n14936), .ZN(n14937) );
  AOI211_X1 U18300 ( .C1(n19241), .C2(n14939), .A(n14938), .B(n14937), .ZN(
        n14940) );
  OAI21_X1 U18301 ( .B1(n19333), .B2(n19207), .A(n14940), .ZN(n14941) );
  AOI21_X1 U18302 ( .B1(n14942), .B2(n19226), .A(n14941), .ZN(n14943) );
  OAI211_X1 U18303 ( .C1(n19247), .C2(n20143), .A(n14944), .B(n14943), .ZN(
        P2_U2853) );
  NOR2_X1 U18304 ( .A1(n15330), .A2(n14945), .ZN(n14950) );
  AOI21_X1 U18305 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n14945), .A(n14950), .ZN(
        n14951) );
  OAI21_X1 U18306 ( .B1(n14952), .B2(n19289), .A(n14951), .ZN(P2_U2857) );
  INV_X1 U18307 ( .A(n16178), .ZN(n15127) );
  INV_X1 U18308 ( .A(n14953), .ZN(n15022) );
  NAND2_X1 U18309 ( .A1(n14955), .A2(n14954), .ZN(n15021) );
  NAND3_X1 U18310 ( .A1(n15022), .A2(n19278), .A3(n15021), .ZN(n14957) );
  NAND2_X1 U18311 ( .A1(n14945), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14956) );
  OAI211_X1 U18312 ( .C1(n14945), .C2(n15127), .A(n14957), .B(n14956), .ZN(
        P2_U2858) );
  NAND2_X1 U18313 ( .A1(n14958), .A2(n14959), .ZN(n14960) );
  NAND2_X1 U18314 ( .A1(n14961), .A2(n14960), .ZN(n16186) );
  NOR2_X1 U18315 ( .A1(n14963), .A2(n14962), .ZN(n14965) );
  XNOR2_X1 U18316 ( .A(n14965), .B(n14964), .ZN(n15035) );
  NAND2_X1 U18317 ( .A1(n15035), .A2(n19278), .ZN(n14967) );
  NAND2_X1 U18318 ( .A1(n14945), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n14966) );
  OAI211_X1 U18319 ( .C1(n16186), .C2(n14945), .A(n14967), .B(n14966), .ZN(
        P2_U2859) );
  OR2_X1 U18320 ( .A1(n14968), .A2(n14969), .ZN(n14970) );
  NAND2_X1 U18321 ( .A1(n14958), .A2(n14970), .ZN(n16204) );
  AOI21_X1 U18322 ( .B1(n14973), .B2(n14972), .A(n14971), .ZN(n15045) );
  NAND2_X1 U18323 ( .A1(n15045), .A2(n19278), .ZN(n14975) );
  NAND2_X1 U18324 ( .A1(n14945), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n14974) );
  OAI211_X1 U18325 ( .C1(n16204), .C2(n14945), .A(n14975), .B(n14974), .ZN(
        P2_U2860) );
  OAI21_X1 U18326 ( .B1(n14976), .B2(n14978), .A(n14977), .ZN(n15052) );
  NOR2_X1 U18327 ( .A1(n14979), .A2(n14980), .ZN(n14981) );
  OR2_X1 U18328 ( .A1(n14968), .A2(n14981), .ZN(n15157) );
  NOR2_X1 U18329 ( .A1(n15157), .A2(n14945), .ZN(n14982) );
  AOI21_X1 U18330 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n14945), .A(n14982), .ZN(
        n14983) );
  OAI21_X1 U18331 ( .B1(n15052), .B2(n19289), .A(n14983), .ZN(P2_U2861) );
  OAI21_X1 U18332 ( .B1(n14984), .B2(n14986), .A(n14985), .ZN(n15062) );
  INV_X1 U18333 ( .A(n14987), .ZN(n14989) );
  INV_X1 U18334 ( .A(n14997), .ZN(n14988) );
  AOI21_X1 U18335 ( .B1(n14989), .B2(n14988), .A(n14979), .ZN(n16227) );
  NOR2_X1 U18336 ( .A1(n19293), .A2(n16222), .ZN(n14990) );
  AOI21_X1 U18337 ( .B1(n16227), .B2(n19293), .A(n14990), .ZN(n14991) );
  OAI21_X1 U18338 ( .B1(n15062), .B2(n19289), .A(n14991), .ZN(P2_U2862) );
  AOI21_X1 U18339 ( .B1(n14992), .B2(n14993), .A(n9863), .ZN(n14994) );
  XOR2_X1 U18340 ( .A(n14995), .B(n14994), .Z(n15071) );
  AND2_X1 U18341 ( .A1(n15192), .A2(n14996), .ZN(n14998) );
  OR2_X1 U18342 ( .A1(n14998), .A2(n14997), .ZN(n16239) );
  MUX2_X1 U18343 ( .A(n16239), .B(n14999), .S(n14945), .Z(n15000) );
  OAI21_X1 U18344 ( .B1(n15071), .B2(n19289), .A(n15000), .ZN(P2_U2863) );
  INV_X1 U18345 ( .A(n9937), .ZN(n16274) );
  AND2_X1 U18346 ( .A1(n16274), .A2(n15002), .ZN(n16269) );
  OR2_X1 U18347 ( .A1(n16269), .A2(n15003), .ZN(n15004) );
  AND2_X1 U18348 ( .A1(n15001), .A2(n15004), .ZN(n15087) );
  NAND2_X1 U18349 ( .A1(n15087), .A2(n19278), .ZN(n15006) );
  NAND2_X1 U18350 ( .A1(n14945), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n15005) );
  OAI211_X1 U18351 ( .C1(n15428), .C2(n14945), .A(n15006), .B(n15005), .ZN(
        P2_U2866) );
  INV_X1 U18352 ( .A(n15007), .ZN(n15008) );
  OR2_X1 U18353 ( .A1(n9937), .A2(n15007), .ZN(n16270) );
  OAI21_X1 U18354 ( .B1(n16274), .B2(n15008), .A(n16270), .ZN(n15099) );
  AND2_X1 U18355 ( .A1(n9926), .A2(n15009), .ZN(n15010) );
  OR2_X1 U18356 ( .A1(n15010), .A2(n15236), .ZN(n19056) );
  NOR2_X1 U18357 ( .A1(n19056), .A2(n14945), .ZN(n15011) );
  AOI21_X1 U18358 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n14945), .A(n15011), .ZN(
        n15012) );
  OAI21_X1 U18359 ( .B1(n19289), .B2(n15099), .A(n15012), .ZN(P2_U2868) );
  NOR2_X1 U18360 ( .A1(n15014), .A2(n15015), .ZN(n15016) );
  OR2_X1 U18361 ( .A1(n15013), .A2(n15016), .ZN(n15108) );
  OR2_X1 U18362 ( .A1(n14904), .A2(n15017), .ZN(n15018) );
  NAND2_X1 U18363 ( .A1(n15265), .A2(n15018), .ZN(n15484) );
  NOR2_X1 U18364 ( .A1(n15484), .A2(n14945), .ZN(n15019) );
  AOI21_X1 U18365 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n14945), .A(n15019), .ZN(
        n15020) );
  OAI21_X1 U18366 ( .B1(n15108), .B2(n19289), .A(n15020), .ZN(P2_U2870) );
  NAND3_X1 U18367 ( .A1(n15022), .A2(n19342), .A3(n15021), .ZN(n15027) );
  AOI22_X1 U18368 ( .A1(n19298), .A2(n15023), .B1(n19356), .B2(
        P2_EAX_REG_29__SCAN_IN), .ZN(n15026) );
  AOI22_X1 U18369 ( .A1(n19299), .A2(BUF1_REG_29__SCAN_IN), .B1(n19300), .B2(
        BUF2_REG_29__SCAN_IN), .ZN(n15025) );
  NAND2_X1 U18370 ( .A1(n19357), .A2(n16177), .ZN(n15024) );
  NAND4_X1 U18371 ( .A1(n15027), .A2(n15026), .A3(n15025), .A4(n15024), .ZN(
        P2_U2890) );
  OR2_X1 U18372 ( .A1(n15040), .A2(n15028), .ZN(n15029) );
  NAND2_X1 U18373 ( .A1(n15030), .A2(n15029), .ZN(n16197) );
  AOI22_X1 U18374 ( .A1(n19299), .A2(BUF1_REG_28__SCAN_IN), .B1(n19300), .B2(
        BUF2_REG_28__SCAN_IN), .ZN(n15033) );
  AOI22_X1 U18375 ( .A1(n19298), .A2(n15031), .B1(n19356), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n15032) );
  OAI211_X1 U18376 ( .C1(n19348), .C2(n16197), .A(n15033), .B(n15032), .ZN(
        n15034) );
  AOI21_X1 U18377 ( .B1(n15035), .B2(n19342), .A(n15034), .ZN(n15036) );
  INV_X1 U18378 ( .A(n15036), .ZN(P2_U2891) );
  NOR2_X1 U18379 ( .A1(n15037), .A2(n15038), .ZN(n15039) );
  AOI22_X1 U18380 ( .A1(n19299), .A2(BUF1_REG_27__SCAN_IN), .B1(n19300), .B2(
        BUF2_REG_27__SCAN_IN), .ZN(n15043) );
  AOI22_X1 U18381 ( .A1(n19298), .A2(n15041), .B1(n19356), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n15042) );
  OAI211_X1 U18382 ( .C1(n19348), .C2(n16211), .A(n15043), .B(n15042), .ZN(
        n15044) );
  AOI21_X1 U18383 ( .B1(n15045), .B2(n19342), .A(n15044), .ZN(n15046) );
  INV_X1 U18384 ( .A(n15046), .ZN(P2_U2892) );
  INV_X1 U18385 ( .A(n15037), .ZN(n15047) );
  OAI21_X1 U18386 ( .B1(n15053), .B2(n15048), .A(n15047), .ZN(n15354) );
  OAI22_X1 U18387 ( .A1(n19348), .A2(n15354), .B1(n19347), .B2(n13567), .ZN(
        n15049) );
  AOI21_X1 U18388 ( .B1(n19298), .B2(n19319), .A(n15049), .ZN(n15051) );
  AOI22_X1 U18389 ( .A1(n19299), .A2(BUF1_REG_26__SCAN_IN), .B1(n19300), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n15050) );
  OAI211_X1 U18390 ( .C1(n15052), .C2(n19361), .A(n15051), .B(n15050), .ZN(
        P2_U2893) );
  INV_X1 U18391 ( .A(n15053), .ZN(n15056) );
  NAND2_X1 U18392 ( .A1(n15066), .A2(n15054), .ZN(n15055) );
  NAND2_X1 U18393 ( .A1(n15056), .A2(n15055), .ZN(n16225) );
  AOI22_X1 U18394 ( .A1(n19299), .A2(BUF1_REG_25__SCAN_IN), .B1(n19300), .B2(
        BUF2_REG_25__SCAN_IN), .ZN(n15059) );
  AOI22_X1 U18395 ( .A1(n19298), .A2(n15057), .B1(n19356), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n15058) );
  OAI211_X1 U18396 ( .C1(n19348), .C2(n16225), .A(n15059), .B(n15058), .ZN(
        n15060) );
  INV_X1 U18397 ( .A(n15060), .ZN(n15061) );
  OAI21_X1 U18398 ( .B1(n15062), .B2(n19361), .A(n15061), .ZN(P2_U2894) );
  NAND2_X1 U18399 ( .A1(n15063), .A2(n15064), .ZN(n15065) );
  AND2_X1 U18400 ( .A1(n15066), .A2(n15065), .ZN(n16237) );
  INV_X1 U18401 ( .A(n19298), .ZN(n15103) );
  INV_X1 U18402 ( .A(n19326), .ZN(n15067) );
  OAI22_X1 U18403 ( .A1(n15103), .A2(n15067), .B1(n19347), .B2(n13581), .ZN(
        n15068) );
  AOI21_X1 U18404 ( .B1(n19357), .B2(n16237), .A(n15068), .ZN(n15070) );
  AOI22_X1 U18405 ( .A1(n19299), .A2(BUF1_REG_24__SCAN_IN), .B1(n19300), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n15069) );
  OAI211_X1 U18406 ( .C1(n15071), .C2(n19361), .A(n15070), .B(n15069), .ZN(
        P2_U2895) );
  AOI21_X1 U18407 ( .B1(n15072), .B2(n15074), .A(n15073), .ZN(n16263) );
  OR2_X1 U18408 ( .A1(n15415), .A2(n15075), .ZN(n15076) );
  NAND2_X1 U18409 ( .A1(n15063), .A2(n15076), .ZN(n16259) );
  AOI22_X1 U18410 ( .A1(n19299), .A2(BUF1_REG_23__SCAN_IN), .B1(n19300), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n15079) );
  AOI22_X1 U18411 ( .A1(n19298), .A2(n15077), .B1(n19356), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n15078) );
  OAI211_X1 U18412 ( .C1(n19348), .C2(n16259), .A(n15079), .B(n15078), .ZN(
        n15080) );
  AOI21_X1 U18413 ( .B1(n16263), .B2(n19342), .A(n15080), .ZN(n15081) );
  INV_X1 U18414 ( .A(n15081), .ZN(P2_U2896) );
  OAI22_X1 U18415 ( .A1(n15103), .A2(n19471), .B1(n19347), .B2(n15082), .ZN(
        n15086) );
  INV_X1 U18416 ( .A(n19300), .ZN(n15084) );
  INV_X1 U18417 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n15083) );
  NOR2_X1 U18418 ( .A1(n15084), .A2(n15083), .ZN(n15085) );
  AOI211_X1 U18419 ( .C1(BUF1_REG_21__SCAN_IN), .C2(n19299), .A(n15086), .B(
        n15085), .ZN(n15089) );
  NAND2_X1 U18420 ( .A1(n15087), .A2(n19342), .ZN(n15088) );
  OAI211_X1 U18421 ( .C1(n15429), .C2(n19348), .A(n15089), .B(n15088), .ZN(
        P2_U2898) );
  AND2_X1 U18422 ( .A1(n15465), .A2(n15091), .ZN(n15092) );
  NOR2_X1 U18423 ( .A1(n15090), .A2(n15092), .ZN(n19058) );
  NAND2_X1 U18424 ( .A1(n19299), .A2(BUF1_REG_19__SCAN_IN), .ZN(n15096) );
  NAND2_X1 U18425 ( .A1(n19300), .A2(BUF2_REG_19__SCAN_IN), .ZN(n15095) );
  AOI22_X1 U18426 ( .A1(n19298), .A2(n15093), .B1(n19356), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n15094) );
  NAND3_X1 U18427 ( .A1(n15096), .A2(n15095), .A3(n15094), .ZN(n15097) );
  AOI21_X1 U18428 ( .B1(n19058), .B2(n19357), .A(n15097), .ZN(n15098) );
  OAI21_X1 U18429 ( .B1(n19361), .B2(n15099), .A(n15098), .ZN(P2_U2900) );
  OAI21_X1 U18430 ( .B1(n15101), .B2(n15100), .A(n15463), .ZN(n15488) );
  INV_X1 U18431 ( .A(n15488), .ZN(n19081) );
  NAND2_X1 U18432 ( .A1(n19081), .A2(n19357), .ZN(n15107) );
  OAI22_X1 U18433 ( .A1(n15103), .A2(n19448), .B1(n19347), .B2(n15102), .ZN(
        n15105) );
  AND2_X1 U18434 ( .A1(n19300), .A2(BUF2_REG_17__SCAN_IN), .ZN(n15104) );
  AOI211_X1 U18435 ( .C1(BUF1_REG_17__SCAN_IN), .C2(n19299), .A(n15105), .B(
        n15104), .ZN(n15106) );
  OAI211_X1 U18436 ( .C1(n15108), .C2(n19361), .A(n15107), .B(n15106), .ZN(
        P2_U2902) );
  NAND2_X1 U18437 ( .A1(n15110), .A2(n15109), .ZN(n15113) );
  NOR2_X1 U18438 ( .A1(n15111), .A2(n9862), .ZN(n15112) );
  XNOR2_X1 U18439 ( .A(n15113), .B(n15112), .ZN(n15333) );
  XNOR2_X1 U18440 ( .A(n15122), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16171) );
  NAND2_X1 U18441 ( .A1(n19414), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n15320) );
  NAND2_X1 U18442 ( .A1(n16316), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15114) );
  OAI211_X1 U18443 ( .C1(n16355), .C2(n16171), .A(n15320), .B(n15114), .ZN(
        n15118) );
  OAI21_X1 U18444 ( .B1(n15116), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n15115), .ZN(n15328) );
  NOR2_X1 U18445 ( .A1(n15328), .A2(n16371), .ZN(n15117) );
  AOI211_X1 U18446 ( .C1(n16363), .C2(n16169), .A(n15118), .B(n15117), .ZN(
        n15119) );
  OAI21_X1 U18447 ( .B1(n15333), .B2(n19417), .A(n15119), .ZN(P2_U2984) );
  AOI21_X1 U18448 ( .B1(n16316), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15120), .ZN(n15126) );
  INV_X1 U18449 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15124) );
  INV_X1 U18450 ( .A(n15121), .ZN(n15123) );
  AOI21_X1 U18451 ( .B1(n15124), .B2(n15123), .A(n15122), .ZN(n16152) );
  NAND2_X1 U18452 ( .A1(n19413), .A2(n16152), .ZN(n15125) );
  OAI211_X1 U18453 ( .C1(n15127), .C2(n19416), .A(n15126), .B(n15125), .ZN(
        n15128) );
  AOI21_X1 U18454 ( .B1(n19421), .B2(n15129), .A(n15128), .ZN(n15130) );
  OAI21_X1 U18455 ( .B1(n15131), .B2(n19417), .A(n15130), .ZN(P2_U2985) );
  INV_X1 U18456 ( .A(n15134), .ZN(n15136) );
  OAI22_X1 U18457 ( .A1(n15146), .A2(n15148), .B1(n15136), .B2(n15135), .ZN(
        n15139) );
  XNOR2_X1 U18458 ( .A(n15137), .B(n10961), .ZN(n15138) );
  XNOR2_X1 U18459 ( .A(n15139), .B(n15138), .ZN(n15344) );
  XNOR2_X1 U18460 ( .A(n15140), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15342) );
  INV_X1 U18461 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n20102) );
  NOR2_X1 U18462 ( .A1(n19176), .A2(n20102), .ZN(n15334) );
  NOR2_X1 U18463 ( .A1(n15149), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15141) );
  OR2_X1 U18464 ( .A1(n15121), .A2(n15141), .ZN(n16194) );
  NOR2_X1 U18465 ( .A1(n16355), .A2(n16194), .ZN(n15142) );
  AOI211_X1 U18466 ( .C1(n16316), .C2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15334), .B(n15142), .ZN(n15143) );
  OAI21_X1 U18467 ( .B1(n16186), .B2(n19416), .A(n15143), .ZN(n15144) );
  AOI21_X1 U18468 ( .B1(n15342), .B2(n19421), .A(n15144), .ZN(n15145) );
  OAI21_X1 U18469 ( .B1(n15344), .B2(n19417), .A(n15145), .ZN(P2_U2986) );
  XNOR2_X1 U18470 ( .A(n15146), .B(n15148), .ZN(n15353) );
  AOI21_X1 U18471 ( .B1(n15148), .B2(n15161), .A(n15147), .ZN(n15351) );
  AOI21_X1 U18472 ( .B1(n16198), .B2(n9966), .A(n15149), .ZN(n16153) );
  NAND2_X1 U18473 ( .A1(n19414), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15345) );
  OAI21_X1 U18474 ( .B1(n19425), .B2(n16198), .A(n15345), .ZN(n15150) );
  AOI21_X1 U18475 ( .B1(n19413), .B2(n16153), .A(n15150), .ZN(n15151) );
  OAI21_X1 U18476 ( .B1(n16204), .B2(n19416), .A(n15151), .ZN(n15152) );
  AOI21_X1 U18477 ( .B1(n15351), .B2(n19421), .A(n15152), .ZN(n15153) );
  OAI21_X1 U18478 ( .B1(n15353), .B2(n19417), .A(n15153), .ZN(P2_U2987) );
  OAI21_X1 U18479 ( .B1(n15154), .B2(n15166), .A(n15165), .ZN(n15155) );
  XOR2_X1 U18480 ( .A(n15156), .B(n15155), .Z(n15364) );
  NAND2_X1 U18481 ( .A1(n15168), .A2(n15158), .ZN(n15159) );
  NAND2_X1 U18482 ( .A1(n9966), .A2(n15159), .ZN(n16217) );
  NOR2_X1 U18483 ( .A1(n19176), .A2(n20098), .ZN(n15355) );
  AOI21_X1 U18484 ( .B1(n16316), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15355), .ZN(n15160) );
  OAI21_X1 U18485 ( .B1(n16355), .B2(n16217), .A(n15160), .ZN(n15163) );
  NOR2_X1 U18486 ( .A1(n15172), .A2(n15369), .ZN(n15370) );
  OAI21_X1 U18487 ( .B1(n15370), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15161), .ZN(n15360) );
  NOR2_X1 U18488 ( .A1(n15360), .A2(n16371), .ZN(n15162) );
  AOI211_X1 U18489 ( .C1(n16363), .C2(n16214), .A(n15163), .B(n15162), .ZN(
        n15164) );
  OAI21_X1 U18490 ( .B1(n15364), .B2(n19417), .A(n15164), .ZN(P2_U2988) );
  NOR2_X1 U18491 ( .A1(n15166), .A2(n10954), .ZN(n15167) );
  XNOR2_X1 U18492 ( .A(n15154), .B(n15167), .ZN(n15375) );
  INV_X1 U18493 ( .A(n15168), .ZN(n15169) );
  AOI21_X1 U18494 ( .B1(n15171), .B2(n15182), .A(n15169), .ZN(n16154) );
  NAND2_X1 U18495 ( .A1(n19413), .A2(n16154), .ZN(n15170) );
  NAND2_X1 U18496 ( .A1(n19414), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15365) );
  OAI211_X1 U18497 ( .C1(n19425), .C2(n15171), .A(n15170), .B(n15365), .ZN(
        n15174) );
  NOR2_X1 U18498 ( .A1(n11081), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15371) );
  NOR3_X1 U18499 ( .A1(n15371), .A2(n15370), .A3(n16371), .ZN(n15173) );
  AOI211_X1 U18500 ( .C1(n16363), .C2(n16227), .A(n15174), .B(n15173), .ZN(
        n15175) );
  OAI21_X1 U18501 ( .B1(n15375), .B2(n19417), .A(n15175), .ZN(P2_U2989) );
  XNOR2_X1 U18502 ( .A(n15178), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15179) );
  XNOR2_X1 U18503 ( .A(n15177), .B(n15179), .ZN(n15385) );
  INV_X1 U18504 ( .A(n9908), .ZN(n15180) );
  AOI21_X1 U18505 ( .B1(n15377), .B2(n15180), .A(n11081), .ZN(n15383) );
  INV_X1 U18506 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20094) );
  NOR2_X1 U18507 ( .A1(n19176), .A2(n20094), .ZN(n15380) );
  OR2_X1 U18508 ( .A1(n15193), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15181) );
  NAND2_X1 U18509 ( .A1(n15182), .A2(n15181), .ZN(n16243) );
  NOR2_X1 U18510 ( .A1(n16355), .A2(n16243), .ZN(n15183) );
  AOI211_X1 U18511 ( .C1(n16316), .C2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15380), .B(n15183), .ZN(n15184) );
  OAI21_X1 U18512 ( .B1(n16239), .B2(n19416), .A(n15184), .ZN(n15185) );
  AOI21_X1 U18513 ( .B1(n15383), .B2(n19421), .A(n15185), .ZN(n15186) );
  OAI21_X1 U18514 ( .B1(n15385), .B2(n19417), .A(n15186), .ZN(P2_U2990) );
  XNOR2_X1 U18515 ( .A(n9830), .B(n15188), .ZN(n15405) );
  AOI21_X1 U18516 ( .B1(n15395), .B2(n15419), .A(n9908), .ZN(n15402) );
  NAND2_X1 U18517 ( .A1(n15204), .A2(n15190), .ZN(n15191) );
  NAND2_X1 U18518 ( .A1(n15192), .A2(n15191), .ZN(n15386) );
  AOI21_X1 U18519 ( .B1(n16249), .B2(n15205), .A(n15193), .ZN(n16156) );
  NAND2_X1 U18520 ( .A1(n19414), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n15399) );
  OAI21_X1 U18521 ( .B1(n19425), .B2(n16249), .A(n15399), .ZN(n15194) );
  AOI21_X1 U18522 ( .B1(n19413), .B2(n16156), .A(n15194), .ZN(n15195) );
  OAI21_X1 U18523 ( .B1(n15386), .B2(n19416), .A(n15195), .ZN(n15196) );
  AOI21_X1 U18524 ( .B1(n15402), .B2(n19421), .A(n15196), .ZN(n15197) );
  OAI21_X1 U18525 ( .B1(n15405), .B2(n19417), .A(n15197), .ZN(P2_U2991) );
  NAND2_X1 U18526 ( .A1(n10367), .A2(n15200), .ZN(n15201) );
  XNOR2_X1 U18527 ( .A(n15198), .B(n15201), .ZN(n15423) );
  NAND2_X1 U18528 ( .A1(n9857), .A2(n15202), .ZN(n15203) );
  NAND2_X1 U18529 ( .A1(n15204), .A2(n15203), .ZN(n16268) );
  INV_X1 U18530 ( .A(n16268), .ZN(n15418) );
  OAI21_X1 U18531 ( .B1(n15206), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15205), .ZN(n15796) );
  AOI22_X1 U18532 ( .A1(n16316), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19414), .ZN(n15207) );
  OAI21_X1 U18533 ( .B1(n16355), .B2(n15796), .A(n15207), .ZN(n15208) );
  AOI21_X1 U18534 ( .B1(n15418), .B2(n16363), .A(n15208), .ZN(n15210) );
  OR2_X1 U18535 ( .A1(n9909), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15420) );
  NAND3_X1 U18536 ( .A1(n15420), .A2(n19421), .A3(n15419), .ZN(n15209) );
  OAI211_X1 U18537 ( .C1(n15423), .C2(n19417), .A(n15210), .B(n15209), .ZN(
        P2_U2992) );
  NOR2_X1 U18538 ( .A1(n15212), .A2(n15211), .ZN(n15219) );
  INV_X1 U18539 ( .A(n15533), .ZN(n15214) );
  INV_X1 U18540 ( .A(n15272), .ZN(n15215) );
  INV_X1 U18541 ( .A(n15217), .ZN(n15218) );
  NAND2_X1 U18542 ( .A1(n15220), .A2(n15391), .ZN(n15229) );
  AOI21_X1 U18543 ( .B1(n15221), .B2(n15229), .A(n9909), .ZN(n15432) );
  AND2_X1 U18544 ( .A1(n19414), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15424) );
  NOR2_X1 U18545 ( .A1(n19425), .A2(n15222), .ZN(n15223) );
  AOI211_X1 U18546 ( .C1(n15224), .C2(n19413), .A(n15424), .B(n15223), .ZN(
        n15225) );
  OAI21_X1 U18547 ( .B1(n15428), .B2(n19416), .A(n15225), .ZN(n15226) );
  AOI21_X1 U18548 ( .B1(n15432), .B2(n19421), .A(n15226), .ZN(n15227) );
  OAI21_X1 U18549 ( .B1(n15434), .B2(n19417), .A(n15227), .ZN(P2_U2993) );
  NAND2_X1 U18550 ( .A1(n15220), .A2(n15478), .ZN(n15519) );
  INV_X1 U18551 ( .A(n15437), .ZN(n15228) );
  NOR2_X1 U18552 ( .A1(n15519), .A2(n15228), .ZN(n15250) );
  OAI21_X1 U18553 ( .B1(n15250), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15229), .ZN(n15452) );
  INV_X1 U18554 ( .A(n15230), .ZN(n15232) );
  NOR2_X1 U18555 ( .A1(n15236), .A2(n15235), .ZN(n15237) );
  OR2_X1 U18556 ( .A1(n15238), .A2(n15237), .ZN(n19043) );
  INV_X1 U18557 ( .A(n19043), .ZN(n15449) );
  NAND2_X1 U18558 ( .A1(n19414), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n15442) );
  NAND2_X1 U18559 ( .A1(n16316), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15239) );
  OAI211_X1 U18560 ( .C1(n16355), .C2(n15240), .A(n15442), .B(n15239), .ZN(
        n15241) );
  AOI21_X1 U18561 ( .B1(n15449), .B2(n16363), .A(n15241), .ZN(n15242) );
  OAI211_X1 U18562 ( .C1(n16371), .C2(n15452), .A(n15243), .B(n15242), .ZN(
        P2_U2994) );
  NOR2_X1 U18563 ( .A1(n15244), .A2(n15258), .ZN(n15249) );
  INV_X1 U18564 ( .A(n15245), .ZN(n15246) );
  NOR2_X1 U18565 ( .A1(n15247), .A2(n15246), .ZN(n15248) );
  XNOR2_X1 U18566 ( .A(n15249), .B(n15248), .ZN(n15461) );
  OR2_X1 U18567 ( .A1(n15519), .A2(n15438), .ZN(n15261) );
  AOI21_X1 U18568 ( .B1(n15251), .B2(n15261), .A(n15250), .ZN(n15459) );
  INV_X1 U18569 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n20085) );
  NOR2_X1 U18570 ( .A1(n19176), .A2(n20085), .ZN(n15454) );
  NOR2_X1 U18571 ( .A1(n16355), .A2(n15252), .ZN(n15253) );
  AOI211_X1 U18572 ( .C1(n16316), .C2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n15454), .B(n15253), .ZN(n15254) );
  OAI21_X1 U18573 ( .B1(n19056), .B2(n19416), .A(n15254), .ZN(n15255) );
  AOI21_X1 U18574 ( .B1(n15459), .B2(n19421), .A(n15255), .ZN(n15256) );
  OAI21_X1 U18575 ( .B1(n15461), .B2(n19417), .A(n15256), .ZN(P2_U2995) );
  NOR2_X1 U18576 ( .A1(n15258), .A2(n15257), .ZN(n15259) );
  XNOR2_X1 U18577 ( .A(n15260), .B(n15259), .ZN(n15477) );
  INV_X1 U18578 ( .A(n15519), .ZN(n15514) );
  AOI21_X1 U18579 ( .B1(n15479), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15263) );
  INV_X1 U18580 ( .A(n15261), .ZN(n15262) );
  NOR2_X1 U18581 ( .A1(n15263), .A2(n15262), .ZN(n15475) );
  NAND2_X1 U18582 ( .A1(n15265), .A2(n15264), .ZN(n15266) );
  NAND2_X1 U18583 ( .A1(n9926), .A2(n15266), .ZN(n19067) );
  INV_X1 U18584 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n20083) );
  NOR2_X1 U18585 ( .A1(n19176), .A2(n20083), .ZN(n15470) );
  NOR2_X1 U18586 ( .A1(n16355), .A2(n19063), .ZN(n15267) );
  AOI211_X1 U18587 ( .C1(n16316), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15470), .B(n15267), .ZN(n15268) );
  OAI21_X1 U18588 ( .B1(n19067), .B2(n19416), .A(n15268), .ZN(n15269) );
  AOI21_X1 U18589 ( .B1(n15475), .B2(n19421), .A(n15269), .ZN(n15270) );
  OAI21_X1 U18590 ( .B1(n15477), .B2(n19417), .A(n15270), .ZN(P2_U2996) );
  NAND2_X1 U18591 ( .A1(n15272), .A2(n15271), .ZN(n15275) );
  NAND2_X1 U18592 ( .A1(n15498), .A2(n15273), .ZN(n15274) );
  XOR2_X1 U18593 ( .A(n15275), .B(n15274), .Z(n15492) );
  XNOR2_X1 U18594 ( .A(n15479), .B(n15483), .ZN(n15279) );
  NOR2_X1 U18595 ( .A1(n19176), .A2(n20081), .ZN(n15485) );
  NOR2_X1 U18596 ( .A1(n16355), .A2(n19085), .ZN(n15276) );
  AOI211_X1 U18597 ( .C1(n16316), .C2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n15485), .B(n15276), .ZN(n15277) );
  OAI21_X1 U18598 ( .B1(n15484), .B2(n19416), .A(n15277), .ZN(n15278) );
  AOI21_X1 U18599 ( .B1(n15279), .B2(n19421), .A(n15278), .ZN(n15280) );
  OAI21_X1 U18600 ( .B1(n15492), .B2(n19417), .A(n15280), .ZN(P2_U2997) );
  NAND2_X1 U18601 ( .A1(n19414), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n15493) );
  NAND2_X1 U18602 ( .A1(n16316), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15281) );
  OAI211_X1 U18603 ( .C1(n16355), .C2(n15282), .A(n15493), .B(n15281), .ZN(
        n15284) );
  AOI211_X1 U18604 ( .C1(n15501), .C2(n15513), .A(n16371), .B(n15479), .ZN(
        n15283) );
  AOI211_X1 U18605 ( .C1(n16363), .C2(n15285), .A(n15284), .B(n15283), .ZN(
        n15289) );
  OR2_X1 U18606 ( .A1(n15287), .A2(n15286), .ZN(n15497) );
  NAND3_X1 U18607 ( .A1(n15498), .A2(n15497), .A3(n16366), .ZN(n15288) );
  NAND2_X1 U18608 ( .A1(n15289), .A2(n15288), .ZN(P2_U2998) );
  NAND2_X1 U18609 ( .A1(n15220), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16328) );
  NAND2_X1 U18610 ( .A1(n16327), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15570) );
  XNOR2_X1 U18611 ( .A(n15556), .B(n15545), .ZN(n15554) );
  NAND2_X1 U18612 ( .A1(n15292), .A2(n15291), .ZN(n15293) );
  XNOR2_X1 U18613 ( .A(n15290), .B(n15293), .ZN(n15552) );
  NAND2_X1 U18614 ( .A1(n19414), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n15542) );
  OAI21_X1 U18615 ( .B1(n19425), .B2(n19107), .A(n15542), .ZN(n15294) );
  AOI21_X1 U18616 ( .B1(n19413), .B2(n15295), .A(n15294), .ZN(n15296) );
  OAI21_X1 U18617 ( .B1(n19113), .B2(n19416), .A(n15296), .ZN(n15297) );
  AOI21_X1 U18618 ( .B1(n15552), .B2(n16366), .A(n15297), .ZN(n15298) );
  OAI21_X1 U18619 ( .B1(n15554), .B2(n16371), .A(n15298), .ZN(P2_U3001) );
  XNOR2_X1 U18620 ( .A(n15300), .B(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15301) );
  XNOR2_X1 U18621 ( .A(n15299), .B(n15301), .ZN(n15569) );
  NAND2_X1 U18622 ( .A1(n15570), .A2(n15546), .ZN(n15555) );
  NAND3_X1 U18623 ( .A1(n15556), .A2(n19421), .A3(n15555), .ZN(n15309) );
  AND2_X1 U18624 ( .A1(n15303), .A2(n15302), .ZN(n15304) );
  NOR2_X1 U18625 ( .A1(n15305), .A2(n15304), .ZN(n19271) );
  AND2_X1 U18626 ( .A1(n19414), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n15561) );
  AOI21_X1 U18627 ( .B1(n16316), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n15561), .ZN(n15306) );
  OAI21_X1 U18628 ( .B1(n16355), .B2(n19121), .A(n15306), .ZN(n15307) );
  AOI21_X1 U18629 ( .B1(n19271), .B2(n16363), .A(n15307), .ZN(n15308) );
  OAI211_X1 U18630 ( .C1(n15569), .C2(n19417), .A(n15309), .B(n15308), .ZN(
        P2_U3002) );
  XNOR2_X1 U18631 ( .A(n9832), .B(n15311), .ZN(n15635) );
  AND2_X1 U18632 ( .A1(n19414), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n15626) );
  OAI22_X1 U18633 ( .A1(n19425), .A2(n10181), .B1(n16355), .B2(n19194), .ZN(
        n15312) );
  AOI211_X1 U18634 ( .C1(n19195), .C2(n16363), .A(n15626), .B(n15312), .ZN(
        n15318) );
  NAND2_X1 U18635 ( .A1(n15314), .A2(n15313), .ZN(n15315) );
  XNOR2_X1 U18636 ( .A(n15316), .B(n15315), .ZN(n15633) );
  NAND2_X1 U18637 ( .A1(n15633), .A2(n19421), .ZN(n15317) );
  OAI211_X1 U18638 ( .C1(n15635), .C2(n19417), .A(n15318), .B(n15317), .ZN(
        P2_U3009) );
  INV_X1 U18639 ( .A(n15319), .ZN(n15323) );
  OAI21_X1 U18640 ( .B1(n15321), .B2(n16412), .A(n15320), .ZN(n15322) );
  OAI21_X1 U18641 ( .B1(n15326), .B2(n15325), .A(n15324), .ZN(n15327) );
  INV_X1 U18642 ( .A(n15327), .ZN(n15329) );
  INV_X1 U18643 ( .A(n15331), .ZN(n15332) );
  OAI21_X1 U18644 ( .B1(n15333), .B2(n16425), .A(n15332), .ZN(P2_U3016) );
  INV_X1 U18645 ( .A(n16197), .ZN(n15335) );
  AOI21_X1 U18646 ( .B1(n16387), .B2(n15335), .A(n15334), .ZN(n15338) );
  NAND3_X1 U18647 ( .A1(n15336), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n10961), .ZN(n15337) );
  OAI211_X1 U18648 ( .C1(n15339), .C2(n10961), .A(n15338), .B(n15337), .ZN(
        n15341) );
  NOR2_X1 U18649 ( .A1(n16186), .A2(n16413), .ZN(n15340) );
  AOI211_X1 U18650 ( .C1(n15342), .C2(n16390), .A(n15341), .B(n15340), .ZN(
        n15343) );
  OAI21_X1 U18651 ( .B1(n15344), .B2(n16425), .A(n15343), .ZN(P2_U3018) );
  OAI21_X1 U18652 ( .B1(n16412), .B2(n16211), .A(n15345), .ZN(n15347) );
  AOI211_X1 U18653 ( .C1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n15348), .A(
        n15347), .B(n15346), .ZN(n15349) );
  OAI21_X1 U18654 ( .B1(n16204), .B2(n16413), .A(n15349), .ZN(n15350) );
  AOI21_X1 U18655 ( .B1(n15351), .B2(n16390), .A(n15350), .ZN(n15352) );
  OAI21_X1 U18656 ( .B1(n15353), .B2(n16425), .A(n15352), .ZN(P2_U3019) );
  INV_X1 U18657 ( .A(n15354), .ZN(n16213) );
  AOI21_X1 U18658 ( .B1(n16387), .B2(n16213), .A(n15355), .ZN(n15358) );
  NOR2_X1 U18659 ( .A1(n15378), .A2(n15377), .ZN(n15367) );
  OAI211_X1 U18660 ( .C1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n15367), .B(n15356), .ZN(
        n15357) );
  OAI211_X1 U18661 ( .C1(n15376), .C2(n15359), .A(n15358), .B(n15357), .ZN(
        n15362) );
  NOR2_X1 U18662 ( .A1(n15360), .A2(n16416), .ZN(n15361) );
  AOI211_X1 U18663 ( .C1(n16214), .C2(n16406), .A(n15362), .B(n15361), .ZN(
        n15363) );
  OAI21_X1 U18664 ( .B1(n15364), .B2(n16425), .A(n15363), .ZN(P2_U3020) );
  OAI21_X1 U18665 ( .B1(n16412), .B2(n16225), .A(n15365), .ZN(n15366) );
  AOI21_X1 U18666 ( .B1(n15367), .B2(n15369), .A(n15366), .ZN(n15368) );
  OAI21_X1 U18667 ( .B1(n15376), .B2(n15369), .A(n15368), .ZN(n15373) );
  NOR3_X1 U18668 ( .A1(n15371), .A2(n15370), .A3(n16416), .ZN(n15372) );
  AOI211_X1 U18669 ( .C1(n16227), .C2(n16406), .A(n15373), .B(n15372), .ZN(
        n15374) );
  OAI21_X1 U18670 ( .B1(n15375), .B2(n16425), .A(n15374), .ZN(P2_U3021) );
  AOI21_X1 U18671 ( .B1(n15378), .B2(n15377), .A(n15376), .ZN(n15379) );
  AOI211_X1 U18672 ( .C1(n16387), .C2(n16237), .A(n15380), .B(n15379), .ZN(
        n15381) );
  OAI21_X1 U18673 ( .B1(n16239), .B2(n16413), .A(n15381), .ZN(n15382) );
  AOI21_X1 U18674 ( .B1(n15383), .B2(n16390), .A(n15382), .ZN(n15384) );
  OAI21_X1 U18675 ( .B1(n15385), .B2(n16425), .A(n15384), .ZN(P2_U3022) );
  NAND2_X1 U18676 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15597), .ZN(
        n16377) );
  INV_X1 U18677 ( .A(n15580), .ZN(n15387) );
  NOR2_X1 U18678 ( .A1(n16377), .A2(n15387), .ZN(n15543) );
  INV_X1 U18679 ( .A(n15388), .ZN(n15528) );
  NAND2_X1 U18680 ( .A1(n15543), .A2(n15528), .ZN(n15512) );
  INV_X1 U18681 ( .A(n15389), .ZN(n15390) );
  OR3_X1 U18682 ( .A1(n15512), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n15390), .ZN(n15426) );
  INV_X1 U18683 ( .A(n15391), .ZN(n15392) );
  NAND2_X1 U18684 ( .A1(n16420), .A2(n15392), .ZN(n15393) );
  NAND2_X1 U18685 ( .A1(n15579), .A2(n15393), .ZN(n15425) );
  INV_X1 U18686 ( .A(n15425), .ZN(n15394) );
  AND2_X1 U18687 ( .A1(n15426), .A2(n15394), .ZN(n15409) );
  NOR2_X1 U18688 ( .A1(n15409), .A2(n15395), .ZN(n15401) );
  XNOR2_X1 U18689 ( .A(n15395), .B(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15396) );
  NAND3_X1 U18690 ( .A1(n15397), .A2(n15396), .A3(n15597), .ZN(n15398) );
  OAI211_X1 U18691 ( .C1(n16412), .C2(n16259), .A(n15399), .B(n15398), .ZN(
        n15400) );
  AOI211_X1 U18692 ( .C1(n16262), .C2(n16406), .A(n15401), .B(n15400), .ZN(
        n15404) );
  NAND2_X1 U18693 ( .A1(n15402), .A2(n16390), .ZN(n15403) );
  OAI211_X1 U18694 ( .C1(n15405), .C2(n16425), .A(n15404), .B(n15403), .ZN(
        P2_U3023) );
  OR2_X1 U18695 ( .A1(n15407), .A2(n15406), .ZN(n15411) );
  INV_X1 U18696 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15410) );
  NAND2_X1 U18697 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19414), .ZN(n15408) );
  OAI221_X1 U18698 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n15411), 
        .C1(n15410), .C2(n15409), .A(n15408), .ZN(n15417) );
  NOR2_X1 U18699 ( .A1(n15413), .A2(n15412), .ZN(n15414) );
  OR2_X1 U18700 ( .A1(n15415), .A2(n15414), .ZN(n16279) );
  NOR2_X1 U18701 ( .A1(n16412), .A2(n16279), .ZN(n15416) );
  AOI211_X1 U18702 ( .C1(n15418), .C2(n16406), .A(n15417), .B(n15416), .ZN(
        n15422) );
  NAND3_X1 U18703 ( .A1(n15420), .A2(n16390), .A3(n15419), .ZN(n15421) );
  OAI211_X1 U18704 ( .C1(n15423), .C2(n16425), .A(n15422), .B(n15421), .ZN(
        P2_U3024) );
  AOI21_X1 U18705 ( .B1(n15425), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15424), .ZN(n15427) );
  OAI211_X1 U18706 ( .C1(n15428), .C2(n16413), .A(n15427), .B(n15426), .ZN(
        n15431) );
  NOR2_X1 U18707 ( .A1(n15429), .A2(n16412), .ZN(n15430) );
  AOI211_X1 U18708 ( .C1(n15432), .C2(n16390), .A(n15431), .B(n15430), .ZN(
        n15433) );
  OAI21_X1 U18709 ( .B1(n15434), .B2(n16425), .A(n15433), .ZN(P2_U3025) );
  NAND2_X1 U18710 ( .A1(n15435), .A2(n16407), .ZN(n15451) );
  NAND2_X1 U18711 ( .A1(n15437), .A2(n15436), .ZN(n15444) );
  NOR3_X1 U18712 ( .A1(n15512), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n15438), .ZN(n15453) );
  NAND3_X1 U18713 ( .A1(n15579), .A2(n15478), .A3(n15467), .ZN(n15441) );
  NOR2_X1 U18714 ( .A1(n15439), .A2(n16420), .ZN(n15578) );
  INV_X1 U18715 ( .A(n15578), .ZN(n15440) );
  NAND2_X1 U18716 ( .A1(n15441), .A2(n15440), .ZN(n15466) );
  OAI21_X1 U18717 ( .B1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n16386), .A(
        n15466), .ZN(n15455) );
  OAI21_X1 U18718 ( .B1(n15453), .B2(n15455), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15443) );
  OAI211_X1 U18719 ( .C1(n15512), .C2(n15444), .A(n15443), .B(n15442), .ZN(
        n15448) );
  NOR2_X1 U18720 ( .A1(n15090), .A2(n15445), .ZN(n15446) );
  OR2_X1 U18721 ( .A1(n14854), .A2(n15446), .ZN(n19044) );
  NOR2_X1 U18722 ( .A1(n19044), .A2(n16412), .ZN(n15447) );
  AOI211_X1 U18723 ( .C1(n15449), .C2(n16406), .A(n15448), .B(n15447), .ZN(
        n15450) );
  OAI211_X1 U18724 ( .C1(n15452), .C2(n16416), .A(n15451), .B(n15450), .ZN(
        P2_U3026) );
  NAND2_X1 U18725 ( .A1(n19058), .A2(n16387), .ZN(n15457) );
  AOI211_X1 U18726 ( .C1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15455), .A(
        n15454), .B(n15453), .ZN(n15456) );
  OAI211_X1 U18727 ( .C1(n19056), .C2(n16413), .A(n15457), .B(n15456), .ZN(
        n15458) );
  AOI21_X1 U18728 ( .B1(n15459), .B2(n16390), .A(n15458), .ZN(n15460) );
  OAI21_X1 U18729 ( .B1(n15461), .B2(n16425), .A(n15460), .ZN(P2_U3027) );
  NAND2_X1 U18730 ( .A1(n15463), .A2(n15462), .ZN(n15464) );
  NAND2_X1 U18731 ( .A1(n15465), .A2(n15464), .ZN(n19068) );
  NOR2_X1 U18732 ( .A1(n19068), .A2(n16412), .ZN(n15474) );
  INV_X1 U18733 ( .A(n15466), .ZN(n15471) );
  INV_X1 U18734 ( .A(n15467), .ZN(n15468) );
  NOR3_X1 U18735 ( .A1(n15512), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15468), .ZN(n15469) );
  AOI211_X1 U18736 ( .C1(n15471), .C2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15470), .B(n15469), .ZN(n15472) );
  OAI21_X1 U18737 ( .B1(n16413), .B2(n19067), .A(n15472), .ZN(n15473) );
  AOI211_X1 U18738 ( .C1(n15475), .C2(n16390), .A(n15474), .B(n15473), .ZN(
        n15476) );
  OAI21_X1 U18739 ( .B1(n15477), .B2(n16425), .A(n15476), .ZN(P2_U3028) );
  AOI21_X1 U18740 ( .B1(n15579), .B2(n15478), .A(n15578), .ZN(n15509) );
  OAI21_X1 U18741 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n16386), .A(
        n15502), .ZN(n15490) );
  OAI22_X1 U18742 ( .A1(n15513), .A2(n16416), .B1(n15482), .B2(n15512), .ZN(
        n15496) );
  NAND3_X1 U18743 ( .A1(n15496), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n15483), .ZN(n15487) );
  INV_X1 U18744 ( .A(n15484), .ZN(n19080) );
  AOI21_X1 U18745 ( .B1(n19080), .B2(n16406), .A(n15485), .ZN(n15486) );
  OAI211_X1 U18746 ( .C1(n16412), .C2(n15488), .A(n15487), .B(n15486), .ZN(
        n15489) );
  AOI21_X1 U18747 ( .B1(n15490), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n15489), .ZN(n15491) );
  OAI21_X1 U18748 ( .B1(n15492), .B2(n16425), .A(n15491), .ZN(P2_U3029) );
  NOR2_X1 U18749 ( .A1(n19302), .A2(n16412), .ZN(n15495) );
  OAI21_X1 U18750 ( .B1(n19262), .B2(n16413), .A(n15493), .ZN(n15494) );
  AOI211_X1 U18751 ( .C1(n15496), .C2(n15501), .A(n15495), .B(n15494), .ZN(
        n15500) );
  NAND3_X1 U18752 ( .A1(n15498), .A2(n15497), .A3(n16407), .ZN(n15499) );
  OAI211_X1 U18753 ( .C1(n15502), .C2(n15501), .A(n15500), .B(n15499), .ZN(
        P2_U3030) );
  NAND2_X1 U18754 ( .A1(n15504), .A2(n15503), .ZN(n15505) );
  XNOR2_X1 U18755 ( .A(n15506), .B(n15505), .ZN(n16297) );
  XOR2_X1 U18756 ( .A(n15507), .B(n15508), .Z(n19307) );
  NAND2_X1 U18757 ( .A1(n19093), .A2(n16406), .ZN(n15511) );
  AOI22_X1 U18758 ( .A1(n15509), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B1(
        P2_REIP_REG_15__SCAN_IN), .B2(n19414), .ZN(n15510) );
  OAI211_X1 U18759 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15512), .A(
        n15511), .B(n15510), .ZN(n15516) );
  OAI21_X1 U18760 ( .B1(n15514), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15513), .ZN(n16298) );
  NOR2_X1 U18761 ( .A1(n16298), .A2(n16416), .ZN(n15515) );
  AOI211_X1 U18762 ( .C1(n16387), .C2(n19307), .A(n15516), .B(n15515), .ZN(
        n15517) );
  OAI21_X1 U18763 ( .B1(n16297), .B2(n16425), .A(n15517), .ZN(P2_U3031) );
  OAI21_X1 U18764 ( .B1(n15556), .B2(n15545), .A(n15518), .ZN(n15520) );
  NAND2_X1 U18765 ( .A1(n15520), .A2(n15519), .ZN(n16303) );
  AND2_X1 U18766 ( .A1(n15540), .A2(n15521), .ZN(n15522) );
  OR2_X1 U18767 ( .A1(n15522), .A2(n15507), .ZN(n19311) );
  INV_X1 U18768 ( .A(n19311), .ZN(n15532) );
  NAND2_X1 U18769 ( .A1(n14097), .A2(n15523), .ZN(n15524) );
  NAND2_X1 U18770 ( .A1(n9855), .A2(n15524), .ZN(n19268) );
  AOI21_X1 U18771 ( .B1(n15525), .B2(n16420), .A(n15595), .ZN(n15526) );
  INV_X1 U18772 ( .A(n15526), .ZN(n15566) );
  INV_X1 U18773 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n20076) );
  OAI21_X1 U18774 ( .B1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n15544), .A(
        n15543), .ZN(n15527) );
  OAI22_X1 U18775 ( .A1(n19176), .A2(n20076), .B1(n15528), .B2(n15527), .ZN(
        n15529) );
  AOI21_X1 U18776 ( .B1(n15566), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n15529), .ZN(n15530) );
  OAI21_X1 U18777 ( .B1(n16413), .B2(n19268), .A(n15530), .ZN(n15531) );
  AOI21_X1 U18778 ( .B1(n15532), .B2(n16387), .A(n15531), .ZN(n15538) );
  NAND2_X1 U18779 ( .A1(n15534), .A2(n15533), .ZN(n15535) );
  XNOR2_X1 U18780 ( .A(n15536), .B(n15535), .ZN(n16304) );
  NAND2_X1 U18781 ( .A1(n16304), .A2(n16407), .ZN(n15537) );
  OAI211_X1 U18782 ( .C1(n16303), .C2(n16416), .A(n15538), .B(n15537), .ZN(
        P2_U3032) );
  OAI21_X1 U18783 ( .B1(n15539), .B2(n15541), .A(n15540), .ZN(n19313) );
  NOR2_X1 U18784 ( .A1(n19313), .A2(n16412), .ZN(n15551) );
  INV_X1 U18785 ( .A(n15542), .ZN(n15548) );
  INV_X1 U18786 ( .A(n15543), .ZN(n15564) );
  AOI211_X1 U18787 ( .C1(n15546), .C2(n15545), .A(n15544), .B(n15564), .ZN(
        n15547) );
  AOI211_X1 U18788 ( .C1(n15566), .C2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n15548), .B(n15547), .ZN(n15549) );
  OAI21_X1 U18789 ( .B1(n16413), .B2(n19113), .A(n15549), .ZN(n15550) );
  AOI211_X1 U18790 ( .C1(n15552), .C2(n16407), .A(n15551), .B(n15550), .ZN(
        n15553) );
  OAI21_X1 U18791 ( .B1(n15554), .B2(n16416), .A(n15553), .ZN(P2_U3033) );
  NAND3_X1 U18792 ( .A1(n15556), .A2(n16390), .A3(n15555), .ZN(n15568) );
  INV_X1 U18793 ( .A(n15557), .ZN(n15558) );
  NOR2_X1 U18794 ( .A1(n15558), .A2(n15559), .ZN(n15560) );
  NOR2_X1 U18795 ( .A1(n15539), .A2(n15560), .ZN(n19314) );
  AOI21_X1 U18796 ( .B1(n16387), .B2(n19314), .A(n15561), .ZN(n15563) );
  NAND2_X1 U18797 ( .A1(n19271), .A2(n16406), .ZN(n15562) );
  OAI211_X1 U18798 ( .C1(n15564), .C2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15563), .B(n15562), .ZN(n15565) );
  AOI21_X1 U18799 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n15566), .A(
        n15565), .ZN(n15567) );
  OAI211_X1 U18800 ( .C1(n15569), .C2(n16425), .A(n15568), .B(n15567), .ZN(
        P2_U3034) );
  OAI21_X1 U18801 ( .B1(n16327), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n15570), .ZN(n16312) );
  AND2_X1 U18802 ( .A1(n16318), .A2(n16319), .ZN(n15572) );
  NAND2_X1 U18803 ( .A1(n15571), .A2(n15572), .ZN(n15577) );
  INV_X1 U18804 ( .A(n15573), .ZN(n15574) );
  NOR2_X1 U18805 ( .A1(n15575), .A2(n15574), .ZN(n15576) );
  XNOR2_X1 U18806 ( .A(n15577), .B(n15576), .ZN(n16311) );
  AOI21_X1 U18807 ( .B1(n15579), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15578), .ZN(n16380) );
  INV_X1 U18808 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n20071) );
  NOR2_X1 U18809 ( .A1(n20071), .A2(n19176), .ZN(n15583) );
  INV_X1 U18810 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15581) );
  AOI211_X1 U18811 ( .C1(n16329), .C2(n15581), .A(n15580), .B(n16377), .ZN(
        n15582) );
  AOI211_X1 U18812 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n16380), .A(
        n15583), .B(n15582), .ZN(n15589) );
  NOR2_X1 U18813 ( .A1(n15585), .A2(n15584), .ZN(n15586) );
  OR2_X1 U18814 ( .A1(n15558), .A2(n15586), .ZN(n19318) );
  NOR2_X1 U18815 ( .A1(n16412), .A2(n19318), .ZN(n15587) );
  AOI21_X1 U18816 ( .B1(n19135), .B2(n16406), .A(n15587), .ZN(n15588) );
  OAI211_X1 U18817 ( .C1(n16311), .C2(n16425), .A(n15589), .B(n15588), .ZN(
        n15590) );
  INV_X1 U18818 ( .A(n15590), .ZN(n15591) );
  OAI21_X1 U18819 ( .B1(n16312), .B2(n16416), .A(n15591), .ZN(P2_U3035) );
  OAI21_X1 U18820 ( .B1(n15220), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n16328), .ZN(n16336) );
  AND2_X1 U18821 ( .A1(n15592), .A2(n16318), .ZN(n15593) );
  XNOR2_X1 U18822 ( .A(n9861), .B(n15593), .ZN(n16335) );
  INV_X1 U18823 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15596) );
  NOR2_X1 U18824 ( .A1(n11142), .A2(n19176), .ZN(n15594) );
  AOI221_X1 U18825 ( .B1(n15597), .B2(n15596), .C1(n15595), .C2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n15594), .ZN(n15603) );
  OR2_X1 U18826 ( .A1(n15598), .A2(n9972), .ZN(n15600) );
  NAND2_X1 U18827 ( .A1(n15600), .A2(n15599), .ZN(n19323) );
  NOR2_X1 U18828 ( .A1(n16412), .A2(n19323), .ZN(n15601) );
  AOI21_X1 U18829 ( .B1(n19159), .B2(n16406), .A(n15601), .ZN(n15602) );
  OAI211_X1 U18830 ( .C1(n16335), .C2(n16425), .A(n15603), .B(n15602), .ZN(
        n15604) );
  INV_X1 U18831 ( .A(n15604), .ZN(n15605) );
  OAI21_X1 U18832 ( .B1(n16336), .B2(n16416), .A(n15605), .ZN(P2_U3037) );
  OAI21_X1 U18833 ( .B1(n15607), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n15606), .ZN(n16372) );
  AOI21_X1 U18834 ( .B1(n16420), .B2(n16393), .A(n15608), .ZN(n16385) );
  NOR2_X1 U18835 ( .A1(n16394), .A2(n16393), .ZN(n15610) );
  INV_X1 U18836 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n20063) );
  NOR2_X1 U18837 ( .A1(n20063), .A2(n19176), .ZN(n15609) );
  AOI21_X1 U18838 ( .B1(n16392), .B2(n15610), .A(n15609), .ZN(n15611) );
  OAI21_X1 U18839 ( .B1(n16385), .B2(n16392), .A(n15611), .ZN(n15615) );
  XNOR2_X1 U18840 ( .A(n15613), .B(n15612), .ZN(n19330) );
  NOR2_X1 U18841 ( .A1(n19330), .A2(n16412), .ZN(n15614) );
  AOI211_X1 U18842 ( .C1(n19185), .C2(n16406), .A(n15615), .B(n15614), .ZN(
        n15620) );
  INV_X1 U18843 ( .A(n15617), .ZN(n15618) );
  XNOR2_X1 U18844 ( .A(n15616), .B(n15618), .ZN(n16367) );
  NAND2_X1 U18845 ( .A1(n16367), .A2(n16407), .ZN(n15619) );
  OAI211_X1 U18846 ( .C1(n16372), .C2(n16416), .A(n15620), .B(n15619), .ZN(
        P2_U3040) );
  AOI221_X1 U18847 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C1(n15622), .C2(n15629), .A(
        n15621), .ZN(n15632) );
  OAI21_X1 U18848 ( .B1(n14104), .B2(n15624), .A(n15623), .ZN(n19337) );
  INV_X1 U18849 ( .A(n19337), .ZN(n15625) );
  NAND2_X1 U18850 ( .A1(n15625), .A2(n16387), .ZN(n15628) );
  AOI21_X1 U18851 ( .B1(n19195), .B2(n16406), .A(n15626), .ZN(n15627) );
  OAI211_X1 U18852 ( .C1(n15630), .C2(n15629), .A(n15628), .B(n15627), .ZN(
        n15631) );
  AOI211_X1 U18853 ( .C1(n15633), .C2(n16390), .A(n15632), .B(n15631), .ZN(
        n15634) );
  OAI21_X1 U18854 ( .B1(n15635), .B2(n16425), .A(n15634), .ZN(P2_U3041) );
  INV_X1 U18855 ( .A(n16449), .ZN(n15667) );
  INV_X1 U18856 ( .A(n15636), .ZN(n15637) );
  NOR2_X1 U18857 ( .A1(n15638), .A2(n15637), .ZN(n15654) );
  INV_X1 U18858 ( .A(n16437), .ZN(n15639) );
  MUX2_X1 U18859 ( .A(n15654), .B(n15639), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n15640) );
  OAI21_X1 U18860 ( .B1(n19245), .B2(n15667), .A(n15640), .ZN(n16455) );
  NAND2_X1 U18861 ( .A1(n15641), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20121) );
  INV_X1 U18862 ( .A(n20121), .ZN(n15668) );
  INV_X1 U18863 ( .A(n19256), .ZN(n15642) );
  AOI22_X1 U18864 ( .A1(n19192), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n15642), .B2(n19182), .ZN(n15646) );
  AOI222_X1 U18865 ( .A1(n16455), .A2(n20029), .B1(n15643), .B2(n15668), .C1(
        P2_STATE2_REG_1__SCAN_IN), .C2(n15646), .ZN(n15645) );
  NAND2_X1 U18866 ( .A1(n20123), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15644) );
  OAI21_X1 U18867 ( .B1(n15645), .B2(n20123), .A(n15644), .ZN(P2_U3601) );
  NOR2_X1 U18868 ( .A1(n15646), .A2(n16479), .ZN(n15669) );
  INV_X1 U18869 ( .A(n15669), .ZN(n15656) );
  OAI211_X1 U18870 ( .C1(n19256), .C2(n15648), .A(n19182), .B(n15647), .ZN(
        n19236) );
  OAI21_X1 U18871 ( .B1(n19182), .B2(n15649), .A(n19236), .ZN(n15670) );
  INV_X1 U18872 ( .A(n20029), .ZN(n20128) );
  NOR2_X1 U18873 ( .A1(n10639), .A2(n15650), .ZN(n15653) );
  NAND2_X1 U18874 ( .A1(n16437), .A2(n15651), .ZN(n15652) );
  OAI21_X1 U18875 ( .B1(n15654), .B2(n15653), .A(n15652), .ZN(n15655) );
  AOI21_X1 U18876 ( .B1(n19227), .B2(n16449), .A(n15655), .ZN(n16452) );
  OAI222_X1 U18877 ( .A1(n20130), .A2(n20121), .B1(n15656), .B2(n15670), .C1(
        n20128), .C2(n16452), .ZN(n15657) );
  MUX2_X1 U18878 ( .A(n15657), .B(n15662), .S(n20123), .Z(P2_U3600) );
  OR2_X1 U18879 ( .A1(n15658), .A2(n16430), .ZN(n16439) );
  INV_X1 U18880 ( .A(n15659), .ZN(n15660) );
  NAND2_X1 U18881 ( .A1(n15660), .A2(n16432), .ZN(n16442) );
  NAND2_X1 U18882 ( .A1(n16440), .A2(n16442), .ZN(n15665) );
  NOR2_X1 U18883 ( .A1(n15661), .A2(n11096), .ZN(n16445) );
  NAND2_X1 U18884 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n15662), .ZN(
        n16435) );
  NAND2_X1 U18885 ( .A1(n16437), .A2(n16435), .ZN(n16443) );
  NOR2_X1 U18886 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n15662), .ZN(
        n15663) );
  OAI22_X1 U18887 ( .A1(n16445), .A2(n15665), .B1(n16443), .B2(n15663), .ZN(
        n15664) );
  AOI21_X1 U18888 ( .B1(n16439), .B2(n15665), .A(n15664), .ZN(n15666) );
  OAI21_X1 U18889 ( .B1(n10596), .B2(n15667), .A(n15666), .ZN(n16434) );
  AOI222_X1 U18890 ( .A1(n20029), .A2(n16434), .B1(n15670), .B2(n15669), .C1(
        n15668), .C2(n19611), .ZN(n15672) );
  NAND2_X1 U18891 ( .A1(n20123), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15671) );
  OAI21_X1 U18892 ( .B1(n15672), .B2(n20123), .A(n15671), .ZN(P2_U3599) );
  INV_X1 U18893 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n17040) );
  INV_X1 U18894 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n17038) );
  INV_X1 U18895 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16802) );
  NAND2_X1 U18896 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n17101), .ZN(n17097) );
  INV_X1 U18897 ( .A(n17088), .ZN(n17091) );
  NAND2_X1 U18898 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n17091), .ZN(n15746) );
  INV_X1 U18899 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n16704) );
  INV_X1 U18900 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16718) );
  AOI22_X1 U18901 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17285), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15673) );
  OAI21_X1 U18902 ( .B1(n11479), .B2(n17347), .A(n15673), .ZN(n15682) );
  AOI22_X1 U18903 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17310), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15680) );
  AOI22_X1 U18904 ( .A1(n17292), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15674) );
  OAI21_X1 U18905 ( .B1(n11447), .B2(n17254), .A(n15674), .ZN(n15678) );
  AOI22_X1 U18906 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15676) );
  AOI22_X1 U18907 ( .A1(n17304), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17309), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15675) );
  OAI211_X1 U18908 ( .C1(n17237), .C2(n17252), .A(n15676), .B(n15675), .ZN(
        n15677) );
  AOI211_X1 U18909 ( .C1(n17293), .C2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n15678), .B(n15677), .ZN(n15679) );
  OAI211_X1 U18910 ( .C1(n11498), .C2(n17153), .A(n15680), .B(n15679), .ZN(
        n15681) );
  AOI211_X1 U18911 ( .C1(n17291), .C2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A(
        n15682), .B(n15681), .ZN(n17089) );
  AOI22_X1 U18912 ( .A1(n17309), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n15683) );
  OAI21_X1 U18913 ( .B1(n11523), .B2(n17290), .A(n15683), .ZN(n15691) );
  AOI22_X1 U18914 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17310), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15689) );
  INV_X1 U18915 ( .A(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17289) );
  OAI22_X1 U18916 ( .A1(n11447), .A2(n17287), .B1(n17312), .B2(n17289), .ZN(
        n15688) );
  AOI22_X1 U18917 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17285), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15686) );
  AOI22_X1 U18918 ( .A1(n17304), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n15685) );
  AOI22_X1 U18919 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n15684) );
  NAND3_X1 U18920 ( .A1(n15686), .A2(n15685), .A3(n15684), .ZN(n15687) );
  OAI211_X1 U18921 ( .C1(n11479), .C2(n17359), .A(n15689), .B(n9985), .ZN(
        n15690) );
  AOI211_X1 U18922 ( .C1(n17291), .C2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A(
        n15691), .B(n15690), .ZN(n17098) );
  AOI22_X1 U18923 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n17291), .B1(
        P3_INSTQUEUE_REG_4__0__SCAN_IN), .B2(n9811), .ZN(n15701) );
  AOI22_X1 U18924 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n17325), .B1(
        P3_INSTQUEUE_REG_0__0__SCAN_IN), .B2(n17211), .ZN(n15693) );
  AOI22_X1 U18925 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17200), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15692) );
  OAI211_X1 U18926 ( .C1(n11448), .C2(n18396), .A(n15693), .B(n15692), .ZN(
        n15699) );
  AOI22_X1 U18927 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n17309), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15697) );
  AOI22_X1 U18928 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15696) );
  AOI22_X1 U18929 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17292), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15695) );
  NAND2_X1 U18930 ( .A1(n11444), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n15694) );
  NAND4_X1 U18931 ( .A1(n15697), .A2(n15696), .A3(n15695), .A4(n15694), .ZN(
        n15698) );
  AOI211_X1 U18932 ( .C1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .C2(n17268), .A(
        n15699), .B(n15698), .ZN(n15700) );
  OAI211_X1 U18933 ( .C1(n17197), .C2(n18373), .A(n15701), .B(n15700), .ZN(
        n17103) );
  AOI22_X1 U18934 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15711) );
  INV_X1 U18935 ( .A(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17218) );
  AOI22_X1 U18936 ( .A1(n11497), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15703) );
  AOI22_X1 U18937 ( .A1(n17313), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15702) );
  OAI211_X1 U18938 ( .C1(n11448), .C2(n17218), .A(n15703), .B(n15702), .ZN(
        n15709) );
  AOI22_X1 U18939 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17285), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15707) );
  AOI22_X1 U18940 ( .A1(n17309), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15706) );
  AOI22_X1 U18941 ( .A1(n17310), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17292), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15705) );
  NAND2_X1 U18942 ( .A1(n17268), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n15704) );
  NAND4_X1 U18943 ( .A1(n15707), .A2(n15706), .A3(n15705), .A4(n15704), .ZN(
        n15708) );
  OAI211_X1 U18944 ( .C1(n11479), .C2(n17063), .A(n15711), .B(n15710), .ZN(
        n17104) );
  NAND2_X1 U18945 ( .A1(n17103), .A2(n17104), .ZN(n17102) );
  NOR2_X1 U18946 ( .A1(n17098), .A2(n17102), .ZN(n17094) );
  AOI22_X1 U18947 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n15721) );
  AOI22_X1 U18948 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15720) );
  AOI22_X1 U18949 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17292), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15719) );
  OAI22_X1 U18950 ( .A1(n17197), .A2(n17272), .B1(n11467), .B2(n15712), .ZN(
        n15718) );
  AOI22_X1 U18951 ( .A1(n17304), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15716) );
  AOI22_X1 U18952 ( .A1(n17313), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17309), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15715) );
  AOI22_X1 U18953 ( .A1(n9811), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15714) );
  NAND2_X1 U18954 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n15713) );
  NAND4_X1 U18955 ( .A1(n15716), .A2(n15715), .A3(n15714), .A4(n15713), .ZN(
        n15717) );
  NAND4_X1 U18956 ( .A1(n15721), .A2(n15720), .A3(n15719), .A4(n9987), .ZN(
        n17093) );
  NAND2_X1 U18957 ( .A1(n17094), .A2(n17093), .ZN(n17092) );
  NOR2_X1 U18958 ( .A1(n17089), .A2(n17092), .ZN(n17086) );
  AOI22_X1 U18959 ( .A1(n17310), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15731) );
  INV_X1 U18960 ( .A(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17242) );
  AOI22_X1 U18961 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17200), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15723) );
  AOI22_X1 U18962 ( .A1(n17309), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15722) );
  OAI211_X1 U18963 ( .C1(n11467), .C2(n17242), .A(n15723), .B(n15722), .ZN(
        n15729) );
  AOI22_X1 U18964 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15727) );
  AOI22_X1 U18965 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15726) );
  NAND2_X1 U18966 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n15724) );
  NAND4_X1 U18967 ( .A1(n15727), .A2(n15726), .A3(n15725), .A4(n15724), .ZN(
        n15728) );
  AOI211_X1 U18968 ( .C1(n17292), .C2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n15729), .B(n15728), .ZN(n15730) );
  OAI211_X1 U18969 ( .C1(n17170), .C2(n15732), .A(n15731), .B(n15730), .ZN(
        n17085) );
  NAND2_X1 U18970 ( .A1(n17086), .A2(n17085), .ZN(n17084) );
  AOI22_X1 U18971 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15743) );
  INV_X1 U18972 ( .A(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15735) );
  AOI22_X1 U18973 ( .A1(n17313), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17309), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15734) );
  AOI22_X1 U18974 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15733) );
  OAI211_X1 U18975 ( .C1(n11467), .C2(n15735), .A(n15734), .B(n15733), .ZN(
        n15741) );
  AOI22_X1 U18976 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17291), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15739) );
  AOI22_X1 U18977 ( .A1(n17304), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15738) );
  NAND2_X1 U18978 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n15736) );
  NAND4_X1 U18979 ( .A1(n15739), .A2(n15738), .A3(n15737), .A4(n15736), .ZN(
        n15740) );
  AOI211_X1 U18980 ( .C1(n17292), .C2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n15741), .B(n15740), .ZN(n15742) );
  OAI211_X1 U18981 ( .C1(n11447), .C2(n15744), .A(n15743), .B(n15742), .ZN(
        n17079) );
  XNOR2_X1 U18982 ( .A(n17084), .B(n17079), .ZN(n17380) );
  AOI22_X1 U18983 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17083), .B1(n17361), 
        .B2(n17380), .ZN(n15745) );
  OAI21_X1 U18984 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n15746), .A(n15745), .ZN(
        P3_U2675) );
  INV_X1 U18985 ( .A(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17123) );
  AOI22_X1 U18986 ( .A1(n17285), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15747) );
  OAI21_X1 U18987 ( .B1(n9888), .B2(n17123), .A(n15747), .ZN(n15756) );
  AOI22_X1 U18988 ( .A1(n17313), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15754) );
  OAI22_X1 U18989 ( .A1(n11448), .A2(n17339), .B1(n17197), .B2(n17122), .ZN(
        n15752) );
  AOI22_X1 U18990 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15750) );
  AOI22_X1 U18991 ( .A1(n17309), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15749) );
  AOI22_X1 U18992 ( .A1(n17292), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15748) );
  NAND3_X1 U18993 ( .A1(n15750), .A2(n15749), .A3(n15748), .ZN(n15751) );
  AOI211_X1 U18994 ( .C1(n11444), .C2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A(
        n15752), .B(n15751), .ZN(n15753) );
  OAI211_X1 U18995 ( .C1(n11498), .C2(n17124), .A(n15754), .B(n15753), .ZN(
        n15755) );
  AOI211_X1 U18996 ( .C1(n17245), .C2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A(
        n15756), .B(n15755), .ZN(n17459) );
  AND2_X1 U18997 ( .A1(n17358), .A2(n15757), .ZN(n17246) );
  AOI22_X1 U18998 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17246), .B1(n15758), 
        .B2(n16875), .ZN(n15759) );
  OAI21_X1 U18999 ( .B1(n17459), .B2(n17358), .A(n15759), .ZN(P3_U2690) );
  NOR2_X1 U19000 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18942), .ZN(
        n18370) );
  NOR2_X1 U19001 ( .A1(n18996), .A2(n18965), .ZN(n18844) );
  NAND2_X1 U19002 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18844), .ZN(n18941) );
  INV_X1 U19003 ( .A(n18941), .ZN(n18847) );
  INV_X1 U19004 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16981) );
  NAND2_X1 U19005 ( .A1(n15775), .A2(n16981), .ZN(n15760) );
  OR2_X1 U19006 ( .A1(n17310), .A2(n15760), .ZN(n18321) );
  INV_X1 U19007 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n19005) );
  NAND2_X1 U19008 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n16981), .ZN(n18954) );
  INV_X1 U19009 ( .A(n18486), .ZN(n18536) );
  INV_X1 U19010 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18322) );
  NOR2_X1 U19011 ( .A1(n18322), .A2(n18941), .ZN(n15773) );
  AOI211_X1 U19012 ( .C1(n18847), .C2(n18321), .A(n18536), .B(n15773), .ZN(
        n15761) );
  NOR2_X1 U19013 ( .A1(n18370), .A2(n15761), .ZN(n15763) );
  NOR2_X1 U19014 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n16625) );
  NAND2_X1 U19015 ( .A1(P3_STATEBS16_REG_SCAN_IN), .A2(n16625), .ZN(n18627) );
  INV_X1 U19016 ( .A(n15761), .ZN(n18327) );
  OAI21_X1 U19017 ( .B1(n19005), .B2(n18965), .A(n18942), .ZN(n18990) );
  INV_X1 U19018 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n16655) );
  NOR2_X1 U19019 ( .A1(n18965), .A2(n16655), .ZN(n18845) );
  INV_X1 U19020 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18800) );
  OAI22_X1 U19021 ( .A1(n18990), .A2(n18845), .B1(n18942), .B2(n18800), .ZN(
        n15766) );
  NAND3_X1 U19022 ( .A1(n18801), .A2(n18327), .A3(n15766), .ZN(n15762) );
  OAI221_X1 U19023 ( .B1(n18801), .B2(n15763), .C1(n18801), .C2(n18627), .A(
        n15762), .ZN(P3_U2864) );
  NAND2_X1 U19024 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18511) );
  NOR2_X1 U19025 ( .A1(n18990), .A2(n18845), .ZN(n15765) );
  INV_X1 U19026 ( .A(n15763), .ZN(n15764) );
  AOI221_X1 U19027 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18511), .C1(n15765), 
        .C2(n18511), .A(n15764), .ZN(n18326) );
  INV_X1 U19028 ( .A(n18627), .ZN(n18679) );
  OAI221_X1 U19029 ( .B1(n18679), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n18679), .C2(n15766), .A(n18327), .ZN(n18324) );
  AOI22_X1 U19030 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18326), .B1(
        n18324), .B2(n18330), .ZN(P3_U2865) );
  INV_X1 U19031 ( .A(n18988), .ZN(n18994) );
  NOR2_X1 U19032 ( .A1(n18994), .A2(n18777), .ZN(n15772) );
  INV_X1 U19033 ( .A(n18777), .ZN(n16631) );
  INV_X1 U19034 ( .A(n15767), .ZN(n15774) );
  OAI21_X1 U19035 ( .B1(n15774), .B2(n16648), .A(n16647), .ZN(n15768) );
  NAND3_X1 U19036 ( .A1(n16631), .A2(n18988), .A3(n15768), .ZN(n15870) );
  OAI211_X1 U19037 ( .C1(n18782), .C2(n15770), .A(n15769), .B(n15870), .ZN(
        n15771) );
  AOI21_X1 U19038 ( .B1(n15772), .B2(n17515), .A(n15771), .ZN(n18816) );
  NOR2_X1 U19039 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18942), .ZN(n18335) );
  INV_X1 U19040 ( .A(n18973), .ZN(n18970) );
  INV_X1 U19041 ( .A(n18944), .ZN(n19006) );
  AOI211_X1 U19042 ( .C1(n15775), .C2(n16981), .A(n15774), .B(n16648), .ZN(
        n18784) );
  NAND3_X1 U19043 ( .A1(n18970), .A2(n19006), .A3(n18784), .ZN(n15776) );
  OAI21_X1 U19044 ( .B1(n18970), .B2(n16981), .A(n15776), .ZN(P3_U3284) );
  NAND2_X1 U19045 ( .A1(n15778), .A2(n15777), .ZN(n15779) );
  XNOR2_X1 U19046 ( .A(n15779), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16533) );
  AOI21_X1 U19047 ( .B1(n18268), .B2(n15781), .A(n15780), .ZN(n15784) );
  INV_X1 U19048 ( .A(n17997), .ZN(n17634) );
  OAI21_X1 U19049 ( .B1(n16510), .B2(n17634), .A(n17484), .ZN(n15782) );
  OAI22_X1 U19050 ( .A1(n16528), .A2(n18304), .B1(n18311), .B2(n15782), .ZN(
        n15843) );
  INV_X1 U19051 ( .A(n15843), .ZN(n15783) );
  OAI21_X1 U19052 ( .B1(n18308), .B2(n15784), .A(n15783), .ZN(n15785) );
  AOI22_X1 U19053 ( .A1(n9822), .A2(P3_REIP_REG_29__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15785), .ZN(n15790) );
  INV_X1 U19054 ( .A(n17633), .ZN(n17998) );
  AOI22_X1 U19055 ( .A1(n18231), .A2(n17998), .B1(n18229), .B2(n17997), .ZN(
        n15787) );
  AOI21_X1 U19056 ( .B1(n15787), .B2(n15786), .A(n10081), .ZN(n15842) );
  NAND3_X1 U19057 ( .A1(n15788), .A2(n15842), .A3(n16519), .ZN(n15789) );
  OAI211_X1 U19058 ( .C1(n16533), .C2(n18237), .A(n15790), .B(n15789), .ZN(
        P3_U2833) );
  AOI22_X1 U19059 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19252), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19242), .ZN(n15800) );
  AOI22_X1 U19060 ( .A1(n15791), .A2(n19241), .B1(P2_EBX_REG_22__SCAN_IN), 
        .B2(n19250), .ZN(n15799) );
  OAI22_X1 U19061 ( .A1(n16268), .A2(n19246), .B1(n16279), .B2(n19207), .ZN(
        n15792) );
  INV_X1 U19062 ( .A(n15792), .ZN(n15798) );
  NAND2_X1 U19063 ( .A1(n15793), .A2(n19037), .ZN(n15794) );
  NAND2_X1 U19064 ( .A1(n15794), .A2(n19182), .ZN(n15795) );
  OAI211_X1 U19065 ( .C1(n15796), .C2(n15795), .A(n19198), .B(n16155), .ZN(
        n15797) );
  NAND4_X1 U19066 ( .A1(n15800), .A2(n15799), .A3(n15798), .A4(n15797), .ZN(
        P2_U2833) );
  INV_X1 U19067 ( .A(n15801), .ZN(n15813) );
  AOI211_X1 U19068 ( .C1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n15803), .A(
        n20843), .B(n15802), .ZN(n15809) );
  INV_X1 U19069 ( .A(n15809), .ZN(n15807) );
  INV_X1 U19070 ( .A(n15804), .ZN(n15806) );
  OAI211_X1 U19071 ( .C1(n20791), .C2(n15807), .A(n15806), .B(n15805), .ZN(
        n15808) );
  OAI21_X1 U19072 ( .B1(n15809), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n15808), .ZN(n15810) );
  AOI222_X1 U19073 ( .A1(n12753), .A2(n15811), .B1(n12753), .B2(n15810), .C1(
        n15811), .C2(n15810), .ZN(n15812) );
  AOI222_X1 U19074 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n15813), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15812), .C1(n15813), 
        .C2(n15812), .ZN(n15814) );
  NAND2_X1 U19075 ( .A1(n15814), .A2(n20371), .ZN(n15823) );
  OAI21_X1 U19076 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n15815), .ZN(n15818) );
  AND4_X1 U19077 ( .A1(n15818), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n15817), 
        .A4(n15816), .ZN(n15821) );
  INV_X1 U19078 ( .A(n15819), .ZN(n15820) );
  NAND4_X1 U19079 ( .A1(n15823), .A2(n15822), .A3(n15821), .A4(n15820), .ZN(
        n15831) );
  NAND2_X1 U19080 ( .A1(n15824), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n15830) );
  NOR3_X1 U19081 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20991), .A3(n21064), 
        .ZN(n15827) );
  OAI22_X1 U19082 ( .A1(n15828), .A2(n15827), .B1(n15826), .B2(n15825), .ZN(
        n16150) );
  AOI21_X1 U19083 ( .B1(n15831), .B2(n16145), .A(n16150), .ZN(n16147) );
  AOI211_X1 U19084 ( .C1(n15831), .C2(n15830), .A(n15829), .B(n16147), .ZN(
        n15837) );
  AOI21_X1 U19085 ( .B1(n16146), .B2(n20991), .A(n15832), .ZN(n16148) );
  INV_X1 U19086 ( .A(n16147), .ZN(n15833) );
  OAI21_X1 U19087 ( .B1(n15835), .B2(n15834), .A(n15833), .ZN(n15836) );
  AOI22_X1 U19088 ( .A1(n15837), .A2(n16148), .B1(n21075), .B2(n15836), .ZN(
        P1_U3161) );
  NOR2_X1 U19089 ( .A1(n15839), .A2(n15838), .ZN(n15841) );
  XNOR2_X1 U19090 ( .A(n15841), .B(n15840), .ZN(n16516) );
  NOR2_X1 U19091 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16510), .ZN(
        n16512) );
  AOI22_X1 U19092 ( .A1(n9822), .A2(P3_REIP_REG_30__SCAN_IN), .B1(n16512), 
        .B2(n15842), .ZN(n15846) );
  OAI21_X1 U19093 ( .B1(n15844), .B2(n15843), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15845) );
  OAI211_X1 U19094 ( .C1(n16516), .C2(n18237), .A(n15846), .B(n15845), .ZN(
        P3_U2832) );
  NAND2_X1 U19095 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n16146), .ZN(n20998) );
  NAND3_X1 U19096 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .A3(n21007), .ZN(
        n15848) );
  INV_X1 U19097 ( .A(HOLD), .ZN(n21002) );
  OAI211_X1 U19098 ( .C1(n21007), .C2(n21002), .A(P1_STATE_REG_0__SCAN_IN), 
        .B(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n15847) );
  NAND4_X1 U19099 ( .A1(n21073), .A2(n20998), .A3(n15848), .A4(n15847), .ZN(
        P1_U3195) );
  AND2_X1 U19100 ( .A1(n15849), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR2_X1 U19101 ( .A1(n15851), .A2(n15850), .ZN(n15852) );
  XNOR2_X1 U19102 ( .A(n15852), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15980) );
  INV_X1 U19103 ( .A(n15853), .ZN(n15854) );
  AOI21_X1 U19104 ( .B1(n15856), .B2(n15855), .A(n15854), .ZN(n15967) );
  AOI22_X1 U19105 ( .A1(n15980), .A2(n20357), .B1(n16135), .B2(n15967), .ZN(
        n15863) );
  NAND2_X1 U19106 ( .A1(n16106), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15862) );
  OAI221_X1 U19107 ( .B1(n15858), .B2(n15857), .C1(n15858), .C2(n16097), .A(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15861) );
  NAND3_X1 U19108 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n15859), .A3(
        n12717), .ZN(n15860) );
  NAND4_X1 U19109 ( .A1(n15863), .A2(n15862), .A3(n15861), .A4(n15860), .ZN(
        P1_U3011) );
  NOR2_X1 U19110 ( .A1(n20047), .A2(n16491), .ZN(n20028) );
  AOI22_X1 U19111 ( .A1(n20148), .A2(n16491), .B1(n20028), .B2(n15864), .ZN(
        n15865) );
  AOI21_X1 U19112 ( .B1(n15865), .B2(n20158), .A(n16490), .ZN(P2_U3178) );
  INV_X1 U19113 ( .A(n16477), .ZN(n20170) );
  NAND2_X1 U19114 ( .A1(n16483), .A2(n15866), .ZN(n15867) );
  AOI221_X1 U19115 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16490), .C1(n20170), .C2(
        n16490), .A(n19974), .ZN(n20163) );
  INV_X1 U19116 ( .A(n20163), .ZN(n20164) );
  NOR2_X1 U19117 ( .A1(n16463), .A2(n20164), .ZN(P2_U3047) );
  NAND3_X1 U19118 ( .A1(n18339), .A2(n18336), .A3(n15868), .ZN(n15869) );
  NAND2_X1 U19119 ( .A1(n18366), .A2(n17514), .ZN(n17501) );
  INV_X1 U19120 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17587) );
  NAND2_X2 U19121 ( .A1(n17514), .A2(n17409), .ZN(n17494) );
  AOI22_X1 U19122 ( .A1(n17509), .A2(BUF2_REG_0__SCAN_IN), .B1(n17508), .B2(
        n17978), .ZN(n15871) );
  OAI221_X1 U19123 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17501), .C1(n17587), 
        .C2(n17514), .A(n15871), .ZN(P3_U2735) );
  INV_X1 U19124 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n21162) );
  NOR2_X1 U19125 ( .A1(n21162), .A2(n21378), .ZN(n15886) );
  AOI21_X1 U19126 ( .B1(n15877), .B2(n15886), .A(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n15876) );
  INV_X1 U19127 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n21397) );
  OAI22_X1 U19128 ( .A1(n15984), .A2(n20289), .B1(n21397), .B2(n20218), .ZN(
        n15872) );
  AOI21_X1 U19129 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20255), .A(
        n15872), .ZN(n15874) );
  AOI22_X1 U19130 ( .A1(n15981), .A2(n20245), .B1(n20272), .B2(n15967), .ZN(
        n15873) );
  OAI211_X1 U19131 ( .C1(n15876), .C2(n15875), .A(n15874), .B(n15873), .ZN(
        P1_U2820) );
  OAI21_X1 U19132 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(P1_REIP_REG_18__SCAN_IN), 
        .A(n15877), .ZN(n15885) );
  AOI22_X1 U19133 ( .A1(n15887), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_EBX_REG_19__SCAN_IN), .B2(n20292), .ZN(n15878) );
  OAI211_X1 U19134 ( .C1(n20288), .C2(n14642), .A(n15878), .B(n20256), .ZN(
        n15882) );
  OAI22_X1 U19135 ( .A1(n15880), .A2(n15960), .B1(n20295), .B2(n15879), .ZN(
        n15881) );
  AOI211_X1 U19136 ( .C1(n15883), .C2(n20254), .A(n15882), .B(n15881), .ZN(
        n15884) );
  OAI21_X1 U19137 ( .B1(n15886), .B2(n15885), .A(n15884), .ZN(P1_U2821) );
  INV_X1 U19138 ( .A(n20256), .ZN(n20270) );
  AOI22_X1 U19139 ( .A1(n15887), .A2(P1_REIP_REG_18__SCAN_IN), .B1(n20292), 
        .B2(P1_EBX_REG_18__SCAN_IN), .ZN(n15888) );
  OAI21_X1 U19140 ( .B1(n15889), .B2(n20289), .A(n15888), .ZN(n15890) );
  AOI211_X1 U19141 ( .C1(n20255), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n20270), .B(n15890), .ZN(n15892) );
  AOI22_X1 U19142 ( .A1(n15970), .A2(n20245), .B1(n20272), .B2(n15969), .ZN(
        n15891) );
  OAI211_X1 U19143 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n15893), .A(n15892), 
        .B(n15891), .ZN(P1_U2822) );
  OAI21_X1 U19144 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(P1_REIP_REG_16__SCAN_IN), 
        .A(n15894), .ZN(n15905) );
  NOR2_X1 U19145 ( .A1(n15895), .A2(n15951), .ZN(n15922) );
  AOI21_X1 U19146 ( .B1(n15898), .B2(n15897), .A(n15896), .ZN(n15899) );
  OR2_X1 U19147 ( .A1(n15899), .A2(n9958), .ZN(n15972) );
  INV_X1 U19148 ( .A(n15972), .ZN(n16071) );
  AOI22_X1 U19149 ( .A1(n15922), .A2(P1_REIP_REG_16__SCAN_IN), .B1(n20272), 
        .B2(n16071), .ZN(n15904) );
  NAND2_X1 U19150 ( .A1(n20255), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15900) );
  OAI211_X1 U19151 ( .C1(n20289), .C2(n15996), .A(n20256), .B(n15900), .ZN(
        n15902) );
  NOR2_X1 U19152 ( .A1(n15985), .A2(n15960), .ZN(n15901) );
  AOI211_X1 U19153 ( .C1(n20292), .C2(P1_EBX_REG_16__SCAN_IN), .A(n15902), .B(
        n15901), .ZN(n15903) );
  OAI211_X1 U19154 ( .C1(n15915), .C2(n15905), .A(n15904), .B(n15903), .ZN(
        P1_U2824) );
  INV_X1 U19155 ( .A(n15906), .ZN(n16079) );
  INV_X1 U19156 ( .A(n15907), .ZN(n15908) );
  AOI22_X1 U19157 ( .A1(n16079), .A2(n20272), .B1(n20254), .B2(n15908), .ZN(
        n15914) );
  NAND2_X1 U19158 ( .A1(n20292), .A2(P1_EBX_REG_15__SCAN_IN), .ZN(n15909) );
  OAI211_X1 U19159 ( .C1(n12339), .C2(n20288), .A(n15909), .B(n20256), .ZN(
        n15912) );
  NOR2_X1 U19160 ( .A1(n15910), .A2(n15960), .ZN(n15911) );
  AOI211_X1 U19161 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(n15922), .A(n15912), 
        .B(n15911), .ZN(n15913) );
  OAI211_X1 U19162 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(n15915), .A(n15914), 
        .B(n15913), .ZN(P1_U2825) );
  AOI22_X1 U19163 ( .A1(n20292), .A2(P1_EBX_REG_14__SCAN_IN), .B1(n20254), 
        .B2(n16003), .ZN(n15925) );
  OR2_X1 U19164 ( .A1(n15917), .A2(n15916), .ZN(n15918) );
  AND2_X1 U19165 ( .A1(n15919), .A2(n15918), .ZN(n16086) );
  AOI22_X1 U19166 ( .A1(n16086), .A2(n20272), .B1(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n20255), .ZN(n15924) );
  OR2_X1 U19167 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n15920), .ZN(n15921) );
  AOI22_X1 U19168 ( .A1(n16004), .A2(n20245), .B1(n15922), .B2(n15921), .ZN(
        n15923) );
  NAND4_X1 U19169 ( .A1(n15925), .A2(n15924), .A3(n15923), .A4(n20256), .ZN(
        P1_U2826) );
  NAND2_X1 U19170 ( .A1(n20250), .A2(n15926), .ZN(n15940) );
  NOR2_X1 U19171 ( .A1(n16092), .A2(n20295), .ZN(n15931) );
  AOI21_X1 U19172 ( .B1(n20255), .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n20270), .ZN(n15928) );
  NAND2_X1 U19173 ( .A1(n20292), .A2(P1_EBX_REG_13__SCAN_IN), .ZN(n15927) );
  OAI211_X1 U19174 ( .C1(n20289), .C2(n15929), .A(n15928), .B(n15927), .ZN(
        n15930) );
  AOI211_X1 U19175 ( .C1(n15932), .C2(n20245), .A(n15931), .B(n15930), .ZN(
        n15933) );
  OAI221_X1 U19176 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n15934), .C1(n21382), 
        .C2(n15940), .A(n15933), .ZN(P1_U2827) );
  AOI22_X1 U19177 ( .A1(n20292), .A2(P1_EBX_REG_12__SCAN_IN), .B1(n20254), 
        .B2(n16014), .ZN(n15945) );
  AND2_X1 U19178 ( .A1(n15936), .A2(n15935), .ZN(n15937) );
  NOR2_X1 U19179 ( .A1(n15938), .A2(n15937), .ZN(n16107) );
  AOI22_X1 U19180 ( .A1(n16107), .A2(n20272), .B1(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n20255), .ZN(n15944) );
  INV_X1 U19181 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n21349) );
  INV_X1 U19182 ( .A(n15939), .ZN(n15941) );
  AOI21_X1 U19183 ( .B1(n21349), .B2(n15941), .A(n15940), .ZN(n15942) );
  AOI21_X1 U19184 ( .B1(n16015), .B2(n20245), .A(n15942), .ZN(n15943) );
  NAND4_X1 U19185 ( .A1(n15945), .A2(n15944), .A3(n15943), .A4(n20256), .ZN(
        P1_U2828) );
  INV_X1 U19186 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15948) );
  INV_X1 U19187 ( .A(n16026), .ZN(n15946) );
  AOI21_X1 U19188 ( .B1(n20254), .B2(n15946), .A(n20270), .ZN(n15947) );
  OAI21_X1 U19189 ( .B1(n15948), .B2(n20288), .A(n15947), .ZN(n15950) );
  NOR2_X1 U19190 ( .A1(n16116), .A2(n20295), .ZN(n15949) );
  AOI211_X1 U19191 ( .C1(n20292), .C2(P1_EBX_REG_11__SCAN_IN), .A(n15950), .B(
        n15949), .ZN(n15954) );
  NOR2_X1 U19192 ( .A1(n15952), .A2(n15951), .ZN(n15964) );
  AOI22_X1 U19193 ( .A1(n16023), .A2(n20245), .B1(n15964), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n15953) );
  OAI211_X1 U19194 ( .C1(P1_REIP_REG_11__SCAN_IN), .C2(n15955), .A(n15954), 
        .B(n15953), .ZN(P1_U2829) );
  INV_X1 U19195 ( .A(n15956), .ZN(n15957) );
  AOI22_X1 U19196 ( .A1(n20292), .A2(P1_EBX_REG_10__SCAN_IN), .B1(n15957), 
        .B2(n20254), .ZN(n15966) );
  AOI21_X1 U19197 ( .B1(n20255), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n20270), .ZN(n15959) );
  NAND2_X1 U19198 ( .A1(n16123), .A2(n20272), .ZN(n15958) );
  OAI211_X1 U19199 ( .C1(n15961), .C2(n15960), .A(n15959), .B(n15958), .ZN(
        n15962) );
  AOI221_X1 U19200 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(n15964), .C1(n15963), 
        .C2(n15964), .A(n15962), .ZN(n15965) );
  NAND2_X1 U19201 ( .A1(n15966), .A2(n15965), .ZN(P1_U2830) );
  AOI22_X1 U19202 ( .A1(n15981), .A2(n20303), .B1(n13038), .B2(n15967), .ZN(
        n15968) );
  OAI21_X1 U19203 ( .B1(n20306), .B2(n21397), .A(n15968), .ZN(P1_U2852) );
  INV_X1 U19204 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n21120) );
  AOI22_X1 U19205 ( .A1(n15970), .A2(n20303), .B1(n13038), .B2(n15969), .ZN(
        n15971) );
  OAI21_X1 U19206 ( .B1(n20306), .B2(n21120), .A(n15971), .ZN(P1_U2854) );
  OAI22_X1 U19207 ( .A1(n15985), .A2(n15974), .B1(n15973), .B2(n15972), .ZN(
        n15975) );
  INV_X1 U19208 ( .A(n15975), .ZN(n15976) );
  OAI21_X1 U19209 ( .B1(n20306), .B2(n21197), .A(n15976), .ZN(P1_U2856) );
  INV_X1 U19210 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n15978) );
  AOI22_X1 U19211 ( .A1(n16004), .A2(n20303), .B1(n13038), .B2(n16086), .ZN(
        n15977) );
  OAI21_X1 U19212 ( .B1(n20306), .B2(n15978), .A(n15977), .ZN(P1_U2858) );
  INV_X1 U19213 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n21131) );
  AOI22_X1 U19214 ( .A1(n16015), .A2(n20303), .B1(n13038), .B2(n16107), .ZN(
        n15979) );
  OAI21_X1 U19215 ( .B1(n20306), .B2(n21131), .A(n15979), .ZN(P1_U2860) );
  AOI22_X1 U19216 ( .A1(n16027), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(
        n16106), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n15983) );
  AOI22_X1 U19217 ( .A1(n15981), .A2(n20374), .B1(n16034), .B2(n15980), .ZN(
        n15982) );
  OAI211_X1 U19218 ( .C1(n16031), .C2(n15984), .A(n15983), .B(n15982), .ZN(
        P1_U2979) );
  AOI22_X1 U19219 ( .A1(n16027), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n16106), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n15995) );
  INV_X1 U19220 ( .A(n15985), .ZN(n15993) );
  NAND2_X1 U19221 ( .A1(n15987), .A2(n15986), .ZN(n15989) );
  NAND2_X1 U19222 ( .A1(n15989), .A2(n15988), .ZN(n15992) );
  INV_X1 U19223 ( .A(n15990), .ZN(n15991) );
  XNOR2_X1 U19224 ( .A(n15992), .B(n15991), .ZN(n16074) );
  AOI22_X1 U19225 ( .A1(n15993), .A2(n20374), .B1(n16034), .B2(n16074), .ZN(
        n15994) );
  OAI211_X1 U19226 ( .C1(n16031), .C2(n15996), .A(n15995), .B(n15994), .ZN(
        P1_U2983) );
  OAI21_X1 U19227 ( .B1(n10119), .B2(n15998), .A(n15997), .ZN(n16000) );
  NAND2_X1 U19228 ( .A1(n16000), .A2(n15999), .ZN(n16002) );
  XNOR2_X1 U19229 ( .A(n14680), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16001) );
  XNOR2_X1 U19230 ( .A(n16002), .B(n16001), .ZN(n16091) );
  AOI22_X1 U19231 ( .A1(n16027), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n16106), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16006) );
  AOI22_X1 U19232 ( .A1(n16004), .A2(n20374), .B1(n16033), .B2(n16003), .ZN(
        n16005) );
  OAI211_X1 U19233 ( .C1(n16091), .C2(n20187), .A(n16006), .B(n16005), .ZN(
        P1_U2985) );
  INV_X1 U19234 ( .A(n16007), .ZN(n16008) );
  NOR2_X1 U19235 ( .A1(n16009), .A2(n16008), .ZN(n16013) );
  NAND2_X1 U19236 ( .A1(n16011), .A2(n16010), .ZN(n16012) );
  XNOR2_X1 U19237 ( .A(n16013), .B(n16012), .ZN(n16113) );
  AOI22_X1 U19238 ( .A1(n16027), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n16106), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16017) );
  AOI22_X1 U19239 ( .A1(n16015), .A2(n20374), .B1(n16033), .B2(n16014), .ZN(
        n16016) );
  OAI211_X1 U19240 ( .C1(n16113), .C2(n20187), .A(n16017), .B(n16016), .ZN(
        P1_U2987) );
  AOI22_X1 U19241 ( .A1(n16027), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n16106), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16025) );
  INV_X1 U19242 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16132) );
  NOR3_X1 U19243 ( .A1(n16019), .A2(n16132), .A3(n16018), .ZN(n16021) );
  NOR2_X1 U19244 ( .A1(n16021), .A2(n16020), .ZN(n16022) );
  XOR2_X1 U19245 ( .A(n12710), .B(n16022), .Z(n16118) );
  AOI22_X1 U19246 ( .A1(n16118), .A2(n16034), .B1(n20374), .B2(n16023), .ZN(
        n16024) );
  OAI211_X1 U19247 ( .C1(n16031), .C2(n16026), .A(n16025), .B(n16024), .ZN(
        P1_U2988) );
  AOI22_X1 U19248 ( .A1(n16027), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n16106), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16030) );
  AOI22_X1 U19249 ( .A1(n16028), .A2(n16034), .B1(n20374), .B2(n20237), .ZN(
        n16029) );
  OAI211_X1 U19250 ( .C1(n16031), .C2(n20228), .A(n16030), .B(n16029), .ZN(
        P1_U2992) );
  INV_X1 U19251 ( .A(n16032), .ZN(n16035) );
  AOI222_X1 U19252 ( .A1(n16035), .A2(n16034), .B1(n20253), .B2(n16033), .C1(
        n20265), .C2(n20374), .ZN(n16037) );
  OAI211_X1 U19253 ( .C1(n16039), .C2(n16038), .A(n16037), .B(n16036), .ZN(
        P1_U2994) );
  AOI22_X1 U19254 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n16106), .B1(n16041), 
        .B2(n16040), .ZN(n16046) );
  INV_X1 U19255 ( .A(n16042), .ZN(n16044) );
  AOI22_X1 U19256 ( .A1(n16044), .A2(n16135), .B1(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n16043), .ZN(n16045) );
  OAI211_X1 U19257 ( .C1(n16112), .C2(n16047), .A(n16046), .B(n16045), .ZN(
        P1_U3006) );
  INV_X1 U19258 ( .A(n16048), .ZN(n16051) );
  INV_X1 U19259 ( .A(n16049), .ZN(n16050) );
  AOI22_X1 U19260 ( .A1(n16051), .A2(n20357), .B1(n16135), .B2(n16050), .ZN(
        n16059) );
  INV_X1 U19261 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16056) );
  OAI21_X1 U19262 ( .B1(n16105), .B2(n16053), .A(n16052), .ZN(n16055) );
  NOR2_X1 U19263 ( .A1(n20369), .A2(n21413), .ZN(n16054) );
  AOI221_X1 U19264 ( .B1(n16057), .B2(n16056), .C1(n16055), .C2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A(n16054), .ZN(n16058) );
  NAND2_X1 U19265 ( .A1(n16059), .A2(n16058), .ZN(P1_U3007) );
  INV_X1 U19266 ( .A(n16060), .ZN(n16064) );
  NOR3_X1 U19267 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n16061), .A3(
        n16065), .ZN(n16062) );
  AOI211_X1 U19268 ( .C1(n16064), .C2(n16135), .A(n16063), .B(n16062), .ZN(
        n16069) );
  NOR2_X1 U19269 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n16065), .ZN(
        n16066) );
  OAI21_X1 U19270 ( .B1(n16067), .B2(n16066), .A(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16068) );
  OAI211_X1 U19271 ( .C1(n16070), .C2(n16112), .A(n16069), .B(n16068), .ZN(
        P1_U3009) );
  AOI22_X1 U19272 ( .A1(n16071), .A2(n16135), .B1(n16106), .B2(
        P1_REIP_REG_16__SCAN_IN), .ZN(n16076) );
  AOI21_X1 U19273 ( .B1(n16084), .B2(n16077), .A(n16072), .ZN(n16073) );
  AOI22_X1 U19274 ( .A1(n20357), .A2(n16074), .B1(n16080), .B2(n16073), .ZN(
        n16075) );
  OAI211_X1 U19275 ( .C1(n16085), .C2(n16077), .A(n16076), .B(n16075), .ZN(
        P1_U3015) );
  AOI21_X1 U19276 ( .B1(n16079), .B2(n16135), .A(n16078), .ZN(n16083) );
  AOI22_X1 U19277 ( .A1(n20357), .A2(n16081), .B1(n16080), .B2(n16084), .ZN(
        n16082) );
  OAI211_X1 U19278 ( .C1(n16085), .C2(n16084), .A(n16083), .B(n16082), .ZN(
        P1_U3016) );
  AOI22_X1 U19279 ( .A1(n16086), .A2(n16135), .B1(n16106), .B2(
        P1_REIP_REG_14__SCAN_IN), .ZN(n16090) );
  OAI222_X1 U19280 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16088), 
        .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16114), .C1(n16087), 
        .C2(n16096), .ZN(n16089) );
  OAI211_X1 U19281 ( .C1(n16091), .C2(n16112), .A(n16090), .B(n16089), .ZN(
        P1_U3017) );
  INV_X1 U19282 ( .A(n16092), .ZN(n16095) );
  INV_X1 U19283 ( .A(n16093), .ZN(n16094) );
  AOI222_X1 U19284 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n16106), .B1(n16135), 
        .B2(n16095), .C1(n20357), .C2(n16094), .ZN(n16099) );
  OAI21_X1 U19285 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16097), .A(
        n16096), .ZN(n16098) );
  OAI211_X1 U19286 ( .C1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n16100), .A(
        n16099), .B(n16098), .ZN(P1_U3018) );
  OAI21_X1 U19287 ( .B1(n16109), .B2(n20361), .A(n16101), .ZN(n16102) );
  AOI21_X1 U19288 ( .B1(n16104), .B2(n16103), .A(n16102), .ZN(n16120) );
  OAI21_X1 U19289 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16105), .A(
        n16120), .ZN(n16108) );
  AOI222_X1 U19290 ( .A1(n16108), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), 
        .B1(n16107), .B2(n16135), .C1(P1_REIP_REG_12__SCAN_IN), .C2(n16106), 
        .ZN(n16111) );
  NAND3_X1 U19291 ( .A1(n16109), .A2(n12703), .A3(n16114), .ZN(n16110) );
  OAI211_X1 U19292 ( .C1(n16113), .C2(n16112), .A(n16111), .B(n16110), .ZN(
        P1_U3019) );
  NAND2_X1 U19293 ( .A1(n16115), .A2(n16114), .ZN(n16121) );
  OAI22_X1 U19294 ( .A1(n16116), .A2(n20355), .B1(n21302), .B2(n20369), .ZN(
        n16117) );
  AOI21_X1 U19295 ( .B1(n20357), .B2(n16118), .A(n16117), .ZN(n16119) );
  OAI221_X1 U19296 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16121), 
        .C1(n12710), .C2(n16120), .A(n16119), .ZN(P1_U3020) );
  AOI21_X1 U19297 ( .B1(n16123), .B2(n16135), .A(n16122), .ZN(n16131) );
  AOI211_X1 U19298 ( .C1(n16132), .C2(n16126), .A(n16125), .B(n16124), .ZN(
        n16128) );
  AOI22_X1 U19299 ( .A1(n16129), .A2(n20357), .B1(n16128), .B2(n16127), .ZN(
        n16130) );
  OAI211_X1 U19300 ( .C1(n16133), .C2(n16132), .A(n16131), .B(n16130), .ZN(
        P1_U3021) );
  INV_X1 U19301 ( .A(n20215), .ZN(n16136) );
  AOI21_X1 U19302 ( .B1(n16136), .B2(n16135), .A(n16134), .ZN(n16144) );
  AOI22_X1 U19303 ( .A1(n16138), .A2(n20357), .B1(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n16137), .ZN(n16143) );
  OAI221_X1 U19304 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16141), .C2(n16140), .A(
        n16139), .ZN(n16142) );
  NAND3_X1 U19305 ( .A1(n16144), .A2(n16143), .A3(n16142), .ZN(P1_U3023) );
  AOI221_X1 U19306 ( .B1(n16146), .B2(P1_STATE2_REG_0__SCAN_IN), .C1(n20848), 
        .C2(n21075), .A(n16145), .ZN(n20988) );
  NOR2_X1 U19307 ( .A1(n16147), .A2(n21075), .ZN(n20990) );
  AOI21_X1 U19308 ( .B1(n20990), .B2(n16148), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n16149) );
  AOI221_X1 U19309 ( .B1(n20989), .B2(n16150), .C1(n20988), .C2(n16150), .A(
        n16149), .ZN(P1_U3162) );
  OAI21_X1 U19310 ( .B1(n20990), .B2(n20799), .A(n16151), .ZN(P1_U3466) );
  NAND2_X1 U19311 ( .A1(n19198), .A2(n19182), .ZN(n19255) );
  INV_X1 U19312 ( .A(n16152), .ZN(n16181) );
  INV_X1 U19313 ( .A(n16153), .ZN(n16208) );
  INV_X1 U19314 ( .A(n16154), .ZN(n16230) );
  INV_X1 U19315 ( .A(n16156), .ZN(n16256) );
  NAND2_X1 U19316 ( .A1(n19182), .A2(n16254), .ZN(n16242) );
  NAND2_X1 U19317 ( .A1(n16243), .A2(n16242), .ZN(n16241) );
  NAND2_X1 U19318 ( .A1(n19182), .A2(n16241), .ZN(n16229) );
  NAND2_X1 U19319 ( .A1(n16230), .A2(n16229), .ZN(n16228) );
  NAND2_X1 U19320 ( .A1(n16194), .A2(n16193), .ZN(n16192) );
  INV_X1 U19321 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n16162) );
  NAND2_X1 U19322 ( .A1(n16157), .A2(n19241), .ZN(n16161) );
  INV_X1 U19323 ( .A(n16158), .ZN(n16159) );
  NAND3_X1 U19324 ( .A1(n19409), .A2(P2_EBX_REG_31__SCAN_IN), .A3(n16159), 
        .ZN(n16160) );
  OAI211_X1 U19325 ( .C1(n19222), .C2(n16162), .A(n16161), .B(n16160), .ZN(
        n16163) );
  AOI21_X1 U19326 ( .B1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19252), .A(
        n16163), .ZN(n16166) );
  INV_X1 U19327 ( .A(n16164), .ZN(n19294) );
  AOI22_X1 U19328 ( .A1(n16260), .A2(n19226), .B1(n19239), .B2(n19294), .ZN(
        n16165) );
  OAI211_X1 U19329 ( .C1(n19255), .C2(n16170), .A(n16166), .B(n16165), .ZN(
        P2_U2824) );
  AOI22_X1 U19330 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19252), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19242), .ZN(n16175) );
  AOI22_X1 U19331 ( .A1(n16167), .A2(n19241), .B1(P2_EBX_REG_30__SCAN_IN), 
        .B2(n19250), .ZN(n16174) );
  INV_X1 U19332 ( .A(n15321), .ZN(n16168) );
  AOI22_X1 U19333 ( .A1(n16169), .A2(n19226), .B1(n16168), .B2(n19239), .ZN(
        n16173) );
  NAND4_X1 U19334 ( .A1(n16175), .A2(n16174), .A3(n16173), .A4(n16172), .ZN(
        P2_U2825) );
  AOI22_X1 U19335 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19252), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n19242), .ZN(n16185) );
  AOI22_X1 U19336 ( .A1(n16176), .A2(n19241), .B1(P2_EBX_REG_29__SCAN_IN), 
        .B2(n19250), .ZN(n16184) );
  AOI22_X1 U19337 ( .A1(n16178), .A2(n19226), .B1(n16177), .B2(n19239), .ZN(
        n16183) );
  OAI211_X1 U19338 ( .C1(n16181), .C2(n16180), .A(n19198), .B(n16179), .ZN(
        n16182) );
  NAND4_X1 U19339 ( .A1(n16185), .A2(n16184), .A3(n16183), .A4(n16182), .ZN(
        P2_U2826) );
  INV_X1 U19340 ( .A(n16186), .ZN(n16191) );
  AOI22_X1 U19341 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19252), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n19242), .ZN(n16188) );
  NAND2_X1 U19342 ( .A1(n19250), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n16187) );
  OAI211_X1 U19343 ( .C1(n16189), .C2(n19204), .A(n16188), .B(n16187), .ZN(
        n16190) );
  AOI21_X1 U19344 ( .B1(n16191), .B2(n19226), .A(n16190), .ZN(n16196) );
  OAI211_X1 U19345 ( .C1(n16194), .C2(n16193), .A(n19198), .B(n16192), .ZN(
        n16195) );
  OAI211_X1 U19346 ( .C1(n19207), .C2(n16197), .A(n16196), .B(n16195), .ZN(
        P2_U2827) );
  OAI22_X1 U19347 ( .A1(n16198), .A2(n19223), .B1(n20101), .B2(n19222), .ZN(
        n16201) );
  INV_X1 U19348 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n16199) );
  NOR2_X1 U19349 ( .A1(n19203), .A2(n16199), .ZN(n16200) );
  AOI211_X1 U19350 ( .C1(n16202), .C2(n19241), .A(n16201), .B(n16200), .ZN(
        n16203) );
  OAI21_X1 U19351 ( .B1(n16204), .B2(n19246), .A(n16203), .ZN(n16205) );
  INV_X1 U19352 ( .A(n16205), .ZN(n16210) );
  OAI211_X1 U19353 ( .C1(n16208), .C2(n16207), .A(n19198), .B(n16206), .ZN(
        n16209) );
  OAI211_X1 U19354 ( .C1(n19207), .C2(n16211), .A(n16210), .B(n16209), .ZN(
        P2_U2828) );
  AOI22_X1 U19355 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19252), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n19242), .ZN(n16221) );
  AOI22_X1 U19356 ( .A1(n16212), .A2(n19241), .B1(P2_EBX_REG_26__SCAN_IN), 
        .B2(n19250), .ZN(n16220) );
  AOI22_X1 U19357 ( .A1(n16214), .A2(n19226), .B1(n16213), .B2(n19239), .ZN(
        n16219) );
  OAI211_X1 U19358 ( .C1(n16217), .C2(n16216), .A(n19198), .B(n16215), .ZN(
        n16218) );
  NAND4_X1 U19359 ( .A1(n16221), .A2(n16220), .A3(n16219), .A4(n16218), .ZN(
        P2_U2829) );
  AOI22_X1 U19360 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19252), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n19242), .ZN(n16234) );
  OAI22_X1 U19361 ( .A1(n16223), .A2(n19204), .B1(n19203), .B2(n16222), .ZN(
        n16224) );
  INV_X1 U19362 ( .A(n16224), .ZN(n16233) );
  INV_X1 U19363 ( .A(n16225), .ZN(n16226) );
  AOI22_X1 U19364 ( .A1(n16227), .A2(n19226), .B1(n16226), .B2(n19239), .ZN(
        n16232) );
  OAI211_X1 U19365 ( .C1(n16230), .C2(n16229), .A(n19198), .B(n16228), .ZN(
        n16231) );
  NAND4_X1 U19366 ( .A1(n16234), .A2(n16233), .A3(n16232), .A4(n16231), .ZN(
        P2_U2830) );
  AOI22_X1 U19367 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19252), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19242), .ZN(n16247) );
  INV_X1 U19368 ( .A(n16235), .ZN(n16236) );
  AOI22_X1 U19369 ( .A1(n16236), .A2(n19241), .B1(P2_EBX_REG_24__SCAN_IN), 
        .B2(n19250), .ZN(n16246) );
  INV_X1 U19370 ( .A(n16237), .ZN(n16238) );
  OAI22_X1 U19371 ( .A1(n16239), .A2(n19246), .B1(n16238), .B2(n19207), .ZN(
        n16240) );
  INV_X1 U19372 ( .A(n16240), .ZN(n16245) );
  OAI211_X1 U19373 ( .C1(n16243), .C2(n16242), .A(n19198), .B(n16241), .ZN(
        n16244) );
  NAND4_X1 U19374 ( .A1(n16247), .A2(n16246), .A3(n16245), .A4(n16244), .ZN(
        P2_U2831) );
  NAND2_X1 U19375 ( .A1(n16248), .A2(n19241), .ZN(n16252) );
  OAI22_X1 U19376 ( .A1(n16249), .A2(n19223), .B1(n20092), .B2(n19222), .ZN(
        n16250) );
  AOI21_X1 U19377 ( .B1(n19250), .B2(P2_EBX_REG_23__SCAN_IN), .A(n16250), .ZN(
        n16251) );
  NAND2_X1 U19378 ( .A1(n16252), .A2(n16251), .ZN(n16253) );
  AOI21_X1 U19379 ( .B1(n16262), .B2(n19226), .A(n16253), .ZN(n16258) );
  OAI211_X1 U19380 ( .C1(n16256), .C2(n16255), .A(n19198), .B(n16254), .ZN(
        n16257) );
  OAI211_X1 U19381 ( .C1(n19207), .C2(n16259), .A(n16258), .B(n16257), .ZN(
        P2_U2832) );
  OAI22_X1 U19382 ( .A1(n14945), .A2(n16260), .B1(P2_EBX_REG_31__SCAN_IN), 
        .B2(n19293), .ZN(n16261) );
  INV_X1 U19383 ( .A(n16261), .ZN(P2_U2856) );
  INV_X1 U19384 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n16265) );
  AOI22_X1 U19385 ( .A1(n16263), .A2(n19278), .B1(n19293), .B2(n16262), .ZN(
        n16264) );
  OAI21_X1 U19386 ( .B1(n19293), .B2(n16265), .A(n16264), .ZN(P2_U2864) );
  AOI21_X1 U19387 ( .B1(n16266), .B2(n15001), .A(n13240), .ZN(n16281) );
  AOI22_X1 U19388 ( .A1(n16281), .A2(n19278), .B1(P2_EBX_REG_22__SCAN_IN), 
        .B2(n14945), .ZN(n16267) );
  OAI21_X1 U19389 ( .B1(n14945), .B2(n16268), .A(n16267), .ZN(P2_U2865) );
  AOI21_X1 U19390 ( .B1(n16271), .B2(n16270), .A(n16269), .ZN(n16286) );
  AOI22_X1 U19391 ( .A1(n16286), .A2(n19278), .B1(P2_EBX_REG_20__SCAN_IN), 
        .B2(n14945), .ZN(n16272) );
  OAI21_X1 U19392 ( .B1(n14945), .B2(n19043), .A(n16272), .ZN(P2_U2867) );
  INV_X1 U19393 ( .A(n16273), .ZN(n16276) );
  INV_X1 U19394 ( .A(n15013), .ZN(n16275) );
  AOI21_X1 U19395 ( .B1(n16276), .B2(n16275), .A(n16274), .ZN(n16293) );
  AOI22_X1 U19396 ( .A1(n16293), .A2(n19278), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n14945), .ZN(n16277) );
  OAI21_X1 U19397 ( .B1(n14945), .B2(n19067), .A(n16277), .ZN(P2_U2869) );
  AOI22_X1 U19398 ( .A1(n19298), .A2(n16278), .B1(n19356), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16284) );
  AOI22_X1 U19399 ( .A1(n19300), .A2(BUF2_REG_22__SCAN_IN), .B1(n19299), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n16283) );
  INV_X1 U19400 ( .A(n16279), .ZN(n16280) );
  AOI22_X1 U19401 ( .A1(n16281), .A2(n19342), .B1(n19357), .B2(n16280), .ZN(
        n16282) );
  NAND3_X1 U19402 ( .A1(n16284), .A2(n16283), .A3(n16282), .ZN(P2_U2897) );
  AOI22_X1 U19403 ( .A1(n19298), .A2(n16285), .B1(n19356), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16290) );
  AOI22_X1 U19404 ( .A1(n19300), .A2(BUF2_REG_20__SCAN_IN), .B1(n19299), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n16289) );
  INV_X1 U19405 ( .A(n19044), .ZN(n16287) );
  AOI22_X1 U19406 ( .A1(n16287), .A2(n19357), .B1(n19342), .B2(n16286), .ZN(
        n16288) );
  NAND3_X1 U19407 ( .A1(n16290), .A2(n16289), .A3(n16288), .ZN(P2_U2899) );
  AOI22_X1 U19408 ( .A1(n19298), .A2(n16291), .B1(n19356), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n16296) );
  AOI22_X1 U19409 ( .A1(n19300), .A2(BUF2_REG_18__SCAN_IN), .B1(n19299), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n16295) );
  INV_X1 U19410 ( .A(n19068), .ZN(n16292) );
  AOI22_X1 U19411 ( .A1(n19342), .A2(n16293), .B1(n16292), .B2(n19357), .ZN(
        n16294) );
  NAND3_X1 U19412 ( .A1(n16296), .A2(n16295), .A3(n16294), .ZN(P2_U2901) );
  AOI22_X1 U19413 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19414), .B1(n19413), 
        .B2(n19088), .ZN(n16302) );
  INV_X1 U19414 ( .A(n16297), .ZN(n16300) );
  INV_X1 U19415 ( .A(n16298), .ZN(n16299) );
  AOI222_X1 U19416 ( .A1(n16300), .A2(n16366), .B1(n16363), .B2(n19093), .C1(
        n19421), .C2(n16299), .ZN(n16301) );
  OAI211_X1 U19417 ( .C1(n19425), .C2(n19091), .A(n16302), .B(n16301), .ZN(
        P2_U2999) );
  AOI22_X1 U19418 ( .A1(n16316), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19414), .ZN(n16309) );
  OR2_X1 U19419 ( .A1(n16303), .A2(n16371), .ZN(n16306) );
  NAND2_X1 U19420 ( .A1(n16304), .A2(n16366), .ZN(n16305) );
  OAI211_X1 U19421 ( .C1(n19416), .C2(n19268), .A(n16306), .B(n16305), .ZN(
        n16307) );
  INV_X1 U19422 ( .A(n16307), .ZN(n16308) );
  OAI211_X1 U19423 ( .C1(n16355), .C2(n19099), .A(n16309), .B(n16308), .ZN(
        P2_U3000) );
  AOI22_X1 U19424 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19414), .B1(n19413), 
        .B2(n16310), .ZN(n16315) );
  OAI22_X1 U19425 ( .A1(n16312), .A2(n16371), .B1(n16311), .B2(n19417), .ZN(
        n16313) );
  AOI21_X1 U19426 ( .B1(n16363), .B2(n19135), .A(n16313), .ZN(n16314) );
  OAI211_X1 U19427 ( .C1(n19425), .C2(n19141), .A(n16315), .B(n16314), .ZN(
        P2_U3003) );
  AOI22_X1 U19428 ( .A1(n16316), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19414), .ZN(n16332) );
  NAND2_X1 U19429 ( .A1(n16317), .A2(n16318), .ZN(n16323) );
  INV_X1 U19430 ( .A(n16319), .ZN(n16320) );
  NOR2_X1 U19431 ( .A1(n16321), .A2(n16320), .ZN(n16322) );
  XNOR2_X1 U19432 ( .A(n16323), .B(n16322), .ZN(n16384) );
  INV_X1 U19433 ( .A(n16384), .ZN(n16330) );
  INV_X1 U19434 ( .A(n16324), .ZN(n16325) );
  AOI21_X1 U19435 ( .B1(n16326), .B2(n13977), .A(n16325), .ZN(n19277) );
  AOI21_X1 U19436 ( .B1(n16329), .B2(n16328), .A(n16327), .ZN(n16381) );
  AOI222_X1 U19437 ( .A1(n16330), .A2(n16366), .B1(n16363), .B2(n19277), .C1(
        n19421), .C2(n16381), .ZN(n16331) );
  OAI211_X1 U19438 ( .C1(n16355), .C2(n16333), .A(n16332), .B(n16331), .ZN(
        P2_U3004) );
  AOI22_X1 U19439 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19414), .B1(n19413), 
        .B2(n16334), .ZN(n16339) );
  OAI22_X1 U19440 ( .A1(n16336), .A2(n16371), .B1(n19417), .B2(n16335), .ZN(
        n16337) );
  AOI21_X1 U19441 ( .B1(n16363), .B2(n19159), .A(n16337), .ZN(n16338) );
  OAI211_X1 U19442 ( .C1(n19425), .C2(n19153), .A(n16339), .B(n16338), .ZN(
        P2_U3005) );
  AOI22_X1 U19443 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19414), .B1(n19413), 
        .B2(n16340), .ZN(n16350) );
  AOI21_X1 U19444 ( .B1(n16342), .B2(n16341), .A(n9900), .ZN(n16391) );
  NAND2_X1 U19445 ( .A1(n16344), .A2(n16343), .ZN(n16348) );
  AND2_X1 U19446 ( .A1(n16346), .A2(n16345), .ZN(n16360) );
  NAND2_X1 U19447 ( .A1(n16360), .A2(n16357), .ZN(n16362) );
  NAND2_X1 U19448 ( .A1(n16362), .A2(n16358), .ZN(n16347) );
  XOR2_X1 U19449 ( .A(n16348), .B(n16347), .Z(n16389) );
  INV_X1 U19450 ( .A(n19288), .ZN(n16388) );
  AOI222_X1 U19451 ( .A1(n16391), .A2(n19421), .B1(n16366), .B2(n16389), .C1(
        n16363), .C2(n16388), .ZN(n16349) );
  OAI211_X1 U19452 ( .C1(n19425), .C2(n16351), .A(n16350), .B(n16349), .ZN(
        P2_U3006) );
  XNOR2_X1 U19453 ( .A(n16352), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16353) );
  XNOR2_X1 U19454 ( .A(n16354), .B(n16353), .ZN(n16411) );
  OAI22_X1 U19455 ( .A1(n19425), .A2(n10182), .B1(n16355), .B2(n19168), .ZN(
        n16356) );
  AOI21_X1 U19456 ( .B1(P2_REIP_REG_7__SCAN_IN), .B2(n19414), .A(n16356), .ZN(
        n16365) );
  INV_X1 U19457 ( .A(n16358), .ZN(n16361) );
  AND2_X1 U19458 ( .A1(n16358), .A2(n16357), .ZN(n16359) );
  OAI22_X1 U19459 ( .A1(n16362), .A2(n16361), .B1(n16360), .B2(n16359), .ZN(
        n16408) );
  INV_X1 U19460 ( .A(n19171), .ZN(n16405) );
  AOI22_X1 U19461 ( .A1(n16408), .A2(n16366), .B1(n16363), .B2(n16405), .ZN(
        n16364) );
  OAI211_X1 U19462 ( .C1(n16371), .C2(n16411), .A(n16365), .B(n16364), .ZN(
        P2_U3007) );
  AOI22_X1 U19463 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n19414), .B1(n19413), 
        .B2(n19184), .ZN(n16375) );
  NAND2_X1 U19464 ( .A1(n16367), .A2(n16366), .ZN(n16370) );
  OR2_X1 U19465 ( .A1(n16368), .A2(n19416), .ZN(n16369) );
  OAI211_X1 U19466 ( .C1(n16372), .C2(n16371), .A(n16370), .B(n16369), .ZN(
        n16373) );
  INV_X1 U19467 ( .A(n16373), .ZN(n16374) );
  OAI211_X1 U19468 ( .C1(n19425), .C2(n19177), .A(n16375), .B(n16374), .ZN(
        P2_U3008) );
  INV_X1 U19469 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n20069) );
  NOR2_X1 U19470 ( .A1(n20069), .A2(n19176), .ZN(n16379) );
  XNOR2_X1 U19471 ( .A(n15599), .B(n16376), .ZN(n19321) );
  OAI22_X1 U19472 ( .A1(n16377), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n19321), .B2(n16412), .ZN(n16378) );
  AOI211_X1 U19473 ( .C1(n16380), .C2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n16379), .B(n16378), .ZN(n16383) );
  AOI22_X1 U19474 ( .A1(n16381), .A2(n16390), .B1(n16406), .B2(n19277), .ZN(
        n16382) );
  OAI211_X1 U19475 ( .C1(n16384), .C2(n16425), .A(n16383), .B(n16382), .ZN(
        P2_U3036) );
  OAI21_X1 U19476 ( .B1(n16386), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n16385), .ZN(n16403) );
  AOI22_X1 U19477 ( .A1(n16403), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n16387), .B2(n19324), .ZN(n16399) );
  AOI222_X1 U19478 ( .A1(n16391), .A2(n16390), .B1(n16407), .B2(n16389), .C1(
        n16406), .C2(n16388), .ZN(n16398) );
  NAND2_X1 U19479 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19414), .ZN(n16397) );
  NOR3_X1 U19480 ( .A1(n16394), .A2(n16393), .A3(n16392), .ZN(n16404) );
  OAI221_X1 U19481 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C1(n11076), .C2(n16395), .A(
        n16404), .ZN(n16396) );
  NAND4_X1 U19482 ( .A1(n16399), .A2(n16398), .A3(n16397), .A4(n16396), .ZN(
        P2_U3038) );
  OAI21_X1 U19483 ( .B1(n16401), .B2(n16400), .A(n14923), .ZN(n19329) );
  OAI22_X1 U19484 ( .A1(n19329), .A2(n16412), .B1(n20065), .B2(n19176), .ZN(
        n16402) );
  AOI221_X1 U19485 ( .B1(n16404), .B2(n11076), .C1(n16403), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16402), .ZN(n16410) );
  AOI22_X1 U19486 ( .A1(n16408), .A2(n16407), .B1(n16406), .B2(n16405), .ZN(
        n16409) );
  OAI211_X1 U19487 ( .C1(n16416), .C2(n16411), .A(n16410), .B(n16409), .ZN(
        P2_U3039) );
  OAI22_X1 U19488 ( .A1(n19245), .A2(n16413), .B1(n16412), .B2(n19237), .ZN(
        n16419) );
  INV_X1 U19489 ( .A(n16414), .ZN(n16415) );
  OAI22_X1 U19490 ( .A1(n16417), .A2(n16421), .B1(n16416), .B2(n16415), .ZN(
        n16418) );
  AOI211_X1 U19491 ( .C1(n16421), .C2(n16420), .A(n16419), .B(n16418), .ZN(
        n16423) );
  OAI211_X1 U19492 ( .C1(n16425), .C2(n16424), .A(n16423), .B(n16422), .ZN(
        P2_U3046) );
  OAI22_X1 U19493 ( .A1(n16431), .A2(n16428), .B1(n16427), .B2(n16426), .ZN(
        n16429) );
  AOI21_X1 U19494 ( .B1(n16431), .B2(n16430), .A(n16429), .ZN(n20171) );
  NAND2_X1 U19495 ( .A1(n16474), .A2(n16432), .ZN(n16433) );
  OAI21_X1 U19496 ( .B1(n16434), .B2(n16474), .A(n16433), .ZN(n16470) );
  OR2_X1 U19497 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n16470), .ZN(
        n16461) );
  INV_X1 U19498 ( .A(n16435), .ZN(n16436) );
  AND2_X1 U19499 ( .A1(n16437), .A2(n16436), .ZN(n16438) );
  OAI21_X1 U19500 ( .B1(n16439), .B2(n16438), .A(n16442), .ZN(n16441) );
  NAND2_X1 U19501 ( .A1(n16441), .A2(n16440), .ZN(n16447) );
  OAI211_X1 U19502 ( .C1(n16445), .C2(n9814), .A(n16443), .B(n16442), .ZN(
        n16446) );
  MUX2_X1 U19503 ( .A(n16447), .B(n16446), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n16448) );
  AOI21_X1 U19504 ( .B1(n13821), .B2(n16449), .A(n16448), .ZN(n20120) );
  MUX2_X1 U19505 ( .A(n20120), .B(n10444), .S(n16474), .Z(n16471) );
  INV_X1 U19506 ( .A(n16471), .ZN(n16459) );
  INV_X1 U19507 ( .A(n16474), .ZN(n16454) );
  OAI21_X1 U19508 ( .B1(n20165), .B2(n16455), .A(n16450), .ZN(n16451) );
  NAND2_X1 U19509 ( .A1(n16452), .A2(n16451), .ZN(n16453) );
  OAI211_X1 U19510 ( .C1(n16455), .C2(n19829), .A(n16454), .B(n16453), .ZN(
        n16456) );
  AOI21_X1 U19511 ( .B1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n16461), .A(
        n16456), .ZN(n16458) );
  NOR2_X1 U19512 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n16471), .ZN(
        n16457) );
  OAI22_X1 U19513 ( .A1(n16459), .A2(n20140), .B1(n16458), .B2(n16457), .ZN(
        n16460) );
  OAI21_X1 U19514 ( .B1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n16461), .A(
        n16460), .ZN(n16462) );
  AOI22_X1 U19515 ( .A1(n16464), .A2(n19437), .B1(n16463), .B2(n16462), .ZN(
        n16469) );
  INV_X1 U19516 ( .A(n16465), .ZN(n16468) );
  OAI21_X1 U19517 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n16466), .ZN(n16467) );
  NAND4_X1 U19518 ( .A1(n20171), .A2(n16469), .A3(n16468), .A4(n16467), .ZN(
        n16473) );
  NOR2_X1 U19519 ( .A1(n16471), .A2(n16470), .ZN(n16472) );
  AOI211_X1 U19520 ( .C1(n16474), .C2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n16473), .B(n16472), .ZN(n16489) );
  NOR2_X1 U19521 ( .A1(n16491), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20030) );
  AND2_X1 U19522 ( .A1(n20047), .A2(n20030), .ZN(n16476) );
  AOI211_X1 U19523 ( .C1(n16490), .C2(n16477), .A(n16476), .B(n16475), .ZN(
        n16487) );
  NAND2_X1 U19524 ( .A1(n16478), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n16481) );
  AOI21_X1 U19525 ( .B1(n16489), .B2(n16479), .A(n16491), .ZN(n16480) );
  AOI211_X1 U19526 ( .C1(n16482), .C2(n11017), .A(n16481), .B(n16480), .ZN(
        n20034) );
  AOI21_X1 U19527 ( .B1(n16491), .B2(n20121), .A(n16483), .ZN(n16484) );
  AOI21_X1 U19528 ( .B1(n20047), .B2(n20034), .A(n16484), .ZN(n16485) );
  AOI21_X1 U19529 ( .B1(n20034), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n16485), 
        .ZN(n16486) );
  OAI211_X1 U19530 ( .C1(n16489), .C2(n16488), .A(n16487), .B(n16486), .ZN(
        P2_U3176) );
  AOI221_X1 U19531 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n16491), .C1(
        P2_STATE2_REG_3__SCAN_IN), .C2(n20034), .A(n16490), .ZN(n16492) );
  INV_X1 U19532 ( .A(n16492), .ZN(P2_U3593) );
  INV_X1 U19533 ( .A(n16493), .ZN(n18780) );
  NOR2_X2 U19534 ( .A1(n16495), .A2(n17992), .ZN(n17895) );
  NOR2_X2 U19535 ( .A1(n18993), .A2(n16632), .ZN(n17917) );
  INV_X1 U19536 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16692) );
  NAND2_X1 U19537 ( .A1(n17919), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16925) );
  INV_X1 U19538 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17844) );
  NOR2_X1 U19539 ( .A1(n17844), .A2(n16868), .ZN(n17811) );
  NAND2_X1 U19540 ( .A1(n17811), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16668) );
  NAND3_X1 U19541 ( .A1(n17713), .A2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17686) );
  INV_X1 U19542 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17666) );
  NOR2_X1 U19543 ( .A1(n17676), .A2(n17666), .ZN(n17662) );
  NAND2_X1 U19544 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17627) );
  NAND2_X1 U19545 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16520), .ZN(
        n16506) );
  NAND2_X1 U19546 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18996), .ZN(n17989) );
  INV_X1 U19547 ( .A(n17734), .ZN(n17703) );
  NAND2_X1 U19548 ( .A1(n16526), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16496) );
  AND2_X1 U19549 ( .A1(n16496), .A2(n18719), .ZN(n16527) );
  AOI211_X1 U19550 ( .C1(n17824), .C2(n16657), .A(n17975), .B(n16527), .ZN(
        n16523) );
  OAI21_X1 U19551 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n17703), .A(
        n16523), .ZN(n16508) );
  NOR2_X1 U19552 ( .A1(n17834), .A2(n16496), .ZN(n16509) );
  INV_X1 U19553 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16682) );
  XNOR2_X1 U19554 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n16682), .ZN(
        n16497) );
  AOI22_X1 U19555 ( .A1(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n16508), .B1(
        n16509), .B2(n16497), .ZN(n16498) );
  OAI21_X1 U19556 ( .B1(n17841), .B2(n16991), .A(n16498), .ZN(n16499) );
  NAND2_X1 U19557 ( .A1(n18308), .A2(P3_REIP_REG_31__SCAN_IN), .ZN(n16500) );
  OAI21_X1 U19558 ( .B1(n16505), .B2(n17860), .A(n16504), .ZN(P3_U2799) );
  INV_X1 U19559 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18923) );
  OAI21_X1 U19560 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16520), .A(
        n16506), .ZN(n16679) );
  OAI22_X1 U19561 ( .A1(n18312), .A2(n18923), .B1(n17841), .B2(n16679), .ZN(
        n16507) );
  AOI221_X1 U19562 ( .B1(n16509), .B2(n16682), .C1(n16508), .C2(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A(n16507), .ZN(n16515) );
  OAI21_X1 U19563 ( .B1(n16510), .B2(n17634), .A(n17895), .ZN(n16517) );
  OAI21_X1 U19564 ( .B1(n16528), .B2(n17993), .A(n16517), .ZN(n16513) );
  NOR2_X2 U19565 ( .A1(n18099), .A2(n17885), .ZN(n17794) );
  NOR2_X1 U19566 ( .A1(n16511), .A2(n17774), .ZN(n17646) );
  AOI22_X1 U19567 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16513), .B1(
        n16512), .B2(n17646), .ZN(n16514) );
  OAI211_X1 U19568 ( .C1(n16516), .C2(n17898), .A(n16515), .B(n16514), .ZN(
        P3_U2800) );
  AOI21_X1 U19569 ( .B1(n16519), .B2(n16518), .A(n16517), .ZN(n16525) );
  NAND2_X1 U19570 ( .A1(n18308), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16522) );
  AOI21_X1 U19571 ( .B1(n16692), .B2(n16657), .A(n16520), .ZN(n16691) );
  OAI21_X1 U19572 ( .B1(n17734), .B2(n17827), .A(n16691), .ZN(n16521) );
  OAI211_X1 U19573 ( .C1(n16523), .C2(n16692), .A(n16522), .B(n16521), .ZN(
        n16524) );
  AOI211_X1 U19574 ( .C1(n16527), .C2(n16526), .A(n16525), .B(n16524), .ZN(
        n16532) );
  NOR2_X1 U19575 ( .A1(n16528), .A2(n17993), .ZN(n16529) );
  OAI21_X1 U19576 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16530), .A(
        n16529), .ZN(n16531) );
  OAI211_X1 U19577 ( .C1(n16533), .C2(n17898), .A(n16532), .B(n16531), .ZN(
        P3_U2801) );
  NOR3_X1 U19578 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16535) );
  NOR4_X1 U19579 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16534) );
  INV_X2 U19580 ( .A(n16617), .ZN(U215) );
  NAND4_X1 U19581 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16535), .A3(n16534), .A4(
        U215), .ZN(U213) );
  INV_X1 U19582 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19366) );
  INV_X2 U19583 ( .A(U214), .ZN(n16582) );
  INV_X1 U19584 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16620) );
  OAI222_X1 U19585 ( .A1(U212), .A2(n19366), .B1(n16584), .B2(n13065), .C1(
        U214), .C2(n16620), .ZN(U216) );
  INV_X1 U19586 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n19371) );
  INV_X1 U19587 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20434) );
  INV_X1 U19588 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n16537) );
  OAI222_X1 U19589 ( .A1(U212), .A2(n19371), .B1(n16584), .B2(n20434), .C1(
        U214), .C2(n16537), .ZN(U217) );
  INV_X1 U19590 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20427) );
  INV_X2 U19591 ( .A(U212), .ZN(n16581) );
  AOI22_X1 U19592 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16582), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16581), .ZN(n16538) );
  OAI21_X1 U19593 ( .B1(n20427), .B2(n16584), .A(n16538), .ZN(U218) );
  INV_X1 U19594 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n20420) );
  AOI22_X1 U19595 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16582), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16581), .ZN(n16539) );
  OAI21_X1 U19596 ( .B1(n20420), .B2(n16584), .A(n16539), .ZN(U219) );
  INV_X1 U19597 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n20412) );
  AOI22_X1 U19598 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16582), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16581), .ZN(n16540) );
  OAI21_X1 U19599 ( .B1(n20412), .B2(n16584), .A(n16540), .ZN(U220) );
  INV_X1 U19600 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20404) );
  AOI22_X1 U19601 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16582), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16581), .ZN(n16541) );
  OAI21_X1 U19602 ( .B1(n20404), .B2(n16584), .A(n16541), .ZN(U221) );
  INV_X1 U19603 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20395) );
  AOI22_X1 U19604 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16582), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16581), .ZN(n16542) );
  OAI21_X1 U19605 ( .B1(n20395), .B2(n16584), .A(n16542), .ZN(U222) );
  INV_X1 U19606 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n20378) );
  AOI22_X1 U19607 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16582), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16581), .ZN(n16543) );
  OAI21_X1 U19608 ( .B1(n20378), .B2(n16584), .A(n16543), .ZN(U223) );
  INV_X1 U19609 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n20439) );
  AOI22_X1 U19610 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16582), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16581), .ZN(n16544) );
  OAI21_X1 U19611 ( .B1(n20439), .B2(n16584), .A(n16544), .ZN(U224) );
  INV_X1 U19612 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n20432) );
  AOI22_X1 U19613 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16582), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16581), .ZN(n16545) );
  OAI21_X1 U19614 ( .B1(n20432), .B2(n16584), .A(n16545), .ZN(U225) );
  INV_X1 U19615 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20425) );
  AOI22_X1 U19616 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16582), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16581), .ZN(n16546) );
  OAI21_X1 U19617 ( .B1(n20425), .B2(n16584), .A(n16546), .ZN(U226) );
  INV_X1 U19618 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n20418) );
  AOI22_X1 U19619 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16582), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16581), .ZN(n16547) );
  OAI21_X1 U19620 ( .B1(n20418), .B2(n16584), .A(n16547), .ZN(U227) );
  INV_X1 U19621 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n20410) );
  AOI22_X1 U19622 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16582), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16581), .ZN(n16548) );
  OAI21_X1 U19623 ( .B1(n20410), .B2(n16584), .A(n16548), .ZN(U228) );
  INV_X1 U19624 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n20401) );
  AOI22_X1 U19625 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16582), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16581), .ZN(n16549) );
  OAI21_X1 U19626 ( .B1(n20401), .B2(n16584), .A(n16549), .ZN(U229) );
  INV_X1 U19627 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20394) );
  AOI22_X1 U19628 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16582), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16581), .ZN(n16550) );
  OAI21_X1 U19629 ( .B1(n20394), .B2(n16584), .A(n16550), .ZN(U230) );
  INV_X1 U19630 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n20375) );
  AOI22_X1 U19631 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16582), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16581), .ZN(n16551) );
  OAI21_X1 U19632 ( .B1(n20375), .B2(n16584), .A(n16551), .ZN(U231) );
  AOI22_X1 U19633 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16582), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16581), .ZN(n16552) );
  OAI21_X1 U19634 ( .B1(n13743), .B2(n16584), .A(n16552), .ZN(U232) );
  AOI22_X1 U19635 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16582), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16581), .ZN(n16553) );
  OAI21_X1 U19636 ( .B1(n16554), .B2(n16584), .A(n16553), .ZN(U233) );
  AOI22_X1 U19637 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16582), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16581), .ZN(n16555) );
  OAI21_X1 U19638 ( .B1(n16556), .B2(n16584), .A(n16555), .ZN(U234) );
  AOI22_X1 U19639 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16582), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16581), .ZN(n16557) );
  OAI21_X1 U19640 ( .B1(n16558), .B2(n16584), .A(n16557), .ZN(U235) );
  AOI22_X1 U19641 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16582), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16581), .ZN(n16559) );
  OAI21_X1 U19642 ( .B1(n16560), .B2(n16584), .A(n16559), .ZN(U236) );
  AOI22_X1 U19643 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16582), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16581), .ZN(n16561) );
  OAI21_X1 U19644 ( .B1(n16562), .B2(n16584), .A(n16561), .ZN(U237) );
  AOI22_X1 U19645 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16582), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16581), .ZN(n16563) );
  OAI21_X1 U19646 ( .B1(n16564), .B2(n16584), .A(n16563), .ZN(U238) );
  INV_X1 U19647 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16566) );
  AOI22_X1 U19648 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16582), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16581), .ZN(n16565) );
  OAI21_X1 U19649 ( .B1(n16566), .B2(n16584), .A(n16565), .ZN(U239) );
  INV_X1 U19650 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16568) );
  AOI22_X1 U19651 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16582), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16581), .ZN(n16567) );
  OAI21_X1 U19652 ( .B1(n16568), .B2(n16584), .A(n16567), .ZN(U240) );
  AOI22_X1 U19653 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16582), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16581), .ZN(n16569) );
  OAI21_X1 U19654 ( .B1(n16570), .B2(n16584), .A(n16569), .ZN(U241) );
  AOI22_X1 U19655 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16582), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16581), .ZN(n16571) );
  OAI21_X1 U19656 ( .B1(n16572), .B2(n16584), .A(n16571), .ZN(U242) );
  AOI22_X1 U19657 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16582), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16581), .ZN(n16573) );
  OAI21_X1 U19658 ( .B1(n16574), .B2(n16584), .A(n16573), .ZN(U243) );
  AOI22_X1 U19659 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16582), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16581), .ZN(n16575) );
  OAI21_X1 U19660 ( .B1(n16576), .B2(n16584), .A(n16575), .ZN(U244) );
  AOI22_X1 U19661 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16582), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16581), .ZN(n16577) );
  OAI21_X1 U19662 ( .B1(n16578), .B2(n16584), .A(n16577), .ZN(U245) );
  AOI22_X1 U19663 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16582), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16581), .ZN(n16579) );
  OAI21_X1 U19664 ( .B1(n16580), .B2(n16584), .A(n16579), .ZN(U246) );
  AOI22_X1 U19665 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16582), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16581), .ZN(n16583) );
  OAI21_X1 U19666 ( .B1(n16585), .B2(n16584), .A(n16583), .ZN(U247) );
  INV_X1 U19667 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n16586) );
  AOI22_X1 U19668 ( .A1(n16617), .A2(n16586), .B1(n18329), .B2(U215), .ZN(U251) );
  OAI22_X1 U19669 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16617), .ZN(n16587) );
  INV_X1 U19670 ( .A(n16587), .ZN(U252) );
  INV_X1 U19671 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16588) );
  AOI22_X1 U19672 ( .A1(n16617), .A2(n16588), .B1(n18342), .B2(U215), .ZN(U253) );
  INV_X1 U19673 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16589) );
  INV_X1 U19674 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18346) );
  AOI22_X1 U19675 ( .A1(n16617), .A2(n16589), .B1(n18346), .B2(U215), .ZN(U254) );
  INV_X1 U19676 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16590) );
  INV_X1 U19677 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18350) );
  AOI22_X1 U19678 ( .A1(n16617), .A2(n16590), .B1(n18350), .B2(U215), .ZN(U255) );
  INV_X1 U19679 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16591) );
  INV_X1 U19680 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18354) );
  AOI22_X1 U19681 ( .A1(n16618), .A2(n16591), .B1(n18354), .B2(U215), .ZN(U256) );
  INV_X1 U19682 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16592) );
  INV_X1 U19683 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18358) );
  AOI22_X1 U19684 ( .A1(n16618), .A2(n16592), .B1(n18358), .B2(U215), .ZN(U257) );
  INV_X1 U19685 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16593) );
  INV_X1 U19686 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18363) );
  AOI22_X1 U19687 ( .A1(n16617), .A2(n16593), .B1(n18363), .B2(U215), .ZN(U258) );
  INV_X1 U19688 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16594) );
  INV_X1 U19689 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17483) );
  AOI22_X1 U19690 ( .A1(n16618), .A2(n16594), .B1(n17483), .B2(U215), .ZN(U259) );
  INV_X1 U19691 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16595) );
  INV_X1 U19692 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17478) );
  AOI22_X1 U19693 ( .A1(n16617), .A2(n16595), .B1(n17478), .B2(U215), .ZN(U260) );
  OAI22_X1 U19694 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16617), .ZN(n16596) );
  INV_X1 U19695 ( .A(n16596), .ZN(U261) );
  OAI22_X1 U19696 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16617), .ZN(n16597) );
  INV_X1 U19697 ( .A(n16597), .ZN(U262) );
  INV_X1 U19698 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16598) );
  INV_X1 U19699 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17467) );
  AOI22_X1 U19700 ( .A1(n16617), .A2(n16598), .B1(n17467), .B2(U215), .ZN(U263) );
  INV_X1 U19701 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16599) );
  INV_X1 U19702 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17462) );
  AOI22_X1 U19703 ( .A1(n16617), .A2(n16599), .B1(n17462), .B2(U215), .ZN(U264) );
  OAI22_X1 U19704 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16617), .ZN(n16600) );
  INV_X1 U19705 ( .A(n16600), .ZN(U265) );
  OAI22_X1 U19706 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16617), .ZN(n16601) );
  INV_X1 U19707 ( .A(n16601), .ZN(U266) );
  INV_X1 U19708 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n16602) );
  INV_X1 U19709 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n19443) );
  AOI22_X1 U19710 ( .A1(n16618), .A2(n16602), .B1(n19443), .B2(U215), .ZN(U267) );
  INV_X1 U19711 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n16603) );
  INV_X1 U19712 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n19449) );
  AOI22_X1 U19713 ( .A1(n16617), .A2(n16603), .B1(n19449), .B2(U215), .ZN(U268) );
  INV_X1 U19714 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n16604) );
  INV_X1 U19715 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n19454) );
  AOI22_X1 U19716 ( .A1(n16617), .A2(n16604), .B1(n19454), .B2(U215), .ZN(U269) );
  OAI22_X1 U19717 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16618), .ZN(n16605) );
  INV_X1 U19718 ( .A(n16605), .ZN(U270) );
  OAI22_X1 U19719 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16618), .ZN(n16606) );
  INV_X1 U19720 ( .A(n16606), .ZN(U271) );
  INV_X1 U19721 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n16607) );
  AOI22_X1 U19722 ( .A1(n16617), .A2(n16607), .B1(n15083), .B2(U215), .ZN(U272) );
  INV_X1 U19723 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n16608) );
  INV_X1 U19724 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n18359) );
  AOI22_X1 U19725 ( .A1(n16617), .A2(n16608), .B1(n18359), .B2(U215), .ZN(U273) );
  OAI22_X1 U19726 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16617), .ZN(n16609) );
  INV_X1 U19727 ( .A(n16609), .ZN(U274) );
  OAI22_X1 U19728 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16618), .ZN(n16610) );
  INV_X1 U19729 ( .A(n16610), .ZN(U275) );
  OAI22_X1 U19730 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16617), .ZN(n16611) );
  INV_X1 U19731 ( .A(n16611), .ZN(U276) );
  OAI22_X1 U19732 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16617), .ZN(n16612) );
  INV_X1 U19733 ( .A(n16612), .ZN(U277) );
  OAI22_X1 U19734 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16617), .ZN(n16614) );
  INV_X1 U19735 ( .A(n16614), .ZN(U278) );
  INV_X1 U19736 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n16615) );
  INV_X1 U19737 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n19463) );
  AOI22_X1 U19738 ( .A1(n16618), .A2(n16615), .B1(n19463), .B2(U215), .ZN(U279) );
  INV_X1 U19739 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n16616) );
  INV_X1 U19740 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n19469) );
  AOI22_X1 U19741 ( .A1(n16617), .A2(n16616), .B1(n19469), .B2(U215), .ZN(U280) );
  INV_X1 U19742 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n19474) );
  AOI22_X1 U19743 ( .A1(n16618), .A2(n19371), .B1(n19474), .B2(U215), .ZN(U281) );
  INV_X1 U19744 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19483) );
  AOI22_X1 U19745 ( .A1(n16618), .A2(n19366), .B1(n19483), .B2(U215), .ZN(U282) );
  INV_X1 U19746 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16619) );
  AOI222_X1 U19747 ( .A1(n16620), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n19366), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16619), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16621) );
  INV_X2 U19748 ( .A(n16623), .ZN(n16622) );
  INV_X1 U19749 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18883) );
  INV_X1 U19750 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20070) );
  AOI22_X1 U19751 ( .A1(n16622), .A2(n18883), .B1(n20070), .B2(n16623), .ZN(
        U347) );
  INV_X1 U19752 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18881) );
  INV_X1 U19753 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20068) );
  AOI22_X1 U19754 ( .A1(n16622), .A2(n18881), .B1(n20068), .B2(n16623), .ZN(
        U348) );
  INV_X1 U19755 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18878) );
  INV_X1 U19756 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20067) );
  AOI22_X1 U19757 ( .A1(n16622), .A2(n18878), .B1(n20067), .B2(n16623), .ZN(
        U349) );
  INV_X1 U19758 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18877) );
  INV_X1 U19759 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20066) );
  AOI22_X1 U19760 ( .A1(n16622), .A2(n18877), .B1(n20066), .B2(n16623), .ZN(
        U350) );
  INV_X1 U19761 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18875) );
  INV_X1 U19762 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20064) );
  AOI22_X1 U19763 ( .A1(n16622), .A2(n18875), .B1(n20064), .B2(n16623), .ZN(
        U351) );
  INV_X1 U19764 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18873) );
  INV_X1 U19765 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20062) );
  AOI22_X1 U19766 ( .A1(n16622), .A2(n18873), .B1(n20062), .B2(n16623), .ZN(
        U352) );
  INV_X1 U19767 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18871) );
  INV_X1 U19768 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20061) );
  AOI22_X1 U19769 ( .A1(n16622), .A2(n18871), .B1(n20061), .B2(n16623), .ZN(
        U353) );
  INV_X1 U19770 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18869) );
  AOI22_X1 U19771 ( .A1(n16622), .A2(n18869), .B1(n20059), .B2(n16623), .ZN(
        U354) );
  INV_X1 U19772 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18921) );
  INV_X1 U19773 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20105) );
  AOI22_X1 U19774 ( .A1(n16622), .A2(n18921), .B1(n20105), .B2(n16623), .ZN(
        U356) );
  INV_X1 U19775 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18918) );
  INV_X1 U19776 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20103) );
  AOI22_X1 U19777 ( .A1(n16622), .A2(n18918), .B1(n20103), .B2(n16623), .ZN(
        U357) );
  INV_X1 U19778 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18917) );
  INV_X1 U19779 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20100) );
  AOI22_X1 U19780 ( .A1(n16622), .A2(n18917), .B1(n20100), .B2(n16623), .ZN(
        U358) );
  INV_X1 U19781 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18915) );
  INV_X1 U19782 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20099) );
  AOI22_X1 U19783 ( .A1(n16622), .A2(n18915), .B1(n20099), .B2(n16623), .ZN(
        U359) );
  INV_X1 U19784 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18913) );
  INV_X1 U19785 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20097) );
  AOI22_X1 U19786 ( .A1(n16622), .A2(n18913), .B1(n20097), .B2(n16623), .ZN(
        U360) );
  INV_X1 U19787 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18911) );
  INV_X1 U19788 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20095) );
  AOI22_X1 U19789 ( .A1(n16622), .A2(n18911), .B1(n20095), .B2(n16623), .ZN(
        U361) );
  INV_X1 U19790 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18908) );
  INV_X1 U19791 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20093) );
  AOI22_X1 U19792 ( .A1(n16622), .A2(n18908), .B1(n20093), .B2(n16623), .ZN(
        U362) );
  INV_X1 U19793 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18907) );
  INV_X1 U19794 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20091) );
  AOI22_X1 U19795 ( .A1(n16622), .A2(n18907), .B1(n20091), .B2(n16623), .ZN(
        U363) );
  INV_X1 U19796 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18904) );
  INV_X1 U19797 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20089) );
  AOI22_X1 U19798 ( .A1(n16622), .A2(n18904), .B1(n20089), .B2(n16623), .ZN(
        U364) );
  INV_X1 U19799 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18867) );
  INV_X1 U19800 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20058) );
  AOI22_X1 U19801 ( .A1(n16622), .A2(n18867), .B1(n20058), .B2(n16623), .ZN(
        U365) );
  INV_X1 U19802 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18903) );
  INV_X1 U19803 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20087) );
  AOI22_X1 U19804 ( .A1(n16622), .A2(n18903), .B1(n20087), .B2(n16623), .ZN(
        U366) );
  INV_X1 U19805 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18900) );
  INV_X1 U19806 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20086) );
  AOI22_X1 U19807 ( .A1(n16622), .A2(n18900), .B1(n20086), .B2(n16623), .ZN(
        U367) );
  INV_X1 U19808 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18899) );
  INV_X1 U19809 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20084) );
  AOI22_X1 U19810 ( .A1(n16622), .A2(n18899), .B1(n20084), .B2(n16623), .ZN(
        U368) );
  INV_X1 U19811 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18897) );
  INV_X1 U19812 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20082) );
  AOI22_X1 U19813 ( .A1(n16622), .A2(n18897), .B1(n20082), .B2(n16623), .ZN(
        U369) );
  INV_X1 U19814 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18895) );
  INV_X1 U19815 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20080) );
  AOI22_X1 U19816 ( .A1(n16622), .A2(n18895), .B1(n20080), .B2(n16623), .ZN(
        U370) );
  INV_X1 U19817 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18893) );
  INV_X1 U19818 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20079) );
  AOI22_X1 U19819 ( .A1(n16622), .A2(n18893), .B1(n20079), .B2(n16623), .ZN(
        U371) );
  INV_X1 U19820 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18890) );
  INV_X1 U19821 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20077) );
  AOI22_X1 U19822 ( .A1(n16622), .A2(n18890), .B1(n20077), .B2(n16623), .ZN(
        U372) );
  INV_X1 U19823 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18889) );
  INV_X1 U19824 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20075) );
  AOI22_X1 U19825 ( .A1(n16622), .A2(n18889), .B1(n20075), .B2(n16623), .ZN(
        U373) );
  INV_X1 U19826 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18887) );
  INV_X1 U19827 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20074) );
  AOI22_X1 U19828 ( .A1(n16622), .A2(n18887), .B1(n20074), .B2(n16623), .ZN(
        U374) );
  INV_X1 U19829 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18885) );
  INV_X1 U19830 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20072) );
  AOI22_X1 U19831 ( .A1(n16622), .A2(n18885), .B1(n20072), .B2(n16623), .ZN(
        U375) );
  INV_X1 U19832 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18865) );
  INV_X1 U19833 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20057) );
  AOI22_X1 U19834 ( .A1(n16622), .A2(n18865), .B1(n20057), .B2(n16623), .ZN(
        U376) );
  INV_X1 U19835 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16624) );
  INV_X1 U19836 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18864) );
  NAND2_X1 U19837 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18864), .ZN(n18856) );
  AOI22_X1 U19838 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18856), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n18862), .ZN(n18939) );
  OAI21_X1 U19839 ( .B1(n18862), .B2(n16624), .A(n18936), .ZN(P3_U2633) );
  INV_X1 U19840 ( .A(P3_CODEFETCH_REG_SCAN_IN), .ZN(n16627) );
  NAND2_X1 U19841 ( .A1(n18839), .A2(n16625), .ZN(n16626) );
  OAI221_X1 U19842 ( .B1(n16627), .B2(n17553), .C1(n16627), .C2(n16629), .A(
        n16626), .ZN(P3_U2634) );
  AOI21_X1 U19843 ( .B1(n18862), .B2(n18864), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16628) );
  AOI22_X1 U19844 ( .A1(n18933), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16628), 
        .B2(n19003), .ZN(P3_U2635) );
  OAI21_X1 U19845 ( .B1(n18849), .B2(BS16), .A(n18939), .ZN(n18937) );
  OAI21_X1 U19846 ( .B1(n18939), .B2(n16655), .A(n18937), .ZN(P3_U2636) );
  AND3_X1 U19847 ( .A1(n16631), .A2(n16630), .A3(n16629), .ZN(n18824) );
  NOR2_X1 U19848 ( .A1(n18824), .A2(n18828), .ZN(n18984) );
  OAI21_X1 U19849 ( .B1(n18984), .B2(n18322), .A(n16632), .ZN(P3_U2637) );
  NOR4_X1 U19850 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16636) );
  NOR4_X1 U19851 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16635) );
  NOR4_X1 U19852 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16634) );
  NOR4_X1 U19853 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16633) );
  NAND4_X1 U19854 ( .A1(n16636), .A2(n16635), .A3(n16634), .A4(n16633), .ZN(
        n16642) );
  NOR4_X1 U19855 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16640) );
  AOI211_X1 U19856 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16639) );
  NOR4_X1 U19857 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16638) );
  NOR4_X1 U19858 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16637) );
  NAND4_X1 U19859 ( .A1(n16640), .A2(n16639), .A3(n16638), .A4(n16637), .ZN(
        n16641) );
  NOR2_X1 U19860 ( .A1(n16642), .A2(n16641), .ZN(n18978) );
  INV_X1 U19861 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18931) );
  NOR3_X1 U19862 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16644) );
  OAI21_X1 U19863 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16644), .A(n18978), .ZN(
        n16643) );
  OAI21_X1 U19864 ( .B1(n18978), .B2(n18931), .A(n16643), .ZN(P3_U2638) );
  INV_X1 U19865 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18974) );
  INV_X1 U19866 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18938) );
  AOI21_X1 U19867 ( .B1(n18974), .B2(n18938), .A(n16644), .ZN(n16645) );
  INV_X1 U19868 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18928) );
  INV_X1 U19869 ( .A(n18978), .ZN(n18981) );
  AOI22_X1 U19870 ( .A1(n18978), .A2(n16645), .B1(n18928), .B2(n18981), .ZN(
        P3_U2639) );
  NOR2_X1 U19871 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18942), .ZN(n18713) );
  INV_X1 U19872 ( .A(n18842), .ZN(n17012) );
  AOI211_X1 U19873 ( .C1(n18839), .C2(n18713), .A(n9822), .B(n17012), .ZN(
        n16649) );
  NAND3_X1 U19874 ( .A1(n16648), .A2(n16647), .A3(n16646), .ZN(n18778) );
  NAND2_X1 U19875 ( .A1(n17553), .A2(n18778), .ZN(n16650) );
  OAI211_X1 U19876 ( .C1(n18992), .C2(n18993), .A(n18988), .B(n16655), .ZN(
        n18774) );
  INV_X1 U19877 ( .A(n18774), .ZN(n16651) );
  AOI211_X4 U19878 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18993), .A(n16651), .B(
        n16654), .ZN(n17007) );
  AOI22_X1 U19879 ( .A1(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n17018), .B1(
        P3_EBX_REG_31__SCAN_IN), .B2(n17007), .ZN(n16678) );
  INV_X1 U19880 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18925) );
  AOI22_X1 U19881 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(P3_REIP_REG_30__SCAN_IN), 
        .B1(n18923), .B2(n18925), .ZN(n16656) );
  INV_X1 U19882 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18920) );
  INV_X1 U19883 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18898) );
  INV_X1 U19884 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18891) );
  INV_X1 U19885 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18886) );
  INV_X1 U19886 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18879) );
  INV_X1 U19887 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18874) );
  INV_X1 U19888 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18870) );
  NAND3_X1 U19889 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16989) );
  NOR2_X1 U19890 ( .A1(n18870), .A2(n16989), .ZN(n16964) );
  NAND2_X1 U19891 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16964), .ZN(n16958) );
  NOR2_X1 U19892 ( .A1(n18874), .A2(n16958), .ZN(n16934) );
  NAND2_X1 U19893 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n16934), .ZN(n16924) );
  NOR2_X1 U19894 ( .A1(n18879), .A2(n16924), .ZN(n16862) );
  NAND4_X1 U19895 ( .A1(n16862), .A2(P3_REIP_REG_11__SCAN_IN), .A3(
        P3_REIP_REG_10__SCAN_IN), .A4(P3_REIP_REG_9__SCAN_IN), .ZN(n16877) );
  NOR2_X1 U19896 ( .A1(n18886), .A2(n16877), .ZN(n16872) );
  NAND2_X1 U19897 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16872), .ZN(n16670) );
  NAND4_X1 U19898 ( .A1(n16845), .A2(P3_REIP_REG_17__SCAN_IN), .A3(
        P3_REIP_REG_16__SCAN_IN), .A4(P3_REIP_REG_15__SCAN_IN), .ZN(n16816) );
  NAND3_X1 U19899 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n16800), .A3(
        P3_REIP_REG_20__SCAN_IN), .ZN(n16769) );
  INV_X1 U19900 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18905) );
  INV_X1 U19901 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18906) );
  NOR2_X1 U19902 ( .A1(n18905), .A2(n18906), .ZN(n16770) );
  NAND2_X1 U19903 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16770), .ZN(n16669) );
  NAND2_X1 U19904 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16750), .ZN(n16743) );
  NAND2_X1 U19905 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .ZN(n16652) );
  NAND3_X1 U19906 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16712), .ZN(n16698) );
  NOR2_X1 U19907 ( .A1(n18920), .A2(n16698), .ZN(n16684) );
  NAND2_X1 U19908 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18993), .ZN(n16653) );
  AOI211_X4 U19909 ( .C1(n18988), .C2(n16655), .A(n16654), .B(n16653), .ZN(
        n17026) );
  NOR3_X1 U19910 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17003) );
  INV_X1 U19911 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17341) );
  NAND2_X1 U19912 ( .A1(n17003), .A2(n17341), .ZN(n16998) );
  NOR2_X1 U19913 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16998), .ZN(n16974) );
  INV_X1 U19914 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16966) );
  NAND2_X1 U19915 ( .A1(n16974), .A2(n16966), .ZN(n16965) );
  NAND2_X1 U19916 ( .A1(n16946), .A2(n17331), .ZN(n16943) );
  NAND2_X1 U19917 ( .A1(n16915), .A2(n16920), .ZN(n16906) );
  NAND2_X1 U19918 ( .A1(n16905), .A2(n17250), .ZN(n16893) );
  NAND2_X1 U19919 ( .A1(n16876), .A2(n16875), .ZN(n16865) );
  INV_X1 U19920 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16849) );
  NAND2_X1 U19921 ( .A1(n16853), .A2(n16849), .ZN(n16846) );
  INV_X1 U19922 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16819) );
  NAND2_X1 U19923 ( .A1(n16829), .A2(n16819), .ZN(n16818) );
  NAND2_X1 U19924 ( .A1(n16811), .A2(n16802), .ZN(n16801) );
  INV_X1 U19925 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17134) );
  NAND2_X1 U19926 ( .A1(n16786), .A2(n17134), .ZN(n16780) );
  INV_X1 U19927 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n17039) );
  NAND2_X1 U19928 ( .A1(n16763), .A2(n17039), .ZN(n16759) );
  INV_X1 U19929 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17042) );
  NAND2_X1 U19930 ( .A1(n16744), .A2(n17042), .ZN(n16740) );
  NAND2_X1 U19931 ( .A1(n16726), .A2(n16718), .ZN(n16717) );
  NOR2_X1 U19932 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16717), .ZN(n16711) );
  INV_X1 U19933 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17082) );
  NAND2_X1 U19934 ( .A1(n16711), .A2(n17082), .ZN(n16681) );
  NOR2_X1 U19935 ( .A1(n17030), .A2(n16681), .ZN(n16685) );
  INV_X1 U19936 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17049) );
  AOI22_X1 U19937 ( .A1(n16656), .A2(n16684), .B1(n16685), .B2(n17049), .ZN(
        n16677) );
  INV_X1 U19938 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17643) );
  NAND2_X1 U19939 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17714) );
  NAND2_X1 U19940 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17713), .ZN(
        n16665) );
  NAND2_X1 U19941 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17664), .ZN(
        n16663) );
  INV_X1 U19942 ( .A(n16663), .ZN(n16659) );
  NAND3_X1 U19943 ( .A1(n17662), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A3(
        n16659), .ZN(n16660) );
  NOR2_X1 U19944 ( .A1(n17643), .A2(n16660), .ZN(n16658) );
  OAI21_X1 U19945 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16658), .A(
        n16657), .ZN(n17630) );
  INV_X1 U19946 ( .A(n17630), .ZN(n16702) );
  AOI21_X1 U19947 ( .B1(n17643), .B2(n16660), .A(n16658), .ZN(n17638) );
  NAND2_X1 U19948 ( .A1(n17662), .A2(n16659), .ZN(n16661) );
  INV_X1 U19949 ( .A(n16661), .ZN(n17621) );
  OAI21_X1 U19950 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17621), .A(
        n16660), .ZN(n17654) );
  INV_X1 U19951 ( .A(n17654), .ZN(n16725) );
  NOR2_X1 U19952 ( .A1(n17676), .A2(n16663), .ZN(n16662) );
  OAI21_X1 U19953 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16662), .A(
        n16661), .ZN(n17665) );
  INV_X1 U19954 ( .A(n17665), .ZN(n16735) );
  AOI21_X1 U19955 ( .B1(n17676), .B2(n16663), .A(n16662), .ZN(n17679) );
  OAI21_X1 U19956 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17664), .A(
        n16663), .ZN(n17700) );
  INV_X1 U19957 ( .A(n17700), .ZN(n16755) );
  INV_X1 U19958 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16775) );
  INV_X1 U19959 ( .A(n16665), .ZN(n16666) );
  NAND2_X1 U19960 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16666), .ZN(
        n16664) );
  AOI21_X1 U19961 ( .B1(n16775), .B2(n16664), .A(n17664), .ZN(n17704) );
  INV_X1 U19962 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17720) );
  OAI22_X1 U19963 ( .A1(n17720), .A2(n16666), .B1(n16665), .B2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17718) );
  INV_X1 U19964 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17983) );
  NOR2_X1 U19965 ( .A1(n17983), .A2(n17737), .ZN(n17701) );
  INV_X1 U19966 ( .A(n17701), .ZN(n16795) );
  AOI21_X1 U19967 ( .B1(n17736), .B2(n16795), .A(n16666), .ZN(n17740) );
  AND2_X1 U19968 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17889), .ZN(
        n16935) );
  NAND2_X1 U19969 ( .A1(n16667), .A2(n16935), .ZN(n17823) );
  NOR2_X1 U19970 ( .A1(n16668), .A2(n17823), .ZN(n17787) );
  NAND2_X1 U19971 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17787), .ZN(
        n16839) );
  NOR2_X1 U19972 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16839), .ZN(
        n16807) );
  AOI21_X1 U19973 ( .B1(n17701), .B2(n16807), .A(n9847), .ZN(n16785) );
  NOR2_X1 U19974 ( .A1(n17740), .A2(n16785), .ZN(n16784) );
  NOR2_X1 U19975 ( .A1(n16767), .A2(n16991), .ZN(n16754) );
  NOR2_X1 U19976 ( .A1(n16755), .A2(n16754), .ZN(n16753) );
  NOR2_X1 U19977 ( .A1(n16753), .A2(n16991), .ZN(n16748) );
  NOR2_X1 U19978 ( .A1(n17679), .A2(n16748), .ZN(n16747) );
  NOR2_X1 U19979 ( .A1(n17638), .A2(n16714), .ZN(n16713) );
  NOR2_X1 U19980 ( .A1(n16713), .A2(n16991), .ZN(n16701) );
  NOR2_X1 U19981 ( .A1(n16702), .A2(n16701), .ZN(n16700) );
  NAND4_X1 U19982 ( .A1(n16959), .A2(n17012), .A3(n16689), .A4(n16679), .ZN(
        n16676) );
  NAND2_X1 U19983 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16707) );
  INV_X1 U19984 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18910) );
  INV_X1 U19985 ( .A(n16669), .ZN(n16673) );
  NAND2_X1 U19986 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_20__SCAN_IN), 
        .ZN(n16672) );
  INV_X1 U19987 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18896) );
  NAND2_X1 U19988 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16836) );
  NOR2_X1 U19989 ( .A1(n18896), .A2(n16836), .ZN(n16671) );
  NOR2_X1 U19990 ( .A1(n18891), .A2(n16670), .ZN(n16827) );
  NAND3_X1 U19991 ( .A1(n16671), .A2(n16827), .A3(n17034), .ZN(n16793) );
  NOR3_X1 U19992 ( .A1(n18898), .A2(n16672), .A3(n16793), .ZN(n16765) );
  NAND2_X1 U19993 ( .A1(n16673), .A2(n16765), .ZN(n16746) );
  NOR2_X1 U19994 ( .A1(n18910), .A2(n16746), .ZN(n16737) );
  NAND3_X1 U19995 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .A3(n16737), .ZN(n16703) );
  NOR2_X1 U19996 ( .A1(n16707), .A2(n16703), .ZN(n16674) );
  NOR2_X1 U19997 ( .A1(n17009), .A2(n16973), .ZN(n16766) );
  AOI21_X1 U19998 ( .B1(P3_REIP_REG_29__SCAN_IN), .B2(n16674), .A(n16766), 
        .ZN(n16694) );
  NAND2_X1 U19999 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n16694), .ZN(n16675) );
  NAND4_X1 U20000 ( .A1(n16678), .A2(n16677), .A3(n16676), .A4(n16675), .ZN(
        P3_U2640) );
  NOR2_X1 U20001 ( .A1(n16689), .A2(n16991), .ZN(n16680) );
  XOR2_X1 U20002 ( .A(n16680), .B(n16679), .Z(n16688) );
  NAND2_X1 U20003 ( .A1(n17026), .A2(n16681), .ZN(n16695) );
  OAI22_X1 U20004 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16695), .B1(n16682), 
        .B2(n16969), .ZN(n16683) );
  AOI221_X1 U20005 ( .B1(n16694), .B2(P3_REIP_REG_30__SCAN_IN), .C1(n16684), 
        .C2(n18923), .A(n16683), .ZN(n16687) );
  OAI21_X1 U20006 ( .B1(n17007), .B2(n16685), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16686) );
  OAI211_X1 U20007 ( .C1(n18842), .C2(n16688), .A(n16687), .B(n16686), .ZN(
        P3_U2641) );
  OAI22_X1 U20008 ( .A1(n16692), .A2(n16969), .B1(n17031), .B2(n17082), .ZN(
        n16693) );
  INV_X1 U20009 ( .A(n16695), .ZN(n16696) );
  OAI21_X1 U20010 ( .B1(n16711), .B2(n17082), .A(n16696), .ZN(n16697) );
  INV_X1 U20011 ( .A(n16717), .ZN(n16699) );
  OAI21_X1 U20012 ( .B1(n16699), .B2(n16704), .A(n17026), .ZN(n16710) );
  AOI211_X1 U20013 ( .C1(n16702), .C2(n16701), .A(n16700), .B(n18842), .ZN(
        n16706) );
  INV_X1 U20014 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18919) );
  NAND2_X1 U20015 ( .A1(n17032), .A2(n16703), .ZN(n16731) );
  OAI22_X1 U20016 ( .A1(n18919), .A2(n16731), .B1(n17031), .B2(n16704), .ZN(
        n16705) );
  AOI211_X1 U20017 ( .C1(n17018), .C2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16706), .B(n16705), .ZN(n16709) );
  OAI211_X1 U20018 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16712), .B(n16707), .ZN(n16708) );
  OAI211_X1 U20019 ( .C1(n16711), .C2(n16710), .A(n16709), .B(n16708), .ZN(
        P3_U2643) );
  INV_X1 U20020 ( .A(n16712), .ZN(n16721) );
  AOI211_X1 U20021 ( .C1(n17638), .C2(n16714), .A(n16713), .B(n18842), .ZN(
        n16716) );
  INV_X1 U20022 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18916) );
  OAI22_X1 U20023 ( .A1(n18916), .A2(n16731), .B1(n17031), .B2(n16718), .ZN(
        n16715) );
  AOI211_X1 U20024 ( .C1(n17018), .C2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16716), .B(n16715), .ZN(n16720) );
  OAI211_X1 U20025 ( .C1(n16726), .C2(n16718), .A(n17026), .B(n16717), .ZN(
        n16719) );
  OAI211_X1 U20026 ( .C1(P3_REIP_REG_27__SCAN_IN), .C2(n16721), .A(n16720), 
        .B(n16719), .ZN(P3_U2644) );
  INV_X1 U20027 ( .A(n16743), .ZN(n16722) );
  AOI21_X1 U20028 ( .B1(P3_REIP_REG_25__SCAN_IN), .B2(n16722), .A(
        P3_REIP_REG_26__SCAN_IN), .ZN(n16732) );
  AOI211_X1 U20029 ( .C1(n16725), .C2(n16724), .A(n16723), .B(n18842), .ZN(
        n16729) );
  AOI211_X1 U20030 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16740), .A(n16726), .B(
        n17030), .ZN(n16728) );
  INV_X1 U20031 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n17043) );
  OAI22_X1 U20032 ( .A1(n10073), .A2(n16969), .B1(n17031), .B2(n17043), .ZN(
        n16727) );
  NOR3_X1 U20033 ( .A1(n16729), .A2(n16728), .A3(n16727), .ZN(n16730) );
  OAI21_X1 U20034 ( .B1(n16732), .B2(n16731), .A(n16730), .ZN(P3_U2645) );
  AOI211_X1 U20035 ( .C1(n16735), .C2(n16734), .A(n16733), .B(n18842), .ZN(
        n16739) );
  NAND2_X1 U20036 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n17032), .ZN(n16736) );
  OAI22_X1 U20037 ( .A1(n16737), .A2(n16736), .B1(n17031), .B2(n17042), .ZN(
        n16738) );
  AOI211_X1 U20038 ( .C1(n17018), .C2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16739), .B(n16738), .ZN(n16742) );
  OAI211_X1 U20039 ( .C1(n16744), .C2(n17042), .A(n17026), .B(n16740), .ZN(
        n16741) );
  OAI211_X1 U20040 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n16743), .A(n16742), 
        .B(n16741), .ZN(P3_U2646) );
  AOI211_X1 U20041 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16759), .A(n16744), .B(
        n17030), .ZN(n16745) );
  AOI21_X1 U20042 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17007), .A(n16745), .ZN(
        n16752) );
  AND2_X1 U20043 ( .A1(n17032), .A2(n16746), .ZN(n16758) );
  AOI211_X1 U20044 ( .C1(n17679), .C2(n16748), .A(n16747), .B(n18842), .ZN(
        n16749) );
  AOI221_X1 U20045 ( .B1(n16758), .B2(P3_REIP_REG_24__SCAN_IN), .C1(n16750), 
        .C2(n18910), .A(n16749), .ZN(n16751) );
  OAI211_X1 U20046 ( .C1(n17676), .C2(n16969), .A(n16752), .B(n16751), .ZN(
        P3_U2647) );
  AOI22_X1 U20047 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17018), .B1(
        n17007), .B2(P3_EBX_REG_23__SCAN_IN), .ZN(n16762) );
  INV_X1 U20048 ( .A(n16769), .ZN(n16779) );
  AND2_X1 U20049 ( .A1(n16779), .A2(n16770), .ZN(n16757) );
  INV_X1 U20050 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18909) );
  AOI211_X1 U20051 ( .C1(n16755), .C2(n16754), .A(n16753), .B(n18842), .ZN(
        n16756) );
  AOI221_X1 U20052 ( .B1(n16758), .B2(P3_REIP_REG_23__SCAN_IN), .C1(n16757), 
        .C2(n18909), .A(n16756), .ZN(n16761) );
  OAI211_X1 U20053 ( .C1(n16763), .C2(n17039), .A(n17026), .B(n16759), .ZN(
        n16760) );
  NAND3_X1 U20054 ( .A1(n16762), .A2(n16761), .A3(n16760), .ZN(P3_U2648) );
  AOI211_X1 U20055 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16780), .A(n16763), .B(
        n17030), .ZN(n16764) );
  AOI21_X1 U20056 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17007), .A(n16764), .ZN(
        n16774) );
  NOR2_X1 U20057 ( .A1(n16766), .A2(n16765), .ZN(n16789) );
  AOI211_X1 U20058 ( .C1(n17704), .C2(n16768), .A(n16767), .B(n18842), .ZN(
        n16772) );
  AOI211_X1 U20059 ( .C1(n18905), .C2(n18906), .A(n16770), .B(n16769), .ZN(
        n16771) );
  AOI211_X1 U20060 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n16789), .A(n16772), 
        .B(n16771), .ZN(n16773) );
  OAI211_X1 U20061 ( .C1(n16775), .C2(n16969), .A(n16774), .B(n16773), .ZN(
        P3_U2649) );
  AOI22_X1 U20062 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n17018), .B1(
        n17007), .B2(P3_EBX_REG_21__SCAN_IN), .ZN(n16783) );
  AOI211_X1 U20063 ( .C1(n17718), .C2(n16777), .A(n16776), .B(n18842), .ZN(
        n16778) );
  AOI221_X1 U20064 ( .B1(n16789), .B2(P3_REIP_REG_21__SCAN_IN), .C1(n16779), 
        .C2(n18905), .A(n16778), .ZN(n16782) );
  OAI211_X1 U20065 ( .C1(n16786), .C2(n17134), .A(n17026), .B(n16780), .ZN(
        n16781) );
  NAND3_X1 U20066 ( .A1(n16783), .A2(n16782), .A3(n16781), .ZN(P3_U2650) );
  AOI22_X1 U20067 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17018), .B1(
        n17007), .B2(P3_EBX_REG_20__SCAN_IN), .ZN(n16792) );
  AOI211_X1 U20068 ( .C1(n17740), .C2(n16785), .A(n16784), .B(n18842), .ZN(
        n16788) );
  AOI211_X1 U20069 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16801), .A(n16786), .B(
        n17030), .ZN(n16787) );
  AOI211_X1 U20070 ( .C1(n16789), .C2(P3_REIP_REG_20__SCAN_IN), .A(n16788), 
        .B(n16787), .ZN(n16791) );
  INV_X1 U20071 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18902) );
  NAND3_X1 U20072 ( .A1(n16800), .A2(P3_REIP_REG_19__SCAN_IN), .A3(n18902), 
        .ZN(n16790) );
  NAND3_X1 U20073 ( .A1(n16792), .A2(n16791), .A3(n16790), .ZN(P3_U2651) );
  AOI22_X1 U20074 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n17018), .B1(
        n17007), .B2(P3_EBX_REG_19__SCAN_IN), .ZN(n16805) );
  INV_X1 U20075 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18901) );
  NAND2_X1 U20076 ( .A1(n17032), .A2(n16793), .ZN(n16826) );
  OAI21_X1 U20077 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n16816), .A(n16826), 
        .ZN(n16799) );
  INV_X1 U20078 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17759) );
  NOR2_X1 U20079 ( .A1(n17983), .A2(n17770), .ZN(n16830) );
  NAND2_X1 U20080 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n16830), .ZN(
        n17747) );
  NOR2_X1 U20081 ( .A1(n17759), .A2(n17747), .ZN(n16806) );
  NOR2_X1 U20082 ( .A1(n16807), .A2(n16991), .ZN(n16841) );
  INV_X1 U20083 ( .A(n16841), .ZN(n16831) );
  OAI21_X1 U20084 ( .B1(n16991), .B2(n16806), .A(n16831), .ZN(n16794) );
  INV_X1 U20085 ( .A(n16794), .ZN(n16797) );
  OAI21_X1 U20086 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16806), .A(
        n16795), .ZN(n17748) );
  OAI21_X1 U20087 ( .B1(n16797), .B2(n17748), .A(n17012), .ZN(n16796) );
  AOI21_X1 U20088 ( .B1(n16797), .B2(n17748), .A(n16796), .ZN(n16798) );
  AOI221_X1 U20089 ( .B1(n16800), .B2(n18901), .C1(n16799), .C2(
        P3_REIP_REG_19__SCAN_IN), .A(n16798), .ZN(n16804) );
  OAI211_X1 U20090 ( .C1(n16811), .C2(n16802), .A(n17026), .B(n16801), .ZN(
        n16803) );
  NAND4_X1 U20091 ( .A1(n16805), .A2(n16804), .A3(n18312), .A4(n16803), .ZN(
        P3_U2652) );
  AOI21_X1 U20092 ( .B1(n17759), .B2(n17747), .A(n16806), .ZN(n17767) );
  INV_X1 U20093 ( .A(n17747), .ZN(n16808) );
  AOI21_X1 U20094 ( .B1(n16808), .B2(n16807), .A(n16991), .ZN(n16810) );
  OAI21_X1 U20095 ( .B1(n17767), .B2(n16810), .A(n17012), .ZN(n16809) );
  AOI21_X1 U20096 ( .B1(n17767), .B2(n16810), .A(n16809), .ZN(n16814) );
  AOI211_X1 U20097 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16818), .A(n16811), .B(
        n17030), .ZN(n16813) );
  INV_X1 U20098 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17182) );
  OAI22_X1 U20099 ( .A1(n17759), .A2(n16969), .B1(n17031), .B2(n17182), .ZN(
        n16812) );
  NOR4_X1 U20100 ( .A1(n9822), .A2(n16814), .A3(n16813), .A4(n16812), .ZN(
        n16815) );
  OAI221_X1 U20101 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n16816), .C1(n18898), 
        .C2(n16826), .A(n16815), .ZN(P3_U2653) );
  AOI22_X1 U20102 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n17018), .B1(
        n17007), .B2(P3_EBX_REG_17__SCAN_IN), .ZN(n16825) );
  NOR2_X1 U20103 ( .A1(n16836), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n16823) );
  OAI21_X1 U20104 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16830), .A(
        n17747), .ZN(n17771) );
  INV_X1 U20105 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16992) );
  NAND2_X1 U20106 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16992), .ZN(
        n16977) );
  OAI21_X1 U20107 ( .B1(n17770), .B2(n16977), .A(n16959), .ZN(n16817) );
  XNOR2_X1 U20108 ( .A(n17771), .B(n16817), .ZN(n16821) );
  OAI211_X1 U20109 ( .C1(n16829), .C2(n16819), .A(n17026), .B(n16818), .ZN(
        n16820) );
  OAI211_X1 U20110 ( .C1(n18842), .C2(n16821), .A(n18312), .B(n16820), .ZN(
        n16822) );
  AOI21_X1 U20111 ( .B1(n16823), .B2(n16845), .A(n16822), .ZN(n16824) );
  OAI211_X1 U20112 ( .C1(n18896), .C2(n16826), .A(n16825), .B(n16824), .ZN(
        P3_U2654) );
  INV_X1 U20113 ( .A(n16827), .ZN(n16828) );
  AOI21_X1 U20114 ( .B1(n17009), .B2(n16828), .A(n16973), .ZN(n16851) );
  INV_X1 U20115 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18894) );
  AOI211_X1 U20116 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16846), .A(n16829), .B(
        n17030), .ZN(n16835) );
  INV_X1 U20117 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17784) );
  AOI21_X1 U20118 ( .B1(n17784), .B2(n16839), .A(n16830), .ZN(n17788) );
  INV_X1 U20119 ( .A(n17788), .ZN(n16832) );
  OAI221_X1 U20120 ( .B1(n17788), .B2(n16841), .C1(n16832), .C2(n16831), .A(
        n17012), .ZN(n16833) );
  OAI211_X1 U20121 ( .C1(n17784), .C2(n16969), .A(n18312), .B(n16833), .ZN(
        n16834) );
  AOI211_X1 U20122 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17007), .A(n16835), .B(
        n16834), .ZN(n16838) );
  OAI211_X1 U20123 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(P3_REIP_REG_15__SCAN_IN), .A(n16845), .B(n16836), .ZN(n16837) );
  OAI211_X1 U20124 ( .C1(n16851), .C2(n18894), .A(n16838), .B(n16837), .ZN(
        P3_U2655) );
  INV_X1 U20125 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18892) );
  OAI21_X1 U20126 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17787), .A(
        n16839), .ZN(n17800) );
  NAND2_X1 U20127 ( .A1(n16959), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16911) );
  NAND2_X1 U20128 ( .A1(n17012), .A2(n16911), .ZN(n17028) );
  AOI211_X1 U20129 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n16959), .A(
        n17800), .B(n17028), .ZN(n16840) );
  AOI211_X1 U20130 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n17018), .A(
        n9822), .B(n16840), .ZN(n16843) );
  NAND3_X1 U20131 ( .A1(n17012), .A2(n16841), .A3(n17800), .ZN(n16842) );
  OAI211_X1 U20132 ( .C1(n16851), .C2(n18892), .A(n16843), .B(n16842), .ZN(
        n16844) );
  AOI21_X1 U20133 ( .B1(n16845), .B2(n18892), .A(n16844), .ZN(n16848) );
  OAI211_X1 U20134 ( .C1(n16853), .C2(n16849), .A(n17026), .B(n16846), .ZN(
        n16847) );
  OAI211_X1 U20135 ( .C1(n16849), .C2(n17031), .A(n16848), .B(n16847), .ZN(
        P3_U2656) );
  INV_X1 U20136 ( .A(n17811), .ZN(n17835) );
  NOR2_X1 U20137 ( .A1(n17835), .A2(n17823), .ZN(n16859) );
  AOI21_X1 U20138 ( .B1(n16859), .B2(n16992), .A(n16991), .ZN(n16860) );
  INV_X1 U20139 ( .A(n17787), .ZN(n16850) );
  OAI21_X1 U20140 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16859), .A(
        n16850), .ZN(n17812) );
  XOR2_X1 U20141 ( .A(n16860), .B(n17812), .Z(n16858) );
  AOI21_X1 U20142 ( .B1(n17007), .B2(P3_EBX_REG_14__SCAN_IN), .A(n9822), .ZN(
        n16857) );
  AOI21_X1 U20143 ( .B1(n18891), .B2(n16852), .A(n16851), .ZN(n16855) );
  AOI211_X1 U20144 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16865), .A(n16853), .B(
        n17030), .ZN(n16854) );
  AOI211_X1 U20145 ( .C1(n17018), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16855), .B(n16854), .ZN(n16856) );
  OAI211_X1 U20146 ( .C1(n18842), .C2(n16858), .A(n16857), .B(n16856), .ZN(
        P3_U2657) );
  INV_X1 U20147 ( .A(n17823), .ZN(n16879) );
  NAND2_X1 U20148 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16879), .ZN(
        n16878) );
  AOI21_X1 U20149 ( .B1(n16868), .B2(n16878), .A(n16859), .ZN(n17826) );
  INV_X1 U20150 ( .A(n17826), .ZN(n16861) );
  AND3_X1 U20151 ( .A1(n16861), .A2(n17012), .A3(n16860), .ZN(n16871) );
  AOI211_X1 U20152 ( .C1(n16959), .C2(n16878), .A(n16861), .B(n17028), .ZN(
        n16870) );
  NAND3_X1 U20153 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(P3_REIP_REG_10__SCAN_IN), 
        .A3(P3_REIP_REG_9__SCAN_IN), .ZN(n16863) );
  NAND2_X1 U20154 ( .A1(n16862), .A2(n17034), .ZN(n16896) );
  OAI21_X1 U20155 ( .B1(n16863), .B2(n16896), .A(n17032), .ZN(n16890) );
  INV_X1 U20156 ( .A(n16890), .ZN(n16864) );
  NOR2_X1 U20157 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17023), .ZN(n16882) );
  OAI21_X1 U20158 ( .B1(n16864), .B2(n16882), .A(P3_REIP_REG_13__SCAN_IN), 
        .ZN(n16867) );
  OAI211_X1 U20159 ( .C1(n16876), .C2(n16875), .A(n17026), .B(n16865), .ZN(
        n16866) );
  OAI211_X1 U20160 ( .C1(n16969), .C2(n16868), .A(n16867), .B(n16866), .ZN(
        n16869) );
  NOR4_X1 U20161 ( .A1(n9822), .A2(n16871), .A3(n16870), .A4(n16869), .ZN(
        n16874) );
  INV_X1 U20162 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18888) );
  NAND3_X1 U20163 ( .A1(n17009), .A2(n16872), .A3(n18888), .ZN(n16873) );
  OAI211_X1 U20164 ( .C1(n16875), .C2(n17031), .A(n16874), .B(n16873), .ZN(
        P3_U2658) );
  AOI211_X1 U20165 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16893), .A(n16876), .B(
        n17030), .ZN(n16886) );
  INV_X1 U20166 ( .A(n16877), .ZN(n16883) );
  OAI21_X1 U20167 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n16879), .A(
        n16878), .ZN(n17840) );
  OAI21_X1 U20168 ( .B1(n17833), .B2(n16977), .A(n16959), .ZN(n16880) );
  XOR2_X1 U20169 ( .A(n17840), .B(n16880), .Z(n16881) );
  AOI22_X1 U20170 ( .A1(n16883), .A2(n16882), .B1(n17012), .B2(n16881), .ZN(
        n16884) );
  OAI211_X1 U20171 ( .C1(n17844), .C2(n16969), .A(n16884), .B(n18312), .ZN(
        n16885) );
  AOI211_X1 U20172 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17007), .A(n16886), .B(
        n16885), .ZN(n16887) );
  OAI21_X1 U20173 ( .B1(n18886), .B2(n16890), .A(n16887), .ZN(P3_U2659) );
  INV_X1 U20174 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18882) );
  INV_X1 U20175 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18880) );
  NOR2_X1 U20176 ( .A1(n18882), .A2(n18880), .ZN(n16904) );
  NOR3_X1 U20177 ( .A1(n17023), .A2(n18879), .A3(n16924), .ZN(n16903) );
  AOI21_X1 U20178 ( .B1(n16904), .B2(n16903), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16891) );
  NAND3_X1 U20179 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(n16935), .ZN(n16898) );
  NOR2_X1 U20180 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16898), .ZN(
        n16899) );
  AOI21_X1 U20181 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16899), .A(
        n16991), .ZN(n16888) );
  INV_X1 U20182 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17865) );
  NOR2_X1 U20183 ( .A1(n17865), .A2(n16898), .ZN(n16897) );
  OAI21_X1 U20184 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16897), .A(
        n17823), .ZN(n17856) );
  XOR2_X1 U20185 ( .A(n16888), .B(n17856), .Z(n16889) );
  OAI22_X1 U20186 ( .A1(n16891), .A2(n16890), .B1(n18842), .B2(n16889), .ZN(
        n16892) );
  AOI211_X1 U20187 ( .C1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n17018), .A(
        n9822), .B(n16892), .ZN(n16895) );
  OAI211_X1 U20188 ( .C1(n16905), .C2(n17250), .A(n17026), .B(n16893), .ZN(
        n16894) );
  OAI211_X1 U20189 ( .C1(n17250), .C2(n17031), .A(n16895), .B(n16894), .ZN(
        P3_U2660) );
  NAND2_X1 U20190 ( .A1(n17032), .A2(n16896), .ZN(n16923) );
  AOI21_X1 U20191 ( .B1(n17865), .B2(n16898), .A(n16897), .ZN(n17868) );
  NOR2_X1 U20192 ( .A1(n16899), .A2(n16991), .ZN(n16901) );
  INV_X1 U20193 ( .A(n17868), .ZN(n16900) );
  INV_X1 U20194 ( .A(n16901), .ZN(n16914) );
  AOI221_X1 U20195 ( .B1(n17868), .B2(n16901), .C1(n16900), .C2(n16914), .A(
        n18842), .ZN(n16902) );
  AOI211_X1 U20196 ( .C1(n17007), .C2(P3_EBX_REG_10__SCAN_IN), .A(n9822), .B(
        n16902), .ZN(n16910) );
  INV_X1 U20197 ( .A(n16903), .ZN(n16922) );
  AOI211_X1 U20198 ( .C1(n18882), .C2(n18880), .A(n16904), .B(n16922), .ZN(
        n16908) );
  AOI211_X1 U20199 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16906), .A(n16905), .B(
        n17030), .ZN(n16907) );
  AOI211_X1 U20200 ( .C1(n17018), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16908), .B(n16907), .ZN(n16909) );
  OAI211_X1 U20201 ( .C1(n18882), .C2(n16923), .A(n16910), .B(n16909), .ZN(
        P3_U2661) );
  NOR2_X1 U20202 ( .A1(n16915), .A2(n17030), .ZN(n16931) );
  NAND2_X1 U20203 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16935), .ZN(
        n16926) );
  XOR2_X1 U20204 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n16926), .Z(n17880) );
  INV_X1 U20205 ( .A(n16926), .ZN(n16912) );
  NOR2_X1 U20206 ( .A1(n16959), .A2(n18842), .ZN(n17002) );
  INV_X1 U20207 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16917) );
  OAI33_X1 U20208 ( .A1(n16912), .A2(n17002), .A3(n16917), .B1(n16926), .B2(
        n16911), .B3(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16913) );
  AOI211_X1 U20209 ( .C1(n17880), .C2(n16914), .A(n18842), .B(n16913), .ZN(
        n16919) );
  OAI221_X1 U20210 ( .B1(n17007), .B2(n17026), .C1(n17007), .C2(n16915), .A(
        P3_EBX_REG_9__SCAN_IN), .ZN(n16916) );
  OAI211_X1 U20211 ( .C1(n16917), .C2(n16969), .A(n18312), .B(n16916), .ZN(
        n16918) );
  AOI211_X1 U20212 ( .C1(n16931), .C2(n16920), .A(n16919), .B(n16918), .ZN(
        n16921) );
  OAI221_X1 U20213 ( .B1(P3_REIP_REG_9__SCAN_IN), .B2(n16922), .C1(n18880), 
        .C2(n16923), .A(n16921), .ZN(P3_U2662) );
  NAND2_X1 U20214 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16943), .ZN(n16930) );
  AOI221_X1 U20215 ( .B1(n17023), .B2(n18879), .C1(n16924), .C2(n18879), .A(
        n16923), .ZN(n16929) );
  INV_X1 U20216 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17888) );
  INV_X1 U20217 ( .A(n16925), .ZN(n17887) );
  INV_X1 U20218 ( .A(n16977), .ZN(n17013) );
  NAND2_X1 U20219 ( .A1(n17887), .A2(n17013), .ZN(n16936) );
  INV_X1 U20220 ( .A(n16936), .ZN(n16951) );
  AOI21_X1 U20221 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16951), .A(
        n16991), .ZN(n16938) );
  OAI21_X1 U20222 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16935), .A(
        n16926), .ZN(n17891) );
  XOR2_X1 U20223 ( .A(n16938), .B(n17891), .Z(n16927) );
  OAI22_X1 U20224 ( .A1(n17888), .A2(n16969), .B1(n18842), .B2(n16927), .ZN(
        n16928) );
  AOI211_X1 U20225 ( .C1(n16931), .C2(n16930), .A(n16929), .B(n16928), .ZN(
        n16932) );
  OAI211_X1 U20226 ( .C1(n17031), .C2(n16933), .A(n16932), .B(n18312), .ZN(
        P3_U2663) );
  INV_X1 U20227 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18876) );
  AND3_X1 U20228 ( .A1(n17009), .A2(n16934), .A3(n18876), .ZN(n16942) );
  AOI221_X1 U20229 ( .B1(n18874), .B2(n17009), .C1(n16958), .C2(n17009), .A(
        n16973), .ZN(n16940) );
  NAND2_X1 U20230 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17919), .ZN(
        n16961) );
  INV_X1 U20231 ( .A(n16961), .ZN(n16948) );
  NAND2_X1 U20232 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16948), .ZN(
        n16947) );
  AOI21_X1 U20233 ( .B1(n17903), .B2(n16947), .A(n16935), .ZN(n17909) );
  AOI21_X1 U20234 ( .B1(n17909), .B2(n16936), .A(n18842), .ZN(n16937) );
  OAI22_X1 U20235 ( .A1(n17909), .A2(n16938), .B1(n17002), .B2(n16937), .ZN(
        n16939) );
  OAI211_X1 U20236 ( .C1(n16940), .C2(n18876), .A(n18312), .B(n16939), .ZN(
        n16941) );
  AOI211_X1 U20237 ( .C1(n17018), .C2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n16942), .B(n16941), .ZN(n16945) );
  OAI211_X1 U20238 ( .C1(n16946), .C2(n17331), .A(n17026), .B(n16943), .ZN(
        n16944) );
  OAI211_X1 U20239 ( .C1(n17331), .C2(n17031), .A(n16945), .B(n16944), .ZN(
        P3_U2664) );
  AOI21_X1 U20240 ( .B1(n17009), .B2(n16958), .A(n16973), .ZN(n16972) );
  AOI22_X1 U20241 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17018), .B1(
        n17007), .B2(P3_EBX_REG_6__SCAN_IN), .ZN(n16957) );
  NOR3_X1 U20242 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n17023), .A3(n16958), .ZN(
        n16955) );
  AOI211_X1 U20243 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16965), .A(n16946), .B(
        n17030), .ZN(n16954) );
  OAI21_X1 U20244 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16948), .A(
        n16947), .ZN(n17923) );
  AOI211_X1 U20245 ( .C1(n16959), .C2(n16961), .A(n17923), .B(n17028), .ZN(
        n16953) );
  NOR2_X1 U20246 ( .A1(n16991), .A2(n18842), .ZN(n17019) );
  NAND2_X1 U20247 ( .A1(n17923), .A2(n17019), .ZN(n16950) );
  OAI21_X1 U20248 ( .B1(n16951), .B2(n16950), .A(n18312), .ZN(n16952) );
  NOR4_X1 U20249 ( .A1(n16955), .A2(n16954), .A3(n16953), .A4(n16952), .ZN(
        n16956) );
  OAI211_X1 U20250 ( .C1(n16972), .C2(n18874), .A(n16957), .B(n16956), .ZN(
        P3_U2665) );
  INV_X1 U20251 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18872) );
  AND2_X1 U20252 ( .A1(n16958), .A2(n17009), .ZN(n16963) );
  NOR2_X1 U20253 ( .A1(n17983), .A2(n17931), .ZN(n16975) );
  INV_X1 U20254 ( .A(n16975), .ZN(n16960) );
  OAI21_X1 U20255 ( .B1(n16960), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n16959), .ZN(n16978) );
  OAI21_X1 U20256 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n16975), .A(
        n16961), .ZN(n17935) );
  XOR2_X1 U20257 ( .A(n16978), .B(n17935), .Z(n16962) );
  AOI22_X1 U20258 ( .A1(n16964), .A2(n16963), .B1(n17012), .B2(n16962), .ZN(
        n16968) );
  OAI211_X1 U20259 ( .C1(n16974), .C2(n16966), .A(n17026), .B(n16965), .ZN(
        n16967) );
  OAI211_X1 U20260 ( .C1(n16969), .C2(n17930), .A(n16968), .B(n16967), .ZN(
        n16970) );
  AOI211_X1 U20261 ( .C1(n17007), .C2(P3_EBX_REG_5__SCAN_IN), .A(n9822), .B(
        n16970), .ZN(n16971) );
  OAI21_X1 U20262 ( .B1(n16972), .B2(n18872), .A(n16971), .ZN(P3_U2666) );
  AOI21_X1 U20263 ( .B1(n17009), .B2(n16989), .A(n16973), .ZN(n16987) );
  AOI22_X1 U20264 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17018), .B1(
        n17007), .B2(P3_EBX_REG_4__SCAN_IN), .ZN(n16986) );
  AOI211_X1 U20265 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16998), .A(n16974), .B(
        n17030), .ZN(n16984) );
  NOR3_X1 U20266 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17023), .A3(n16989), .ZN(
        n16983) );
  NAND2_X1 U20267 ( .A1(n18336), .A2(n19008), .ZN(n17037) );
  INV_X1 U20268 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n16976) );
  NAND2_X1 U20269 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17949), .ZN(
        n16990) );
  AOI21_X1 U20270 ( .B1(n16976), .B2(n16990), .A(n16975), .ZN(n17950) );
  NAND2_X1 U20271 ( .A1(n17949), .A2(n16976), .ZN(n17946) );
  OAI22_X1 U20272 ( .A1(n17950), .A2(n16978), .B1(n16977), .B2(n17946), .ZN(
        n16979) );
  AOI22_X1 U20273 ( .A1(n17012), .A2(n16979), .B1(n17950), .B2(n17002), .ZN(
        n16980) );
  OAI221_X1 U20274 ( .B1(n17037), .B2(n17312), .C1(n17037), .C2(n16981), .A(
        n16980), .ZN(n16982) );
  NOR4_X1 U20275 ( .A1(n9822), .A2(n16984), .A3(n16983), .A4(n16982), .ZN(
        n16985) );
  OAI211_X1 U20276 ( .C1(n16987), .C2(n18870), .A(n16986), .B(n16985), .ZN(
        P3_U2667) );
  INV_X1 U20277 ( .A(n16987), .ZN(n16997) );
  INV_X1 U20278 ( .A(n17037), .ZN(n19010) );
  INV_X1 U20279 ( .A(n18789), .ZN(n17004) );
  AOI21_X1 U20280 ( .B1(n11435), .B2(n17004), .A(n17292), .ZN(n18947) );
  AOI22_X1 U20281 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n17018), .B1(
        n19010), .B2(n18947), .ZN(n16988) );
  INV_X1 U20282 ( .A(n16988), .ZN(n16996) );
  NAND2_X1 U20283 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n17008) );
  NAND2_X1 U20284 ( .A1(n17009), .A2(n16989), .ZN(n16994) );
  INV_X1 U20285 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17976) );
  NOR2_X1 U20286 ( .A1(n17983), .A2(n17976), .ZN(n17001) );
  OAI21_X1 U20287 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17001), .A(
        n16990), .ZN(n17961) );
  AOI21_X1 U20288 ( .B1(n16992), .B2(n17001), .A(n16991), .ZN(n17011) );
  XOR2_X1 U20289 ( .A(n17961), .B(n17011), .Z(n16993) );
  OAI22_X1 U20290 ( .A1(n17008), .A2(n16994), .B1(n18842), .B2(n16993), .ZN(
        n16995) );
  AOI211_X1 U20291 ( .C1(P3_REIP_REG_3__SCAN_IN), .C2(n16997), .A(n16996), .B(
        n16995), .ZN(n17000) );
  OAI211_X1 U20292 ( .C1(n17003), .C2(n17341), .A(n17026), .B(n16998), .ZN(
        n16999) );
  OAI211_X1 U20293 ( .C1(n17341), .C2(n17031), .A(n17000), .B(n16999), .ZN(
        P3_U2668) );
  AOI21_X1 U20294 ( .B1(n17983), .B2(n17976), .A(n17001), .ZN(n17010) );
  AOI22_X1 U20295 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n17018), .B1(
        n17002), .B2(n17010), .ZN(n17017) );
  OR2_X1 U20296 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), .ZN(
        n17020) );
  AOI211_X1 U20297 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17020), .A(n17003), .B(
        n17030), .ZN(n17006) );
  INV_X1 U20298 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18866) );
  NAND2_X1 U20299 ( .A1(n10256), .A2(n18807), .ZN(n18790) );
  NAND2_X1 U20300 ( .A1(n17004), .A2(n18790), .ZN(n18953) );
  OAI22_X1 U20301 ( .A1(n18866), .A2(n17034), .B1(n18953), .B2(n17037), .ZN(
        n17005) );
  AOI211_X1 U20302 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17007), .A(n17006), .B(
        n17005), .ZN(n17016) );
  OAI211_X1 U20303 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n17009), .B(n17008), .ZN(n17015) );
  INV_X1 U20304 ( .A(n17010), .ZN(n17972) );
  OAI211_X1 U20305 ( .C1(n17013), .C2(n17972), .A(n17012), .B(n17011), .ZN(
        n17014) );
  NAND4_X1 U20306 ( .A1(n17017), .A2(n17016), .A3(n17015), .A4(n17014), .ZN(
        P3_U2669) );
  AOI211_X1 U20307 ( .C1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n17019), .A(
        n17018), .B(n17983), .ZN(n17029) );
  AND2_X1 U20308 ( .A1(n17020), .A2(n17350), .ZN(n17356) );
  NAND2_X1 U20309 ( .A1(n17021), .A2(n18807), .ZN(n18958) );
  OAI22_X1 U20310 ( .A1(n18974), .A2(n17034), .B1(n18958), .B2(n17037), .ZN(
        n17025) );
  INV_X1 U20311 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17022) );
  OAI22_X1 U20312 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17023), .B1(n17031), 
        .B2(n17022), .ZN(n17024) );
  AOI211_X1 U20313 ( .C1(n17026), .C2(n17356), .A(n17025), .B(n17024), .ZN(
        n17027) );
  OAI221_X1 U20314 ( .B1(n17029), .B2(n17983), .C1(n17029), .C2(n17028), .A(
        n17027), .ZN(P3_U2670) );
  NAND2_X1 U20315 ( .A1(n17031), .A2(n17030), .ZN(n17033) );
  AOI22_X1 U20316 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n17033), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n17032), .ZN(n17036) );
  NAND3_X1 U20317 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18944), .A3(
        n17034), .ZN(n17035) );
  OAI211_X1 U20318 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n17037), .A(
        n17036), .B(n17035), .ZN(P3_U2671) );
  NOR4_X1 U20319 ( .A1(n17040), .A2(n17039), .A3(n17038), .A4(n17134), .ZN(
        n17045) );
  NAND2_X1 U20320 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n17041) );
  NOR4_X1 U20321 ( .A1(n17082), .A2(n17043), .A3(n17042), .A4(n17041), .ZN(
        n17044) );
  NAND4_X1 U20322 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17166), .A3(n17045), 
        .A4(n17044), .ZN(n17048) );
  NOR2_X1 U20323 ( .A1(n17049), .A2(n17048), .ZN(n17077) );
  NAND2_X1 U20324 ( .A1(n17358), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17047) );
  NAND2_X1 U20325 ( .A1(n17077), .A2(n18366), .ZN(n17046) );
  OAI22_X1 U20326 ( .A1(n17077), .A2(n17047), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17046), .ZN(P3_U2672) );
  NAND2_X1 U20327 ( .A1(n17049), .A2(n17048), .ZN(n17050) );
  NAND2_X1 U20328 ( .A1(n17050), .A2(n17358), .ZN(n17076) );
  INV_X1 U20329 ( .A(n17084), .ZN(n17078) );
  AOI22_X1 U20330 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17292), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17061) );
  AOI22_X1 U20331 ( .A1(n17309), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17052) );
  AOI22_X1 U20332 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17051) );
  OAI211_X1 U20333 ( .C1(n11467), .C2(n17053), .A(n17052), .B(n17051), .ZN(
        n17059) );
  AOI22_X1 U20334 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17057) );
  AOI22_X1 U20335 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17056) );
  AOI22_X1 U20336 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17273), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17055) );
  NAND2_X1 U20337 ( .A1(n11474), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n17054) );
  NAND4_X1 U20338 ( .A1(n17057), .A2(n17056), .A3(n17055), .A4(n17054), .ZN(
        n17058) );
  AOI211_X1 U20339 ( .C1(n11444), .C2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A(
        n17059), .B(n17058), .ZN(n17060) );
  OAI211_X1 U20340 ( .C1(n17197), .C2(n18387), .A(n17061), .B(n17060), .ZN(
        n17081) );
  NAND3_X1 U20341 ( .A1(n17079), .A2(n17078), .A3(n17081), .ZN(n17075) );
  AOI22_X1 U20342 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17062) );
  OAI21_X1 U20343 ( .B1(n11523), .B2(n17063), .A(n17062), .ZN(n17073) );
  AOI22_X1 U20344 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17309), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17070) );
  AOI22_X1 U20345 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17292), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17064) );
  OAI21_X1 U20346 ( .B1(n17197), .B2(n17218), .A(n17064), .ZN(n17068) );
  INV_X1 U20347 ( .A(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17216) );
  AOI22_X1 U20348 ( .A1(n17285), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17273), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17066) );
  AOI22_X1 U20349 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17065) );
  OAI211_X1 U20350 ( .C1(n11467), .C2(n17216), .A(n17066), .B(n17065), .ZN(
        n17067) );
  AOI211_X1 U20351 ( .C1(n11444), .C2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n17068), .B(n17067), .ZN(n17069) );
  OAI211_X1 U20352 ( .C1(n11447), .C2(n17071), .A(n17070), .B(n17069), .ZN(
        n17072) );
  AOI211_X1 U20353 ( .C1(n17245), .C2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n17073), .B(n17072), .ZN(n17074) );
  XNOR2_X1 U20354 ( .A(n17075), .B(n17074), .ZN(n17375) );
  OAI22_X1 U20355 ( .A1(n17077), .A2(n17076), .B1(n17375), .B2(n17358), .ZN(
        P3_U2673) );
  NAND2_X1 U20356 ( .A1(n17079), .A2(n17078), .ZN(n17080) );
  XOR2_X1 U20357 ( .A(n17081), .B(n17080), .Z(n17379) );
  OAI21_X1 U20358 ( .B1(n17086), .B2(n17085), .A(n17084), .ZN(n17388) );
  NAND3_X1 U20359 ( .A1(n17088), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n17358), 
        .ZN(n17087) );
  OAI221_X1 U20360 ( .B1(n17088), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n17358), 
        .C2(n17388), .A(n17087), .ZN(P3_U2676) );
  AOI21_X1 U20361 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17358), .A(n17096), .ZN(
        n17090) );
  XNOR2_X1 U20362 ( .A(n17089), .B(n17092), .ZN(n17393) );
  OAI22_X1 U20363 ( .A1(n17091), .A2(n17090), .B1(n17358), .B2(n17393), .ZN(
        P3_U2677) );
  AOI21_X1 U20364 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17358), .A(n17100), .ZN(
        n17095) );
  OAI21_X1 U20365 ( .B1(n17094), .B2(n17093), .A(n17092), .ZN(n17398) );
  OAI22_X1 U20366 ( .A1(n17096), .A2(n17095), .B1(n17358), .B2(n17398), .ZN(
        P3_U2678) );
  INV_X1 U20367 ( .A(n17097), .ZN(n17106) );
  AOI21_X1 U20368 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17358), .A(n17106), .ZN(
        n17099) );
  XNOR2_X1 U20369 ( .A(n17098), .B(n17102), .ZN(n17403) );
  OAI22_X1 U20370 ( .A1(n17100), .A2(n17099), .B1(n17358), .B2(n17403), .ZN(
        P3_U2679) );
  AOI21_X1 U20371 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17358), .A(n17101), .ZN(
        n17105) );
  OAI21_X1 U20372 ( .B1(n17104), .B2(n17103), .A(n17102), .ZN(n17408) );
  OAI22_X1 U20373 ( .A1(n17106), .A2(n17105), .B1(n17358), .B2(n17408), .ZN(
        P3_U2680) );
  AOI22_X1 U20374 ( .A1(n17304), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17107) );
  OAI21_X1 U20375 ( .B1(n17288), .B2(n17108), .A(n17107), .ZN(n17118) );
  AOI22_X1 U20376 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17116) );
  OAI21_X1 U20377 ( .B1(n11447), .B2(n17110), .A(n17109), .ZN(n17114) );
  AOI22_X1 U20378 ( .A1(n17309), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17112) );
  AOI22_X1 U20379 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17273), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17111) );
  OAI211_X1 U20380 ( .C1(n11448), .C2(n18387), .A(n17112), .B(n17111), .ZN(
        n17113) );
  AOI211_X1 U20381 ( .C1(n17292), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n17114), .B(n17113), .ZN(n17115) );
  OAI211_X1 U20382 ( .C1(n17197), .C2(n17333), .A(n17116), .B(n17115), .ZN(
        n17117) );
  AOI211_X1 U20383 ( .C1(n17245), .C2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n17118), .B(n17117), .ZN(n17411) );
  NAND3_X1 U20384 ( .A1(n17120), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n17358), 
        .ZN(n17119) );
  OAI221_X1 U20385 ( .B1(n17120), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n17358), 
        .C2(n17411), .A(n17119), .ZN(P3_U2681) );
  AOI22_X1 U20386 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17285), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17121) );
  OAI21_X1 U20387 ( .B1(n11479), .B2(n17122), .A(n17121), .ZN(n17133) );
  OAI22_X1 U20388 ( .A1(n11447), .A2(n17124), .B1(n9856), .B2(n17123), .ZN(
        n17129) );
  AOI22_X1 U20389 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17127) );
  AOI22_X1 U20390 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17126) );
  AOI22_X1 U20391 ( .A1(n17292), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17125) );
  NAND3_X1 U20392 ( .A1(n17127), .A2(n17126), .A3(n17125), .ZN(n17128) );
  AOI211_X1 U20393 ( .C1(n17245), .C2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A(
        n17129), .B(n17128), .ZN(n17130) );
  OAI211_X1 U20394 ( .C1(n17197), .C2(n17339), .A(n17131), .B(n17130), .ZN(
        n17132) );
  AOI211_X1 U20395 ( .C1(n17219), .C2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A(
        n17133), .B(n17132), .ZN(n17417) );
  AOI21_X1 U20396 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17166), .A(n17361), .ZN(
        n17148) );
  AOI22_X1 U20397 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17148), .B1(n17135), 
        .B2(n17134), .ZN(n17136) );
  OAI21_X1 U20398 ( .B1(n17417), .B2(n17358), .A(n17136), .ZN(P3_U2682) );
  AOI22_X1 U20399 ( .A1(n9811), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17137) );
  OAI21_X1 U20400 ( .B1(n9890), .B2(n17236), .A(n17137), .ZN(n17147) );
  AOI22_X1 U20401 ( .A1(n17309), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17145) );
  OAI22_X1 U20402 ( .A1(n11447), .A2(n17232), .B1(n11467), .B2(n17138), .ZN(
        n17143) );
  AOI22_X1 U20403 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17141) );
  AOI22_X1 U20404 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17140) );
  AOI22_X1 U20405 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17292), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17139) );
  NAND3_X1 U20406 ( .A1(n17141), .A2(n17140), .A3(n17139), .ZN(n17142) );
  AOI211_X1 U20407 ( .C1(n11444), .C2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n17143), .B(n17142), .ZN(n17144) );
  OAI211_X1 U20408 ( .C1(n17197), .C2(n17343), .A(n17145), .B(n17144), .ZN(
        n17146) );
  AOI211_X1 U20409 ( .C1(n17219), .C2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n17147), .B(n17146), .ZN(n17420) );
  OAI21_X1 U20410 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17149), .A(n17148), .ZN(
        n17150) );
  OAI21_X1 U20411 ( .B1(n17420), .B2(n17358), .A(n17150), .ZN(P3_U2683) );
  INV_X1 U20412 ( .A(n17167), .ZN(n17151) );
  OAI21_X1 U20413 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17151), .A(n17358), .ZN(
        n17165) );
  AOI22_X1 U20414 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17309), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17152) );
  OAI21_X1 U20415 ( .B1(n17288), .B2(n17153), .A(n17152), .ZN(n17164) );
  AOI22_X1 U20416 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17162) );
  INV_X1 U20417 ( .A(n17155), .ZN(n17160) );
  AOI22_X1 U20418 ( .A1(n17304), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17273), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17158) );
  AOI22_X1 U20419 ( .A1(n17211), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17157) );
  AOI22_X1 U20420 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17292), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17156) );
  NAND3_X1 U20421 ( .A1(n17158), .A2(n17157), .A3(n17156), .ZN(n17159) );
  AOI211_X1 U20422 ( .C1(n11474), .C2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A(
        n17160), .B(n17159), .ZN(n17161) );
  OAI211_X1 U20423 ( .C1(n17197), .C2(n17347), .A(n17162), .B(n17161), .ZN(
        n17163) );
  AOI211_X1 U20424 ( .C1(n17245), .C2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A(
        n17164), .B(n17163), .ZN(n17430) );
  OAI22_X1 U20425 ( .A1(n17166), .A2(n17165), .B1(n17430), .B2(n17358), .ZN(
        P3_U2684) );
  NAND2_X1 U20426 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17167), .ZN(n17184) );
  AOI22_X1 U20427 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17168) );
  OAI21_X1 U20428 ( .B1(n17170), .B2(n17169), .A(n17168), .ZN(n17181) );
  AOI22_X1 U20429 ( .A1(n17310), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17309), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17178) );
  INV_X1 U20430 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17172) );
  OAI21_X1 U20431 ( .B1(n11467), .B2(n17172), .A(n17171), .ZN(n17176) );
  AOI22_X1 U20432 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17285), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17174) );
  AOI22_X1 U20433 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17173) );
  OAI211_X1 U20434 ( .C1(n11448), .C2(n17272), .A(n17174), .B(n17173), .ZN(
        n17175) );
  AOI211_X1 U20435 ( .C1(n17292), .C2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n17176), .B(n17175), .ZN(n17177) );
  OAI211_X1 U20436 ( .C1(n17288), .C2(n17179), .A(n17178), .B(n17177), .ZN(
        n17180) );
  AOI211_X1 U20437 ( .C1(n17245), .C2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n17181), .B(n17180), .ZN(n17435) );
  NAND4_X1 U20438 ( .A1(n18366), .A2(P3_EBX_REG_17__SCAN_IN), .A3(n17185), 
        .A4(n17182), .ZN(n17183) );
  OAI221_X1 U20439 ( .B1(n17361), .B2(n17184), .C1(n17358), .C2(n17435), .A(
        n17183), .ZN(P3_U2685) );
  NAND2_X1 U20440 ( .A1(n18366), .A2(n17185), .ZN(n17199) );
  NOR2_X1 U20441 ( .A1(n17361), .A2(n17185), .ZN(n17212) );
  AOI22_X1 U20442 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17200), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17196) );
  INV_X1 U20443 ( .A(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17188) );
  AOI22_X1 U20444 ( .A1(n17309), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17187) );
  AOI22_X1 U20445 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17291), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17186) );
  OAI211_X1 U20446 ( .C1(n11467), .C2(n17188), .A(n17187), .B(n17186), .ZN(
        n17194) );
  AOI22_X1 U20447 ( .A1(n17285), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17192) );
  AOI22_X1 U20448 ( .A1(n17304), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17273), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17191) );
  AOI22_X1 U20449 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17292), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17190) );
  NAND4_X1 U20450 ( .A1(n17192), .A2(n17191), .A3(n17190), .A4(n17189), .ZN(
        n17193) );
  AOI211_X1 U20451 ( .C1(n17293), .C2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A(
        n17194), .B(n17193), .ZN(n17195) );
  OAI211_X1 U20452 ( .C1(n17197), .C2(n17359), .A(n17196), .B(n17195), .ZN(
        n17436) );
  AOI22_X1 U20453 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17212), .B1(n17361), 
        .B2(n17436), .ZN(n17198) );
  OAI21_X1 U20454 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n17199), .A(n17198), .ZN(
        P3_U2686) );
  INV_X1 U20455 ( .A(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17322) );
  OAI22_X1 U20456 ( .A1(n17322), .A2(n9888), .B1(n17317), .B2(n17197), .ZN(
        n17210) );
  AOI22_X1 U20457 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17200), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17208) );
  AOI22_X1 U20458 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__0__SCAN_IN), .B2(n17325), .ZN(n17207) );
  OAI22_X1 U20459 ( .A1(n11448), .A2(n18373), .B1(n17312), .B2(n18396), .ZN(
        n17205) );
  AOI22_X1 U20460 ( .A1(n17304), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17309), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17203) );
  AOI22_X1 U20461 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n17284), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17202) );
  NAND3_X1 U20462 ( .A1(n17203), .A2(n17202), .A3(n17201), .ZN(n17204) );
  AOI211_X1 U20463 ( .C1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .C2(n11474), .A(
        n17205), .B(n17204), .ZN(n17206) );
  NAND3_X1 U20464 ( .A1(n17208), .A2(n17207), .A3(n17206), .ZN(n17209) );
  AOI211_X1 U20465 ( .C1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .C2(n17211), .A(
        n17210), .B(n17209), .ZN(n17447) );
  OAI21_X1 U20466 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17213), .A(n17212), .ZN(
        n17214) );
  OAI21_X1 U20467 ( .B1(n17447), .B2(n17358), .A(n17214), .ZN(P3_U2687) );
  AOI22_X1 U20468 ( .A1(n9811), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17215) );
  OAI21_X1 U20469 ( .B1(n9856), .B2(n17216), .A(n17215), .ZN(n17228) );
  INV_X1 U20470 ( .A(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17226) );
  AOI22_X1 U20471 ( .A1(n11474), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17273), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17225) );
  AOI22_X1 U20472 ( .A1(n17310), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17217) );
  OAI21_X1 U20473 ( .B1(n17312), .B2(n17218), .A(n17217), .ZN(n17224) );
  AOI22_X1 U20474 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17221) );
  AOI22_X1 U20475 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17220) );
  OAI211_X1 U20476 ( .C1(n11448), .C2(n17222), .A(n17221), .B(n17220), .ZN(
        n17223) );
  OAI211_X1 U20477 ( .C1(n11523), .C2(n17226), .A(n17225), .B(n9994), .ZN(
        n17227) );
  AOI211_X1 U20478 ( .C1(n17245), .C2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A(
        n17228), .B(n17227), .ZN(n17452) );
  OAI21_X1 U20479 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n9951), .A(n17229), .ZN(
        n17230) );
  AOI22_X1 U20480 ( .A1(n17361), .A2(n17452), .B1(n17230), .B2(n17358), .ZN(
        P3_U2688) );
  AOI22_X1 U20481 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17231) );
  OAI21_X1 U20482 ( .B1(n11498), .B2(n17232), .A(n17231), .ZN(n17244) );
  AOI22_X1 U20483 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17241) );
  AOI22_X1 U20484 ( .A1(n17310), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17233) );
  OAI21_X1 U20485 ( .B1(n11448), .B2(n17343), .A(n17233), .ZN(n17239) );
  AOI22_X1 U20486 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17235) );
  AOI22_X1 U20487 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17234) );
  OAI211_X1 U20488 ( .C1(n17237), .C2(n17236), .A(n17235), .B(n17234), .ZN(
        n17238) );
  AOI211_X1 U20489 ( .C1(n17292), .C2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A(
        n17239), .B(n17238), .ZN(n17240) );
  OAI211_X1 U20490 ( .C1(n9856), .C2(n17242), .A(n17241), .B(n17240), .ZN(
        n17243) );
  AOI211_X1 U20491 ( .C1(n17245), .C2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n17244), .B(n17243), .ZN(n17464) );
  OAI21_X1 U20492 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17247), .A(n17246), .ZN(
        n17248) );
  OAI21_X1 U20493 ( .B1(n17464), .B2(n17358), .A(n17248), .ZN(P3_U2691) );
  NAND2_X1 U20494 ( .A1(n17250), .A2(n17249), .ZN(n17265) );
  AOI22_X1 U20495 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17292), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17263) );
  AOI22_X1 U20496 ( .A1(n17273), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17251) );
  OAI21_X1 U20497 ( .B1(n11523), .B2(n17252), .A(n17251), .ZN(n17261) );
  OAI22_X1 U20498 ( .A1(n17288), .A2(n17254), .B1(n17197), .B2(n17253), .ZN(
        n17255) );
  AOI21_X1 U20499 ( .B1(n17309), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n17255), .ZN(n17259) );
  AOI22_X1 U20500 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17258) );
  AOI22_X1 U20501 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17257) );
  NAND4_X1 U20502 ( .A1(n17259), .A2(n17258), .A3(n17257), .A4(n17256), .ZN(
        n17260) );
  AOI211_X1 U20503 ( .C1(n9812), .C2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n17261), .B(n17260), .ZN(n17262) );
  OAI211_X1 U20504 ( .C1(n11448), .C2(n17347), .A(n17263), .B(n17262), .ZN(
        n17468) );
  OAI221_X1 U20505 ( .B1(n17361), .B2(n17265), .C1(n17358), .C2(n17468), .A(
        n17264), .ZN(n17266) );
  INV_X1 U20506 ( .A(n17266), .ZN(P3_U2692) );
  NAND2_X1 U20507 ( .A1(n18366), .A2(n17267), .ZN(n17283) );
  NOR2_X1 U20508 ( .A1(n17361), .A2(n17267), .ZN(n17305) );
  AOI22_X1 U20509 ( .A1(n17310), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17268), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17281) );
  AOI22_X1 U20510 ( .A1(n9812), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17271) );
  AOI22_X1 U20511 ( .A1(n9811), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17270) );
  OAI211_X1 U20512 ( .C1(n17312), .C2(n17272), .A(n17271), .B(n17270), .ZN(
        n17280) );
  AOI22_X1 U20513 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17273), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17278) );
  AOI22_X1 U20514 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17309), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17277) );
  AOI22_X1 U20515 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17291), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17276) );
  NAND2_X1 U20516 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n17275) );
  NAND4_X1 U20517 ( .A1(n17278), .A2(n17277), .A3(n17276), .A4(n17275), .ZN(
        n17279) );
  OAI211_X1 U20518 ( .C1(n11448), .C2(n17354), .A(n17281), .B(n9995), .ZN(
        n17471) );
  AOI22_X1 U20519 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17305), .B1(n17361), 
        .B2(n17471), .ZN(n17282) );
  OAI21_X1 U20520 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17283), .A(n17282), .ZN(
        P3_U2693) );
  AOI22_X1 U20521 ( .A1(n9811), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17286) );
  OAI21_X1 U20522 ( .B1(n17288), .B2(n17287), .A(n17286), .ZN(n17303) );
  INV_X1 U20523 ( .A(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17301) );
  AOI22_X1 U20524 ( .A1(n17309), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17300) );
  OAI22_X1 U20525 ( .A1(n17197), .A2(n17290), .B1(n11467), .B2(n17289), .ZN(
        n17298) );
  AOI22_X1 U20526 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17291), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17296) );
  AOI22_X1 U20527 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17211), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17295) );
  AOI22_X1 U20528 ( .A1(n17293), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17292), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17294) );
  NAND3_X1 U20529 ( .A1(n17296), .A2(n17295), .A3(n17294), .ZN(n17297) );
  OAI211_X1 U20530 ( .C1(n11447), .C2(n17301), .A(n17300), .B(n17299), .ZN(
        n17302) );
  AOI211_X1 U20531 ( .C1(n17304), .C2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A(
        n17303), .B(n17302), .ZN(n17475) );
  OAI21_X1 U20532 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17306), .A(n17305), .ZN(
        n17307) );
  OAI21_X1 U20533 ( .B1(n17475), .B2(n17358), .A(n17307), .ZN(P3_U2694) );
  INV_X1 U20534 ( .A(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18491) );
  AOI22_X1 U20535 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__0__SCAN_IN), .B2(n17284), .ZN(n17308) );
  OAI21_X1 U20536 ( .B1(n9888), .B2(n18491), .A(n17308), .ZN(n17324) );
  AOI22_X1 U20537 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n17309), .B1(
        P3_INSTQUEUE_REG_14__0__SCAN_IN), .B2(n17211), .ZN(n17321) );
  OAI21_X1 U20538 ( .B1(n17312), .B2(n18373), .A(n17311), .ZN(n17319) );
  AOI22_X1 U20539 ( .A1(n17313), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17304), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17316) );
  AOI22_X1 U20540 ( .A1(n17314), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17315) );
  OAI211_X1 U20541 ( .C1(n17317), .C2(n11448), .A(n17316), .B(n17315), .ZN(
        n17318) );
  AOI211_X1 U20542 ( .C1(n17268), .C2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n17319), .B(n17318), .ZN(n17320) );
  OAI211_X1 U20543 ( .C1(n17322), .C2(n11447), .A(n17321), .B(n17320), .ZN(
        n17323) );
  AOI211_X1 U20544 ( .C1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .C2(n17325), .A(
        n17324), .B(n17323), .ZN(n17480) );
  NOR2_X1 U20545 ( .A1(n17409), .A2(n17328), .ZN(n17329) );
  OAI221_X1 U20546 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(P3_EBX_REG_7__SCAN_IN), 
        .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17329), .A(n17326), .ZN(n17327) );
  AOI22_X1 U20547 ( .A1(n17361), .A2(n17480), .B1(n17327), .B2(n17358), .ZN(
        P3_U2695) );
  NAND2_X1 U20548 ( .A1(n17358), .A2(n17328), .ZN(n17334) );
  AOI22_X1 U20549 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n17361), .B1(
        n17329), .B2(n17331), .ZN(n17330) );
  OAI21_X1 U20550 ( .B1(n17331), .B2(n17334), .A(n17330), .ZN(P3_U2696) );
  AND2_X1 U20551 ( .A1(n17332), .A2(n17336), .ZN(n17335) );
  OAI22_X1 U20552 ( .A1(n17335), .A2(n17334), .B1(n17333), .B2(n17358), .ZN(
        P3_U2697) );
  OAI21_X1 U20553 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17337), .A(n17336), .ZN(
        n17338) );
  AOI22_X1 U20554 ( .A1(n17361), .A2(n17339), .B1(n17338), .B2(n17358), .ZN(
        P3_U2698) );
  NOR2_X1 U20555 ( .A1(n17409), .A2(n17360), .ZN(n17355) );
  NAND2_X1 U20556 ( .A1(n17340), .A2(n17355), .ZN(n17346) );
  NOR2_X1 U20557 ( .A1(n17341), .A2(n17346), .ZN(n17349) );
  AOI21_X1 U20558 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17358), .A(n17349), .ZN(
        n17345) );
  INV_X1 U20559 ( .A(n17355), .ZN(n17363) );
  NOR2_X1 U20560 ( .A1(n17342), .A2(n17363), .ZN(n17344) );
  OAI22_X1 U20561 ( .A1(n17345), .A2(n17344), .B1(n17343), .B2(n17358), .ZN(
        P3_U2699) );
  INV_X1 U20562 ( .A(n17346), .ZN(n17352) );
  AOI21_X1 U20563 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17358), .A(n17352), .ZN(
        n17348) );
  OAI22_X1 U20564 ( .A1(n17349), .A2(n17348), .B1(n17347), .B2(n17358), .ZN(
        P3_U2700) );
  AOI21_X1 U20565 ( .B1(n18366), .B2(n17350), .A(n17360), .ZN(n17351) );
  NOR2_X1 U20566 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n17351), .ZN(n17353) );
  AOI211_X1 U20567 ( .C1(n17361), .C2(n17354), .A(n17353), .B(n17352), .ZN(
        P3_U2701) );
  AOI22_X1 U20568 ( .A1(P3_EBX_REG_1__SCAN_IN), .A2(n17360), .B1(n17356), .B2(
        n17355), .ZN(n17357) );
  OAI21_X1 U20569 ( .B1(n17359), .B2(n17358), .A(n17357), .ZN(P3_U2702) );
  AOI22_X1 U20570 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17361), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17360), .ZN(n17362) );
  OAI21_X1 U20571 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17363), .A(n17362), .ZN(
        P3_U2703) );
  INV_X1 U20572 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17581) );
  INV_X1 U20573 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17576) );
  INV_X1 U20574 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17568) );
  INV_X1 U20575 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17558) );
  INV_X1 U20576 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17620) );
  NAND4_X1 U20577 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(P3_EAX_REG_9__SCAN_IN), .ZN(n17366)
         );
  NAND4_X1 U20578 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(P3_EAX_REG_7__SCAN_IN), 
        .A3(P3_EAX_REG_6__SCAN_IN), .A4(P3_EAX_REG_3__SCAN_IN), .ZN(n17365) );
  NAND2_X1 U20579 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .ZN(n17453) );
  INV_X1 U20580 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17589) );
  NOR2_X1 U20581 ( .A1(n17589), .A2(n17587), .ZN(n17502) );
  NAND4_X1 U20582 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17502), .A3(
        P3_EAX_REG_14__SCAN_IN), .A4(P3_EAX_REG_13__SCAN_IN), .ZN(n17364) );
  NOR4_X1 U20583 ( .A1(n17366), .A2(n17365), .A3(n17453), .A4(n17364), .ZN(
        n17367) );
  NAND2_X1 U20584 ( .A1(n17514), .A2(n17367), .ZN(n17455) );
  NAND4_X1 U20585 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .A3(P3_EAX_REG_20__SCAN_IN), .A4(P3_EAX_REG_19__SCAN_IN), .ZN(n17410)
         );
  NAND2_X1 U20586 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17405), .ZN(n17404) );
  NAND2_X1 U20587 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17400), .ZN(n17399) );
  NAND2_X1 U20588 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17389), .ZN(n17385) );
  NAND2_X1 U20589 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17381), .ZN(n17376) );
  NAND2_X1 U20590 ( .A1(n17372), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17371) );
  NOR2_X2 U20591 ( .A1(n18360), .A2(n17494), .ZN(n17442) );
  OAI22_X1 U20592 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17501), .B1(n17449), 
        .B2(n17372), .ZN(n17368) );
  AOI22_X1 U20593 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17442), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17368), .ZN(n17369) );
  OAI21_X1 U20594 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17371), .A(n17369), .ZN(
        P3_U2704) );
  NOR2_X2 U20595 ( .A1(n17370), .A2(n17494), .ZN(n17443) );
  AOI22_X1 U20596 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17443), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17442), .ZN(n17374) );
  OAI211_X1 U20597 ( .C1(n17372), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17494), .B(
        n17371), .ZN(n17373) );
  OAI211_X1 U20598 ( .C1(n17375), .C2(n17504), .A(n17374), .B(n17373), .ZN(
        P3_U2705) );
  AOI22_X1 U20599 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17443), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17442), .ZN(n17378) );
  OAI211_X1 U20600 ( .C1(n17381), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17494), .B(
        n17376), .ZN(n17377) );
  OAI211_X1 U20601 ( .C1(n17504), .C2(n17379), .A(n17378), .B(n17377), .ZN(
        P3_U2706) );
  INV_X1 U20602 ( .A(n17442), .ZN(n17441) );
  AOI22_X1 U20603 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17443), .B1(n17380), .B2(
        n17508), .ZN(n17384) );
  AOI211_X1 U20604 ( .C1(n17581), .C2(n17385), .A(n17381), .B(n17449), .ZN(
        n17382) );
  INV_X1 U20605 ( .A(n17382), .ZN(n17383) );
  OAI211_X1 U20606 ( .C1(n17441), .C2(n19463), .A(n17384), .B(n17383), .ZN(
        P3_U2707) );
  AOI22_X1 U20607 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17443), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17442), .ZN(n17387) );
  OAI211_X1 U20608 ( .C1(n17389), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17494), .B(
        n17385), .ZN(n17386) );
  OAI211_X1 U20609 ( .C1(n17504), .C2(n17388), .A(n17387), .B(n17386), .ZN(
        P3_U2708) );
  AOI22_X1 U20610 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17443), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17442), .ZN(n17392) );
  AOI211_X1 U20611 ( .C1(n17576), .C2(n17394), .A(n17389), .B(n17449), .ZN(
        n17390) );
  INV_X1 U20612 ( .A(n17390), .ZN(n17391) );
  OAI211_X1 U20613 ( .C1(n17504), .C2(n17393), .A(n17392), .B(n17391), .ZN(
        P3_U2709) );
  AOI22_X1 U20614 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17443), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17442), .ZN(n17397) );
  OAI211_X1 U20615 ( .C1(n17395), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17494), .B(
        n17394), .ZN(n17396) );
  OAI211_X1 U20616 ( .C1(n17504), .C2(n17398), .A(n17397), .B(n17396), .ZN(
        P3_U2710) );
  AOI22_X1 U20617 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17443), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17442), .ZN(n17402) );
  OAI211_X1 U20618 ( .C1(n17400), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17494), .B(
        n17399), .ZN(n17401) );
  OAI211_X1 U20619 ( .C1(n17504), .C2(n17403), .A(n17402), .B(n17401), .ZN(
        P3_U2711) );
  AOI22_X1 U20620 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17443), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17442), .ZN(n17407) );
  OAI211_X1 U20621 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17405), .A(n17494), .B(
        n17404), .ZN(n17406) );
  OAI211_X1 U20622 ( .C1(n17504), .C2(n17408), .A(n17407), .B(n17406), .ZN(
        P3_U2712) );
  INV_X1 U20623 ( .A(n17443), .ZN(n17416) );
  NOR2_X1 U20624 ( .A1(n17409), .A2(n17444), .ZN(n17438) );
  NAND2_X1 U20625 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n17438), .ZN(n17437) );
  NOR2_X1 U20626 ( .A1(n17410), .A2(n17437), .ZN(n17414) );
  INV_X1 U20627 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17560) );
  NAND3_X1 U20628 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(n17431), .ZN(n17422) );
  NAND2_X1 U20629 ( .A1(n17494), .A2(n17422), .ZN(n17426) );
  OAI21_X1 U20630 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17501), .A(n17426), .ZN(
        n17413) );
  OAI22_X1 U20631 ( .A1(n17411), .A2(n17504), .B1(n18359), .B2(n17441), .ZN(
        n17412) );
  AOI221_X1 U20632 ( .B1(n17414), .B2(n17568), .C1(n17413), .C2(
        P3_EAX_REG_22__SCAN_IN), .A(n17412), .ZN(n17415) );
  OAI21_X1 U20633 ( .B1(n18358), .B2(n17416), .A(n17415), .ZN(P3_U2713) );
  INV_X1 U20634 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17566) );
  OAI22_X1 U20635 ( .A1(n17417), .A2(n17504), .B1(n15083), .B2(n17441), .ZN(
        n17418) );
  AOI21_X1 U20636 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17443), .A(n17418), .ZN(
        n17419) );
  OAI221_X1 U20637 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17422), .C1(n17566), 
        .C2(n17426), .A(n17419), .ZN(P3_U2714) );
  INV_X1 U20638 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17564) );
  INV_X1 U20639 ( .A(n17420), .ZN(n17421) );
  AOI22_X1 U20640 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17443), .B1(n17508), .B2(
        n17421), .ZN(n17425) );
  NAND2_X1 U20641 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17431), .ZN(n17427) );
  INV_X1 U20642 ( .A(n17427), .ZN(n17423) );
  AOI22_X1 U20643 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n17442), .B1(n17423), .B2(
        n17422), .ZN(n17424) );
  OAI211_X1 U20644 ( .C1(n17564), .C2(n17426), .A(n17425), .B(n17424), .ZN(
        P3_U2715) );
  AOI22_X1 U20645 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17443), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17442), .ZN(n17429) );
  OAI211_X1 U20646 ( .C1(n17431), .C2(P3_EAX_REG_19__SCAN_IN), .A(n17494), .B(
        n17427), .ZN(n17428) );
  OAI211_X1 U20647 ( .C1(n17430), .C2(n17504), .A(n17429), .B(n17428), .ZN(
        P3_U2716) );
  AOI22_X1 U20648 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17443), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17442), .ZN(n17434) );
  AOI211_X1 U20649 ( .C1(n17560), .C2(n17437), .A(n17431), .B(n17449), .ZN(
        n17432) );
  INV_X1 U20650 ( .A(n17432), .ZN(n17433) );
  OAI211_X1 U20651 ( .C1(n17435), .C2(n17504), .A(n17434), .B(n17433), .ZN(
        P3_U2717) );
  AOI22_X1 U20652 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17443), .B1(n17508), .B2(
        n17436), .ZN(n17440) );
  OAI211_X1 U20653 ( .C1(n17438), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17494), .B(
        n17437), .ZN(n17439) );
  OAI211_X1 U20654 ( .C1(n17441), .C2(n19449), .A(n17440), .B(n17439), .ZN(
        P3_U2718) );
  AOI22_X1 U20655 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17443), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17442), .ZN(n17446) );
  OAI211_X1 U20656 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17448), .A(n17494), .B(
        n17444), .ZN(n17445) );
  OAI211_X1 U20657 ( .C1(n17447), .C2(n17504), .A(n17446), .B(n17445), .ZN(
        P3_U2719) );
  AOI211_X1 U20658 ( .C1(n17620), .C2(n17455), .A(n17449), .B(n17448), .ZN(
        n17450) );
  AOI21_X1 U20659 ( .B1(n17509), .B2(BUF2_REG_15__SCAN_IN), .A(n17450), .ZN(
        n17451) );
  OAI21_X1 U20660 ( .B1(n17452), .B2(n17504), .A(n17451), .ZN(P3_U2720) );
  INV_X1 U20661 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17610) );
  INV_X1 U20662 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17603) );
  INV_X1 U20663 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17591) );
  INV_X1 U20664 ( .A(n17502), .ZN(n17510) );
  NAND2_X1 U20665 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17506), .ZN(n17493) );
  NAND2_X1 U20666 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17489), .ZN(n17479) );
  NAND2_X1 U20667 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17482), .ZN(n17473) );
  NAND2_X1 U20668 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17477), .ZN(n17470) );
  NOR2_X1 U20669 ( .A1(n17610), .A2(n17470), .ZN(n17463) );
  NAND2_X1 U20670 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17466), .ZN(n17458) );
  AOI22_X1 U20671 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17509), .B1(n17508), .B2(
        n17454), .ZN(n17457) );
  NAND3_X1 U20672 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17494), .A3(n17455), 
        .ZN(n17456) );
  OAI211_X1 U20673 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n17458), .A(n17457), .B(
        n17456), .ZN(P3_U2721) );
  INV_X1 U20674 ( .A(n17458), .ZN(n17461) );
  AOI21_X1 U20675 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17494), .A(n17466), .ZN(
        n17460) );
  OAI222_X1 U20676 ( .A1(n17507), .A2(n17462), .B1(n17461), .B2(n17460), .C1(
        n17504), .C2(n17459), .ZN(P3_U2722) );
  AOI21_X1 U20677 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17494), .A(n17463), .ZN(
        n17465) );
  OAI222_X1 U20678 ( .A1(n17507), .A2(n17467), .B1(n17466), .B2(n17465), .C1(
        n17504), .C2(n17464), .ZN(P3_U2723) );
  NAND2_X1 U20679 ( .A1(n17494), .A2(n17470), .ZN(n17474) );
  AOI22_X1 U20680 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17509), .B1(n17508), .B2(
        n17468), .ZN(n17469) );
  OAI221_X1 U20681 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17470), .C1(n17610), 
        .C2(n17474), .A(n17469), .ZN(P3_U2724) );
  INV_X1 U20682 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17608) );
  AOI22_X1 U20683 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17509), .B1(n17508), .B2(
        n17471), .ZN(n17472) );
  OAI221_X1 U20684 ( .B1(n17474), .B2(n17608), .C1(n17474), .C2(n17473), .A(
        n17472), .ZN(P3_U2725) );
  AOI21_X1 U20685 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17494), .A(n17482), .ZN(
        n17476) );
  OAI222_X1 U20686 ( .A1(n17507), .A2(n17478), .B1(n17477), .B2(n17476), .C1(
        n17504), .C2(n17475), .ZN(P3_U2726) );
  INV_X1 U20687 ( .A(n17479), .ZN(n17486) );
  AOI21_X1 U20688 ( .B1(P3_EAX_REG_8__SCAN_IN), .B2(n17494), .A(n17486), .ZN(
        n17481) );
  OAI222_X1 U20689 ( .A1(n17507), .A2(n17483), .B1(n17482), .B2(n17481), .C1(
        n17504), .C2(n17480), .ZN(P3_U2727) );
  AOI21_X1 U20690 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17494), .A(n17489), .ZN(
        n17485) );
  OAI222_X1 U20691 ( .A1(n17507), .A2(n18363), .B1(n17486), .B2(n17485), .C1(
        n17504), .C2(n17484), .ZN(P3_U2728) );
  AOI21_X1 U20692 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17494), .A(n17492), .ZN(
        n17488) );
  OAI222_X1 U20693 ( .A1(n18358), .A2(n17507), .B1(n17489), .B2(n17488), .C1(
        n17504), .C2(n17487), .ZN(P3_U2729) );
  INV_X1 U20694 ( .A(n17493), .ZN(n17500) );
  AOI22_X1 U20695 ( .A1(n17500), .A2(P3_EAX_REG_4__SCAN_IN), .B1(
        P3_EAX_REG_5__SCAN_IN), .B2(n17494), .ZN(n17491) );
  OAI222_X1 U20696 ( .A1(n18354), .A2(n17507), .B1(n17492), .B2(n17491), .C1(
        n17504), .C2(n17490), .ZN(P3_U2730) );
  INV_X1 U20697 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17595) );
  NOR2_X1 U20698 ( .A1(n17595), .A2(n17493), .ZN(n17497) );
  AOI21_X1 U20699 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17494), .A(n17500), .ZN(
        n17496) );
  OAI222_X1 U20700 ( .A1(n18350), .A2(n17507), .B1(n17497), .B2(n17496), .C1(
        n17504), .C2(n17495), .ZN(P3_U2731) );
  AOI21_X1 U20701 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17494), .A(n17506), .ZN(
        n17499) );
  OAI222_X1 U20702 ( .A1(n18346), .A2(n17507), .B1(n17500), .B2(n17499), .C1(
        n17504), .C2(n17498), .ZN(P3_U2732) );
  INV_X1 U20703 ( .A(n17501), .ZN(n17511) );
  AOI22_X1 U20704 ( .A1(n17511), .A2(n17502), .B1(P3_EAX_REG_2__SCAN_IN), .B2(
        n17494), .ZN(n17505) );
  OAI222_X1 U20705 ( .A1(n18342), .A2(n17507), .B1(n17506), .B2(n17505), .C1(
        n17504), .C2(n17503), .ZN(P3_U2733) );
  AOI22_X1 U20706 ( .A1(n17509), .A2(BUF2_REG_1__SCAN_IN), .B1(n17508), .B2(
        n11533), .ZN(n17513) );
  OAI211_X1 U20707 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(P3_EAX_REG_0__SCAN_IN), 
        .A(n17511), .B(n17510), .ZN(n17512) );
  OAI211_X1 U20708 ( .C1(n17514), .C2(n17589), .A(n17513), .B(n17512), .ZN(
        P3_U2734) );
  NAND2_X1 U20709 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17824), .ZN(n18773) );
  INV_X2 U20710 ( .A(n18773), .ZN(n17550) );
  NOR2_X4 U20711 ( .A1(n17550), .A2(n17517), .ZN(n17530) );
  AND2_X1 U20712 ( .A1(n17530), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20713 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17585) );
  AOI22_X1 U20714 ( .A1(n17550), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(n17530), .ZN(n17518) );
  OAI21_X1 U20715 ( .B1(n17585), .B2(n17534), .A(n17518), .ZN(P3_U2737) );
  INV_X1 U20716 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17583) );
  AOI22_X1 U20717 ( .A1(n17550), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17530), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17519) );
  OAI21_X1 U20718 ( .B1(n17583), .B2(n17534), .A(n17519), .ZN(P3_U2738) );
  AOI22_X1 U20719 ( .A1(n17550), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17530), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17520) );
  OAI21_X1 U20720 ( .B1(n17581), .B2(n17534), .A(n17520), .ZN(P3_U2739) );
  INV_X1 U20721 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17579) );
  AOI22_X1 U20722 ( .A1(n17550), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17530), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17521) );
  OAI21_X1 U20723 ( .B1(n17579), .B2(n17534), .A(n17521), .ZN(P3_U2740) );
  AOI22_X1 U20724 ( .A1(n17550), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17530), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17522) );
  OAI21_X1 U20725 ( .B1(n17576), .B2(n17534), .A(n17522), .ZN(P3_U2741) );
  INV_X1 U20726 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17574) );
  AOI22_X1 U20727 ( .A1(n17550), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17530), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17523) );
  OAI21_X1 U20728 ( .B1(n17574), .B2(n17534), .A(n17523), .ZN(P3_U2742) );
  INV_X1 U20729 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17572) );
  AOI22_X1 U20730 ( .A1(n17550), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17530), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17524) );
  OAI21_X1 U20731 ( .B1(n17572), .B2(n17534), .A(n17524), .ZN(P3_U2743) );
  INV_X1 U20732 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17570) );
  AOI22_X1 U20733 ( .A1(n17550), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17530), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17525) );
  OAI21_X1 U20734 ( .B1(n17570), .B2(n17534), .A(n17525), .ZN(P3_U2744) );
  AOI22_X1 U20735 ( .A1(n17550), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17530), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17526) );
  OAI21_X1 U20736 ( .B1(n17568), .B2(n17534), .A(n17526), .ZN(P3_U2745) );
  AOI22_X1 U20737 ( .A1(n17550), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17530), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17527) );
  OAI21_X1 U20738 ( .B1(n17566), .B2(n17534), .A(n17527), .ZN(P3_U2746) );
  AOI22_X1 U20739 ( .A1(n17550), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17530), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17528) );
  OAI21_X1 U20740 ( .B1(n17564), .B2(n17534), .A(n17528), .ZN(P3_U2747) );
  INV_X1 U20741 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17562) );
  AOI22_X1 U20742 ( .A1(n17550), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17530), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17529) );
  OAI21_X1 U20743 ( .B1(n17562), .B2(n17534), .A(n17529), .ZN(P3_U2748) );
  AOI22_X1 U20744 ( .A1(n17550), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17530), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17531) );
  OAI21_X1 U20745 ( .B1(n17560), .B2(n17534), .A(n17531), .ZN(P3_U2749) );
  AOI22_X1 U20746 ( .A1(n17550), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17530), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17532) );
  OAI21_X1 U20747 ( .B1(n17558), .B2(n17534), .A(n17532), .ZN(P3_U2750) );
  INV_X1 U20748 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17556) );
  AOI22_X1 U20749 ( .A1(n17550), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17530), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17533) );
  OAI21_X1 U20750 ( .B1(n17556), .B2(n17534), .A(n17533), .ZN(P3_U2751) );
  AOI22_X1 U20751 ( .A1(n17550), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17530), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17535) );
  OAI21_X1 U20752 ( .B1(n17620), .B2(n17552), .A(n17535), .ZN(P3_U2752) );
  INV_X1 U20753 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17616) );
  AOI22_X1 U20754 ( .A1(n17550), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17530), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17536) );
  OAI21_X1 U20755 ( .B1(n17616), .B2(n17552), .A(n17536), .ZN(P3_U2753) );
  INV_X1 U20756 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17614) );
  AOI22_X1 U20757 ( .A1(n17550), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17530), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17537) );
  OAI21_X1 U20758 ( .B1(n17614), .B2(n17552), .A(n17537), .ZN(P3_U2754) );
  INV_X1 U20759 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17612) );
  AOI22_X1 U20760 ( .A1(n17550), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17530), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17538) );
  OAI21_X1 U20761 ( .B1(n17612), .B2(n17552), .A(n17538), .ZN(P3_U2755) );
  AOI22_X1 U20762 ( .A1(n17550), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17530), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17539) );
  OAI21_X1 U20763 ( .B1(n17610), .B2(n17552), .A(n17539), .ZN(P3_U2756) );
  AOI22_X1 U20764 ( .A1(n17550), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17530), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17540) );
  OAI21_X1 U20765 ( .B1(n17608), .B2(n17552), .A(n17540), .ZN(P3_U2757) );
  INV_X1 U20766 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17606) );
  AOI22_X1 U20767 ( .A1(n17550), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17530), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17541) );
  OAI21_X1 U20768 ( .B1(n17606), .B2(n17552), .A(n17541), .ZN(P3_U2758) );
  AOI22_X1 U20769 ( .A1(n17550), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17530), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17542) );
  OAI21_X1 U20770 ( .B1(n17603), .B2(n17552), .A(n17542), .ZN(P3_U2759) );
  INV_X1 U20771 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17601) );
  AOI22_X1 U20772 ( .A1(n17550), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17530), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17543) );
  OAI21_X1 U20773 ( .B1(n17601), .B2(n17552), .A(n17543), .ZN(P3_U2760) );
  INV_X1 U20774 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17599) );
  AOI22_X1 U20775 ( .A1(n17550), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17530), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17544) );
  OAI21_X1 U20776 ( .B1(n17599), .B2(n17552), .A(n17544), .ZN(P3_U2761) );
  INV_X1 U20777 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17597) );
  AOI22_X1 U20778 ( .A1(n17550), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17530), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17545) );
  OAI21_X1 U20779 ( .B1(n17597), .B2(n17552), .A(n17545), .ZN(P3_U2762) );
  AOI22_X1 U20780 ( .A1(n17550), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17530), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17546) );
  OAI21_X1 U20781 ( .B1(n17595), .B2(n17552), .A(n17546), .ZN(P3_U2763) );
  INV_X1 U20782 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17593) );
  AOI22_X1 U20783 ( .A1(n17550), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17530), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17547) );
  OAI21_X1 U20784 ( .B1(n17593), .B2(n17552), .A(n17547), .ZN(P3_U2764) );
  AOI22_X1 U20785 ( .A1(n17550), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17530), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17548) );
  OAI21_X1 U20786 ( .B1(n17591), .B2(n17552), .A(n17548), .ZN(P3_U2765) );
  AOI22_X1 U20787 ( .A1(n17550), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17530), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17549) );
  OAI21_X1 U20788 ( .B1(n17589), .B2(n17552), .A(n17549), .ZN(P3_U2766) );
  AOI22_X1 U20789 ( .A1(n17550), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17530), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17551) );
  OAI21_X1 U20790 ( .B1(n17587), .B2(n17552), .A(n17551), .ZN(P3_U2767) );
  NOR2_X4 U20791 ( .A1(n18339), .A2(n17604), .ZN(n17577) );
  AOI22_X1 U20792 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17577), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17604), .ZN(n17555) );
  OAI21_X1 U20793 ( .B1(n17556), .B2(n17619), .A(n17555), .ZN(P3_U2768) );
  AOI22_X1 U20794 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17577), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17604), .ZN(n17557) );
  OAI21_X1 U20795 ( .B1(n17558), .B2(n17619), .A(n17557), .ZN(P3_U2769) );
  AOI22_X1 U20796 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17577), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17604), .ZN(n17559) );
  OAI21_X1 U20797 ( .B1(n17560), .B2(n17619), .A(n17559), .ZN(P3_U2770) );
  AOI22_X1 U20798 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17577), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17604), .ZN(n17561) );
  OAI21_X1 U20799 ( .B1(n17562), .B2(n17619), .A(n17561), .ZN(P3_U2771) );
  AOI22_X1 U20800 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17577), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17604), .ZN(n17563) );
  OAI21_X1 U20801 ( .B1(n17564), .B2(n17619), .A(n17563), .ZN(P3_U2772) );
  AOI22_X1 U20802 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17577), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17604), .ZN(n17565) );
  OAI21_X1 U20803 ( .B1(n17566), .B2(n17619), .A(n17565), .ZN(P3_U2773) );
  AOI22_X1 U20804 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17577), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17604), .ZN(n17567) );
  OAI21_X1 U20805 ( .B1(n17568), .B2(n17619), .A(n17567), .ZN(P3_U2774) );
  AOI22_X1 U20806 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17577), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17604), .ZN(n17569) );
  OAI21_X1 U20807 ( .B1(n17570), .B2(n17619), .A(n17569), .ZN(P3_U2775) );
  AOI22_X1 U20808 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17577), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17604), .ZN(n17571) );
  OAI21_X1 U20809 ( .B1(n17572), .B2(n17619), .A(n17571), .ZN(P3_U2776) );
  AOI22_X1 U20810 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17577), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17604), .ZN(n17573) );
  OAI21_X1 U20811 ( .B1(n17574), .B2(n17619), .A(n17573), .ZN(P3_U2777) );
  AOI22_X1 U20812 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17577), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17604), .ZN(n17575) );
  OAI21_X1 U20813 ( .B1(n17576), .B2(n17619), .A(n17575), .ZN(P3_U2778) );
  AOI22_X1 U20814 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17577), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17604), .ZN(n17578) );
  OAI21_X1 U20815 ( .B1(n17579), .B2(n17619), .A(n17578), .ZN(P3_U2779) );
  AOI22_X1 U20816 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17577), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17604), .ZN(n17580) );
  OAI21_X1 U20817 ( .B1(n17581), .B2(n17619), .A(n17580), .ZN(P3_U2780) );
  AOI22_X1 U20818 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17577), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17604), .ZN(n17582) );
  OAI21_X1 U20819 ( .B1(n17583), .B2(n17619), .A(n17582), .ZN(P3_U2781) );
  AOI22_X1 U20820 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17577), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17604), .ZN(n17584) );
  OAI21_X1 U20821 ( .B1(n17585), .B2(n17619), .A(n17584), .ZN(P3_U2782) );
  AOI22_X1 U20822 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17577), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17604), .ZN(n17586) );
  OAI21_X1 U20823 ( .B1(n17587), .B2(n17619), .A(n17586), .ZN(P3_U2783) );
  AOI22_X1 U20824 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17577), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17604), .ZN(n17588) );
  OAI21_X1 U20825 ( .B1(n17589), .B2(n17619), .A(n17588), .ZN(P3_U2784) );
  AOI22_X1 U20826 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17577), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17604), .ZN(n17590) );
  OAI21_X1 U20827 ( .B1(n17591), .B2(n17619), .A(n17590), .ZN(P3_U2785) );
  AOI22_X1 U20828 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17577), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17604), .ZN(n17592) );
  OAI21_X1 U20829 ( .B1(n17593), .B2(n17619), .A(n17592), .ZN(P3_U2786) );
  AOI22_X1 U20830 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17577), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17604), .ZN(n17594) );
  OAI21_X1 U20831 ( .B1(n17595), .B2(n17619), .A(n17594), .ZN(P3_U2787) );
  AOI22_X1 U20832 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17577), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17617), .ZN(n17596) );
  OAI21_X1 U20833 ( .B1(n17597), .B2(n17619), .A(n17596), .ZN(P3_U2788) );
  AOI22_X1 U20834 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17577), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17617), .ZN(n17598) );
  OAI21_X1 U20835 ( .B1(n17599), .B2(n17619), .A(n17598), .ZN(P3_U2789) );
  AOI22_X1 U20836 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17577), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17617), .ZN(n17600) );
  OAI21_X1 U20837 ( .B1(n17601), .B2(n17619), .A(n17600), .ZN(P3_U2790) );
  AOI22_X1 U20838 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17577), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17617), .ZN(n17602) );
  OAI21_X1 U20839 ( .B1(n17603), .B2(n17619), .A(n17602), .ZN(P3_U2791) );
  AOI22_X1 U20840 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17577), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17604), .ZN(n17605) );
  OAI21_X1 U20841 ( .B1(n17606), .B2(n17619), .A(n17605), .ZN(P3_U2792) );
  AOI22_X1 U20842 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17577), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17617), .ZN(n17607) );
  OAI21_X1 U20843 ( .B1(n17608), .B2(n17619), .A(n17607), .ZN(P3_U2793) );
  AOI22_X1 U20844 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17577), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17617), .ZN(n17609) );
  OAI21_X1 U20845 ( .B1(n17610), .B2(n17619), .A(n17609), .ZN(P3_U2794) );
  AOI22_X1 U20846 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17577), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17617), .ZN(n17611) );
  OAI21_X1 U20847 ( .B1(n17612), .B2(n17619), .A(n17611), .ZN(P3_U2795) );
  AOI22_X1 U20848 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17577), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17617), .ZN(n17613) );
  OAI21_X1 U20849 ( .B1(n17614), .B2(n17619), .A(n17613), .ZN(P3_U2796) );
  AOI22_X1 U20850 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17577), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17617), .ZN(n17615) );
  OAI21_X1 U20851 ( .B1(n17616), .B2(n17619), .A(n17615), .ZN(P3_U2797) );
  AOI22_X1 U20852 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17577), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17617), .ZN(n17618) );
  OAI21_X1 U20853 ( .B1(n17620), .B2(n17619), .A(n17618), .ZN(P3_U2798) );
  OAI21_X1 U20854 ( .B1(n17621), .B2(n17989), .A(n17988), .ZN(n17622) );
  AOI21_X1 U20855 ( .B1(n18845), .B2(n17626), .A(n17622), .ZN(n17652) );
  OAI21_X1 U20856 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17703), .A(
        n17652), .ZN(n17639) );
  AOI211_X1 U20857 ( .C1(n17625), .C2(n17624), .A(n17623), .B(n17898), .ZN(
        n17632) );
  NOR2_X1 U20858 ( .A1(n17834), .A2(n17626), .ZN(n17644) );
  OAI211_X1 U20859 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17644), .B(n17627), .ZN(n17629) );
  OAI211_X1 U20860 ( .C1(n17841), .C2(n17630), .A(n17629), .B(n17628), .ZN(
        n17631) );
  AOI211_X1 U20861 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n17639), .A(
        n17632), .B(n17631), .ZN(n17636) );
  NAND2_X1 U20862 ( .A1(n17860), .A2(n17993), .ZN(n17733) );
  AOI22_X1 U20863 ( .A1(n17895), .A2(n17634), .B1(n17917), .B2(n17633), .ZN(
        n17658) );
  NAND2_X1 U20864 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17658), .ZN(
        n17645) );
  NAND3_X1 U20865 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17733), .A3(
        n17645), .ZN(n17635) );
  OAI211_X1 U20866 ( .C1(n17774), .C2(n17637), .A(n17636), .B(n17635), .ZN(
        P3_U2802) );
  AOI22_X1 U20867 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17639), .B1(
        n17827), .B2(n17638), .ZN(n17649) );
  NOR2_X1 U20868 ( .A1(n17641), .A2(n17640), .ZN(n17642) );
  XNOR2_X1 U20869 ( .A(n17797), .B(n17642), .ZN(n18004) );
  AOI22_X1 U20870 ( .A1(n17882), .A2(n18004), .B1(n17644), .B2(n17643), .ZN(
        n17648) );
  OAI21_X1 U20871 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17646), .A(
        n17645), .ZN(n17647) );
  NAND2_X1 U20872 ( .A1(n18308), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n18006) );
  NAND4_X1 U20873 ( .A1(n17649), .A2(n17648), .A3(n17647), .A4(n18006), .ZN(
        P3_U2803) );
  NAND3_X1 U20874 ( .A1(n17994), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n17794), .ZN(n17659) );
  OAI21_X1 U20875 ( .B1(n17651), .B2(n18015), .A(n17650), .ZN(n18012) );
  NAND3_X1 U20876 ( .A1(n18719), .A2(n17663), .A3(n17662), .ZN(n17653) );
  AOI21_X1 U20877 ( .B1(n10073), .B2(n17653), .A(n17652), .ZN(n17656) );
  NAND2_X1 U20878 ( .A1(n18308), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n18013) );
  OAI221_X1 U20879 ( .B1(n17654), .B2(n17841), .C1(n17654), .C2(n17703), .A(
        n18013), .ZN(n17655) );
  AOI211_X1 U20880 ( .C1(n17882), .C2(n18012), .A(n17656), .B(n17655), .ZN(
        n17657) );
  OAI221_X1 U20881 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17659), 
        .C1(n18015), .C2(n17658), .A(n17657), .ZN(P3_U2804) );
  OAI21_X1 U20882 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17661), .A(
        n17660), .ZN(n18024) );
  NAND2_X1 U20883 ( .A1(n17663), .A2(n17785), .ZN(n17677) );
  AOI211_X1 U20884 ( .C1(n17676), .C2(n17666), .A(n17662), .B(n17677), .ZN(
        n17668) );
  OR2_X1 U20885 ( .A1(n18463), .A2(n17663), .ZN(n17688) );
  OAI211_X1 U20886 ( .C1(n17664), .C2(n17989), .A(n17988), .B(n17688), .ZN(
        n17690) );
  AOI21_X1 U20887 ( .B1(n17734), .B2(n17685), .A(n17690), .ZN(n17675) );
  OAI22_X1 U20888 ( .A1(n17675), .A2(n17666), .B1(n17841), .B2(n17665), .ZN(
        n17667) );
  AOI211_X1 U20889 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n18308), .A(n17668), 
        .B(n17667), .ZN(n17674) );
  XNOR2_X1 U20890 ( .A(n17669), .B(n18029), .ZN(n18017) );
  OAI21_X1 U20891 ( .B1(n17797), .B2(n17671), .A(n17670), .ZN(n17672) );
  XNOR2_X1 U20892 ( .A(n17672), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n18025) );
  AOI22_X1 U20893 ( .A1(n17917), .A2(n18017), .B1(n17882), .B2(n18025), .ZN(
        n17673) );
  OAI211_X1 U20894 ( .C1(n17860), .C2(n18024), .A(n17674), .B(n17673), .ZN(
        P3_U2805) );
  AOI22_X1 U20895 ( .A1(n17895), .A2(n18030), .B1(n17917), .B2(n18031), .ZN(
        n17694) );
  NAND2_X1 U20896 ( .A1(n18308), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n18039) );
  OAI221_X1 U20897 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n17677), .C1(
        n17676), .C2(n17675), .A(n18039), .ZN(n17678) );
  AOI21_X1 U20898 ( .B1(n17827), .B2(n17679), .A(n17678), .ZN(n17683) );
  OAI21_X1 U20899 ( .B1(n17680), .B2(n17684), .A(n11560), .ZN(n18038) );
  NOR2_X1 U20900 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17681), .ZN(
        n18036) );
  AOI22_X1 U20901 ( .A1(n17882), .A2(n18038), .B1(n17794), .B2(n18036), .ZN(
        n17682) );
  OAI211_X1 U20902 ( .C1(n17694), .C2(n17684), .A(n17683), .B(n17682), .ZN(
        P3_U2806) );
  NOR2_X1 U20903 ( .A1(n18312), .A2(n18909), .ZN(n18044) );
  NAND2_X1 U20904 ( .A1(n17734), .A2(n17685), .ZN(n17687) );
  AOI221_X1 U20905 ( .B1(n17983), .B2(n17688), .C1(n17687), .C2(n17688), .A(
        n17686), .ZN(n17689) );
  AOI211_X1 U20906 ( .C1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .C2(n17690), .A(
        n18044), .B(n17689), .ZN(n17699) );
  OAI22_X1 U20907 ( .A1(n17797), .A2(n18060), .B1(n17691), .B2(n17705), .ZN(
        n17692) );
  NOR2_X1 U20908 ( .A1(n17692), .A2(n17741), .ZN(n17693) );
  XNOR2_X1 U20909 ( .A(n17693), .B(n18048), .ZN(n18045) );
  NOR2_X1 U20910 ( .A1(n17996), .A2(n17774), .ZN(n17696) );
  INV_X1 U20911 ( .A(n17694), .ZN(n17695) );
  MUX2_X1 U20912 ( .A(n17696), .B(n17695), .S(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .Z(n17697) );
  AOI21_X1 U20913 ( .B1(n17882), .B2(n18045), .A(n17697), .ZN(n17698) );
  OAI211_X1 U20914 ( .C1(n17841), .C2(n17700), .A(n17699), .B(n17698), .ZN(
        P3_U2807) );
  INV_X1 U20915 ( .A(n18845), .ZN(n17948) );
  OAI22_X1 U20916 ( .A1(n17713), .A2(n17948), .B1(n17701), .B2(n17989), .ZN(
        n17702) );
  NOR2_X1 U20917 ( .A1(n17975), .A2(n17702), .ZN(n17735) );
  OAI21_X1 U20918 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17703), .A(
        n17735), .ZN(n17724) );
  AOI22_X1 U20919 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17724), .B1(
        n17827), .B2(n17704), .ZN(n17717) );
  INV_X1 U20920 ( .A(n17705), .ZN(n17707) );
  OR2_X1 U20921 ( .A1(n17757), .A2(n17706), .ZN(n18059) );
  AOI221_X1 U20922 ( .B1(n17708), .B2(n17707), .C1(n18059), .C2(n17707), .A(
        n17741), .ZN(n17709) );
  XNOR2_X1 U20923 ( .A(n17709), .B(n18060), .ZN(n18063) );
  NOR2_X1 U20924 ( .A1(n17774), .A2(n18059), .ZN(n17711) );
  OAI22_X1 U20925 ( .A1(n18135), .A2(n17860), .B1(n18140), .B2(n17993), .ZN(
        n17793) );
  AOI21_X1 U20926 ( .B1(n17733), .B2(n18059), .A(n17793), .ZN(n17732) );
  INV_X1 U20927 ( .A(n17732), .ZN(n17710) );
  MUX2_X1 U20928 ( .A(n17711), .B(n17710), .S(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(n17712) );
  AOI21_X1 U20929 ( .B1(n17882), .B2(n18063), .A(n17712), .ZN(n17716) );
  NAND2_X1 U20930 ( .A1(n18308), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18064) );
  AND2_X1 U20931 ( .A1(n17713), .A2(n17785), .ZN(n17719) );
  OAI211_X1 U20932 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17719), .B(n17714), .ZN(n17715) );
  NAND4_X1 U20933 ( .A1(n17717), .A2(n17716), .A3(n18064), .A4(n17715), .ZN(
        P3_U2808) );
  INV_X1 U20934 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17731) );
  NAND2_X1 U20935 ( .A1(n18308), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n18077) );
  INV_X1 U20936 ( .A(n18077), .ZN(n17723) );
  AOI22_X1 U20937 ( .A1(n17720), .A2(n17719), .B1(n17718), .B2(n17827), .ZN(
        n17721) );
  INV_X1 U20938 ( .A(n17721), .ZN(n17722) );
  AOI211_X1 U20939 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(n17724), .A(
        n17723), .B(n17722), .ZN(n17730) );
  INV_X1 U20940 ( .A(n18074), .ZN(n18057) );
  NAND3_X1 U20941 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17797), .A3(
        n17725), .ZN(n17751) );
  INV_X1 U20942 ( .A(n17726), .ZN(n17762) );
  OAI22_X1 U20943 ( .A1(n18057), .A2(n17751), .B1(n17762), .B2(n17727), .ZN(
        n17728) );
  XOR2_X1 U20944 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17728), .Z(
        n18070) );
  NOR2_X1 U20945 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18057), .ZN(
        n18069) );
  NAND2_X1 U20946 ( .A1(n18104), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18067) );
  NOR2_X1 U20947 ( .A1(n17774), .A2(n18067), .ZN(n17753) );
  AOI22_X1 U20948 ( .A1(n17882), .A2(n18070), .B1(n18069), .B2(n17753), .ZN(
        n17729) );
  OAI211_X1 U20949 ( .C1(n17732), .C2(n17731), .A(n17730), .B(n17729), .ZN(
        P3_U2809) );
  INV_X1 U20950 ( .A(n18067), .ZN(n18071) );
  NAND2_X1 U20951 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18071), .ZN(
        n18081) );
  AOI21_X1 U20952 ( .B1(n17733), .B2(n18081), .A(n17793), .ZN(n17756) );
  INV_X1 U20953 ( .A(n17973), .ZN(n17739) );
  AOI221_X1 U20954 ( .B1(n17737), .B2(n17736), .C1(n18463), .C2(n17736), .A(
        n17735), .ZN(n17738) );
  NOR2_X1 U20955 ( .A1(n18312), .A2(n18902), .ZN(n18087) );
  AOI211_X1 U20956 ( .C1(n17740), .C2(n17739), .A(n17738), .B(n18087), .ZN(
        n17745) );
  AOI221_X1 U20957 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17751), 
        .C1(n18096), .C2(n17761), .A(n17741), .ZN(n17742) );
  XOR2_X1 U20958 ( .A(n17742), .B(n18084), .Z(n18090) );
  INV_X1 U20959 ( .A(n18090), .ZN(n17743) );
  NOR2_X1 U20960 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18096), .ZN(
        n18088) );
  AOI22_X1 U20961 ( .A1(n17882), .A2(n17743), .B1(n17753), .B2(n18088), .ZN(
        n17744) );
  OAI211_X1 U20962 ( .C1(n17756), .C2(n18084), .A(n17745), .B(n17744), .ZN(
        P3_U2810) );
  INV_X1 U20963 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17749) );
  OAI21_X1 U20964 ( .B1(n17746), .B2(n17948), .A(n17988), .ZN(n17778) );
  AOI21_X1 U20965 ( .B1(n17824), .B2(n17747), .A(n17778), .ZN(n17758) );
  OAI22_X1 U20966 ( .A1(n17758), .A2(n17749), .B1(n17841), .B2(n17748), .ZN(
        n17750) );
  OAI21_X1 U20967 ( .B1(n17762), .B2(n17761), .A(n17751), .ZN(n17752) );
  XNOR2_X1 U20968 ( .A(n17752), .B(n18096), .ZN(n18092) );
  AOI22_X1 U20969 ( .A1(n17882), .A2(n18092), .B1(n17753), .B2(n18096), .ZN(
        n17754) );
  OAI211_X1 U20970 ( .C1(n17756), .C2(n18096), .A(n17755), .B(n17754), .ZN(
        P3_U2811) );
  AOI21_X1 U20971 ( .B1(n17794), .B2(n17757), .A(n17793), .ZN(n17780) );
  NAND2_X1 U20972 ( .A1(n18308), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18110) );
  OAI221_X1 U20973 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17760), .C1(
        n17759), .C2(n17758), .A(n18110), .ZN(n17766) );
  OAI21_X1 U20974 ( .B1(n17886), .B2(n18107), .A(n17761), .ZN(n17763) );
  XOR2_X1 U20975 ( .A(n17763), .B(n17762), .Z(n18109) );
  INV_X1 U20976 ( .A(n18109), .ZN(n17764) );
  NAND2_X1 U20977 ( .A1(n18104), .A2(n18107), .ZN(n18112) );
  OAI22_X1 U20978 ( .A1(n17898), .A2(n17764), .B1(n17774), .B2(n18112), .ZN(
        n17765) );
  AOI211_X1 U20979 ( .C1(n17827), .C2(n17767), .A(n17766), .B(n17765), .ZN(
        n17768) );
  OAI21_X1 U20980 ( .B1(n17780), .B2(n18107), .A(n17768), .ZN(P3_U2812) );
  OAI21_X1 U20981 ( .B1(n17770), .B2(n18463), .A(n17769), .ZN(n17777) );
  OAI22_X1 U20982 ( .A1(n17973), .A2(n17771), .B1(n18312), .B2(n18896), .ZN(
        n17776) );
  AOI21_X1 U20983 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17773), .A(
        n17772), .ZN(n18117) );
  NAND2_X1 U20984 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18113), .ZN(
        n18115) );
  OAI22_X1 U20985 ( .A1(n18117), .A2(n17898), .B1(n17774), .B2(n18115), .ZN(
        n17775) );
  AOI211_X1 U20986 ( .C1(n17778), .C2(n17777), .A(n17776), .B(n17775), .ZN(
        n17779) );
  OAI21_X1 U20987 ( .B1(n17780), .B2(n18113), .A(n17779), .ZN(P3_U2813) );
  OAI21_X1 U20988 ( .B1(n17886), .B2(n17782), .A(n17781), .ZN(n17783) );
  XNOR2_X1 U20989 ( .A(n17783), .B(n18127), .ZN(n18132) );
  INV_X1 U20990 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17803) );
  NOR2_X1 U20991 ( .A1(n17803), .A2(n17784), .ZN(n17791) );
  OAI211_X1 U20992 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17786), .B(n17785), .ZN(n17790) );
  INV_X1 U20993 ( .A(n17786), .ZN(n17799) );
  AOI21_X1 U20994 ( .B1(n18845), .B2(n17799), .A(n17975), .ZN(n17814) );
  OAI21_X1 U20995 ( .B1(n17787), .B2(n17989), .A(n17814), .ZN(n17802) );
  AOI22_X1 U20996 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17802), .B1(
        n17827), .B2(n17788), .ZN(n17789) );
  NAND2_X1 U20997 ( .A1(n18308), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n18130) );
  OAI211_X1 U20998 ( .C1(n17791), .C2(n17790), .A(n17789), .B(n18130), .ZN(
        n17792) );
  AOI221_X1 U20999 ( .B1(n17794), .B2(n18127), .C1(n17793), .C2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n17792), .ZN(n17795) );
  OAI21_X1 U21000 ( .B1(n17898), .B2(n18132), .A(n17795), .ZN(P3_U2814) );
  NAND2_X1 U21001 ( .A1(n17797), .A2(n18186), .ZN(n17875) );
  NOR2_X1 U21002 ( .A1(n18163), .A2(n17875), .ZN(n17846) );
  NAND2_X1 U21003 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17846), .ZN(
        n17819) );
  NOR2_X1 U21004 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17851), .ZN(
        n18162) );
  AOI221_X1 U21005 ( .B1(n11554), .B2(n17796), .C1(n17819), .C2(n17796), .A(
        n18162), .ZN(n17798) );
  XNOR2_X1 U21006 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17798), .ZN(
        n18146) );
  NOR2_X1 U21007 ( .A1(n17834), .A2(n17799), .ZN(n17804) );
  OAI22_X1 U21008 ( .A1(n18312), .A2(n18892), .B1(n17841), .B2(n17800), .ZN(
        n17801) );
  AOI221_X1 U21009 ( .B1(n17804), .B2(n17803), .C1(n17802), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17801), .ZN(n17808) );
  NOR2_X1 U21010 ( .A1(n18135), .A2(n17860), .ZN(n17806) );
  NAND2_X1 U21011 ( .A1(n11555), .A2(n17809), .ZN(n18134) );
  NOR2_X1 U21012 ( .A1(n18140), .A2(n17993), .ZN(n17805) );
  INV_X1 U21013 ( .A(n18122), .ZN(n18124) );
  OAI21_X1 U21014 ( .B1(n17817), .B2(n18124), .A(n11555), .ZN(n18141) );
  AOI22_X1 U21015 ( .A1(n17806), .A2(n18134), .B1(n17805), .B2(n18141), .ZN(
        n17807) );
  OAI211_X1 U21016 ( .C1(n17898), .C2(n18146), .A(n17808), .B(n17807), .ZN(
        P3_U2815) );
  OAI21_X1 U21017 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17810), .A(
        n17809), .ZN(n18153) );
  NOR2_X1 U21018 ( .A1(n18463), .A2(n17833), .ZN(n17858) );
  AOI21_X1 U21019 ( .B1(n17811), .B2(n17858), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17813) );
  OAI22_X1 U21020 ( .A1(n17814), .A2(n17813), .B1(n17973), .B2(n17812), .ZN(
        n17815) );
  AOI21_X1 U21021 ( .B1(n18308), .B2(P3_REIP_REG_14__SCAN_IN), .A(n17815), 
        .ZN(n17822) );
  NOR2_X1 U21022 ( .A1(n17817), .A2(n18124), .ZN(n17816) );
  AOI221_X1 U21023 ( .B1(n17817), .B2(n11554), .C1(n18148), .C2(n11554), .A(
        n17816), .ZN(n18158) );
  AOI21_X1 U21024 ( .B1(n17819), .B2(n17818), .A(n18162), .ZN(n17820) );
  XNOR2_X1 U21025 ( .A(n17820), .B(n11554), .ZN(n18157) );
  AOI22_X1 U21026 ( .A1(n17917), .A2(n18158), .B1(n17882), .B2(n18157), .ZN(
        n17821) );
  OAI211_X1 U21027 ( .C1(n17860), .C2(n18153), .A(n17822), .B(n17821), .ZN(
        P3_U2816) );
  AOI22_X1 U21028 ( .A1(n17824), .A2(n17823), .B1(n18845), .B2(n17833), .ZN(
        n17825) );
  NAND2_X1 U21029 ( .A1(n17825), .A2(n17988), .ZN(n17843) );
  AOI22_X1 U21030 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17843), .B1(
        n17827), .B2(n17826), .ZN(n17839) );
  NOR2_X1 U21031 ( .A1(n17885), .A2(n18163), .ZN(n17848) );
  NAND2_X1 U21032 ( .A1(n18176), .A2(n18186), .ZN(n18165) );
  NAND2_X1 U21033 ( .A1(n18176), .A2(n18184), .ZN(n18169) );
  AOI22_X1 U21034 ( .A1(n17895), .A2(n18165), .B1(n17917), .B2(n18169), .ZN(
        n17852) );
  NAND2_X1 U21035 ( .A1(n17851), .A2(n17886), .ZN(n17830) );
  INV_X1 U21036 ( .A(n17828), .ZN(n17829) );
  AOI22_X1 U21037 ( .A1(n17830), .A2(n18165), .B1(n17829), .B2(n17886), .ZN(
        n17831) );
  XNOR2_X1 U21038 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n17831), .ZN(
        n18174) );
  OAI22_X1 U21039 ( .A1(n17852), .A2(n18152), .B1(n17898), .B2(n18174), .ZN(
        n17832) );
  AOI21_X1 U21040 ( .B1(n18162), .B2(n17848), .A(n17832), .ZN(n17838) );
  NAND2_X1 U21041 ( .A1(n9822), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n17837) );
  NOR2_X1 U21042 ( .A1(n17834), .A2(n17833), .ZN(n17845) );
  OAI211_X1 U21043 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17845), .B(n17835), .ZN(n17836) );
  NAND4_X1 U21044 ( .A1(n17839), .A2(n17838), .A3(n17837), .A4(n17836), .ZN(
        P3_U2817) );
  OAI22_X1 U21045 ( .A1(n18312), .A2(n18886), .B1(n17841), .B2(n17840), .ZN(
        n17842) );
  AOI221_X1 U21046 ( .B1(n17845), .B2(n17844), .C1(n17843), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n17842), .ZN(n17850) );
  NOR2_X1 U21047 ( .A1(n17846), .A2(n17828), .ZN(n17847) );
  XNOR2_X1 U21048 ( .A(n17847), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n18175) );
  AOI22_X1 U21049 ( .A1(n17882), .A2(n18175), .B1(n17848), .B2(n17851), .ZN(
        n17849) );
  OAI211_X1 U21050 ( .C1(n17852), .C2(n17851), .A(n17850), .B(n17849), .ZN(
        P3_U2818) );
  NAND2_X1 U21051 ( .A1(n18189), .A2(n18193), .ZN(n18199) );
  INV_X1 U21052 ( .A(n17875), .ZN(n17854) );
  AOI21_X1 U21053 ( .B1(n18189), .B2(n17854), .A(n17853), .ZN(n17855) );
  XNOR2_X1 U21054 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n17855), .ZN(
        n18197) );
  INV_X1 U21055 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18884) );
  NOR2_X1 U21056 ( .A1(n18312), .A2(n18884), .ZN(n18196) );
  NAND2_X1 U21057 ( .A1(n17988), .A2(n17948), .ZN(n17984) );
  NAND3_X1 U21058 ( .A1(n18719), .A2(n17919), .A3(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17901) );
  NOR3_X1 U21059 ( .A1(n17903), .A2(n17888), .A3(n17901), .ZN(n17878) );
  NAND2_X1 U21060 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17878), .ZN(
        n17877) );
  NOR2_X1 U21061 ( .A1(n17865), .A2(n17877), .ZN(n17864) );
  AOI21_X1 U21062 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17984), .A(
        n17864), .ZN(n17857) );
  OAI22_X1 U21063 ( .A1(n17858), .A2(n17857), .B1(n17973), .B2(n17856), .ZN(
        n17859) );
  AOI211_X1 U21064 ( .C1(n17882), .C2(n18197), .A(n18196), .B(n17859), .ZN(
        n17862) );
  NOR2_X1 U21065 ( .A1(n18189), .A2(n17885), .ZN(n17872) );
  OAI22_X1 U21066 ( .A1(n18186), .A2(n17860), .B1(n18184), .B2(n17993), .ZN(
        n17863) );
  OAI21_X1 U21067 ( .B1(n17872), .B2(n17863), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17861) );
  OAI211_X1 U21068 ( .C1(n17885), .C2(n18199), .A(n17862), .B(n17861), .ZN(
        P3_U2819) );
  INV_X1 U21069 ( .A(n17863), .ZN(n17884) );
  INV_X1 U21070 ( .A(n17984), .ZN(n17918) );
  AOI211_X1 U21071 ( .C1(n17877), .C2(n17865), .A(n17918), .B(n17864), .ZN(
        n17867) );
  NOR2_X1 U21072 ( .A1(n18312), .A2(n18882), .ZN(n17866) );
  AOI211_X1 U21073 ( .C1(n17868), .C2(n17739), .A(n17867), .B(n17866), .ZN(
        n17874) );
  AOI22_X1 U21074 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17875), .B1(
        n17869), .B2(n18214), .ZN(n17870) );
  XNOR2_X1 U21075 ( .A(n18205), .B(n17870), .ZN(n18200) );
  NAND2_X1 U21076 ( .A1(n18214), .A2(n18205), .ZN(n17871) );
  AOI22_X1 U21077 ( .A1(n17882), .A2(n18200), .B1(n17872), .B2(n17871), .ZN(
        n17873) );
  OAI211_X1 U21078 ( .C1(n17884), .C2(n18205), .A(n17874), .B(n17873), .ZN(
        P3_U2820) );
  NAND2_X1 U21079 ( .A1(n17875), .A2(n17869), .ZN(n17876) );
  XNOR2_X1 U21080 ( .A(n17876), .B(n18214), .ZN(n18218) );
  OAI211_X1 U21081 ( .C1(n17878), .C2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n17984), .B(n17877), .ZN(n17879) );
  NAND2_X1 U21082 ( .A1(n18308), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n18220) );
  OAI211_X1 U21083 ( .C1(n17973), .C2(n17880), .A(n17879), .B(n18220), .ZN(
        n17881) );
  AOI21_X1 U21084 ( .B1(n17882), .B2(n18218), .A(n17881), .ZN(n17883) );
  OAI221_X1 U21085 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17885), .C1(
        n18214), .C2(n17884), .A(n17883), .ZN(P3_U2821) );
  NOR2_X1 U21086 ( .A1(n18186), .A2(n9975), .ZN(n18228) );
  XNOR2_X1 U21087 ( .A(n18228), .B(n17886), .ZN(n18238) );
  OAI21_X1 U21088 ( .B1(n17887), .B2(n17948), .A(n17988), .ZN(n17902) );
  OAI221_X1 U21089 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n17889), .C1(
        n17888), .C2(n17903), .A(n18719), .ZN(n17890) );
  NAND2_X1 U21090 ( .A1(n18308), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n18235) );
  OAI211_X1 U21091 ( .C1(n17973), .C2(n17891), .A(n17890), .B(n18235), .ZN(
        n17892) );
  AOI21_X1 U21092 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n17902), .A(
        n17892), .ZN(n17897) );
  AOI21_X1 U21093 ( .B1(n17894), .B2(n10241), .A(n17893), .ZN(n18230) );
  AOI22_X1 U21094 ( .A1(n17895), .A2(n18228), .B1(n17917), .B2(n18230), .ZN(
        n17896) );
  OAI211_X1 U21095 ( .C1(n18238), .C2(n17898), .A(n17897), .B(n17896), .ZN(
        P3_U2822) );
  OAI21_X1 U21096 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17900), .A(
        n17899), .ZN(n18247) );
  INV_X1 U21097 ( .A(n17901), .ZN(n17904) );
  NOR2_X1 U21098 ( .A1(n18312), .A2(n18876), .ZN(n18243) );
  AOI221_X1 U21099 ( .B1(n17904), .B2(n17903), .C1(n17902), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18243), .ZN(n17911) );
  OAI21_X1 U21100 ( .B1(n17907), .B2(n17906), .A(n17905), .ZN(n17908) );
  XNOR2_X1 U21101 ( .A(n17908), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18244) );
  AOI22_X1 U21102 ( .A1(n17917), .A2(n18244), .B1(n17909), .B2(n17739), .ZN(
        n17910) );
  OAI211_X1 U21103 ( .C1(n17992), .C2(n18247), .A(n17911), .B(n17910), .ZN(
        P3_U2823) );
  NAND2_X1 U21104 ( .A1(n18719), .A2(n17919), .ZN(n17927) );
  AOI22_X1 U21105 ( .A1(n17914), .A2(n17932), .B1(n17913), .B2(n17912), .ZN(
        n17915) );
  XNOR2_X1 U21106 ( .A(n17916), .B(n17915), .ZN(n18250) );
  AOI22_X1 U21107 ( .A1(n9822), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n17917), .B2(
        n18250), .ZN(n17926) );
  AOI21_X1 U21108 ( .B1(n17919), .B2(n18719), .A(n17918), .ZN(n17938) );
  OAI21_X1 U21109 ( .B1(n17922), .B2(n17921), .A(n17920), .ZN(n18255) );
  OAI22_X1 U21110 ( .A1(n17973), .A2(n17923), .B1(n17992), .B2(n18255), .ZN(
        n17924) );
  AOI21_X1 U21111 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17938), .A(
        n17924), .ZN(n17925) );
  OAI211_X1 U21112 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n17927), .A(
        n17926), .B(n17925), .ZN(P3_U2824) );
  OAI21_X1 U21113 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n17929), .A(
        n17928), .ZN(n18256) );
  OAI21_X1 U21114 ( .B1(n17975), .B2(n17931), .A(n17930), .ZN(n17937) );
  OAI21_X1 U21115 ( .B1(n17934), .B2(n17933), .A(n17932), .ZN(n18263) );
  OAI22_X1 U21116 ( .A1(n17973), .A2(n17935), .B1(n17993), .B2(n18263), .ZN(
        n17936) );
  AOI21_X1 U21117 ( .B1(n17938), .B2(n17937), .A(n17936), .ZN(n17939) );
  NAND2_X1 U21118 ( .A1(n9822), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n18261) );
  OAI211_X1 U21119 ( .C1(n17992), .C2(n18256), .A(n17939), .B(n18261), .ZN(
        P3_U2825) );
  OAI21_X1 U21120 ( .B1(n17942), .B2(n17941), .A(n17940), .ZN(n18269) );
  OAI21_X1 U21121 ( .B1(n17945), .B2(n17944), .A(n17943), .ZN(n18275) );
  OAI22_X1 U21122 ( .A1(n17992), .A2(n18275), .B1(n18463), .B2(n17946), .ZN(
        n17947) );
  AOI21_X1 U21123 ( .B1(n18308), .B2(P3_REIP_REG_4__SCAN_IN), .A(n17947), .ZN(
        n17952) );
  OAI21_X1 U21124 ( .B1(n17949), .B2(n17948), .A(n17988), .ZN(n17964) );
  AOI22_X1 U21125 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17964), .B1(
        n17950), .B2(n17739), .ZN(n17951) );
  OAI211_X1 U21126 ( .C1(n17993), .C2(n18269), .A(n17952), .B(n17951), .ZN(
        P3_U2826) );
  OAI21_X1 U21127 ( .B1(n17955), .B2(n17954), .A(n17953), .ZN(n17957) );
  XNOR2_X1 U21128 ( .A(n17957), .B(n17956), .ZN(n18283) );
  NOR2_X1 U21129 ( .A1(n17975), .A2(n17976), .ZN(n17963) );
  OAI21_X1 U21130 ( .B1(n17960), .B2(n17959), .A(n17958), .ZN(n18277) );
  OAI22_X1 U21131 ( .A1(n17973), .A2(n17961), .B1(n17993), .B2(n18277), .ZN(
        n17962) );
  AOI221_X1 U21132 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17964), .C1(
        n17963), .C2(n17964), .A(n17962), .ZN(n17965) );
  NAND2_X1 U21133 ( .A1(n18308), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18281) );
  OAI211_X1 U21134 ( .C1(n17992), .C2(n18283), .A(n17965), .B(n18281), .ZN(
        P3_U2827) );
  OAI21_X1 U21135 ( .B1(n17968), .B2(n17967), .A(n17966), .ZN(n18298) );
  OAI21_X1 U21136 ( .B1(n17971), .B2(n17970), .A(n17969), .ZN(n18290) );
  OAI22_X1 U21137 ( .A1(n17973), .A2(n17972), .B1(n17993), .B2(n18290), .ZN(
        n17974) );
  AOI221_X1 U21138 ( .B1(n18719), .B2(n17976), .C1(n17975), .C2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n17974), .ZN(n17977) );
  NAND2_X1 U21139 ( .A1(n9822), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18296) );
  OAI211_X1 U21140 ( .C1(n17992), .C2(n18298), .A(n17977), .B(n18296), .ZN(
        P3_U2828) );
  NOR2_X1 U21141 ( .A1(n17978), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17979) );
  XNOR2_X1 U21142 ( .A(n17979), .B(n17981), .ZN(n18305) );
  OAI21_X1 U21143 ( .B1(n17981), .B2(n17986), .A(n17980), .ZN(n18303) );
  OAI22_X1 U21144 ( .A1(n18312), .A2(n18974), .B1(n17992), .B2(n18303), .ZN(
        n17982) );
  AOI221_X1 U21145 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17984), .C1(
        n17983), .C2(n17739), .A(n17982), .ZN(n17985) );
  OAI21_X1 U21146 ( .B1(n18305), .B2(n17993), .A(n17985), .ZN(P3_U2829) );
  AOI21_X1 U21147 ( .B1(n17987), .B2(n18300), .A(n17986), .ZN(n18316) );
  INV_X1 U21148 ( .A(n18316), .ZN(n18314) );
  NAND3_X1 U21149 ( .A1(n18965), .A2(n17989), .A3(n17988), .ZN(n17990) );
  AOI22_X1 U21150 ( .A1(n9822), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17990), .ZN(n17991) );
  OAI221_X1 U21151 ( .B1(n18316), .B2(n17993), .C1(n18314), .C2(n17992), .A(
        n17991), .ZN(P3_U2830) );
  NAND3_X1 U21152 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17994), .A3(
        n18042), .ZN(n18010) );
  NOR2_X1 U21153 ( .A1(n18015), .A2(n18010), .ZN(n18003) );
  NOR2_X1 U21154 ( .A1(n17995), .A2(n18285), .ZN(n18000) );
  NAND2_X1 U21155 ( .A1(n18300), .A2(n18797), .ZN(n18286) );
  NAND2_X1 U21156 ( .A1(n18050), .A2(n18286), .ZN(n18102) );
  NOR2_X1 U21157 ( .A1(n17996), .A2(n18102), .ZN(n18055) );
  AOI21_X1 U21158 ( .B1(n18019), .B2(n18055), .A(n18285), .ZN(n18021) );
  OAI22_X1 U21159 ( .A1(n17998), .A2(n18776), .B1(n17997), .B2(n18185), .ZN(
        n17999) );
  NOR4_X1 U21160 ( .A1(n18001), .A2(n18000), .A3(n18021), .A4(n17999), .ZN(
        n18009) );
  INV_X1 U21161 ( .A(n18009), .ZN(n18002) );
  MUX2_X1 U21162 ( .A(n18003), .B(n18002), .S(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .Z(n18005) );
  AOI22_X1 U21163 ( .A1(n9802), .A2(n18005), .B1(n18219), .B2(n18004), .ZN(
        n18007) );
  OAI211_X1 U21164 ( .C1(n18008), .C2(n18310), .A(n18007), .B(n18006), .ZN(
        P3_U2835) );
  AOI211_X1 U21165 ( .C1(n18015), .C2(n18010), .A(n18009), .B(n10081), .ZN(
        n18011) );
  AOI21_X1 U21166 ( .B1(n18219), .B2(n18012), .A(n18011), .ZN(n18014) );
  OAI211_X1 U21167 ( .C1(n18310), .C2(n18015), .A(n18014), .B(n18013), .ZN(
        P3_U2836) );
  AOI22_X1 U21168 ( .A1(n18017), .A2(n18231), .B1(n18016), .B2(n18029), .ZN(
        n18023) );
  NAND2_X1 U21169 ( .A1(n18053), .A2(n18104), .ZN(n18106) );
  OAI21_X1 U21170 ( .B1(n18018), .B2(n18106), .A(n18811), .ZN(n18033) );
  OAI21_X1 U21171 ( .B1(n18019), .B2(n18792), .A(n18033), .ZN(n18020) );
  OAI21_X1 U21172 ( .B1(n18021), .B2(n18020), .A(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18022) );
  OAI211_X1 U21173 ( .C1(n18024), .C2(n18185), .A(n18023), .B(n18022), .ZN(
        n18026) );
  AOI22_X1 U21174 ( .A1(n9802), .A2(n18026), .B1(n18219), .B2(n18025), .ZN(
        n18028) );
  NAND2_X1 U21175 ( .A1(n18308), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n18027) );
  OAI211_X1 U21176 ( .C1(n18310), .C2(n18029), .A(n18028), .B(n18027), .ZN(
        P3_U2837) );
  AOI22_X1 U21177 ( .A1(n18231), .A2(n18031), .B1(n18229), .B2(n18030), .ZN(
        n18032) );
  OAI211_X1 U21178 ( .C1(n18285), .C2(n18055), .A(n18032), .B(n18310), .ZN(
        n18035) );
  NAND2_X1 U21179 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n18033), .ZN(
        n18034) );
  OAI21_X1 U21180 ( .B1(n18035), .B2(n18034), .A(n18312), .ZN(n18049) );
  OAI21_X1 U21181 ( .B1(n18268), .B2(n18035), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18041) );
  INV_X1 U21182 ( .A(n18068), .ZN(n18037) );
  AOI22_X1 U21183 ( .A1(n18219), .A2(n18038), .B1(n18037), .B2(n18036), .ZN(
        n18040) );
  OAI211_X1 U21184 ( .C1(n18049), .C2(n18041), .A(n18040), .B(n18039), .ZN(
        P3_U2838) );
  NAND3_X1 U21185 ( .A1(n18043), .A2(n18042), .A3(n18310), .ZN(n18047) );
  AOI21_X1 U21186 ( .B1(n18045), .B2(n18219), .A(n18044), .ZN(n18046) );
  OAI221_X1 U21187 ( .B1(n18049), .B2(n18048), .C1(n18049), .C2(n18047), .A(
        n18046), .ZN(P3_U2839) );
  NAND2_X1 U21188 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18312), .ZN(
        n18066) );
  NAND2_X1 U21189 ( .A1(n18776), .A2(n18185), .ZN(n18100) );
  NOR2_X1 U21190 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18799), .ZN(
        n18054) );
  INV_X1 U21191 ( .A(n18050), .ZN(n18051) );
  OAI22_X1 U21192 ( .A1(n18140), .A2(n18776), .B1(n18135), .B2(n18185), .ZN(
        n18101) );
  AOI221_X1 U21193 ( .B1(n18051), .B2(n18791), .C1(n18081), .C2(n18791), .A(
        n18101), .ZN(n18052) );
  OAI221_X1 U21194 ( .B1(n18792), .B2(n18053), .C1(n18792), .C2(n18071), .A(
        n18052), .ZN(n18079) );
  AOI211_X1 U21195 ( .C1(n18059), .C2(n18100), .A(n18054), .B(n18079), .ZN(
        n18073) );
  AOI21_X1 U21196 ( .B1(n18190), .B2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n18055), .ZN(n18056) );
  AOI21_X1 U21197 ( .B1(n18811), .B2(n18057), .A(n18056), .ZN(n18058) );
  OAI211_X1 U21198 ( .C1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n18202), .A(
        n18073), .B(n18058), .ZN(n18062) );
  OAI22_X1 U21199 ( .A1(n9822), .A2(n18060), .B1(n18059), .B2(n18068), .ZN(
        n18061) );
  AOI22_X1 U21200 ( .A1(n18219), .A2(n18063), .B1(n18062), .B2(n18061), .ZN(
        n18065) );
  OAI211_X1 U21201 ( .C1(n9802), .C2(n18066), .A(n18065), .B(n18064), .ZN(
        P3_U2840) );
  NOR2_X1 U21202 ( .A1(n18068), .A2(n18067), .ZN(n18091) );
  AOI22_X1 U21203 ( .A1(n18219), .A2(n18070), .B1(n18069), .B2(n18091), .ZN(
        n18078) );
  OAI221_X1 U21204 ( .B1(n18190), .B2(n18072), .C1(n18190), .C2(n18071), .A(
        n9802), .ZN(n18080) );
  NOR2_X1 U21205 ( .A1(n18811), .A2(n18797), .ZN(n18083) );
  OAI21_X1 U21206 ( .B1(n18074), .B2(n18083), .A(n18073), .ZN(n18075) );
  OAI211_X1 U21207 ( .C1(n18080), .C2(n18075), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18312), .ZN(n18076) );
  NAND3_X1 U21208 ( .A1(n18078), .A2(n18077), .A3(n18076), .ZN(P3_U2841) );
  AOI211_X1 U21209 ( .C1(n18081), .C2(n18100), .A(n18080), .B(n18079), .ZN(
        n18082) );
  OR2_X1 U21210 ( .A1(n9822), .A2(n18082), .ZN(n18095) );
  INV_X1 U21211 ( .A(n18083), .ZN(n18299) );
  NAND3_X1 U21212 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18096), .A3(n18299), 
        .ZN(n18085) );
  AOI21_X1 U21213 ( .B1(n18095), .B2(n18085), .A(n18084), .ZN(n18086) );
  AOI211_X1 U21214 ( .C1(n18088), .C2(n18091), .A(n18087), .B(n18086), .ZN(
        n18089) );
  OAI21_X1 U21215 ( .B1(n18237), .B2(n18090), .A(n18089), .ZN(P3_U2842) );
  AOI22_X1 U21216 ( .A1(n18219), .A2(n18092), .B1(n18091), .B2(n18096), .ZN(
        n18094) );
  NAND2_X1 U21217 ( .A1(n18308), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18093) );
  OAI211_X1 U21218 ( .C1(n18096), .C2(n18095), .A(n18094), .B(n18093), .ZN(
        P3_U2843) );
  INV_X1 U21219 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18241) );
  NAND2_X1 U21220 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18267) );
  INV_X1 U21221 ( .A(n18097), .ZN(n18287) );
  OAI22_X1 U21222 ( .A1(n18264), .A2(n18792), .B1(n18267), .B2(n18287), .ZN(
        n18276) );
  NAND3_X1 U21223 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18252), .A3(
        n18276), .ZN(n18240) );
  NOR2_X1 U21224 ( .A1(n18241), .A2(n18240), .ZN(n18223) );
  NAND2_X1 U21225 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18223), .ZN(
        n18133) );
  AOI21_X1 U21226 ( .B1(n18098), .B2(n18133), .A(n10081), .ZN(n18206) );
  INV_X1 U21227 ( .A(n18206), .ZN(n18222) );
  NOR2_X1 U21228 ( .A1(n18099), .A2(n18222), .ZN(n18128) );
  INV_X1 U21229 ( .A(n18128), .ZN(n18116) );
  INV_X1 U21230 ( .A(n18100), .ZN(n18188) );
  NOR2_X1 U21231 ( .A1(n10081), .A2(n18101), .ZN(n18125) );
  INV_X1 U21232 ( .A(n18285), .ZN(n18266) );
  OAI21_X1 U21233 ( .B1(n18127), .B2(n18102), .A(n18266), .ZN(n18103) );
  OAI211_X1 U21234 ( .C1(n18104), .C2(n18188), .A(n18125), .B(n18103), .ZN(
        n18105) );
  AOI21_X1 U21235 ( .B1(n18811), .B2(n18106), .A(n18105), .ZN(n18114) );
  AOI221_X1 U21236 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18114), 
        .C1(n18285), .C2(n18114), .A(n18107), .ZN(n18108) );
  AOI22_X1 U21237 ( .A1(n18109), .A2(n18219), .B1(n18108), .B2(n18312), .ZN(
        n18111) );
  OAI211_X1 U21238 ( .C1(n18112), .C2(n18116), .A(n18111), .B(n18110), .ZN(
        P3_U2844) );
  NOR2_X1 U21239 ( .A1(n18312), .A2(n18896), .ZN(n18120) );
  NOR3_X1 U21240 ( .A1(n9822), .A2(n18114), .A3(n18113), .ZN(n18119) );
  OAI22_X1 U21241 ( .A1(n18117), .A2(n18237), .B1(n18116), .B2(n18115), .ZN(
        n18118) );
  OR3_X1 U21242 ( .A1(n18120), .A2(n18119), .A3(n18118), .ZN(P3_U2845) );
  NAND2_X1 U21243 ( .A1(n18811), .A2(n18121), .ZN(n18166) );
  NAND2_X1 U21244 ( .A1(n18190), .A2(n18166), .ZN(n18212) );
  NAND2_X1 U21245 ( .A1(n18149), .A2(n18791), .ZN(n18210) );
  OAI211_X1 U21246 ( .C1(n18122), .C2(n18202), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n18210), .ZN(n18123) );
  AOI221_X1 U21247 ( .B1(n18124), .B2(n18212), .C1(n18211), .C2(n18212), .A(
        n18123), .ZN(n18139) );
  AOI221_X1 U21248 ( .B1(n18126), .B2(n18125), .C1(n18139), .C2(n18125), .A(
        n9822), .ZN(n18129) );
  AOI22_X1 U21249 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18129), .B1(
        n18128), .B2(n18127), .ZN(n18131) );
  OAI211_X1 U21250 ( .C1(n18132), .C2(n18237), .A(n18131), .B(n18130), .ZN(
        P3_U2846) );
  AOI22_X1 U21251 ( .A1(n9822), .A2(P3_REIP_REG_15__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18294), .ZN(n18145) );
  NOR2_X1 U21252 ( .A1(n18148), .A2(n18133), .ZN(n18156) );
  AOI21_X1 U21253 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18156), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18138) );
  INV_X1 U21254 ( .A(n18134), .ZN(n18137) );
  OR2_X1 U21255 ( .A1(n18185), .A2(n18135), .ZN(n18136) );
  OAI22_X1 U21256 ( .A1(n18139), .A2(n18138), .B1(n18137), .B2(n18136), .ZN(
        n18143) );
  NOR2_X1 U21257 ( .A1(n18140), .A2(n18304), .ZN(n18142) );
  AOI22_X1 U21258 ( .A1(n9802), .A2(n18143), .B1(n18142), .B2(n18141), .ZN(
        n18144) );
  OAI211_X1 U21259 ( .C1(n18237), .C2(n18146), .A(n18145), .B(n18144), .ZN(
        P3_U2847) );
  AOI21_X1 U21260 ( .B1(n18176), .B2(n18147), .A(n18190), .ZN(n18171) );
  OAI21_X1 U21261 ( .B1(n18149), .B2(n18148), .A(n18791), .ZN(n18150) );
  OAI211_X1 U21262 ( .C1(n18176), .C2(n18792), .A(n18166), .B(n18150), .ZN(
        n18151) );
  AOI211_X1 U21263 ( .C1(n18152), .C2(n18299), .A(n18171), .B(n18151), .ZN(
        n18154) );
  OAI22_X1 U21264 ( .A1(n18154), .A2(n11554), .B1(n18185), .B2(n18153), .ZN(
        n18155) );
  AOI21_X1 U21265 ( .B1(n18156), .B2(n11554), .A(n18155), .ZN(n18161) );
  AOI22_X1 U21266 ( .A1(n9822), .A2(P3_REIP_REG_14__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18294), .ZN(n18160) );
  INV_X1 U21267 ( .A(n18304), .ZN(n18315) );
  AOI22_X1 U21268 ( .A1(n18315), .A2(n18158), .B1(n18219), .B2(n18157), .ZN(
        n18159) );
  OAI211_X1 U21269 ( .C1(n18161), .C2(n10081), .A(n18160), .B(n18159), .ZN(
        P3_U2848) );
  NOR2_X1 U21270 ( .A1(n18163), .A2(n18222), .ZN(n18181) );
  AOI22_X1 U21271 ( .A1(n9822), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18162), 
        .B2(n18181), .ZN(n18173) );
  INV_X1 U21272 ( .A(n18163), .ZN(n18164) );
  AOI21_X1 U21273 ( .B1(n18164), .B2(n18210), .A(n18202), .ZN(n18192) );
  INV_X1 U21274 ( .A(n18165), .ZN(n18167) );
  OAI21_X1 U21275 ( .B1(n18167), .B2(n18185), .A(n18166), .ZN(n18168) );
  AOI211_X1 U21276 ( .C1(n18231), .C2(n18169), .A(n18192), .B(n18168), .ZN(
        n18178) );
  OAI211_X1 U21277 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n18202), .A(
        n9802), .B(n18178), .ZN(n18170) );
  OAI211_X1 U21278 ( .C1(n18171), .C2(n18170), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18312), .ZN(n18172) );
  OAI211_X1 U21279 ( .C1(n18237), .C2(n18174), .A(n18173), .B(n18172), .ZN(
        P3_U2849) );
  AOI22_X1 U21280 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18294), .B1(
        n18219), .B2(n18175), .ZN(n18183) );
  INV_X1 U21281 ( .A(n18176), .ZN(n18177) );
  NOR2_X1 U21282 ( .A1(n18177), .A2(n18211), .ZN(n18179) );
  OAI211_X1 U21283 ( .C1(n18179), .C2(n18190), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n18178), .ZN(n18180) );
  OAI211_X1 U21284 ( .C1(n18181), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n9802), .B(n18180), .ZN(n18182) );
  OAI211_X1 U21285 ( .C1(n18886), .C2(n18312), .A(n18183), .B(n18182), .ZN(
        P3_U2850) );
  OAI22_X1 U21286 ( .A1(n18186), .A2(n18185), .B1(n18776), .B2(n18184), .ZN(
        n18201) );
  OAI21_X1 U21287 ( .B1(n18211), .B2(n18214), .A(n18212), .ZN(n18187) );
  OAI21_X1 U21288 ( .B1(n18189), .B2(n18188), .A(n18187), .ZN(n18204) );
  OAI21_X1 U21289 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n18190), .A(
        n9802), .ZN(n18191) );
  NOR4_X1 U21290 ( .A1(n18192), .A2(n18201), .A3(n18204), .A4(n18191), .ZN(
        n18194) );
  NOR3_X1 U21291 ( .A1(n9822), .A2(n18194), .A3(n18193), .ZN(n18195) );
  AOI211_X1 U21292 ( .C1(n18219), .C2(n18197), .A(n18196), .B(n18195), .ZN(
        n18198) );
  OAI21_X1 U21293 ( .B1(n18222), .B2(n18199), .A(n18198), .ZN(P3_U2851) );
  AOI22_X1 U21294 ( .A1(n9822), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18219), 
        .B2(n18200), .ZN(n18209) );
  NOR2_X1 U21295 ( .A1(n18294), .A2(n18201), .ZN(n18216) );
  OAI211_X1 U21296 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18202), .A(
        n18216), .B(n18210), .ZN(n18203) );
  OAI211_X1 U21297 ( .C1(n18204), .C2(n18203), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n18312), .ZN(n18208) );
  NAND3_X1 U21298 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18206), .A3(
        n18205), .ZN(n18207) );
  NAND3_X1 U21299 ( .A1(n18209), .A2(n18208), .A3(n18207), .ZN(P3_U2852) );
  INV_X1 U21300 ( .A(n18210), .ZN(n18213) );
  OAI21_X1 U21301 ( .B1(n18213), .B2(n18212), .A(n18211), .ZN(n18215) );
  AOI211_X1 U21302 ( .C1(n18216), .C2(n18215), .A(n9822), .B(n18214), .ZN(
        n18217) );
  AOI21_X1 U21303 ( .B1(n18219), .B2(n18218), .A(n18217), .ZN(n18221) );
  OAI211_X1 U21304 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18222), .A(
        n18221), .B(n18220), .ZN(P3_U2853) );
  INV_X1 U21305 ( .A(n18223), .ZN(n18233) );
  NAND2_X1 U21306 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18227) );
  NAND2_X1 U21307 ( .A1(n18224), .A2(n18266), .ZN(n18225) );
  OAI211_X1 U21308 ( .C1(n18226), .C2(n18792), .A(n18286), .B(n18225), .ZN(
        n18248) );
  AOI21_X1 U21309 ( .B1(n18227), .B2(n18268), .A(n18248), .ZN(n18239) );
  AOI22_X1 U21310 ( .A1(n18231), .A2(n18230), .B1(n18229), .B2(n18228), .ZN(
        n18232) );
  OAI221_X1 U21311 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n18233), .C1(
        n10241), .C2(n18239), .A(n18232), .ZN(n18234) );
  AOI22_X1 U21312 ( .A1(n9802), .A2(n18234), .B1(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n18294), .ZN(n18236) );
  OAI211_X1 U21313 ( .C1(n18238), .C2(n18237), .A(n18236), .B(n18235), .ZN(
        P3_U2854) );
  AOI211_X1 U21314 ( .C1(n18241), .C2(n18240), .A(n18239), .B(n10081), .ZN(
        n18242) );
  AOI211_X1 U21315 ( .C1(n18294), .C2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18243), .B(n18242), .ZN(n18246) );
  NAND2_X1 U21316 ( .A1(n18315), .A2(n18244), .ZN(n18245) );
  OAI211_X1 U21317 ( .C1(n18247), .C2(n18311), .A(n18246), .B(n18245), .ZN(
        P3_U2855) );
  AOI21_X1 U21318 ( .B1(n9802), .B2(n18248), .A(n18294), .ZN(n18258) );
  OAI22_X1 U21319 ( .A1(n18258), .A2(n18251), .B1(n18312), .B2(n18874), .ZN(
        n18249) );
  AOI21_X1 U21320 ( .B1(n18315), .B2(n18250), .A(n18249), .ZN(n18254) );
  NAND4_X1 U21321 ( .A1(n18252), .A2(n9802), .A3(n18251), .A4(n18276), .ZN(
        n18253) );
  OAI211_X1 U21322 ( .C1(n18255), .C2(n18311), .A(n18254), .B(n18253), .ZN(
        P3_U2856) );
  NAND3_X1 U21323 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n9802), .A3(
        n18276), .ZN(n18270) );
  NOR2_X1 U21324 ( .A1(n18270), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18260) );
  OAI22_X1 U21325 ( .A1(n18258), .A2(n18257), .B1(n18311), .B2(n18256), .ZN(
        n18259) );
  AOI21_X1 U21326 ( .B1(n18260), .B2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n18259), .ZN(n18262) );
  OAI211_X1 U21327 ( .C1(n18263), .C2(n18304), .A(n18262), .B(n18261), .ZN(
        P3_U2857) );
  NAND2_X1 U21328 ( .A1(n18811), .A2(n18264), .ZN(n18289) );
  NAND3_X1 U21329 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18286), .A3(
        n18289), .ZN(n18265) );
  AOI21_X1 U21330 ( .B1(n18267), .B2(n18266), .A(n18265), .ZN(n18279) );
  NAND2_X1 U21331 ( .A1(n9802), .A2(n18268), .ZN(n18301) );
  OAI21_X1 U21332 ( .B1(n18279), .B2(n18301), .A(n18310), .ZN(n18272) );
  OAI22_X1 U21333 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18270), .B1(
        n18269), .B2(n18304), .ZN(n18271) );
  AOI21_X1 U21334 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18272), .A(
        n18271), .ZN(n18274) );
  NAND2_X1 U21335 ( .A1(n18308), .A2(P3_REIP_REG_4__SCAN_IN), .ZN(n18273) );
  OAI211_X1 U21336 ( .C1(n18311), .C2(n18275), .A(n18274), .B(n18273), .ZN(
        P3_U2858) );
  OAI21_X1 U21337 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18276), .A(
        n9802), .ZN(n18278) );
  OAI22_X1 U21338 ( .A1(n18279), .A2(n18278), .B1(n18304), .B2(n18277), .ZN(
        n18280) );
  AOI21_X1 U21339 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18294), .A(
        n18280), .ZN(n18282) );
  OAI211_X1 U21340 ( .C1(n18311), .C2(n18283), .A(n18282), .B(n18281), .ZN(
        P3_U2859) );
  AOI211_X1 U21341 ( .C1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n18286), .A(
        n18285), .B(n18284), .ZN(n18293) );
  INV_X1 U21342 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18952) );
  NOR3_X1 U21343 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18952), .A3(
        n18287), .ZN(n18292) );
  NAND4_X1 U21344 ( .A1(n18811), .A2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18288) );
  OAI211_X1 U21345 ( .C1(n18290), .C2(n18776), .A(n18289), .B(n18288), .ZN(
        n18291) );
  OR3_X1 U21346 ( .A1(n18293), .A2(n18292), .A3(n18291), .ZN(n18295) );
  AOI22_X1 U21347 ( .A1(n9802), .A2(n18295), .B1(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n18294), .ZN(n18297) );
  OAI211_X1 U21348 ( .C1(n18311), .C2(n18298), .A(n18297), .B(n18296), .ZN(
        P3_U2860) );
  NAND3_X1 U21349 ( .A1(n9802), .A2(n18300), .A3(n18299), .ZN(n18319) );
  NOR3_X1 U21350 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18302), .A3(
        n18301), .ZN(n18307) );
  OAI22_X1 U21351 ( .A1(n18305), .A2(n18304), .B1(n18311), .B2(n18303), .ZN(
        n18306) );
  AOI211_X1 U21352 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(n18308), .A(n18307), .B(
        n18306), .ZN(n18309) );
  OAI221_X1 U21353 ( .B1(n18952), .B2(n18310), .C1(n18952), .C2(n18319), .A(
        n18309), .ZN(P3_U2861) );
  INV_X1 U21354 ( .A(n18311), .ZN(n18317) );
  INV_X1 U21355 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n18980) );
  NOR2_X1 U21356 ( .A1(n18312), .A2(n18980), .ZN(n18313) );
  AOI221_X1 U21357 ( .B1(n18317), .B2(n18316), .C1(n18315), .C2(n18314), .A(
        n18313), .ZN(n18320) );
  OAI211_X1 U21358 ( .C1(n10081), .C2(n18791), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n18312), .ZN(n18318) );
  NAND3_X1 U21359 ( .A1(n18320), .A2(n18319), .A3(n18318), .ZN(P3_U2862) );
  AOI211_X1 U21360 ( .C1(n18322), .C2(n18321), .A(n18965), .B(n19005), .ZN(
        n18830) );
  OAI21_X1 U21361 ( .B1(n18830), .B2(n18370), .A(n18327), .ZN(n18323) );
  OAI221_X1 U21362 ( .B1(n18800), .B2(n18990), .C1(n18800), .C2(n18327), .A(
        n18323), .ZN(P3_U2863) );
  NOR2_X1 U21363 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18820), .ZN(
        n18583) );
  NOR2_X1 U21364 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18330), .ZN(
        n18513) );
  NOR2_X1 U21365 ( .A1(n18583), .A2(n18513), .ZN(n18325) );
  OAI22_X1 U21366 ( .A1(n18326), .A2(n18820), .B1(n18325), .B2(n18324), .ZN(
        P3_U2866) );
  NOR2_X1 U21367 ( .A1(n18328), .A2(n18327), .ZN(P3_U2867) );
  NAND2_X1 U21368 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18332) );
  NOR2_X1 U21369 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18332), .ZN(
        n18718) );
  NAND2_X1 U21370 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18718), .ZN(
        n18755) );
  NAND2_X1 U21371 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18719), .ZN(n18723) );
  NOR2_X2 U21372 ( .A1(n18486), .A2(n18329), .ZN(n18714) );
  NOR2_X1 U21373 ( .A1(n18820), .A2(n18511), .ZN(n18717) );
  INV_X1 U21374 ( .A(n18717), .ZN(n18712) );
  NOR2_X2 U21375 ( .A1(n18800), .A2(n18712), .ZN(n18767) );
  NOR2_X1 U21376 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18805) );
  NAND2_X1 U21377 ( .A1(n18330), .A2(n18820), .ZN(n18416) );
  INV_X1 U21378 ( .A(n18416), .ZN(n18415) );
  NAND2_X1 U21379 ( .A1(n18805), .A2(n18415), .ZN(n18437) );
  NOR2_X1 U21380 ( .A1(n18767), .A2(n18426), .ZN(n18392) );
  NOR2_X1 U21381 ( .A1(n18713), .A2(n18392), .ZN(n18364) );
  NOR2_X2 U21382 ( .A1(n18463), .A2(n19443), .ZN(n18715) );
  NAND2_X1 U21383 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18800), .ZN(
        n18331) );
  NOR2_X2 U21384 ( .A1(n18332), .A2(n18331), .ZN(n18707) );
  AOI22_X1 U21385 ( .A1(n18714), .A2(n18364), .B1(n18715), .B2(n18707), .ZN(
        n18338) );
  NOR2_X1 U21386 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18800), .ZN(
        n18557) );
  NOR2_X1 U21387 ( .A1(n18582), .A2(n18557), .ZN(n18629) );
  NOR2_X1 U21388 ( .A1(n18629), .A2(n18332), .ZN(n18680) );
  AOI21_X1 U21389 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n18486), .ZN(n18677) );
  INV_X1 U21390 ( .A(n18392), .ZN(n18333) );
  AOI22_X1 U21391 ( .A1(n18719), .A2(n18680), .B1(n18677), .B2(n18333), .ZN(
        n18367) );
  NAND2_X1 U21392 ( .A1(n18335), .A2(n18334), .ZN(n18365) );
  NOR2_X1 U21393 ( .A1(n18336), .A2(n18365), .ZN(n18720) );
  AOI22_X1 U21394 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18367), .B1(
        n18426), .B2(n18720), .ZN(n18337) );
  OAI211_X1 U21395 ( .C1(n18755), .C2(n18723), .A(n18338), .B(n18337), .ZN(
        P3_U2868) );
  NAND2_X1 U21396 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18719), .ZN(n18688) );
  NOR2_X2 U21397 ( .A1(n18463), .A2(n19449), .ZN(n18685) );
  AOI22_X1 U21398 ( .A1(n18364), .A2(n18724), .B1(n18707), .B2(n18685), .ZN(
        n18341) );
  NOR2_X2 U21399 ( .A1(n18339), .A2(n18365), .ZN(n18726) );
  AOI22_X1 U21400 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18367), .B1(
        n18426), .B2(n18726), .ZN(n18340) );
  OAI211_X1 U21401 ( .C1(n18755), .C2(n18688), .A(n18341), .B(n18340), .ZN(
        P3_U2869) );
  INV_X1 U21402 ( .A(n18707), .ZN(n18683) );
  NAND2_X1 U21403 ( .A1(n18719), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18735) );
  INV_X1 U21404 ( .A(n18755), .ZN(n18765) );
  NAND2_X1 U21405 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18719), .ZN(n18567) );
  INV_X1 U21406 ( .A(n18567), .ZN(n18731) );
  NOR2_X2 U21407 ( .A1(n18486), .A2(n18342), .ZN(n18730) );
  AOI22_X1 U21408 ( .A1(n18765), .A2(n18731), .B1(n18364), .B2(n18730), .ZN(
        n18345) );
  NOR2_X2 U21409 ( .A1(n18343), .A2(n18365), .ZN(n18732) );
  AOI22_X1 U21410 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18367), .B1(
        n18426), .B2(n18732), .ZN(n18344) );
  OAI211_X1 U21411 ( .C1(n18683), .C2(n18735), .A(n18345), .B(n18344), .ZN(
        P3_U2870) );
  NAND2_X1 U21412 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18719), .ZN(n18741) );
  NOR2_X2 U21413 ( .A1(n18486), .A2(n18346), .ZN(n18736) );
  NAND2_X1 U21414 ( .A1(n18719), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18694) );
  INV_X1 U21415 ( .A(n18694), .ZN(n18737) );
  AOI22_X1 U21416 ( .A1(n18364), .A2(n18736), .B1(n18707), .B2(n18737), .ZN(
        n18349) );
  AOI22_X1 U21417 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18367), .B1(
        n18426), .B2(n18738), .ZN(n18348) );
  OAI211_X1 U21418 ( .C1(n18755), .C2(n18741), .A(n18349), .B(n18348), .ZN(
        P3_U2871) );
  NAND2_X1 U21419 ( .A1(n18719), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18747) );
  NOR2_X2 U21420 ( .A1(n18486), .A2(n18350), .ZN(n18742) );
  AOI22_X1 U21421 ( .A1(n18765), .A2(n18743), .B1(n18364), .B2(n18742), .ZN(
        n18353) );
  NOR2_X2 U21422 ( .A1(n18351), .A2(n18365), .ZN(n18744) );
  AOI22_X1 U21423 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18367), .B1(
        n18426), .B2(n18744), .ZN(n18352) );
  OAI211_X1 U21424 ( .C1(n18683), .C2(n18747), .A(n18353), .B(n18352), .ZN(
        P3_U2872) );
  NAND2_X1 U21425 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18719), .ZN(n18700) );
  NOR2_X2 U21426 ( .A1(n18486), .A2(n18354), .ZN(n18748) );
  NOR2_X1 U21427 ( .A1(n18463), .A2(n15083), .ZN(n18697) );
  AOI22_X1 U21428 ( .A1(n18364), .A2(n18748), .B1(n18707), .B2(n18697), .ZN(
        n18357) );
  NOR2_X2 U21429 ( .A1(n18355), .A2(n18365), .ZN(n18751) );
  AOI22_X1 U21430 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18367), .B1(
        n18426), .B2(n18751), .ZN(n18356) );
  OAI211_X1 U21431 ( .C1(n18755), .C2(n18700), .A(n18357), .B(n18356), .ZN(
        P3_U2873) );
  NAND2_X1 U21432 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18719), .ZN(n18761) );
  NOR2_X2 U21433 ( .A1(n18358), .A2(n18486), .ZN(n18756) );
  NOR2_X1 U21434 ( .A1(n18359), .A2(n18463), .ZN(n18757) );
  AOI22_X1 U21435 ( .A1(n18364), .A2(n18756), .B1(n18707), .B2(n18757), .ZN(
        n18362) );
  NOR2_X2 U21436 ( .A1(n18360), .A2(n18365), .ZN(n18758) );
  AOI22_X1 U21437 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18367), .B1(
        n18426), .B2(n18758), .ZN(n18361) );
  OAI211_X1 U21438 ( .C1(n18755), .C2(n18761), .A(n18362), .B(n18361), .ZN(
        P3_U2874) );
  NAND2_X1 U21439 ( .A1(n18719), .A2(BUF2_REG_31__SCAN_IN), .ZN(n18772) );
  NOR2_X2 U21440 ( .A1(n18363), .A2(n18486), .ZN(n18763) );
  NAND2_X1 U21441 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18719), .ZN(n18675) );
  INV_X1 U21442 ( .A(n18675), .ZN(n18764) );
  AOI22_X1 U21443 ( .A1(n18364), .A2(n18763), .B1(n18707), .B2(n18764), .ZN(
        n18369) );
  NOR2_X2 U21444 ( .A1(n18366), .A2(n18365), .ZN(n18766) );
  AOI22_X1 U21445 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18367), .B1(
        n18426), .B2(n18766), .ZN(n18368) );
  OAI211_X1 U21446 ( .C1(n18755), .C2(n18772), .A(n18369), .B(n18368), .ZN(
        P3_U2875) );
  NOR2_X1 U21447 ( .A1(n18370), .A2(n18486), .ZN(n18716) );
  NAND2_X1 U21448 ( .A1(n18716), .A2(n18801), .ZN(n18460) );
  OAI22_X1 U21449 ( .A1(n18463), .A2(n18712), .B1(n18416), .B2(n18460), .ZN(
        n18386) );
  INV_X1 U21450 ( .A(n18723), .ZN(n18676) );
  INV_X1 U21451 ( .A(n18713), .ZN(n18837) );
  NAND2_X1 U21452 ( .A1(n18801), .A2(n18837), .ZN(n18558) );
  NOR2_X1 U21453 ( .A1(n18416), .A2(n18558), .ZN(n18388) );
  AOI22_X1 U21454 ( .A1(n18676), .A2(n18707), .B1(n18714), .B2(n18388), .ZN(
        n18372) );
  NAND2_X1 U21455 ( .A1(n18415), .A2(n18557), .ZN(n18459) );
  INV_X1 U21456 ( .A(n18459), .ZN(n18452) );
  AOI22_X1 U21457 ( .A1(n18767), .A2(n18715), .B1(n18720), .B2(n18452), .ZN(
        n18371) );
  OAI211_X1 U21458 ( .C1(n18373), .C2(n18386), .A(n18372), .B(n18371), .ZN(
        P3_U2876) );
  AOI22_X1 U21459 ( .A1(n18767), .A2(n18685), .B1(n18724), .B2(n18388), .ZN(
        n18375) );
  INV_X1 U21460 ( .A(n18386), .ZN(n18389) );
  AOI22_X1 U21461 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18389), .B1(
        n18726), .B2(n18452), .ZN(n18374) );
  OAI211_X1 U21462 ( .C1(n18683), .C2(n18688), .A(n18375), .B(n18374), .ZN(
        P3_U2877) );
  INV_X1 U21463 ( .A(n18767), .ZN(n18414) );
  AOI22_X1 U21464 ( .A1(n18707), .A2(n18731), .B1(n18730), .B2(n18388), .ZN(
        n18377) );
  AOI22_X1 U21465 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18389), .B1(
        n18732), .B2(n18452), .ZN(n18376) );
  OAI211_X1 U21466 ( .C1(n18414), .C2(n18735), .A(n18377), .B(n18376), .ZN(
        P3_U2878) );
  AOI22_X1 U21467 ( .A1(n18767), .A2(n18737), .B1(n18736), .B2(n18388), .ZN(
        n18379) );
  AOI22_X1 U21468 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18389), .B1(
        n18738), .B2(n18452), .ZN(n18378) );
  OAI211_X1 U21469 ( .C1(n18683), .C2(n18741), .A(n18379), .B(n18378), .ZN(
        P3_U2879) );
  INV_X1 U21470 ( .A(n18743), .ZN(n18642) );
  INV_X1 U21471 ( .A(n18747), .ZN(n18639) );
  AOI22_X1 U21472 ( .A1(n18767), .A2(n18639), .B1(n18742), .B2(n18388), .ZN(
        n18381) );
  AOI22_X1 U21473 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18389), .B1(
        n18744), .B2(n18452), .ZN(n18380) );
  OAI211_X1 U21474 ( .C1(n18683), .C2(n18642), .A(n18381), .B(n18380), .ZN(
        P3_U2880) );
  INV_X1 U21475 ( .A(n18697), .ZN(n18754) );
  INV_X1 U21476 ( .A(n18700), .ZN(n18750) );
  AOI22_X1 U21477 ( .A1(n18707), .A2(n18750), .B1(n18748), .B2(n18388), .ZN(
        n18383) );
  AOI22_X1 U21478 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18389), .B1(
        n18751), .B2(n18452), .ZN(n18382) );
  OAI211_X1 U21479 ( .C1(n18414), .C2(n18754), .A(n18383), .B(n18382), .ZN(
        P3_U2881) );
  INV_X1 U21480 ( .A(n18761), .ZN(n18702) );
  AOI22_X1 U21481 ( .A1(n18707), .A2(n18702), .B1(n18756), .B2(n18388), .ZN(
        n18385) );
  AOI22_X1 U21482 ( .A1(n18767), .A2(n18757), .B1(n18758), .B2(n18452), .ZN(
        n18384) );
  OAI211_X1 U21483 ( .C1(n18387), .C2(n18386), .A(n18385), .B(n18384), .ZN(
        P3_U2882) );
  AOI22_X1 U21484 ( .A1(n18767), .A2(n18764), .B1(n18763), .B2(n18388), .ZN(
        n18391) );
  AOI22_X1 U21485 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18389), .B1(
        n18766), .B2(n18452), .ZN(n18390) );
  OAI211_X1 U21486 ( .C1(n18683), .C2(n18772), .A(n18391), .B(n18390), .ZN(
        P3_U2883) );
  NAND2_X1 U21487 ( .A1(n18415), .A2(n18582), .ZN(n18484) );
  NOR2_X1 U21488 ( .A1(n18452), .A2(n18473), .ZN(n18438) );
  OAI21_X1 U21489 ( .B1(n18627), .B2(n18392), .A(n18438), .ZN(n18393) );
  OAI211_X1 U21490 ( .C1(n18942), .C2(n18473), .A(n18393), .B(n18536), .ZN(
        n18411) );
  INV_X1 U21491 ( .A(n18411), .ZN(n18397) );
  NOR2_X1 U21492 ( .A1(n18713), .A2(n18438), .ZN(n18410) );
  AOI22_X1 U21493 ( .A1(n18676), .A2(n18767), .B1(n18714), .B2(n18410), .ZN(
        n18395) );
  AOI22_X1 U21494 ( .A1(n18426), .A2(n18715), .B1(n18720), .B2(n18473), .ZN(
        n18394) );
  OAI211_X1 U21495 ( .C1(n18397), .C2(n18396), .A(n18395), .B(n18394), .ZN(
        P3_U2884) );
  AOI22_X1 U21496 ( .A1(n18426), .A2(n18685), .B1(n18724), .B2(n18410), .ZN(
        n18399) );
  AOI22_X1 U21497 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18411), .B1(
        n18726), .B2(n18473), .ZN(n18398) );
  OAI211_X1 U21498 ( .C1(n18414), .C2(n18688), .A(n18399), .B(n18398), .ZN(
        P3_U2885) );
  INV_X1 U21499 ( .A(n18735), .ZN(n18564) );
  AOI22_X1 U21500 ( .A1(n18426), .A2(n18564), .B1(n18730), .B2(n18410), .ZN(
        n18401) );
  AOI22_X1 U21501 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18411), .B1(
        n18732), .B2(n18473), .ZN(n18400) );
  OAI211_X1 U21502 ( .C1(n18414), .C2(n18567), .A(n18401), .B(n18400), .ZN(
        P3_U2886) );
  AOI22_X1 U21503 ( .A1(n18426), .A2(n18737), .B1(n18736), .B2(n18410), .ZN(
        n18403) );
  AOI22_X1 U21504 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18411), .B1(
        n18738), .B2(n18473), .ZN(n18402) );
  OAI211_X1 U21505 ( .C1(n18414), .C2(n18741), .A(n18403), .B(n18402), .ZN(
        P3_U2887) );
  AOI22_X1 U21506 ( .A1(n18767), .A2(n18743), .B1(n18742), .B2(n18410), .ZN(
        n18405) );
  AOI22_X1 U21507 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18411), .B1(
        n18744), .B2(n18473), .ZN(n18404) );
  OAI211_X1 U21508 ( .C1(n18437), .C2(n18747), .A(n18405), .B(n18404), .ZN(
        P3_U2888) );
  AOI22_X1 U21509 ( .A1(n18426), .A2(n18697), .B1(n18748), .B2(n18410), .ZN(
        n18407) );
  AOI22_X1 U21510 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18411), .B1(
        n18751), .B2(n18473), .ZN(n18406) );
  OAI211_X1 U21511 ( .C1(n18414), .C2(n18700), .A(n18407), .B(n18406), .ZN(
        P3_U2889) );
  INV_X1 U21512 ( .A(n18757), .ZN(n18705) );
  AOI22_X1 U21513 ( .A1(n18767), .A2(n18702), .B1(n18756), .B2(n18410), .ZN(
        n18409) );
  AOI22_X1 U21514 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18411), .B1(
        n18758), .B2(n18473), .ZN(n18408) );
  OAI211_X1 U21515 ( .C1(n18437), .C2(n18705), .A(n18409), .B(n18408), .ZN(
        P3_U2890) );
  AOI22_X1 U21516 ( .A1(n18426), .A2(n18764), .B1(n18763), .B2(n18410), .ZN(
        n18413) );
  AOI22_X1 U21517 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18411), .B1(
        n18766), .B2(n18473), .ZN(n18412) );
  OAI211_X1 U21518 ( .C1(n18414), .C2(n18772), .A(n18413), .B(n18412), .ZN(
        P3_U2891) );
  NAND2_X1 U21519 ( .A1(n18801), .A2(n18627), .ZN(n18512) );
  NAND2_X1 U21520 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18415), .ZN(
        n18462) );
  NOR2_X2 U21521 ( .A1(n18800), .A2(n18462), .ZN(n18507) );
  OAI21_X1 U21522 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18416), .A(n18505), 
        .ZN(n18417) );
  NAND3_X1 U21523 ( .A1(n18536), .A2(n18512), .A3(n18417), .ZN(n18434) );
  NOR2_X1 U21524 ( .A1(n18713), .A2(n18462), .ZN(n18433) );
  AOI22_X1 U21525 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18434), .B1(
        n18714), .B2(n18433), .ZN(n18419) );
  AOI22_X1 U21526 ( .A1(n18720), .A2(n18507), .B1(n18715), .B2(n18452), .ZN(
        n18418) );
  OAI211_X1 U21527 ( .C1(n18723), .C2(n18437), .A(n18419), .B(n18418), .ZN(
        P3_U2892) );
  INV_X1 U21528 ( .A(n18685), .ZN(n18729) );
  INV_X1 U21529 ( .A(n18688), .ZN(n18725) );
  AOI22_X1 U21530 ( .A1(n18426), .A2(n18725), .B1(n18724), .B2(n18433), .ZN(
        n18421) );
  AOI22_X1 U21531 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18434), .B1(
        n18726), .B2(n18507), .ZN(n18420) );
  OAI211_X1 U21532 ( .C1(n18729), .C2(n18459), .A(n18421), .B(n18420), .ZN(
        P3_U2893) );
  AOI22_X1 U21533 ( .A1(n18426), .A2(n18731), .B1(n18730), .B2(n18433), .ZN(
        n18423) );
  AOI22_X1 U21534 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18434), .B1(
        n18732), .B2(n18507), .ZN(n18422) );
  OAI211_X1 U21535 ( .C1(n18735), .C2(n18459), .A(n18423), .B(n18422), .ZN(
        P3_U2894) );
  AOI22_X1 U21536 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18434), .B1(
        n18736), .B2(n18433), .ZN(n18425) );
  AOI22_X1 U21537 ( .A1(n18738), .A2(n18507), .B1(n18737), .B2(n18452), .ZN(
        n18424) );
  OAI211_X1 U21538 ( .C1(n18437), .C2(n18741), .A(n18425), .B(n18424), .ZN(
        P3_U2895) );
  AOI22_X1 U21539 ( .A1(n18426), .A2(n18743), .B1(n18742), .B2(n18433), .ZN(
        n18428) );
  AOI22_X1 U21540 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18434), .B1(
        n18744), .B2(n18507), .ZN(n18427) );
  OAI211_X1 U21541 ( .C1(n18747), .C2(n18459), .A(n18428), .B(n18427), .ZN(
        P3_U2896) );
  AOI22_X1 U21542 ( .A1(n18697), .A2(n18452), .B1(n18748), .B2(n18433), .ZN(
        n18430) );
  AOI22_X1 U21543 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18434), .B1(
        n18751), .B2(n18507), .ZN(n18429) );
  OAI211_X1 U21544 ( .C1(n18437), .C2(n18700), .A(n18430), .B(n18429), .ZN(
        P3_U2897) );
  AOI22_X1 U21545 ( .A1(n18757), .A2(n18452), .B1(n18756), .B2(n18433), .ZN(
        n18432) );
  AOI22_X1 U21546 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18434), .B1(
        n18758), .B2(n18507), .ZN(n18431) );
  OAI211_X1 U21547 ( .C1(n18437), .C2(n18761), .A(n18432), .B(n18431), .ZN(
        P3_U2898) );
  AOI22_X1 U21548 ( .A1(n18764), .A2(n18452), .B1(n18763), .B2(n18433), .ZN(
        n18436) );
  AOI22_X1 U21549 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18434), .B1(
        n18766), .B2(n18507), .ZN(n18435) );
  OAI211_X1 U21550 ( .C1(n18437), .C2(n18772), .A(n18436), .B(n18435), .ZN(
        P3_U2899) );
  NAND2_X1 U21551 ( .A1(n18805), .A2(n18513), .ZN(n18533) );
  AOI21_X1 U21552 ( .B1(n18505), .B2(n18533), .A(n18713), .ZN(n18455) );
  AOI22_X1 U21553 ( .A1(n18676), .A2(n18452), .B1(n18714), .B2(n18455), .ZN(
        n18441) );
  AOI221_X1 U21554 ( .B1(n18438), .B2(n18505), .C1(n18627), .C2(n18505), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18439) );
  OAI21_X1 U21555 ( .B1(n18526), .B2(n18439), .A(n18536), .ZN(n18456) );
  AOI22_X1 U21556 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18456), .B1(
        n18715), .B2(n18473), .ZN(n18440) );
  OAI211_X1 U21557 ( .C1(n18684), .C2(n18533), .A(n18441), .B(n18440), .ZN(
        P3_U2900) );
  AOI22_X1 U21558 ( .A1(n18685), .A2(n18473), .B1(n18724), .B2(n18455), .ZN(
        n18443) );
  AOI22_X1 U21559 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18456), .B1(
        n18726), .B2(n18526), .ZN(n18442) );
  OAI211_X1 U21560 ( .C1(n18688), .C2(n18459), .A(n18443), .B(n18442), .ZN(
        P3_U2901) );
  AOI22_X1 U21561 ( .A1(n18731), .A2(n18452), .B1(n18730), .B2(n18455), .ZN(
        n18445) );
  AOI22_X1 U21562 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18456), .B1(
        n18732), .B2(n18526), .ZN(n18444) );
  OAI211_X1 U21563 ( .C1(n18735), .C2(n18484), .A(n18445), .B(n18444), .ZN(
        P3_U2902) );
  AOI22_X1 U21564 ( .A1(n18737), .A2(n18473), .B1(n18736), .B2(n18455), .ZN(
        n18447) );
  AOI22_X1 U21565 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18456), .B1(
        n18738), .B2(n18526), .ZN(n18446) );
  OAI211_X1 U21566 ( .C1(n18741), .C2(n18459), .A(n18447), .B(n18446), .ZN(
        P3_U2903) );
  AOI22_X1 U21567 ( .A1(n18743), .A2(n18452), .B1(n18742), .B2(n18455), .ZN(
        n18449) );
  AOI22_X1 U21568 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18456), .B1(
        n18744), .B2(n18526), .ZN(n18448) );
  OAI211_X1 U21569 ( .C1(n18747), .C2(n18484), .A(n18449), .B(n18448), .ZN(
        P3_U2904) );
  AOI22_X1 U21570 ( .A1(n18750), .A2(n18452), .B1(n18748), .B2(n18455), .ZN(
        n18451) );
  AOI22_X1 U21571 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18456), .B1(
        n18751), .B2(n18526), .ZN(n18450) );
  OAI211_X1 U21572 ( .C1(n18754), .C2(n18484), .A(n18451), .B(n18450), .ZN(
        P3_U2905) );
  AOI22_X1 U21573 ( .A1(n18702), .A2(n18452), .B1(n18756), .B2(n18455), .ZN(
        n18454) );
  AOI22_X1 U21574 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18456), .B1(
        n18758), .B2(n18526), .ZN(n18453) );
  OAI211_X1 U21575 ( .C1(n18705), .C2(n18484), .A(n18454), .B(n18453), .ZN(
        P3_U2906) );
  AOI22_X1 U21576 ( .A1(n18764), .A2(n18473), .B1(n18763), .B2(n18455), .ZN(
        n18458) );
  AOI22_X1 U21577 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18456), .B1(
        n18766), .B2(n18526), .ZN(n18457) );
  OAI211_X1 U21578 ( .C1(n18772), .C2(n18459), .A(n18458), .B(n18457), .ZN(
        P3_U2907) );
  NAND2_X1 U21579 ( .A1(n18513), .A2(n18557), .ZN(n18549) );
  INV_X1 U21580 ( .A(n18513), .ZN(n18461) );
  NOR2_X1 U21581 ( .A1(n18461), .A2(n18558), .ZN(n18480) );
  AOI22_X1 U21582 ( .A1(n18714), .A2(n18480), .B1(n18715), .B2(n18507), .ZN(
        n18466) );
  OAI22_X1 U21583 ( .A1(n18463), .A2(n18462), .B1(n18461), .B2(n18460), .ZN(
        n18464) );
  INV_X1 U21584 ( .A(n18464), .ZN(n18481) );
  AOI22_X1 U21585 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18481), .B1(
        n18676), .B2(n18473), .ZN(n18465) );
  OAI211_X1 U21586 ( .C1(n18684), .C2(n18549), .A(n18466), .B(n18465), .ZN(
        P3_U2908) );
  AOI22_X1 U21587 ( .A1(n18685), .A2(n18507), .B1(n18724), .B2(n18480), .ZN(
        n18468) );
  AOI22_X1 U21588 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18481), .B1(
        n18726), .B2(n18553), .ZN(n18467) );
  OAI211_X1 U21589 ( .C1(n18688), .C2(n18484), .A(n18468), .B(n18467), .ZN(
        P3_U2909) );
  AOI22_X1 U21590 ( .A1(n18731), .A2(n18473), .B1(n18730), .B2(n18480), .ZN(
        n18470) );
  AOI22_X1 U21591 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18481), .B1(
        n18732), .B2(n18553), .ZN(n18469) );
  OAI211_X1 U21592 ( .C1(n18735), .C2(n18505), .A(n18470), .B(n18469), .ZN(
        P3_U2910) );
  AOI22_X1 U21593 ( .A1(n18737), .A2(n18507), .B1(n18736), .B2(n18480), .ZN(
        n18472) );
  AOI22_X1 U21594 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18481), .B1(
        n18738), .B2(n18553), .ZN(n18471) );
  OAI211_X1 U21595 ( .C1(n18741), .C2(n18484), .A(n18472), .B(n18471), .ZN(
        P3_U2911) );
  AOI22_X1 U21596 ( .A1(n18743), .A2(n18473), .B1(n18742), .B2(n18480), .ZN(
        n18475) );
  AOI22_X1 U21597 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18481), .B1(
        n18744), .B2(n18553), .ZN(n18474) );
  OAI211_X1 U21598 ( .C1(n18747), .C2(n18505), .A(n18475), .B(n18474), .ZN(
        P3_U2912) );
  AOI22_X1 U21599 ( .A1(n18697), .A2(n18507), .B1(n18748), .B2(n18480), .ZN(
        n18477) );
  AOI22_X1 U21600 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18481), .B1(
        n18751), .B2(n18553), .ZN(n18476) );
  OAI211_X1 U21601 ( .C1(n18700), .C2(n18484), .A(n18477), .B(n18476), .ZN(
        P3_U2913) );
  AOI22_X1 U21602 ( .A1(n18757), .A2(n18507), .B1(n18756), .B2(n18480), .ZN(
        n18479) );
  AOI22_X1 U21603 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18481), .B1(
        n18758), .B2(n18553), .ZN(n18478) );
  OAI211_X1 U21604 ( .C1(n18761), .C2(n18484), .A(n18479), .B(n18478), .ZN(
        P3_U2914) );
  AOI22_X1 U21605 ( .A1(n18764), .A2(n18507), .B1(n18763), .B2(n18480), .ZN(
        n18483) );
  AOI22_X1 U21606 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18481), .B1(
        n18766), .B2(n18553), .ZN(n18482) );
  OAI211_X1 U21607 ( .C1(n18772), .C2(n18484), .A(n18483), .B(n18482), .ZN(
        P3_U2915) );
  NAND2_X1 U21608 ( .A1(n18513), .A2(n18582), .ZN(n18581) );
  NAND2_X1 U21609 ( .A1(n18505), .A2(n18533), .ZN(n18485) );
  NAND2_X1 U21610 ( .A1(n18549), .A2(n18581), .ZN(n18488) );
  AOI21_X1 U21611 ( .B1(n18679), .B2(n18485), .A(n18488), .ZN(n18487) );
  AOI211_X1 U21612 ( .C1(P3_STATE2_REG_3__SCAN_IN), .C2(n18581), .A(n18487), 
        .B(n18486), .ZN(n18492) );
  INV_X1 U21613 ( .A(n18488), .ZN(n18534) );
  NOR2_X1 U21614 ( .A1(n18713), .A2(n18534), .ZN(n18506) );
  AOI22_X1 U21615 ( .A1(n18714), .A2(n18506), .B1(n18715), .B2(n18526), .ZN(
        n18490) );
  INV_X1 U21616 ( .A(n18581), .ZN(n18572) );
  AOI22_X1 U21617 ( .A1(n18676), .A2(n18507), .B1(n18720), .B2(n18572), .ZN(
        n18489) );
  OAI211_X1 U21618 ( .C1(n18492), .C2(n18491), .A(n18490), .B(n18489), .ZN(
        P3_U2916) );
  AOI22_X1 U21619 ( .A1(n18685), .A2(n18526), .B1(n18724), .B2(n18506), .ZN(
        n18494) );
  INV_X1 U21620 ( .A(n18492), .ZN(n18508) );
  AOI22_X1 U21621 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18508), .B1(
        n18726), .B2(n18572), .ZN(n18493) );
  OAI211_X1 U21622 ( .C1(n18688), .C2(n18505), .A(n18494), .B(n18493), .ZN(
        P3_U2917) );
  AOI22_X1 U21623 ( .A1(n18731), .A2(n18507), .B1(n18730), .B2(n18506), .ZN(
        n18496) );
  AOI22_X1 U21624 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18508), .B1(
        n18732), .B2(n18572), .ZN(n18495) );
  OAI211_X1 U21625 ( .C1(n18735), .C2(n18533), .A(n18496), .B(n18495), .ZN(
        P3_U2918) );
  AOI22_X1 U21626 ( .A1(n18737), .A2(n18526), .B1(n18736), .B2(n18506), .ZN(
        n18498) );
  AOI22_X1 U21627 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18508), .B1(
        n18738), .B2(n18572), .ZN(n18497) );
  OAI211_X1 U21628 ( .C1(n18741), .C2(n18505), .A(n18498), .B(n18497), .ZN(
        P3_U2919) );
  AOI22_X1 U21629 ( .A1(n18639), .A2(n18526), .B1(n18742), .B2(n18506), .ZN(
        n18500) );
  AOI22_X1 U21630 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18508), .B1(
        n18744), .B2(n18572), .ZN(n18499) );
  OAI211_X1 U21631 ( .C1(n18642), .C2(n18505), .A(n18500), .B(n18499), .ZN(
        P3_U2920) );
  AOI22_X1 U21632 ( .A1(n18697), .A2(n18526), .B1(n18748), .B2(n18506), .ZN(
        n18502) );
  AOI22_X1 U21633 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18508), .B1(
        n18751), .B2(n18572), .ZN(n18501) );
  OAI211_X1 U21634 ( .C1(n18700), .C2(n18505), .A(n18502), .B(n18501), .ZN(
        P3_U2921) );
  AOI22_X1 U21635 ( .A1(n18757), .A2(n18526), .B1(n18756), .B2(n18506), .ZN(
        n18504) );
  AOI22_X1 U21636 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18508), .B1(
        n18758), .B2(n18572), .ZN(n18503) );
  OAI211_X1 U21637 ( .C1(n18761), .C2(n18505), .A(n18504), .B(n18503), .ZN(
        P3_U2922) );
  INV_X1 U21638 ( .A(n18772), .ZN(n18671) );
  AOI22_X1 U21639 ( .A1(n18671), .A2(n18507), .B1(n18763), .B2(n18506), .ZN(
        n18510) );
  AOI22_X1 U21640 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18508), .B1(
        n18766), .B2(n18572), .ZN(n18509) );
  OAI211_X1 U21641 ( .C1(n18675), .C2(n18533), .A(n18510), .B(n18509), .ZN(
        P3_U2923) );
  NOR2_X1 U21642 ( .A1(n18511), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18559) );
  AND2_X1 U21643 ( .A1(n18837), .A2(n18559), .ZN(n18529) );
  AOI22_X1 U21644 ( .A1(n18714), .A2(n18529), .B1(n18715), .B2(n18553), .ZN(
        n18515) );
  NAND3_X1 U21645 ( .A1(n18513), .A2(n18716), .A3(n18512), .ZN(n18530) );
  NAND2_X1 U21646 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18559), .ZN(
        n18600) );
  AOI22_X1 U21647 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18530), .B1(
        n18720), .B2(n18602), .ZN(n18514) );
  OAI211_X1 U21648 ( .C1(n18723), .C2(n18533), .A(n18515), .B(n18514), .ZN(
        P3_U2924) );
  AOI22_X1 U21649 ( .A1(n18725), .A2(n18526), .B1(n18724), .B2(n18529), .ZN(
        n18517) );
  AOI22_X1 U21650 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18530), .B1(
        n18726), .B2(n18602), .ZN(n18516) );
  OAI211_X1 U21651 ( .C1(n18729), .C2(n18549), .A(n18517), .B(n18516), .ZN(
        P3_U2925) );
  AOI22_X1 U21652 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18530), .B1(
        n18730), .B2(n18529), .ZN(n18519) );
  AOI22_X1 U21653 ( .A1(n18732), .A2(n18602), .B1(n18731), .B2(n18526), .ZN(
        n18518) );
  OAI211_X1 U21654 ( .C1(n18735), .C2(n18549), .A(n18519), .B(n18518), .ZN(
        P3_U2926) );
  AOI22_X1 U21655 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18530), .B1(
        n18736), .B2(n18529), .ZN(n18521) );
  AOI22_X1 U21656 ( .A1(n18738), .A2(n18602), .B1(n18737), .B2(n18553), .ZN(
        n18520) );
  OAI211_X1 U21657 ( .C1(n18741), .C2(n18533), .A(n18521), .B(n18520), .ZN(
        P3_U2927) );
  AOI22_X1 U21658 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18530), .B1(
        n18742), .B2(n18529), .ZN(n18523) );
  AOI22_X1 U21659 ( .A1(n18744), .A2(n18602), .B1(n18743), .B2(n18526), .ZN(
        n18522) );
  OAI211_X1 U21660 ( .C1(n18747), .C2(n18549), .A(n18523), .B(n18522), .ZN(
        P3_U2928) );
  AOI22_X1 U21661 ( .A1(n18697), .A2(n18553), .B1(n18748), .B2(n18529), .ZN(
        n18525) );
  AOI22_X1 U21662 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18530), .B1(
        n18751), .B2(n18602), .ZN(n18524) );
  OAI211_X1 U21663 ( .C1(n18700), .C2(n18533), .A(n18525), .B(n18524), .ZN(
        P3_U2929) );
  AOI22_X1 U21664 ( .A1(n18702), .A2(n18526), .B1(n18756), .B2(n18529), .ZN(
        n18528) );
  AOI22_X1 U21665 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18530), .B1(
        n18758), .B2(n18602), .ZN(n18527) );
  OAI211_X1 U21666 ( .C1(n18705), .C2(n18549), .A(n18528), .B(n18527), .ZN(
        P3_U2930) );
  AOI22_X1 U21667 ( .A1(n18764), .A2(n18553), .B1(n18763), .B2(n18529), .ZN(
        n18532) );
  AOI22_X1 U21668 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18530), .B1(
        n18766), .B2(n18602), .ZN(n18531) );
  OAI211_X1 U21669 ( .C1(n18772), .C2(n18533), .A(n18532), .B(n18531), .ZN(
        P3_U2931) );
  NAND2_X1 U21670 ( .A1(n18805), .A2(n18583), .ZN(n18626) );
  NOR2_X1 U21671 ( .A1(n18602), .A2(n18619), .ZN(n18584) );
  NOR2_X1 U21672 ( .A1(n18713), .A2(n18584), .ZN(n18552) );
  AOI22_X1 U21673 ( .A1(n18676), .A2(n18553), .B1(n18714), .B2(n18552), .ZN(
        n18538) );
  OAI21_X1 U21674 ( .B1(n18534), .B2(n18627), .A(n18584), .ZN(n18535) );
  OAI211_X1 U21675 ( .C1(n18619), .C2(n18942), .A(n18536), .B(n18535), .ZN(
        n18554) );
  AOI22_X1 U21676 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18554), .B1(
        n18715), .B2(n18572), .ZN(n18537) );
  OAI211_X1 U21677 ( .C1(n18684), .C2(n18626), .A(n18538), .B(n18537), .ZN(
        P3_U2932) );
  AOI22_X1 U21678 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18554), .B1(
        n18724), .B2(n18552), .ZN(n18540) );
  AOI22_X1 U21679 ( .A1(n18726), .A2(n18619), .B1(n18685), .B2(n18572), .ZN(
        n18539) );
  OAI211_X1 U21680 ( .C1(n18688), .C2(n18549), .A(n18540), .B(n18539), .ZN(
        P3_U2933) );
  AOI22_X1 U21681 ( .A1(n18564), .A2(n18572), .B1(n18730), .B2(n18552), .ZN(
        n18542) );
  AOI22_X1 U21682 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18554), .B1(
        n18732), .B2(n18619), .ZN(n18541) );
  OAI211_X1 U21683 ( .C1(n18567), .C2(n18549), .A(n18542), .B(n18541), .ZN(
        P3_U2934) );
  INV_X1 U21684 ( .A(n18741), .ZN(n18691) );
  AOI22_X1 U21685 ( .A1(n18691), .A2(n18553), .B1(n18736), .B2(n18552), .ZN(
        n18544) );
  AOI22_X1 U21686 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18554), .B1(
        n18738), .B2(n18619), .ZN(n18543) );
  OAI211_X1 U21687 ( .C1(n18694), .C2(n18581), .A(n18544), .B(n18543), .ZN(
        P3_U2935) );
  AOI22_X1 U21688 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18554), .B1(
        n18742), .B2(n18552), .ZN(n18546) );
  AOI22_X1 U21689 ( .A1(n18639), .A2(n18572), .B1(n18744), .B2(n18619), .ZN(
        n18545) );
  OAI211_X1 U21690 ( .C1(n18642), .C2(n18549), .A(n18546), .B(n18545), .ZN(
        P3_U2936) );
  AOI22_X1 U21691 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18554), .B1(
        n18748), .B2(n18552), .ZN(n18548) );
  AOI22_X1 U21692 ( .A1(n18751), .A2(n18619), .B1(n18697), .B2(n18572), .ZN(
        n18547) );
  OAI211_X1 U21693 ( .C1(n18700), .C2(n18549), .A(n18548), .B(n18547), .ZN(
        P3_U2937) );
  AOI22_X1 U21694 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18554), .B1(
        n18756), .B2(n18552), .ZN(n18551) );
  AOI22_X1 U21695 ( .A1(n18702), .A2(n18553), .B1(n18758), .B2(n18619), .ZN(
        n18550) );
  OAI211_X1 U21696 ( .C1(n18705), .C2(n18581), .A(n18551), .B(n18550), .ZN(
        P3_U2938) );
  AOI22_X1 U21697 ( .A1(n18671), .A2(n18553), .B1(n18763), .B2(n18552), .ZN(
        n18556) );
  AOI22_X1 U21698 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18554), .B1(
        n18766), .B2(n18619), .ZN(n18555) );
  OAI211_X1 U21699 ( .C1(n18675), .C2(n18581), .A(n18556), .B(n18555), .ZN(
        P3_U2939) );
  NAND2_X1 U21700 ( .A1(n18583), .A2(n18557), .ZN(n18652) );
  INV_X1 U21701 ( .A(n18583), .ZN(n18628) );
  NOR2_X1 U21702 ( .A1(n18628), .A2(n18558), .ZN(n18577) );
  AOI22_X1 U21703 ( .A1(n18714), .A2(n18577), .B1(n18715), .B2(n18602), .ZN(
        n18561) );
  NOR2_X1 U21704 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18628), .ZN(
        n18606) );
  AOI22_X1 U21705 ( .A1(n18719), .A2(n18559), .B1(n18716), .B2(n18606), .ZN(
        n18578) );
  AOI22_X1 U21706 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18578), .B1(
        n18676), .B2(n18572), .ZN(n18560) );
  OAI211_X1 U21707 ( .C1(n18684), .C2(n18652), .A(n18561), .B(n18560), .ZN(
        P3_U2940) );
  AOI22_X1 U21708 ( .A1(n18685), .A2(n18602), .B1(n18724), .B2(n18577), .ZN(
        n18563) );
  AOI22_X1 U21709 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18578), .B1(
        n18726), .B2(n18643), .ZN(n18562) );
  OAI211_X1 U21710 ( .C1(n18688), .C2(n18581), .A(n18563), .B(n18562), .ZN(
        P3_U2941) );
  AOI22_X1 U21711 ( .A1(n18564), .A2(n18602), .B1(n18730), .B2(n18577), .ZN(
        n18566) );
  AOI22_X1 U21712 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18578), .B1(
        n18732), .B2(n18643), .ZN(n18565) );
  OAI211_X1 U21713 ( .C1(n18567), .C2(n18581), .A(n18566), .B(n18565), .ZN(
        P3_U2942) );
  AOI22_X1 U21714 ( .A1(n18691), .A2(n18572), .B1(n18736), .B2(n18577), .ZN(
        n18569) );
  AOI22_X1 U21715 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18578), .B1(
        n18738), .B2(n18643), .ZN(n18568) );
  OAI211_X1 U21716 ( .C1(n18694), .C2(n18600), .A(n18569), .B(n18568), .ZN(
        P3_U2943) );
  AOI22_X1 U21717 ( .A1(n18743), .A2(n18572), .B1(n18742), .B2(n18577), .ZN(
        n18571) );
  AOI22_X1 U21718 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18578), .B1(
        n18744), .B2(n18643), .ZN(n18570) );
  OAI211_X1 U21719 ( .C1(n18747), .C2(n18600), .A(n18571), .B(n18570), .ZN(
        P3_U2944) );
  AOI22_X1 U21720 ( .A1(n18750), .A2(n18572), .B1(n18748), .B2(n18577), .ZN(
        n18574) );
  AOI22_X1 U21721 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18578), .B1(
        n18751), .B2(n18643), .ZN(n18573) );
  OAI211_X1 U21722 ( .C1(n18754), .C2(n18600), .A(n18574), .B(n18573), .ZN(
        P3_U2945) );
  AOI22_X1 U21723 ( .A1(n18757), .A2(n18602), .B1(n18756), .B2(n18577), .ZN(
        n18576) );
  AOI22_X1 U21724 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18578), .B1(
        n18758), .B2(n18643), .ZN(n18575) );
  OAI211_X1 U21725 ( .C1(n18761), .C2(n18581), .A(n18576), .B(n18575), .ZN(
        P3_U2946) );
  AOI22_X1 U21726 ( .A1(n18764), .A2(n18602), .B1(n18763), .B2(n18577), .ZN(
        n18580) );
  AOI22_X1 U21727 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18578), .B1(
        n18766), .B2(n18643), .ZN(n18579) );
  OAI211_X1 U21728 ( .C1(n18772), .C2(n18581), .A(n18580), .B(n18579), .ZN(
        P3_U2947) );
  NAND2_X1 U21729 ( .A1(n18583), .A2(n18582), .ZN(n18666) );
  AOI21_X1 U21730 ( .B1(n18652), .B2(n18666), .A(n18713), .ZN(n18601) );
  AOI22_X1 U21731 ( .A1(n18676), .A2(n18602), .B1(n18714), .B2(n18601), .ZN(
        n18587) );
  OAI211_X1 U21732 ( .C1(n18584), .C2(n18627), .A(n18652), .B(n18666), .ZN(
        n18585) );
  NAND2_X1 U21733 ( .A1(n18677), .A2(n18585), .ZN(n18603) );
  AOI22_X1 U21734 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18603), .B1(
        n18715), .B2(n18619), .ZN(n18586) );
  OAI211_X1 U21735 ( .C1(n18684), .C2(n18666), .A(n18587), .B(n18586), .ZN(
        P3_U2948) );
  AOI22_X1 U21736 ( .A1(n18685), .A2(n18619), .B1(n18724), .B2(n18601), .ZN(
        n18589) );
  INV_X1 U21737 ( .A(n18666), .ZN(n18670) );
  AOI22_X1 U21738 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18603), .B1(
        n18726), .B2(n18670), .ZN(n18588) );
  OAI211_X1 U21739 ( .C1(n18688), .C2(n18600), .A(n18589), .B(n18588), .ZN(
        P3_U2949) );
  AOI22_X1 U21740 ( .A1(n18731), .A2(n18602), .B1(n18730), .B2(n18601), .ZN(
        n18591) );
  AOI22_X1 U21741 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18603), .B1(
        n18732), .B2(n18670), .ZN(n18590) );
  OAI211_X1 U21742 ( .C1(n18735), .C2(n18626), .A(n18591), .B(n18590), .ZN(
        P3_U2950) );
  AOI22_X1 U21743 ( .A1(n18691), .A2(n18602), .B1(n18736), .B2(n18601), .ZN(
        n18593) );
  AOI22_X1 U21744 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18603), .B1(
        n18738), .B2(n18670), .ZN(n18592) );
  OAI211_X1 U21745 ( .C1(n18694), .C2(n18626), .A(n18593), .B(n18592), .ZN(
        P3_U2951) );
  AOI22_X1 U21746 ( .A1(n18639), .A2(n18619), .B1(n18742), .B2(n18601), .ZN(
        n18595) );
  AOI22_X1 U21747 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18603), .B1(
        n18744), .B2(n18670), .ZN(n18594) );
  OAI211_X1 U21748 ( .C1(n18642), .C2(n18600), .A(n18595), .B(n18594), .ZN(
        P3_U2952) );
  AOI22_X1 U21749 ( .A1(n18750), .A2(n18602), .B1(n18748), .B2(n18601), .ZN(
        n18597) );
  AOI22_X1 U21750 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18603), .B1(
        n18751), .B2(n18670), .ZN(n18596) );
  OAI211_X1 U21751 ( .C1(n18754), .C2(n18626), .A(n18597), .B(n18596), .ZN(
        P3_U2953) );
  AOI22_X1 U21752 ( .A1(n18757), .A2(n18619), .B1(n18756), .B2(n18601), .ZN(
        n18599) );
  AOI22_X1 U21753 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18603), .B1(
        n18758), .B2(n18670), .ZN(n18598) );
  OAI211_X1 U21754 ( .C1(n18761), .C2(n18600), .A(n18599), .B(n18598), .ZN(
        P3_U2954) );
  AOI22_X1 U21755 ( .A1(n18671), .A2(n18602), .B1(n18763), .B2(n18601), .ZN(
        n18605) );
  AOI22_X1 U21756 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18603), .B1(
        n18766), .B2(n18670), .ZN(n18604) );
  OAI211_X1 U21757 ( .C1(n18675), .C2(n18626), .A(n18605), .B(n18604), .ZN(
        P3_U2955) );
  NOR2_X1 U21758 ( .A1(n18801), .A2(n18628), .ZN(n18653) );
  NAND2_X1 U21759 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18653), .ZN(
        n18711) );
  AND2_X1 U21760 ( .A1(n18837), .A2(n18653), .ZN(n18622) );
  AOI22_X1 U21761 ( .A1(n18676), .A2(n18619), .B1(n18714), .B2(n18622), .ZN(
        n18608) );
  AOI22_X1 U21762 ( .A1(n18719), .A2(n18606), .B1(n18716), .B2(n18653), .ZN(
        n18623) );
  AOI22_X1 U21763 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18623), .B1(
        n18715), .B2(n18643), .ZN(n18607) );
  OAI211_X1 U21764 ( .C1(n18684), .C2(n18711), .A(n18608), .B(n18607), .ZN(
        P3_U2956) );
  AOI22_X1 U21765 ( .A1(n18685), .A2(n18643), .B1(n18724), .B2(n18622), .ZN(
        n18610) );
  AOI22_X1 U21766 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18623), .B1(
        n18726), .B2(n18701), .ZN(n18609) );
  OAI211_X1 U21767 ( .C1(n18688), .C2(n18626), .A(n18610), .B(n18609), .ZN(
        P3_U2957) );
  AOI22_X1 U21768 ( .A1(n18731), .A2(n18619), .B1(n18730), .B2(n18622), .ZN(
        n18612) );
  AOI22_X1 U21769 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18623), .B1(
        n18732), .B2(n18701), .ZN(n18611) );
  OAI211_X1 U21770 ( .C1(n18735), .C2(n18652), .A(n18612), .B(n18611), .ZN(
        P3_U2958) );
  AOI22_X1 U21771 ( .A1(n18737), .A2(n18643), .B1(n18736), .B2(n18622), .ZN(
        n18614) );
  AOI22_X1 U21772 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18623), .B1(
        n18738), .B2(n18701), .ZN(n18613) );
  OAI211_X1 U21773 ( .C1(n18741), .C2(n18626), .A(n18614), .B(n18613), .ZN(
        P3_U2959) );
  AOI22_X1 U21774 ( .A1(n18743), .A2(n18619), .B1(n18742), .B2(n18622), .ZN(
        n18616) );
  AOI22_X1 U21775 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18623), .B1(
        n18744), .B2(n18701), .ZN(n18615) );
  OAI211_X1 U21776 ( .C1(n18747), .C2(n18652), .A(n18616), .B(n18615), .ZN(
        P3_U2960) );
  AOI22_X1 U21777 ( .A1(n18697), .A2(n18643), .B1(n18748), .B2(n18622), .ZN(
        n18618) );
  AOI22_X1 U21778 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18623), .B1(
        n18751), .B2(n18701), .ZN(n18617) );
  OAI211_X1 U21779 ( .C1(n18700), .C2(n18626), .A(n18618), .B(n18617), .ZN(
        P3_U2961) );
  AOI22_X1 U21780 ( .A1(n18702), .A2(n18619), .B1(n18756), .B2(n18622), .ZN(
        n18621) );
  AOI22_X1 U21781 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18623), .B1(
        n18758), .B2(n18701), .ZN(n18620) );
  OAI211_X1 U21782 ( .C1(n18705), .C2(n18652), .A(n18621), .B(n18620), .ZN(
        P3_U2962) );
  AOI22_X1 U21783 ( .A1(n18764), .A2(n18643), .B1(n18763), .B2(n18622), .ZN(
        n18625) );
  AOI22_X1 U21784 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18623), .B1(
        n18766), .B2(n18701), .ZN(n18624) );
  OAI211_X1 U21785 ( .C1(n18772), .C2(n18626), .A(n18625), .B(n18624), .ZN(
        P3_U2963) );
  NAND2_X1 U21786 ( .A1(n18718), .A2(n18800), .ZN(n18771) );
  NOR3_X1 U21787 ( .A1(n18629), .A2(n18628), .A3(n18627), .ZN(n18630) );
  NAND2_X1 U21788 ( .A1(n18711), .A2(n18771), .ZN(n18678) );
  OAI21_X1 U21789 ( .B1(n18630), .B2(n18678), .A(n18677), .ZN(n18649) );
  AND2_X1 U21790 ( .A1(n18837), .A2(n18678), .ZN(n18648) );
  AOI22_X1 U21791 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18649), .B1(
        n18714), .B2(n18648), .ZN(n18632) );
  AOI22_X1 U21792 ( .A1(n18676), .A2(n18643), .B1(n18715), .B2(n18670), .ZN(
        n18631) );
  OAI211_X1 U21793 ( .C1(n18684), .C2(n18771), .A(n18632), .B(n18631), .ZN(
        P3_U2964) );
  AOI22_X1 U21794 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18649), .B1(
        n18724), .B2(n18648), .ZN(n18634) );
  INV_X1 U21795 ( .A(n18771), .ZN(n18749) );
  AOI22_X1 U21796 ( .A1(n18726), .A2(n18749), .B1(n18685), .B2(n18670), .ZN(
        n18633) );
  OAI211_X1 U21797 ( .C1(n18688), .C2(n18652), .A(n18634), .B(n18633), .ZN(
        P3_U2965) );
  AOI22_X1 U21798 ( .A1(n18731), .A2(n18643), .B1(n18730), .B2(n18648), .ZN(
        n18636) );
  AOI22_X1 U21799 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18649), .B1(
        n18732), .B2(n18749), .ZN(n18635) );
  OAI211_X1 U21800 ( .C1(n18735), .C2(n18666), .A(n18636), .B(n18635), .ZN(
        P3_U2966) );
  AOI22_X1 U21801 ( .A1(n18737), .A2(n18670), .B1(n18736), .B2(n18648), .ZN(
        n18638) );
  AOI22_X1 U21802 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18649), .B1(
        n18738), .B2(n18749), .ZN(n18637) );
  OAI211_X1 U21803 ( .C1(n18741), .C2(n18652), .A(n18638), .B(n18637), .ZN(
        P3_U2967) );
  AOI22_X1 U21804 ( .A1(n18639), .A2(n18670), .B1(n18742), .B2(n18648), .ZN(
        n18641) );
  AOI22_X1 U21805 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18649), .B1(
        n18744), .B2(n18749), .ZN(n18640) );
  OAI211_X1 U21806 ( .C1(n18642), .C2(n18652), .A(n18641), .B(n18640), .ZN(
        P3_U2968) );
  AOI22_X1 U21807 ( .A1(n18750), .A2(n18643), .B1(n18748), .B2(n18648), .ZN(
        n18645) );
  AOI22_X1 U21808 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18649), .B1(
        n18751), .B2(n18749), .ZN(n18644) );
  OAI211_X1 U21809 ( .C1(n18754), .C2(n18666), .A(n18645), .B(n18644), .ZN(
        P3_U2969) );
  AOI22_X1 U21810 ( .A1(n18757), .A2(n18670), .B1(n18756), .B2(n18648), .ZN(
        n18647) );
  AOI22_X1 U21811 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18649), .B1(
        n18758), .B2(n18749), .ZN(n18646) );
  OAI211_X1 U21812 ( .C1(n18761), .C2(n18652), .A(n18647), .B(n18646), .ZN(
        P3_U2970) );
  AOI22_X1 U21813 ( .A1(n18764), .A2(n18670), .B1(n18763), .B2(n18648), .ZN(
        n18651) );
  AOI22_X1 U21814 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18649), .B1(
        n18766), .B2(n18749), .ZN(n18650) );
  OAI211_X1 U21815 ( .C1(n18772), .C2(n18652), .A(n18651), .B(n18650), .ZN(
        P3_U2971) );
  AND2_X1 U21816 ( .A1(n18837), .A2(n18718), .ZN(n18669) );
  AOI22_X1 U21817 ( .A1(n18676), .A2(n18670), .B1(n18714), .B2(n18669), .ZN(
        n18655) );
  AOI22_X1 U21818 ( .A1(n18719), .A2(n18653), .B1(n18718), .B2(n18716), .ZN(
        n18672) );
  AOI22_X1 U21819 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18672), .B1(
        n18715), .B2(n18701), .ZN(n18654) );
  OAI211_X1 U21820 ( .C1(n18755), .C2(n18684), .A(n18655), .B(n18654), .ZN(
        P3_U2972) );
  AOI22_X1 U21821 ( .A1(n18725), .A2(n18670), .B1(n18724), .B2(n18669), .ZN(
        n18657) );
  AOI22_X1 U21822 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18672), .B1(
        n18765), .B2(n18726), .ZN(n18656) );
  OAI211_X1 U21823 ( .C1(n18729), .C2(n18711), .A(n18657), .B(n18656), .ZN(
        P3_U2973) );
  AOI22_X1 U21824 ( .A1(n18731), .A2(n18670), .B1(n18730), .B2(n18669), .ZN(
        n18659) );
  AOI22_X1 U21825 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18672), .B1(
        n18765), .B2(n18732), .ZN(n18658) );
  OAI211_X1 U21826 ( .C1(n18735), .C2(n18711), .A(n18659), .B(n18658), .ZN(
        P3_U2974) );
  AOI22_X1 U21827 ( .A1(n18737), .A2(n18701), .B1(n18736), .B2(n18669), .ZN(
        n18661) );
  AOI22_X1 U21828 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18672), .B1(
        n18765), .B2(n18738), .ZN(n18660) );
  OAI211_X1 U21829 ( .C1(n18741), .C2(n18666), .A(n18661), .B(n18660), .ZN(
        P3_U2975) );
  AOI22_X1 U21830 ( .A1(n18743), .A2(n18670), .B1(n18742), .B2(n18669), .ZN(
        n18663) );
  AOI22_X1 U21831 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18672), .B1(
        n18765), .B2(n18744), .ZN(n18662) );
  OAI211_X1 U21832 ( .C1(n18747), .C2(n18711), .A(n18663), .B(n18662), .ZN(
        P3_U2976) );
  AOI22_X1 U21833 ( .A1(n18697), .A2(n18701), .B1(n18748), .B2(n18669), .ZN(
        n18665) );
  AOI22_X1 U21834 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18672), .B1(
        n18765), .B2(n18751), .ZN(n18664) );
  OAI211_X1 U21835 ( .C1(n18700), .C2(n18666), .A(n18665), .B(n18664), .ZN(
        P3_U2977) );
  AOI22_X1 U21836 ( .A1(n18702), .A2(n18670), .B1(n18756), .B2(n18669), .ZN(
        n18668) );
  AOI22_X1 U21837 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18672), .B1(
        n18765), .B2(n18758), .ZN(n18667) );
  OAI211_X1 U21838 ( .C1(n18705), .C2(n18711), .A(n18668), .B(n18667), .ZN(
        P3_U2978) );
  AOI22_X1 U21839 ( .A1(n18671), .A2(n18670), .B1(n18763), .B2(n18669), .ZN(
        n18674) );
  AOI22_X1 U21840 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18672), .B1(
        n18765), .B2(n18766), .ZN(n18673) );
  OAI211_X1 U21841 ( .C1(n18675), .C2(n18711), .A(n18674), .B(n18673), .ZN(
        P3_U2979) );
  AND2_X1 U21842 ( .A1(n18837), .A2(n18680), .ZN(n18706) );
  AOI22_X1 U21843 ( .A1(n18676), .A2(n18701), .B1(n18714), .B2(n18706), .ZN(
        n18682) );
  OAI221_X1 U21844 ( .B1(n18680), .B2(n18679), .C1(n18680), .C2(n18678), .A(
        n18677), .ZN(n18708) );
  AOI22_X1 U21845 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18708), .B1(
        n18715), .B2(n18749), .ZN(n18681) );
  OAI211_X1 U21846 ( .C1(n18684), .C2(n18683), .A(n18682), .B(n18681), .ZN(
        P3_U2980) );
  AOI22_X1 U21847 ( .A1(n18685), .A2(n18749), .B1(n18724), .B2(n18706), .ZN(
        n18687) );
  AOI22_X1 U21848 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18708), .B1(
        n18707), .B2(n18726), .ZN(n18686) );
  OAI211_X1 U21849 ( .C1(n18688), .C2(n18711), .A(n18687), .B(n18686), .ZN(
        P3_U2981) );
  AOI22_X1 U21850 ( .A1(n18731), .A2(n18701), .B1(n18730), .B2(n18706), .ZN(
        n18690) );
  AOI22_X1 U21851 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18708), .B1(
        n18707), .B2(n18732), .ZN(n18689) );
  OAI211_X1 U21852 ( .C1(n18735), .C2(n18771), .A(n18690), .B(n18689), .ZN(
        P3_U2982) );
  AOI22_X1 U21853 ( .A1(n18691), .A2(n18701), .B1(n18736), .B2(n18706), .ZN(
        n18693) );
  AOI22_X1 U21854 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18708), .B1(
        n18707), .B2(n18738), .ZN(n18692) );
  OAI211_X1 U21855 ( .C1(n18694), .C2(n18771), .A(n18693), .B(n18692), .ZN(
        P3_U2983) );
  AOI22_X1 U21856 ( .A1(n18743), .A2(n18701), .B1(n18742), .B2(n18706), .ZN(
        n18696) );
  AOI22_X1 U21857 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18708), .B1(
        n18707), .B2(n18744), .ZN(n18695) );
  OAI211_X1 U21858 ( .C1(n18747), .C2(n18771), .A(n18696), .B(n18695), .ZN(
        P3_U2984) );
  AOI22_X1 U21859 ( .A1(n18697), .A2(n18749), .B1(n18748), .B2(n18706), .ZN(
        n18699) );
  AOI22_X1 U21860 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18708), .B1(
        n18707), .B2(n18751), .ZN(n18698) );
  OAI211_X1 U21861 ( .C1(n18700), .C2(n18711), .A(n18699), .B(n18698), .ZN(
        P3_U2985) );
  AOI22_X1 U21862 ( .A1(n18702), .A2(n18701), .B1(n18756), .B2(n18706), .ZN(
        n18704) );
  AOI22_X1 U21863 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18708), .B1(
        n18707), .B2(n18758), .ZN(n18703) );
  OAI211_X1 U21864 ( .C1(n18705), .C2(n18771), .A(n18704), .B(n18703), .ZN(
        P3_U2986) );
  AOI22_X1 U21865 ( .A1(n18764), .A2(n18749), .B1(n18763), .B2(n18706), .ZN(
        n18710) );
  AOI22_X1 U21866 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18708), .B1(
        n18707), .B2(n18766), .ZN(n18709) );
  OAI211_X1 U21867 ( .C1(n18772), .C2(n18711), .A(n18710), .B(n18709), .ZN(
        P3_U2987) );
  NOR2_X1 U21868 ( .A1(n18713), .A2(n18712), .ZN(n18762) );
  AOI22_X1 U21869 ( .A1(n18765), .A2(n18715), .B1(n18714), .B2(n18762), .ZN(
        n18722) );
  AOI22_X1 U21870 ( .A1(n18719), .A2(n18718), .B1(n18717), .B2(n18716), .ZN(
        n18768) );
  AOI22_X1 U21871 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18768), .B1(
        n18767), .B2(n18720), .ZN(n18721) );
  OAI211_X1 U21872 ( .C1(n18723), .C2(n18771), .A(n18722), .B(n18721), .ZN(
        P3_U2988) );
  AOI22_X1 U21873 ( .A1(n18725), .A2(n18749), .B1(n18724), .B2(n18762), .ZN(
        n18728) );
  AOI22_X1 U21874 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18768), .B1(
        n18767), .B2(n18726), .ZN(n18727) );
  OAI211_X1 U21875 ( .C1(n18755), .C2(n18729), .A(n18728), .B(n18727), .ZN(
        P3_U2989) );
  AOI22_X1 U21876 ( .A1(n18731), .A2(n18749), .B1(n18730), .B2(n18762), .ZN(
        n18734) );
  AOI22_X1 U21877 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18768), .B1(
        n18767), .B2(n18732), .ZN(n18733) );
  OAI211_X1 U21878 ( .C1(n18755), .C2(n18735), .A(n18734), .B(n18733), .ZN(
        P3_U2990) );
  AOI22_X1 U21879 ( .A1(n18765), .A2(n18737), .B1(n18736), .B2(n18762), .ZN(
        n18740) );
  AOI22_X1 U21880 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18768), .B1(
        n18767), .B2(n18738), .ZN(n18739) );
  OAI211_X1 U21881 ( .C1(n18741), .C2(n18771), .A(n18740), .B(n18739), .ZN(
        P3_U2991) );
  AOI22_X1 U21882 ( .A1(n18743), .A2(n18749), .B1(n18742), .B2(n18762), .ZN(
        n18746) );
  AOI22_X1 U21883 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18768), .B1(
        n18767), .B2(n18744), .ZN(n18745) );
  OAI211_X1 U21884 ( .C1(n18755), .C2(n18747), .A(n18746), .B(n18745), .ZN(
        P3_U2992) );
  AOI22_X1 U21885 ( .A1(n18750), .A2(n18749), .B1(n18748), .B2(n18762), .ZN(
        n18753) );
  AOI22_X1 U21886 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18768), .B1(
        n18767), .B2(n18751), .ZN(n18752) );
  OAI211_X1 U21887 ( .C1(n18755), .C2(n18754), .A(n18753), .B(n18752), .ZN(
        P3_U2993) );
  AOI22_X1 U21888 ( .A1(n18765), .A2(n18757), .B1(n18756), .B2(n18762), .ZN(
        n18760) );
  AOI22_X1 U21889 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18768), .B1(
        n18767), .B2(n18758), .ZN(n18759) );
  OAI211_X1 U21890 ( .C1(n18761), .C2(n18771), .A(n18760), .B(n18759), .ZN(
        P3_U2994) );
  AOI22_X1 U21891 ( .A1(n18765), .A2(n18764), .B1(n18763), .B2(n18762), .ZN(
        n18770) );
  AOI22_X1 U21892 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18768), .B1(
        n18767), .B2(n18766), .ZN(n18769) );
  OAI211_X1 U21893 ( .C1(n18772), .C2(n18771), .A(n18770), .B(n18769), .ZN(
        P3_U2995) );
  NOR2_X1 U21894 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n18999) );
  NAND2_X1 U21895 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18999), .ZN(n18832) );
  OAI22_X1 U21896 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18832), .B1(
        n18773), .B2(n18988), .ZN(n18836) );
  NOR3_X1 U21897 ( .A1(n18993), .A2(n18775), .A3(n18774), .ZN(n18829) );
  NAND2_X1 U21898 ( .A1(n18792), .A2(n18776), .ZN(n18781) );
  AOI222_X1 U21899 ( .A1(n18782), .A2(n18781), .B1(n18780), .B2(n18779), .C1(
        n18778), .C2(n18777), .ZN(n18986) );
  AOI211_X1 U21900 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n18816), .A(
        n18784), .B(n18783), .ZN(n18827) );
  AOI21_X1 U21901 ( .B1(n18787), .B2(n18786), .A(n18785), .ZN(n18814) );
  AOI22_X1 U21902 ( .A1(n10256), .A2(n18807), .B1(n18809), .B2(n18791), .ZN(
        n18788) );
  OAI21_X1 U21903 ( .B1(n18789), .B2(n18814), .A(n18788), .ZN(n18948) );
  NOR2_X1 U21904 ( .A1(n11435), .A2(n18948), .ZN(n18795) );
  INV_X1 U21905 ( .A(n18790), .ZN(n18793) );
  AOI21_X1 U21906 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18797), .A(
        n18791), .ZN(n18808) );
  OAI22_X1 U21907 ( .A1(n18793), .A2(n18792), .B1(n18808), .B2(n18809), .ZN(
        n18945) );
  AOI21_X1 U21908 ( .B1(n18945), .B2(n18815), .A(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18794) );
  AOI21_X1 U21909 ( .B1(n18815), .B2(n18795), .A(n18794), .ZN(n18823) );
  NOR2_X1 U21910 ( .A1(n18797), .A2(n18796), .ZN(n18798) );
  OAI22_X1 U21911 ( .A1(n18958), .A2(n18798), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18808), .ZN(n18962) );
  INV_X1 U21912 ( .A(n18962), .ZN(n18804) );
  OAI22_X1 U21913 ( .A1(n18972), .A2(n18799), .B1(n18798), .B2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18802) );
  NOR3_X1 U21914 ( .A1(n18801), .A2(n18800), .A3(n18802), .ZN(n18803) );
  INV_X1 U21915 ( .A(n18802), .ZN(n18966) );
  OAI22_X1 U21916 ( .A1(n18804), .A2(n18803), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18966), .ZN(n18806) );
  AOI21_X1 U21917 ( .B1(n18806), .B2(n18815), .A(n18805), .ZN(n18818) );
  NAND2_X1 U21918 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18807), .ZN(
        n18813) );
  AOI21_X1 U21919 ( .B1(n18964), .B2(n10256), .A(n18808), .ZN(n18810) );
  AOI22_X1 U21920 ( .A1(n18811), .A2(n18953), .B1(n18810), .B2(n18809), .ZN(
        n18812) );
  OAI21_X1 U21921 ( .B1(n18814), .B2(n18813), .A(n18812), .ZN(n18956) );
  AOI22_X1 U21922 ( .A1(n18816), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n18956), .B2(n18815), .ZN(n18819) );
  OR2_X1 U21923 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18819), .ZN(
        n18817) );
  AOI221_X1 U21924 ( .B1(n18818), .B2(n18817), .C1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C2(n18819), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18822) );
  OAI21_X1 U21925 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n18819), .ZN(n18821) );
  AOI222_X1 U21926 ( .A1(n18823), .A2(n18822), .B1(n18823), .B2(n18821), .C1(
        n18822), .C2(n18820), .ZN(n18826) );
  OAI21_X1 U21927 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18824), .ZN(n18825) );
  NAND4_X1 U21928 ( .A1(n18986), .A2(n18827), .A3(n18826), .A4(n18825), .ZN(
        n18833) );
  NOR3_X1 U21929 ( .A1(n18829), .A2(n18833), .A3(n18828), .ZN(n18940) );
  AOI21_X1 U21930 ( .B1(n18994), .B2(n19005), .A(n18940), .ZN(n18838) );
  INV_X1 U21931 ( .A(n18830), .ZN(n18831) );
  NAND3_X1 U21932 ( .A1(n18838), .A2(n18832), .A3(n18831), .ZN(n18834) );
  AOI22_X1 U21933 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18834), .B1(n18991), 
        .B2(n18833), .ZN(n18835) );
  OAI21_X1 U21934 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18836), .A(n18835), 
        .ZN(P3_U2996) );
  NAND2_X1 U21935 ( .A1(n18994), .A2(n17550), .ZN(n18841) );
  NAND3_X1 U21936 ( .A1(n18994), .A2(n18844), .A3(n19005), .ZN(n18843) );
  NAND3_X1 U21937 ( .A1(n18839), .A2(n18838), .A3(n18837), .ZN(n18840) );
  NAND4_X1 U21938 ( .A1(n18842), .A2(n18841), .A3(n18843), .A4(n18840), .ZN(
        P3_U2997) );
  INV_X1 U21939 ( .A(n18843), .ZN(n18848) );
  NOR3_X1 U21940 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18845), .A3(n18844), 
        .ZN(n18846) );
  NOR3_X1 U21941 ( .A1(n18848), .A2(n18847), .A3(n18846), .ZN(P3_U2998) );
  AND2_X1 U21942 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18936), .ZN(
        P3_U2999) );
  AND2_X1 U21943 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18936), .ZN(
        P3_U3000) );
  AND2_X1 U21944 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18936), .ZN(
        P3_U3001) );
  AND2_X1 U21945 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18936), .ZN(
        P3_U3002) );
  AND2_X1 U21946 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18936), .ZN(
        P3_U3003) );
  AND2_X1 U21947 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18936), .ZN(
        P3_U3004) );
  AND2_X1 U21948 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18936), .ZN(
        P3_U3005) );
  AND2_X1 U21949 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18936), .ZN(
        P3_U3006) );
  AND2_X1 U21950 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18936), .ZN(
        P3_U3007) );
  AND2_X1 U21951 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18936), .ZN(
        P3_U3008) );
  AND2_X1 U21952 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18936), .ZN(
        P3_U3009) );
  AND2_X1 U21953 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18936), .ZN(
        P3_U3010) );
  AND2_X1 U21954 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18936), .ZN(
        P3_U3011) );
  AND2_X1 U21955 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18936), .ZN(
        P3_U3012) );
  AND2_X1 U21956 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18936), .ZN(
        P3_U3013) );
  AND2_X1 U21957 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18936), .ZN(
        P3_U3014) );
  AND2_X1 U21958 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18936), .ZN(
        P3_U3015) );
  AND2_X1 U21959 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18936), .ZN(
        P3_U3016) );
  AND2_X1 U21960 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18936), .ZN(
        P3_U3017) );
  AND2_X1 U21961 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18936), .ZN(
        P3_U3018) );
  AND2_X1 U21962 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18936), .ZN(
        P3_U3019) );
  AND2_X1 U21963 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18936), .ZN(
        P3_U3020) );
  AND2_X1 U21964 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18936), .ZN(P3_U3021) );
  AND2_X1 U21965 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18936), .ZN(P3_U3022) );
  AND2_X1 U21966 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18936), .ZN(P3_U3023) );
  AND2_X1 U21967 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18936), .ZN(P3_U3024) );
  AND2_X1 U21968 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18936), .ZN(P3_U3025) );
  AND2_X1 U21969 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18936), .ZN(P3_U3026) );
  AND2_X1 U21970 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18936), .ZN(P3_U3027) );
  AND2_X1 U21971 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18936), .ZN(P3_U3028) );
  OAI21_X1 U21972 ( .B1(n18849), .B2(n21002), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18850) );
  AOI22_X1 U21973 ( .A1(n18862), .A2(n18864), .B1(n19003), .B2(n18850), .ZN(
        n18852) );
  INV_X1 U21974 ( .A(NA), .ZN(n21132) );
  OR3_X1 U21975 ( .A1(n21132), .A2(P3_STATE_REG_0__SCAN_IN), .A3(
        P3_STATE_REG_1__SCAN_IN), .ZN(n18851) );
  OAI211_X1 U21976 ( .C1(n18988), .C2(n18856), .A(n18852), .B(n18851), .ZN(
        P3_U3029) );
  NOR2_X1 U21977 ( .A1(n18864), .A2(n21002), .ZN(n18860) );
  INV_X1 U21978 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19001) );
  NOR3_X1 U21979 ( .A1(n18860), .A2(n19001), .A3(n18862), .ZN(n18853) );
  NAND2_X1 U21980 ( .A1(n18994), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18858) );
  INV_X1 U21981 ( .A(n18858), .ZN(n18857) );
  NOR2_X1 U21982 ( .A1(n18853), .A2(n18857), .ZN(n18855) );
  OAI211_X1 U21983 ( .C1(n21002), .C2(n18856), .A(n18855), .B(n18854), .ZN(
        P3_U3030) );
  AOI221_X1 U21984 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n18862), .C1(n21132), 
        .C2(n18862), .A(n18857), .ZN(n18863) );
  OAI22_X1 U21985 ( .A1(NA), .A2(n18858), .B1(P3_STATE_REG_1__SCAN_IN), .B2(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18859) );
  OAI22_X1 U21986 ( .A1(n18860), .A2(n18859), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18861) );
  OAI22_X1 U21987 ( .A1(n18863), .A2(n18864), .B1(n18862), .B2(n18861), .ZN(
        P3_U3031) );
  OAI222_X1 U21988 ( .A1(n18974), .A2(n18922), .B1(n18865), .B2(n18933), .C1(
        n18866), .C2(n18926), .ZN(P3_U3032) );
  INV_X1 U21989 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18868) );
  OAI222_X1 U21990 ( .A1(n18926), .A2(n18868), .B1(n18867), .B2(n18933), .C1(
        n18866), .C2(n18922), .ZN(P3_U3033) );
  OAI222_X1 U21991 ( .A1(n18926), .A2(n18870), .B1(n18869), .B2(n18933), .C1(
        n18868), .C2(n18922), .ZN(P3_U3034) );
  OAI222_X1 U21992 ( .A1(n18926), .A2(n18872), .B1(n18871), .B2(n18933), .C1(
        n18870), .C2(n18922), .ZN(P3_U3035) );
  OAI222_X1 U21993 ( .A1(n18926), .A2(n18874), .B1(n18873), .B2(n18933), .C1(
        n18872), .C2(n18922), .ZN(P3_U3036) );
  OAI222_X1 U21994 ( .A1(n18926), .A2(n18876), .B1(n18875), .B2(n18933), .C1(
        n18874), .C2(n18922), .ZN(P3_U3037) );
  OAI222_X1 U21995 ( .A1(n18926), .A2(n18879), .B1(n18877), .B2(n18933), .C1(
        n18876), .C2(n18922), .ZN(P3_U3038) );
  OAI222_X1 U21996 ( .A1(n18879), .A2(n18922), .B1(n18878), .B2(n18933), .C1(
        n18880), .C2(n18926), .ZN(P3_U3039) );
  OAI222_X1 U21997 ( .A1(n18926), .A2(n18882), .B1(n18881), .B2(n18933), .C1(
        n18880), .C2(n18922), .ZN(P3_U3040) );
  OAI222_X1 U21998 ( .A1(n18926), .A2(n18884), .B1(n18883), .B2(n18933), .C1(
        n18882), .C2(n18922), .ZN(P3_U3041) );
  OAI222_X1 U21999 ( .A1(n18926), .A2(n18886), .B1(n18885), .B2(n18933), .C1(
        n18884), .C2(n18922), .ZN(P3_U3042) );
  OAI222_X1 U22000 ( .A1(n18926), .A2(n18888), .B1(n18887), .B2(n18933), .C1(
        n18886), .C2(n18922), .ZN(P3_U3043) );
  OAI222_X1 U22001 ( .A1(n18926), .A2(n18891), .B1(n18889), .B2(n18933), .C1(
        n18888), .C2(n18922), .ZN(P3_U3044) );
  OAI222_X1 U22002 ( .A1(n18891), .A2(n18922), .B1(n18890), .B2(n18933), .C1(
        n18892), .C2(n18926), .ZN(P3_U3045) );
  OAI222_X1 U22003 ( .A1(n18926), .A2(n18894), .B1(n18893), .B2(n18933), .C1(
        n18892), .C2(n18922), .ZN(P3_U3046) );
  OAI222_X1 U22004 ( .A1(n18926), .A2(n18896), .B1(n18895), .B2(n18933), .C1(
        n18894), .C2(n18922), .ZN(P3_U3047) );
  OAI222_X1 U22005 ( .A1(n18926), .A2(n18898), .B1(n18897), .B2(n18933), .C1(
        n18896), .C2(n18922), .ZN(P3_U3048) );
  OAI222_X1 U22006 ( .A1(n18926), .A2(n18901), .B1(n18899), .B2(n18933), .C1(
        n18898), .C2(n18922), .ZN(P3_U3049) );
  OAI222_X1 U22007 ( .A1(n18901), .A2(n18922), .B1(n18900), .B2(n18933), .C1(
        n18902), .C2(n18926), .ZN(P3_U3050) );
  OAI222_X1 U22008 ( .A1(n18926), .A2(n18905), .B1(n18903), .B2(n18933), .C1(
        n18902), .C2(n18922), .ZN(P3_U3051) );
  OAI222_X1 U22009 ( .A1(n18905), .A2(n18922), .B1(n18904), .B2(n18933), .C1(
        n18906), .C2(n18926), .ZN(P3_U3052) );
  OAI222_X1 U22010 ( .A1(n18926), .A2(n18909), .B1(n18907), .B2(n18933), .C1(
        n18906), .C2(n18922), .ZN(P3_U3053) );
  OAI222_X1 U22011 ( .A1(n18909), .A2(n18922), .B1(n18908), .B2(n18933), .C1(
        n18910), .C2(n18926), .ZN(P3_U3054) );
  INV_X1 U22012 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18912) );
  OAI222_X1 U22013 ( .A1(n18926), .A2(n18912), .B1(n18911), .B2(n18933), .C1(
        n18910), .C2(n18922), .ZN(P3_U3055) );
  INV_X1 U22014 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18914) );
  OAI222_X1 U22015 ( .A1(n18926), .A2(n18914), .B1(n18913), .B2(n18933), .C1(
        n18912), .C2(n18922), .ZN(P3_U3056) );
  OAI222_X1 U22016 ( .A1(n18926), .A2(n18916), .B1(n18915), .B2(n18933), .C1(
        n18914), .C2(n18922), .ZN(P3_U3057) );
  OAI222_X1 U22017 ( .A1(n18926), .A2(n18919), .B1(n18917), .B2(n18933), .C1(
        n18916), .C2(n18922), .ZN(P3_U3058) );
  OAI222_X1 U22018 ( .A1(n18919), .A2(n18922), .B1(n18918), .B2(n18933), .C1(
        n18920), .C2(n18926), .ZN(P3_U3059) );
  OAI222_X1 U22019 ( .A1(n18926), .A2(n18923), .B1(n18921), .B2(n18933), .C1(
        n18920), .C2(n18922), .ZN(P3_U3060) );
  INV_X1 U22020 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18924) );
  OAI222_X1 U22021 ( .A1(n18926), .A2(n18925), .B1(n18924), .B2(n18933), .C1(
        n18923), .C2(n18922), .ZN(P3_U3061) );
  INV_X1 U22022 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n18927) );
  AOI22_X1 U22023 ( .A1(n18933), .A2(n18928), .B1(n18927), .B2(n19003), .ZN(
        P3_U3274) );
  INV_X1 U22024 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18976) );
  INV_X1 U22025 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n18929) );
  AOI22_X1 U22026 ( .A1(n18933), .A2(n18976), .B1(n18929), .B2(n19003), .ZN(
        P3_U3275) );
  INV_X1 U22027 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n18930) );
  AOI22_X1 U22028 ( .A1(n18933), .A2(n18931), .B1(n18930), .B2(n19003), .ZN(
        P3_U3276) );
  INV_X1 U22029 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18982) );
  INV_X1 U22030 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n18932) );
  AOI22_X1 U22031 ( .A1(n18933), .A2(n18982), .B1(n18932), .B2(n19003), .ZN(
        P3_U3277) );
  INV_X1 U22032 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18935) );
  INV_X1 U22033 ( .A(n18937), .ZN(n18934) );
  AOI21_X1 U22034 ( .B1(n18936), .B2(n18935), .A(n18934), .ZN(P3_U3280) );
  OAI21_X1 U22035 ( .B1(n18939), .B2(n18938), .A(n18937), .ZN(P3_U3281) );
  NOR2_X1 U22036 ( .A1(n18940), .A2(n18996), .ZN(n18943) );
  OAI21_X1 U22037 ( .B1(n18943), .B2(n18942), .A(n18941), .ZN(P3_U3282) );
  INV_X1 U22038 ( .A(n18954), .ZN(n18969) );
  NOR2_X1 U22039 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18944), .ZN(
        n18946) );
  AOI22_X1 U22040 ( .A1(n18969), .A2(n18947), .B1(n18946), .B2(n18945), .ZN(
        n18950) );
  AOI21_X1 U22041 ( .B1(n19006), .B2(n18948), .A(n18973), .ZN(n18949) );
  OAI22_X1 U22042 ( .A1(n18973), .A2(n18950), .B1(n18949), .B2(n11435), .ZN(
        P3_U3285) );
  NAND2_X1 U22043 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18968) );
  AOI22_X1 U22044 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n18952), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n18951), .ZN(n18960) );
  OAI22_X1 U22045 ( .A1(n18954), .A2(n18953), .B1(n18968), .B2(n18960), .ZN(
        n18955) );
  AOI21_X1 U22046 ( .B1(n19006), .B2(n18956), .A(n18955), .ZN(n18957) );
  AOI22_X1 U22047 ( .A1(n18973), .A2(n10256), .B1(n18957), .B2(n18970), .ZN(
        P3_U3288) );
  INV_X1 U22048 ( .A(n18958), .ZN(n18961) );
  INV_X1 U22049 ( .A(n18968), .ZN(n18959) );
  AOI222_X1 U22050 ( .A1(n18962), .A2(n19006), .B1(n18969), .B2(n18961), .C1(
        n18960), .C2(n18959), .ZN(n18963) );
  AOI22_X1 U22051 ( .A1(n18973), .A2(n18964), .B1(n18963), .B2(n18970), .ZN(
        P3_U3289) );
  OAI21_X1 U22052 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18966), .A(n18965), 
        .ZN(n18967) );
  AOI22_X1 U22053 ( .A1(n18969), .A2(n18972), .B1(n18968), .B2(n18967), .ZN(
        n18971) );
  AOI22_X1 U22054 ( .A1(n18973), .A2(n18972), .B1(n18971), .B2(n18970), .ZN(
        P3_U3290) );
  AOI21_X1 U22055 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18975) );
  AOI22_X1 U22056 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18975), .B2(n18974), .ZN(n18977) );
  AOI22_X1 U22057 ( .A1(n18978), .A2(n18977), .B1(n18976), .B2(n18981), .ZN(
        P3_U3292) );
  NOR2_X1 U22058 ( .A1(n18981), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18979) );
  AOI22_X1 U22059 ( .A1(n18982), .A2(n18981), .B1(n18980), .B2(n18979), .ZN(
        P3_U3293) );
  INV_X1 U22060 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18983) );
  AOI22_X1 U22061 ( .A1(n18933), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18983), 
        .B2(n19003), .ZN(P3_U3294) );
  INV_X1 U22062 ( .A(n18984), .ZN(n18987) );
  NAND2_X1 U22063 ( .A1(n18987), .A2(P3_MORE_REG_SCAN_IN), .ZN(n18985) );
  OAI21_X1 U22064 ( .B1(n18987), .B2(n18986), .A(n18985), .ZN(P3_U3295) );
  AOI21_X1 U22065 ( .B1(n17550), .B2(n18988), .A(n19008), .ZN(n18989) );
  OAI21_X1 U22066 ( .B1(n18991), .B2(n18990), .A(n18989), .ZN(n19002) );
  OAI21_X1 U22067 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n18993), .A(n18992), 
        .ZN(n18995) );
  AOI211_X1 U22068 ( .C1(n19007), .C2(n18995), .A(n18994), .B(n19005), .ZN(
        n18997) );
  NOR2_X1 U22069 ( .A1(n18997), .A2(n18996), .ZN(n18998) );
  OAI21_X1 U22070 ( .B1(n18999), .B2(n18998), .A(n19002), .ZN(n19000) );
  OAI21_X1 U22071 ( .B1(n19002), .B2(n19001), .A(n19000), .ZN(P3_U3296) );
  INV_X1 U22072 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n19011) );
  INV_X1 U22073 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n19004) );
  AOI22_X1 U22074 ( .A1(n18933), .A2(n19011), .B1(n19004), .B2(n19003), .ZN(
        P3_U3297) );
  AOI21_X1 U22075 ( .B1(n19006), .B2(n19005), .A(n19008), .ZN(n19012) );
  INV_X1 U22076 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n19009) );
  AOI22_X1 U22077 ( .A1(n19012), .A2(n19009), .B1(n19008), .B2(n19007), .ZN(
        P3_U3298) );
  AOI21_X1 U22078 ( .B1(n19012), .B2(n19011), .A(n19010), .ZN(P3_U3299) );
  INV_X1 U22079 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19018) );
  INV_X1 U22080 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n19013) );
  NAND2_X1 U22081 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20055), .ZN(n20045) );
  NAND2_X1 U22082 ( .A1(n19018), .A2(n19017), .ZN(n20042) );
  OAI21_X1 U22083 ( .B1(n19018), .B2(n20045), .A(n20042), .ZN(n20119) );
  OAI21_X1 U22084 ( .B1(n19018), .B2(n19013), .A(n20035), .ZN(P2_U2815) );
  INV_X1 U22085 ( .A(n19014), .ZN(n19015) );
  AOI22_X1 U22086 ( .A1(n19015), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n20029), 
        .B2(n20030), .ZN(n19016) );
  INV_X1 U22087 ( .A(n19016), .ZN(P2_U2816) );
  INV_X2 U22088 ( .A(n20175), .ZN(n20178) );
  AOI21_X1 U22089 ( .B1(n19018), .B2(n20055), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n19019) );
  AOI22_X1 U22090 ( .A1(n20178), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n19019), 
        .B2(n20175), .ZN(P2_U2817) );
  OAI21_X1 U22091 ( .B1(n20036), .B2(BS16), .A(n20119), .ZN(n20117) );
  OAI21_X1 U22092 ( .B1(n20119), .B2(n19612), .A(n20117), .ZN(P2_U2818) );
  NOR4_X1 U22093 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19023) );
  NOR4_X1 U22094 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19022) );
  NOR4_X1 U22095 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19021) );
  NOR4_X1 U22096 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19020) );
  NAND4_X1 U22097 ( .A1(n19023), .A2(n19022), .A3(n19021), .A4(n19020), .ZN(
        n19029) );
  NOR4_X1 U22098 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19027) );
  AOI211_X1 U22099 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19026) );
  NOR4_X1 U22100 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19025) );
  NOR4_X1 U22101 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19024) );
  NAND4_X1 U22102 ( .A1(n19027), .A2(n19026), .A3(n19025), .A4(n19024), .ZN(
        n19028) );
  NOR2_X1 U22103 ( .A1(n19029), .A2(n19028), .ZN(n19036) );
  INV_X1 U22104 ( .A(n19036), .ZN(n19035) );
  NOR2_X1 U22105 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19035), .ZN(n19030) );
  INV_X1 U22106 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20115) );
  AOI22_X1 U22107 ( .A1(n19030), .A2(n10562), .B1(n19035), .B2(n20115), .ZN(
        P2_U2820) );
  OR3_X1 U22108 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19034) );
  INV_X1 U22109 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20113) );
  AOI22_X1 U22110 ( .A1(n19030), .A2(n19034), .B1(n19035), .B2(n20113), .ZN(
        P2_U2821) );
  INV_X1 U22111 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20118) );
  NAND2_X1 U22112 ( .A1(n19030), .A2(n20118), .ZN(n19033) );
  INV_X1 U22113 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n20056) );
  OAI21_X1 U22114 ( .B1(n10562), .B2(n20056), .A(n19036), .ZN(n19031) );
  OAI21_X1 U22115 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19036), .A(n19031), 
        .ZN(n19032) );
  OAI221_X1 U22116 ( .B1(n19033), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19033), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19032), .ZN(P2_U2822) );
  INV_X1 U22117 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20111) );
  OAI221_X1 U22118 ( .B1(n19036), .B2(n20111), .C1(n19035), .C2(n19034), .A(
        n19033), .ZN(P2_U2823) );
  AOI211_X1 U22119 ( .C1(n19042), .C2(n19038), .A(n20032), .B(n19037), .ZN(
        n19041) );
  NOR2_X1 U22120 ( .A1(n19039), .A2(n19204), .ZN(n19040) );
  NOR2_X1 U22121 ( .A1(n19041), .A2(n19040), .ZN(n19049) );
  AOI22_X1 U22122 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19252), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n19242), .ZN(n19048) );
  AOI22_X1 U22123 ( .A1(P2_EBX_REG_20__SCAN_IN), .A2(n19250), .B1(n19042), 
        .B2(n19251), .ZN(n19047) );
  OAI22_X1 U22124 ( .A1(n19044), .A2(n19207), .B1(n19043), .B2(n19246), .ZN(
        n19045) );
  INV_X1 U22125 ( .A(n19045), .ZN(n19046) );
  NAND4_X1 U22126 ( .A1(n19049), .A2(n19048), .A3(n19047), .A4(n19046), .ZN(
        P2_U2835) );
  NOR2_X1 U22127 ( .A1(n19192), .A2(n19050), .ZN(n19051) );
  XNOR2_X1 U22128 ( .A(n19052), .B(n19051), .ZN(n19061) );
  AOI22_X1 U22129 ( .A1(n19053), .A2(n19241), .B1(P2_EBX_REG_19__SCAN_IN), 
        .B2(n19250), .ZN(n19054) );
  OAI211_X1 U22130 ( .C1(n20085), .C2(n19222), .A(n19054), .B(n19176), .ZN(
        n19055) );
  AOI21_X1 U22131 ( .B1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n19252), .A(
        n19055), .ZN(n19060) );
  NOR2_X1 U22132 ( .A1(n19056), .A2(n19246), .ZN(n19057) );
  AOI21_X1 U22133 ( .B1(n19058), .B2(n19239), .A(n19057), .ZN(n19059) );
  OAI211_X1 U22134 ( .C1(n20032), .C2(n19061), .A(n19060), .B(n19059), .ZN(
        P2_U2836) );
  NAND2_X1 U22135 ( .A1(n19182), .A2(n19062), .ZN(n19073) );
  XNOR2_X1 U22136 ( .A(n19063), .B(n19073), .ZN(n19072) );
  AOI22_X1 U22137 ( .A1(P2_EBX_REG_18__SCAN_IN), .A2(n19250), .B1(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n19252), .ZN(n19064) );
  OAI21_X1 U22138 ( .B1(n19065), .B2(n19204), .A(n19064), .ZN(n19066) );
  AOI211_X1 U22139 ( .C1(P2_REIP_REG_18__SCAN_IN), .C2(n19242), .A(n19414), 
        .B(n19066), .ZN(n19071) );
  OAI22_X1 U22140 ( .A1(n19068), .A2(n19207), .B1(n19067), .B2(n19246), .ZN(
        n19069) );
  INV_X1 U22141 ( .A(n19069), .ZN(n19070) );
  OAI211_X1 U22142 ( .C1(n20032), .C2(n19072), .A(n19071), .B(n19070), .ZN(
        P2_U2837) );
  INV_X1 U22143 ( .A(n19251), .ZN(n19084) );
  INV_X1 U22144 ( .A(n19073), .ZN(n19074) );
  OAI211_X1 U22145 ( .C1(n19075), .C2(n19085), .A(n19074), .B(n19198), .ZN(
        n19077) );
  AOI22_X1 U22146 ( .A1(P2_EBX_REG_17__SCAN_IN), .A2(n19250), .B1(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n19252), .ZN(n19076) );
  OAI211_X1 U22147 ( .C1(n19204), .C2(n19078), .A(n19077), .B(n19076), .ZN(
        n19079) );
  AOI211_X1 U22148 ( .C1(P2_REIP_REG_17__SCAN_IN), .C2(n19242), .A(n19414), 
        .B(n19079), .ZN(n19083) );
  AOI22_X1 U22149 ( .A1(n19081), .A2(n19239), .B1(n19080), .B2(n19226), .ZN(
        n19082) );
  OAI211_X1 U22150 ( .C1(n19085), .C2(n19084), .A(n19083), .B(n19082), .ZN(
        P2_U2838) );
  NOR2_X1 U22151 ( .A1(n19192), .A2(n19086), .ZN(n19087) );
  XNOR2_X1 U22152 ( .A(n19088), .B(n19087), .ZN(n19096) );
  AOI22_X1 U22153 ( .A1(n19089), .A2(n19241), .B1(P2_EBX_REG_15__SCAN_IN), 
        .B2(n19250), .ZN(n19090) );
  OAI21_X1 U22154 ( .B1(n19091), .B2(n19223), .A(n19090), .ZN(n19092) );
  AOI211_X1 U22155 ( .C1(P2_REIP_REG_15__SCAN_IN), .C2(n19242), .A(n19414), 
        .B(n19092), .ZN(n19095) );
  AOI22_X1 U22156 ( .A1(n19307), .A2(n19239), .B1(n19093), .B2(n19226), .ZN(
        n19094) );
  OAI211_X1 U22157 ( .C1(n20032), .C2(n19096), .A(n19095), .B(n19094), .ZN(
        P2_U2840) );
  NAND2_X1 U22158 ( .A1(n19182), .A2(n19097), .ZN(n19098) );
  XNOR2_X1 U22159 ( .A(n19099), .B(n19098), .ZN(n19106) );
  AOI22_X1 U22160 ( .A1(n19100), .A2(n19241), .B1(P2_EBX_REG_14__SCAN_IN), 
        .B2(n19250), .ZN(n19101) );
  OAI211_X1 U22161 ( .C1(n20076), .C2(n19222), .A(n19101), .B(n19176), .ZN(
        n19102) );
  AOI21_X1 U22162 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19252), .A(
        n19102), .ZN(n19105) );
  OAI22_X1 U22163 ( .A1(n19311), .A2(n19207), .B1(n19268), .B2(n19246), .ZN(
        n19103) );
  INV_X1 U22164 ( .A(n19103), .ZN(n19104) );
  OAI211_X1 U22165 ( .C1(n20032), .C2(n19106), .A(n19105), .B(n19104), .ZN(
        P2_U2841) );
  OAI22_X1 U22166 ( .A1(n19108), .A2(n19204), .B1(n19107), .B2(n19223), .ZN(
        n19109) );
  AOI211_X1 U22167 ( .C1(P2_REIP_REG_13__SCAN_IN), .C2(n19242), .A(n19414), 
        .B(n19109), .ZN(n19117) );
  NOR2_X1 U22168 ( .A1(n19192), .A2(n19110), .ZN(n19111) );
  XNOR2_X1 U22169 ( .A(n19112), .B(n19111), .ZN(n19115) );
  OAI22_X1 U22170 ( .A1(n19313), .A2(n19207), .B1(n19113), .B2(n19246), .ZN(
        n19114) );
  AOI21_X1 U22171 ( .B1(n19115), .B2(n19198), .A(n19114), .ZN(n19116) );
  OAI211_X1 U22172 ( .C1(n19203), .C2(n19118), .A(n19117), .B(n19116), .ZN(
        P2_U2842) );
  NAND2_X1 U22173 ( .A1(n19182), .A2(n19119), .ZN(n19120) );
  XNOR2_X1 U22174 ( .A(n19121), .B(n19120), .ZN(n19127) );
  INV_X1 U22175 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n19275) );
  AOI22_X1 U22176 ( .A1(n19122), .A2(n19241), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19252), .ZN(n19123) );
  OAI21_X1 U22177 ( .B1(n19203), .B2(n19275), .A(n19123), .ZN(n19124) );
  AOI211_X1 U22178 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n19242), .A(n19414), 
        .B(n19124), .ZN(n19126) );
  AOI22_X1 U22179 ( .A1(n19271), .A2(n19226), .B1(n19314), .B2(n19239), .ZN(
        n19125) );
  OAI211_X1 U22180 ( .C1(n20032), .C2(n19127), .A(n19126), .B(n19125), .ZN(
        P2_U2843) );
  INV_X1 U22181 ( .A(n19128), .ZN(n19130) );
  OAI22_X1 U22182 ( .A1(n19130), .A2(n19204), .B1(n19203), .B2(n19129), .ZN(
        n19131) );
  AOI211_X1 U22183 ( .C1(P2_REIP_REG_11__SCAN_IN), .C2(n19242), .A(n19414), 
        .B(n19131), .ZN(n19140) );
  NOR2_X1 U22184 ( .A1(n19192), .A2(n19132), .ZN(n19133) );
  XNOR2_X1 U22185 ( .A(n19134), .B(n19133), .ZN(n19138) );
  INV_X1 U22186 ( .A(n19135), .ZN(n19136) );
  OAI22_X1 U22187 ( .A1(n19136), .A2(n19246), .B1(n19318), .B2(n19207), .ZN(
        n19137) );
  AOI21_X1 U22188 ( .B1(n19138), .B2(n19198), .A(n19137), .ZN(n19139) );
  OAI211_X1 U22189 ( .C1(n19141), .C2(n19223), .A(n19140), .B(n19139), .ZN(
        P2_U2844) );
  NAND2_X1 U22190 ( .A1(n19182), .A2(n19142), .ZN(n19144) );
  XOR2_X1 U22191 ( .A(n19144), .B(n19143), .Z(n19151) );
  AOI22_X1 U22192 ( .A1(n19145), .A2(n19241), .B1(P2_EBX_REG_10__SCAN_IN), 
        .B2(n19250), .ZN(n19146) );
  OAI211_X1 U22193 ( .C1(n20069), .C2(n19222), .A(n19146), .B(n19176), .ZN(
        n19149) );
  INV_X1 U22194 ( .A(n19277), .ZN(n19147) );
  OAI22_X1 U22195 ( .A1(n19147), .A2(n19246), .B1(n19207), .B2(n19321), .ZN(
        n19148) );
  AOI211_X1 U22196 ( .C1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n19252), .A(
        n19149), .B(n19148), .ZN(n19150) );
  OAI21_X1 U22197 ( .B1(n19151), .B2(n20032), .A(n19150), .ZN(P2_U2845) );
  INV_X1 U22198 ( .A(n19152), .ZN(n19154) );
  OAI22_X1 U22199 ( .A1(n19154), .A2(n19204), .B1(n19153), .B2(n19223), .ZN(
        n19155) );
  AOI211_X1 U22200 ( .C1(P2_REIP_REG_9__SCAN_IN), .C2(n19242), .A(n19414), .B(
        n19155), .ZN(n19164) );
  NOR2_X1 U22201 ( .A1(n19192), .A2(n19156), .ZN(n19157) );
  XNOR2_X1 U22202 ( .A(n19158), .B(n19157), .ZN(n19162) );
  INV_X1 U22203 ( .A(n19159), .ZN(n19160) );
  OAI22_X1 U22204 ( .A1(n19160), .A2(n19246), .B1(n19207), .B2(n19323), .ZN(
        n19161) );
  AOI21_X1 U22205 ( .B1(n19162), .B2(n19198), .A(n19161), .ZN(n19163) );
  OAI211_X1 U22206 ( .C1(n19203), .C2(n19165), .A(n19164), .B(n19163), .ZN(
        P2_U2846) );
  NOR2_X1 U22207 ( .A1(n19192), .A2(n19166), .ZN(n19167) );
  XOR2_X1 U22208 ( .A(n19168), .B(n19167), .Z(n19175) );
  AOI22_X1 U22209 ( .A1(n19169), .A2(n19241), .B1(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n19252), .ZN(n19170) );
  OAI211_X1 U22210 ( .C1(n20065), .C2(n19222), .A(n19170), .B(n19176), .ZN(
        n19173) );
  OAI22_X1 U22211 ( .A1(n19329), .A2(n19207), .B1(n19246), .B2(n19171), .ZN(
        n19172) );
  AOI211_X1 U22212 ( .C1(P2_EBX_REG_7__SCAN_IN), .C2(n19250), .A(n19173), .B(
        n19172), .ZN(n19174) );
  OAI21_X1 U22213 ( .B1(n20032), .B2(n19175), .A(n19174), .ZN(P2_U2848) );
  OAI21_X1 U22214 ( .B1(n20063), .B2(n19222), .A(n19176), .ZN(n19180) );
  OAI22_X1 U22215 ( .A1(n19178), .A2(n19204), .B1(n19177), .B2(n19223), .ZN(
        n19179) );
  AOI211_X1 U22216 ( .C1(P2_EBX_REG_6__SCAN_IN), .C2(n19250), .A(n19180), .B(
        n19179), .ZN(n19188) );
  NAND2_X1 U22217 ( .A1(n19182), .A2(n19181), .ZN(n19183) );
  XNOR2_X1 U22218 ( .A(n19184), .B(n19183), .ZN(n19186) );
  AOI22_X1 U22219 ( .A1(n19186), .A2(n19198), .B1(n19226), .B2(n19185), .ZN(
        n19187) );
  OAI211_X1 U22220 ( .C1(n19207), .C2(n19330), .A(n19188), .B(n19187), .ZN(
        P2_U2849) );
  OAI22_X1 U22221 ( .A1(n19204), .A2(n19189), .B1(n10181), .B2(n19223), .ZN(
        n19190) );
  AOI211_X1 U22222 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n19242), .A(n19414), .B(
        n19190), .ZN(n19201) );
  NOR2_X1 U22223 ( .A1(n19192), .A2(n19191), .ZN(n19193) );
  XNOR2_X1 U22224 ( .A(n19194), .B(n19193), .ZN(n19199) );
  INV_X1 U22225 ( .A(n19195), .ZN(n19196) );
  OAI22_X1 U22226 ( .A1(n19337), .A2(n19207), .B1(n19246), .B2(n19196), .ZN(
        n19197) );
  AOI21_X1 U22227 ( .B1(n19199), .B2(n19198), .A(n19197), .ZN(n19200) );
  OAI211_X1 U22228 ( .C1(n19203), .C2(n19202), .A(n19201), .B(n19200), .ZN(
        P2_U2850) );
  AOI22_X1 U22229 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n19250), .B1(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n19252), .ZN(n19220) );
  INV_X1 U22230 ( .A(n19339), .ZN(n19206) );
  OAI22_X1 U22231 ( .A1(n19207), .A2(n19206), .B1(n19205), .B2(n19204), .ZN(
        n19208) );
  AOI211_X1 U22232 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n19242), .A(n19414), .B(
        n19208), .ZN(n19219) );
  OR2_X1 U22233 ( .A1(n19209), .A2(n19210), .ZN(n19211) );
  NAND2_X1 U22234 ( .A1(n19212), .A2(n19211), .ZN(n19341) );
  OAI22_X1 U22235 ( .A1(n19341), .A2(n19247), .B1(n19246), .B2(n19415), .ZN(
        n19213) );
  INV_X1 U22236 ( .A(n19213), .ZN(n19218) );
  AND2_X1 U22237 ( .A1(n19182), .A2(n19214), .ZN(n19216) );
  AOI21_X1 U22238 ( .B1(n19412), .B2(n19216), .A(n20032), .ZN(n19215) );
  OAI21_X1 U22239 ( .B1(n19412), .B2(n19216), .A(n19215), .ZN(n19217) );
  NAND4_X1 U22240 ( .A1(n19220), .A2(n19219), .A3(n19218), .A4(n19217), .ZN(
        P2_U2851) );
  NAND2_X1 U22241 ( .A1(n19250), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n19231) );
  INV_X1 U22242 ( .A(n19221), .ZN(n19225) );
  OAI22_X1 U22243 ( .A1(n19233), .A2(n19223), .B1(n20056), .B2(n19222), .ZN(
        n19224) );
  AOI21_X1 U22244 ( .B1(n19241), .B2(n19225), .A(n19224), .ZN(n19230) );
  NAND2_X1 U22245 ( .A1(n19227), .A2(n19226), .ZN(n19229) );
  NAND2_X1 U22246 ( .A1(n19239), .A2(n20154), .ZN(n19228) );
  AND4_X1 U22247 ( .A1(n19231), .A2(n19230), .A3(n19229), .A4(n19228), .ZN(
        n19235) );
  AOI22_X1 U22248 ( .A1(n19251), .A2(n19233), .B1(n20152), .B2(n19232), .ZN(
        n19234) );
  OAI211_X1 U22249 ( .C1(n20032), .C2(n19236), .A(n19235), .B(n19234), .ZN(
        P2_U2854) );
  INV_X1 U22250 ( .A(n19237), .ZN(n19238) );
  AOI22_X1 U22251 ( .A1(n19241), .A2(n19240), .B1(n19239), .B2(n19238), .ZN(
        n19244) );
  NAND2_X1 U22252 ( .A1(n19242), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n19243) );
  OAI211_X1 U22253 ( .C1(n19246), .C2(n19245), .A(n19244), .B(n19243), .ZN(
        n19249) );
  NOR2_X1 U22254 ( .A1(n20160), .A2(n19247), .ZN(n19248) );
  AOI211_X1 U22255 ( .C1(P2_EBX_REG_0__SCAN_IN), .C2(n19250), .A(n19249), .B(
        n19248), .ZN(n19254) );
  OAI21_X1 U22256 ( .B1(n19252), .B2(n19251), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19253) );
  OAI211_X1 U22257 ( .C1(n19256), .C2(n19255), .A(n19254), .B(n19253), .ZN(
        P2_U2855) );
  AND2_X1 U22258 ( .A1(n14174), .A2(n19257), .ZN(n19258) );
  OR2_X1 U22259 ( .A1(n19258), .A2(n15014), .ZN(n19301) );
  INV_X1 U22260 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n19259) );
  OAI22_X1 U22261 ( .A1(n19301), .A2(n19289), .B1(n19293), .B2(n19259), .ZN(
        n19260) );
  INV_X1 U22262 ( .A(n19260), .ZN(n19261) );
  OAI21_X1 U22263 ( .B1(n14945), .B2(n19262), .A(n19261), .ZN(P2_U2871) );
  AOI21_X1 U22264 ( .B1(n14096), .B2(n19264), .A(n19263), .ZN(n19265) );
  NOR3_X1 U22265 ( .A1(n9949), .A2(n19265), .A3(n19289), .ZN(n19266) );
  AOI21_X1 U22266 ( .B1(P2_EBX_REG_14__SCAN_IN), .B2(n14945), .A(n19266), .ZN(
        n19267) );
  OAI21_X1 U22267 ( .B1(n19268), .B2(n14945), .A(n19267), .ZN(P2_U2873) );
  OAI21_X1 U22268 ( .B1(n14003), .B2(n19269), .A(n19278), .ZN(n19270) );
  OR2_X1 U22269 ( .A1(n19270), .A2(n14096), .ZN(n19273) );
  NAND2_X1 U22270 ( .A1(n19271), .A2(n19293), .ZN(n19272) );
  AND2_X1 U22271 ( .A1(n19273), .A2(n19272), .ZN(n19274) );
  OAI21_X1 U22272 ( .B1(n19293), .B2(n19275), .A(n19274), .ZN(P2_U2875) );
  XNOR2_X1 U22273 ( .A(n13975), .B(n19276), .ZN(n19279) );
  AOI22_X1 U22274 ( .A1(n19279), .A2(n19278), .B1(n19293), .B2(n19277), .ZN(
        n19280) );
  OAI21_X1 U22275 ( .B1(n19293), .B2(n19281), .A(n19280), .ZN(P2_U2877) );
  AOI211_X1 U22276 ( .C1(n19285), .C2(n9969), .A(n19289), .B(n19284), .ZN(
        n19286) );
  AOI21_X1 U22277 ( .B1(P2_EBX_REG_8__SCAN_IN), .B2(n14945), .A(n19286), .ZN(
        n19287) );
  OAI21_X1 U22278 ( .B1(n19288), .B2(n14945), .A(n19287), .ZN(P2_U2879) );
  OAI22_X1 U22279 ( .A1(n19341), .A2(n19289), .B1(n14945), .B2(n19415), .ZN(
        n19290) );
  INV_X1 U22280 ( .A(n19290), .ZN(n19291) );
  OAI21_X1 U22281 ( .B1(n19293), .B2(n19292), .A(n19291), .ZN(P2_U2883) );
  AOI22_X1 U22282 ( .A1(n19300), .A2(BUF2_REG_31__SCAN_IN), .B1(n19294), .B2(
        n19357), .ZN(n19296) );
  AOI22_X1 U22283 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19356), .B1(n19299), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19295) );
  NAND2_X1 U22284 ( .A1(n19296), .A2(n19295), .ZN(P2_U2888) );
  AOI22_X1 U22285 ( .A1(n19298), .A2(n19297), .B1(n19356), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n19306) );
  AOI22_X1 U22286 ( .A1(n19300), .A2(BUF2_REG_16__SCAN_IN), .B1(n19299), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n19305) );
  OAI22_X1 U22287 ( .A1(n19302), .A2(n19348), .B1(n19361), .B2(n19301), .ZN(
        n19303) );
  INV_X1 U22288 ( .A(n19303), .ZN(n19304) );
  NAND3_X1 U22289 ( .A1(n19306), .A2(n19305), .A3(n19304), .ZN(P2_U2903) );
  INV_X1 U22290 ( .A(n19307), .ZN(n19309) );
  OAI222_X1 U22291 ( .A1(n19309), .A2(n19338), .B1(n13451), .B2(n19347), .C1(
        n19308), .C2(n19365), .ZN(P2_U2904) );
  AOI22_X1 U22292 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19356), .B1(n19406), 
        .B2(n19325), .ZN(n19310) );
  OAI21_X1 U22293 ( .B1(n19338), .B2(n19311), .A(n19310), .ZN(P2_U2905) );
  INV_X1 U22294 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19377) );
  OAI222_X1 U22295 ( .A1(n19313), .A2(n19338), .B1(n19377), .B2(n19347), .C1(
        n19365), .C2(n19312), .ZN(P2_U2906) );
  INV_X1 U22296 ( .A(n19314), .ZN(n19316) );
  INV_X1 U22297 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19379) );
  OAI222_X1 U22298 ( .A1(n19316), .A2(n19338), .B1(n19379), .B2(n19347), .C1(
        n19365), .C2(n19315), .ZN(P2_U2907) );
  INV_X1 U22299 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19381) );
  OAI222_X1 U22300 ( .A1(n19318), .A2(n19338), .B1(n19381), .B2(n19347), .C1(
        n19365), .C2(n19317), .ZN(P2_U2908) );
  AOI22_X1 U22301 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19356), .B1(n19319), 
        .B2(n19325), .ZN(n19320) );
  OAI21_X1 U22302 ( .B1(n19338), .B2(n19321), .A(n19320), .ZN(P2_U2909) );
  INV_X1 U22303 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19384) );
  OAI222_X1 U22304 ( .A1(n19323), .A2(n19338), .B1(n19384), .B2(n19347), .C1(
        n19365), .C2(n19322), .ZN(P2_U2910) );
  INV_X1 U22305 ( .A(n19324), .ZN(n19328) );
  AOI22_X1 U22306 ( .A1(P2_EAX_REG_8__SCAN_IN), .A2(n19356), .B1(n19326), .B2(
        n19325), .ZN(n19327) );
  OAI21_X1 U22307 ( .B1(n19338), .B2(n19328), .A(n19327), .ZN(P2_U2911) );
  OAI222_X1 U22308 ( .A1(n19329), .A2(n19338), .B1(n19388), .B2(n19347), .C1(
        n19365), .C2(n19488), .ZN(P2_U2912) );
  INV_X1 U22309 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19390) );
  OAI222_X1 U22310 ( .A1(n19330), .A2(n19338), .B1(n19390), .B2(n19347), .C1(
        n19365), .C2(n19476), .ZN(P2_U2913) );
  INV_X1 U22311 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19392) );
  OAI22_X1 U22312 ( .A1(n19392), .A2(n19347), .B1(n19471), .B2(n19365), .ZN(
        n19331) );
  INV_X1 U22313 ( .A(n19331), .ZN(n19336) );
  AOI21_X1 U22314 ( .B1(n19333), .B2(n20143), .A(n19332), .ZN(n19352) );
  XNOR2_X1 U22315 ( .A(n20122), .B(n20137), .ZN(n19351) );
  NOR2_X1 U22316 ( .A1(n19352), .A2(n19351), .ZN(n19350) );
  AOI21_X1 U22317 ( .B1(n20122), .B2(n20137), .A(n19350), .ZN(n19334) );
  NOR2_X1 U22318 ( .A1(n19334), .A2(n19339), .ZN(n19340) );
  OR3_X1 U22319 ( .A1(n19340), .A2(n19341), .A3(n19361), .ZN(n19335) );
  OAI211_X1 U22320 ( .C1(n19338), .C2(n19337), .A(n19336), .B(n19335), .ZN(
        P2_U2914) );
  AOI22_X1 U22321 ( .A1(n19357), .A2(n19339), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19356), .ZN(n19345) );
  XOR2_X1 U22322 ( .A(n19341), .B(n19340), .Z(n19343) );
  NAND2_X1 U22323 ( .A1(n19343), .A2(n19342), .ZN(n19344) );
  OAI211_X1 U22324 ( .C1(n19465), .C2(n19365), .A(n19345), .B(n19344), .ZN(
        P2_U2915) );
  INV_X1 U22325 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19346) );
  OAI22_X1 U22326 ( .A1(n20137), .A2(n19348), .B1(n19347), .B2(n19346), .ZN(
        n19349) );
  INV_X1 U22327 ( .A(n19349), .ZN(n19355) );
  AOI21_X1 U22328 ( .B1(n19352), .B2(n19351), .A(n19350), .ZN(n19353) );
  OR2_X1 U22329 ( .A1(n19353), .A2(n19361), .ZN(n19354) );
  OAI211_X1 U22330 ( .C1(n19459), .C2(n19365), .A(n19355), .B(n19354), .ZN(
        P2_U2916) );
  AOI22_X1 U22331 ( .A1(n19357), .A2(n20154), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19356), .ZN(n19364) );
  AOI21_X1 U22332 ( .B1(n19360), .B2(n19359), .A(n19358), .ZN(n19362) );
  OR2_X1 U22333 ( .A1(n19362), .A2(n19361), .ZN(n19363) );
  OAI211_X1 U22334 ( .C1(n19448), .C2(n19365), .A(n19364), .B(n19363), .ZN(
        P2_U2918) );
  NOR2_X1 U22335 ( .A1(n19370), .A2(n19366), .ZN(P2_U2920) );
  INV_X1 U22336 ( .A(n19367), .ZN(n19368) );
  AOI22_X1 U22337 ( .A1(n19368), .A2(P2_EAX_REG_30__SCAN_IN), .B1(
        P2_UWORD_REG_14__SCAN_IN), .B2(n19402), .ZN(n19369) );
  OAI21_X1 U22338 ( .B1(n19371), .B2(n19370), .A(n19369), .ZN(P2_U2921) );
  AOI22_X1 U22339 ( .A1(n19402), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19396), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19373) );
  OAI21_X1 U22340 ( .B1(n13451), .B2(n19404), .A(n19373), .ZN(P2_U2936) );
  INV_X1 U22341 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19375) );
  AOI22_X1 U22342 ( .A1(n19402), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19396), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19374) );
  OAI21_X1 U22343 ( .B1(n19375), .B2(n19404), .A(n19374), .ZN(P2_U2937) );
  AOI22_X1 U22344 ( .A1(n19402), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19396), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19376) );
  OAI21_X1 U22345 ( .B1(n19377), .B2(n19404), .A(n19376), .ZN(P2_U2938) );
  AOI22_X1 U22346 ( .A1(n19402), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19396), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19378) );
  OAI21_X1 U22347 ( .B1(n19379), .B2(n19404), .A(n19378), .ZN(P2_U2939) );
  AOI22_X1 U22348 ( .A1(n19397), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19396), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19380) );
  OAI21_X1 U22349 ( .B1(n19381), .B2(n19404), .A(n19380), .ZN(P2_U2940) );
  AOI22_X1 U22350 ( .A1(n19397), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19396), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19382) );
  OAI21_X1 U22351 ( .B1(n11298), .B2(n19404), .A(n19382), .ZN(P2_U2941) );
  AOI22_X1 U22352 ( .A1(n19397), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19396), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19383) );
  OAI21_X1 U22353 ( .B1(n19384), .B2(n19404), .A(n19383), .ZN(P2_U2942) );
  AOI22_X1 U22354 ( .A1(n19397), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19396), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19385) );
  OAI21_X1 U22355 ( .B1(n19386), .B2(n19404), .A(n19385), .ZN(P2_U2943) );
  AOI22_X1 U22356 ( .A1(n19397), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19396), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19387) );
  OAI21_X1 U22357 ( .B1(n19388), .B2(n19404), .A(n19387), .ZN(P2_U2944) );
  AOI22_X1 U22358 ( .A1(n19397), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19396), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19389) );
  OAI21_X1 U22359 ( .B1(n19390), .B2(n19404), .A(n19389), .ZN(P2_U2945) );
  AOI22_X1 U22360 ( .A1(n19397), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19396), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19391) );
  OAI21_X1 U22361 ( .B1(n19392), .B2(n19404), .A(n19391), .ZN(P2_U2946) );
  INV_X1 U22362 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19394) );
  AOI22_X1 U22363 ( .A1(n19397), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19396), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19393) );
  OAI21_X1 U22364 ( .B1(n19394), .B2(n19404), .A(n19393), .ZN(P2_U2947) );
  AOI22_X1 U22365 ( .A1(n19397), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19396), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19395) );
  OAI21_X1 U22366 ( .B1(n19346), .B2(n19404), .A(n19395), .ZN(P2_U2948) );
  INV_X1 U22367 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19399) );
  AOI22_X1 U22368 ( .A1(n19397), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19396), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19398) );
  OAI21_X1 U22369 ( .B1(n19399), .B2(n19404), .A(n19398), .ZN(P2_U2949) );
  INV_X1 U22370 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19401) );
  AOI22_X1 U22371 ( .A1(n19402), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19396), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19400) );
  OAI21_X1 U22372 ( .B1(n19401), .B2(n19404), .A(n19400), .ZN(P2_U2950) );
  AOI22_X1 U22373 ( .A1(n19402), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19396), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19403) );
  OAI21_X1 U22374 ( .B1(n13682), .B2(n19404), .A(n19403), .ZN(P2_U2951) );
  AOI22_X1 U22375 ( .A1(P2_UWORD_REG_14__SCAN_IN), .A2(n19405), .B1(n19409), 
        .B2(P2_EAX_REG_30__SCAN_IN), .ZN(n19408) );
  NAND2_X1 U22376 ( .A1(n19407), .A2(n19406), .ZN(n19410) );
  NAND2_X1 U22377 ( .A1(n19408), .A2(n19410), .ZN(P2_U2966) );
  AOI22_X1 U22378 ( .A1(P2_LWORD_REG_14__SCAN_IN), .A2(n19405), .B1(n19409), 
        .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n19411) );
  NAND2_X1 U22379 ( .A1(n19411), .A2(n19410), .ZN(P2_U2981) );
  AOI22_X1 U22380 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19414), .B1(n19413), 
        .B2(n19412), .ZN(n19423) );
  OAI22_X1 U22381 ( .A1(n19418), .A2(n19417), .B1(n19416), .B2(n19415), .ZN(
        n19419) );
  AOI21_X1 U22382 ( .B1(n19421), .B2(n19420), .A(n19419), .ZN(n19422) );
  OAI211_X1 U22383 ( .C1(n19425), .C2(n19424), .A(n19423), .B(n19422), .ZN(
        P2_U3010) );
  NAND2_X1 U22384 ( .A1(n20126), .A2(n19528), .ZN(n19426) );
  NAND2_X1 U22385 ( .A1(n20126), .A2(n19612), .ZN(n19922) );
  NAND2_X1 U22386 ( .A1(n19427), .A2(n19922), .ZN(n19439) );
  INV_X1 U22387 ( .A(n20017), .ZN(n19428) );
  NAND2_X1 U22388 ( .A1(n19439), .A2(n19428), .ZN(n19431) );
  NAND2_X1 U22389 ( .A1(n19440), .A2(n20136), .ZN(n19429) );
  INV_X1 U22390 ( .A(n20126), .ZN(n19765) );
  NAND2_X1 U22391 ( .A1(n19429), .A2(n19765), .ZN(n19430) );
  NAND2_X1 U22392 ( .A1(n19431), .A2(n19430), .ZN(n19433) );
  NAND2_X1 U22393 ( .A1(n20140), .A2(n20147), .ZN(n19577) );
  OR2_X1 U22394 ( .A1(n19577), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19502) );
  NOR2_X1 U22395 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19502), .ZN(
        n19486) );
  INV_X1 U22396 ( .A(n19486), .ZN(n19432) );
  NAND2_X1 U22397 ( .A1(n19433), .A2(n19432), .ZN(n19434) );
  AOI22_X1 U22398 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19481), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19480), .ZN(n19979) );
  INV_X1 U22399 ( .A(n19979), .ZN(n19929) );
  NAND2_X1 U22400 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19974), .ZN(n19475) );
  INV_X1 U22401 ( .A(n19475), .ZN(n19485) );
  AND2_X1 U22402 ( .A1(n19437), .A2(n19485), .ZN(n19967) );
  AOI22_X1 U22403 ( .A1(n19929), .A2(n20021), .B1(n19967), .B2(n19486), .ZN(
        n19445) );
  NOR2_X2 U22404 ( .A1(n19438), .A2(n19673), .ZN(n19968) );
  OAI21_X1 U22405 ( .B1(n20017), .B2(n19486), .A(n19439), .ZN(n19442) );
  OAI21_X1 U22406 ( .B1(n19440), .B2(n19486), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19441) );
  NAND2_X1 U22407 ( .A1(n19442), .A2(n19441), .ZN(n19489) );
  OAI22_X2 U22408 ( .A1(n20375), .A2(n19484), .B1(n19443), .B2(n19482), .ZN(
        n19976) );
  AOI22_X1 U22409 ( .A1(n19968), .A2(n19489), .B1(n19544), .B2(n19976), .ZN(
        n19444) );
  OAI211_X1 U22410 ( .C1(n19487), .C2(n19446), .A(n19445), .B(n19444), .ZN(
        P2_U3048) );
  AOI22_X1 U22411 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19481), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19480), .ZN(n19985) );
  INV_X1 U22412 ( .A(n19985), .ZN(n19937) );
  AOI22_X1 U22413 ( .A1(n19937), .A2(n20021), .B1(n19980), .B2(n19486), .ZN(
        n19451) );
  NOR2_X2 U22414 ( .A1(n19448), .A2(n19673), .ZN(n19981) );
  OAI22_X2 U22415 ( .A1(n20394), .A2(n19484), .B1(n19449), .B2(n19482), .ZN(
        n19982) );
  AOI22_X1 U22416 ( .A1(n19981), .A2(n19489), .B1(n19544), .B2(n19982), .ZN(
        n19450) );
  OAI211_X1 U22417 ( .C1(n19487), .C2(n19452), .A(n19451), .B(n19450), .ZN(
        P2_U3049) );
  AOI22_X2 U22418 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19481), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19480), .ZN(n19991) );
  INV_X1 U22419 ( .A(n19991), .ZN(n19941) );
  NOR2_X2 U22420 ( .A1(n10502), .A2(n19475), .ZN(n19986) );
  AOI22_X1 U22421 ( .A1(n19941), .A2(n20021), .B1(n19986), .B2(n19486), .ZN(
        n19456) );
  NOR2_X2 U22422 ( .A1(n19453), .A2(n19673), .ZN(n19987) );
  OAI22_X2 U22423 ( .A1(n20401), .A2(n19484), .B1(n19454), .B2(n19482), .ZN(
        n19988) );
  AOI22_X1 U22424 ( .A1(n19987), .A2(n19489), .B1(n19544), .B2(n19988), .ZN(
        n19455) );
  OAI211_X1 U22425 ( .C1(n19487), .C2(n19457), .A(n19456), .B(n19455), .ZN(
        P2_U3050) );
  AOI22_X1 U22426 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19481), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19480), .ZN(n19997) );
  INV_X1 U22427 ( .A(n19997), .ZN(n19944) );
  AOI22_X1 U22428 ( .A1(n19944), .A2(n20021), .B1(n19992), .B2(n19486), .ZN(
        n19461) );
  NOR2_X2 U22429 ( .A1(n19459), .A2(n19673), .ZN(n19993) );
  AOI22_X1 U22430 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19481), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19480), .ZN(n19782) );
  AOI22_X1 U22431 ( .A1(n19993), .A2(n19489), .B1(n19544), .B2(n19994), .ZN(
        n19460) );
  OAI211_X1 U22432 ( .C1(n19487), .C2(n19462), .A(n19461), .B(n19460), .ZN(
        P2_U3051) );
  OR2_X1 U22433 ( .A1(n19464), .A2(n19475), .ZN(n19523) );
  AOI22_X1 U22434 ( .A1(n19947), .A2(n20021), .B1(n19998), .B2(n19486), .ZN(
        n19467) );
  NOR2_X2 U22435 ( .A1(n19465), .A2(n19673), .ZN(n19999) );
  AOI22_X1 U22436 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19481), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19480), .ZN(n19814) );
  INV_X1 U22437 ( .A(n19814), .ZN(n20000) );
  AOI22_X1 U22438 ( .A1(n19999), .A2(n19489), .B1(n19544), .B2(n20000), .ZN(
        n19466) );
  OAI211_X1 U22439 ( .C1(n19487), .C2(n19468), .A(n19467), .B(n19466), .ZN(
        P2_U3052) );
  NOR2_X2 U22440 ( .A1(n19470), .A2(n19475), .ZN(n20004) );
  AOI22_X1 U22441 ( .A1(n19950), .A2(n20021), .B1(n20004), .B2(n19486), .ZN(
        n19473) );
  NOR2_X2 U22442 ( .A1(n19471), .A2(n19673), .ZN(n20005) );
  AOI22_X1 U22443 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19481), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19480), .ZN(n19817) );
  AOI22_X1 U22444 ( .A1(n20005), .A2(n19489), .B1(n19544), .B2(n20006), .ZN(
        n19472) );
  OAI211_X1 U22445 ( .C1(n19487), .C2(n13871), .A(n19473), .B(n19472), .ZN(
        P2_U3053) );
  NOR2_X2 U22446 ( .A1(n13076), .A2(n19475), .ZN(n20010) );
  AOI22_X1 U22447 ( .A1(n19954), .A2(n20021), .B1(n20010), .B2(n19486), .ZN(
        n19478) );
  NOR2_X2 U22448 ( .A1(n19476), .A2(n19673), .ZN(n20011) );
  AOI22_X1 U22449 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19481), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19480), .ZN(n19820) );
  AOI22_X1 U22450 ( .A1(n20011), .A2(n19489), .B1(n19544), .B2(n20012), .ZN(
        n19477) );
  OAI211_X1 U22451 ( .C1(n19487), .C2(n19479), .A(n19478), .B(n19477), .ZN(
        P2_U3054) );
  AOI22_X1 U22452 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19481), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19480), .ZN(n19827) );
  AOI22_X1 U22453 ( .A1(n19958), .A2(n20021), .B1(n20016), .B2(n19486), .ZN(
        n19492) );
  INV_X1 U22454 ( .A(n19487), .ZN(n19490) );
  NOR2_X2 U22455 ( .A1(n19488), .A2(n19673), .ZN(n20018) );
  AOI22_X1 U22456 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19490), .B1(
        n20018), .B2(n19489), .ZN(n19491) );
  OAI211_X1 U22457 ( .C1(n19827), .C2(n19528), .A(n19492), .B(n19491), .ZN(
        P2_U3055) );
  INV_X1 U22458 ( .A(n19764), .ZN(n19500) );
  NOR2_X1 U22459 ( .A1(n19763), .A2(n19577), .ZN(n19505) );
  INV_X1 U22460 ( .A(n19505), .ZN(n19539) );
  NAND2_X1 U22461 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19539), .ZN(n19493) );
  NOR2_X1 U22462 ( .A1(n19494), .A2(n19493), .ZN(n19501) );
  INV_X1 U22463 ( .A(n19502), .ZN(n19495) );
  AOI21_X1 U22464 ( .B1(n20136), .B2(n19495), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19496) );
  INV_X1 U22465 ( .A(n19968), .ZN(n19498) );
  INV_X1 U22466 ( .A(n19967), .ZN(n19497) );
  OAI22_X1 U22467 ( .A1(n19542), .A2(n19498), .B1(n19497), .B2(n19539), .ZN(
        n19499) );
  INV_X1 U22468 ( .A(n19499), .ZN(n19507) );
  AND2_X1 U22469 ( .A1(n20122), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19698) );
  NAND2_X1 U22470 ( .A1(n19698), .A2(n19500), .ZN(n19503) );
  AOI21_X1 U22471 ( .B1(n19503), .B2(n19502), .A(n19501), .ZN(n19504) );
  OAI211_X1 U22472 ( .C1(n19505), .C2(n20136), .A(n19504), .B(n19974), .ZN(
        n19545) );
  AOI22_X1 U22473 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19545), .B1(
        n19544), .B2(n19929), .ZN(n19506) );
  OAI211_X1 U22474 ( .C1(n19839), .C2(n19563), .A(n19507), .B(n19506), .ZN(
        P2_U3056) );
  INV_X1 U22475 ( .A(n19981), .ZN(n19509) );
  INV_X1 U22476 ( .A(n19980), .ZN(n19508) );
  OAI22_X1 U22477 ( .A1(n19542), .A2(n19509), .B1(n19508), .B2(n19539), .ZN(
        n19510) );
  INV_X1 U22478 ( .A(n19510), .ZN(n19512) );
  AOI22_X1 U22479 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19545), .B1(
        n19572), .B2(n19982), .ZN(n19511) );
  OAI211_X1 U22480 ( .C1(n19985), .C2(n19528), .A(n19512), .B(n19511), .ZN(
        P2_U3057) );
  INV_X1 U22481 ( .A(n19987), .ZN(n19514) );
  INV_X1 U22482 ( .A(n19986), .ZN(n19513) );
  OAI22_X1 U22483 ( .A1(n19542), .A2(n19514), .B1(n19513), .B2(n19539), .ZN(
        n19515) );
  INV_X1 U22484 ( .A(n19515), .ZN(n19517) );
  AOI22_X1 U22485 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19545), .B1(
        n19572), .B2(n19988), .ZN(n19516) );
  OAI211_X1 U22486 ( .C1(n19991), .C2(n19528), .A(n19517), .B(n19516), .ZN(
        P2_U3058) );
  INV_X1 U22487 ( .A(n19993), .ZN(n19519) );
  INV_X1 U22488 ( .A(n19992), .ZN(n19518) );
  OAI22_X1 U22489 ( .A1(n19542), .A2(n19519), .B1(n19518), .B2(n19539), .ZN(
        n19520) );
  INV_X1 U22490 ( .A(n19520), .ZN(n19522) );
  AOI22_X1 U22491 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19545), .B1(
        n19572), .B2(n19994), .ZN(n19521) );
  OAI211_X1 U22492 ( .C1(n19997), .C2(n19528), .A(n19522), .B(n19521), .ZN(
        P2_U3059) );
  INV_X1 U22493 ( .A(n19999), .ZN(n19524) );
  OAI22_X1 U22494 ( .A1(n19542), .A2(n19524), .B1(n19523), .B2(n19539), .ZN(
        n19525) );
  INV_X1 U22495 ( .A(n19525), .ZN(n19527) );
  AOI22_X1 U22496 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19545), .B1(
        n19572), .B2(n20000), .ZN(n19526) );
  OAI211_X1 U22497 ( .C1(n20003), .C2(n19528), .A(n19527), .B(n19526), .ZN(
        P2_U3060) );
  INV_X1 U22498 ( .A(n20005), .ZN(n19530) );
  INV_X1 U22499 ( .A(n20004), .ZN(n19529) );
  OAI22_X1 U22500 ( .A1(n19542), .A2(n19530), .B1(n19529), .B2(n19539), .ZN(
        n19531) );
  INV_X1 U22501 ( .A(n19531), .ZN(n19533) );
  AOI22_X1 U22502 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19545), .B1(
        n19544), .B2(n19950), .ZN(n19532) );
  OAI211_X1 U22503 ( .C1(n19817), .C2(n19563), .A(n19533), .B(n19532), .ZN(
        P2_U3061) );
  INV_X1 U22504 ( .A(n20011), .ZN(n19535) );
  INV_X1 U22505 ( .A(n20010), .ZN(n19534) );
  OAI22_X1 U22506 ( .A1(n19542), .A2(n19535), .B1(n19534), .B2(n19539), .ZN(
        n19536) );
  INV_X1 U22507 ( .A(n19536), .ZN(n19538) );
  AOI22_X1 U22508 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19545), .B1(
        n19544), .B2(n19954), .ZN(n19537) );
  OAI211_X1 U22509 ( .C1(n19820), .C2(n19563), .A(n19538), .B(n19537), .ZN(
        P2_U3062) );
  INV_X1 U22510 ( .A(n20018), .ZN(n19541) );
  INV_X1 U22511 ( .A(n20016), .ZN(n19540) );
  OAI22_X1 U22512 ( .A1(n19542), .A2(n19541), .B1(n19540), .B2(n19539), .ZN(
        n19543) );
  INV_X1 U22513 ( .A(n19543), .ZN(n19547) );
  AOI22_X1 U22514 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19545), .B1(
        n19544), .B2(n19958), .ZN(n19546) );
  OAI211_X1 U22515 ( .C1(n19827), .C2(n19563), .A(n19547), .B(n19546), .ZN(
        P2_U3063) );
  NOR2_X1 U22516 ( .A1(n19795), .A2(n19577), .ZN(n19570) );
  OAI21_X1 U22517 ( .B1(n10703), .B2(n19570), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19549) );
  NOR2_X1 U22518 ( .A1(n19797), .A2(n19577), .ZN(n19550) );
  INV_X1 U22519 ( .A(n19550), .ZN(n19548) );
  NAND2_X1 U22520 ( .A1(n19549), .A2(n19548), .ZN(n19571) );
  AOI22_X1 U22521 ( .A1(n19571), .A2(n19968), .B1(n19967), .B2(n19570), .ZN(
        n19556) );
  NAND2_X1 U22522 ( .A1(n19606), .A2(n19563), .ZN(n19551) );
  AOI21_X1 U22523 ( .B1(n19551), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19550), 
        .ZN(n19553) );
  AOI21_X1 U22524 ( .B1(n10703), .B2(n20136), .A(n19570), .ZN(n19552) );
  MUX2_X1 U22525 ( .A(n19553), .B(n19552), .S(n19765), .Z(n19554) );
  AOI22_X1 U22526 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19573), .B1(
        n19592), .B2(n19976), .ZN(n19555) );
  OAI211_X1 U22527 ( .C1(n19979), .C2(n19563), .A(n19556), .B(n19555), .ZN(
        P2_U3064) );
  AOI22_X1 U22528 ( .A1(n19571), .A2(n19981), .B1(n19980), .B2(n19570), .ZN(
        n19558) );
  AOI22_X1 U22529 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19573), .B1(
        n19592), .B2(n19982), .ZN(n19557) );
  OAI211_X1 U22530 ( .C1(n19985), .C2(n19563), .A(n19558), .B(n19557), .ZN(
        P2_U3065) );
  AOI22_X1 U22531 ( .A1(n19571), .A2(n19987), .B1(n19986), .B2(n19570), .ZN(
        n19560) );
  AOI22_X1 U22532 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19573), .B1(
        n19592), .B2(n19988), .ZN(n19559) );
  OAI211_X1 U22533 ( .C1(n19991), .C2(n19563), .A(n19560), .B(n19559), .ZN(
        P2_U3066) );
  AOI22_X1 U22534 ( .A1(n19571), .A2(n19993), .B1(n19992), .B2(n19570), .ZN(
        n19562) );
  AOI22_X1 U22535 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19573), .B1(
        n19592), .B2(n19994), .ZN(n19561) );
  OAI211_X1 U22536 ( .C1(n19997), .C2(n19563), .A(n19562), .B(n19561), .ZN(
        P2_U3067) );
  AOI22_X1 U22537 ( .A1(n19571), .A2(n19999), .B1(n19998), .B2(n19570), .ZN(
        n19565) );
  AOI22_X1 U22538 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19573), .B1(
        n19572), .B2(n19947), .ZN(n19564) );
  OAI211_X1 U22539 ( .C1(n19814), .C2(n19606), .A(n19565), .B(n19564), .ZN(
        P2_U3068) );
  AOI22_X1 U22540 ( .A1(n19571), .A2(n20005), .B1(n20004), .B2(n19570), .ZN(
        n19567) );
  AOI22_X1 U22541 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19573), .B1(
        n19572), .B2(n19950), .ZN(n19566) );
  OAI211_X1 U22542 ( .C1(n19817), .C2(n19606), .A(n19567), .B(n19566), .ZN(
        P2_U3069) );
  AOI22_X1 U22543 ( .A1(n19571), .A2(n20011), .B1(n20010), .B2(n19570), .ZN(
        n19569) );
  AOI22_X1 U22544 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19573), .B1(
        n19572), .B2(n19954), .ZN(n19568) );
  OAI211_X1 U22545 ( .C1(n19820), .C2(n19606), .A(n19569), .B(n19568), .ZN(
        P2_U3070) );
  AOI22_X1 U22546 ( .A1(n19571), .A2(n20018), .B1(n20016), .B2(n19570), .ZN(
        n19575) );
  AOI22_X1 U22547 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19573), .B1(
        n19572), .B2(n19958), .ZN(n19574) );
  OAI211_X1 U22548 ( .C1(n19827), .C2(n19606), .A(n19575), .B(n19574), .ZN(
        P2_U3071) );
  INV_X1 U22549 ( .A(n19576), .ZN(n19709) );
  NOR2_X1 U22550 ( .A1(n19829), .A2(n19577), .ZN(n19601) );
  AOI22_X1 U22551 ( .A1(n19628), .A2(n19976), .B1(n19601), .B2(n19967), .ZN(
        n19587) );
  INV_X1 U22552 ( .A(n19698), .ZN(n19639) );
  OAI21_X1 U22553 ( .B1(n19639), .B2(n20127), .A(n20126), .ZN(n19585) );
  NOR2_X1 U22554 ( .A1(n16450), .A2(n19577), .ZN(n19581) );
  INV_X1 U22555 ( .A(n19582), .ZN(n19579) );
  INV_X1 U22556 ( .A(n19601), .ZN(n19578) );
  OAI211_X1 U22557 ( .C1(n19579), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19578), 
        .B(n19765), .ZN(n19580) );
  OAI211_X1 U22558 ( .C1(n19585), .C2(n19581), .A(n19974), .B(n19580), .ZN(
        n19603) );
  INV_X1 U22559 ( .A(n19581), .ZN(n19584) );
  OAI21_X1 U22560 ( .B1(n19582), .B2(n19601), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19583) );
  OAI21_X1 U22561 ( .B1(n19585), .B2(n19584), .A(n19583), .ZN(n19602) );
  AOI22_X1 U22562 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19603), .B1(
        n19968), .B2(n19602), .ZN(n19586) );
  OAI211_X1 U22563 ( .C1(n19979), .C2(n19606), .A(n19587), .B(n19586), .ZN(
        P2_U3072) );
  INV_X1 U22564 ( .A(n19982), .ZN(n19843) );
  AOI22_X1 U22565 ( .A1(n19937), .A2(n19592), .B1(n19601), .B2(n19980), .ZN(
        n19589) );
  AOI22_X1 U22566 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19603), .B1(
        n19981), .B2(n19602), .ZN(n19588) );
  OAI211_X1 U22567 ( .C1(n19843), .C2(n19638), .A(n19589), .B(n19588), .ZN(
        P2_U3073) );
  AOI22_X1 U22568 ( .A1(n19628), .A2(n19988), .B1(n19601), .B2(n19986), .ZN(
        n19591) );
  AOI22_X1 U22569 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19603), .B1(
        n19987), .B2(n19602), .ZN(n19590) );
  OAI211_X1 U22570 ( .C1(n19991), .C2(n19606), .A(n19591), .B(n19590), .ZN(
        P2_U3074) );
  AOI22_X1 U22571 ( .A1(n19944), .A2(n19592), .B1(n19601), .B2(n19992), .ZN(
        n19594) );
  AOI22_X1 U22572 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19603), .B1(
        n19993), .B2(n19602), .ZN(n19593) );
  OAI211_X1 U22573 ( .C1(n19782), .C2(n19638), .A(n19594), .B(n19593), .ZN(
        P2_U3075) );
  AOI22_X1 U22574 ( .A1(n19628), .A2(n20000), .B1(n19601), .B2(n19998), .ZN(
        n19596) );
  AOI22_X1 U22575 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19603), .B1(
        n19999), .B2(n19602), .ZN(n19595) );
  OAI211_X1 U22576 ( .C1(n20003), .C2(n19606), .A(n19596), .B(n19595), .ZN(
        P2_U3076) );
  AOI22_X1 U22577 ( .A1(n19628), .A2(n20006), .B1(n19601), .B2(n20004), .ZN(
        n19598) );
  AOI22_X1 U22578 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19603), .B1(
        n20005), .B2(n19602), .ZN(n19597) );
  OAI211_X1 U22579 ( .C1(n20009), .C2(n19606), .A(n19598), .B(n19597), .ZN(
        P2_U3077) );
  AOI22_X1 U22580 ( .A1(n19628), .A2(n20012), .B1(n19601), .B2(n20010), .ZN(
        n19600) );
  AOI22_X1 U22581 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19603), .B1(
        n20011), .B2(n19602), .ZN(n19599) );
  OAI211_X1 U22582 ( .C1(n20015), .C2(n19606), .A(n19600), .B(n19599), .ZN(
        P2_U3078) );
  INV_X1 U22583 ( .A(n19827), .ZN(n20020) );
  AOI22_X1 U22584 ( .A1(n19628), .A2(n20020), .B1(n19601), .B2(n20016), .ZN(
        n19605) );
  AOI22_X1 U22585 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19603), .B1(
        n20018), .B2(n19602), .ZN(n19604) );
  OAI211_X1 U22586 ( .C1(n20026), .C2(n19606), .A(n19605), .B(n19604), .ZN(
        P2_U3079) );
  NOR2_X1 U22587 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20147), .ZN(
        n19699) );
  NAND2_X1 U22588 ( .A1(n19699), .A2(n16450), .ZN(n19645) );
  NOR2_X1 U22589 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19645), .ZN(
        n19633) );
  NOR3_X1 U22590 ( .A1(n19607), .A2(n19633), .A3(n20158), .ZN(n19613) );
  INV_X1 U22591 ( .A(n19671), .ZN(n19608) );
  NAND2_X1 U22592 ( .A1(n19609), .A2(n19608), .ZN(n19867) );
  NOR2_X1 U22593 ( .A1(n19867), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19617) );
  AOI21_X1 U22594 ( .B1(n20136), .B2(n19617), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19610) );
  AOI22_X1 U22595 ( .A1(n19634), .A2(n19968), .B1(n19967), .B2(n19633), .ZN(
        n19619) );
  AOI21_X1 U22596 ( .B1(n19638), .B2(n19661), .A(n19612), .ZN(n19616) );
  INV_X1 U22597 ( .A(n19633), .ZN(n19614) );
  AOI211_X1 U22598 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19614), .A(n19673), 
        .B(n19613), .ZN(n19615) );
  AOI22_X1 U22599 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19635), .B1(
        n19663), .B2(n19976), .ZN(n19618) );
  OAI211_X1 U22600 ( .C1(n19979), .C2(n19638), .A(n19619), .B(n19618), .ZN(
        P2_U3080) );
  AOI22_X1 U22601 ( .A1(n19634), .A2(n19981), .B1(n19980), .B2(n19633), .ZN(
        n19621) );
  AOI22_X1 U22602 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19635), .B1(
        n19663), .B2(n19982), .ZN(n19620) );
  OAI211_X1 U22603 ( .C1(n19985), .C2(n19638), .A(n19621), .B(n19620), .ZN(
        P2_U3081) );
  AOI22_X1 U22604 ( .A1(n19634), .A2(n19987), .B1(n19986), .B2(n19633), .ZN(
        n19623) );
  AOI22_X1 U22605 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19635), .B1(
        n19663), .B2(n19988), .ZN(n19622) );
  OAI211_X1 U22606 ( .C1(n19991), .C2(n19638), .A(n19623), .B(n19622), .ZN(
        P2_U3082) );
  AOI22_X1 U22607 ( .A1(n19634), .A2(n19993), .B1(n19992), .B2(n19633), .ZN(
        n19625) );
  AOI22_X1 U22608 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19635), .B1(
        n19628), .B2(n19944), .ZN(n19624) );
  OAI211_X1 U22609 ( .C1(n19782), .C2(n19661), .A(n19625), .B(n19624), .ZN(
        P2_U3083) );
  AOI22_X1 U22610 ( .A1(n19634), .A2(n19999), .B1(n19998), .B2(n19633), .ZN(
        n19627) );
  AOI22_X1 U22611 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19635), .B1(
        n19628), .B2(n19947), .ZN(n19626) );
  OAI211_X1 U22612 ( .C1(n19814), .C2(n19661), .A(n19627), .B(n19626), .ZN(
        P2_U3084) );
  AOI22_X1 U22613 ( .A1(n19634), .A2(n20005), .B1(n20004), .B2(n19633), .ZN(
        n19630) );
  AOI22_X1 U22614 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19635), .B1(
        n19628), .B2(n19950), .ZN(n19629) );
  OAI211_X1 U22615 ( .C1(n19817), .C2(n19661), .A(n19630), .B(n19629), .ZN(
        P2_U3085) );
  AOI22_X1 U22616 ( .A1(n19634), .A2(n20011), .B1(n20010), .B2(n19633), .ZN(
        n19632) );
  AOI22_X1 U22617 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19635), .B1(
        n19663), .B2(n20012), .ZN(n19631) );
  OAI211_X1 U22618 ( .C1(n20015), .C2(n19638), .A(n19632), .B(n19631), .ZN(
        P2_U3086) );
  AOI22_X1 U22619 ( .A1(n19634), .A2(n20018), .B1(n20016), .B2(n19633), .ZN(
        n19637) );
  AOI22_X1 U22620 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19635), .B1(
        n19663), .B2(n20020), .ZN(n19636) );
  OAI211_X1 U22621 ( .C1(n20026), .C2(n19638), .A(n19637), .B(n19636), .ZN(
        P2_U3087) );
  INV_X1 U22622 ( .A(n19699), .ZN(n19670) );
  NOR2_X1 U22623 ( .A1(n19763), .A2(n19670), .ZN(n19662) );
  AOI22_X1 U22624 ( .A1(n19929), .A2(n19663), .B1(n19662), .B2(n19967), .ZN(
        n19648) );
  OAI21_X1 U22625 ( .B1(n19639), .B2(n19898), .A(n20126), .ZN(n19646) );
  INV_X1 U22626 ( .A(n19645), .ZN(n19643) );
  INV_X1 U22627 ( .A(n10705), .ZN(n19641) );
  INV_X1 U22628 ( .A(n19662), .ZN(n19640) );
  OAI211_X1 U22629 ( .C1(n19641), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19640), 
        .B(n19765), .ZN(n19642) );
  OAI211_X1 U22630 ( .C1(n19646), .C2(n19643), .A(n19974), .B(n19642), .ZN(
        n19665) );
  OAI21_X1 U22631 ( .B1(n10705), .B2(n19662), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19644) );
  OAI21_X1 U22632 ( .B1(n19646), .B2(n19645), .A(n19644), .ZN(n19664) );
  AOI22_X1 U22633 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19665), .B1(
        n19968), .B2(n19664), .ZN(n19647) );
  OAI211_X1 U22634 ( .C1(n19839), .C2(n19697), .A(n19648), .B(n19647), .ZN(
        P2_U3088) );
  AOI22_X1 U22635 ( .A1(n19937), .A2(n19663), .B1(n19662), .B2(n19980), .ZN(
        n19650) );
  AOI22_X1 U22636 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19665), .B1(
        n19981), .B2(n19664), .ZN(n19649) );
  OAI211_X1 U22637 ( .C1(n19843), .C2(n19697), .A(n19650), .B(n19649), .ZN(
        P2_U3089) );
  AOI22_X1 U22638 ( .A1(n19685), .A2(n19988), .B1(n19986), .B2(n19662), .ZN(
        n19652) );
  AOI22_X1 U22639 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19665), .B1(
        n19987), .B2(n19664), .ZN(n19651) );
  OAI211_X1 U22640 ( .C1(n19991), .C2(n19661), .A(n19652), .B(n19651), .ZN(
        P2_U3090) );
  AOI22_X1 U22641 ( .A1(n19944), .A2(n19663), .B1(n19662), .B2(n19992), .ZN(
        n19654) );
  AOI22_X1 U22642 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19665), .B1(
        n19993), .B2(n19664), .ZN(n19653) );
  OAI211_X1 U22643 ( .C1(n19782), .C2(n19697), .A(n19654), .B(n19653), .ZN(
        P2_U3091) );
  AOI22_X1 U22644 ( .A1(n19947), .A2(n19663), .B1(n19662), .B2(n19998), .ZN(
        n19656) );
  AOI22_X1 U22645 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19665), .B1(
        n19999), .B2(n19664), .ZN(n19655) );
  OAI211_X1 U22646 ( .C1(n19814), .C2(n19697), .A(n19656), .B(n19655), .ZN(
        P2_U3092) );
  AOI22_X1 U22647 ( .A1(n19685), .A2(n20006), .B1(n19662), .B2(n20004), .ZN(
        n19658) );
  AOI22_X1 U22648 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19665), .B1(
        n20005), .B2(n19664), .ZN(n19657) );
  OAI211_X1 U22649 ( .C1(n20009), .C2(n19661), .A(n19658), .B(n19657), .ZN(
        P2_U3093) );
  AOI22_X1 U22650 ( .A1(n19685), .A2(n20012), .B1(n19662), .B2(n20010), .ZN(
        n19660) );
  AOI22_X1 U22651 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19665), .B1(
        n20011), .B2(n19664), .ZN(n19659) );
  OAI211_X1 U22652 ( .C1(n20015), .C2(n19661), .A(n19660), .B(n19659), .ZN(
        P2_U3094) );
  AOI22_X1 U22653 ( .A1(n19958), .A2(n19663), .B1(n19662), .B2(n20016), .ZN(
        n19667) );
  AOI22_X1 U22654 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19665), .B1(
        n20018), .B2(n19664), .ZN(n19666) );
  OAI211_X1 U22655 ( .C1(n19827), .C2(n19697), .A(n19667), .B(n19666), .ZN(
        P2_U3095) );
  NOR2_X2 U22656 ( .A1(n19920), .A2(n19668), .ZN(n19723) );
  NOR2_X1 U22657 ( .A1(n19795), .A2(n19670), .ZN(n19692) );
  OAI21_X1 U22658 ( .B1(n10707), .B2(n19692), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19669) );
  OAI21_X1 U22659 ( .B1(n19670), .B2(n19797), .A(n19669), .ZN(n19693) );
  AOI22_X1 U22660 ( .A1(n19693), .A2(n19968), .B1(n19967), .B2(n19692), .ZN(
        n19678) );
  OAI21_X1 U22661 ( .B1(n19685), .B2(n19723), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19675) );
  NAND2_X1 U22662 ( .A1(n19671), .A2(n19699), .ZN(n19674) );
  AOI211_X1 U22663 ( .C1(n19675), .C2(n19674), .A(n19673), .B(n19672), .ZN(
        n19676) );
  AOI22_X1 U22664 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19694), .B1(
        n19685), .B2(n19929), .ZN(n19677) );
  OAI211_X1 U22665 ( .C1(n19839), .C2(n19732), .A(n19678), .B(n19677), .ZN(
        P2_U3096) );
  AOI22_X1 U22666 ( .A1(n19693), .A2(n19981), .B1(n19980), .B2(n19692), .ZN(
        n19680) );
  AOI22_X1 U22667 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19694), .B1(
        n19685), .B2(n19937), .ZN(n19679) );
  OAI211_X1 U22668 ( .C1(n19843), .C2(n19732), .A(n19680), .B(n19679), .ZN(
        P2_U3097) );
  AOI22_X1 U22669 ( .A1(n19693), .A2(n19987), .B1(n19986), .B2(n19692), .ZN(
        n19682) );
  AOI22_X1 U22670 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19694), .B1(
        n19723), .B2(n19988), .ZN(n19681) );
  OAI211_X1 U22671 ( .C1(n19991), .C2(n19697), .A(n19682), .B(n19681), .ZN(
        P2_U3098) );
  AOI22_X1 U22672 ( .A1(n19693), .A2(n19993), .B1(n19992), .B2(n19692), .ZN(
        n19684) );
  AOI22_X1 U22673 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19694), .B1(
        n19723), .B2(n19994), .ZN(n19683) );
  OAI211_X1 U22674 ( .C1(n19997), .C2(n19697), .A(n19684), .B(n19683), .ZN(
        P2_U3099) );
  AOI22_X1 U22675 ( .A1(n19693), .A2(n19999), .B1(n19998), .B2(n19692), .ZN(
        n19687) );
  AOI22_X1 U22676 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19694), .B1(
        n19685), .B2(n19947), .ZN(n19686) );
  OAI211_X1 U22677 ( .C1(n19814), .C2(n19732), .A(n19687), .B(n19686), .ZN(
        P2_U3100) );
  AOI22_X1 U22678 ( .A1(n19693), .A2(n20005), .B1(n20004), .B2(n19692), .ZN(
        n19689) );
  AOI22_X1 U22679 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19694), .B1(
        n19723), .B2(n20006), .ZN(n19688) );
  OAI211_X1 U22680 ( .C1(n20009), .C2(n19697), .A(n19689), .B(n19688), .ZN(
        P2_U3101) );
  AOI22_X1 U22681 ( .A1(n19693), .A2(n20011), .B1(n20010), .B2(n19692), .ZN(
        n19691) );
  AOI22_X1 U22682 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19694), .B1(
        n19723), .B2(n20012), .ZN(n19690) );
  OAI211_X1 U22683 ( .C1(n20015), .C2(n19697), .A(n19691), .B(n19690), .ZN(
        P2_U3102) );
  AOI22_X1 U22684 ( .A1(n19693), .A2(n20018), .B1(n20016), .B2(n19692), .ZN(
        n19696) );
  AOI22_X1 U22685 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19694), .B1(
        n19723), .B2(n20020), .ZN(n19695) );
  OAI211_X1 U22686 ( .C1(n20026), .C2(n19697), .A(n19696), .B(n19695), .ZN(
        P2_U3103) );
  INV_X1 U22687 ( .A(n19920), .ZN(n19969) );
  AND2_X1 U22688 ( .A1(n19698), .A2(n19969), .ZN(n20125) );
  NOR2_X1 U22689 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19924), .ZN(
        n19705) );
  OAI21_X1 U22690 ( .B1(n20125), .B2(n19705), .A(n19974), .ZN(n19704) );
  INV_X1 U22691 ( .A(n19829), .ZN(n19700) );
  NAND2_X1 U22692 ( .A1(n19700), .A2(n19699), .ZN(n19735) );
  INV_X1 U22693 ( .A(n19735), .ZN(n19738) );
  NAND2_X1 U22694 ( .A1(n19735), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19701) );
  OAI21_X1 U22695 ( .B1(n19738), .B2(n20136), .A(n19708), .ZN(n19703) );
  INV_X1 U22696 ( .A(n19729), .ZN(n19727) );
  INV_X1 U22697 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n19712) );
  INV_X1 U22698 ( .A(n19705), .ZN(n19706) );
  OAI21_X1 U22699 ( .B1(n19706), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20158), 
        .ZN(n19707) );
  AND2_X1 U22700 ( .A1(n19708), .A2(n19707), .ZN(n19728) );
  AOI22_X1 U22701 ( .A1(n19728), .A2(n19968), .B1(n19738), .B2(n19967), .ZN(
        n19711) );
  AOI22_X1 U22702 ( .A1(n19758), .A2(n19976), .B1(n19723), .B2(n19929), .ZN(
        n19710) );
  OAI211_X1 U22703 ( .C1(n19727), .C2(n19712), .A(n19711), .B(n19710), .ZN(
        P2_U3104) );
  AOI22_X1 U22704 ( .A1(n19728), .A2(n19981), .B1(n19738), .B2(n19980), .ZN(
        n19714) );
  AOI22_X1 U22705 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19729), .B1(
        n19723), .B2(n19937), .ZN(n19713) );
  OAI211_X1 U22706 ( .C1(n19843), .C2(n19750), .A(n19714), .B(n19713), .ZN(
        P2_U3105) );
  INV_X1 U22707 ( .A(n19988), .ZN(n19779) );
  AOI22_X1 U22708 ( .A1(n19728), .A2(n19987), .B1(n19738), .B2(n19986), .ZN(
        n19716) );
  AOI22_X1 U22709 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19729), .B1(
        n19723), .B2(n19941), .ZN(n19715) );
  OAI211_X1 U22710 ( .C1(n19779), .C2(n19750), .A(n19716), .B(n19715), .ZN(
        P2_U3106) );
  AOI22_X1 U22711 ( .A1(n19728), .A2(n19993), .B1(n19738), .B2(n19992), .ZN(
        n19718) );
  AOI22_X1 U22712 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19729), .B1(
        n19723), .B2(n19944), .ZN(n19717) );
  OAI211_X1 U22713 ( .C1(n19782), .C2(n19750), .A(n19718), .B(n19717), .ZN(
        P2_U3107) );
  AOI22_X1 U22714 ( .A1(n19728), .A2(n19999), .B1(n19738), .B2(n19998), .ZN(
        n19720) );
  AOI22_X1 U22715 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19729), .B1(
        n19723), .B2(n19947), .ZN(n19719) );
  OAI211_X1 U22716 ( .C1(n19814), .C2(n19750), .A(n19720), .B(n19719), .ZN(
        P2_U3108) );
  AOI22_X1 U22717 ( .A1(n19728), .A2(n20005), .B1(n19738), .B2(n20004), .ZN(
        n19722) );
  AOI22_X1 U22718 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19729), .B1(
        n19758), .B2(n20006), .ZN(n19721) );
  OAI211_X1 U22719 ( .C1(n20009), .C2(n19732), .A(n19722), .B(n19721), .ZN(
        P2_U3109) );
  INV_X1 U22720 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n19726) );
  AOI22_X1 U22721 ( .A1(n19728), .A2(n20011), .B1(n19738), .B2(n20010), .ZN(
        n19725) );
  AOI22_X1 U22722 ( .A1(n19758), .A2(n20012), .B1(n19723), .B2(n19954), .ZN(
        n19724) );
  OAI211_X1 U22723 ( .C1(n19727), .C2(n19726), .A(n19725), .B(n19724), .ZN(
        P2_U3110) );
  AOI22_X1 U22724 ( .A1(n19728), .A2(n20018), .B1(n19738), .B2(n20016), .ZN(
        n19731) );
  AOI22_X1 U22725 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19729), .B1(
        n19758), .B2(n20020), .ZN(n19730) );
  OAI211_X1 U22726 ( .C1(n20026), .C2(n19732), .A(n19731), .B(n19730), .ZN(
        P2_U3111) );
  NAND2_X1 U22727 ( .A1(n20147), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19828) );
  NOR2_X1 U22728 ( .A1(n19828), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19769) );
  INV_X1 U22729 ( .A(n19769), .ZN(n19771) );
  NOR2_X1 U22730 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19771), .ZN(
        n19757) );
  AOI22_X1 U22731 ( .A1(n19976), .A2(n19790), .B1(n19967), .B2(n19757), .ZN(
        n19743) );
  NAND2_X1 U22732 ( .A1(n19750), .A2(n20126), .ZN(n19733) );
  OAI21_X1 U22733 ( .B1(n19733), .B2(n19790), .A(n19922), .ZN(n19737) );
  AOI21_X1 U22734 ( .B1(n19739), .B2(n20136), .A(n20126), .ZN(n19734) );
  AOI21_X1 U22735 ( .B1(n19737), .B2(n19735), .A(n19734), .ZN(n19736) );
  OAI21_X1 U22736 ( .B1(n19757), .B2(n19736), .A(n19974), .ZN(n19760) );
  OAI21_X1 U22737 ( .B1(n19738), .B2(n19757), .A(n19737), .ZN(n19741) );
  OAI21_X1 U22738 ( .B1(n19739), .B2(n19757), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19740) );
  NAND2_X1 U22739 ( .A1(n19741), .A2(n19740), .ZN(n19759) );
  AOI22_X1 U22740 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19760), .B1(
        n19968), .B2(n19759), .ZN(n19742) );
  OAI211_X1 U22741 ( .C1(n19979), .C2(n19750), .A(n19743), .B(n19742), .ZN(
        P2_U3112) );
  AOI22_X1 U22742 ( .A1(n19982), .A2(n19790), .B1(n19980), .B2(n19757), .ZN(
        n19745) );
  AOI22_X1 U22743 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19760), .B1(
        n19759), .B2(n19981), .ZN(n19744) );
  OAI211_X1 U22744 ( .C1(n19985), .C2(n19750), .A(n19745), .B(n19744), .ZN(
        P2_U3113) );
  AOI22_X1 U22745 ( .A1(n19988), .A2(n19790), .B1(n19986), .B2(n19757), .ZN(
        n19747) );
  AOI22_X1 U22746 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19760), .B1(
        n19759), .B2(n19987), .ZN(n19746) );
  OAI211_X1 U22747 ( .C1(n19991), .C2(n19750), .A(n19747), .B(n19746), .ZN(
        P2_U3114) );
  AOI22_X1 U22748 ( .A1(n19790), .A2(n19994), .B1(n19992), .B2(n19757), .ZN(
        n19749) );
  AOI22_X1 U22749 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19760), .B1(
        n19759), .B2(n19993), .ZN(n19748) );
  OAI211_X1 U22750 ( .C1(n19997), .C2(n19750), .A(n19749), .B(n19748), .ZN(
        P2_U3115) );
  AOI22_X1 U22751 ( .A1(n19758), .A2(n19947), .B1(n19998), .B2(n19757), .ZN(
        n19752) );
  AOI22_X1 U22752 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19760), .B1(
        n19759), .B2(n19999), .ZN(n19751) );
  OAI211_X1 U22753 ( .C1(n19814), .C2(n19789), .A(n19752), .B(n19751), .ZN(
        P2_U3116) );
  AOI22_X1 U22754 ( .A1(n19758), .A2(n19950), .B1(n20004), .B2(n19757), .ZN(
        n19754) );
  AOI22_X1 U22755 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19760), .B1(
        n19759), .B2(n20005), .ZN(n19753) );
  OAI211_X1 U22756 ( .C1(n19817), .C2(n19789), .A(n19754), .B(n19753), .ZN(
        P2_U3117) );
  AOI22_X1 U22757 ( .A1(n19758), .A2(n19954), .B1(n20010), .B2(n19757), .ZN(
        n19756) );
  AOI22_X1 U22758 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19760), .B1(
        n19759), .B2(n20011), .ZN(n19755) );
  OAI211_X1 U22759 ( .C1(n19820), .C2(n19789), .A(n19756), .B(n19755), .ZN(
        P2_U3118) );
  AOI22_X1 U22760 ( .A1(n19758), .A2(n19958), .B1(n20016), .B2(n19757), .ZN(
        n19762) );
  AOI22_X1 U22761 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19760), .B1(
        n19759), .B2(n20018), .ZN(n19761) );
  OAI211_X1 U22762 ( .C1(n19827), .C2(n19789), .A(n19762), .B(n19761), .ZN(
        P2_U3119) );
  NOR2_X1 U22763 ( .A1(n19763), .A2(n19828), .ZN(n19799) );
  AOI22_X1 U22764 ( .A1(n19929), .A2(n19790), .B1(n19967), .B2(n19799), .ZN(
        n19774) );
  NAND2_X1 U22765 ( .A1(n20132), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19831) );
  OAI21_X1 U22766 ( .B1(n19831), .B2(n19764), .A(n20126), .ZN(n19772) );
  INV_X1 U22767 ( .A(n10818), .ZN(n19767) );
  INV_X1 U22768 ( .A(n19799), .ZN(n19766) );
  OAI211_X1 U22769 ( .C1(n19767), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19766), 
        .B(n19765), .ZN(n19768) );
  OAI211_X1 U22770 ( .C1(n19772), .C2(n19769), .A(n19974), .B(n19768), .ZN(
        n19792) );
  OAI21_X1 U22771 ( .B1(n10818), .B2(n19799), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19770) );
  OAI21_X1 U22772 ( .B1(n19772), .B2(n19771), .A(n19770), .ZN(n19791) );
  AOI22_X1 U22773 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19792), .B1(
        n19968), .B2(n19791), .ZN(n19773) );
  OAI211_X1 U22774 ( .C1(n19839), .C2(n19811), .A(n19774), .B(n19773), .ZN(
        P2_U3120) );
  AOI22_X1 U22775 ( .A1(n19982), .A2(n19823), .B1(n19980), .B2(n19799), .ZN(
        n19776) );
  AOI22_X1 U22776 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19792), .B1(
        n19981), .B2(n19791), .ZN(n19775) );
  OAI211_X1 U22777 ( .C1(n19985), .C2(n19789), .A(n19776), .B(n19775), .ZN(
        P2_U3121) );
  AOI22_X1 U22778 ( .A1(n19941), .A2(n19790), .B1(n19986), .B2(n19799), .ZN(
        n19778) );
  AOI22_X1 U22779 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19792), .B1(
        n19987), .B2(n19791), .ZN(n19777) );
  OAI211_X1 U22780 ( .C1(n19779), .C2(n19811), .A(n19778), .B(n19777), .ZN(
        P2_U3122) );
  AOI22_X1 U22781 ( .A1(n19944), .A2(n19790), .B1(n19992), .B2(n19799), .ZN(
        n19781) );
  AOI22_X1 U22782 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19792), .B1(
        n19993), .B2(n19791), .ZN(n19780) );
  OAI211_X1 U22783 ( .C1(n19782), .C2(n19811), .A(n19781), .B(n19780), .ZN(
        P2_U3123) );
  AOI22_X1 U22784 ( .A1(n20000), .A2(n19823), .B1(n19998), .B2(n19799), .ZN(
        n19784) );
  AOI22_X1 U22785 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19792), .B1(
        n19999), .B2(n19791), .ZN(n19783) );
  OAI211_X1 U22786 ( .C1(n20003), .C2(n19789), .A(n19784), .B(n19783), .ZN(
        P2_U3124) );
  AOI22_X1 U22787 ( .A1(n20006), .A2(n19823), .B1(n20004), .B2(n19799), .ZN(
        n19786) );
  AOI22_X1 U22788 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19792), .B1(
        n20005), .B2(n19791), .ZN(n19785) );
  OAI211_X1 U22789 ( .C1(n20009), .C2(n19789), .A(n19786), .B(n19785), .ZN(
        P2_U3125) );
  AOI22_X1 U22790 ( .A1(n20012), .A2(n19823), .B1(n20010), .B2(n19799), .ZN(
        n19788) );
  AOI22_X1 U22791 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19792), .B1(
        n20011), .B2(n19791), .ZN(n19787) );
  OAI211_X1 U22792 ( .C1(n20015), .C2(n19789), .A(n19788), .B(n19787), .ZN(
        P2_U3126) );
  AOI22_X1 U22793 ( .A1(n19958), .A2(n19790), .B1(n20016), .B2(n19799), .ZN(
        n19794) );
  AOI22_X1 U22794 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19792), .B1(
        n20018), .B2(n19791), .ZN(n19793) );
  OAI211_X1 U22795 ( .C1(n19827), .C2(n19811), .A(n19794), .B(n19793), .ZN(
        P2_U3127) );
  NOR2_X1 U22796 ( .A1(n19795), .A2(n19828), .ZN(n19821) );
  OAI21_X1 U22797 ( .B1(n19798), .B2(n19821), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19796) );
  OAI21_X1 U22798 ( .B1(n19828), .B2(n19797), .A(n19796), .ZN(n19822) );
  AOI22_X1 U22799 ( .A1(n19822), .A2(n19968), .B1(n19967), .B2(n19821), .ZN(
        n19804) );
  INV_X1 U22800 ( .A(n19798), .ZN(n19801) );
  AOI221_X1 U22801 ( .B1(n19823), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19840), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19799), .ZN(n19800) );
  AOI211_X1 U22802 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19801), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19800), .ZN(n19802) );
  OAI21_X1 U22803 ( .B1(n19802), .B2(n19821), .A(n19974), .ZN(n19824) );
  AOI22_X1 U22804 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19824), .B1(
        n19840), .B2(n19976), .ZN(n19803) );
  OAI211_X1 U22805 ( .C1(n19979), .C2(n19811), .A(n19804), .B(n19803), .ZN(
        P2_U3128) );
  AOI22_X1 U22806 ( .A1(n19822), .A2(n19981), .B1(n19980), .B2(n19821), .ZN(
        n19806) );
  AOI22_X1 U22807 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19824), .B1(
        n19840), .B2(n19982), .ZN(n19805) );
  OAI211_X1 U22808 ( .C1(n19985), .C2(n19811), .A(n19806), .B(n19805), .ZN(
        P2_U3129) );
  AOI22_X1 U22809 ( .A1(n19822), .A2(n19987), .B1(n19986), .B2(n19821), .ZN(
        n19808) );
  AOI22_X1 U22810 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19824), .B1(
        n19840), .B2(n19988), .ZN(n19807) );
  OAI211_X1 U22811 ( .C1(n19991), .C2(n19811), .A(n19808), .B(n19807), .ZN(
        P2_U3130) );
  AOI22_X1 U22812 ( .A1(n19822), .A2(n19993), .B1(n19992), .B2(n19821), .ZN(
        n19810) );
  AOI22_X1 U22813 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19824), .B1(
        n19840), .B2(n19994), .ZN(n19809) );
  OAI211_X1 U22814 ( .C1(n19997), .C2(n19811), .A(n19810), .B(n19809), .ZN(
        P2_U3131) );
  AOI22_X1 U22815 ( .A1(n19822), .A2(n19999), .B1(n19998), .B2(n19821), .ZN(
        n19813) );
  AOI22_X1 U22816 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19824), .B1(
        n19823), .B2(n19947), .ZN(n19812) );
  OAI211_X1 U22817 ( .C1(n19814), .C2(n19859), .A(n19813), .B(n19812), .ZN(
        P2_U3132) );
  AOI22_X1 U22818 ( .A1(n19822), .A2(n20005), .B1(n20004), .B2(n19821), .ZN(
        n19816) );
  AOI22_X1 U22819 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19824), .B1(
        n19823), .B2(n19950), .ZN(n19815) );
  OAI211_X1 U22820 ( .C1(n19817), .C2(n19859), .A(n19816), .B(n19815), .ZN(
        P2_U3133) );
  AOI22_X1 U22821 ( .A1(n19822), .A2(n20011), .B1(n20010), .B2(n19821), .ZN(
        n19819) );
  AOI22_X1 U22822 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19824), .B1(
        n19823), .B2(n19954), .ZN(n19818) );
  OAI211_X1 U22823 ( .C1(n19820), .C2(n19859), .A(n19819), .B(n19818), .ZN(
        P2_U3134) );
  AOI22_X1 U22824 ( .A1(n19822), .A2(n20018), .B1(n20016), .B2(n19821), .ZN(
        n19826) );
  AOI22_X1 U22825 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19824), .B1(
        n19823), .B2(n19958), .ZN(n19825) );
  OAI211_X1 U22826 ( .C1(n19827), .C2(n19859), .A(n19826), .B(n19825), .ZN(
        P2_U3135) );
  OR2_X1 U22827 ( .A1(n16450), .A2(n19828), .ZN(n19834) );
  OR2_X1 U22828 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19834), .ZN(n19830) );
  NOR2_X1 U22829 ( .A1(n19829), .A2(n19828), .ZN(n19854) );
  NOR3_X1 U22830 ( .A1(n10817), .A2(n19854), .A3(n20158), .ZN(n19833) );
  AOI21_X1 U22831 ( .B1(n20158), .B2(n19830), .A(n19833), .ZN(n19855) );
  AOI22_X1 U22832 ( .A1(n19855), .A2(n19968), .B1(n19967), .B2(n19854), .ZN(
        n19838) );
  INV_X1 U22833 ( .A(n19831), .ZN(n19970) );
  INV_X1 U22834 ( .A(n20127), .ZN(n19832) );
  NAND2_X1 U22835 ( .A1(n19970), .A2(n19832), .ZN(n19835) );
  AOI21_X1 U22836 ( .B1(n19835), .B2(n19834), .A(n19833), .ZN(n19836) );
  OAI211_X1 U22837 ( .C1(n19854), .C2(n20136), .A(n19836), .B(n19974), .ZN(
        n19856) );
  AOI22_X1 U22838 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19856), .B1(
        n19840), .B2(n19929), .ZN(n19837) );
  OAI211_X1 U22839 ( .C1(n19839), .C2(n19889), .A(n19838), .B(n19837), .ZN(
        P2_U3136) );
  AOI22_X1 U22840 ( .A1(n19855), .A2(n19981), .B1(n19980), .B2(n19854), .ZN(
        n19842) );
  AOI22_X1 U22841 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19856), .B1(
        n19840), .B2(n19937), .ZN(n19841) );
  OAI211_X1 U22842 ( .C1(n19843), .C2(n19889), .A(n19842), .B(n19841), .ZN(
        P2_U3137) );
  AOI22_X1 U22843 ( .A1(n19855), .A2(n19987), .B1(n19986), .B2(n19854), .ZN(
        n19845) );
  AOI22_X1 U22844 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19856), .B1(
        n19865), .B2(n19988), .ZN(n19844) );
  OAI211_X1 U22845 ( .C1(n19991), .C2(n19859), .A(n19845), .B(n19844), .ZN(
        P2_U3138) );
  AOI22_X1 U22846 ( .A1(n19855), .A2(n19993), .B1(n19992), .B2(n19854), .ZN(
        n19847) );
  AOI22_X1 U22847 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19856), .B1(
        n19865), .B2(n19994), .ZN(n19846) );
  OAI211_X1 U22848 ( .C1(n19997), .C2(n19859), .A(n19847), .B(n19846), .ZN(
        P2_U3139) );
  AOI22_X1 U22849 ( .A1(n19855), .A2(n19999), .B1(n19998), .B2(n19854), .ZN(
        n19849) );
  AOI22_X1 U22850 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19856), .B1(
        n19865), .B2(n20000), .ZN(n19848) );
  OAI211_X1 U22851 ( .C1(n20003), .C2(n19859), .A(n19849), .B(n19848), .ZN(
        P2_U3140) );
  AOI22_X1 U22852 ( .A1(n19855), .A2(n20005), .B1(n20004), .B2(n19854), .ZN(
        n19851) );
  AOI22_X1 U22853 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19856), .B1(
        n19865), .B2(n20006), .ZN(n19850) );
  OAI211_X1 U22854 ( .C1(n20009), .C2(n19859), .A(n19851), .B(n19850), .ZN(
        P2_U3141) );
  AOI22_X1 U22855 ( .A1(n19855), .A2(n20011), .B1(n20010), .B2(n19854), .ZN(
        n19853) );
  AOI22_X1 U22856 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19856), .B1(
        n19865), .B2(n20012), .ZN(n19852) );
  OAI211_X1 U22857 ( .C1(n20015), .C2(n19859), .A(n19853), .B(n19852), .ZN(
        P2_U3142) );
  AOI22_X1 U22858 ( .A1(n19855), .A2(n20018), .B1(n20016), .B2(n19854), .ZN(
        n19858) );
  AOI22_X1 U22859 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19856), .B1(
        n19865), .B2(n20020), .ZN(n19857) );
  OAI211_X1 U22860 ( .C1(n20026), .C2(n19859), .A(n19858), .B(n19857), .ZN(
        P2_U3143) );
  INV_X1 U22861 ( .A(n19860), .ZN(n19862) );
  NAND3_X1 U22862 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n16450), .ZN(n19895) );
  NOR2_X1 U22863 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19895), .ZN(
        n19884) );
  OAI21_X1 U22864 ( .B1(n19863), .B2(n19884), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19861) );
  OAI21_X1 U22865 ( .B1(n19862), .B2(n19867), .A(n19861), .ZN(n19885) );
  AOI22_X1 U22866 ( .A1(n19885), .A2(n19968), .B1(n19967), .B2(n19884), .ZN(
        n19871) );
  INV_X1 U22867 ( .A(n19863), .ZN(n19864) );
  AOI21_X1 U22868 ( .B1(n19864), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19869) );
  OAI21_X1 U22869 ( .B1(n19865), .B2(n19890), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19866) );
  OAI21_X1 U22870 ( .B1(n19867), .B2(n20140), .A(n19866), .ZN(n19868) );
  OAI211_X1 U22871 ( .C1(n19884), .C2(n19869), .A(n19868), .B(n19974), .ZN(
        n19886) );
  AOI22_X1 U22872 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19886), .B1(
        n19890), .B2(n19976), .ZN(n19870) );
  OAI211_X1 U22873 ( .C1(n19979), .C2(n19889), .A(n19871), .B(n19870), .ZN(
        P2_U3144) );
  AOI22_X1 U22874 ( .A1(n19885), .A2(n19981), .B1(n19980), .B2(n19884), .ZN(
        n19873) );
  AOI22_X1 U22875 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19886), .B1(
        n19890), .B2(n19982), .ZN(n19872) );
  OAI211_X1 U22876 ( .C1(n19985), .C2(n19889), .A(n19873), .B(n19872), .ZN(
        P2_U3145) );
  AOI22_X1 U22877 ( .A1(n19885), .A2(n19987), .B1(n19986), .B2(n19884), .ZN(
        n19875) );
  AOI22_X1 U22878 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19886), .B1(
        n19890), .B2(n19988), .ZN(n19874) );
  OAI211_X1 U22879 ( .C1(n19991), .C2(n19889), .A(n19875), .B(n19874), .ZN(
        P2_U3146) );
  AOI22_X1 U22880 ( .A1(n19885), .A2(n19993), .B1(n19992), .B2(n19884), .ZN(
        n19877) );
  AOI22_X1 U22881 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19886), .B1(
        n19890), .B2(n19994), .ZN(n19876) );
  OAI211_X1 U22882 ( .C1(n19997), .C2(n19889), .A(n19877), .B(n19876), .ZN(
        P2_U3147) );
  AOI22_X1 U22883 ( .A1(n19885), .A2(n19999), .B1(n19998), .B2(n19884), .ZN(
        n19879) );
  AOI22_X1 U22884 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19886), .B1(
        n19890), .B2(n20000), .ZN(n19878) );
  OAI211_X1 U22885 ( .C1(n20003), .C2(n19889), .A(n19879), .B(n19878), .ZN(
        P2_U3148) );
  AOI22_X1 U22886 ( .A1(n19885), .A2(n20005), .B1(n20004), .B2(n19884), .ZN(
        n19881) );
  AOI22_X1 U22887 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19886), .B1(
        n19890), .B2(n20006), .ZN(n19880) );
  OAI211_X1 U22888 ( .C1(n20009), .C2(n19889), .A(n19881), .B(n19880), .ZN(
        P2_U3149) );
  AOI22_X1 U22889 ( .A1(n19885), .A2(n20011), .B1(n20010), .B2(n19884), .ZN(
        n19883) );
  AOI22_X1 U22890 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19886), .B1(
        n19890), .B2(n20012), .ZN(n19882) );
  OAI211_X1 U22891 ( .C1(n20015), .C2(n19889), .A(n19883), .B(n19882), .ZN(
        P2_U3150) );
  AOI22_X1 U22892 ( .A1(n19885), .A2(n20018), .B1(n20016), .B2(n19884), .ZN(
        n19888) );
  AOI22_X1 U22893 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19886), .B1(
        n19890), .B2(n20020), .ZN(n19887) );
  OAI211_X1 U22894 ( .C1(n20026), .C2(n19889), .A(n19888), .B(n19887), .ZN(
        P2_U3151) );
  NOR2_X1 U22895 ( .A1(n20165), .A2(n19895), .ZN(n19925) );
  NOR3_X1 U22896 ( .A1(n10708), .A2(n19925), .A3(n20158), .ZN(n19894) );
  INV_X1 U22897 ( .A(n19895), .ZN(n19891) );
  AOI21_X1 U22898 ( .B1(n20136), .B2(n19891), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19892) );
  NOR2_X1 U22899 ( .A1(n19894), .A2(n19892), .ZN(n19914) );
  AOI22_X1 U22900 ( .A1(n19914), .A2(n19968), .B1(n19967), .B2(n19925), .ZN(
        n19901) );
  INV_X1 U22901 ( .A(n19898), .ZN(n19893) );
  NAND2_X1 U22902 ( .A1(n19970), .A2(n19893), .ZN(n19896) );
  AOI21_X1 U22903 ( .B1(n19896), .B2(n19895), .A(n19894), .ZN(n19897) );
  OAI211_X1 U22904 ( .C1(n19925), .C2(n20136), .A(n19897), .B(n19974), .ZN(
        n19915) );
  AOI22_X1 U22905 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19915), .B1(
        n19959), .B2(n19976), .ZN(n19900) );
  OAI211_X1 U22906 ( .C1(n19979), .C2(n19918), .A(n19901), .B(n19900), .ZN(
        P2_U3152) );
  AOI22_X1 U22907 ( .A1(n19914), .A2(n19981), .B1(n19980), .B2(n19925), .ZN(
        n19903) );
  AOI22_X1 U22908 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19915), .B1(
        n19959), .B2(n19982), .ZN(n19902) );
  OAI211_X1 U22909 ( .C1(n19985), .C2(n19918), .A(n19903), .B(n19902), .ZN(
        P2_U3153) );
  AOI22_X1 U22910 ( .A1(n19914), .A2(n19987), .B1(n19986), .B2(n19925), .ZN(
        n19905) );
  AOI22_X1 U22911 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19915), .B1(
        n19959), .B2(n19988), .ZN(n19904) );
  OAI211_X1 U22912 ( .C1(n19991), .C2(n19918), .A(n19905), .B(n19904), .ZN(
        P2_U3154) );
  AOI22_X1 U22913 ( .A1(n19914), .A2(n19993), .B1(n19992), .B2(n19925), .ZN(
        n19907) );
  AOI22_X1 U22914 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19915), .B1(
        n19959), .B2(n19994), .ZN(n19906) );
  OAI211_X1 U22915 ( .C1(n19997), .C2(n19918), .A(n19907), .B(n19906), .ZN(
        P2_U3155) );
  AOI22_X1 U22916 ( .A1(n19914), .A2(n19999), .B1(n19998), .B2(n19925), .ZN(
        n19909) );
  AOI22_X1 U22917 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19915), .B1(
        n19959), .B2(n20000), .ZN(n19908) );
  OAI211_X1 U22918 ( .C1(n20003), .C2(n19918), .A(n19909), .B(n19908), .ZN(
        P2_U3156) );
  AOI22_X1 U22919 ( .A1(n19914), .A2(n20005), .B1(n20004), .B2(n19925), .ZN(
        n19911) );
  AOI22_X1 U22920 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19915), .B1(
        n19959), .B2(n20006), .ZN(n19910) );
  OAI211_X1 U22921 ( .C1(n20009), .C2(n19918), .A(n19911), .B(n19910), .ZN(
        P2_U3157) );
  AOI22_X1 U22922 ( .A1(n19914), .A2(n20011), .B1(n20010), .B2(n19925), .ZN(
        n19913) );
  AOI22_X1 U22923 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19915), .B1(
        n19959), .B2(n20012), .ZN(n19912) );
  OAI211_X1 U22924 ( .C1(n20015), .C2(n19918), .A(n19913), .B(n19912), .ZN(
        P2_U3158) );
  AOI22_X1 U22925 ( .A1(n19914), .A2(n20018), .B1(n20016), .B2(n19925), .ZN(
        n19917) );
  AOI22_X1 U22926 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19915), .B1(
        n19959), .B2(n20020), .ZN(n19916) );
  OAI211_X1 U22927 ( .C1(n20026), .C2(n19918), .A(n19917), .B(n19916), .ZN(
        P2_U3159) );
  INV_X1 U22928 ( .A(n19959), .ZN(n19919) );
  NAND2_X1 U22929 ( .A1(n19919), .A2(n20126), .ZN(n19923) );
  OAI21_X1 U22930 ( .B1(n19923), .B2(n19964), .A(n19922), .ZN(n19930) );
  NOR3_X2 U22931 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20140), .A3(
        n19924), .ZN(n19957) );
  NOR2_X1 U22932 ( .A1(n19957), .A2(n19925), .ZN(n19932) );
  AOI21_X1 U22933 ( .B1(n19926), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19927) );
  OAI21_X1 U22934 ( .B1(n19927), .B2(n19957), .A(n19974), .ZN(n19928) );
  AOI22_X1 U22935 ( .A1(n19929), .A2(n19959), .B1(n19967), .B2(n19957), .ZN(
        n19935) );
  INV_X1 U22936 ( .A(n19930), .ZN(n19933) );
  OAI21_X1 U22937 ( .B1(n10823), .B2(n19957), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19931) );
  AOI22_X1 U22938 ( .A1(n19968), .A2(n19960), .B1(n19964), .B2(n19976), .ZN(
        n19934) );
  OAI211_X1 U22939 ( .C1(n19963), .C2(n19936), .A(n19935), .B(n19934), .ZN(
        P2_U3160) );
  INV_X1 U22940 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n19940) );
  AOI22_X1 U22941 ( .A1(n19982), .A2(n19964), .B1(n19980), .B2(n19957), .ZN(
        n19939) );
  AOI22_X1 U22942 ( .A1(n19981), .A2(n19960), .B1(n19959), .B2(n19937), .ZN(
        n19938) );
  OAI211_X1 U22943 ( .C1(n19963), .C2(n19940), .A(n19939), .B(n19938), .ZN(
        P2_U3161) );
  AOI22_X1 U22944 ( .A1(n19988), .A2(n19964), .B1(n19986), .B2(n19957), .ZN(
        n19943) );
  AOI22_X1 U22945 ( .A1(n19987), .A2(n19960), .B1(n19959), .B2(n19941), .ZN(
        n19942) );
  OAI211_X1 U22946 ( .C1(n19963), .C2(n10663), .A(n19943), .B(n19942), .ZN(
        P2_U3162) );
  AOI22_X1 U22947 ( .A1(n19944), .A2(n19959), .B1(n19992), .B2(n19957), .ZN(
        n19946) );
  AOI22_X1 U22948 ( .A1(n19993), .A2(n19960), .B1(n19964), .B2(n19994), .ZN(
        n19945) );
  OAI211_X1 U22949 ( .C1(n19963), .C2(n10771), .A(n19946), .B(n19945), .ZN(
        P2_U3163) );
  AOI22_X1 U22950 ( .A1(n20000), .A2(n19964), .B1(n19998), .B2(n19957), .ZN(
        n19949) );
  AOI22_X1 U22951 ( .A1(n19999), .A2(n19960), .B1(n19959), .B2(n19947), .ZN(
        n19948) );
  OAI211_X1 U22952 ( .C1(n19963), .C2(n10695), .A(n19949), .B(n19948), .ZN(
        P2_U3164) );
  INV_X1 U22953 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n19953) );
  AOI22_X1 U22954 ( .A1(n19964), .A2(n20006), .B1(n20004), .B2(n19957), .ZN(
        n19952) );
  AOI22_X1 U22955 ( .A1(n20005), .A2(n19960), .B1(n19959), .B2(n19950), .ZN(
        n19951) );
  OAI211_X1 U22956 ( .C1(n19963), .C2(n19953), .A(n19952), .B(n19951), .ZN(
        P2_U3165) );
  AOI22_X1 U22957 ( .A1(n19964), .A2(n20012), .B1(n20010), .B2(n19957), .ZN(
        n19956) );
  AOI22_X1 U22958 ( .A1(n20011), .A2(n19960), .B1(n19959), .B2(n19954), .ZN(
        n19955) );
  OAI211_X1 U22959 ( .C1(n19963), .C2(n10834), .A(n19956), .B(n19955), .ZN(
        P2_U3166) );
  AOI22_X1 U22960 ( .A1(n20020), .A2(n19964), .B1(n20016), .B2(n19957), .ZN(
        n19962) );
  AOI22_X1 U22961 ( .A1(n20018), .A2(n19960), .B1(n19959), .B2(n19958), .ZN(
        n19961) );
  OAI211_X1 U22962 ( .C1(n19963), .C2(n10746), .A(n19962), .B(n19961), .ZN(
        P2_U3167) );
  NAND2_X1 U22963 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19965), .ZN(
        n19972) );
  OR2_X1 U22964 ( .A1(n19972), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19966) );
  NOR3_X1 U22965 ( .A1(n10716), .A2(n20017), .A3(n20158), .ZN(n19971) );
  AOI21_X1 U22966 ( .B1(n20158), .B2(n19966), .A(n19971), .ZN(n20019) );
  AOI22_X1 U22967 ( .A1(n20019), .A2(n19968), .B1(n20017), .B2(n19967), .ZN(
        n19978) );
  NAND2_X1 U22968 ( .A1(n19970), .A2(n19969), .ZN(n19973) );
  AOI21_X1 U22969 ( .B1(n19973), .B2(n19972), .A(n19971), .ZN(n19975) );
  OAI211_X1 U22970 ( .C1(n20017), .C2(n20136), .A(n19975), .B(n19974), .ZN(
        n20022) );
  AOI22_X1 U22971 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20022), .B1(
        n20021), .B2(n19976), .ZN(n19977) );
  OAI211_X1 U22972 ( .C1(n19979), .C2(n20025), .A(n19978), .B(n19977), .ZN(
        P2_U3168) );
  AOI22_X1 U22973 ( .A1(n20019), .A2(n19981), .B1(n20017), .B2(n19980), .ZN(
        n19984) );
  AOI22_X1 U22974 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20022), .B1(
        n20021), .B2(n19982), .ZN(n19983) );
  OAI211_X1 U22975 ( .C1(n19985), .C2(n20025), .A(n19984), .B(n19983), .ZN(
        P2_U3169) );
  AOI22_X1 U22976 ( .A1(n20019), .A2(n19987), .B1(n20017), .B2(n19986), .ZN(
        n19990) );
  AOI22_X1 U22977 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20022), .B1(
        n20021), .B2(n19988), .ZN(n19989) );
  OAI211_X1 U22978 ( .C1(n19991), .C2(n20025), .A(n19990), .B(n19989), .ZN(
        P2_U3170) );
  AOI22_X1 U22979 ( .A1(n20019), .A2(n19993), .B1(n20017), .B2(n19992), .ZN(
        n19996) );
  AOI22_X1 U22980 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20022), .B1(
        n20021), .B2(n19994), .ZN(n19995) );
  OAI211_X1 U22981 ( .C1(n19997), .C2(n20025), .A(n19996), .B(n19995), .ZN(
        P2_U3171) );
  AOI22_X1 U22982 ( .A1(n20019), .A2(n19999), .B1(n20017), .B2(n19998), .ZN(
        n20002) );
  AOI22_X1 U22983 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20022), .B1(
        n20021), .B2(n20000), .ZN(n20001) );
  OAI211_X1 U22984 ( .C1(n20003), .C2(n20025), .A(n20002), .B(n20001), .ZN(
        P2_U3172) );
  AOI22_X1 U22985 ( .A1(n20019), .A2(n20005), .B1(n20017), .B2(n20004), .ZN(
        n20008) );
  AOI22_X1 U22986 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20022), .B1(
        n20021), .B2(n20006), .ZN(n20007) );
  OAI211_X1 U22987 ( .C1(n20009), .C2(n20025), .A(n20008), .B(n20007), .ZN(
        P2_U3173) );
  AOI22_X1 U22988 ( .A1(n20019), .A2(n20011), .B1(n20017), .B2(n20010), .ZN(
        n20014) );
  AOI22_X1 U22989 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20022), .B1(
        n20021), .B2(n20012), .ZN(n20013) );
  OAI211_X1 U22990 ( .C1(n20015), .C2(n20025), .A(n20014), .B(n20013), .ZN(
        P2_U3174) );
  AOI22_X1 U22991 ( .A1(n20019), .A2(n20018), .B1(n20017), .B2(n20016), .ZN(
        n20024) );
  AOI22_X1 U22992 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20022), .B1(
        n20021), .B2(n20020), .ZN(n20023) );
  OAI211_X1 U22993 ( .C1(n20026), .C2(n20025), .A(n20024), .B(n20023), .ZN(
        P2_U3175) );
  AOI21_X1 U22994 ( .B1(n20029), .B2(n20028), .A(n20027), .ZN(n20033) );
  OAI211_X1 U22995 ( .C1(n20034), .C2(n20030), .A(n20047), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n20031) );
  OAI211_X1 U22996 ( .C1(n20034), .C2(n20033), .A(n20032), .B(n20031), .ZN(
        P2_U3177) );
  AND2_X1 U22997 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20035), .ZN(
        P2_U3179) );
  AND2_X1 U22998 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20035), .ZN(
        P2_U3180) );
  AND2_X1 U22999 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20035), .ZN(
        P2_U3181) );
  AND2_X1 U23000 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20035), .ZN(
        P2_U3182) );
  AND2_X1 U23001 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20035), .ZN(
        P2_U3183) );
  AND2_X1 U23002 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20035), .ZN(
        P2_U3184) );
  AND2_X1 U23003 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20035), .ZN(
        P2_U3185) );
  AND2_X1 U23004 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20035), .ZN(
        P2_U3186) );
  AND2_X1 U23005 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20035), .ZN(
        P2_U3187) );
  AND2_X1 U23006 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20035), .ZN(
        P2_U3188) );
  AND2_X1 U23007 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20035), .ZN(
        P2_U3189) );
  AND2_X1 U23008 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20035), .ZN(
        P2_U3190) );
  AND2_X1 U23009 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20035), .ZN(
        P2_U3191) );
  AND2_X1 U23010 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20035), .ZN(
        P2_U3192) );
  AND2_X1 U23011 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20035), .ZN(
        P2_U3193) );
  AND2_X1 U23012 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20035), .ZN(
        P2_U3194) );
  AND2_X1 U23013 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20035), .ZN(
        P2_U3195) );
  AND2_X1 U23014 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20035), .ZN(
        P2_U3196) );
  AND2_X1 U23015 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20035), .ZN(
        P2_U3197) );
  AND2_X1 U23016 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20035), .ZN(
        P2_U3198) );
  AND2_X1 U23017 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20035), .ZN(
        P2_U3199) );
  AND2_X1 U23018 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20035), .ZN(
        P2_U3200) );
  AND2_X1 U23019 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20035), .ZN(P2_U3201) );
  AND2_X1 U23020 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20035), .ZN(P2_U3202) );
  AND2_X1 U23021 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20035), .ZN(P2_U3203) );
  AND2_X1 U23022 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20035), .ZN(P2_U3204) );
  AND2_X1 U23023 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20035), .ZN(P2_U3205) );
  AND2_X1 U23024 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20035), .ZN(P2_U3206) );
  AND2_X1 U23025 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20035), .ZN(P2_U3207) );
  AND2_X1 U23026 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20035), .ZN(P2_U3208) );
  NAND2_X1 U23027 ( .A1(n20047), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n20049) );
  NAND3_X1 U23028 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n20049), .ZN(n20038) );
  AOI211_X1 U23029 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n21002), .A(
        n20036), .B(n20178), .ZN(n20037) );
  NOR2_X1 U23030 ( .A1(n21132), .A2(n20042), .ZN(n20054) );
  AOI211_X1 U23031 ( .C1(n20055), .C2(n20038), .A(n20037), .B(n20054), .ZN(
        n20039) );
  INV_X1 U23032 ( .A(n20039), .ZN(P2_U3209) );
  INV_X1 U23033 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20040) );
  AOI21_X1 U23034 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21002), .A(n20055), 
        .ZN(n20046) );
  NOR2_X1 U23035 ( .A1(n20040), .A2(n20046), .ZN(n20043) );
  AOI21_X1 U23036 ( .B1(n20043), .B2(n20042), .A(n20041), .ZN(n20044) );
  OAI211_X1 U23037 ( .C1(n21002), .C2(n20045), .A(n20044), .B(n20049), .ZN(
        P2_U3210) );
  AOI21_X1 U23038 ( .B1(n20048), .B2(n20047), .A(n20046), .ZN(n20053) );
  OAI22_X1 U23039 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n20050), .B1(NA), 
        .B2(n20049), .ZN(n20051) );
  OAI211_X1 U23040 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n20051), .ZN(n20052) );
  OAI21_X1 U23041 ( .B1(n20054), .B2(n20053), .A(n20052), .ZN(P2_U3211) );
  OAI222_X1 U23042 ( .A1(n20109), .A2(n10580), .B1(n20057), .B2(n20178), .C1(
        n20056), .C2(n20106), .ZN(P2_U3212) );
  OAI222_X1 U23043 ( .A1(n20106), .A2(n10580), .B1(n20058), .B2(n20178), .C1(
        n20060), .C2(n20109), .ZN(P2_U3213) );
  OAI222_X1 U23044 ( .A1(n20106), .A2(n20060), .B1(n20059), .B2(n20178), .C1(
        n11123), .C2(n20109), .ZN(P2_U3214) );
  OAI222_X1 U23045 ( .A1(n20109), .A2(n11127), .B1(n20061), .B2(n20178), .C1(
        n11123), .C2(n20106), .ZN(P2_U3215) );
  OAI222_X1 U23046 ( .A1(n20109), .A2(n20063), .B1(n20062), .B2(n20178), .C1(
        n11127), .C2(n20106), .ZN(P2_U3216) );
  OAI222_X1 U23047 ( .A1(n20109), .A2(n20065), .B1(n20064), .B2(n20178), .C1(
        n20063), .C2(n20106), .ZN(P2_U3217) );
  OAI222_X1 U23048 ( .A1(n20109), .A2(n14928), .B1(n20066), .B2(n20178), .C1(
        n20065), .C2(n20106), .ZN(P2_U3218) );
  OAI222_X1 U23049 ( .A1(n20109), .A2(n11142), .B1(n20067), .B2(n20178), .C1(
        n14928), .C2(n20106), .ZN(P2_U3219) );
  OAI222_X1 U23050 ( .A1(n20109), .A2(n20069), .B1(n20068), .B2(n20178), .C1(
        n11142), .C2(n20106), .ZN(P2_U3220) );
  OAI222_X1 U23051 ( .A1(n20109), .A2(n20071), .B1(n20070), .B2(n20178), .C1(
        n20069), .C2(n20106), .ZN(P2_U3221) );
  INV_X1 U23052 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n20073) );
  OAI222_X1 U23053 ( .A1(n20109), .A2(n20073), .B1(n20072), .B2(n20178), .C1(
        n20071), .C2(n20106), .ZN(P2_U3222) );
  OAI222_X1 U23054 ( .A1(n20109), .A2(n11157), .B1(n20074), .B2(n20178), .C1(
        n20073), .C2(n20106), .ZN(P2_U3223) );
  OAI222_X1 U23055 ( .A1(n20109), .A2(n20076), .B1(n20075), .B2(n20178), .C1(
        n11157), .C2(n20106), .ZN(P2_U3224) );
  INV_X1 U23056 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n20078) );
  OAI222_X1 U23057 ( .A1(n20109), .A2(n20078), .B1(n20077), .B2(n20178), .C1(
        n20076), .C2(n20106), .ZN(P2_U3225) );
  OAI222_X1 U23058 ( .A1(n20109), .A2(n14910), .B1(n20079), .B2(n20178), .C1(
        n20078), .C2(n20106), .ZN(P2_U3226) );
  OAI222_X1 U23059 ( .A1(n20109), .A2(n20081), .B1(n20080), .B2(n20178), .C1(
        n14910), .C2(n20106), .ZN(P2_U3227) );
  OAI222_X1 U23060 ( .A1(n20109), .A2(n20083), .B1(n20082), .B2(n20178), .C1(
        n20081), .C2(n20106), .ZN(P2_U3228) );
  OAI222_X1 U23061 ( .A1(n20109), .A2(n20085), .B1(n20084), .B2(n20178), .C1(
        n20083), .C2(n20106), .ZN(P2_U3229) );
  OAI222_X1 U23062 ( .A1(n20109), .A2(n11180), .B1(n20086), .B2(n20178), .C1(
        n20085), .C2(n20106), .ZN(P2_U3230) );
  OAI222_X1 U23063 ( .A1(n20109), .A2(n20088), .B1(n20087), .B2(n20178), .C1(
        n11180), .C2(n20106), .ZN(P2_U3231) );
  INV_X1 U23064 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n20090) );
  OAI222_X1 U23065 ( .A1(n20109), .A2(n20090), .B1(n20089), .B2(n20178), .C1(
        n20088), .C2(n20106), .ZN(P2_U3232) );
  OAI222_X1 U23066 ( .A1(n20109), .A2(n20092), .B1(n20091), .B2(n20178), .C1(
        n20090), .C2(n20106), .ZN(P2_U3233) );
  OAI222_X1 U23067 ( .A1(n20109), .A2(n20094), .B1(n20093), .B2(n20178), .C1(
        n20092), .C2(n20106), .ZN(P2_U3234) );
  OAI222_X1 U23068 ( .A1(n20109), .A2(n20096), .B1(n20095), .B2(n20178), .C1(
        n20094), .C2(n20106), .ZN(P2_U3235) );
  OAI222_X1 U23069 ( .A1(n20109), .A2(n20098), .B1(n20097), .B2(n20178), .C1(
        n20096), .C2(n20106), .ZN(P2_U3236) );
  OAI222_X1 U23070 ( .A1(n20109), .A2(n20101), .B1(n20099), .B2(n20178), .C1(
        n20098), .C2(n20106), .ZN(P2_U3237) );
  OAI222_X1 U23071 ( .A1(n20106), .A2(n20101), .B1(n20100), .B2(n20178), .C1(
        n20102), .C2(n20109), .ZN(P2_U3238) );
  OAI222_X1 U23072 ( .A1(n20109), .A2(n20104), .B1(n20103), .B2(n20178), .C1(
        n20102), .C2(n20106), .ZN(P2_U3239) );
  OAI222_X1 U23073 ( .A1(n20109), .A2(n20107), .B1(n20105), .B2(n20178), .C1(
        n20104), .C2(n20106), .ZN(P2_U3240) );
  INV_X1 U23074 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20108) );
  OAI222_X1 U23075 ( .A1(n20109), .A2(n16162), .B1(n20108), .B2(n20178), .C1(
        n20107), .C2(n20106), .ZN(P2_U3241) );
  INV_X1 U23076 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n20110) );
  AOI22_X1 U23077 ( .A1(n20178), .A2(n20111), .B1(n20110), .B2(n20175), .ZN(
        P2_U3585) );
  MUX2_X1 U23078 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n20178), .Z(P2_U3586) );
  INV_X1 U23079 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n20112) );
  AOI22_X1 U23080 ( .A1(n20178), .A2(n20113), .B1(n20112), .B2(n20175), .ZN(
        P2_U3587) );
  INV_X1 U23081 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n20114) );
  AOI22_X1 U23082 ( .A1(n20178), .A2(n20115), .B1(n20114), .B2(n20175), .ZN(
        P2_U3588) );
  OAI21_X1 U23083 ( .B1(n20119), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20117), 
        .ZN(n20116) );
  INV_X1 U23084 ( .A(n20116), .ZN(P2_U3591) );
  OAI21_X1 U23085 ( .B1(n20119), .B2(n20118), .A(n20117), .ZN(P2_U3592) );
  OAI22_X1 U23086 ( .A1(n20122), .A2(n20121), .B1(n20128), .B2(n20120), .ZN(
        n20124) );
  MUX2_X1 U23087 ( .A(n20124), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n20123), .Z(P2_U3596) );
  NAND2_X1 U23088 ( .A1(n20125), .A2(n20126), .ZN(n20135) );
  NAND2_X1 U23089 ( .A1(n20126), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20151) );
  OR2_X1 U23090 ( .A1(n20127), .A2(n20151), .ZN(n20141) );
  NAND2_X1 U23091 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n20128), .ZN(n20129) );
  OR2_X1 U23092 ( .A1(n20130), .A2(n20129), .ZN(n20131) );
  NAND2_X1 U23093 ( .A1(n20131), .A2(n20156), .ZN(n20142) );
  NAND2_X1 U23094 ( .A1(n20141), .A2(n20142), .ZN(n20133) );
  NAND2_X1 U23095 ( .A1(n20133), .A2(n20132), .ZN(n20134) );
  OAI211_X1 U23096 ( .C1(n20137), .C2(n20136), .A(n20135), .B(n20134), .ZN(
        n20138) );
  INV_X1 U23097 ( .A(n20138), .ZN(n20139) );
  AOI22_X1 U23098 ( .A1(n20163), .A2(n20140), .B1(n20139), .B2(n20164), .ZN(
        P2_U3602) );
  OAI21_X1 U23099 ( .B1(n20143), .B2(n20142), .A(n20141), .ZN(n20144) );
  AOI21_X1 U23100 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20145), .A(n20144), 
        .ZN(n20146) );
  AOI22_X1 U23101 ( .A1(n20163), .A2(n20147), .B1(n20146), .B2(n20164), .ZN(
        P2_U3603) );
  INV_X1 U23102 ( .A(n20148), .ZN(n20149) );
  NAND3_X1 U23103 ( .A1(n20152), .A2(n20156), .A3(n20149), .ZN(n20150) );
  OAI21_X1 U23104 ( .B1(n20152), .B2(n20151), .A(n20150), .ZN(n20153) );
  AOI21_X1 U23105 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20154), .A(n20153), 
        .ZN(n20155) );
  AOI22_X1 U23106 ( .A1(n20163), .A2(n16450), .B1(n20155), .B2(n20164), .ZN(
        P2_U3604) );
  INV_X1 U23107 ( .A(n20156), .ZN(n20159) );
  OAI22_X1 U23108 ( .A1(n20160), .A2(n20159), .B1(n20158), .B2(n20157), .ZN(
        n20161) );
  AOI21_X1 U23109 ( .B1(n20165), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20161), 
        .ZN(n20162) );
  OAI22_X1 U23110 ( .A1(n20165), .A2(n20164), .B1(n20163), .B2(n20162), .ZN(
        P2_U3605) );
  INV_X1 U23111 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20166) );
  AOI22_X1 U23112 ( .A1(n20178), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20166), 
        .B2(n20175), .ZN(P2_U3608) );
  AOI22_X1 U23113 ( .A1(n20170), .A2(n20169), .B1(n20168), .B2(n20167), .ZN(
        n20172) );
  OAI21_X1 U23114 ( .B1(n20172), .B2(n11015), .A(n20171), .ZN(n20174) );
  MUX2_X1 U23115 ( .A(P2_MORE_REG_SCAN_IN), .B(n20174), .S(n20173), .Z(
        P2_U3609) );
  INV_X1 U23116 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n20176) );
  AOI22_X1 U23117 ( .A1(n20178), .A2(n20177), .B1(n20176), .B2(n20175), .ZN(
        P2_U3611) );
  NAND2_X1 U23118 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20999), .ZN(n21081) );
  INV_X1 U23119 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n21312) );
  INV_X1 U23120 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20179) );
  OAI21_X1 U23121 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n20179), .A(
        P1_STATE_REG_0__SCAN_IN), .ZN(n21000) );
  NAND2_X1 U23122 ( .A1(n21000), .A2(n21081), .ZN(n21054) );
  OAI21_X1 U23123 ( .B1(n21038), .B2(n21312), .A(n21054), .ZN(P1_U2802) );
  OAI21_X1 U23124 ( .B1(n20181), .B2(n20180), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20182) );
  OAI21_X1 U23125 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20183), .A(n20182), 
        .ZN(P1_U2803) );
  NOR2_X1 U23126 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20185) );
  OAI21_X1 U23127 ( .B1(n20185), .B2(P1_D_C_N_REG_SCAN_IN), .A(n21081), .ZN(
        n20184) );
  OAI21_X1 U23128 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21081), .A(n20184), 
        .ZN(P1_U2804) );
  OAI21_X1 U23129 ( .B1(BS16), .B2(n20185), .A(n21058), .ZN(n21056) );
  OAI21_X1 U23130 ( .B1(n21058), .B2(n20848), .A(n21056), .ZN(P1_U2805) );
  INV_X1 U23131 ( .A(n20186), .ZN(n20188) );
  OAI21_X1 U23132 ( .B1(n20188), .B2(n21319), .A(n20187), .ZN(P1_U2806) );
  NOR4_X1 U23133 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20192) );
  NOR4_X1 U23134 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20191) );
  NOR4_X1 U23135 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20190) );
  NOR4_X1 U23136 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20189) );
  NAND4_X1 U23137 ( .A1(n20192), .A2(n20191), .A3(n20190), .A4(n20189), .ZN(
        n20198) );
  NOR4_X1 U23138 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20196) );
  AOI211_X1 U23139 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20195) );
  NOR4_X1 U23140 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20194) );
  NOR4_X1 U23141 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20193) );
  NAND4_X1 U23142 ( .A1(n20196), .A2(n20195), .A3(n20194), .A4(n20193), .ZN(
        n20197) );
  NOR2_X1 U23143 ( .A1(n20198), .A2(n20197), .ZN(n21061) );
  INV_X1 U23144 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21362) );
  NOR3_X1 U23145 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20200) );
  OAI21_X1 U23146 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20200), .A(n21061), .ZN(
        n20199) );
  OAI21_X1 U23147 ( .B1(n21061), .B2(n21362), .A(n20199), .ZN(P1_U2807) );
  INV_X1 U23148 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21057) );
  AOI21_X1 U23149 ( .B1(n21391), .B2(n21057), .A(n20200), .ZN(n20201) );
  INV_X1 U23150 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21163) );
  INV_X1 U23151 ( .A(n21061), .ZN(n21063) );
  AOI22_X1 U23152 ( .A1(n21061), .A2(n20201), .B1(n21163), .B2(n21063), .ZN(
        P1_U2808) );
  NAND2_X1 U23153 ( .A1(n20250), .A2(n20202), .ZN(n20225) );
  INV_X1 U23154 ( .A(n20203), .ZN(n20212) );
  AOI21_X1 U23155 ( .B1(n20255), .B2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n20270), .ZN(n20205) );
  NAND2_X1 U23156 ( .A1(n20292), .A2(P1_EBX_REG_9__SCAN_IN), .ZN(n20204) );
  OAI211_X1 U23157 ( .C1(n20206), .C2(n20289), .A(n20205), .B(n20204), .ZN(
        n20207) );
  AOI21_X1 U23158 ( .B1(n20208), .B2(n20272), .A(n20207), .ZN(n20209) );
  OAI21_X1 U23159 ( .B1(n20210), .B2(P1_REIP_REG_9__SCAN_IN), .A(n20209), .ZN(
        n20211) );
  AOI21_X1 U23160 ( .B1(n20212), .B2(n20245), .A(n20211), .ZN(n20213) );
  OAI21_X1 U23161 ( .B1(n21381), .B2(n20225), .A(n20213), .ZN(P1_U2831) );
  NOR2_X1 U23162 ( .A1(n20276), .A2(n20227), .ZN(n20230) );
  AOI21_X1 U23163 ( .B1(P1_REIP_REG_7__SCAN_IN), .B2(n20230), .A(
        P1_REIP_REG_8__SCAN_IN), .ZN(n20226) );
  OAI22_X1 U23164 ( .A1(n20215), .A2(n20295), .B1(n20214), .B2(n20289), .ZN(
        n20216) );
  INV_X1 U23165 ( .A(n20216), .ZN(n20224) );
  INV_X1 U23166 ( .A(n20217), .ZN(n20222) );
  NOR2_X1 U23167 ( .A1(n20218), .A2(n10036), .ZN(n20221) );
  OAI21_X1 U23168 ( .B1(n20288), .B2(n20219), .A(n20256), .ZN(n20220) );
  AOI211_X1 U23169 ( .C1(n20222), .C2(n20245), .A(n20221), .B(n20220), .ZN(
        n20223) );
  OAI211_X1 U23170 ( .C1(n20226), .C2(n20225), .A(n20224), .B(n20223), .ZN(
        P1_U2832) );
  OAI21_X1 U23171 ( .B1(n20252), .B2(n20227), .A(n20250), .ZN(n20243) );
  INV_X1 U23172 ( .A(n20228), .ZN(n20229) );
  AOI22_X1 U23173 ( .A1(n20229), .A2(n20254), .B1(n20255), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20233) );
  NAND2_X1 U23174 ( .A1(n20292), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n20232) );
  NAND2_X1 U23175 ( .A1(n21379), .A2(n20230), .ZN(n20231) );
  AND4_X1 U23176 ( .A1(n20233), .A2(n20232), .A3(n20256), .A4(n20231), .ZN(
        n20234) );
  OAI21_X1 U23177 ( .B1(n20235), .B2(n20295), .A(n20234), .ZN(n20236) );
  AOI21_X1 U23178 ( .B1(n20237), .B2(n20245), .A(n20236), .ZN(n20238) );
  OAI21_X1 U23179 ( .B1(n20243), .B2(n21379), .A(n20238), .ZN(P1_U2833) );
  AOI22_X1 U23180 ( .A1(n20239), .A2(n20272), .B1(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n20255), .ZN(n20249) );
  INV_X1 U23181 ( .A(n20240), .ZN(n20241) );
  AOI22_X1 U23182 ( .A1(n20292), .A2(P1_EBX_REG_6__SCAN_IN), .B1(n20241), .B2(
        n20254), .ZN(n20242) );
  OAI21_X1 U23183 ( .B1(n20243), .B2(n21365), .A(n20242), .ZN(n20244) );
  AOI21_X1 U23184 ( .B1(n20246), .B2(n20245), .A(n20244), .ZN(n20248) );
  NAND4_X1 U23185 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n20285), .A3(n20275), 
        .A4(n21365), .ZN(n20247) );
  NAND4_X1 U23186 ( .A1(n20249), .A2(n20248), .A3(n20256), .A4(n20247), .ZN(
        P1_U2834) );
  INV_X1 U23187 ( .A(n20275), .ZN(n20251) );
  OAI21_X1 U23188 ( .B1(n20252), .B2(n20251), .A(n20250), .ZN(n20280) );
  INV_X1 U23189 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n21014) );
  AOI22_X1 U23190 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n20255), .B1(
        n20254), .B2(n20253), .ZN(n20261) );
  NAND2_X1 U23191 ( .A1(n20292), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n20260) );
  NAND2_X1 U23192 ( .A1(n20285), .A2(n20275), .ZN(n20257) );
  OAI21_X1 U23193 ( .B1(P1_REIP_REG_5__SCAN_IN), .B2(n20257), .A(n20256), .ZN(
        n20258) );
  INV_X1 U23194 ( .A(n20258), .ZN(n20259) );
  AND3_X1 U23195 ( .A1(n20261), .A2(n20260), .A3(n20259), .ZN(n20262) );
  OAI21_X1 U23196 ( .B1(n20263), .B2(n20295), .A(n20262), .ZN(n20264) );
  AOI21_X1 U23197 ( .B1(n20265), .B2(n20297), .A(n20264), .ZN(n20266) );
  OAI21_X1 U23198 ( .B1(n20280), .B2(n21014), .A(n20266), .ZN(P1_U2835) );
  OAI22_X1 U23199 ( .A1(n20268), .A2(n20288), .B1(n20267), .B2(n20289), .ZN(
        n20269) );
  AOI211_X1 U23200 ( .C1(n20271), .C2(n20286), .A(n20270), .B(n20269), .ZN(
        n20284) );
  NAND2_X1 U23201 ( .A1(n20273), .A2(n20272), .ZN(n20279) );
  NOR3_X1 U23202 ( .A1(n20276), .A2(n20275), .A3(n20274), .ZN(n20277) );
  AOI21_X1 U23203 ( .B1(n20292), .B2(P1_EBX_REG_4__SCAN_IN), .A(n20277), .ZN(
        n20278) );
  OAI211_X1 U23204 ( .C1(n21332), .C2(n20280), .A(n20279), .B(n20278), .ZN(
        n20281) );
  AOI21_X1 U23205 ( .B1(n20282), .B2(n20297), .A(n20281), .ZN(n20283) );
  NAND2_X1 U23206 ( .A1(n20284), .A2(n20283), .ZN(P1_U2836) );
  AOI21_X1 U23207 ( .B1(n20285), .B2(P1_REIP_REG_1__SCAN_IN), .A(
        P1_REIP_REG_2__SCAN_IN), .ZN(n20300) );
  NAND2_X1 U23208 ( .A1(n20384), .A2(n20286), .ZN(n20294) );
  INV_X1 U23209 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n20287) );
  OAI22_X1 U23210 ( .A1(n20290), .A2(n20289), .B1(n20288), .B2(n20287), .ZN(
        n20291) );
  AOI21_X1 U23211 ( .B1(P1_EBX_REG_2__SCAN_IN), .B2(n20292), .A(n20291), .ZN(
        n20293) );
  OAI211_X1 U23212 ( .C1(n20301), .C2(n20295), .A(n20294), .B(n20293), .ZN(
        n20296) );
  AOI21_X1 U23213 ( .B1(n20304), .B2(n20297), .A(n20296), .ZN(n20298) );
  OAI21_X1 U23214 ( .B1(n20300), .B2(n20299), .A(n20298), .ZN(P1_U2838) );
  INV_X1 U23215 ( .A(n20301), .ZN(n20302) );
  AOI22_X1 U23216 ( .A1(n20304), .A2(n20303), .B1(n13038), .B2(n20302), .ZN(
        n20305) );
  OAI21_X1 U23217 ( .B1(n20306), .B2(n10033), .A(n20305), .ZN(P1_U2870) );
  AOI22_X1 U23218 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20310), .B1(n15849), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20307) );
  OAI21_X1 U23219 ( .B1(n20309), .B2(n20308), .A(n20307), .ZN(P1_U2921) );
  INV_X1 U23220 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20312) );
  AOI22_X1 U23221 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20319), .B1(n15849), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20311) );
  OAI21_X1 U23222 ( .B1(n20312), .B2(n20338), .A(n20311), .ZN(P1_U2922) );
  INV_X1 U23223 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20314) );
  AOI22_X1 U23224 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20319), .B1(n15849), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20313) );
  OAI21_X1 U23225 ( .B1(n20314), .B2(n20338), .A(n20313), .ZN(P1_U2923) );
  AOI22_X1 U23226 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20319), .B1(n15849), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20315) );
  OAI21_X1 U23227 ( .B1(n14528), .B2(n20338), .A(n20315), .ZN(P1_U2924) );
  INV_X1 U23228 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20317) );
  AOI22_X1 U23229 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20319), .B1(n15849), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20316) );
  OAI21_X1 U23230 ( .B1(n20317), .B2(n20338), .A(n20316), .ZN(P1_U2925) );
  AOI22_X1 U23231 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20319), .B1(n15849), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20318) );
  OAI21_X1 U23232 ( .B1(n14217), .B2(n20338), .A(n20318), .ZN(P1_U2926) );
  INV_X1 U23233 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20321) );
  AOI22_X1 U23234 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20319), .B1(n15849), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20320) );
  OAI21_X1 U23235 ( .B1(n20321), .B2(n20338), .A(n20320), .ZN(P1_U2927) );
  AOI22_X1 U23236 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20336), .B1(n15849), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20322) );
  OAI21_X1 U23237 ( .B1(n20323), .B2(n20338), .A(n20322), .ZN(P1_U2928) );
  AOI22_X1 U23238 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20336), .B1(n15849), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20324) );
  OAI21_X1 U23239 ( .B1(n12206), .B2(n20338), .A(n20324), .ZN(P1_U2929) );
  AOI22_X1 U23240 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20336), .B1(n15849), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20325) );
  OAI21_X1 U23241 ( .B1(n12197), .B2(n20338), .A(n20325), .ZN(P1_U2930) );
  AOI22_X1 U23242 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20336), .B1(n15849), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20326) );
  OAI21_X1 U23243 ( .B1(n20327), .B2(n20338), .A(n20326), .ZN(P1_U2931) );
  AOI22_X1 U23244 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20336), .B1(n15849), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20328) );
  OAI21_X1 U23245 ( .B1(n20329), .B2(n20338), .A(n20328), .ZN(P1_U2932) );
  AOI22_X1 U23246 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20336), .B1(n15849), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20330) );
  OAI21_X1 U23247 ( .B1(n20331), .B2(n20338), .A(n20330), .ZN(P1_U2933) );
  AOI22_X1 U23248 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20336), .B1(n15849), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20332) );
  OAI21_X1 U23249 ( .B1(n20333), .B2(n20338), .A(n20332), .ZN(P1_U2934) );
  AOI22_X1 U23250 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20336), .B1(n15849), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20334) );
  OAI21_X1 U23251 ( .B1(n20335), .B2(n20338), .A(n20334), .ZN(P1_U2935) );
  AOI22_X1 U23252 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20336), .B1(n15849), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20337) );
  OAI21_X1 U23253 ( .B1(n20339), .B2(n20338), .A(n20337), .ZN(P1_U2936) );
  AOI22_X1 U23254 ( .A1(n20351), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20348), .ZN(n20341) );
  NAND2_X1 U23255 ( .A1(n20341), .A2(n20340), .ZN(P1_U2961) );
  AOI22_X1 U23256 ( .A1(n20351), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20348), .ZN(n20343) );
  NAND2_X1 U23257 ( .A1(n20343), .A2(n20342), .ZN(P1_U2962) );
  AOI22_X1 U23258 ( .A1(n20351), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20348), .ZN(n20345) );
  NAND2_X1 U23259 ( .A1(n20345), .A2(n20344), .ZN(P1_U2963) );
  AOI22_X1 U23260 ( .A1(n20351), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20348), .ZN(n20347) );
  NAND2_X1 U23261 ( .A1(n20347), .A2(n20346), .ZN(P1_U2964) );
  AOI22_X1 U23262 ( .A1(n20351), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20348), .ZN(n20350) );
  NAND2_X1 U23263 ( .A1(n20350), .A2(n20349), .ZN(P1_U2965) );
  AOI22_X1 U23264 ( .A1(n20351), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20348), .ZN(n20353) );
  NAND2_X1 U23265 ( .A1(n20353), .A2(n20352), .ZN(P1_U2966) );
  NOR2_X1 U23266 ( .A1(n20355), .A2(n20354), .ZN(n20356) );
  AOI21_X1 U23267 ( .B1(n20358), .B2(n20357), .A(n20356), .ZN(n20368) );
  INV_X1 U23268 ( .A(n20359), .ZN(n20365) );
  INV_X1 U23269 ( .A(n20360), .ZN(n20363) );
  NAND3_X1 U23270 ( .A1(n20363), .A2(n20362), .A3(n20361), .ZN(n20364) );
  OAI21_X1 U23271 ( .B1(n20366), .B2(n20365), .A(n20364), .ZN(n20367) );
  OAI211_X1 U23272 ( .C1(n13697), .C2(n20369), .A(n20368), .B(n20367), .ZN(
        P1_U3031) );
  NOR2_X1 U23273 ( .A1(n20371), .A2(n20370), .ZN(P1_U3032) );
  INV_X1 U23274 ( .A(DATAI_16_), .ZN(n21347) );
  OAI22_X1 U23275 ( .A1(n21347), .A2(n20441), .B1(n20375), .B2(n20440), .ZN(
        n20852) );
  INV_X1 U23276 ( .A(n20479), .ZN(n20377) );
  INV_X1 U23277 ( .A(DATAI_24_), .ZN(n21366) );
  OAI22_X1 U23278 ( .A1(n21366), .A2(n20441), .B1(n20378), .B2(n20440), .ZN(
        n20935) );
  INV_X1 U23279 ( .A(n20935), .ZN(n20855) );
  NAND2_X1 U23280 ( .A1(n20444), .A2(n20380), .ZN(n20792) );
  NAND3_X1 U23281 ( .A1(n12729), .A2(n12753), .A3(n20791), .ZN(n20453) );
  OR2_X1 U23282 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20453), .ZN(
        n20445) );
  OAI22_X1 U23283 ( .A1(n20986), .A2(n20855), .B1(n20792), .B2(n20445), .ZN(
        n20381) );
  INV_X1 U23284 ( .A(n20381), .ZN(n20393) );
  INV_X1 U23285 ( .A(n20477), .ZN(n20382) );
  OAI21_X1 U23286 ( .B1(n20382), .B2(n20966), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20383) );
  NAND2_X1 U23287 ( .A1(n20383), .A2(n20933), .ZN(n20391) );
  OR2_X1 U23288 ( .A1(n20659), .A2(n20384), .ZN(n20509) );
  NOR2_X1 U23289 ( .A1(n20509), .A2(n20881), .ZN(n20388) );
  INV_X1 U23290 ( .A(n20389), .ZN(n20385) );
  NOR2_X1 U23291 ( .A1(n20385), .A2(n20991), .ZN(n20790) );
  NAND2_X1 U23292 ( .A1(n20719), .A2(n20661), .ZN(n20538) );
  AOI22_X1 U23293 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20538), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n20445), .ZN(n20386) );
  OAI211_X1 U23294 ( .C1(n20391), .C2(n20388), .A(n20721), .B(n20386), .ZN(
        n20449) );
  INV_X1 U23295 ( .A(n20388), .ZN(n20390) );
  NOR2_X1 U23296 ( .A1(n20389), .A2(n20991), .ZN(n20714) );
  INV_X1 U23297 ( .A(n20714), .ZN(n20663) );
  AOI22_X1 U23298 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20449), .B1(
        n20923), .B2(n20448), .ZN(n20392) );
  OAI211_X1 U23299 ( .C1(n20938), .C2(n20477), .A(n20393), .B(n20392), .ZN(
        P1_U3033) );
  INV_X1 U23300 ( .A(DATAI_17_), .ZN(n21160) );
  OAI22_X1 U23301 ( .A1(n20394), .A2(n20440), .B1(n21160), .B2(n20441), .ZN(
        n20941) );
  INV_X1 U23302 ( .A(n20941), .ZN(n20895) );
  INV_X1 U23303 ( .A(DATAI_25_), .ZN(n20396) );
  OAI22_X1 U23304 ( .A1(n20396), .A2(n20441), .B1(n20395), .B2(n20440), .ZN(
        n20892) );
  INV_X1 U23305 ( .A(n20892), .ZN(n20944) );
  NAND2_X1 U23306 ( .A1(n20444), .A2(n11917), .ZN(n20804) );
  OAI22_X1 U23307 ( .A1(n20986), .A2(n20944), .B1(n20804), .B2(n20445), .ZN(
        n20397) );
  INV_X1 U23308 ( .A(n20397), .ZN(n20400) );
  AOI22_X1 U23309 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20449), .B1(
        n20939), .B2(n20448), .ZN(n20399) );
  OAI211_X1 U23310 ( .C1(n20895), .C2(n20477), .A(n20400), .B(n20399), .ZN(
        P1_U3034) );
  INV_X1 U23311 ( .A(DATAI_18_), .ZN(n20402) );
  OAI22_X1 U23312 ( .A1(n20402), .A2(n20441), .B1(n20401), .B2(n20440), .ZN(
        n20947) );
  INV_X1 U23313 ( .A(n20947), .ZN(n20899) );
  INV_X1 U23314 ( .A(DATAI_26_), .ZN(n20403) );
  OAI22_X1 U23315 ( .A1(n20404), .A2(n20440), .B1(n20403), .B2(n20441), .ZN(
        n20896) );
  INV_X1 U23316 ( .A(n20896), .ZN(n20950) );
  NAND2_X1 U23317 ( .A1(n20444), .A2(n20405), .ZN(n20809) );
  OAI22_X1 U23318 ( .A1(n20986), .A2(n20950), .B1(n20809), .B2(n20445), .ZN(
        n20406) );
  INV_X1 U23319 ( .A(n20406), .ZN(n20409) );
  AOI22_X1 U23320 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20449), .B1(
        n20945), .B2(n20448), .ZN(n20408) );
  OAI211_X1 U23321 ( .C1(n20899), .C2(n20477), .A(n20409), .B(n20408), .ZN(
        P1_U3035) );
  INV_X1 U23322 ( .A(DATAI_19_), .ZN(n21331) );
  OAI22_X1 U23323 ( .A1(n21331), .A2(n20441), .B1(n20410), .B2(n20440), .ZN(
        n20860) );
  INV_X1 U23324 ( .A(DATAI_27_), .ZN(n20411) );
  OAI22_X1 U23325 ( .A1(n20412), .A2(n20440), .B1(n20411), .B2(n20441), .ZN(
        n20953) );
  INV_X1 U23326 ( .A(n20953), .ZN(n20863) );
  NAND2_X1 U23327 ( .A1(n20444), .A2(n20413), .ZN(n20814) );
  OAI22_X1 U23328 ( .A1(n20986), .A2(n20863), .B1(n20814), .B2(n20445), .ZN(
        n20414) );
  INV_X1 U23329 ( .A(n20414), .ZN(n20417) );
  AOI22_X1 U23330 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20449), .B1(
        n20951), .B2(n20448), .ZN(n20416) );
  OAI211_X1 U23331 ( .C1(n20956), .C2(n20477), .A(n20417), .B(n20416), .ZN(
        P1_U3036) );
  INV_X1 U23332 ( .A(DATAI_20_), .ZN(n20419) );
  OAI22_X1 U23333 ( .A1(n20419), .A2(n20441), .B1(n20418), .B2(n20440), .ZN(
        n20959) );
  INV_X1 U23334 ( .A(n20959), .ZN(n20905) );
  INV_X1 U23335 ( .A(DATAI_28_), .ZN(n21146) );
  OAI22_X1 U23336 ( .A1(n20420), .A2(n20440), .B1(n21146), .B2(n20441), .ZN(
        n20902) );
  INV_X1 U23337 ( .A(n20902), .ZN(n20962) );
  NAND2_X1 U23338 ( .A1(n20444), .A2(n13773), .ZN(n20819) );
  OAI22_X1 U23339 ( .A1(n20986), .A2(n20962), .B1(n20819), .B2(n20445), .ZN(
        n20421) );
  INV_X1 U23340 ( .A(n20421), .ZN(n20424) );
  AOI22_X1 U23341 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20449), .B1(
        n20957), .B2(n20448), .ZN(n20423) );
  OAI211_X1 U23342 ( .C1(n20905), .C2(n20477), .A(n20424), .B(n20423), .ZN(
        P1_U3037) );
  INV_X1 U23343 ( .A(DATAI_21_), .ZN(n20426) );
  OAI22_X1 U23344 ( .A1(n20426), .A2(n20441), .B1(n20425), .B2(n20440), .ZN(
        n20965) );
  INV_X1 U23345 ( .A(DATAI_29_), .ZN(n21275) );
  OAI22_X1 U23346 ( .A1(n20427), .A2(n20440), .B1(n21275), .B2(n20441), .ZN(
        n20906) );
  INV_X1 U23347 ( .A(n20906), .ZN(n20970) );
  NAND2_X1 U23348 ( .A1(n20444), .A2(n11926), .ZN(n20824) );
  OAI22_X1 U23349 ( .A1(n20986), .A2(n20970), .B1(n20824), .B2(n20445), .ZN(
        n20428) );
  INV_X1 U23350 ( .A(n20428), .ZN(n20431) );
  AOI22_X1 U23351 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20449), .B1(
        n20963), .B2(n20448), .ZN(n20430) );
  OAI211_X1 U23352 ( .C1(n20909), .C2(n20477), .A(n20431), .B(n20430), .ZN(
        P1_U3038) );
  INV_X1 U23353 ( .A(DATAI_22_), .ZN(n20433) );
  OAI22_X1 U23354 ( .A1(n20433), .A2(n20441), .B1(n20432), .B2(n20440), .ZN(
        n20868) );
  INV_X1 U23355 ( .A(n20868), .ZN(n20976) );
  INV_X1 U23356 ( .A(DATAI_30_), .ZN(n21178) );
  OAI22_X1 U23357 ( .A1(n20434), .A2(n20440), .B1(n21178), .B2(n20441), .ZN(
        n20973) );
  INV_X1 U23358 ( .A(n20973), .ZN(n20871) );
  NAND2_X1 U23359 ( .A1(n20444), .A2(n11928), .ZN(n20829) );
  OAI22_X1 U23360 ( .A1(n20986), .A2(n20871), .B1(n20829), .B2(n20445), .ZN(
        n20435) );
  INV_X1 U23361 ( .A(n20435), .ZN(n20438) );
  AOI22_X1 U23362 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20449), .B1(
        n20971), .B2(n20448), .ZN(n20437) );
  OAI211_X1 U23363 ( .C1(n20976), .C2(n20477), .A(n20438), .B(n20437), .ZN(
        P1_U3039) );
  INV_X1 U23364 ( .A(DATAI_23_), .ZN(n21122) );
  OAI22_X1 U23365 ( .A1(n21122), .A2(n20441), .B1(n20439), .B2(n20440), .ZN(
        n20874) );
  INV_X1 U23366 ( .A(n20874), .ZN(n20987) );
  INV_X1 U23367 ( .A(DATAI_31_), .ZN(n20442) );
  OAI22_X1 U23368 ( .A1(n20442), .A2(n20441), .B1(n13065), .B2(n20440), .ZN(
        n20981) );
  INV_X1 U23369 ( .A(n20981), .ZN(n20879) );
  NAND2_X1 U23370 ( .A1(n20444), .A2(n20443), .ZN(n20835) );
  OAI22_X1 U23371 ( .A1(n20986), .A2(n20879), .B1(n20835), .B2(n20445), .ZN(
        n20446) );
  INV_X1 U23372 ( .A(n20446), .ZN(n20451) );
  AOI22_X1 U23373 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20449), .B1(
        n20978), .B2(n20448), .ZN(n20450) );
  OAI211_X1 U23374 ( .C1(n20987), .C2(n20477), .A(n20451), .B(n20450), .ZN(
        P1_U3040) );
  NOR2_X1 U23375 ( .A1(n20843), .A2(n20453), .ZN(n20473) );
  INV_X1 U23376 ( .A(n20509), .ZN(n20452) );
  INV_X1 U23377 ( .A(n20565), .ZN(n20845) );
  AOI21_X1 U23378 ( .B1(n20452), .B2(n20845), .A(n20473), .ZN(n20454) );
  OAI22_X1 U23379 ( .A1(n20454), .A2(n20926), .B1(n20453), .B2(n20991), .ZN(
        n20472) );
  AOI22_X1 U23380 ( .A1(n20924), .A2(n20473), .B1(n20472), .B2(n20923), .ZN(
        n20459) );
  INV_X1 U23381 ( .A(n20453), .ZN(n20456) );
  INV_X1 U23382 ( .A(n20480), .ZN(n20512) );
  OAI211_X1 U23383 ( .C1(n20512), .C2(n20848), .A(n20933), .B(n20454), .ZN(
        n20455) );
  OAI211_X1 U23384 ( .C1(n20933), .C2(n20456), .A(n20932), .B(n20455), .ZN(
        n20474) );
  INV_X1 U23385 ( .A(n20851), .ZN(n20457) );
  AOI22_X1 U23386 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20474), .B1(
        n20502), .B2(n20852), .ZN(n20458) );
  OAI211_X1 U23387 ( .C1(n20855), .C2(n20477), .A(n20459), .B(n20458), .ZN(
        P1_U3041) );
  AOI22_X1 U23388 ( .A1(n20940), .A2(n20473), .B1(n20472), .B2(n20939), .ZN(
        n20461) );
  AOI22_X1 U23389 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20474), .B1(
        n20502), .B2(n20941), .ZN(n20460) );
  OAI211_X1 U23390 ( .C1(n20944), .C2(n20477), .A(n20461), .B(n20460), .ZN(
        P1_U3042) );
  AOI22_X1 U23391 ( .A1(n20946), .A2(n20473), .B1(n20472), .B2(n20945), .ZN(
        n20463) );
  AOI22_X1 U23392 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20474), .B1(
        n20502), .B2(n20947), .ZN(n20462) );
  OAI211_X1 U23393 ( .C1(n20950), .C2(n20477), .A(n20463), .B(n20462), .ZN(
        P1_U3043) );
  AOI22_X1 U23394 ( .A1(n20952), .A2(n20473), .B1(n20472), .B2(n20951), .ZN(
        n20465) );
  AOI22_X1 U23395 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20474), .B1(
        n20502), .B2(n20860), .ZN(n20464) );
  OAI211_X1 U23396 ( .C1(n20863), .C2(n20477), .A(n20465), .B(n20464), .ZN(
        P1_U3044) );
  AOI22_X1 U23397 ( .A1(n20958), .A2(n20473), .B1(n20472), .B2(n20957), .ZN(
        n20467) );
  AOI22_X1 U23398 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20474), .B1(
        n20502), .B2(n20959), .ZN(n20466) );
  OAI211_X1 U23399 ( .C1(n20962), .C2(n20477), .A(n20467), .B(n20466), .ZN(
        P1_U3045) );
  AOI22_X1 U23400 ( .A1(n20964), .A2(n20473), .B1(n20472), .B2(n20963), .ZN(
        n20469) );
  AOI22_X1 U23401 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20474), .B1(
        n20502), .B2(n20965), .ZN(n20468) );
  OAI211_X1 U23402 ( .C1(n20970), .C2(n20477), .A(n20469), .B(n20468), .ZN(
        P1_U3046) );
  AOI22_X1 U23403 ( .A1(n20972), .A2(n20473), .B1(n20472), .B2(n20971), .ZN(
        n20471) );
  AOI22_X1 U23404 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20474), .B1(
        n20502), .B2(n20868), .ZN(n20470) );
  OAI211_X1 U23405 ( .C1(n20871), .C2(n20477), .A(n20471), .B(n20470), .ZN(
        P1_U3047) );
  AOI22_X1 U23406 ( .A1(n20980), .A2(n20473), .B1(n20978), .B2(n20472), .ZN(
        n20476) );
  AOI22_X1 U23407 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20474), .B1(
        n20502), .B2(n20874), .ZN(n20475) );
  OAI211_X1 U23408 ( .C1(n20879), .C2(n20477), .A(n20476), .B(n20475), .ZN(
        P1_U3048) );
  INV_X1 U23409 ( .A(n20502), .ZN(n20478) );
  NAND2_X1 U23410 ( .A1(n20478), .A2(n20933), .ZN(n20481) );
  OAI21_X1 U23411 ( .B1(n20481), .B2(n20532), .A(n20786), .ZN(n20482) );
  NOR2_X1 U23412 ( .A1(n20509), .A2(n20660), .ZN(n20485) );
  NAND3_X1 U23413 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n12729), .A3(
        n12753), .ZN(n20513) );
  NOR2_X1 U23414 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20513), .ZN(
        n20501) );
  AOI22_X1 U23415 ( .A1(n20502), .A2(n20935), .B1(n20924), .B2(n20501), .ZN(
        n20488) );
  INV_X1 U23416 ( .A(n20482), .ZN(n20486) );
  INV_X1 U23417 ( .A(n20501), .ZN(n20483) );
  NOR2_X1 U23418 ( .A1(n10383), .A2(n20991), .ZN(n20595) );
  AOI21_X1 U23419 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20483), .A(n20595), 
        .ZN(n20484) );
  OAI211_X1 U23420 ( .C1(n20486), .C2(n20485), .A(n20721), .B(n20484), .ZN(
        n20503) );
  AOI22_X1 U23421 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20503), .B1(
        n20532), .B2(n20852), .ZN(n20487) );
  OAI211_X1 U23422 ( .C1(n20506), .C2(n20803), .A(n20488), .B(n20487), .ZN(
        P1_U3049) );
  INV_X1 U23423 ( .A(n20939), .ZN(n20808) );
  AOI22_X1 U23424 ( .A1(n20502), .A2(n20892), .B1(n20940), .B2(n20501), .ZN(
        n20490) );
  AOI22_X1 U23425 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20503), .B1(
        n20532), .B2(n20941), .ZN(n20489) );
  OAI211_X1 U23426 ( .C1(n20506), .C2(n20808), .A(n20490), .B(n20489), .ZN(
        P1_U3050) );
  INV_X1 U23427 ( .A(n20945), .ZN(n20813) );
  AOI22_X1 U23428 ( .A1(n20502), .A2(n20896), .B1(n20946), .B2(n20501), .ZN(
        n20492) );
  AOI22_X1 U23429 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20503), .B1(
        n20532), .B2(n20947), .ZN(n20491) );
  OAI211_X1 U23430 ( .C1(n20506), .C2(n20813), .A(n20492), .B(n20491), .ZN(
        P1_U3051) );
  INV_X1 U23431 ( .A(n20951), .ZN(n20818) );
  AOI22_X1 U23432 ( .A1(n20502), .A2(n20953), .B1(n20952), .B2(n20501), .ZN(
        n20494) );
  AOI22_X1 U23433 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20503), .B1(
        n20532), .B2(n20860), .ZN(n20493) );
  OAI211_X1 U23434 ( .C1(n20506), .C2(n20818), .A(n20494), .B(n20493), .ZN(
        P1_U3052) );
  INV_X1 U23435 ( .A(n20957), .ZN(n20823) );
  AOI22_X1 U23436 ( .A1(n20532), .A2(n20959), .B1(n20958), .B2(n20501), .ZN(
        n20496) );
  AOI22_X1 U23437 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20503), .B1(
        n20502), .B2(n20902), .ZN(n20495) );
  OAI211_X1 U23438 ( .C1(n20506), .C2(n20823), .A(n20496), .B(n20495), .ZN(
        P1_U3053) );
  AOI22_X1 U23439 ( .A1(n20532), .A2(n20965), .B1(n20964), .B2(n20501), .ZN(
        n20498) );
  AOI22_X1 U23440 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20503), .B1(
        n20502), .B2(n20906), .ZN(n20497) );
  OAI211_X1 U23441 ( .C1(n20506), .C2(n20828), .A(n20498), .B(n20497), .ZN(
        P1_U3054) );
  INV_X1 U23442 ( .A(n20971), .ZN(n20833) );
  AOI22_X1 U23443 ( .A1(n20532), .A2(n20868), .B1(n20972), .B2(n20501), .ZN(
        n20500) );
  AOI22_X1 U23444 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20503), .B1(
        n20502), .B2(n20973), .ZN(n20499) );
  OAI211_X1 U23445 ( .C1(n20506), .C2(n20833), .A(n20500), .B(n20499), .ZN(
        P1_U3055) );
  INV_X1 U23446 ( .A(n20978), .ZN(n20841) );
  AOI22_X1 U23447 ( .A1(n20502), .A2(n20981), .B1(n20980), .B2(n20501), .ZN(
        n20505) );
  AOI22_X1 U23448 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20503), .B1(
        n20532), .B2(n20874), .ZN(n20504) );
  OAI211_X1 U23449 ( .C1(n20506), .C2(n20841), .A(n20505), .B(n20504), .ZN(
        P1_U3056) );
  INV_X1 U23450 ( .A(n20513), .ZN(n20511) );
  NAND2_X1 U23451 ( .A1(n12075), .A2(n20507), .ZN(n20919) );
  NOR2_X1 U23452 ( .A1(n20752), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20531) );
  INV_X1 U23453 ( .A(n20531), .ZN(n20508) );
  OAI21_X1 U23454 ( .B1(n20509), .B2(n20919), .A(n20508), .ZN(n20515) );
  AOI21_X1 U23455 ( .B1(n20512), .B2(n20933), .A(n20929), .ZN(n20516) );
  INV_X1 U23456 ( .A(n20516), .ZN(n20510) );
  AOI22_X1 U23457 ( .A1(n20560), .A2(n20852), .B1(n20924), .B2(n20531), .ZN(
        n20518) );
  INV_X1 U23458 ( .A(n20932), .ZN(n20757) );
  AOI21_X1 U23459 ( .B1(n20926), .B2(n20513), .A(n20757), .ZN(n20514) );
  OAI21_X1 U23460 ( .B1(n20516), .B2(n20515), .A(n20514), .ZN(n20533) );
  AOI22_X1 U23461 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20533), .B1(
        n20532), .B2(n20935), .ZN(n20517) );
  OAI211_X1 U23462 ( .C1(n20536), .C2(n20803), .A(n20518), .B(n20517), .ZN(
        P1_U3057) );
  AOI22_X1 U23463 ( .A1(n20560), .A2(n20941), .B1(n20940), .B2(n20531), .ZN(
        n20520) );
  AOI22_X1 U23464 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20533), .B1(
        n20532), .B2(n20892), .ZN(n20519) );
  OAI211_X1 U23465 ( .C1(n20536), .C2(n20808), .A(n20520), .B(n20519), .ZN(
        P1_U3058) );
  AOI22_X1 U23466 ( .A1(n20560), .A2(n20947), .B1(n20946), .B2(n20531), .ZN(
        n20522) );
  AOI22_X1 U23467 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20533), .B1(
        n20532), .B2(n20896), .ZN(n20521) );
  OAI211_X1 U23468 ( .C1(n20536), .C2(n20813), .A(n20522), .B(n20521), .ZN(
        P1_U3059) );
  AOI22_X1 U23469 ( .A1(n20560), .A2(n20860), .B1(n20952), .B2(n20531), .ZN(
        n20524) );
  AOI22_X1 U23470 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20533), .B1(
        n20532), .B2(n20953), .ZN(n20523) );
  OAI211_X1 U23471 ( .C1(n20536), .C2(n20818), .A(n20524), .B(n20523), .ZN(
        P1_U3060) );
  AOI22_X1 U23472 ( .A1(n20560), .A2(n20959), .B1(n20958), .B2(n20531), .ZN(
        n20526) );
  AOI22_X1 U23473 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20533), .B1(
        n20532), .B2(n20902), .ZN(n20525) );
  OAI211_X1 U23474 ( .C1(n20536), .C2(n20823), .A(n20526), .B(n20525), .ZN(
        P1_U3061) );
  AOI22_X1 U23475 ( .A1(n20560), .A2(n20965), .B1(n20964), .B2(n20531), .ZN(
        n20528) );
  AOI22_X1 U23476 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20533), .B1(
        n20532), .B2(n20906), .ZN(n20527) );
  OAI211_X1 U23477 ( .C1(n20536), .C2(n20828), .A(n20528), .B(n20527), .ZN(
        P1_U3062) );
  AOI22_X1 U23478 ( .A1(n20532), .A2(n20973), .B1(n20972), .B2(n20531), .ZN(
        n20530) );
  AOI22_X1 U23479 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20533), .B1(
        n20560), .B2(n20868), .ZN(n20529) );
  OAI211_X1 U23480 ( .C1(n20536), .C2(n20833), .A(n20530), .B(n20529), .ZN(
        P1_U3063) );
  AOI22_X1 U23481 ( .A1(n20532), .A2(n20981), .B1(n20980), .B2(n20531), .ZN(
        n20535) );
  AOI22_X1 U23482 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20533), .B1(
        n20560), .B2(n20874), .ZN(n20534) );
  OAI211_X1 U23483 ( .C1(n20536), .C2(n20841), .A(n20535), .B(n20534), .ZN(
        P1_U3064) );
  NAND3_X1 U23484 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n12729), .A3(
        n20791), .ZN(n20567) );
  NOR2_X1 U23485 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20567), .ZN(
        n20559) );
  NOR2_X1 U23486 ( .A1(n13909), .A2(n20537), .ZN(n20592) );
  NAND2_X1 U23487 ( .A1(n20592), .A2(n20933), .ZN(n20632) );
  INV_X1 U23488 ( .A(n20790), .ZN(n20883) );
  OAI22_X1 U23489 ( .A1(n20632), .A2(n20881), .B1(n20538), .B2(n20883), .ZN(
        n20558) );
  AOI22_X1 U23490 ( .A1(n20924), .A2(n20559), .B1(n20923), .B2(n20558), .ZN(
        n20545) );
  INV_X1 U23491 ( .A(n20560), .ZN(n20539) );
  AOI21_X1 U23492 ( .B1(n20539), .B2(n20589), .A(n20848), .ZN(n20540) );
  AOI21_X1 U23493 ( .B1(n20592), .B2(n20660), .A(n20540), .ZN(n20541) );
  NOR2_X1 U23494 ( .A1(n20541), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20543) );
  AOI22_X1 U23495 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20561), .B1(
        n20560), .B2(n20935), .ZN(n20544) );
  OAI211_X1 U23496 ( .C1(n20938), .C2(n20589), .A(n20545), .B(n20544), .ZN(
        P1_U3065) );
  AOI22_X1 U23497 ( .A1(n20940), .A2(n20559), .B1(n20939), .B2(n20558), .ZN(
        n20547) );
  AOI22_X1 U23498 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20561), .B1(
        n20560), .B2(n20892), .ZN(n20546) );
  OAI211_X1 U23499 ( .C1(n20895), .C2(n20589), .A(n20547), .B(n20546), .ZN(
        P1_U3066) );
  AOI22_X1 U23500 ( .A1(n20946), .A2(n20559), .B1(n20945), .B2(n20558), .ZN(
        n20549) );
  AOI22_X1 U23501 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20561), .B1(
        n20560), .B2(n20896), .ZN(n20548) );
  OAI211_X1 U23502 ( .C1(n20899), .C2(n20589), .A(n20549), .B(n20548), .ZN(
        P1_U3067) );
  AOI22_X1 U23503 ( .A1(n20952), .A2(n20559), .B1(n20951), .B2(n20558), .ZN(
        n20551) );
  AOI22_X1 U23504 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20561), .B1(
        n20560), .B2(n20953), .ZN(n20550) );
  OAI211_X1 U23505 ( .C1(n20956), .C2(n20589), .A(n20551), .B(n20550), .ZN(
        P1_U3068) );
  AOI22_X1 U23506 ( .A1(n20958), .A2(n20559), .B1(n20957), .B2(n20558), .ZN(
        n20553) );
  AOI22_X1 U23507 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20561), .B1(
        n20560), .B2(n20902), .ZN(n20552) );
  OAI211_X1 U23508 ( .C1(n20905), .C2(n20589), .A(n20553), .B(n20552), .ZN(
        P1_U3069) );
  AOI22_X1 U23509 ( .A1(n20964), .A2(n20559), .B1(n20963), .B2(n20558), .ZN(
        n20555) );
  AOI22_X1 U23510 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20561), .B1(
        n20560), .B2(n20906), .ZN(n20554) );
  OAI211_X1 U23511 ( .C1(n20909), .C2(n20589), .A(n20555), .B(n20554), .ZN(
        P1_U3070) );
  AOI22_X1 U23512 ( .A1(n20972), .A2(n20559), .B1(n20971), .B2(n20558), .ZN(
        n20557) );
  AOI22_X1 U23513 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20561), .B1(
        n20560), .B2(n20973), .ZN(n20556) );
  OAI211_X1 U23514 ( .C1(n20976), .C2(n20589), .A(n20557), .B(n20556), .ZN(
        P1_U3071) );
  AOI22_X1 U23515 ( .A1(n20980), .A2(n20559), .B1(n20978), .B2(n20558), .ZN(
        n20563) );
  AOI22_X1 U23516 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20561), .B1(
        n20560), .B2(n20981), .ZN(n20562) );
  OAI211_X1 U23517 ( .C1(n20987), .C2(n20589), .A(n20563), .B(n20562), .ZN(
        P1_U3072) );
  NOR2_X1 U23518 ( .A1(n20843), .A2(n20567), .ZN(n20585) );
  INV_X1 U23519 ( .A(n20585), .ZN(n20564) );
  OAI222_X1 U23520 ( .A1(n20632), .A2(n20565), .B1(n20564), .B2(n20926), .C1(
        n20991), .C2(n20567), .ZN(n20584) );
  AOI22_X1 U23521 ( .A1(n20924), .A2(n20585), .B1(n20923), .B2(n20584), .ZN(
        n20571) );
  INV_X1 U23522 ( .A(n20629), .ZN(n20566) );
  NAND2_X1 U23523 ( .A1(n20566), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20634) );
  NOR2_X1 U23524 ( .A1(n20634), .A2(n20926), .ZN(n20569) );
  INV_X1 U23525 ( .A(n20567), .ZN(n20568) );
  OAI21_X1 U23526 ( .B1(n20569), .B2(n20568), .A(n20932), .ZN(n20586) );
  AOI22_X1 U23527 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20586), .B1(
        n20618), .B2(n20852), .ZN(n20570) );
  OAI211_X1 U23528 ( .C1(n20855), .C2(n20589), .A(n20571), .B(n20570), .ZN(
        P1_U3073) );
  AOI22_X1 U23529 ( .A1(n20940), .A2(n20585), .B1(n20939), .B2(n20584), .ZN(
        n20573) );
  AOI22_X1 U23530 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20586), .B1(
        n20618), .B2(n20941), .ZN(n20572) );
  OAI211_X1 U23531 ( .C1(n20944), .C2(n20589), .A(n20573), .B(n20572), .ZN(
        P1_U3074) );
  AOI22_X1 U23532 ( .A1(n20946), .A2(n20585), .B1(n20945), .B2(n20584), .ZN(
        n20575) );
  AOI22_X1 U23533 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20586), .B1(
        n20618), .B2(n20947), .ZN(n20574) );
  OAI211_X1 U23534 ( .C1(n20950), .C2(n20589), .A(n20575), .B(n20574), .ZN(
        P1_U3075) );
  AOI22_X1 U23535 ( .A1(n20952), .A2(n20585), .B1(n20951), .B2(n20584), .ZN(
        n20577) );
  AOI22_X1 U23536 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20586), .B1(
        n20618), .B2(n20860), .ZN(n20576) );
  OAI211_X1 U23537 ( .C1(n20863), .C2(n20589), .A(n20577), .B(n20576), .ZN(
        P1_U3076) );
  AOI22_X1 U23538 ( .A1(n20958), .A2(n20585), .B1(n20957), .B2(n20584), .ZN(
        n20579) );
  AOI22_X1 U23539 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20586), .B1(
        n20618), .B2(n20959), .ZN(n20578) );
  OAI211_X1 U23540 ( .C1(n20962), .C2(n20589), .A(n20579), .B(n20578), .ZN(
        P1_U3077) );
  AOI22_X1 U23541 ( .A1(n20964), .A2(n20585), .B1(n20963), .B2(n20584), .ZN(
        n20581) );
  AOI22_X1 U23542 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20586), .B1(
        n20618), .B2(n20965), .ZN(n20580) );
  OAI211_X1 U23543 ( .C1(n20970), .C2(n20589), .A(n20581), .B(n20580), .ZN(
        P1_U3078) );
  AOI22_X1 U23544 ( .A1(n20972), .A2(n20585), .B1(n20971), .B2(n20584), .ZN(
        n20583) );
  AOI22_X1 U23545 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20586), .B1(
        n20618), .B2(n20868), .ZN(n20582) );
  OAI211_X1 U23546 ( .C1(n20871), .C2(n20589), .A(n20583), .B(n20582), .ZN(
        P1_U3079) );
  AOI22_X1 U23547 ( .A1(n20980), .A2(n20585), .B1(n20978), .B2(n20584), .ZN(
        n20588) );
  AOI22_X1 U23548 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20586), .B1(
        n20618), .B2(n20874), .ZN(n20587) );
  OAI211_X1 U23549 ( .C1(n20879), .C2(n20589), .A(n20588), .B(n20587), .ZN(
        P1_U3080) );
  NAND3_X1 U23550 ( .A1(n20624), .A2(n20622), .A3(n20933), .ZN(n20591) );
  NAND2_X1 U23551 ( .A1(n20591), .A2(n20786), .ZN(n20597) );
  AND2_X1 U23552 ( .A1(n20592), .A2(n20881), .ZN(n20594) );
  INV_X1 U23553 ( .A(n20635), .ZN(n20630) );
  NOR2_X1 U23554 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20630), .ZN(
        n20599) );
  INV_X1 U23555 ( .A(n20599), .ZN(n20621) );
  OAI22_X1 U23556 ( .A1(n20624), .A2(n20938), .B1(n20621), .B2(n20792), .ZN(
        n20593) );
  INV_X1 U23557 ( .A(n20593), .ZN(n20601) );
  INV_X1 U23558 ( .A(n20594), .ZN(n20596) );
  AOI21_X1 U23559 ( .B1(n20597), .B2(n20596), .A(n20595), .ZN(n20598) );
  OAI211_X1 U23560 ( .C1(n20599), .C2(n20799), .A(n20888), .B(n20598), .ZN(
        n20625) );
  AOI22_X1 U23561 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20625), .B1(
        n20618), .B2(n20935), .ZN(n20600) );
  OAI211_X1 U23562 ( .C1(n20628), .C2(n20803), .A(n20601), .B(n20600), .ZN(
        P1_U3081) );
  OAI22_X1 U23563 ( .A1(n20624), .A2(n20895), .B1(n20621), .B2(n20804), .ZN(
        n20602) );
  INV_X1 U23564 ( .A(n20602), .ZN(n20604) );
  AOI22_X1 U23565 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20625), .B1(
        n20618), .B2(n20892), .ZN(n20603) );
  OAI211_X1 U23566 ( .C1(n20628), .C2(n20808), .A(n20604), .B(n20603), .ZN(
        P1_U3082) );
  OAI22_X1 U23567 ( .A1(n20624), .A2(n20899), .B1(n20621), .B2(n20809), .ZN(
        n20605) );
  INV_X1 U23568 ( .A(n20605), .ZN(n20607) );
  AOI22_X1 U23569 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20625), .B1(
        n20618), .B2(n20896), .ZN(n20606) );
  OAI211_X1 U23570 ( .C1(n20628), .C2(n20813), .A(n20607), .B(n20606), .ZN(
        P1_U3083) );
  OAI22_X1 U23571 ( .A1(n20624), .A2(n20956), .B1(n20621), .B2(n20814), .ZN(
        n20608) );
  INV_X1 U23572 ( .A(n20608), .ZN(n20610) );
  AOI22_X1 U23573 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20625), .B1(
        n20618), .B2(n20953), .ZN(n20609) );
  OAI211_X1 U23574 ( .C1(n20628), .C2(n20818), .A(n20610), .B(n20609), .ZN(
        P1_U3084) );
  OAI22_X1 U23575 ( .A1(n20624), .A2(n20905), .B1(n20621), .B2(n20819), .ZN(
        n20611) );
  INV_X1 U23576 ( .A(n20611), .ZN(n20613) );
  AOI22_X1 U23577 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20625), .B1(
        n20618), .B2(n20902), .ZN(n20612) );
  OAI211_X1 U23578 ( .C1(n20628), .C2(n20823), .A(n20613), .B(n20612), .ZN(
        P1_U3085) );
  OAI22_X1 U23579 ( .A1(n20624), .A2(n20909), .B1(n20621), .B2(n20824), .ZN(
        n20614) );
  INV_X1 U23580 ( .A(n20614), .ZN(n20616) );
  AOI22_X1 U23581 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20625), .B1(
        n20618), .B2(n20906), .ZN(n20615) );
  OAI211_X1 U23582 ( .C1(n20628), .C2(n20828), .A(n20616), .B(n20615), .ZN(
        P1_U3086) );
  OAI22_X1 U23583 ( .A1(n20624), .A2(n20976), .B1(n20621), .B2(n20829), .ZN(
        n20617) );
  INV_X1 U23584 ( .A(n20617), .ZN(n20620) );
  AOI22_X1 U23585 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20625), .B1(
        n20618), .B2(n20973), .ZN(n20619) );
  OAI211_X1 U23586 ( .C1(n20628), .C2(n20833), .A(n20620), .B(n20619), .ZN(
        P1_U3087) );
  OAI22_X1 U23587 ( .A1(n20622), .A2(n20879), .B1(n20835), .B2(n20621), .ZN(
        n20623) );
  INV_X1 U23588 ( .A(n20623), .ZN(n20627) );
  AOI22_X1 U23589 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20625), .B1(
        n20653), .B2(n20874), .ZN(n20626) );
  OAI211_X1 U23590 ( .C1(n20628), .C2(n20841), .A(n20627), .B(n20626), .ZN(
        P1_U3088) );
  INV_X1 U23591 ( .A(n20631), .ZN(n20652) );
  OAI222_X1 U23592 ( .A1(n20919), .A2(n20632), .B1(n20631), .B2(n20926), .C1(
        n20991), .C2(n20630), .ZN(n20651) );
  AOI22_X1 U23593 ( .A1(n20924), .A2(n20652), .B1(n20923), .B2(n20651), .ZN(
        n20638) );
  NOR3_X1 U23594 ( .A1(n20634), .A2(n20633), .A3(n20926), .ZN(n20636) );
  OAI21_X1 U23595 ( .B1(n20636), .B2(n20635), .A(n20932), .ZN(n20654) );
  AOI22_X1 U23596 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20654), .B1(
        n20653), .B2(n20935), .ZN(n20637) );
  OAI211_X1 U23597 ( .C1(n20938), .C2(n20664), .A(n20638), .B(n20637), .ZN(
        P1_U3089) );
  AOI22_X1 U23598 ( .A1(n20940), .A2(n20652), .B1(n20939), .B2(n20651), .ZN(
        n20640) );
  AOI22_X1 U23599 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20654), .B1(
        n20653), .B2(n20892), .ZN(n20639) );
  OAI211_X1 U23600 ( .C1(n20895), .C2(n20664), .A(n20640), .B(n20639), .ZN(
        P1_U3090) );
  AOI22_X1 U23601 ( .A1(n20946), .A2(n20652), .B1(n20945), .B2(n20651), .ZN(
        n20642) );
  AOI22_X1 U23602 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20654), .B1(
        n20653), .B2(n20896), .ZN(n20641) );
  OAI211_X1 U23603 ( .C1(n20899), .C2(n20664), .A(n20642), .B(n20641), .ZN(
        P1_U3091) );
  AOI22_X1 U23604 ( .A1(n20952), .A2(n20652), .B1(n20951), .B2(n20651), .ZN(
        n20644) );
  AOI22_X1 U23605 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20654), .B1(
        n20653), .B2(n20953), .ZN(n20643) );
  OAI211_X1 U23606 ( .C1(n20956), .C2(n20664), .A(n20644), .B(n20643), .ZN(
        P1_U3092) );
  AOI22_X1 U23607 ( .A1(n20958), .A2(n20652), .B1(n20957), .B2(n20651), .ZN(
        n20646) );
  AOI22_X1 U23608 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20654), .B1(
        n20653), .B2(n20902), .ZN(n20645) );
  OAI211_X1 U23609 ( .C1(n20905), .C2(n20664), .A(n20646), .B(n20645), .ZN(
        P1_U3093) );
  AOI22_X1 U23610 ( .A1(n20964), .A2(n20652), .B1(n20963), .B2(n20651), .ZN(
        n20648) );
  AOI22_X1 U23611 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20654), .B1(
        n20653), .B2(n20906), .ZN(n20647) );
  OAI211_X1 U23612 ( .C1(n20909), .C2(n20664), .A(n20648), .B(n20647), .ZN(
        P1_U3094) );
  AOI22_X1 U23613 ( .A1(n20972), .A2(n20652), .B1(n20971), .B2(n20651), .ZN(
        n20650) );
  AOI22_X1 U23614 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20654), .B1(
        n20653), .B2(n20973), .ZN(n20649) );
  OAI211_X1 U23615 ( .C1(n20976), .C2(n20664), .A(n20650), .B(n20649), .ZN(
        P1_U3095) );
  AOI22_X1 U23616 ( .A1(n20980), .A2(n20652), .B1(n20978), .B2(n20651), .ZN(
        n20656) );
  AOI22_X1 U23617 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20654), .B1(
        n20653), .B2(n20981), .ZN(n20655) );
  OAI211_X1 U23618 ( .C1(n20987), .C2(n20664), .A(n20656), .B(n20655), .ZN(
        P1_U3096) );
  INV_X1 U23619 ( .A(n20763), .ZN(n20658) );
  NAND3_X1 U23620 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12753), .A3(
        n20791), .ZN(n20689) );
  NOR2_X1 U23621 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20689), .ZN(
        n20684) );
  AND2_X1 U23622 ( .A1(n20659), .A2(n13909), .ZN(n20751) );
  AOI21_X1 U23623 ( .B1(n20751), .B2(n20660), .A(n20684), .ZN(n20666) );
  INV_X1 U23624 ( .A(n20719), .ZN(n20662) );
  NOR2_X1 U23625 ( .A1(n20662), .A2(n20661), .ZN(n20789) );
  INV_X1 U23626 ( .A(n20789), .ZN(n20795) );
  OAI22_X1 U23627 ( .A1(n20666), .A2(n20926), .B1(n20663), .B2(n20795), .ZN(
        n20683) );
  AOI22_X1 U23628 ( .A1(n20924), .A2(n20684), .B1(n20923), .B2(n20683), .ZN(
        n20670) );
  INV_X1 U23629 ( .A(n20712), .ZN(n20665) );
  OAI21_X1 U23630 ( .B1(n20665), .B2(n20685), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20667) );
  NAND2_X1 U23631 ( .A1(n20667), .A2(n20666), .ZN(n20668) );
  AOI22_X1 U23632 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20686), .B1(
        n20685), .B2(n20935), .ZN(n20669) );
  OAI211_X1 U23633 ( .C1(n20938), .C2(n20712), .A(n20670), .B(n20669), .ZN(
        P1_U3097) );
  AOI22_X1 U23634 ( .A1(n20940), .A2(n20684), .B1(n20939), .B2(n20683), .ZN(
        n20672) );
  AOI22_X1 U23635 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20686), .B1(
        n20685), .B2(n20892), .ZN(n20671) );
  OAI211_X1 U23636 ( .C1(n20895), .C2(n20712), .A(n20672), .B(n20671), .ZN(
        P1_U3098) );
  AOI22_X1 U23637 ( .A1(n20946), .A2(n20684), .B1(n20945), .B2(n20683), .ZN(
        n20674) );
  AOI22_X1 U23638 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20686), .B1(
        n20685), .B2(n20896), .ZN(n20673) );
  OAI211_X1 U23639 ( .C1(n20899), .C2(n20712), .A(n20674), .B(n20673), .ZN(
        P1_U3099) );
  AOI22_X1 U23640 ( .A1(n20952), .A2(n20684), .B1(n20951), .B2(n20683), .ZN(
        n20676) );
  AOI22_X1 U23641 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20686), .B1(
        n20685), .B2(n20953), .ZN(n20675) );
  OAI211_X1 U23642 ( .C1(n20956), .C2(n20712), .A(n20676), .B(n20675), .ZN(
        P1_U3100) );
  AOI22_X1 U23643 ( .A1(n20958), .A2(n20684), .B1(n20957), .B2(n20683), .ZN(
        n20678) );
  AOI22_X1 U23644 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20686), .B1(
        n20685), .B2(n20902), .ZN(n20677) );
  OAI211_X1 U23645 ( .C1(n20905), .C2(n20712), .A(n20678), .B(n20677), .ZN(
        P1_U3101) );
  AOI22_X1 U23646 ( .A1(n20964), .A2(n20684), .B1(n20963), .B2(n20683), .ZN(
        n20680) );
  AOI22_X1 U23647 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20686), .B1(
        n20685), .B2(n20906), .ZN(n20679) );
  OAI211_X1 U23648 ( .C1(n20909), .C2(n20712), .A(n20680), .B(n20679), .ZN(
        P1_U3102) );
  AOI22_X1 U23649 ( .A1(n20972), .A2(n20684), .B1(n20971), .B2(n20683), .ZN(
        n20682) );
  AOI22_X1 U23650 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20686), .B1(
        n20685), .B2(n20973), .ZN(n20681) );
  OAI211_X1 U23651 ( .C1(n20976), .C2(n20712), .A(n20682), .B(n20681), .ZN(
        P1_U3103) );
  AOI22_X1 U23652 ( .A1(n20980), .A2(n20684), .B1(n20978), .B2(n20683), .ZN(
        n20688) );
  AOI22_X1 U23653 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20686), .B1(
        n20685), .B2(n20981), .ZN(n20687) );
  OAI211_X1 U23654 ( .C1(n20987), .C2(n20712), .A(n20688), .B(n20687), .ZN(
        P1_U3104) );
  NOR2_X1 U23655 ( .A1(n20843), .A2(n20689), .ZN(n20708) );
  AOI21_X1 U23656 ( .B1(n20751), .B2(n20845), .A(n20708), .ZN(n20690) );
  OAI22_X1 U23657 ( .A1(n20690), .A2(n20926), .B1(n20689), .B2(n20991), .ZN(
        n20707) );
  AOI22_X1 U23658 ( .A1(n20924), .A2(n20708), .B1(n20923), .B2(n20707), .ZN(
        n20694) );
  INV_X1 U23659 ( .A(n20689), .ZN(n20692) );
  OAI211_X1 U23660 ( .C1(n20763), .C2(n20848), .A(n20933), .B(n20690), .ZN(
        n20691) );
  OAI211_X1 U23661 ( .C1(n20933), .C2(n20692), .A(n20932), .B(n20691), .ZN(
        n20709) );
  AOI22_X1 U23662 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20709), .B1(
        n20746), .B2(n20852), .ZN(n20693) );
  OAI211_X1 U23663 ( .C1(n20855), .C2(n20712), .A(n20694), .B(n20693), .ZN(
        P1_U3105) );
  AOI22_X1 U23664 ( .A1(n20940), .A2(n20708), .B1(n20939), .B2(n20707), .ZN(
        n20696) );
  AOI22_X1 U23665 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20709), .B1(
        n20746), .B2(n20941), .ZN(n20695) );
  OAI211_X1 U23666 ( .C1(n20944), .C2(n20712), .A(n20696), .B(n20695), .ZN(
        P1_U3106) );
  AOI22_X1 U23667 ( .A1(n20946), .A2(n20708), .B1(n20945), .B2(n20707), .ZN(
        n20698) );
  AOI22_X1 U23668 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20709), .B1(
        n20746), .B2(n20947), .ZN(n20697) );
  OAI211_X1 U23669 ( .C1(n20950), .C2(n20712), .A(n20698), .B(n20697), .ZN(
        P1_U3107) );
  AOI22_X1 U23670 ( .A1(n20952), .A2(n20708), .B1(n20951), .B2(n20707), .ZN(
        n20700) );
  AOI22_X1 U23671 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20709), .B1(
        n20746), .B2(n20860), .ZN(n20699) );
  OAI211_X1 U23672 ( .C1(n20863), .C2(n20712), .A(n20700), .B(n20699), .ZN(
        P1_U3108) );
  AOI22_X1 U23673 ( .A1(n20958), .A2(n20708), .B1(n20957), .B2(n20707), .ZN(
        n20702) );
  AOI22_X1 U23674 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20709), .B1(
        n20746), .B2(n20959), .ZN(n20701) );
  OAI211_X1 U23675 ( .C1(n20962), .C2(n20712), .A(n20702), .B(n20701), .ZN(
        P1_U3109) );
  AOI22_X1 U23676 ( .A1(n20964), .A2(n20708), .B1(n20963), .B2(n20707), .ZN(
        n20704) );
  AOI22_X1 U23677 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20709), .B1(
        n20746), .B2(n20965), .ZN(n20703) );
  OAI211_X1 U23678 ( .C1(n20970), .C2(n20712), .A(n20704), .B(n20703), .ZN(
        P1_U3110) );
  AOI22_X1 U23679 ( .A1(n20972), .A2(n20708), .B1(n20971), .B2(n20707), .ZN(
        n20706) );
  AOI22_X1 U23680 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20709), .B1(
        n20746), .B2(n20868), .ZN(n20705) );
  OAI211_X1 U23681 ( .C1(n20871), .C2(n20712), .A(n20706), .B(n20705), .ZN(
        P1_U3111) );
  AOI22_X1 U23682 ( .A1(n20980), .A2(n20708), .B1(n20978), .B2(n20707), .ZN(
        n20711) );
  AOI22_X1 U23683 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20709), .B1(
        n20746), .B2(n20874), .ZN(n20710) );
  OAI211_X1 U23684 ( .C1(n20879), .C2(n20712), .A(n20711), .B(n20710), .ZN(
        P1_U3112) );
  NAND3_X1 U23685 ( .A1(n20783), .A2(n20739), .A3(n20933), .ZN(n20713) );
  NAND2_X1 U23686 ( .A1(n20713), .A2(n20786), .ZN(n20718) );
  AND2_X1 U23687 ( .A1(n20751), .A2(n20881), .ZN(n20716) );
  NOR2_X1 U23688 ( .A1(n20719), .A2(n12729), .ZN(n20882) );
  NAND3_X1 U23689 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n12753), .ZN(n20758) );
  OR2_X1 U23690 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20758), .ZN(
        n20744) );
  OAI22_X1 U23691 ( .A1(n20739), .A2(n20855), .B1(n20792), .B2(n20744), .ZN(
        n20715) );
  INV_X1 U23692 ( .A(n20715), .ZN(n20723) );
  INV_X1 U23693 ( .A(n20716), .ZN(n20717) );
  AOI22_X1 U23694 ( .A1(n20718), .A2(n20717), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20744), .ZN(n20720) );
  OAI21_X1 U23695 ( .B1(n12729), .B2(n20719), .A(P1_STATE2_REG_2__SCAN_IN), 
        .ZN(n20887) );
  NAND3_X1 U23696 ( .A1(n20721), .A2(n20720), .A3(n20887), .ZN(n20747) );
  AOI22_X1 U23697 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20747), .B1(
        n20741), .B2(n20852), .ZN(n20722) );
  OAI211_X1 U23698 ( .C1(n20750), .C2(n20803), .A(n20723), .B(n20722), .ZN(
        P1_U3113) );
  OAI22_X1 U23699 ( .A1(n20739), .A2(n20944), .B1(n20804), .B2(n20744), .ZN(
        n20724) );
  INV_X1 U23700 ( .A(n20724), .ZN(n20726) );
  AOI22_X1 U23701 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20747), .B1(
        n20741), .B2(n20941), .ZN(n20725) );
  OAI211_X1 U23702 ( .C1(n20750), .C2(n20808), .A(n20726), .B(n20725), .ZN(
        P1_U3114) );
  OAI22_X1 U23703 ( .A1(n20739), .A2(n20950), .B1(n20809), .B2(n20744), .ZN(
        n20727) );
  INV_X1 U23704 ( .A(n20727), .ZN(n20729) );
  AOI22_X1 U23705 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20747), .B1(
        n20741), .B2(n20947), .ZN(n20728) );
  OAI211_X1 U23706 ( .C1(n20750), .C2(n20813), .A(n20729), .B(n20728), .ZN(
        P1_U3115) );
  OAI22_X1 U23707 ( .A1(n20739), .A2(n20863), .B1(n20814), .B2(n20744), .ZN(
        n20730) );
  INV_X1 U23708 ( .A(n20730), .ZN(n20732) );
  AOI22_X1 U23709 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20747), .B1(
        n20741), .B2(n20860), .ZN(n20731) );
  OAI211_X1 U23710 ( .C1(n20750), .C2(n20818), .A(n20732), .B(n20731), .ZN(
        P1_U3116) );
  OAI22_X1 U23711 ( .A1(n20739), .A2(n20962), .B1(n20819), .B2(n20744), .ZN(
        n20733) );
  INV_X1 U23712 ( .A(n20733), .ZN(n20735) );
  AOI22_X1 U23713 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20747), .B1(
        n20741), .B2(n20959), .ZN(n20734) );
  OAI211_X1 U23714 ( .C1(n20750), .C2(n20823), .A(n20735), .B(n20734), .ZN(
        P1_U3117) );
  OAI22_X1 U23715 ( .A1(n20783), .A2(n20909), .B1(n20824), .B2(n20744), .ZN(
        n20736) );
  INV_X1 U23716 ( .A(n20736), .ZN(n20738) );
  AOI22_X1 U23717 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20747), .B1(
        n20746), .B2(n20906), .ZN(n20737) );
  OAI211_X1 U23718 ( .C1(n20750), .C2(n20828), .A(n20738), .B(n20737), .ZN(
        P1_U3118) );
  OAI22_X1 U23719 ( .A1(n20739), .A2(n20871), .B1(n20829), .B2(n20744), .ZN(
        n20740) );
  INV_X1 U23720 ( .A(n20740), .ZN(n20743) );
  AOI22_X1 U23721 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20747), .B1(
        n20741), .B2(n20868), .ZN(n20742) );
  OAI211_X1 U23722 ( .C1(n20750), .C2(n20833), .A(n20743), .B(n20742), .ZN(
        P1_U3119) );
  OAI22_X1 U23723 ( .A1(n20783), .A2(n20987), .B1(n20835), .B2(n20744), .ZN(
        n20745) );
  INV_X1 U23724 ( .A(n20745), .ZN(n20749) );
  AOI22_X1 U23725 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20747), .B1(
        n20746), .B2(n20981), .ZN(n20748) );
  OAI211_X1 U23726 ( .C1(n20750), .C2(n20841), .A(n20749), .B(n20748), .ZN(
        P1_U3120) );
  INV_X1 U23727 ( .A(n20751), .ZN(n20754) );
  INV_X1 U23728 ( .A(n20752), .ZN(n20753) );
  NAND2_X1 U23729 ( .A1(n20753), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20756) );
  OAI21_X1 U23730 ( .B1(n20754), .B2(n20919), .A(n20756), .ZN(n20760) );
  INV_X1 U23731 ( .A(n20760), .ZN(n20755) );
  OAI22_X1 U23732 ( .A1(n20755), .A2(n20926), .B1(n20758), .B2(n20991), .ZN(
        n20779) );
  INV_X1 U23733 ( .A(n20756), .ZN(n20778) );
  AOI22_X1 U23734 ( .A1(n20779), .A2(n20923), .B1(n20924), .B2(n20778), .ZN(
        n20765) );
  AOI21_X1 U23735 ( .B1(n20763), .B2(n20933), .A(n20929), .ZN(n20761) );
  AOI21_X1 U23736 ( .B1(n20926), .B2(n20758), .A(n20757), .ZN(n20759) );
  AOI22_X1 U23737 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20780), .B1(
        n20837), .B2(n20852), .ZN(n20764) );
  OAI211_X1 U23738 ( .C1(n20855), .C2(n20783), .A(n20765), .B(n20764), .ZN(
        P1_U3121) );
  AOI22_X1 U23739 ( .A1(n20779), .A2(n20939), .B1(n20940), .B2(n20778), .ZN(
        n20767) );
  AOI22_X1 U23740 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20780), .B1(
        n20837), .B2(n20941), .ZN(n20766) );
  OAI211_X1 U23741 ( .C1(n20944), .C2(n20783), .A(n20767), .B(n20766), .ZN(
        P1_U3122) );
  AOI22_X1 U23742 ( .A1(n20779), .A2(n20945), .B1(n20946), .B2(n20778), .ZN(
        n20769) );
  AOI22_X1 U23743 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20780), .B1(
        n20837), .B2(n20947), .ZN(n20768) );
  OAI211_X1 U23744 ( .C1(n20950), .C2(n20783), .A(n20769), .B(n20768), .ZN(
        P1_U3123) );
  AOI22_X1 U23745 ( .A1(n20779), .A2(n20951), .B1(n20952), .B2(n20778), .ZN(
        n20771) );
  AOI22_X1 U23746 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20780), .B1(
        n20837), .B2(n20860), .ZN(n20770) );
  OAI211_X1 U23747 ( .C1(n20863), .C2(n20783), .A(n20771), .B(n20770), .ZN(
        P1_U3124) );
  AOI22_X1 U23748 ( .A1(n20779), .A2(n20957), .B1(n20958), .B2(n20778), .ZN(
        n20773) );
  AOI22_X1 U23749 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20780), .B1(
        n20837), .B2(n20959), .ZN(n20772) );
  OAI211_X1 U23750 ( .C1(n20962), .C2(n20783), .A(n20773), .B(n20772), .ZN(
        P1_U3125) );
  AOI22_X1 U23751 ( .A1(n20779), .A2(n20963), .B1(n20964), .B2(n20778), .ZN(
        n20775) );
  AOI22_X1 U23752 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20780), .B1(
        n20837), .B2(n20965), .ZN(n20774) );
  OAI211_X1 U23753 ( .C1(n20970), .C2(n20783), .A(n20775), .B(n20774), .ZN(
        P1_U3126) );
  AOI22_X1 U23754 ( .A1(n20779), .A2(n20971), .B1(n20972), .B2(n20778), .ZN(
        n20777) );
  AOI22_X1 U23755 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20780), .B1(
        n20837), .B2(n20868), .ZN(n20776) );
  OAI211_X1 U23756 ( .C1(n20871), .C2(n20783), .A(n20777), .B(n20776), .ZN(
        P1_U3127) );
  AOI22_X1 U23757 ( .A1(n20779), .A2(n20978), .B1(n20980), .B2(n20778), .ZN(
        n20782) );
  AOI22_X1 U23758 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20780), .B1(
        n20837), .B2(n20874), .ZN(n20781) );
  OAI211_X1 U23759 ( .C1(n20879), .C2(n20783), .A(n20782), .B(n20781), .ZN(
        P1_U3128) );
  NAND3_X1 U23760 ( .A1(n20785), .A2(n20933), .A3(n20878), .ZN(n20787) );
  NAND2_X1 U23761 ( .A1(n20787), .A2(n20786), .ZN(n20797) );
  OR2_X1 U23762 ( .A1(n13909), .A2(n20788), .ZN(n20844) );
  NOR2_X1 U23763 ( .A1(n20844), .A2(n20881), .ZN(n20794) );
  NAND3_X1 U23764 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20791), .ZN(n20846) );
  NOR2_X1 U23765 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20846), .ZN(
        n20800) );
  INV_X1 U23766 ( .A(n20800), .ZN(n20834) );
  OAI22_X1 U23767 ( .A1(n20878), .A2(n20938), .B1(n20792), .B2(n20834), .ZN(
        n20793) );
  INV_X1 U23768 ( .A(n20793), .ZN(n20802) );
  INV_X1 U23769 ( .A(n20794), .ZN(n20796) );
  AOI22_X1 U23770 ( .A1(n20797), .A2(n20796), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20795), .ZN(n20798) );
  OAI211_X1 U23771 ( .C1(n20800), .C2(n20799), .A(n20888), .B(n20798), .ZN(
        n20838) );
  AOI22_X1 U23772 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20838), .B1(
        n20837), .B2(n20935), .ZN(n20801) );
  OAI211_X1 U23773 ( .C1(n20842), .C2(n20803), .A(n20802), .B(n20801), .ZN(
        P1_U3129) );
  OAI22_X1 U23774 ( .A1(n20878), .A2(n20895), .B1(n20834), .B2(n20804), .ZN(
        n20805) );
  INV_X1 U23775 ( .A(n20805), .ZN(n20807) );
  AOI22_X1 U23776 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20838), .B1(
        n20837), .B2(n20892), .ZN(n20806) );
  OAI211_X1 U23777 ( .C1(n20842), .C2(n20808), .A(n20807), .B(n20806), .ZN(
        P1_U3130) );
  OAI22_X1 U23778 ( .A1(n20878), .A2(n20899), .B1(n20834), .B2(n20809), .ZN(
        n20810) );
  INV_X1 U23779 ( .A(n20810), .ZN(n20812) );
  AOI22_X1 U23780 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20838), .B1(
        n20837), .B2(n20896), .ZN(n20811) );
  OAI211_X1 U23781 ( .C1(n20842), .C2(n20813), .A(n20812), .B(n20811), .ZN(
        P1_U3131) );
  OAI22_X1 U23782 ( .A1(n20878), .A2(n20956), .B1(n20834), .B2(n20814), .ZN(
        n20815) );
  INV_X1 U23783 ( .A(n20815), .ZN(n20817) );
  AOI22_X1 U23784 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20838), .B1(
        n20837), .B2(n20953), .ZN(n20816) );
  OAI211_X1 U23785 ( .C1(n20842), .C2(n20818), .A(n20817), .B(n20816), .ZN(
        P1_U3132) );
  OAI22_X1 U23786 ( .A1(n20878), .A2(n20905), .B1(n20834), .B2(n20819), .ZN(
        n20820) );
  INV_X1 U23787 ( .A(n20820), .ZN(n20822) );
  AOI22_X1 U23788 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20838), .B1(
        n20837), .B2(n20902), .ZN(n20821) );
  OAI211_X1 U23789 ( .C1(n20842), .C2(n20823), .A(n20822), .B(n20821), .ZN(
        P1_U3133) );
  OAI22_X1 U23790 ( .A1(n20878), .A2(n20909), .B1(n20834), .B2(n20824), .ZN(
        n20825) );
  INV_X1 U23791 ( .A(n20825), .ZN(n20827) );
  AOI22_X1 U23792 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20838), .B1(
        n20837), .B2(n20906), .ZN(n20826) );
  OAI211_X1 U23793 ( .C1(n20842), .C2(n20828), .A(n20827), .B(n20826), .ZN(
        P1_U3134) );
  OAI22_X1 U23794 ( .A1(n20878), .A2(n20976), .B1(n20834), .B2(n20829), .ZN(
        n20830) );
  INV_X1 U23795 ( .A(n20830), .ZN(n20832) );
  AOI22_X1 U23796 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20838), .B1(
        n20837), .B2(n20973), .ZN(n20831) );
  OAI211_X1 U23797 ( .C1(n20842), .C2(n20833), .A(n20832), .B(n20831), .ZN(
        P1_U3135) );
  OAI22_X1 U23798 ( .A1(n20878), .A2(n20987), .B1(n20835), .B2(n20834), .ZN(
        n20836) );
  INV_X1 U23799 ( .A(n20836), .ZN(n20840) );
  AOI22_X1 U23800 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20838), .B1(
        n20837), .B2(n20981), .ZN(n20839) );
  OAI211_X1 U23801 ( .C1(n20842), .C2(n20841), .A(n20840), .B(n20839), .ZN(
        P1_U3136) );
  NOR2_X1 U23802 ( .A1(n20843), .A2(n20846), .ZN(n20873) );
  INV_X1 U23803 ( .A(n20844), .ZN(n20921) );
  AOI21_X1 U23804 ( .B1(n20921), .B2(n20845), .A(n20873), .ZN(n20847) );
  OAI22_X1 U23805 ( .A1(n20847), .A2(n20926), .B1(n20846), .B2(n20991), .ZN(
        n20872) );
  AOI22_X1 U23806 ( .A1(n20924), .A2(n20873), .B1(n20923), .B2(n20872), .ZN(
        n20854) );
  INV_X1 U23807 ( .A(n20846), .ZN(n20850) );
  OAI211_X1 U23808 ( .C1(n20925), .C2(n20848), .A(n20933), .B(n20847), .ZN(
        n20849) );
  OAI211_X1 U23809 ( .C1(n20933), .C2(n20850), .A(n20932), .B(n20849), .ZN(
        n20875) );
  AOI22_X1 U23810 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20875), .B1(
        n20914), .B2(n20852), .ZN(n20853) );
  OAI211_X1 U23811 ( .C1(n20855), .C2(n20878), .A(n20854), .B(n20853), .ZN(
        P1_U3137) );
  AOI22_X1 U23812 ( .A1(n20940), .A2(n20873), .B1(n20939), .B2(n20872), .ZN(
        n20857) );
  AOI22_X1 U23813 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20875), .B1(
        n20914), .B2(n20941), .ZN(n20856) );
  OAI211_X1 U23814 ( .C1(n20944), .C2(n20878), .A(n20857), .B(n20856), .ZN(
        P1_U3138) );
  AOI22_X1 U23815 ( .A1(n20946), .A2(n20873), .B1(n20945), .B2(n20872), .ZN(
        n20859) );
  AOI22_X1 U23816 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20875), .B1(
        n20914), .B2(n20947), .ZN(n20858) );
  OAI211_X1 U23817 ( .C1(n20950), .C2(n20878), .A(n20859), .B(n20858), .ZN(
        P1_U3139) );
  AOI22_X1 U23818 ( .A1(n20952), .A2(n20873), .B1(n20951), .B2(n20872), .ZN(
        n20862) );
  AOI22_X1 U23819 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20875), .B1(
        n20914), .B2(n20860), .ZN(n20861) );
  OAI211_X1 U23820 ( .C1(n20863), .C2(n20878), .A(n20862), .B(n20861), .ZN(
        P1_U3140) );
  AOI22_X1 U23821 ( .A1(n20958), .A2(n20873), .B1(n20957), .B2(n20872), .ZN(
        n20865) );
  AOI22_X1 U23822 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20875), .B1(
        n20914), .B2(n20959), .ZN(n20864) );
  OAI211_X1 U23823 ( .C1(n20962), .C2(n20878), .A(n20865), .B(n20864), .ZN(
        P1_U3141) );
  AOI22_X1 U23824 ( .A1(n20964), .A2(n20873), .B1(n20963), .B2(n20872), .ZN(
        n20867) );
  AOI22_X1 U23825 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20875), .B1(
        n20914), .B2(n20965), .ZN(n20866) );
  OAI211_X1 U23826 ( .C1(n20970), .C2(n20878), .A(n20867), .B(n20866), .ZN(
        P1_U3142) );
  AOI22_X1 U23827 ( .A1(n20972), .A2(n20873), .B1(n20971), .B2(n20872), .ZN(
        n20870) );
  AOI22_X1 U23828 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20875), .B1(
        n20914), .B2(n20868), .ZN(n20869) );
  OAI211_X1 U23829 ( .C1(n20871), .C2(n20878), .A(n20870), .B(n20869), .ZN(
        P1_U3143) );
  AOI22_X1 U23830 ( .A1(n20980), .A2(n20873), .B1(n20978), .B2(n20872), .ZN(
        n20877) );
  AOI22_X1 U23831 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20875), .B1(
        n20914), .B2(n20874), .ZN(n20876) );
  OAI211_X1 U23832 ( .C1(n20879), .C2(n20878), .A(n20877), .B(n20876), .ZN(
        P1_U3144) );
  NOR2_X1 U23833 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20922), .ZN(
        n20913) );
  NAND2_X1 U23834 ( .A1(n20921), .A2(n20881), .ZN(n20885) );
  INV_X1 U23835 ( .A(n20882), .ZN(n20884) );
  OAI22_X1 U23836 ( .A1(n20885), .A2(n20926), .B1(n20884), .B2(n20883), .ZN(
        n20912) );
  AOI22_X1 U23837 ( .A1(n20924), .A2(n20913), .B1(n20923), .B2(n20912), .ZN(
        n20891) );
  OAI21_X1 U23838 ( .B1(n20982), .B2(n20914), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20886) );
  AOI21_X1 U23839 ( .B1(n20886), .B2(n20885), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20889) );
  AOI22_X1 U23840 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20915), .B1(
        n20914), .B2(n20935), .ZN(n20890) );
  OAI211_X1 U23841 ( .C1(n20938), .C2(n20969), .A(n20891), .B(n20890), .ZN(
        P1_U3145) );
  AOI22_X1 U23842 ( .A1(n20940), .A2(n20913), .B1(n20939), .B2(n20912), .ZN(
        n20894) );
  AOI22_X1 U23843 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20915), .B1(
        n20914), .B2(n20892), .ZN(n20893) );
  OAI211_X1 U23844 ( .C1(n20895), .C2(n20969), .A(n20894), .B(n20893), .ZN(
        P1_U3146) );
  AOI22_X1 U23845 ( .A1(n20946), .A2(n20913), .B1(n20945), .B2(n20912), .ZN(
        n20898) );
  AOI22_X1 U23846 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20915), .B1(
        n20914), .B2(n20896), .ZN(n20897) );
  OAI211_X1 U23847 ( .C1(n20899), .C2(n20969), .A(n20898), .B(n20897), .ZN(
        P1_U3147) );
  AOI22_X1 U23848 ( .A1(n20952), .A2(n20913), .B1(n20951), .B2(n20912), .ZN(
        n20901) );
  AOI22_X1 U23849 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20915), .B1(
        n20914), .B2(n20953), .ZN(n20900) );
  OAI211_X1 U23850 ( .C1(n20956), .C2(n20969), .A(n20901), .B(n20900), .ZN(
        P1_U3148) );
  AOI22_X1 U23851 ( .A1(n20958), .A2(n20913), .B1(n20957), .B2(n20912), .ZN(
        n20904) );
  AOI22_X1 U23852 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20915), .B1(
        n20914), .B2(n20902), .ZN(n20903) );
  OAI211_X1 U23853 ( .C1(n20905), .C2(n20969), .A(n20904), .B(n20903), .ZN(
        P1_U3149) );
  AOI22_X1 U23854 ( .A1(n20964), .A2(n20913), .B1(n20963), .B2(n20912), .ZN(
        n20908) );
  AOI22_X1 U23855 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20915), .B1(
        n20914), .B2(n20906), .ZN(n20907) );
  OAI211_X1 U23856 ( .C1(n20909), .C2(n20969), .A(n20908), .B(n20907), .ZN(
        P1_U3150) );
  AOI22_X1 U23857 ( .A1(n20972), .A2(n20913), .B1(n20971), .B2(n20912), .ZN(
        n20911) );
  AOI22_X1 U23858 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20915), .B1(
        n20914), .B2(n20973), .ZN(n20910) );
  OAI211_X1 U23859 ( .C1(n20976), .C2(n20969), .A(n20911), .B(n20910), .ZN(
        P1_U3151) );
  AOI22_X1 U23860 ( .A1(n20980), .A2(n20913), .B1(n20978), .B2(n20912), .ZN(
        n20917) );
  AOI22_X1 U23861 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20915), .B1(
        n20914), .B2(n20981), .ZN(n20916) );
  OAI211_X1 U23862 ( .C1(n20987), .C2(n20969), .A(n20917), .B(n20916), .ZN(
        P1_U3152) );
  INV_X1 U23863 ( .A(n20918), .ZN(n20979) );
  INV_X1 U23864 ( .A(n20919), .ZN(n20920) );
  AOI21_X1 U23865 ( .B1(n20921), .B2(n20920), .A(n20979), .ZN(n20928) );
  OAI22_X1 U23866 ( .A1(n20928), .A2(n20926), .B1(n20922), .B2(n20991), .ZN(
        n20977) );
  AOI22_X1 U23867 ( .A1(n20924), .A2(n20979), .B1(n20923), .B2(n20977), .ZN(
        n20937) );
  INV_X1 U23868 ( .A(n20925), .ZN(n20927) );
  NOR2_X1 U23869 ( .A1(n20927), .A2(n20926), .ZN(n20930) );
  OAI21_X1 U23870 ( .B1(n20930), .B2(n20929), .A(n20928), .ZN(n20931) );
  OAI211_X1 U23871 ( .C1(n20934), .C2(n20933), .A(n20932), .B(n20931), .ZN(
        n20983) );
  AOI22_X1 U23872 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20983), .B1(
        n20982), .B2(n20935), .ZN(n20936) );
  OAI211_X1 U23873 ( .C1(n20938), .C2(n20986), .A(n20937), .B(n20936), .ZN(
        P1_U3153) );
  AOI22_X1 U23874 ( .A1(n20940), .A2(n20979), .B1(n20939), .B2(n20977), .ZN(
        n20943) );
  AOI22_X1 U23875 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20983), .B1(
        n20966), .B2(n20941), .ZN(n20942) );
  OAI211_X1 U23876 ( .C1(n20944), .C2(n20969), .A(n20943), .B(n20942), .ZN(
        P1_U3154) );
  AOI22_X1 U23877 ( .A1(n20946), .A2(n20979), .B1(n20945), .B2(n20977), .ZN(
        n20949) );
  AOI22_X1 U23878 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20983), .B1(
        n20966), .B2(n20947), .ZN(n20948) );
  OAI211_X1 U23879 ( .C1(n20950), .C2(n20969), .A(n20949), .B(n20948), .ZN(
        P1_U3155) );
  AOI22_X1 U23880 ( .A1(n20952), .A2(n20979), .B1(n20951), .B2(n20977), .ZN(
        n20955) );
  AOI22_X1 U23881 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20983), .B1(
        n20982), .B2(n20953), .ZN(n20954) );
  OAI211_X1 U23882 ( .C1(n20956), .C2(n20986), .A(n20955), .B(n20954), .ZN(
        P1_U3156) );
  AOI22_X1 U23883 ( .A1(n20958), .A2(n20979), .B1(n20957), .B2(n20977), .ZN(
        n20961) );
  AOI22_X1 U23884 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20983), .B1(
        n20966), .B2(n20959), .ZN(n20960) );
  OAI211_X1 U23885 ( .C1(n20962), .C2(n20969), .A(n20961), .B(n20960), .ZN(
        P1_U3157) );
  AOI22_X1 U23886 ( .A1(n20964), .A2(n20979), .B1(n20963), .B2(n20977), .ZN(
        n20968) );
  AOI22_X1 U23887 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20983), .B1(
        n20966), .B2(n20965), .ZN(n20967) );
  OAI211_X1 U23888 ( .C1(n20970), .C2(n20969), .A(n20968), .B(n20967), .ZN(
        P1_U3158) );
  AOI22_X1 U23889 ( .A1(n20972), .A2(n20979), .B1(n20971), .B2(n20977), .ZN(
        n20975) );
  AOI22_X1 U23890 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20983), .B1(
        n20982), .B2(n20973), .ZN(n20974) );
  OAI211_X1 U23891 ( .C1(n20976), .C2(n20986), .A(n20975), .B(n20974), .ZN(
        P1_U3159) );
  AOI22_X1 U23892 ( .A1(n20980), .A2(n20979), .B1(n20978), .B2(n20977), .ZN(
        n20985) );
  AOI22_X1 U23893 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20983), .B1(
        n20982), .B2(n20981), .ZN(n20984) );
  OAI211_X1 U23894 ( .C1(n20987), .C2(n20986), .A(n20985), .B(n20984), .ZN(
        P1_U3160) );
  INV_X1 U23895 ( .A(n20988), .ZN(n20992) );
  AOI22_X1 U23896 ( .A1(n20992), .A2(n20991), .B1(n20990), .B2(n20989), .ZN(
        P1_U3163) );
  AND2_X1 U23897 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n21054), .ZN(
        P1_U3164) );
  AND2_X1 U23898 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n21054), .ZN(
        P1_U3165) );
  AND2_X1 U23899 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20993), .ZN(
        P1_U3166) );
  AND2_X1 U23900 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20993), .ZN(
        P1_U3167) );
  AND2_X1 U23901 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20993), .ZN(
        P1_U3168) );
  AND2_X1 U23902 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20993), .ZN(
        P1_U3169) );
  AND2_X1 U23903 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20993), .ZN(
        P1_U3170) );
  AND2_X1 U23904 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20993), .ZN(
        P1_U3171) );
  AND2_X1 U23905 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20993), .ZN(
        P1_U3172) );
  AND2_X1 U23906 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20993), .ZN(
        P1_U3173) );
  AND2_X1 U23907 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20993), .ZN(
        P1_U3174) );
  AND2_X1 U23908 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20993), .ZN(
        P1_U3175) );
  AND2_X1 U23909 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20993), .ZN(
        P1_U3176) );
  AND2_X1 U23910 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20993), .ZN(
        P1_U3177) );
  AND2_X1 U23911 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20993), .ZN(
        P1_U3178) );
  AND2_X1 U23912 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20993), .ZN(
        P1_U3179) );
  AND2_X1 U23913 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20993), .ZN(
        P1_U3180) );
  AND2_X1 U23914 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20993), .ZN(
        P1_U3181) );
  AND2_X1 U23915 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20993), .ZN(
        P1_U3182) );
  AND2_X1 U23916 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20993), .ZN(
        P1_U3183) );
  AND2_X1 U23917 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n21054), .ZN(
        P1_U3184) );
  AND2_X1 U23918 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n21054), .ZN(
        P1_U3185) );
  AND2_X1 U23919 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20993), .ZN(P1_U3186) );
  AND2_X1 U23920 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n21054), .ZN(P1_U3187) );
  AND2_X1 U23921 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21054), .ZN(P1_U3188) );
  AND2_X1 U23922 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n21054), .ZN(P1_U3189) );
  AND2_X1 U23923 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n21054), .ZN(P1_U3190) );
  AND2_X1 U23924 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21054), .ZN(P1_U3191) );
  AND2_X1 U23925 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n21054), .ZN(P1_U3192) );
  AND2_X1 U23926 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n21054), .ZN(P1_U3193) );
  NAND2_X1 U23927 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20998), .ZN(n21004) );
  INV_X1 U23928 ( .A(n21004), .ZN(n20997) );
  INV_X1 U23929 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21134) );
  NOR2_X1 U23930 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20994) );
  OAI22_X1 U23931 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21132), .B1(n20994), 
        .B2(n21002), .ZN(n20995) );
  OAI21_X1 U23932 ( .B1(n21134), .B2(n20995), .A(n21081), .ZN(n20996) );
  OAI21_X1 U23933 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n20997), .A(n20996), 
        .ZN(P1_U3194) );
  NOR2_X1 U23934 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21134), .ZN(n21001) );
  OAI33_X1 U23935 ( .A1(n21002), .A2(n21001), .A3(n21000), .B1(n20999), .B2(NA), .B3(n20998), .ZN(n21003) );
  OAI21_X1 U23936 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .A(n21003), 
        .ZN(n21006) );
  OAI211_X1 U23937 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n21132), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n21004), .ZN(n21005) );
  NAND2_X1 U23938 ( .A1(n21006), .A2(n21005), .ZN(P1_U3196) );
  NOR2_X1 U23939 ( .A1(n21007), .A2(n21081), .ZN(n21046) );
  AOI22_X1 U23940 ( .A1(P1_ADDRESS_REG_0__SCAN_IN), .A2(n21081), .B1(
        P1_REIP_REG_1__SCAN_IN), .B2(n21046), .ZN(n21008) );
  OAI21_X1 U23941 ( .B1(n21009), .B2(n21042), .A(n21008), .ZN(P1_U3197) );
  AOI22_X1 U23942 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n21081), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n21046), .ZN(n21010) );
  OAI21_X1 U23943 ( .B1(n21012), .B2(n21042), .A(n21010), .ZN(P1_U3198) );
  INV_X1 U23944 ( .A(n21046), .ZN(n21045) );
  OAI222_X1 U23945 ( .A1(n21045), .A2(n21012), .B1(n21011), .B2(n21038), .C1(
        n21332), .C2(n21042), .ZN(P1_U3199) );
  INV_X1 U23946 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n21013) );
  INV_X2 U23947 ( .A(n21043), .ZN(n21042) );
  OAI222_X1 U23948 ( .A1(n21045), .A2(n21332), .B1(n21013), .B2(n21038), .C1(
        n21014), .C2(n21042), .ZN(P1_U3200) );
  INV_X1 U23949 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n21015) );
  OAI222_X1 U23950 ( .A1(n21042), .A2(n21365), .B1(n21015), .B2(n21038), .C1(
        n21014), .C2(n21045), .ZN(P1_U3201) );
  INV_X1 U23951 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n21016) );
  OAI222_X1 U23952 ( .A1(n21045), .A2(n21365), .B1(n21016), .B2(n21038), .C1(
        n21379), .C2(n21042), .ZN(P1_U3202) );
  INV_X1 U23953 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n21017) );
  OAI222_X1 U23954 ( .A1(n21045), .A2(n21379), .B1(n21017), .B2(n21038), .C1(
        n21019), .C2(n21042), .ZN(P1_U3203) );
  INV_X1 U23955 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n21018) );
  OAI222_X1 U23956 ( .A1(n21045), .A2(n21019), .B1(n21018), .B2(n21038), .C1(
        n21381), .C2(n21042), .ZN(P1_U3204) );
  INV_X1 U23957 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n21020) );
  OAI222_X1 U23958 ( .A1(n21045), .A2(n21381), .B1(n21020), .B2(n21038), .C1(
        n21384), .C2(n21042), .ZN(P1_U3205) );
  INV_X1 U23959 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n21021) );
  OAI222_X1 U23960 ( .A1(n21045), .A2(n21384), .B1(n21021), .B2(n21038), .C1(
        n21302), .C2(n21042), .ZN(P1_U3206) );
  INV_X1 U23961 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n21022) );
  OAI222_X1 U23962 ( .A1(n21045), .A2(n21302), .B1(n21022), .B2(n21038), .C1(
        n21349), .C2(n21042), .ZN(P1_U3207) );
  INV_X1 U23963 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n21023) );
  OAI222_X1 U23964 ( .A1(n21045), .A2(n21349), .B1(n21023), .B2(n21038), .C1(
        n21382), .C2(n21042), .ZN(P1_U3208) );
  INV_X1 U23965 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n21024) );
  OAI222_X1 U23966 ( .A1(n21045), .A2(n21382), .B1(n21024), .B2(n21038), .C1(
        n21341), .C2(n21042), .ZN(P1_U3209) );
  INV_X1 U23967 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n21136) );
  INV_X1 U23968 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n21025) );
  OAI222_X1 U23969 ( .A1(n21042), .A2(n21136), .B1(n21025), .B2(n21038), .C1(
        n21341), .C2(n21045), .ZN(P1_U3210) );
  INV_X1 U23970 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n21400) );
  INV_X1 U23971 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n21026) );
  OAI222_X1 U23972 ( .A1(n21042), .A2(n21400), .B1(n21026), .B2(n21038), .C1(
        n21136), .C2(n21045), .ZN(P1_U3211) );
  AOI22_X1 U23973 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n21081), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n21043), .ZN(n21027) );
  OAI21_X1 U23974 ( .B1(n21400), .B2(n21045), .A(n21027), .ZN(P1_U3212) );
  AOI22_X1 U23975 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n21081), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n21046), .ZN(n21028) );
  OAI21_X1 U23976 ( .B1(n21378), .B2(n21042), .A(n21028), .ZN(P1_U3213) );
  INV_X1 U23977 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n21029) );
  OAI222_X1 U23978 ( .A1(n21045), .A2(n21378), .B1(n21029), .B2(n21038), .C1(
        n21162), .C2(n21042), .ZN(P1_U3214) );
  INV_X1 U23979 ( .A(P1_ADDRESS_REG_18__SCAN_IN), .ZN(n21030) );
  INV_X1 U23980 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n21210) );
  OAI222_X1 U23981 ( .A1(n21045), .A2(n21162), .B1(n21030), .B2(n21038), .C1(
        n21210), .C2(n21042), .ZN(P1_U3215) );
  INV_X1 U23982 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n21031) );
  OAI222_X1 U23983 ( .A1(n21042), .A2(n21369), .B1(n21031), .B2(n21038), .C1(
        n21210), .C2(n21045), .ZN(P1_U3216) );
  INV_X1 U23984 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n21032) );
  OAI222_X1 U23985 ( .A1(n21045), .A2(n21369), .B1(n21032), .B2(n21038), .C1(
        n21309), .C2(n21042), .ZN(P1_U3217) );
  INV_X1 U23986 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n21033) );
  INV_X1 U23987 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n21398) );
  OAI222_X1 U23988 ( .A1(n21045), .A2(n21309), .B1(n21033), .B2(n21038), .C1(
        n21398), .C2(n21042), .ZN(P1_U3218) );
  INV_X1 U23989 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n21034) );
  OAI222_X1 U23990 ( .A1(n21042), .A2(n21413), .B1(n21034), .B2(n21038), .C1(
        n21398), .C2(n21045), .ZN(P1_U3219) );
  INV_X1 U23991 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n21035) );
  OAI222_X1 U23992 ( .A1(n21045), .A2(n21413), .B1(n21035), .B2(n21038), .C1(
        n14592), .C2(n21042), .ZN(P1_U3220) );
  INV_X1 U23993 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n21036) );
  OAI222_X1 U23994 ( .A1(n21045), .A2(n14592), .B1(n21036), .B2(n21038), .C1(
        n21037), .C2(n21042), .ZN(P1_U3221) );
  INV_X1 U23995 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n21039) );
  OAI222_X1 U23996 ( .A1(n21042), .A2(n21412), .B1(n21039), .B2(n21038), .C1(
        n21037), .C2(n21045), .ZN(P1_U3222) );
  INV_X1 U23997 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n21040) );
  OAI222_X1 U23998 ( .A1(n21045), .A2(n21412), .B1(n21040), .B2(n21038), .C1(
        n21310), .C2(n21042), .ZN(P1_U3223) );
  INV_X1 U23999 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n21041) );
  OAI222_X1 U24000 ( .A1(n21042), .A2(n21408), .B1(n21041), .B2(n21038), .C1(
        n21310), .C2(n21045), .ZN(P1_U3224) );
  AOI22_X1 U24001 ( .A1(P1_ADDRESS_REG_28__SCAN_IN), .A2(n21081), .B1(
        P1_REIP_REG_30__SCAN_IN), .B2(n21043), .ZN(n21044) );
  OAI21_X1 U24002 ( .B1(n21408), .B2(n21045), .A(n21044), .ZN(P1_U3225) );
  AOI22_X1 U24003 ( .A1(P1_ADDRESS_REG_29__SCAN_IN), .A2(n21081), .B1(
        P1_REIP_REG_30__SCAN_IN), .B2(n21046), .ZN(n21047) );
  OAI21_X1 U24004 ( .B1(n21048), .B2(n21042), .A(n21047), .ZN(P1_U3226) );
  INV_X1 U24005 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n21049) );
  AOI22_X1 U24006 ( .A1(n21038), .A2(n21163), .B1(n21049), .B2(n21081), .ZN(
        P1_U3458) );
  INV_X1 U24007 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21150) );
  INV_X1 U24008 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n21050) );
  AOI22_X1 U24009 ( .A1(n21038), .A2(n21150), .B1(n21050), .B2(n21081), .ZN(
        P1_U3459) );
  INV_X1 U24010 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n21051) );
  AOI22_X1 U24011 ( .A1(n21038), .A2(n21362), .B1(n21051), .B2(n21081), .ZN(
        P1_U3460) );
  INV_X1 U24012 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21156) );
  INV_X1 U24013 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n21052) );
  AOI22_X1 U24014 ( .A1(n21038), .A2(n21156), .B1(n21052), .B2(n21081), .ZN(
        P1_U3461) );
  INV_X1 U24015 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n21055) );
  INV_X1 U24016 ( .A(n21056), .ZN(n21053) );
  AOI21_X1 U24017 ( .B1(n21055), .B2(n21054), .A(n21053), .ZN(P1_U3464) );
  OAI21_X1 U24018 ( .B1(n21058), .B2(n21057), .A(n21056), .ZN(P1_U3465) );
  AOI21_X1 U24019 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n21059) );
  AOI22_X1 U24020 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n21059), .B2(n21391), .ZN(n21060) );
  AOI22_X1 U24021 ( .A1(n21061), .A2(n21060), .B1(n21150), .B2(n21063), .ZN(
        P1_U3481) );
  NOR2_X1 U24022 ( .A1(n21063), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n21062) );
  AOI22_X1 U24023 ( .A1(n21156), .A2(n21063), .B1(n13697), .B2(n21062), .ZN(
        P1_U3482) );
  AOI22_X1 U24024 ( .A1(n21038), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21375), 
        .B2(n21081), .ZN(P1_U3483) );
  NAND2_X1 U24025 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21064), .ZN(n21072) );
  INV_X1 U24026 ( .A(n21065), .ZN(n21066) );
  OAI211_X1 U24027 ( .C1(n21072), .C2(n21068), .A(n21067), .B(n21066), .ZN(
        n21080) );
  AOI21_X1 U24028 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n21070), .A(n21069), 
        .ZN(n21071) );
  AOI211_X1 U24029 ( .C1(n21074), .C2(n21073), .A(n21072), .B(n21071), .ZN(
        n21076) );
  NOR2_X1 U24030 ( .A1(n21076), .A2(n21075), .ZN(n21078) );
  OAI21_X1 U24031 ( .B1(n21078), .B2(n21077), .A(n21080), .ZN(n21079) );
  OAI21_X1 U24032 ( .B1(n21080), .B2(n21134), .A(n21079), .ZN(P1_U3485) );
  INV_X1 U24033 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n21082) );
  AOI22_X1 U24034 ( .A1(n21038), .A2(n21392), .B1(n21082), .B2(n21081), .ZN(
        P1_U3486) );
  AOI22_X1 U24035 ( .A1(n16621), .A2(P3_ADDRESS_REG_29__SCAN_IN), .B1(
        P2_ADDRESS_REG_29__SCAN_IN), .B2(n16623), .ZN(n21470) );
  OAI22_X1 U24036 ( .A1(P1_EBX_REG_27__SCAN_IN), .A2(keyinput_g88), .B1(
        DATAI_21_), .B2(keyinput_g11), .ZN(n21083) );
  AOI221_X1 U24037 ( .B1(P1_EBX_REG_27__SCAN_IN), .B2(keyinput_g88), .C1(
        keyinput_g11), .C2(DATAI_21_), .A(n21083), .ZN(n21090) );
  OAI22_X1 U24038 ( .A1(DATAI_29_), .A2(keyinput_g3), .B1(P1_D_C_N_REG_SCAN_IN), .B2(keyinput_g42), .ZN(n21084) );
  AOI221_X1 U24039 ( .B1(DATAI_29_), .B2(keyinput_g3), .C1(keyinput_g42), .C2(
        P1_D_C_N_REG_SCAN_IN), .A(n21084), .ZN(n21089) );
  OAI22_X1 U24040 ( .A1(P1_EAX_REG_23__SCAN_IN), .A2(keyinput_g124), .B1(
        P1_EBX_REG_25__SCAN_IN), .B2(keyinput_g90), .ZN(n21085) );
  AOI221_X1 U24041 ( .B1(P1_EAX_REG_23__SCAN_IN), .B2(keyinput_g124), .C1(
        keyinput_g90), .C2(P1_EBX_REG_25__SCAN_IN), .A(n21085), .ZN(n21088) );
  OAI22_X1 U24042 ( .A1(DATAI_31_), .A2(keyinput_g1), .B1(keyinput_g32), .B2(
        DATAI_0_), .ZN(n21086) );
  AOI221_X1 U24043 ( .B1(DATAI_31_), .B2(keyinput_g1), .C1(DATAI_0_), .C2(
        keyinput_g32), .A(n21086), .ZN(n21087) );
  NAND4_X1 U24044 ( .A1(n21090), .A2(n21089), .A3(n21088), .A4(n21087), .ZN(
        n21222) );
  OAI22_X1 U24045 ( .A1(READY1), .A2(keyinput_g36), .B1(P1_REIP_REG_5__SCAN_IN), .B2(keyinput_g78), .ZN(n21091) );
  AOI221_X1 U24046 ( .B1(READY1), .B2(keyinput_g36), .C1(keyinput_g78), .C2(
        P1_REIP_REG_5__SCAN_IN), .A(n21091), .ZN(n21117) );
  OAI22_X1 U24047 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(keyinput_g81), .B1(
        keyinput_g20), .B2(DATAI_12_), .ZN(n21092) );
  AOI221_X1 U24048 ( .B1(P1_REIP_REG_2__SCAN_IN), .B2(keyinput_g81), .C1(
        DATAI_12_), .C2(keyinput_g20), .A(n21092), .ZN(n21095) );
  OAI22_X1 U24049 ( .A1(P1_EBX_REG_6__SCAN_IN), .A2(keyinput_g109), .B1(
        keyinput_g83), .B2(P1_REIP_REG_0__SCAN_IN), .ZN(n21093) );
  AOI221_X1 U24050 ( .B1(P1_EBX_REG_6__SCAN_IN), .B2(keyinput_g109), .C1(
        P1_REIP_REG_0__SCAN_IN), .C2(keyinput_g83), .A(n21093), .ZN(n21094) );
  OAI211_X1 U24051 ( .C1(n21097), .C2(keyinput_g98), .A(n21095), .B(n21094), 
        .ZN(n21096) );
  AOI21_X1 U24052 ( .B1(n21097), .B2(keyinput_g98), .A(n21096), .ZN(n21116) );
  AOI22_X1 U24053 ( .A1(READY2), .A2(keyinput_g37), .B1(P1_EAX_REG_25__SCAN_IN), .B2(keyinput_g122), .ZN(n21098) );
  OAI221_X1 U24054 ( .B1(READY2), .B2(keyinput_g37), .C1(
        P1_EAX_REG_25__SCAN_IN), .C2(keyinput_g122), .A(n21098), .ZN(n21105)
         );
  AOI22_X1 U24055 ( .A1(P1_EBX_REG_22__SCAN_IN), .A2(keyinput_g93), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(keyinput_g123), .ZN(n21099) );
  OAI221_X1 U24056 ( .B1(P1_EBX_REG_22__SCAN_IN), .B2(keyinput_g93), .C1(
        P1_EAX_REG_24__SCAN_IN), .C2(keyinput_g123), .A(n21099), .ZN(n21104)
         );
  AOI22_X1 U24057 ( .A1(P1_EBX_REG_14__SCAN_IN), .A2(keyinput_g101), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(keyinput_g126), .ZN(n21100) );
  OAI221_X1 U24058 ( .B1(P1_EBX_REG_14__SCAN_IN), .B2(keyinput_g101), .C1(
        P1_EAX_REG_21__SCAN_IN), .C2(keyinput_g126), .A(n21100), .ZN(n21103)
         );
  AOI22_X1 U24059 ( .A1(DATAI_18_), .A2(keyinput_g14), .B1(
        P1_EBX_REG_11__SCAN_IN), .B2(keyinput_g104), .ZN(n21101) );
  OAI221_X1 U24060 ( .B1(DATAI_18_), .B2(keyinput_g14), .C1(
        P1_EBX_REG_11__SCAN_IN), .C2(keyinput_g104), .A(n21101), .ZN(n21102)
         );
  NOR4_X1 U24061 ( .A1(n21105), .A2(n21104), .A3(n21103), .A4(n21102), .ZN(
        n21115) );
  AOI22_X1 U24062 ( .A1(DATAI_22_), .A2(keyinput_g10), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(keyinput_g66), .ZN(n21106) );
  OAI221_X1 U24063 ( .B1(DATAI_22_), .B2(keyinput_g10), .C1(
        P1_REIP_REG_17__SCAN_IN), .C2(keyinput_g66), .A(n21106), .ZN(n21113)
         );
  AOI22_X1 U24064 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(keyinput_g46), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(keyinput_g67), .ZN(n21107) );
  OAI221_X1 U24065 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(keyinput_g46), .C1(
        P1_REIP_REG_16__SCAN_IN), .C2(keyinput_g67), .A(n21107), .ZN(n21112)
         );
  AOI22_X1 U24066 ( .A1(BS16), .A2(keyinput_g35), .B1(P1_EBX_REG_30__SCAN_IN), 
        .B2(keyinput_g85), .ZN(n21108) );
  OAI221_X1 U24067 ( .B1(BS16), .B2(keyinput_g35), .C1(P1_EBX_REG_30__SCAN_IN), 
        .C2(keyinput_g85), .A(n21108), .ZN(n21111) );
  AOI22_X1 U24068 ( .A1(DATAI_15_), .A2(keyinput_g17), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(keyinput_g118), .ZN(n21109) );
  OAI221_X1 U24069 ( .B1(DATAI_15_), .B2(keyinput_g17), .C1(
        P1_EAX_REG_29__SCAN_IN), .C2(keyinput_g118), .A(n21109), .ZN(n21110)
         );
  NOR4_X1 U24070 ( .A1(n21113), .A2(n21112), .A3(n21111), .A4(n21110), .ZN(
        n21114) );
  NAND4_X1 U24071 ( .A1(n21117), .A2(n21116), .A3(n21115), .A4(n21114), .ZN(
        n21221) );
  INV_X1 U24072 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n21395) );
  AOI22_X1 U24073 ( .A1(DATAI_25_), .A2(keyinput_g7), .B1(n21395), .B2(
        keyinput_g38), .ZN(n21118) );
  OAI221_X1 U24074 ( .B1(DATAI_25_), .B2(keyinput_g7), .C1(n21395), .C2(
        keyinput_g38), .A(n21118), .ZN(n21127) );
  AOI22_X1 U24075 ( .A1(n21120), .A2(keyinput_g97), .B1(n21326), .B2(
        keyinput_g125), .ZN(n21119) );
  OAI221_X1 U24076 ( .B1(n21120), .B2(keyinput_g97), .C1(n21326), .C2(
        keyinput_g125), .A(n21119), .ZN(n21126) );
  AOI22_X1 U24077 ( .A1(n21413), .A2(keyinput_g59), .B1(keyinput_g9), .B2(
        n21122), .ZN(n21121) );
  OAI221_X1 U24078 ( .B1(n21413), .B2(keyinput_g59), .C1(n21122), .C2(
        keyinput_g9), .A(n21121), .ZN(n21125) );
  AOI22_X1 U24079 ( .A1(n21381), .A2(keyinput_g74), .B1(keyinput_g76), .B2(
        n21379), .ZN(n21123) );
  OAI221_X1 U24080 ( .B1(n21381), .B2(keyinput_g74), .C1(n21379), .C2(
        keyinput_g76), .A(n21123), .ZN(n21124) );
  NOR4_X1 U24081 ( .A1(n21127), .A2(n21126), .A3(n21125), .A4(n21124), .ZN(
        n21171) );
  INV_X1 U24082 ( .A(DATAI_11_), .ZN(n21129) );
  AOI22_X1 U24083 ( .A1(n21129), .A2(keyinput_g21), .B1(keyinput_g39), .B2(
        n21312), .ZN(n21128) );
  OAI221_X1 U24084 ( .B1(n21129), .B2(keyinput_g21), .C1(n21312), .C2(
        keyinput_g39), .A(n21128), .ZN(n21140) );
  AOI22_X1 U24085 ( .A1(n21132), .A2(keyinput_g34), .B1(n21131), .B2(
        keyinput_g103), .ZN(n21130) );
  OAI221_X1 U24086 ( .B1(n21132), .B2(keyinput_g34), .C1(n21131), .C2(
        keyinput_g103), .A(n21130), .ZN(n21139) );
  AOI22_X1 U24087 ( .A1(n21391), .A2(keyinput_g82), .B1(keyinput_g43), .B2(
        n21134), .ZN(n21133) );
  OAI221_X1 U24088 ( .B1(n21391), .B2(keyinput_g82), .C1(n21134), .C2(
        keyinput_g43), .A(n21133), .ZN(n21138) );
  AOI22_X1 U24089 ( .A1(n21366), .A2(keyinput_g8), .B1(n21136), .B2(
        keyinput_g68), .ZN(n21135) );
  OAI221_X1 U24090 ( .B1(n21366), .B2(keyinput_g8), .C1(n21136), .C2(
        keyinput_g68), .A(n21135), .ZN(n21137) );
  NOR4_X1 U24091 ( .A1(n21140), .A2(n21139), .A3(n21138), .A4(n21137), .ZN(
        n21170) );
  AOI22_X1 U24092 ( .A1(n21331), .A2(keyinput_g13), .B1(n21142), .B2(
        keyinput_g106), .ZN(n21141) );
  OAI221_X1 U24093 ( .B1(n21331), .B2(keyinput_g13), .C1(n21142), .C2(
        keyinput_g106), .A(n21141), .ZN(n21154) );
  INV_X1 U24094 ( .A(DATAI_6_), .ZN(n21144) );
  AOI22_X1 U24095 ( .A1(n21315), .A2(keyinput_g87), .B1(keyinput_g26), .B2(
        n21144), .ZN(n21143) );
  OAI221_X1 U24096 ( .B1(n21315), .B2(keyinput_g87), .C1(n21144), .C2(
        keyinput_g26), .A(n21143), .ZN(n21153) );
  INV_X1 U24097 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n21147) );
  AOI22_X1 U24098 ( .A1(n21147), .A2(keyinput_g45), .B1(n21146), .B2(
        keyinput_g4), .ZN(n21145) );
  OAI221_X1 U24099 ( .B1(n21147), .B2(keyinput_g45), .C1(n21146), .C2(
        keyinput_g4), .A(n21145), .ZN(n21152) );
  INV_X1 U24100 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n21149) );
  AOI22_X1 U24101 ( .A1(n21150), .A2(keyinput_g50), .B1(n21149), .B2(
        keyinput_g40), .ZN(n21148) );
  OAI221_X1 U24102 ( .B1(n21150), .B2(keyinput_g50), .C1(n21149), .C2(
        keyinput_g40), .A(n21148), .ZN(n21151) );
  NOR4_X1 U24103 ( .A1(n21154), .A2(n21153), .A3(n21152), .A4(n21151), .ZN(
        n21169) );
  AOI22_X1 U24104 ( .A1(n21369), .A2(keyinput_g62), .B1(keyinput_g48), .B2(
        n21156), .ZN(n21155) );
  OAI221_X1 U24105 ( .B1(n21369), .B2(keyinput_g62), .C1(n21156), .C2(
        keyinput_g48), .A(n21155), .ZN(n21167) );
  INV_X1 U24106 ( .A(DATAI_5_), .ZN(n21158) );
  AOI22_X1 U24107 ( .A1(n21300), .A2(keyinput_g84), .B1(keyinput_g27), .B2(
        n21158), .ZN(n21157) );
  OAI221_X1 U24108 ( .B1(n21300), .B2(keyinput_g84), .C1(n21158), .C2(
        keyinput_g27), .A(n21157), .ZN(n21166) );
  AOI22_X1 U24109 ( .A1(n21160), .A2(keyinput_g15), .B1(keyinput_g0), .B2(
        n21392), .ZN(n21159) );
  OAI221_X1 U24110 ( .B1(n21160), .B2(keyinput_g15), .C1(n21392), .C2(
        keyinput_g0), .A(n21159), .ZN(n21165) );
  AOI22_X1 U24111 ( .A1(n21163), .A2(keyinput_g51), .B1(n21162), .B2(
        keyinput_g64), .ZN(n21161) );
  OAI221_X1 U24112 ( .B1(n21163), .B2(keyinput_g51), .C1(n21162), .C2(
        keyinput_g64), .A(n21161), .ZN(n21164) );
  NOR4_X1 U24113 ( .A1(n21167), .A2(n21166), .A3(n21165), .A4(n21164), .ZN(
        n21168) );
  NAND4_X1 U24114 ( .A1(n21171), .A2(n21170), .A3(n21169), .A4(n21168), .ZN(
        n21220) );
  INV_X1 U24115 ( .A(DATAI_13_), .ZN(n21173) );
  AOI22_X1 U24116 ( .A1(n21173), .A2(keyinput_g19), .B1(n21365), .B2(
        keyinput_g77), .ZN(n21172) );
  OAI221_X1 U24117 ( .B1(n21173), .B2(keyinput_g19), .C1(n21365), .C2(
        keyinput_g77), .A(n21172), .ZN(n21183) );
  INV_X1 U24118 ( .A(DATAI_14_), .ZN(n21175) );
  AOI22_X1 U24119 ( .A1(n21175), .A2(keyinput_g18), .B1(n10025), .B2(
        keyinput_g108), .ZN(n21174) );
  OAI221_X1 U24120 ( .B1(n21175), .B2(keyinput_g18), .C1(n10025), .C2(
        keyinput_g108), .A(n21174), .ZN(n21182) );
  AOI22_X1 U24121 ( .A1(n21349), .A2(keyinput_g71), .B1(keyinput_g56), .B2(
        n21412), .ZN(n21176) );
  OAI221_X1 U24122 ( .B1(n21349), .B2(keyinput_g71), .C1(n21412), .C2(
        keyinput_g56), .A(n21176), .ZN(n21181) );
  AOI22_X1 U24123 ( .A1(n21179), .A2(keyinput_g117), .B1(keyinput_g2), .B2(
        n21178), .ZN(n21177) );
  OAI221_X1 U24124 ( .B1(n21179), .B2(keyinput_g117), .C1(n21178), .C2(
        keyinput_g2), .A(n21177), .ZN(n21180) );
  NOR4_X1 U24125 ( .A1(n21183), .A2(n21182), .A3(n21181), .A4(n21180), .ZN(
        n21218) );
  AOI22_X1 U24126 ( .A1(n10033), .A2(keyinput_g113), .B1(keyinput_g49), .B2(
        n21362), .ZN(n21184) );
  OAI221_X1 U24127 ( .B1(n10033), .B2(keyinput_g113), .C1(n21362), .C2(
        keyinput_g49), .A(n21184), .ZN(n21191) );
  INV_X1 U24128 ( .A(DATAI_3_), .ZN(n21342) );
  AOI22_X1 U24129 ( .A1(n21397), .A2(keyinput_g95), .B1(keyinput_g29), .B2(
        n21342), .ZN(n21185) );
  OAI221_X1 U24130 ( .B1(n21397), .B2(keyinput_g95), .C1(n21342), .C2(
        keyinput_g29), .A(n21185), .ZN(n21190) );
  INV_X1 U24131 ( .A(P1_EAX_REG_31__SCAN_IN), .ZN(n21303) );
  AOI22_X1 U24132 ( .A1(n21398), .A2(keyinput_g60), .B1(n21303), .B2(
        keyinput_g116), .ZN(n21186) );
  OAI221_X1 U24133 ( .B1(n21398), .B2(keyinput_g60), .C1(n21303), .C2(
        keyinput_g116), .A(n21186), .ZN(n21189) );
  AOI22_X1 U24134 ( .A1(n21309), .A2(keyinput_g61), .B1(n21341), .B2(
        keyinput_g69), .ZN(n21187) );
  OAI221_X1 U24135 ( .B1(n21309), .B2(keyinput_g61), .C1(n21341), .C2(
        keyinput_g69), .A(n21187), .ZN(n21188) );
  NOR4_X1 U24136 ( .A1(n21191), .A2(n21190), .A3(n21189), .A4(n21188), .ZN(
        n21217) );
  INV_X1 U24137 ( .A(DATAI_4_), .ZN(n21334) );
  AOI22_X1 U24138 ( .A1(n21334), .A2(keyinput_g28), .B1(n21378), .B2(
        keyinput_g65), .ZN(n21192) );
  OAI221_X1 U24139 ( .B1(n21334), .B2(keyinput_g28), .C1(n21378), .C2(
        keyinput_g65), .A(n21192), .ZN(n21203) );
  INV_X1 U24140 ( .A(DATAI_9_), .ZN(n21194) );
  AOI22_X1 U24141 ( .A1(n21195), .A2(keyinput_g92), .B1(keyinput_g23), .B2(
        n21194), .ZN(n21193) );
  OAI221_X1 U24142 ( .B1(n21195), .B2(keyinput_g92), .C1(n21194), .C2(
        keyinput_g23), .A(n21193), .ZN(n21202) );
  AOI22_X1 U24143 ( .A1(n21197), .A2(keyinput_g99), .B1(keyinput_g102), .B2(
        n21299), .ZN(n21196) );
  OAI221_X1 U24144 ( .B1(n21197), .B2(keyinput_g99), .C1(n21299), .C2(
        keyinput_g102), .A(n21196), .ZN(n21201) );
  AOI22_X1 U24145 ( .A1(n21199), .A2(keyinput_g112), .B1(keyinput_g47), .B2(
        n21375), .ZN(n21198) );
  OAI221_X1 U24146 ( .B1(n21199), .B2(keyinput_g112), .C1(n21375), .C2(
        keyinput_g47), .A(n21198), .ZN(n21200) );
  NOR4_X1 U24147 ( .A1(n21203), .A2(n21202), .A3(n21201), .A4(n21200), .ZN(
        n21216) );
  AOI22_X1 U24148 ( .A1(n21310), .A2(keyinput_g55), .B1(n21384), .B2(
        keyinput_g73), .ZN(n21204) );
  OAI221_X1 U24149 ( .B1(n21310), .B2(keyinput_g55), .C1(n21384), .C2(
        keyinput_g73), .A(n21204), .ZN(n21214) );
  AOI22_X1 U24150 ( .A1(n21206), .A2(keyinput_g119), .B1(keyinput_g72), .B2(
        n21302), .ZN(n21205) );
  OAI221_X1 U24151 ( .B1(n21206), .B2(keyinput_g119), .C1(n21302), .C2(
        keyinput_g72), .A(n21205), .ZN(n21213) );
  INV_X1 U24152 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n21208) );
  AOI22_X1 U24153 ( .A1(n21208), .A2(keyinput_g111), .B1(n21316), .B2(
        keyinput_g121), .ZN(n21207) );
  OAI221_X1 U24154 ( .B1(n21208), .B2(keyinput_g111), .C1(n21316), .C2(
        keyinput_g121), .A(n21207), .ZN(n21212) );
  AOI22_X1 U24155 ( .A1(n14592), .A2(keyinput_g58), .B1(n21210), .B2(
        keyinput_g63), .ZN(n21209) );
  OAI221_X1 U24156 ( .B1(n14592), .B2(keyinput_g58), .C1(n21210), .C2(
        keyinput_g63), .A(n21209), .ZN(n21211) );
  NOR4_X1 U24157 ( .A1(n21214), .A2(n21213), .A3(n21212), .A4(n21211), .ZN(
        n21215) );
  NAND4_X1 U24158 ( .A1(n21218), .A2(n21217), .A3(n21216), .A4(n21215), .ZN(
        n21219) );
  NOR4_X1 U24159 ( .A1(n21222), .A2(n21221), .A3(n21220), .A4(n21219), .ZN(
        n21260) );
  OAI22_X1 U24160 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(keyinput_g79), .B1(
        keyinput_g6), .B2(DATAI_26_), .ZN(n21223) );
  AOI221_X1 U24161 ( .B1(P1_REIP_REG_4__SCAN_IN), .B2(keyinput_g79), .C1(
        DATAI_26_), .C2(keyinput_g6), .A(n21223), .ZN(n21230) );
  OAI22_X1 U24162 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(keyinput_g57), .B1(
        DATAI_8_), .B2(keyinput_g24), .ZN(n21224) );
  AOI221_X1 U24163 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(keyinput_g57), .C1(
        keyinput_g24), .C2(DATAI_8_), .A(n21224), .ZN(n21229) );
  OAI22_X1 U24164 ( .A1(P1_EBX_REG_5__SCAN_IN), .A2(keyinput_g110), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(keyinput_g41), .ZN(n21225) );
  AOI221_X1 U24165 ( .B1(P1_EBX_REG_5__SCAN_IN), .B2(keyinput_g110), .C1(
        keyinput_g41), .C2(P1_M_IO_N_REG_SCAN_IN), .A(n21225), .ZN(n21228) );
  OAI22_X1 U24166 ( .A1(DATAI_27_), .A2(keyinput_g5), .B1(DATAI_7_), .B2(
        keyinput_g25), .ZN(n21226) );
  AOI221_X1 U24167 ( .B1(DATAI_27_), .B2(keyinput_g5), .C1(keyinput_g25), .C2(
        DATAI_7_), .A(n21226), .ZN(n21227) );
  NAND4_X1 U24168 ( .A1(n21230), .A2(n21229), .A3(n21228), .A4(n21227), .ZN(
        n21258) );
  OAI22_X1 U24169 ( .A1(P1_EBX_REG_26__SCAN_IN), .A2(keyinput_g89), .B1(
        keyinput_g91), .B2(P1_EBX_REG_24__SCAN_IN), .ZN(n21231) );
  AOI221_X1 U24170 ( .B1(P1_EBX_REG_26__SCAN_IN), .B2(keyinput_g89), .C1(
        P1_EBX_REG_24__SCAN_IN), .C2(keyinput_g91), .A(n21231), .ZN(n21238) );
  OAI22_X1 U24171 ( .A1(P1_EAX_REG_20__SCAN_IN), .A2(keyinput_g127), .B1(
        DATAI_2_), .B2(keyinput_g30), .ZN(n21232) );
  AOI221_X1 U24172 ( .B1(P1_EAX_REG_20__SCAN_IN), .B2(keyinput_g127), .C1(
        keyinput_g30), .C2(DATAI_2_), .A(n21232), .ZN(n21237) );
  OAI22_X1 U24173 ( .A1(P1_EBX_REG_1__SCAN_IN), .A2(keyinput_g114), .B1(
        P1_REIP_REG_29__SCAN_IN), .B2(keyinput_g54), .ZN(n21233) );
  AOI221_X1 U24174 ( .B1(P1_EBX_REG_1__SCAN_IN), .B2(keyinput_g114), .C1(
        keyinput_g54), .C2(P1_REIP_REG_29__SCAN_IN), .A(n21233), .ZN(n21236)
         );
  OAI22_X1 U24175 ( .A1(P1_REIP_REG_31__SCAN_IN), .A2(keyinput_g52), .B1(
        DATAI_20_), .B2(keyinput_g12), .ZN(n21234) );
  AOI221_X1 U24176 ( .B1(P1_REIP_REG_31__SCAN_IN), .B2(keyinput_g52), .C1(
        keyinput_g12), .C2(DATAI_20_), .A(n21234), .ZN(n21235) );
  NAND4_X1 U24177 ( .A1(n21238), .A2(n21237), .A3(n21236), .A4(n21235), .ZN(
        n21257) );
  OAI22_X1 U24178 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(keyinput_g53), .B1(
        keyinput_g16), .B2(DATAI_16_), .ZN(n21239) );
  AOI221_X1 U24179 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(keyinput_g53), .C1(
        DATAI_16_), .C2(keyinput_g16), .A(n21239), .ZN(n21246) );
  OAI22_X1 U24180 ( .A1(P1_EBX_REG_21__SCAN_IN), .A2(keyinput_g94), .B1(
        keyinput_g100), .B2(P1_EBX_REG_15__SCAN_IN), .ZN(n21240) );
  AOI221_X1 U24181 ( .B1(P1_EBX_REG_21__SCAN_IN), .B2(keyinput_g94), .C1(
        P1_EBX_REG_15__SCAN_IN), .C2(keyinput_g100), .A(n21240), .ZN(n21245)
         );
  OAI22_X1 U24182 ( .A1(P1_EBX_REG_29__SCAN_IN), .A2(keyinput_g86), .B1(
        DATAI_1_), .B2(keyinput_g31), .ZN(n21241) );
  AOI221_X1 U24183 ( .B1(P1_EBX_REG_29__SCAN_IN), .B2(keyinput_g86), .C1(
        keyinput_g31), .C2(DATAI_1_), .A(n21241), .ZN(n21244) );
  OAI22_X1 U24184 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(keyinput_g70), .B1(
        keyinput_g22), .B2(DATAI_10_), .ZN(n21242) );
  AOI221_X1 U24185 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(keyinput_g70), .C1(
        DATAI_10_), .C2(keyinput_g22), .A(n21242), .ZN(n21243) );
  NAND4_X1 U24186 ( .A1(n21246), .A2(n21245), .A3(n21244), .A4(n21243), .ZN(
        n21256) );
  OAI22_X1 U24187 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(keyinput_g44), .B1(
        keyinput_g107), .B2(P1_EBX_REG_8__SCAN_IN), .ZN(n21247) );
  AOI221_X1 U24188 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(keyinput_g44), .C1(
        P1_EBX_REG_8__SCAN_IN), .C2(keyinput_g107), .A(n21247), .ZN(n21254) );
  OAI22_X1 U24189 ( .A1(P1_EBX_REG_19__SCAN_IN), .A2(keyinput_g96), .B1(
        keyinput_g33), .B2(HOLD), .ZN(n21248) );
  AOI221_X1 U24190 ( .B1(P1_EBX_REG_19__SCAN_IN), .B2(keyinput_g96), .C1(HOLD), 
        .C2(keyinput_g33), .A(n21248), .ZN(n21253) );
  OAI22_X1 U24191 ( .A1(P1_EAX_REG_27__SCAN_IN), .A2(keyinput_g120), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(keyinput_g80), .ZN(n21249) );
  AOI221_X1 U24192 ( .B1(P1_EAX_REG_27__SCAN_IN), .B2(keyinput_g120), .C1(
        keyinput_g80), .C2(P1_REIP_REG_3__SCAN_IN), .A(n21249), .ZN(n21252) );
  OAI22_X1 U24193 ( .A1(P1_EBX_REG_10__SCAN_IN), .A2(keyinput_g105), .B1(
        keyinput_g75), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n21250) );
  AOI221_X1 U24194 ( .B1(P1_EBX_REG_10__SCAN_IN), .B2(keyinput_g105), .C1(
        P1_REIP_REG_8__SCAN_IN), .C2(keyinput_g75), .A(n21250), .ZN(n21251) );
  NAND4_X1 U24195 ( .A1(n21254), .A2(n21253), .A3(n21252), .A4(n21251), .ZN(
        n21255) );
  NOR4_X1 U24196 ( .A1(n21258), .A2(n21257), .A3(n21256), .A4(n21255), .ZN(
        n21259) );
  AOI22_X1 U24197 ( .A1(n21260), .A2(n21259), .B1(keyinput_g115), .B2(n12903), 
        .ZN(n21468) );
  OAI22_X1 U24198 ( .A1(P1_EAX_REG_20__SCAN_IN), .A2(keyinput_f127), .B1(
        keyinput_f41), .B2(P1_M_IO_N_REG_SCAN_IN), .ZN(n21261) );
  AOI221_X1 U24199 ( .B1(P1_EAX_REG_20__SCAN_IN), .B2(keyinput_f127), .C1(
        P1_M_IO_N_REG_SCAN_IN), .C2(keyinput_f41), .A(n21261), .ZN(n21268) );
  OAI22_X1 U24200 ( .A1(P1_EAX_REG_24__SCAN_IN), .A2(keyinput_f123), .B1(
        keyinput_f19), .B2(DATAI_13_), .ZN(n21262) );
  AOI221_X1 U24201 ( .B1(P1_EAX_REG_24__SCAN_IN), .B2(keyinput_f123), .C1(
        DATAI_13_), .C2(keyinput_f19), .A(n21262), .ZN(n21267) );
  OAI22_X1 U24202 ( .A1(P1_REIP_REG_31__SCAN_IN), .A2(keyinput_f52), .B1(
        DATAI_9_), .B2(keyinput_f23), .ZN(n21263) );
  AOI221_X1 U24203 ( .B1(P1_REIP_REG_31__SCAN_IN), .B2(keyinput_f52), .C1(
        keyinput_f23), .C2(DATAI_9_), .A(n21263), .ZN(n21266) );
  OAI22_X1 U24204 ( .A1(P1_EBX_REG_1__SCAN_IN), .A2(keyinput_f114), .B1(BS16), 
        .B2(keyinput_f35), .ZN(n21264) );
  AOI221_X1 U24205 ( .B1(P1_EBX_REG_1__SCAN_IN), .B2(keyinput_f114), .C1(
        keyinput_f35), .C2(BS16), .A(n21264), .ZN(n21265) );
  NAND4_X1 U24206 ( .A1(n21268), .A2(n21267), .A3(n21266), .A4(n21265), .ZN(
        n21427) );
  OAI22_X1 U24207 ( .A1(P1_EAX_REG_28__SCAN_IN), .A2(keyinput_f119), .B1(NA), 
        .B2(keyinput_f34), .ZN(n21269) );
  AOI221_X1 U24208 ( .B1(P1_EAX_REG_28__SCAN_IN), .B2(keyinput_f119), .C1(
        keyinput_f34), .C2(NA), .A(n21269), .ZN(n21295) );
  OAI22_X1 U24209 ( .A1(P1_EBX_REG_2__SCAN_IN), .A2(keyinput_f113), .B1(
        keyinput_f68), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n21270) );
  AOI221_X1 U24210 ( .B1(P1_EBX_REG_2__SCAN_IN), .B2(keyinput_f113), .C1(
        P1_REIP_REG_15__SCAN_IN), .C2(keyinput_f68), .A(n21270), .ZN(n21273)
         );
  OAI22_X1 U24211 ( .A1(P1_EBX_REG_15__SCAN_IN), .A2(keyinput_f100), .B1(
        keyinput_f57), .B2(P1_REIP_REG_26__SCAN_IN), .ZN(n21271) );
  AOI221_X1 U24212 ( .B1(P1_EBX_REG_15__SCAN_IN), .B2(keyinput_f100), .C1(
        P1_REIP_REG_26__SCAN_IN), .C2(keyinput_f57), .A(n21271), .ZN(n21272)
         );
  OAI211_X1 U24213 ( .C1(n21275), .C2(keyinput_f3), .A(n21273), .B(n21272), 
        .ZN(n21274) );
  AOI21_X1 U24214 ( .B1(n21275), .B2(keyinput_f3), .A(n21274), .ZN(n21294) );
  AOI22_X1 U24215 ( .A1(DATAI_5_), .A2(keyinput_f27), .B1(DATAI_22_), .B2(
        keyinput_f10), .ZN(n21276) );
  OAI221_X1 U24216 ( .B1(DATAI_5_), .B2(keyinput_f27), .C1(DATAI_22_), .C2(
        keyinput_f10), .A(n21276), .ZN(n21283) );
  AOI22_X1 U24217 ( .A1(P1_EBX_REG_16__SCAN_IN), .A2(keyinput_f99), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(keyinput_f117), .ZN(n21277) );
  OAI221_X1 U24218 ( .B1(P1_EBX_REG_16__SCAN_IN), .B2(keyinput_f99), .C1(
        P1_EAX_REG_30__SCAN_IN), .C2(keyinput_f117), .A(n21277), .ZN(n21282)
         );
  AOI22_X1 U24219 ( .A1(DATAI_0_), .A2(keyinput_f32), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(keyinput_f118), .ZN(n21278) );
  OAI221_X1 U24220 ( .B1(DATAI_0_), .B2(keyinput_f32), .C1(
        P1_EAX_REG_29__SCAN_IN), .C2(keyinput_f118), .A(n21278), .ZN(n21281)
         );
  AOI22_X1 U24221 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(keyinput_f40), .B1(
        P1_EBX_REG_23__SCAN_IN), .B2(keyinput_f92), .ZN(n21279) );
  OAI221_X1 U24222 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(keyinput_f40), .C1(
        P1_EBX_REG_23__SCAN_IN), .C2(keyinput_f92), .A(n21279), .ZN(n21280) );
  NOR4_X1 U24223 ( .A1(n21283), .A2(n21282), .A3(n21281), .A4(n21280), .ZN(
        n21293) );
  AOI22_X1 U24224 ( .A1(DATAI_11_), .A2(keyinput_f21), .B1(
        P1_EBX_REG_12__SCAN_IN), .B2(keyinput_f103), .ZN(n21284) );
  OAI221_X1 U24225 ( .B1(DATAI_11_), .B2(keyinput_f21), .C1(
        P1_EBX_REG_12__SCAN_IN), .C2(keyinput_f103), .A(n21284), .ZN(n21291)
         );
  AOI22_X1 U24226 ( .A1(P1_MORE_REG_SCAN_IN), .A2(keyinput_f45), .B1(
        P1_EBX_REG_18__SCAN_IN), .B2(keyinput_f97), .ZN(n21285) );
  OAI221_X1 U24227 ( .B1(P1_MORE_REG_SCAN_IN), .B2(keyinput_f45), .C1(
        P1_EBX_REG_18__SCAN_IN), .C2(keyinput_f97), .A(n21285), .ZN(n21290) );
  AOI22_X1 U24228 ( .A1(DATAI_20_), .A2(keyinput_f12), .B1(
        P1_EBX_REG_26__SCAN_IN), .B2(keyinput_f89), .ZN(n21286) );
  OAI221_X1 U24229 ( .B1(DATAI_20_), .B2(keyinput_f12), .C1(
        P1_EBX_REG_26__SCAN_IN), .C2(keyinput_f89), .A(n21286), .ZN(n21289) );
  AOI22_X1 U24230 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(keyinput_f80), .B1(
        P1_EBX_REG_7__SCAN_IN), .B2(keyinput_f108), .ZN(n21287) );
  OAI221_X1 U24231 ( .B1(P1_REIP_REG_3__SCAN_IN), .B2(keyinput_f80), .C1(
        P1_EBX_REG_7__SCAN_IN), .C2(keyinput_f108), .A(n21287), .ZN(n21288) );
  NOR4_X1 U24232 ( .A1(n21291), .A2(n21290), .A3(n21289), .A4(n21288), .ZN(
        n21292) );
  NAND4_X1 U24233 ( .A1(n21295), .A2(n21294), .A3(n21293), .A4(n21292), .ZN(
        n21426) );
  AOI22_X1 U24234 ( .A1(DATAI_8_), .A2(keyinput_f24), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(keyinput_f66), .ZN(n21296) );
  OAI221_X1 U24235 ( .B1(DATAI_8_), .B2(keyinput_f24), .C1(
        P1_REIP_REG_17__SCAN_IN), .C2(keyinput_f66), .A(n21296), .ZN(n21307)
         );
  AOI22_X1 U24236 ( .A1(DATAI_21_), .A2(keyinput_f11), .B1(DATAI_25_), .B2(
        keyinput_f7), .ZN(n21297) );
  OAI221_X1 U24237 ( .B1(DATAI_21_), .B2(keyinput_f11), .C1(DATAI_25_), .C2(
        keyinput_f7), .A(n21297), .ZN(n21306) );
  AOI22_X1 U24238 ( .A1(n21300), .A2(keyinput_f84), .B1(n21299), .B2(
        keyinput_f102), .ZN(n21298) );
  OAI221_X1 U24239 ( .B1(n21300), .B2(keyinput_f84), .C1(n21299), .C2(
        keyinput_f102), .A(n21298), .ZN(n21305) );
  AOI22_X1 U24240 ( .A1(n21303), .A2(keyinput_f116), .B1(keyinput_f72), .B2(
        n21302), .ZN(n21301) );
  OAI221_X1 U24241 ( .B1(n21303), .B2(keyinput_f116), .C1(n21302), .C2(
        keyinput_f72), .A(n21301), .ZN(n21304) );
  NOR4_X1 U24242 ( .A1(n21307), .A2(n21306), .A3(n21305), .A4(n21304), .ZN(
        n21358) );
  AOI22_X1 U24243 ( .A1(n21310), .A2(keyinput_f55), .B1(n21309), .B2(
        keyinput_f61), .ZN(n21308) );
  OAI221_X1 U24244 ( .B1(n21310), .B2(keyinput_f55), .C1(n21309), .C2(
        keyinput_f61), .A(n21308), .ZN(n21323) );
  AOI22_X1 U24245 ( .A1(n21313), .A2(keyinput_f88), .B1(keyinput_f39), .B2(
        n21312), .ZN(n21311) );
  OAI221_X1 U24246 ( .B1(n21313), .B2(keyinput_f88), .C1(n21312), .C2(
        keyinput_f39), .A(n21311), .ZN(n21322) );
  AOI22_X1 U24247 ( .A1(n21316), .A2(keyinput_f121), .B1(keyinput_f87), .B2(
        n21315), .ZN(n21314) );
  OAI221_X1 U24248 ( .B1(n21316), .B2(keyinput_f121), .C1(n21315), .C2(
        keyinput_f87), .A(n21314), .ZN(n21321) );
  AOI22_X1 U24249 ( .A1(n21319), .A2(keyinput_f46), .B1(n21318), .B2(
        keyinput_f104), .ZN(n21317) );
  OAI221_X1 U24250 ( .B1(n21319), .B2(keyinput_f46), .C1(n21318), .C2(
        keyinput_f104), .A(n21317), .ZN(n21320) );
  NOR4_X1 U24251 ( .A1(n21323), .A2(n21322), .A3(n21321), .A4(n21320), .ZN(
        n21357) );
  AOI22_X1 U24252 ( .A1(n21326), .A2(keyinput_f125), .B1(keyinput_f90), .B2(
        n21325), .ZN(n21324) );
  OAI221_X1 U24253 ( .B1(n21326), .B2(keyinput_f125), .C1(n21325), .C2(
        keyinput_f90), .A(n21324), .ZN(n21339) );
  INV_X1 U24254 ( .A(READY2), .ZN(n21329) );
  INV_X1 U24255 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n21328) );
  AOI22_X1 U24256 ( .A1(n21329), .A2(keyinput_f37), .B1(n21328), .B2(
        keyinput_f109), .ZN(n21327) );
  OAI221_X1 U24257 ( .B1(n21329), .B2(keyinput_f37), .C1(n21328), .C2(
        keyinput_f109), .A(n21327), .ZN(n21338) );
  AOI22_X1 U24258 ( .A1(n21332), .A2(keyinput_f79), .B1(keyinput_f13), .B2(
        n21331), .ZN(n21330) );
  OAI221_X1 U24259 ( .B1(n21332), .B2(keyinput_f79), .C1(n21331), .C2(
        keyinput_f13), .A(n21330), .ZN(n21337) );
  INV_X1 U24260 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n21335) );
  AOI22_X1 U24261 ( .A1(n21335), .A2(keyinput_f105), .B1(keyinput_f28), .B2(
        n21334), .ZN(n21333) );
  OAI221_X1 U24262 ( .B1(n21335), .B2(keyinput_f105), .C1(n21334), .C2(
        keyinput_f28), .A(n21333), .ZN(n21336) );
  NOR4_X1 U24263 ( .A1(n21339), .A2(n21338), .A3(n21337), .A4(n21336), .ZN(
        n21356) );
  AOI22_X1 U24264 ( .A1(n21342), .A2(keyinput_f29), .B1(n21341), .B2(
        keyinput_f69), .ZN(n21340) );
  OAI221_X1 U24265 ( .B1(n21342), .B2(keyinput_f29), .C1(n21341), .C2(
        keyinput_f69), .A(n21340), .ZN(n21354) );
  INV_X1 U24266 ( .A(keyinput_f42), .ZN(n21344) );
  AOI22_X1 U24267 ( .A1(n10036), .A2(keyinput_f107), .B1(P1_D_C_N_REG_SCAN_IN), 
        .B2(n21344), .ZN(n21343) );
  OAI221_X1 U24268 ( .B1(n10036), .B2(keyinput_f107), .C1(n21344), .C2(
        P1_D_C_N_REG_SCAN_IN), .A(n21343), .ZN(n21353) );
  INV_X1 U24269 ( .A(DATAI_10_), .ZN(n21346) );
  AOI22_X1 U24270 ( .A1(n21347), .A2(keyinput_f16), .B1(n21346), .B2(
        keyinput_f22), .ZN(n21345) );
  OAI221_X1 U24271 ( .B1(n21347), .B2(keyinput_f16), .C1(n21346), .C2(
        keyinput_f22), .A(n21345), .ZN(n21352) );
  AOI22_X1 U24272 ( .A1(n21350), .A2(keyinput_f120), .B1(keyinput_f71), .B2(
        n21349), .ZN(n21348) );
  OAI221_X1 U24273 ( .B1(n21350), .B2(keyinput_f120), .C1(n21349), .C2(
        keyinput_f71), .A(n21348), .ZN(n21351) );
  NOR4_X1 U24274 ( .A1(n21354), .A2(n21353), .A3(n21352), .A4(n21351), .ZN(
        n21355) );
  NAND4_X1 U24275 ( .A1(n21358), .A2(n21357), .A3(n21356), .A4(n21355), .ZN(
        n21425) );
  INV_X1 U24276 ( .A(DATAI_2_), .ZN(n21360) );
  AOI22_X1 U24277 ( .A1(n21360), .A2(keyinput_f30), .B1(n10028), .B2(
        keyinput_f96), .ZN(n21359) );
  OAI221_X1 U24278 ( .B1(n21360), .B2(keyinput_f30), .C1(n10028), .C2(
        keyinput_f96), .A(n21359), .ZN(n21373) );
  AOI22_X1 U24279 ( .A1(n21363), .A2(keyinput_f91), .B1(keyinput_f49), .B2(
        n21362), .ZN(n21361) );
  OAI221_X1 U24280 ( .B1(n21363), .B2(keyinput_f91), .C1(n21362), .C2(
        keyinput_f49), .A(n21361), .ZN(n21372) );
  AOI22_X1 U24281 ( .A1(n21366), .A2(keyinput_f8), .B1(n21365), .B2(
        keyinput_f77), .ZN(n21364) );
  OAI221_X1 U24282 ( .B1(n21366), .B2(keyinput_f8), .C1(n21365), .C2(
        keyinput_f77), .A(n21364), .ZN(n21371) );
  INV_X1 U24283 ( .A(DATAI_12_), .ZN(n21368) );
  AOI22_X1 U24284 ( .A1(n21369), .A2(keyinput_f62), .B1(keyinput_f20), .B2(
        n21368), .ZN(n21367) );
  OAI221_X1 U24285 ( .B1(n21369), .B2(keyinput_f62), .C1(n21368), .C2(
        keyinput_f20), .A(n21367), .ZN(n21370) );
  NOR4_X1 U24286 ( .A1(n21373), .A2(n21372), .A3(n21371), .A4(n21370), .ZN(
        n21423) );
  AOI22_X1 U24287 ( .A1(n21376), .A2(keyinput_f110), .B1(keyinput_f47), .B2(
        n21375), .ZN(n21374) );
  OAI221_X1 U24288 ( .B1(n21376), .B2(keyinput_f110), .C1(n21375), .C2(
        keyinput_f47), .A(n21374), .ZN(n21389) );
  AOI22_X1 U24289 ( .A1(n21379), .A2(keyinput_f76), .B1(keyinput_f65), .B2(
        n21378), .ZN(n21377) );
  OAI221_X1 U24290 ( .B1(n21379), .B2(keyinput_f76), .C1(n21378), .C2(
        keyinput_f65), .A(n21377), .ZN(n21388) );
  AOI22_X1 U24291 ( .A1(n21382), .A2(keyinput_f70), .B1(keyinput_f74), .B2(
        n21381), .ZN(n21380) );
  OAI221_X1 U24292 ( .B1(n21382), .B2(keyinput_f70), .C1(n21381), .C2(
        keyinput_f74), .A(n21380), .ZN(n21387) );
  AOI22_X1 U24293 ( .A1(n21385), .A2(keyinput_f85), .B1(keyinput_f73), .B2(
        n21384), .ZN(n21383) );
  OAI221_X1 U24294 ( .B1(n21385), .B2(keyinput_f85), .C1(n21384), .C2(
        keyinput_f73), .A(n21383), .ZN(n21386) );
  NOR4_X1 U24295 ( .A1(n21389), .A2(n21388), .A3(n21387), .A4(n21386), .ZN(
        n21422) );
  AOI22_X1 U24296 ( .A1(n21392), .A2(keyinput_f0), .B1(n21391), .B2(
        keyinput_f82), .ZN(n21390) );
  OAI221_X1 U24297 ( .B1(n21392), .B2(keyinput_f0), .C1(n21391), .C2(
        keyinput_f82), .A(n21390), .ZN(n21405) );
  AOI22_X1 U24298 ( .A1(n21395), .A2(keyinput_f38), .B1(n21394), .B2(
        keyinput_f25), .ZN(n21393) );
  OAI221_X1 U24299 ( .B1(n21395), .B2(keyinput_f38), .C1(n21394), .C2(
        keyinput_f25), .A(n21393), .ZN(n21404) );
  AOI22_X1 U24300 ( .A1(n21398), .A2(keyinput_f60), .B1(n21397), .B2(
        keyinput_f95), .ZN(n21396) );
  OAI221_X1 U24301 ( .B1(n21398), .B2(keyinput_f60), .C1(n21397), .C2(
        keyinput_f95), .A(n21396), .ZN(n21403) );
  INV_X1 U24302 ( .A(DATAI_1_), .ZN(n21401) );
  AOI22_X1 U24303 ( .A1(n21401), .A2(keyinput_f31), .B1(n21400), .B2(
        keyinput_f67), .ZN(n21399) );
  OAI221_X1 U24304 ( .B1(n21401), .B2(keyinput_f31), .C1(n21400), .C2(
        keyinput_f67), .A(n21399), .ZN(n21402) );
  NOR4_X1 U24305 ( .A1(n21405), .A2(n21404), .A3(n21403), .A4(n21402), .ZN(
        n21421) );
  INV_X1 U24306 ( .A(READY1), .ZN(n21407) );
  AOI22_X1 U24307 ( .A1(n21408), .A2(keyinput_f54), .B1(n21407), .B2(
        keyinput_f36), .ZN(n21406) );
  OAI221_X1 U24308 ( .B1(n21408), .B2(keyinput_f54), .C1(n21407), .C2(
        keyinput_f36), .A(n21406), .ZN(n21419) );
  AOI22_X1 U24309 ( .A1(n13744), .A2(keyinput_f17), .B1(n21410), .B2(
        keyinput_f86), .ZN(n21409) );
  OAI221_X1 U24310 ( .B1(n13744), .B2(keyinput_f17), .C1(n21410), .C2(
        keyinput_f86), .A(n21409), .ZN(n21418) );
  AOI22_X1 U24311 ( .A1(n21413), .A2(keyinput_f59), .B1(keyinput_f56), .B2(
        n21412), .ZN(n21411) );
  OAI221_X1 U24312 ( .B1(n21413), .B2(keyinput_f59), .C1(n21412), .C2(
        keyinput_f56), .A(n21411), .ZN(n21417) );
  AOI22_X1 U24313 ( .A1(n14422), .A2(keyinput_f93), .B1(keyinput_f94), .B2(
        n21415), .ZN(n21414) );
  OAI221_X1 U24314 ( .B1(n14422), .B2(keyinput_f93), .C1(n21415), .C2(
        keyinput_f94), .A(n21414), .ZN(n21416) );
  NOR4_X1 U24315 ( .A1(n21419), .A2(n21418), .A3(n21417), .A4(n21416), .ZN(
        n21420) );
  NAND4_X1 U24316 ( .A1(n21423), .A2(n21422), .A3(n21421), .A4(n21420), .ZN(
        n21424) );
  NOR4_X1 U24317 ( .A1(n21427), .A2(n21426), .A3(n21425), .A4(n21424), .ZN(
        n21465) );
  OAI22_X1 U24318 ( .A1(DATAI_14_), .A2(keyinput_f18), .B1(keyinput_f43), .B2(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21428) );
  AOI221_X1 U24319 ( .B1(DATAI_14_), .B2(keyinput_f18), .C1(
        P1_REQUESTPENDING_REG_SCAN_IN), .C2(keyinput_f43), .A(n21428), .ZN(
        n21435) );
  OAI22_X1 U24320 ( .A1(P1_EBX_REG_9__SCAN_IN), .A2(keyinput_f106), .B1(
        DATAI_26_), .B2(keyinput_f6), .ZN(n21429) );
  AOI221_X1 U24321 ( .B1(P1_EBX_REG_9__SCAN_IN), .B2(keyinput_f106), .C1(
        keyinput_f6), .C2(DATAI_26_), .A(n21429), .ZN(n21434) );
  OAI22_X1 U24322 ( .A1(P1_EBX_REG_14__SCAN_IN), .A2(keyinput_f101), .B1(
        keyinput_f15), .B2(DATAI_17_), .ZN(n21430) );
  AOI221_X1 U24323 ( .B1(P1_EBX_REG_14__SCAN_IN), .B2(keyinput_f101), .C1(
        DATAI_17_), .C2(keyinput_f15), .A(n21430), .ZN(n21433) );
  OAI22_X1 U24324 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(keyinput_f75), .B1(
        DATAI_27_), .B2(keyinput_f5), .ZN(n21431) );
  AOI221_X1 U24325 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(keyinput_f75), .C1(
        keyinput_f5), .C2(DATAI_27_), .A(n21431), .ZN(n21432) );
  NAND4_X1 U24326 ( .A1(n21435), .A2(n21434), .A3(n21433), .A4(n21432), .ZN(
        n21463) );
  OAI22_X1 U24327 ( .A1(P1_EBX_REG_4__SCAN_IN), .A2(keyinput_f111), .B1(
        P1_REIP_REG_30__SCAN_IN), .B2(keyinput_f53), .ZN(n21436) );
  AOI221_X1 U24328 ( .B1(P1_EBX_REG_4__SCAN_IN), .B2(keyinput_f111), .C1(
        keyinput_f53), .C2(P1_REIP_REG_30__SCAN_IN), .A(n21436), .ZN(n21443)
         );
  OAI22_X1 U24329 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(keyinput_f58), .B1(
        DATAI_28_), .B2(keyinput_f4), .ZN(n21437) );
  AOI221_X1 U24330 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(keyinput_f58), .C1(
        keyinput_f4), .C2(DATAI_28_), .A(n21437), .ZN(n21442) );
  OAI22_X1 U24331 ( .A1(P1_EAX_REG_25__SCAN_IN), .A2(keyinput_f122), .B1(
        DATAI_6_), .B2(keyinput_f26), .ZN(n21438) );
  AOI221_X1 U24332 ( .B1(P1_EAX_REG_25__SCAN_IN), .B2(keyinput_f122), .C1(
        keyinput_f26), .C2(DATAI_6_), .A(n21438), .ZN(n21441) );
  OAI22_X1 U24333 ( .A1(DATAI_31_), .A2(keyinput_f1), .B1(
        P1_BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_f48), .ZN(n21439) );
  AOI221_X1 U24334 ( .B1(DATAI_31_), .B2(keyinput_f1), .C1(keyinput_f48), .C2(
        P1_BYTEENABLE_REG_0__SCAN_IN), .A(n21439), .ZN(n21440) );
  NAND4_X1 U24335 ( .A1(n21443), .A2(n21442), .A3(n21441), .A4(n21440), .ZN(
        n21462) );
  OAI22_X1 U24336 ( .A1(P1_EBX_REG_17__SCAN_IN), .A2(keyinput_f98), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(keyinput_f78), .ZN(n21444) );
  AOI221_X1 U24337 ( .B1(P1_EBX_REG_17__SCAN_IN), .B2(keyinput_f98), .C1(
        keyinput_f78), .C2(P1_REIP_REG_5__SCAN_IN), .A(n21444), .ZN(n21451) );
  OAI22_X1 U24338 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(keyinput_f81), .B1(
        keyinput_f51), .B2(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21445) );
  AOI221_X1 U24339 ( .B1(P1_REIP_REG_2__SCAN_IN), .B2(keyinput_f81), .C1(
        P1_BYTEENABLE_REG_3__SCAN_IN), .C2(keyinput_f51), .A(n21445), .ZN(
        n21450) );
  OAI22_X1 U24340 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(keyinput_f63), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(keyinput_f64), .ZN(n21446) );
  AOI221_X1 U24341 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(keyinput_f63), .C1(
        keyinput_f64), .C2(P1_REIP_REG_19__SCAN_IN), .A(n21446), .ZN(n21449)
         );
  OAI22_X1 U24342 ( .A1(P1_EBX_REG_3__SCAN_IN), .A2(keyinput_f112), .B1(
        keyinput_f83), .B2(P1_REIP_REG_0__SCAN_IN), .ZN(n21447) );
  AOI221_X1 U24343 ( .B1(P1_EBX_REG_3__SCAN_IN), .B2(keyinput_f112), .C1(
        P1_REIP_REG_0__SCAN_IN), .C2(keyinput_f83), .A(n21447), .ZN(n21448) );
  NAND4_X1 U24344 ( .A1(n21451), .A2(n21450), .A3(n21449), .A4(n21448), .ZN(
        n21461) );
  OAI22_X1 U24345 ( .A1(DATAI_30_), .A2(keyinput_f2), .B1(keyinput_f9), .B2(
        DATAI_23_), .ZN(n21452) );
  AOI221_X1 U24346 ( .B1(DATAI_30_), .B2(keyinput_f2), .C1(DATAI_23_), .C2(
        keyinput_f9), .A(n21452), .ZN(n21459) );
  OAI22_X1 U24347 ( .A1(DATAI_18_), .A2(keyinput_f14), .B1(keyinput_f50), .B2(
        P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21453) );
  AOI221_X1 U24348 ( .B1(DATAI_18_), .B2(keyinput_f14), .C1(
        P1_BYTEENABLE_REG_2__SCAN_IN), .C2(keyinput_f50), .A(n21453), .ZN(
        n21458) );
  OAI22_X1 U24349 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(keyinput_f44), .B1(HOLD), .B2(keyinput_f33), .ZN(n21454) );
  AOI221_X1 U24350 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(keyinput_f44), .C1(
        keyinput_f33), .C2(HOLD), .A(n21454), .ZN(n21457) );
  OAI22_X1 U24351 ( .A1(P1_EAX_REG_21__SCAN_IN), .A2(keyinput_f126), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(keyinput_f124), .ZN(n21455) );
  AOI221_X1 U24352 ( .B1(P1_EAX_REG_21__SCAN_IN), .B2(keyinput_f126), .C1(
        keyinput_f124), .C2(P1_EAX_REG_23__SCAN_IN), .A(n21455), .ZN(n21456)
         );
  NAND4_X1 U24353 ( .A1(n21459), .A2(n21458), .A3(n21457), .A4(n21456), .ZN(
        n21460) );
  NOR4_X1 U24354 ( .A1(n21463), .A2(n21462), .A3(n21461), .A4(n21460), .ZN(
        n21464) );
  AOI22_X1 U24355 ( .A1(n21465), .A2(n21464), .B1(keyinput_f115), .B2(n12903), 
        .ZN(n21466) );
  OAI21_X1 U24356 ( .B1(keyinput_f115), .B2(n12903), .A(n21466), .ZN(n21467)
         );
  OAI211_X1 U24357 ( .C1(keyinput_g115), .C2(n12903), .A(n21468), .B(n21467), 
        .ZN(n21469) );
  XOR2_X1 U24358 ( .A(n21470), .B(n21469), .Z(U355) );
  INV_X2 U11347 ( .A(n14639), .ZN(n16018) );
  CLKBUF_X1 U11276 ( .A(n12344), .Z(n12861) );
  AND2_X1 U11296 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13924) );
  CLKBUF_X1 U11318 ( .A(n11952), .Z(n11953) );
  CLKBUF_X2 U11325 ( .A(n10567), .Z(n10588) );
  INV_X1 U11353 ( .A(n11025), .ZN(n9820) );
  CLKBUF_X1 U11368 ( .A(n10706), .Z(n19440) );
  AND2_X1 U11382 ( .A1(n10617), .A2(n10626), .ZN(n10823) );
  CLKBUF_X3 U11486 ( .A(n10589), .Z(n14253) );
  XNOR2_X1 U11491 ( .A(n10186), .B(n11119), .ZN(n9833) );
  CLKBUF_X1 U11527 ( .A(n10597), .Z(n10607) );
  CLKBUF_X2 U11647 ( .A(n16949), .Z(n16991) );
  CLKBUF_X1 U12366 ( .A(n9887), .Z(n17197) );
  CLKBUF_X1 U12807 ( .A(n11929), .Z(n20443) );
endmodule

