

module b14_C_SARLock_k_128_4 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3352, 
        U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, 
        U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, 
        U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, 
        U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, 
        U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, 
        U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, 
        U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, 
        U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, 
        U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, 
        U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, 
        U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, 
        U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, 
        U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, 
        U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, 
        U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, 
        U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, 
        U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, 
        U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, 
        U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, 
        U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, 
        U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, 
        U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, 
        U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, 
        U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, 
        U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867;

  INV_X2 U2413 ( .A(n4517), .ZN(n4781) );
  CLKBUF_X2 U2414 ( .A(n2804), .Z(n2919) );
  AND2_X1 U2415 ( .A1(n3918), .A2(n4186), .ZN(n4476) );
  CLKBUF_X2 U2416 ( .A(n2804), .Z(n2953) );
  AOI21_X1 U2417 ( .B1(n3063), .B2(REG2_REG_3__SCAN_IN), .A(n2292), .ZN(n3064)
         );
  INV_X2 U2418 ( .A(n2956), .ZN(n2791) );
  INV_X1 U2419 ( .A(IR_REG_31__SCAN_IN), .ZN(n2663) );
  AND2_X1 U2420 ( .A1(n3308), .A2(n3307), .ZN(n3309) );
  NAND2_X1 U2421 ( .A1(n2931), .A2(n2930), .ZN(n3939) );
  AOI21_X1 U2422 ( .B1(n3226), .B2(n3225), .A(n2830), .ZN(n3233) );
  XOR2_X1 U2423 ( .A(n4656), .B(n4655), .Z(n4668) );
  NAND2_X1 U2424 ( .A1(n2214), .A2(n4074), .ZN(n3269) );
  XNOR2_X2 U2425 ( .A(n4266), .B(n4822), .ZN(n4690) );
  NAND2_X2 U2426 ( .A1(n4678), .A2(n4265), .ZN(n4266) );
  NAND2_X2 U2427 ( .A1(n4747), .A2(n4275), .ZN(n4277) );
  XNOR2_X2 U2428 ( .A(n2665), .B(n2664), .ZN(n2677) );
  AOI21_X2 U2429 ( .B1(n3085), .B2(REG2_REG_6__SCAN_IN), .A(n2287), .ZN(n3087)
         );
  NOR2_X2 U2430 ( .A1(n3309), .A2(n2352), .ZN(n3604) );
  BUF_X4 U2431 ( .A(n2413), .Z(n2732) );
  OAI21_X2 U2432 ( .B1(n4264), .B2(n4263), .A(n2283), .ZN(n4679) );
  CLKBUF_X3 U2433 ( .A(n2423), .Z(n2170) );
  AND2_X1 U2434 ( .A1(n2381), .A2(n3023), .ZN(n2423) );
  OAI21_X1 U2435 ( .B1(n3269), .B2(n2708), .A(n4079), .ZN(n3299) );
  INV_X2 U2437 ( .A(n4235), .ZN(U4043) );
  NOR2_X2 U2438 ( .A1(n3257), .A2(n3222), .ZN(n3221) );
  NAND4_X1 U2439 ( .A1(n2408), .A2(n2407), .A3(n2406), .A4(n2405), .ZN(n4236)
         );
  INV_X1 U2440 ( .A(n3255), .ZN(n3118) );
  NAND2_X1 U2441 ( .A1(n2422), .A2(REG3_REG_1__SCAN_IN), .ZN(n2389) );
  NAND2_X1 U2442 ( .A1(n2683), .A2(n2594), .ZN(n4648) );
  NOR2_X1 U2443 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2368)
         );
  NOR2_X1 U2444 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2225)
         );
  AND2_X1 U2445 ( .A1(n2342), .A2(n2196), .ZN(n3000) );
  NAND2_X1 U2446 ( .A1(n3967), .A2(n2945), .ZN(n2344) );
  AND2_X1 U2447 ( .A1(n2211), .A2(n2210), .ZN(n2765) );
  NAND2_X1 U2448 ( .A1(n4005), .A2(n2339), .ZN(n2338) );
  NAND2_X1 U2449 ( .A1(n4755), .A2(n4753), .ZN(n4754) );
  NAND2_X1 U2450 ( .A1(n4327), .A2(n2218), .ZN(n4522) );
  NAND2_X1 U2451 ( .A1(n2207), .A2(n2206), .ZN(n3918) );
  AOI21_X1 U2452 ( .B1(n3917), .B2(n2571), .A(n2570), .ZN(n4497) );
  NAND2_X1 U2453 ( .A1(n4419), .A2(n4408), .ZN(n4407) );
  NAND2_X1 U2454 ( .A1(n4698), .A2(n4268), .ZN(n4269) );
  NAND2_X1 U2455 ( .A1(n2215), .A2(n4080), .ZN(n3664) );
  NAND2_X2 U2456 ( .A1(n2702), .A2(n4420), .ZN(n4517) );
  INV_X2 U2457 ( .A(n2866), .ZN(n2959) );
  CLKBUF_X1 U2458 ( .A(n2866), .Z(n2963) );
  NAND2_X1 U2459 ( .A1(n3596), .A2(n2187), .ZN(n3662) );
  AND2_X1 U2460 ( .A1(n3171), .A2(n2284), .ZN(n3061) );
  NAND2_X1 U2461 ( .A1(n2191), .A2(n2176), .ZN(n3247) );
  NAND4_X2 U2462 ( .A1(n2391), .A2(n2390), .A3(n2389), .A4(n2388), .ZN(n2790)
         );
  INV_X1 U2464 ( .A(n3027), .ZN(n3015) );
  INV_X1 U2465 ( .A(n2736), .ZN(n4212) );
  XNOR2_X1 U2466 ( .A(n2293), .B(n3051), .ZN(n3063) );
  AND2_X1 U2467 ( .A1(n2293), .A2(n3062), .ZN(n2292) );
  NAND2_X1 U2468 ( .A1(n2681), .A2(IR_REG_31__SCAN_IN), .ZN(n2665) );
  OAI21_X1 U2469 ( .B1(n2591), .B2(IR_REG_18__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2593) );
  NAND2_X1 U2470 ( .A1(n3933), .A2(IR_REG_31__SCAN_IN), .ZN(n2377) );
  NAND2_X1 U2471 ( .A1(n2680), .A2(n2682), .ZN(n2681) );
  XNOR2_X1 U2472 ( .A(n2686), .B(IR_REG_22__SCAN_IN), .ZN(n4631) );
  NAND2_X1 U2473 ( .A1(n4247), .A2(n2188), .ZN(n2293) );
  AND2_X1 U2474 ( .A1(n2670), .A2(n2375), .ZN(n2376) );
  AND2_X1 U2475 ( .A1(n2666), .A2(n2374), .ZN(n2670) );
  AND2_X2 U2476 ( .A1(n2393), .A2(n3438), .ZN(n2366) );
  NOR2_X2 U2477 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2666)
         );
  INV_X1 U2478 ( .A(IR_REG_24__SCAN_IN), .ZN(n2664) );
  NOR2_X1 U2479 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2226)
         );
  AND2_X2 U2480 ( .A1(n4378), .A2(n4198), .ZN(n4358) );
  INV_X1 U2481 ( .A(n2778), .ZN(n2171) );
  INV_X1 U2482 ( .A(n2171), .ZN(n2172) );
  NOR2_X2 U2483 ( .A1(n4366), .A2(n4342), .ZN(n4347) );
  NOR2_X2 U2484 ( .A1(n3061), .A2(n3060), .ZN(n3078) );
  NAND2_X2 U2485 ( .A1(n2738), .A2(n4212), .ZN(n2777) );
  XNOR2_X2 U2486 ( .A(n2685), .B(n2684), .ZN(n2738) );
  NOR2_X4 U2487 ( .A1(n3776), .A2(n3794), .ZN(n2227) );
  NAND2_X2 U2488 ( .A1(n3729), .A2(n3799), .ZN(n3776) );
  OAI21_X2 U2489 ( .B1(n2687), .B2(n2345), .A(IR_REG_31__SCAN_IN), .ZN(n2729)
         );
  NAND2_X2 U2490 ( .A1(n2216), .A2(n2182), .ZN(n2687) );
  INV_X1 U2491 ( .A(IR_REG_27__SCAN_IN), .ZN(n2280) );
  AOI21_X1 U2492 ( .B1(n2235), .B2(n2237), .A(n2234), .ZN(n2233) );
  INV_X1 U2493 ( .A(n4132), .ZN(n2234) );
  INV_X1 U2494 ( .A(n2238), .ZN(n2235) );
  NOR2_X1 U2495 ( .A1(n2242), .A2(n2195), .ZN(n2241) );
  OR2_X1 U2496 ( .A1(n4236), .A2(n3214), .ZN(n4069) );
  NOR2_X1 U2497 ( .A1(n2246), .A2(n2358), .ZN(n2245) );
  INV_X1 U2498 ( .A(IR_REG_23__SCAN_IN), .ZN(n2682) );
  INV_X1 U2499 ( .A(n2537), .ZN(n2216) );
  NOR2_X1 U2500 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2372)
         );
  AND2_X1 U2501 ( .A1(n4631), .A2(n4212), .ZN(n3029) );
  NAND2_X1 U2502 ( .A1(n4006), .A2(n4007), .ZN(n4005) );
  XNOR2_X1 U2503 ( .A(n2807), .B(n2956), .ZN(n2809) );
  NAND2_X1 U2504 ( .A1(n4699), .A2(n4700), .ZN(n4698) );
  XNOR2_X1 U2505 ( .A(n4297), .B(n2286), .ZN(n4712) );
  NAND2_X1 U2506 ( .A1(n2255), .A2(n2197), .ZN(n2746) );
  NOR2_X1 U2507 ( .A1(n2647), .A2(n2251), .ZN(n2250) );
  NOR2_X1 U2508 ( .A1(n4332), .A2(n4342), .ZN(n2251) );
  AND2_X1 U2509 ( .A1(n2655), .A2(n2654), .ZN(n4325) );
  NAND2_X1 U2510 ( .A1(n4381), .A2(n4367), .ZN(n2631) );
  NAND2_X1 U2511 ( .A1(n2261), .A2(n2264), .ZN(n2260) );
  OR2_X1 U2512 ( .A1(n4543), .A2(n4408), .ZN(n2264) );
  NAND2_X1 U2513 ( .A1(n2175), .A2(n2353), .ZN(n2261) );
  NAND2_X1 U2514 ( .A1(n2712), .A2(n4082), .ZN(n3649) );
  AND2_X1 U2515 ( .A1(n2738), .A2(n3098), .ZN(n4829) );
  INV_X1 U2516 ( .A(n4133), .ZN(n2231) );
  NAND2_X1 U2517 ( .A1(n4476), .A2(n4188), .ZN(n4454) );
  AND2_X1 U2518 ( .A1(n2194), .A2(n4504), .ZN(n2238) );
  NAND2_X1 U2519 ( .A1(n2178), .A2(n2194), .ZN(n2237) );
  NAND2_X1 U2520 ( .A1(n3701), .A2(n4102), .ZN(n3771) );
  NAND2_X1 U2521 ( .A1(n2790), .A2(n2793), .ZN(n4066) );
  NAND2_X1 U2522 ( .A1(n2376), .A2(n2346), .ZN(n2345) );
  INV_X1 U2523 ( .A(n2347), .ZN(n2346) );
  INV_X1 U2524 ( .A(IR_REG_26__SCAN_IN), .ZN(n2375) );
  NAND2_X1 U2525 ( .A1(n2373), .A2(n2348), .ZN(n2347) );
  INV_X1 U2526 ( .A(IR_REG_22__SCAN_IN), .ZN(n2373) );
  INV_X1 U2527 ( .A(IR_REG_21__SCAN_IN), .ZN(n2348) );
  AOI21_X1 U2528 ( .B1(n2174), .B2(n2173), .A(n2204), .ZN(n2302) );
  XNOR2_X1 U2529 ( .A(n2787), .B(n2791), .ZN(n2818) );
  NAND2_X1 U2530 ( .A1(n2786), .A2(n2785), .ZN(n2787) );
  NAND2_X1 U2531 ( .A1(n2331), .A2(n2330), .ZN(n2329) );
  INV_X1 U2532 ( .A(n4029), .ZN(n2330) );
  INV_X1 U2533 ( .A(n4028), .ZN(n2331) );
  AOI22_X1 U2534 ( .A1(n2790), .A2(n2804), .B1(n2789), .B2(n3256), .ZN(n2792)
         );
  XNOR2_X1 U2535 ( .A(n2781), .B(n2791), .ZN(n2820) );
  NAND2_X1 U2536 ( .A1(n2780), .A2(n2779), .ZN(n2781) );
  INV_X1 U2537 ( .A(n4051), .ZN(n2324) );
  AND2_X1 U2538 ( .A1(n3978), .A2(n2322), .ZN(n2321) );
  OR2_X1 U2539 ( .A1(n2893), .A2(n2324), .ZN(n2322) );
  NOR2_X1 U2540 ( .A1(n2172), .A2(n4826), .ZN(n2795) );
  NOR2_X1 U2541 ( .A1(n2984), .A2(n2969), .ZN(n2988) );
  NOR2_X1 U2542 ( .A1(n4020), .A2(n2337), .ZN(n2336) );
  INV_X1 U2543 ( .A(n3957), .ZN(n2337) );
  AOI21_X1 U2544 ( .B1(n2311), .B2(n2314), .A(n2190), .ZN(n2309) );
  XNOR2_X1 U2545 ( .A(n2826), .B(n2791), .ZN(n2827) );
  NAND2_X1 U2546 ( .A1(n2987), .A2(STATE_REG_SCAN_IN), .ZN(n4021) );
  NAND2_X1 U2547 ( .A1(n2732), .A2(REG0_REG_3__SCAN_IN), .ZN(n2427) );
  INV_X1 U2548 ( .A(n4654), .ZN(n4218) );
  OR2_X1 U2549 ( .A1(n3069), .A2(n3068), .ZN(n2291) );
  NAND2_X1 U2550 ( .A1(n2291), .A2(n2290), .ZN(n2289) );
  NAND2_X1 U2551 ( .A1(n4635), .A2(REG2_REG_5__SCAN_IN), .ZN(n2290) );
  NAND2_X1 U2552 ( .A1(n4679), .A2(n4680), .ZN(n4678) );
  NAND2_X1 U2553 ( .A1(n4681), .A2(n4292), .ZN(n4294) );
  XNOR2_X1 U2554 ( .A(n4304), .B(n4276), .ZN(n4755) );
  NOR2_X1 U2555 ( .A1(n4742), .A2(n2294), .ZN(n4304) );
  AND2_X1 U2556 ( .A1(n4303), .A2(REG2_REG_15__SCAN_IN), .ZN(n2294) );
  NOR2_X1 U2557 ( .A1(n2203), .A2(n2223), .ZN(n3042) );
  INV_X1 U2558 ( .A(n2402), .ZN(n2223) );
  NAND2_X1 U2559 ( .A1(n2632), .A2(n2253), .ZN(n2252) );
  NOR2_X1 U2560 ( .A1(n2641), .A2(n2254), .ZN(n2253) );
  INV_X1 U2561 ( .A(n2355), .ZN(n2254) );
  NOR2_X1 U2562 ( .A1(n2618), .A2(n4000), .ZN(n2624) );
  OR2_X1 U2563 ( .A1(n2260), .A2(n2263), .ZN(n2258) );
  AND2_X1 U2564 ( .A1(n4363), .A2(n4389), .ZN(n2263) );
  AND2_X1 U2565 ( .A1(n4414), .A2(n2175), .ZN(n2259) );
  NOR2_X1 U2566 ( .A1(n2262), .A2(n4171), .ZN(n4416) );
  INV_X1 U2567 ( .A(n4414), .ZN(n2262) );
  NAND2_X1 U2568 ( .A1(n3875), .A2(n2559), .ZN(n3917) );
  AOI21_X1 U2569 ( .B1(n2245), .B2(n2243), .A(n2199), .ZN(n2242) );
  INV_X1 U2570 ( .A(n2359), .ZN(n2243) );
  INV_X1 U2571 ( .A(n2245), .ZN(n2244) );
  AOI21_X1 U2572 ( .B1(n2278), .B2(n2276), .A(n2200), .ZN(n2275) );
  INV_X1 U2573 ( .A(n2278), .ZN(n2277) );
  OAI22_X1 U2574 ( .A1(n3651), .A2(n2486), .B1(n3657), .B2(n3759), .ZN(n3726)
         );
  OAI21_X1 U2575 ( .B1(n3664), .B2(n2710), .A(n4083), .ZN(n3638) );
  OR2_X1 U2576 ( .A1(n4831), .A2(n4212), .ZN(n2983) );
  NAND2_X1 U2577 ( .A1(n3202), .A2(n3200), .ZN(n2214) );
  INV_X1 U2578 ( .A(n4514), .ZN(n4486) );
  AND2_X1 U2579 ( .A1(n3243), .A2(n2403), .ZN(n3211) );
  NOR2_X1 U2580 ( .A1(n3247), .A2(n3118), .ZN(n4068) );
  NAND2_X1 U2581 ( .A1(n4654), .A2(n3029), .ZN(n4482) );
  AND2_X1 U2582 ( .A1(n2737), .A2(n2736), .ZN(n3098) );
  AND2_X1 U2583 ( .A1(n3031), .A2(n2985), .ZN(n3114) );
  NOR2_X2 U2584 ( .A1(n4522), .A2(n4525), .ZN(n4655) );
  NAND2_X1 U2585 ( .A1(n2640), .A2(DATAI_24_), .ZN(n4542) );
  AND2_X1 U2586 ( .A1(n4632), .A2(n3098), .ZN(n4658) );
  AND2_X1 U2587 ( .A1(n3842), .A2(n4831), .ZN(n4590) );
  NAND2_X1 U2588 ( .A1(n2273), .A2(n2272), .ZN(n4848) );
  INV_X1 U2589 ( .A(n4142), .ZN(n2272) );
  INV_X1 U2590 ( .A(n3673), .ZN(n2273) );
  OR2_X1 U2591 ( .A1(n4654), .A2(n2741), .ZN(n4578) );
  OR2_X1 U2592 ( .A1(n4783), .A2(n4631), .ZN(n4831) );
  NAND2_X1 U2593 ( .A1(n2673), .A2(n2678), .ZN(n3025) );
  OR2_X1 U2594 ( .A1(n2378), .A2(n2663), .ZN(n2380) );
  NAND2_X1 U2595 ( .A1(n2683), .A2(IR_REG_31__SCAN_IN), .ZN(n2685) );
  AND3_X1 U2596 ( .A1(n2367), .A2(n2366), .A3(n2332), .ZN(n2528) );
  NOR2_X1 U2597 ( .A1(n2334), .A2(IR_REG_10__SCAN_IN), .ZN(n2332) );
  AND3_X1 U2598 ( .A1(n2621), .A2(n2620), .A3(n2619), .ZN(n4543) );
  INV_X1 U2599 ( .A(n4059), .ZN(n4043) );
  INV_X1 U2600 ( .A(n2810), .ZN(n2811) );
  NAND2_X1 U2601 ( .A1(n2639), .A2(n2638), .ZN(n4332) );
  OAI211_X1 U2602 ( .C1(n4421), .C2(n2630), .A(n2615), .B(n2614), .ZN(n4403)
         );
  XNOR2_X1 U2603 ( .A(n4294), .B(n4822), .ZN(n4692) );
  NAND2_X1 U2604 ( .A1(n4692), .A2(REG2_REG_10__SCAN_IN), .ZN(n4691) );
  AND2_X1 U2605 ( .A1(n4675), .A2(n3043), .ZN(n4711) );
  XNOR2_X1 U2606 ( .A(n4269), .B(n2286), .ZN(n4717) );
  NAND2_X1 U2607 ( .A1(n4710), .A2(n4298), .ZN(n4723) );
  NOR2_X1 U2608 ( .A1(n4744), .A2(n4743), .ZN(n4742) );
  XNOR2_X1 U2609 ( .A(n4277), .B(n4276), .ZN(n4758) );
  NOR2_X1 U2610 ( .A1(n4758), .A2(REG1_REG_16__SCAN_IN), .ZN(n4759) );
  NAND2_X1 U2611 ( .A1(n4768), .A2(ADDR_REG_18__SCAN_IN), .ZN(n2298) );
  INV_X1 U2612 ( .A(n4637), .ZN(n2300) );
  AOI21_X1 U2613 ( .B1(n4307), .B2(n4308), .A(n4762), .ZN(n2299) );
  AND2_X1 U2614 ( .A1(n4675), .A2(n3168), .ZN(n4769) );
  AOI22_X1 U2615 ( .A1(n2746), .A2(n4131), .B1(n2656), .B2(n4228), .ZN(n2661)
         );
  OR2_X1 U2616 ( .A1(n2774), .A2(n4493), .ZN(n2220) );
  NAND2_X1 U2617 ( .A1(n4523), .A2(n4226), .ZN(n2210) );
  NAND2_X1 U2618 ( .A1(n2212), .A2(n4514), .ZN(n2211) );
  XNOR2_X1 U2619 ( .A(n2213), .B(n4165), .ZN(n2212) );
  XNOR2_X1 U2620 ( .A(n2746), .B(n4131), .ZN(n4320) );
  AND2_X1 U2621 ( .A1(n4517), .A2(n4658), .ZN(n4446) );
  NAND2_X1 U2622 ( .A1(n2701), .A2(n3031), .ZN(n4420) );
  INV_X1 U2623 ( .A(n2983), .ZN(n2701) );
  AND2_X1 U2624 ( .A1(n2271), .A2(n2465), .ZN(n2270) );
  NAND2_X1 U2625 ( .A1(n2181), .A2(n2274), .ZN(n2271) );
  AOI21_X1 U2626 ( .B1(n2431), .B2(n3203), .A(n2430), .ZN(n3274) );
  INV_X1 U2627 ( .A(IR_REG_28__SCAN_IN), .ZN(n2387) );
  NAND2_X1 U2628 ( .A1(n2729), .A2(n2387), .ZN(n2281) );
  OR2_X1 U2629 ( .A1(n3618), .A2(n3665), .ZN(n2274) );
  NOR2_X1 U2630 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2370)
         );
  NOR2_X1 U2631 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2371)
         );
  INV_X1 U2632 ( .A(n3828), .ZN(n2303) );
  INV_X1 U2633 ( .A(n2866), .ZN(n2796) );
  AND2_X1 U2634 ( .A1(n4453), .A2(n2724), .ZN(n4191) );
  AOI21_X1 U2635 ( .B1(n4143), .B2(n2509), .A(n2183), .ZN(n2278) );
  INV_X1 U2636 ( .A(n2509), .ZN(n2276) );
  NAND2_X1 U2637 ( .A1(n2270), .A2(n2267), .ZN(n2266) );
  INV_X1 U2638 ( .A(n2274), .ZN(n2267) );
  NAND2_X1 U2639 ( .A1(n2402), .A2(DATAI_30_), .ZN(n4177) );
  OR2_X2 U2640 ( .A1(n3662), .A2(n3678), .ZN(n2360) );
  OAI21_X1 U2641 ( .B1(n3591), .B2(n2181), .A(n2274), .ZN(n3673) );
  INV_X1 U2642 ( .A(IR_REG_20__SCAN_IN), .ZN(n2684) );
  INV_X1 U2643 ( .A(IR_REG_15__SCAN_IN), .ZN(n2554) );
  OR2_X1 U2644 ( .A1(n2568), .A2(n2663), .ZN(n2555) );
  INV_X1 U2645 ( .A(n2368), .ZN(n2334) );
  INV_X1 U2646 ( .A(IR_REG_1__SCAN_IN), .ZN(n3407) );
  INV_X1 U2647 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3941) );
  NOR2_X1 U2648 ( .A1(n2476), .A2(n2363), .ZN(n2487) );
  NAND2_X1 U2649 ( .A1(n2327), .A2(n2325), .ZN(n3947) );
  NOR2_X1 U2650 ( .A1(n3949), .A2(n2326), .ZN(n2325) );
  INV_X1 U2651 ( .A(n2328), .ZN(n2326) );
  INV_X1 U2652 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2584) );
  NAND2_X1 U2653 ( .A1(n2344), .A2(n2343), .ZN(n2342) );
  AND2_X1 U2654 ( .A1(n2201), .A2(n4039), .ZN(n2343) );
  INV_X1 U2655 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2510) );
  NAND2_X1 U2656 ( .A1(n3939), .A2(n2317), .ZN(n3996) );
  NOR2_X1 U2657 ( .A1(n2936), .A2(n2318), .ZN(n2317) );
  INV_X1 U2658 ( .A(n2934), .ZN(n2318) );
  NAND2_X1 U2659 ( .A1(n2845), .A2(n2844), .ZN(n2316) );
  NAND2_X1 U2660 ( .A1(n3606), .A2(n3605), .ZN(n2315) );
  AND2_X1 U2661 ( .A1(n3692), .A2(n2312), .ZN(n2311) );
  NAND2_X1 U2662 ( .A1(n2313), .A2(n2315), .ZN(n2312) );
  INV_X1 U2663 ( .A(n2316), .ZN(n2313) );
  INV_X1 U2664 ( .A(n2315), .ZN(n2314) );
  AOI21_X1 U2665 ( .B1(n2184), .B2(n3788), .A(n2306), .ZN(n2305) );
  AND2_X1 U2666 ( .A1(n3787), .A2(n2307), .ZN(n2306) );
  NOR2_X1 U2667 ( .A1(n3956), .A2(n2340), .ZN(n2339) );
  INV_X1 U2668 ( .A(n4009), .ZN(n2340) );
  INV_X1 U2669 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2500) );
  OAI21_X1 U2670 ( .B1(n2402), .B2(n2412), .A(n2221), .ZN(n3214) );
  NAND2_X1 U2671 ( .A1(n2402), .A2(n2411), .ZN(n2221) );
  OR2_X1 U2672 ( .A1(n2892), .A2(n2893), .ZN(n4049) );
  NAND2_X1 U2673 ( .A1(n2892), .A2(n2893), .ZN(n4048) );
  INV_X1 U2674 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2541) );
  OR2_X1 U2675 ( .A1(n2991), .A2(n4218), .ZN(n4022) );
  OR2_X1 U2676 ( .A1(n2404), .A2(n2799), .ZN(n2398) );
  NAND2_X1 U2677 ( .A1(n4249), .A2(n4248), .ZN(n4247) );
  NAND2_X1 U2678 ( .A1(n3172), .A2(REG1_REG_4__SCAN_IN), .ZN(n3171) );
  OR2_X1 U2679 ( .A1(n3089), .A2(n2285), .ZN(n3155) );
  AND2_X1 U2680 ( .A1(n3090), .A2(n4634), .ZN(n2285) );
  AOI21_X1 U2681 ( .B1(n3154), .B2(REG2_REG_7__SCAN_IN), .A(n3153), .ZN(n4291)
         );
  OR2_X1 U2682 ( .A1(n4262), .A2(n4290), .ZN(n2283) );
  NAND2_X1 U2683 ( .A1(n4689), .A2(n4267), .ZN(n4699) );
  NAND2_X1 U2684 ( .A1(n4701), .A2(n4296), .ZN(n4297) );
  NAND2_X1 U2685 ( .A1(n4712), .A2(REG2_REG_12__SCAN_IN), .ZN(n4710) );
  NAND2_X1 U2686 ( .A1(n4727), .A2(n2205), .ZN(n4273) );
  INV_X1 U2687 ( .A(n2578), .ZN(n2580) );
  AND2_X1 U2688 ( .A1(n2603), .A2(REG3_REG_21__SCAN_IN), .ZN(n2611) );
  AOI21_X1 U2689 ( .B1(n2233), .B2(n2236), .A(n2231), .ZN(n2230) );
  INV_X1 U2690 ( .A(n2237), .ZN(n2236) );
  OR2_X1 U2691 ( .A1(n2585), .A2(n2584), .ZN(n2596) );
  NOR2_X1 U2692 ( .A1(n2596), .A2(n4011), .ZN(n2603) );
  NAND2_X1 U2693 ( .A1(n4497), .A2(n2238), .ZN(n2232) );
  NOR2_X1 U2694 ( .A1(n2561), .A2(n2560), .ZN(n2572) );
  INV_X1 U2695 ( .A(n4138), .ZN(n4504) );
  NAND2_X1 U2696 ( .A1(n4497), .A2(n4504), .ZN(n4498) );
  NAND2_X1 U2697 ( .A1(n2558), .A2(n4187), .ZN(n2206) );
  NAND2_X1 U2698 ( .A1(n2720), .A2(n2198), .ZN(n2207) );
  NAND2_X1 U2699 ( .A1(n2720), .A2(n4088), .ZN(n3876) );
  OR2_X1 U2700 ( .A1(n2542), .A2(n2541), .ZN(n2548) );
  OR2_X1 U2701 ( .A1(n2548), .A2(n3458), .ZN(n2561) );
  NOR2_X1 U2702 ( .A1(n2241), .A2(n2354), .ZN(n2240) );
  NAND2_X1 U2703 ( .A1(n4183), .A2(n2246), .ZN(n3854) );
  NOR2_X1 U2704 ( .A1(n2511), .A2(n2510), .ZN(n2522) );
  OR2_X1 U2705 ( .A1(n3704), .A2(n4143), .ZN(n2356) );
  NAND2_X1 U2706 ( .A1(n3723), .A2(n4101), .ZN(n2713) );
  AND2_X1 U2707 ( .A1(n3770), .A2(n4102), .ZN(n4143) );
  NAND2_X1 U2708 ( .A1(n3592), .A2(n4089), .ZN(n2215) );
  AND2_X1 U2709 ( .A1(n2709), .A2(n4083), .ZN(n4142) );
  AND2_X1 U2710 ( .A1(n2448), .A2(REG3_REG_6__SCAN_IN), .ZN(n2457) );
  NAND2_X1 U2711 ( .A1(n3246), .A2(n4068), .ZN(n3245) );
  NAND2_X1 U2712 ( .A1(n2728), .A2(n2727), .ZN(n4514) );
  INV_X1 U2713 ( .A(n4068), .ZN(n3097) );
  OAI21_X1 U2714 ( .B1(n2402), .B2(n4826), .A(n2222), .ZN(n3255) );
  NAND2_X1 U2715 ( .A1(n2402), .A2(DATAI_0_), .ZN(n2222) );
  NAND2_X1 U2716 ( .A1(n2402), .A2(DATAI_31_), .ZN(n4656) );
  NOR2_X1 U2717 ( .A1(n2656), .A2(n4124), .ZN(n2218) );
  AND2_X1 U2718 ( .A1(n4347), .A2(n2217), .ZN(n2754) );
  AND2_X1 U2719 ( .A1(n2989), .A2(n4527), .ZN(n2217) );
  OR2_X1 U2720 ( .A1(n4383), .A2(n4362), .ZN(n4366) );
  OR2_X2 U2721 ( .A1(n4407), .A2(n4389), .ZN(n4383) );
  INV_X1 U2722 ( .A(n4402), .ZN(n4408) );
  AND2_X1 U2723 ( .A1(n4503), .A2(n4512), .ZN(n4501) );
  INV_X1 U2724 ( .A(n3952), .ZN(n4488) );
  NOR2_X1 U2725 ( .A1(n4587), .A2(n3926), .ZN(n4503) );
  OR2_X1 U2726 ( .A1(n3882), .A2(n3982), .ZN(n4587) );
  NAND2_X1 U2727 ( .A1(n3859), .A2(n4055), .ZN(n3882) );
  INV_X1 U2728 ( .A(n2882), .ZN(n4055) );
  NOR2_X1 U2729 ( .A1(n3902), .A2(n3845), .ZN(n3859) );
  NAND2_X1 U2730 ( .A1(n2247), .A2(n2245), .ZN(n3838) );
  AND2_X1 U2731 ( .A1(n2247), .A2(n2248), .ZN(n3839) );
  NAND2_X1 U2732 ( .A1(n2530), .A2(n2359), .ZN(n2247) );
  NAND2_X1 U2733 ( .A1(n2227), .A2(n3833), .ZN(n3845) );
  INV_X1 U2734 ( .A(n3733), .ZN(n3760) );
  AND2_X1 U2735 ( .A1(n3596), .A2(n3595), .ZN(n3663) );
  INV_X1 U2736 ( .A(n4658), .ZN(n4577) );
  AND3_X1 U2737 ( .A1(n2752), .A2(n2751), .A3(n2966), .ZN(n2759) );
  AND2_X1 U2738 ( .A1(n2172), .A2(n4807), .ZN(n3031) );
  INV_X1 U2739 ( .A(IR_REG_29__SCAN_IN), .ZN(n2379) );
  INV_X1 U2740 ( .A(IR_REG_19__SCAN_IN), .ZN(n2592) );
  INV_X1 U2741 ( .A(IR_REG_5__SCAN_IN), .ZN(n2365) );
  XNOR2_X1 U2742 ( .A(n2485), .B(IR_REG_9__SCAN_IN), .ZN(n4287) );
  OR3_X1 U2743 ( .A1(n2483), .A2(IR_REG_7__SCAN_IN), .A3(IR_REG_8__SCAN_IN), 
        .ZN(n2484) );
  INV_X1 U2744 ( .A(IR_REG_7__SCAN_IN), .ZN(n2470) );
  INV_X1 U2745 ( .A(IR_REG_3__SCAN_IN), .ZN(n2441) );
  INV_X1 U2746 ( .A(IR_REG_4__SCAN_IN), .ZN(n2442) );
  NAND2_X1 U2747 ( .A1(n2296), .A2(n2295), .ZN(n2410) );
  NAND2_X1 U2748 ( .A1(IR_REG_31__SCAN_IN), .A2(n3438), .ZN(n2295) );
  OAI21_X1 U2749 ( .B1(n2393), .B2(n2663), .A(IR_REG_2__SCAN_IN), .ZN(n2296)
         );
  NAND2_X1 U2750 ( .A1(n2342), .A2(n2341), .ZN(n2975) );
  AND2_X1 U2751 ( .A1(n2999), .A2(n2196), .ZN(n2341) );
  NAND2_X1 U2752 ( .A1(n4005), .A2(n4009), .ZN(n3960) );
  INV_X1 U2753 ( .A(n4557), .ZN(n4447) );
  INV_X1 U2754 ( .A(n3879), .ZN(n3982) );
  AOI21_X1 U2755 ( .B1(n2321), .B2(n2323), .A(n2894), .ZN(n2320) );
  AND2_X1 U2756 ( .A1(n2893), .A2(n2324), .ZN(n2323) );
  INV_X1 U2757 ( .A(n4542), .ZN(n4389) );
  INV_X1 U2758 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4000) );
  XNOR2_X1 U2759 ( .A(n2935), .B(n2791), .ZN(n3999) );
  INV_X1 U2760 ( .A(n3271), .ZN(n3193) );
  NAND2_X1 U2761 ( .A1(n2310), .A2(n2315), .ZN(n3691) );
  NAND2_X1 U2762 ( .A1(n3604), .A2(n2316), .ZN(n2310) );
  OAI21_X1 U2763 ( .B1(n3604), .B2(n2314), .A(n2311), .ZN(n3690) );
  AOI21_X1 U2764 ( .B1(n2988), .B2(n4658), .A(n4785), .ZN(n4056) );
  AND2_X1 U2765 ( .A1(n2988), .A2(n2971), .ZN(n3713) );
  AND2_X1 U2766 ( .A1(n2640), .A2(DATAI_20_), .ZN(n4466) );
  NAND2_X1 U2767 ( .A1(n2304), .A2(n2305), .ZN(n3830) );
  OR2_X1 U2768 ( .A1(n2864), .A2(n2173), .ZN(n2304) );
  NAND2_X1 U2769 ( .A1(n2338), .A2(n3957), .ZN(n4019) );
  NAND2_X1 U2770 ( .A1(n2852), .A2(n2854), .ZN(n2855) );
  INV_X1 U2771 ( .A(n3214), .ZN(n3222) );
  AND2_X1 U2772 ( .A1(n2648), .A2(n2634), .ZN(n4351) );
  INV_X1 U2773 ( .A(n4056), .ZN(n4041) );
  INV_X1 U2774 ( .A(n4349), .ZN(n4342) );
  AND2_X1 U2775 ( .A1(n2982), .A2(n4218), .ZN(n4059) );
  INV_X1 U2776 ( .A(n4022), .ZN(n4054) );
  NAND2_X1 U2777 ( .A1(n2646), .A2(n2645), .ZN(n4229) );
  OAI21_X1 U2778 ( .B1(n4385), .B2(n2630), .A(n2386), .ZN(n4363) );
  NAND4_X1 U2779 ( .A1(n2440), .A2(n2439), .A3(n2438), .A4(n2437), .ZN(n4233)
         );
  NAND3_X1 U2780 ( .A1(n2418), .A2(n2417), .A3(n2416), .ZN(n3229) );
  OR2_X1 U2781 ( .A1(n2404), .A2(n2414), .ZN(n2417) );
  NOR2_X1 U2782 ( .A1(n2361), .A2(n2180), .ZN(n2416) );
  OR2_X1 U2783 ( .A1(n2404), .A2(n2424), .ZN(n2425) );
  OR2_X1 U2784 ( .A1(n2404), .A2(n3049), .ZN(n2405) );
  OR2_X1 U2785 ( .A1(n2172), .A2(n3026), .ZN(n4235) );
  OR2_X1 U2786 ( .A1(n2404), .A2(n4861), .ZN(n2391) );
  NAND2_X1 U2787 ( .A1(n3059), .A2(n3066), .ZN(n2284) );
  AOI22_X1 U2788 ( .A1(n3067), .A2(REG2_REG_4__SCAN_IN), .B1(n3066), .B2(n3065), .ZN(n3069) );
  INV_X1 U2789 ( .A(n2291), .ZN(n3075) );
  XNOR2_X1 U2790 ( .A(n2289), .B(n2288), .ZN(n3085) );
  INV_X1 U2791 ( .A(n3155), .ZN(n3157) );
  AND2_X1 U2792 ( .A1(n2289), .A2(n4634), .ZN(n2287) );
  NAND2_X1 U2793 ( .A1(n4691), .A2(n4295), .ZN(n4702) );
  NAND2_X1 U2794 ( .A1(n4716), .A2(n4270), .ZN(n4728) );
  NAND2_X1 U2795 ( .A1(n4728), .A2(n4729), .ZN(n4727) );
  XNOR2_X1 U2796 ( .A(n4273), .B(n4816), .ZN(n4739) );
  NOR2_X1 U2797 ( .A1(n4301), .A2(n4733), .ZN(n4744) );
  NOR2_X1 U2798 ( .A1(n4759), .A2(n4278), .ZN(n4771) );
  NAND2_X1 U2799 ( .A1(n4754), .A2(n4305), .ZN(n4763) );
  NAND2_X1 U2800 ( .A1(n2252), .A2(n2249), .ZN(n4321) );
  INV_X1 U2801 ( .A(n2251), .ZN(n2249) );
  NAND2_X1 U2802 ( .A1(n2632), .A2(n2355), .ZN(n4338) );
  OR2_X1 U2803 ( .A1(n2633), .A2(n2625), .ZN(n4370) );
  NAND2_X1 U2804 ( .A1(n2257), .A2(n2256), .ZN(n4375) );
  INV_X1 U2805 ( .A(n2260), .ZN(n2256) );
  NOR2_X1 U2806 ( .A1(n4416), .A2(n2353), .ZN(n4394) );
  OAI21_X1 U2807 ( .B1(n2530), .B2(n2244), .A(n2242), .ZN(n3853) );
  INV_X1 U2808 ( .A(n3906), .ZN(n3902) );
  NAND2_X1 U2809 ( .A1(n4848), .A2(n2465), .ZN(n3644) );
  INV_X1 U2810 ( .A(n3229), .ZN(n2421) );
  INV_X1 U2811 ( .A(n4648), .ZN(n4516) );
  INV_X1 U2812 ( .A(n4420), .ZN(n4785) );
  AND2_X2 U2813 ( .A1(n2759), .A2(n2967), .ZN(n4867) );
  INV_X1 U2814 ( .A(n4867), .ZN(n4865) );
  INV_X1 U2815 ( .A(n2209), .ZN(n2208) );
  OAI21_X1 U2816 ( .B1(n2766), .B2(n4590), .A(n2764), .ZN(n2209) );
  XNOR2_X1 U2817 ( .A(n2668), .B(n2374), .ZN(n3027) );
  NAND2_X1 U2818 ( .A1(n3025), .A2(n3031), .ZN(n4806) );
  XNOR2_X1 U2819 ( .A(n2731), .B(IR_REG_28__SCAN_IN), .ZN(n4654) );
  NAND2_X1 U2820 ( .A1(n2671), .A2(IR_REG_31__SCAN_IN), .ZN(n2672) );
  INV_X1 U2821 ( .A(n4299), .ZN(n4818) );
  INV_X1 U2822 ( .A(n4285), .ZN(n4820) );
  XNOR2_X1 U2823 ( .A(n2444), .B(IR_REG_5__SCAN_IN), .ZN(n4635) );
  AOI21_X1 U2824 ( .B1(n2300), .B2(n2299), .A(n2297), .ZN(n4310) );
  NAND2_X1 U2825 ( .A1(n2298), .A2(n4309), .ZN(n2297) );
  AOI21_X1 U2826 ( .B1(n2219), .B2(n4517), .A(n2350), .ZN(n2745) );
  OR2_X1 U2827 ( .A1(n4316), .A2(n4585), .ZN(n2756) );
  NOR2_X1 U2828 ( .A1(n3787), .A2(n3788), .ZN(n2173) );
  AND2_X1 U2829 ( .A1(n2305), .A2(n2303), .ZN(n2174) );
  NOR2_X1 U2830 ( .A1(n2622), .A2(n2192), .ZN(n2175) );
  AND2_X1 U2831 ( .A1(n2401), .A2(n2399), .ZN(n2176) );
  OR2_X2 U2832 ( .A1(n2345), .A2(n2189), .ZN(n2177) );
  NAND2_X1 U2833 ( .A1(n4472), .A2(n2595), .ZN(n2178) );
  OR2_X1 U2834 ( .A1(n2244), .A2(n2195), .ZN(n2179) );
  AND2_X1 U2835 ( .A1(n2640), .A2(DATAI_28_), .ZN(n2656) );
  INV_X1 U2836 ( .A(n4634), .ZN(n2288) );
  OR2_X1 U2837 ( .A1(n3023), .A2(n2381), .ZN(n2404) );
  NAND3_X1 U2838 ( .A1(n2679), .A2(n2678), .A3(n3015), .ZN(n2778) );
  NAND2_X1 U2839 ( .A1(n2397), .A2(n3256), .ZN(n2706) );
  AND2_X1 U2840 ( .A1(n2170), .A2(REG2_REG_4__SCAN_IN), .ZN(n2180) );
  AND2_X1 U2841 ( .A1(n3665), .A2(n3618), .ZN(n2181) );
  AND4_X1 U2842 ( .A1(n2372), .A2(n2371), .A3(n2370), .A4(n2554), .ZN(n2182)
         );
  AND2_X1 U2843 ( .A1(n4232), .A2(n3794), .ZN(n2183) );
  XNOR2_X1 U2844 ( .A(n2380), .B(n2379), .ZN(n2381) );
  OR2_X1 U2845 ( .A1(n3787), .A2(n2307), .ZN(n2184) );
  OR2_X1 U2846 ( .A1(n2687), .A2(IR_REG_21__SCAN_IN), .ZN(n2185) );
  AND3_X1 U2847 ( .A1(n2368), .A2(n2369), .A3(n2333), .ZN(n2186) );
  AND2_X1 U2848 ( .A1(n3595), .A2(n3668), .ZN(n2187) );
  OR2_X1 U2849 ( .A1(n4255), .A2(n3040), .ZN(n2188) );
  OR2_X1 U2850 ( .A1(IR_REG_27__SCAN_IN), .A2(IR_REG_28__SCAN_IN), .ZN(n2189)
         );
  NAND2_X1 U2851 ( .A1(n3715), .A2(n3716), .ZN(n2190) );
  AND2_X1 U2852 ( .A1(n2398), .A2(n2400), .ZN(n2191) );
  NOR2_X1 U2853 ( .A1(n4425), .A2(n2353), .ZN(n2192) );
  OR2_X1 U2854 ( .A1(n3695), .A2(n3678), .ZN(n2193) );
  INV_X1 U2855 ( .A(n4146), .ZN(n2246) );
  NAND2_X1 U2856 ( .A1(n4509), .A2(n3952), .ZN(n2194) );
  INV_X1 U2857 ( .A(IR_REG_25__SCAN_IN), .ZN(n2374) );
  NOR2_X1 U2858 ( .A1(n2537), .A2(IR_REG_14__SCAN_IN), .ZN(n2568) );
  AND2_X1 U2859 ( .A1(n4231), .A2(n2882), .ZN(n2195) );
  NAND2_X1 U2860 ( .A1(n2864), .A2(n3751), .ZN(n3786) );
  NAND2_X1 U2861 ( .A1(n2232), .A2(n2237), .ZN(n4452) );
  NAND2_X1 U2862 ( .A1(n2327), .A2(n2328), .ZN(n3946) );
  INV_X1 U2863 ( .A(n2239), .ZN(n3874) );
  OR2_X1 U2864 ( .A1(n2952), .A2(n2951), .ZN(n2196) );
  NAND2_X1 U2865 ( .A1(n2367), .A2(n2366), .ZN(n2494) );
  OR2_X1 U2866 ( .A1(n4346), .A2(n4527), .ZN(n2197) );
  AND2_X1 U2867 ( .A1(n4187), .A2(n4088), .ZN(n2198) );
  INV_X1 U2868 ( .A(n2228), .ZN(n4565) );
  NOR2_X1 U2869 ( .A1(n4490), .A2(n4466), .ZN(n2228) );
  NOR2_X1 U2870 ( .A1(n4058), .A2(n3902), .ZN(n2199) );
  NOR2_X1 U2871 ( .A1(n4232), .A2(n3794), .ZN(n2200) );
  INV_X1 U2872 ( .A(IR_REG_10__SCAN_IN), .ZN(n2333) );
  NAND2_X1 U2873 ( .A1(n2944), .A2(n3968), .ZN(n2201) );
  NAND2_X1 U2874 ( .A1(n2778), .A2(n2777), .ZN(n2926) );
  INV_X4 U2875 ( .A(n2926), .ZN(n2789) );
  XNOR2_X1 U2876 ( .A(n2672), .B(IR_REG_26__SCAN_IN), .ZN(n2678) );
  NAND2_X1 U2877 ( .A1(n2356), .A2(n2509), .ZN(n3775) );
  OR2_X1 U2878 ( .A1(n2662), .A2(n2663), .ZN(n2680) );
  OR2_X1 U2879 ( .A1(n2740), .A2(n4420), .ZN(n2202) );
  INV_X1 U2880 ( .A(n2358), .ZN(n2248) );
  NAND2_X1 U2881 ( .A1(n2640), .A2(DATAI_27_), .ZN(n4527) );
  AND2_X2 U2882 ( .A1(n2759), .A2(n2758), .ZN(n4860) );
  INV_X1 U2883 ( .A(n4860), .ZN(n4858) );
  NAND4_X1 U2884 ( .A1(n2428), .A2(n2427), .A3(n2426), .A4(n2425), .ZN(n4234)
         );
  INV_X1 U2885 ( .A(n4276), .ZN(n4812) );
  INV_X1 U2886 ( .A(n3751), .ZN(n2307) );
  AND2_X1 U2887 ( .A1(n3030), .A2(n3029), .ZN(n2203) );
  AND2_X1 U2888 ( .A1(n2871), .A2(n2870), .ZN(n2204) );
  OR2_X1 U2889 ( .A1(n4818), .A2(n4271), .ZN(n2205) );
  INV_X1 U2890 ( .A(n2656), .ZN(n2989) );
  INV_X1 U2891 ( .A(n4709), .ZN(n2286) );
  INV_X1 U2892 ( .A(IR_REG_13__SCAN_IN), .ZN(n2369) );
  NAND2_X1 U2893 ( .A1(n2765), .A2(n2208), .ZN(n2773) );
  OAI21_X1 U2894 ( .B1(n2747), .B2(n4064), .A(n4123), .ZN(n2213) );
  INV_X1 U2895 ( .A(n3246), .ZN(n2705) );
  AND2_X2 U2896 ( .A1(n2706), .A2(n4066), .ZN(n3246) );
  OAI21_X2 U2897 ( .B1(n3649), .B2(n4099), .A(n4085), .ZN(n3723) );
  OAI21_X2 U2898 ( .B1(n3771), .B2(n2715), .A(n4105), .ZN(n4183) );
  AND2_X2 U2899 ( .A1(n4347), .A2(n4527), .ZN(n4327) );
  NAND3_X1 U2900 ( .A1(n2220), .A2(n2765), .A3(n2202), .ZN(n2219) );
  NOR2_X4 U2901 ( .A1(n2360), .A2(n3657), .ZN(n3727) );
  NOR2_X4 U2902 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2393)
         );
  AND4_X2 U2903 ( .A1(n2226), .A2(n2225), .A3(n2224), .A4(n2365), .ZN(n2367)
         );
  NAND3_X2 U2905 ( .A1(n2367), .A2(n2366), .A3(n2186), .ZN(n2537) );
  NOR3_X4 U2906 ( .A1(n4490), .A2(n4447), .A3(n4466), .ZN(n4439) );
  AND2_X2 U2907 ( .A1(n4439), .A2(n4417), .ZN(n4419) );
  NAND2_X1 U2908 ( .A1(n2281), .A2(n2280), .ZN(n2279) );
  OAI21_X1 U2909 ( .B1(n2729), .B2(n2387), .A(IR_REG_27__SCAN_IN), .ZN(n2282)
         );
  INV_X1 U2910 ( .A(n2366), .ZN(n2409) );
  NAND2_X1 U2911 ( .A1(n4497), .A2(n2233), .ZN(n2229) );
  NAND2_X1 U2912 ( .A1(n2229), .A2(n2230), .ZN(n4434) );
  OAI21_X1 U2913 ( .B1(n2530), .B2(n2179), .A(n2240), .ZN(n2239) );
  NAND2_X1 U2914 ( .A1(n2252), .A2(n2250), .ZN(n2255) );
  INV_X1 U2915 ( .A(n2259), .ZN(n2257) );
  NOR2_X1 U2916 ( .A1(n2259), .A2(n2258), .ZN(n2623) );
  NAND4_X1 U2917 ( .A1(n2268), .A2(n2266), .A3(n2265), .A4(n2193), .ZN(n2475)
         );
  NAND2_X1 U2918 ( .A1(n4142), .A2(n2465), .ZN(n2265) );
  NAND2_X1 U2919 ( .A1(n2269), .A2(n2270), .ZN(n2268) );
  INV_X1 U2920 ( .A(n3591), .ZN(n2269) );
  OAI21_X1 U2921 ( .B1(n3704), .B2(n2277), .A(n2275), .ZN(n3811) );
  NAND2_X2 U2922 ( .A1(n2282), .A2(n2279), .ZN(n2402) );
  MUX2_X1 U2923 ( .A(n2392), .B(IR_REG_31__SCAN_IN), .S(n3407), .Z(n2395) );
  NOR2_X2 U2924 ( .A1(n3080), .A2(n2450), .ZN(n3089) );
  XNOR2_X2 U2925 ( .A(n3088), .B(n2288), .ZN(n3080) );
  NAND2_X1 U2926 ( .A1(n2864), .A2(n2174), .ZN(n2301) );
  NAND2_X1 U2927 ( .A1(n2301), .A2(n2302), .ZN(n3895) );
  NAND2_X1 U2928 ( .A1(n3604), .A2(n2311), .ZN(n2308) );
  NAND2_X1 U2929 ( .A1(n2308), .A2(n2309), .ZN(n3714) );
  NAND2_X1 U2930 ( .A1(n3939), .A2(n2934), .ZN(n2937) );
  NAND2_X1 U2931 ( .A1(n2892), .A2(n2321), .ZN(n2319) );
  NAND2_X1 U2932 ( .A1(n2319), .A2(n2320), .ZN(n3986) );
  NAND2_X1 U2933 ( .A1(n4031), .A2(n2329), .ZN(n2327) );
  NAND2_X1 U2934 ( .A1(n4028), .A2(n4029), .ZN(n2328) );
  NAND3_X1 U2935 ( .A1(n2367), .A2(n2366), .A3(n2333), .ZN(n2335) );
  INV_X1 U2936 ( .A(n2335), .ZN(n2496) );
  NAND2_X1 U2937 ( .A1(n2338), .A2(n2336), .ZN(n4017) );
  AND2_X1 U2938 ( .A1(n2344), .A2(n2201), .ZN(n4038) );
  INV_X1 U2939 ( .A(n2975), .ZN(n3006) );
  NOR2_X1 U2940 ( .A1(n2687), .A2(n2347), .ZN(n2662) );
  NOR2_X2 U2941 ( .A1(n2687), .A2(n2177), .ZN(n2378) );
  AOI21_X2 U2942 ( .B1(n4635), .B2(REG1_REG_5__SCAN_IN), .A(n3078), .ZN(n3088)
         );
  OAI21_X1 U2943 ( .B1(n3007), .B2(n3006), .A(n3005), .ZN(U3211) );
  MUX2_X2 U2944 ( .A(REG0_REG_28__SCAN_IN), .B(n2760), .S(n4860), .Z(n2761) );
  MUX2_X2 U2945 ( .A(REG1_REG_28__SCAN_IN), .B(n2760), .S(n4867), .Z(n2753) );
  AND2_X2 U2946 ( .A1(n3023), .A2(n2382), .ZN(n2422) );
  BUF_X8 U2947 ( .A(n2402), .Z(n2640) );
  AND2_X1 U2948 ( .A1(n4517), .A2(n2739), .ZN(n4776) );
  NOR2_X1 U2949 ( .A1(n4867), .A2(n2767), .ZN(n2349) );
  XNOR2_X1 U2950 ( .A(n2820), .B(n2821), .ZN(n3189) );
  OR2_X1 U2951 ( .A1(n2744), .A2(n2743), .ZN(n2350) );
  AND2_X1 U2952 ( .A1(n2974), .A2(n2973), .ZN(n2351) );
  AND2_X1 U2953 ( .A1(n2842), .A2(n2841), .ZN(n2352) );
  AND2_X1 U2954 ( .A1(n4403), .A2(n4427), .ZN(n2353) );
  NOR2_X1 U2955 ( .A1(n4231), .A2(n2882), .ZN(n2354) );
  OR2_X1 U2956 ( .A1(n4381), .A2(n4367), .ZN(n2355) );
  INV_X1 U2957 ( .A(n4367), .ZN(n4362) );
  NAND2_X1 U2958 ( .A1(n2640), .A2(DATAI_25_), .ZN(n4367) );
  AND2_X1 U2959 ( .A1(n2996), .A2(n2995), .ZN(n2357) );
  INV_X1 U2960 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2771) );
  INV_X1 U2961 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2560) );
  INV_X1 U2962 ( .A(n4255), .ZN(n2412) );
  AND2_X1 U2963 ( .A1(n4184), .A2(n4187), .ZN(n4150) );
  INV_X1 U2964 ( .A(n4150), .ZN(n2558) );
  OAI21_X1 U2965 ( .B1(n4370), .B2(n2630), .A(n2629), .ZN(n4343) );
  AND2_X1 U2966 ( .A1(n3843), .A2(n3817), .ZN(n2358) );
  OR2_X1 U2967 ( .A1(n3843), .A2(n3817), .ZN(n2359) );
  INV_X1 U2968 ( .A(n4829), .ZN(n2782) );
  AND2_X1 U2969 ( .A1(n2422), .A2(n3285), .ZN(n2361) );
  OR2_X1 U2970 ( .A1(n2774), .A2(n4628), .ZN(n2362) );
  INV_X1 U2971 ( .A(n3199), .ZN(n2430) );
  INV_X1 U2972 ( .A(IR_REG_2__SCAN_IN), .ZN(n3438) );
  OR2_X1 U2973 ( .A1(n2924), .A2(n2923), .ZN(n2925) );
  INV_X1 U2974 ( .A(n3275), .ZN(n2432) );
  INV_X1 U2975 ( .A(n3938), .ZN(n2930) );
  INV_X1 U2976 ( .A(n2853), .ZN(n2854) );
  INV_X1 U2977 ( .A(IR_REG_17__SCAN_IN), .ZN(n2579) );
  INV_X1 U2978 ( .A(n4822), .ZN(n4293) );
  INV_X1 U2979 ( .A(n3247), .ZN(n3249) );
  AND2_X1 U2980 ( .A1(n2972), .A2(n3713), .ZN(n2973) );
  INV_X1 U2981 ( .A(REG3_REG_16__SCAN_IN), .ZN(n3458) );
  OR3_X1 U2982 ( .A1(n2648), .A2(n2992), .A3(n3001), .ZN(n2740) );
  NAND2_X1 U2983 ( .A1(n2580), .A2(n2579), .ZN(n2591) );
  AND2_X1 U2984 ( .A1(n2649), .A2(n2740), .ZN(n4314) );
  NAND2_X1 U2985 ( .A1(n2611), .A2(REG3_REG_22__SCAN_IN), .ZN(n2616) );
  AND2_X1 U2986 ( .A1(n4479), .A2(n4477), .ZN(n4138) );
  AND2_X1 U2987 ( .A1(n2522), .A2(REG3_REG_13__SCAN_IN), .ZN(n2531) );
  INV_X1 U2988 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2767) );
  INV_X1 U2989 ( .A(n4578), .ZN(n4506) );
  INV_X1 U2990 ( .A(n3025), .ZN(n2700) );
  NAND2_X1 U2991 ( .A1(n2531), .A2(REG3_REG_14__SCAN_IN), .ZN(n2542) );
  OR2_X1 U2992 ( .A1(n2616), .A2(n3941), .ZN(n2618) );
  NAND2_X1 U2993 ( .A1(n2457), .A2(REG3_REG_7__SCAN_IN), .ZN(n2476) );
  AND2_X1 U2994 ( .A1(n2434), .A2(REG3_REG_5__SCAN_IN), .ZN(n2448) );
  INV_X1 U2995 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4011) );
  OR2_X1 U2996 ( .A1(n2501), .A2(n2500), .ZN(n2511) );
  OAI21_X1 U2997 ( .B1(n3119), .B2(n3120), .A(n2803), .ZN(n3124) );
  NAND2_X1 U2998 ( .A1(n2633), .A2(REG3_REG_26__SCAN_IN), .ZN(n2648) );
  AND2_X1 U2999 ( .A1(n2624), .A2(REG3_REG_25__SCAN_IN), .ZN(n2633) );
  INV_X1 U3000 ( .A(n4332), .ZN(n4528) );
  INV_X1 U3001 ( .A(n4363), .ZN(n4406) );
  AND2_X1 U3002 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2434) );
  INV_X1 U3003 ( .A(n4776), .ZN(n4493) );
  NAND2_X1 U3004 ( .A1(n2640), .A2(DATAI_22_), .ZN(n4417) );
  INV_X1 U3005 ( .A(n3618), .ZN(n3595) );
  AND2_X1 U3006 ( .A1(n3114), .A2(n2983), .ZN(n2752) );
  OR2_X1 U3007 ( .A1(n3031), .A2(n4221), .ZN(n3041) );
  AND2_X1 U3008 ( .A1(n2640), .A2(DATAI_23_), .ZN(n4402) );
  AOI21_X1 U3009 ( .B1(n3986), .B2(n3988), .A(n3987), .ZN(n4031) );
  INV_X1 U3010 ( .A(n4021), .ZN(n4053) );
  INV_X1 U3011 ( .A(n2422), .ZN(n2630) );
  AND2_X1 U3012 ( .A1(n3042), .A2(n3041), .ZN(n4675) );
  INV_X1 U3013 ( .A(n4177), .ZN(n4525) );
  INV_X1 U3014 ( .A(n4482), .ZN(n4508) );
  AND2_X1 U3015 ( .A1(n2676), .A2(n2675), .ZN(n2967) );
  NAND2_X1 U3016 ( .A1(n4858), .A2(n2771), .ZN(n2772) );
  INV_X1 U3017 ( .A(n4590), .ZN(n4856) );
  INV_X1 U3018 ( .A(n2967), .ZN(n2758) );
  OAI21_X1 U3019 ( .B1(n2680), .B2(n2682), .A(n2681), .ZN(n3030) );
  AND2_X1 U3020 ( .A1(n2540), .A2(n2539), .ZN(n4272) );
  AND2_X1 U3021 ( .A1(n3032), .A2(n3041), .ZN(n4768) );
  INV_X1 U3022 ( .A(n3713), .ZN(n4062) );
  INV_X1 U3023 ( .A(n4325), .ZN(n4228) );
  OAI211_X1 U3024 ( .C1(n4441), .C2(n2630), .A(n2608), .B(n2607), .ZN(n4428)
         );
  NAND2_X1 U3025 ( .A1(n4675), .A2(n4654), .ZN(n4775) );
  INV_X1 U3026 ( .A(n4711), .ZN(n4762) );
  NAND2_X1 U3027 ( .A1(n4517), .A2(n2704), .ZN(n4521) );
  NAND2_X1 U3028 ( .A1(n4867), .A2(n4829), .ZN(n4585) );
  OR2_X1 U3029 ( .A1(n4316), .A2(n4628), .ZN(n2762) );
  NAND2_X1 U3030 ( .A1(n4860), .A2(n4829), .ZN(n4628) );
  INV_X1 U3031 ( .A(n4806), .ZN(n4805) );
  AND2_X1 U3032 ( .A1(n3030), .A2(STATE_REG_SCAN_IN), .ZN(n4807) );
  INV_X1 U3033 ( .A(n4272), .ZN(n4816) );
  OAI21_X1 U3034 ( .B1(n2766), .B2(n4521), .A(n2745), .ZN(U3354) );
  NAND2_X1 U3035 ( .A1(n2770), .A2(n2769), .ZN(U3547) );
  NAND2_X1 U3036 ( .A1(REG3_REG_8__SCAN_IN), .A2(REG3_REG_9__SCAN_IN), .ZN(
        n2363) );
  NAND2_X1 U3037 ( .A1(n2487), .A2(REG3_REG_10__SCAN_IN), .ZN(n2501) );
  NAND2_X1 U3038 ( .A1(n2572), .A2(REG3_REG_18__SCAN_IN), .ZN(n2585) );
  AND2_X1 U3039 ( .A1(n2618), .A2(n4000), .ZN(n2364) );
  OR2_X1 U3040 ( .A1(n2364), .A2(n2624), .ZN(n4385) );
  NAND2_X1 U3041 ( .A1(n2378), .A2(n2379), .ZN(n3933) );
  XNOR2_X2 U3042 ( .A(n2377), .B(IR_REG_30__SCAN_IN), .ZN(n3023) );
  INV_X1 U3043 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4547) );
  NAND2_X1 U3044 ( .A1(n2423), .A2(REG2_REG_24__SCAN_IN), .ZN(n2384) );
  INV_X1 U3045 ( .A(n2381), .ZN(n2382) );
  NOR2_X2 U3046 ( .A1(n3023), .A2(n2382), .ZN(n2413) );
  NAND2_X1 U3047 ( .A1(n2413), .A2(REG0_REG_24__SCAN_IN), .ZN(n2383) );
  OAI211_X1 U3048 ( .C1(n3146), .C2(n4547), .A(n2384), .B(n2383), .ZN(n2385)
         );
  INV_X1 U3049 ( .A(n2385), .ZN(n2386) );
  NAND2_X1 U3050 ( .A1(n2423), .A2(REG2_REG_1__SCAN_IN), .ZN(n2390) );
  NAND2_X1 U3051 ( .A1(n2413), .A2(REG0_REG_1__SCAN_IN), .ZN(n2388) );
  NAND2_X1 U3052 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2392)
         );
  INV_X1 U3053 ( .A(n2393), .ZN(n2394) );
  NAND2_X1 U3054 ( .A1(n2395), .A2(n2394), .ZN(n3047) );
  INV_X1 U3055 ( .A(DATAI_1_), .ZN(n2396) );
  MUX2_X1 U3056 ( .A(n3047), .B(n2396), .S(n2402), .Z(n2793) );
  INV_X1 U3057 ( .A(n2790), .ZN(n2397) );
  INV_X1 U3058 ( .A(n2793), .ZN(n3256) );
  NAND2_X1 U3059 ( .A1(n2422), .A2(REG3_REG_0__SCAN_IN), .ZN(n2401) );
  NAND2_X1 U3060 ( .A1(n2423), .A2(REG2_REG_0__SCAN_IN), .ZN(n2400) );
  NAND2_X1 U3061 ( .A1(n2413), .A2(REG0_REG_0__SCAN_IN), .ZN(n2399) );
  INV_X1 U3062 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2799) );
  AND2_X1 U3063 ( .A1(n3247), .A2(n3255), .ZN(n3244) );
  NAND2_X1 U3064 ( .A1(n2705), .A2(n3244), .ZN(n3243) );
  NAND2_X1 U3065 ( .A1(n2790), .A2(n3256), .ZN(n2403) );
  NAND2_X1 U3066 ( .A1(n2422), .A2(REG3_REG_2__SCAN_IN), .ZN(n2408) );
  NAND2_X1 U3067 ( .A1(n2413), .A2(REG0_REG_2__SCAN_IN), .ZN(n2407) );
  NAND2_X1 U3068 ( .A1(n2423), .A2(REG2_REG_2__SCAN_IN), .ZN(n2406) );
  INV_X1 U3069 ( .A(REG1_REG_2__SCAN_IN), .ZN(n3049) );
  NAND2_X1 U3070 ( .A1(n2410), .A2(n2409), .ZN(n4255) );
  INV_X1 U3071 ( .A(DATAI_2_), .ZN(n2411) );
  NAND2_X1 U3072 ( .A1(n4236), .A2(n3214), .ZN(n4072) );
  NAND2_X1 U3073 ( .A1(n4069), .A2(n4072), .ZN(n4145) );
  NAND2_X1 U3074 ( .A1(n3211), .A2(n4145), .ZN(n3198) );
  NAND2_X1 U3075 ( .A1(n2413), .A2(REG0_REG_4__SCAN_IN), .ZN(n2418) );
  INV_X1 U3076 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2414) );
  NOR2_X1 U3077 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2415) );
  NOR2_X1 U3078 ( .A1(n2434), .A2(n2415), .ZN(n3285) );
  NAND2_X1 U3079 ( .A1(n2409), .A2(IR_REG_31__SCAN_IN), .ZN(n2429) );
  NAND2_X1 U3080 ( .A1(n2429), .A2(n2441), .ZN(n2419) );
  NAND2_X1 U3081 ( .A1(n2419), .A2(IR_REG_31__SCAN_IN), .ZN(n2420) );
  XNOR2_X1 U3082 ( .A(n2420), .B(n2442), .ZN(n3176) );
  INV_X1 U3083 ( .A(DATAI_4_), .ZN(n3008) );
  MUX2_X1 U3084 ( .A(n3176), .B(n3008), .S(n2640), .Z(n3271) );
  NAND2_X1 U3085 ( .A1(n2421), .A2(n3193), .ZN(n4075) );
  NAND2_X1 U3086 ( .A1(n3229), .A2(n3271), .ZN(n4079) );
  NAND2_X1 U3087 ( .A1(n4075), .A2(n4079), .ZN(n3267) );
  INV_X1 U3088 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3044) );
  NAND2_X1 U3089 ( .A1(n2422), .A2(n3044), .ZN(n2428) );
  NAND2_X1 U3090 ( .A1(n2170), .A2(REG2_REG_3__SCAN_IN), .ZN(n2426) );
  INV_X1 U3091 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2424) );
  INV_X1 U3092 ( .A(n4234), .ZN(n2431) );
  XNOR2_X1 U3093 ( .A(n2429), .B(IR_REG_3__SCAN_IN), .ZN(n3062) );
  MUX2_X1 U3094 ( .A(n3062), .B(DATAI_3_), .S(n2640), .Z(n3209) );
  OR2_X1 U3095 ( .A1(n4236), .A2(n3222), .ZN(n3199) );
  NAND3_X1 U3096 ( .A1(n3198), .A2(n3267), .A3(n3274), .ZN(n3273) );
  NAND2_X1 U3097 ( .A1(n4234), .A2(n3209), .ZN(n3275) );
  NAND2_X1 U3098 ( .A1(n3267), .A2(n2432), .ZN(n3272) );
  NAND2_X1 U3099 ( .A1(n3229), .A2(n3193), .ZN(n2433) );
  NAND3_X1 U3100 ( .A1(n3273), .A2(n3272), .A3(n2433), .ZN(n3296) );
  NAND2_X1 U3101 ( .A1(n2732), .A2(REG0_REG_5__SCAN_IN), .ZN(n2440) );
  NOR2_X1 U3102 ( .A1(n2434), .A2(REG3_REG_5__SCAN_IN), .ZN(n2435) );
  NOR2_X1 U3103 ( .A1(n2448), .A2(n2435), .ZN(n3627) );
  NAND2_X1 U3104 ( .A1(n2422), .A2(n3627), .ZN(n2439) );
  NAND2_X1 U3105 ( .A1(n2170), .A2(REG2_REG_5__SCAN_IN), .ZN(n2438) );
  INV_X1 U3106 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2436) );
  OR2_X1 U3107 ( .A1(n2404), .A2(n2436), .ZN(n2437) );
  NAND2_X1 U3108 ( .A1(n2442), .A2(n2441), .ZN(n2443) );
  OR2_X1 U3109 ( .A1(n2409), .A2(n2443), .ZN(n2455) );
  NAND2_X1 U3110 ( .A1(n2455), .A2(IR_REG_31__SCAN_IN), .ZN(n2444) );
  MUX2_X1 U3111 ( .A(n4635), .B(DATAI_5_), .S(n2640), .Z(n3631) );
  OR2_X1 U3112 ( .A1(n4233), .A2(n3631), .ZN(n2445) );
  NAND2_X1 U3113 ( .A1(n3296), .A2(n2445), .ZN(n2447) );
  NAND2_X1 U3114 ( .A1(n4233), .A2(n3631), .ZN(n2446) );
  NAND2_X1 U3115 ( .A1(n2447), .A2(n2446), .ZN(n3591) );
  NAND2_X1 U3116 ( .A1(n2170), .A2(REG2_REG_6__SCAN_IN), .ZN(n2454) );
  NOR2_X1 U3117 ( .A1(n2448), .A2(REG3_REG_6__SCAN_IN), .ZN(n2449) );
  NOR2_X1 U3118 ( .A1(n2457), .A2(n2449), .ZN(n3614) );
  NAND2_X1 U3119 ( .A1(n2422), .A2(n3614), .ZN(n2453) );
  NAND2_X1 U3120 ( .A1(n2732), .A2(REG0_REG_6__SCAN_IN), .ZN(n2452) );
  INV_X1 U3121 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2450) );
  OR2_X1 U3122 ( .A1(n2404), .A2(n2450), .ZN(n2451) );
  NAND4_X1 U3123 ( .A1(n2454), .A2(n2453), .A3(n2452), .A4(n2451), .ZN(n3665)
         );
  NOR2_X1 U3124 ( .A1(n2455), .A2(IR_REG_5__SCAN_IN), .ZN(n2464) );
  OR2_X1 U3125 ( .A1(n2464), .A2(n2663), .ZN(n2456) );
  XNOR2_X1 U3126 ( .A(n2456), .B(IR_REG_6__SCAN_IN), .ZN(n4634) );
  MUX2_X1 U3127 ( .A(n4634), .B(DATAI_6_), .S(n2640), .Z(n3618) );
  NAND2_X1 U3128 ( .A1(n2170), .A2(REG2_REG_7__SCAN_IN), .ZN(n2462) );
  OAI21_X1 U3129 ( .B1(n2457), .B2(REG3_REG_7__SCAN_IN), .A(n2476), .ZN(n3671)
         );
  INV_X1 U3130 ( .A(n3671), .ZN(n2458) );
  NAND2_X1 U3131 ( .A1(n2422), .A2(n2458), .ZN(n2461) );
  NAND2_X1 U3132 ( .A1(n2732), .A2(REG0_REG_7__SCAN_IN), .ZN(n2460) );
  INV_X1 U3133 ( .A(REG1_REG_7__SCAN_IN), .ZN(n3156) );
  OR2_X1 U3134 ( .A1(n2404), .A2(n3156), .ZN(n2459) );
  NAND4_X1 U3135 ( .A1(n2462), .A2(n2461), .A3(n2460), .A4(n2459), .ZN(n3679)
         );
  INV_X1 U3136 ( .A(IR_REG_6__SCAN_IN), .ZN(n2463) );
  NAND2_X1 U3137 ( .A1(n2464), .A2(n2463), .ZN(n2483) );
  NAND2_X1 U3138 ( .A1(n2483), .A2(IR_REG_31__SCAN_IN), .ZN(n2471) );
  XNOR2_X1 U3139 ( .A(n2471), .B(n2470), .ZN(n3158) );
  INV_X1 U3140 ( .A(DATAI_7_), .ZN(n3460) );
  MUX2_X1 U3141 ( .A(n3158), .B(n3460), .S(n2640), .Z(n3668) );
  OR2_X1 U3142 ( .A1(n3679), .A2(n3668), .ZN(n2709) );
  NAND2_X1 U3143 ( .A1(n3679), .A2(n3668), .ZN(n4083) );
  INV_X1 U3144 ( .A(n3668), .ZN(n3314) );
  NAND2_X1 U3145 ( .A1(n3679), .A2(n3314), .ZN(n2465) );
  NAND2_X1 U3146 ( .A1(n2732), .A2(REG0_REG_8__SCAN_IN), .ZN(n2469) );
  XNOR2_X1 U3147 ( .A(n2476), .B(REG3_REG_8__SCAN_IN), .ZN(n3640) );
  NAND2_X1 U31480 ( .A1(n2422), .A2(n3640), .ZN(n2468) );
  NAND2_X1 U31490 ( .A1(n2170), .A2(REG2_REG_8__SCAN_IN), .ZN(n2467) );
  INV_X1 U3150 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4263) );
  OR2_X1 U3151 ( .A1(n3146), .A2(n4263), .ZN(n2466) );
  NAND4_X1 U3152 ( .A1(n2469), .A2(n2468), .A3(n2467), .A4(n2466), .ZN(n3695)
         );
  NAND2_X1 U3153 ( .A1(n2471), .A2(n2470), .ZN(n2472) );
  NAND2_X1 U3154 ( .A1(n2472), .A2(IR_REG_31__SCAN_IN), .ZN(n2473) );
  XNOR2_X1 U3155 ( .A(n2473), .B(IR_REG_8__SCAN_IN), .ZN(n4633) );
  MUX2_X1 U3156 ( .A(n4633), .B(DATAI_8_), .S(n2640), .Z(n3678) );
  NAND2_X1 U3157 ( .A1(n3695), .A2(n3678), .ZN(n2474) );
  NAND2_X1 U3158 ( .A1(n2475), .A2(n2474), .ZN(n3651) );
  INV_X1 U3159 ( .A(n2476), .ZN(n2477) );
  AOI21_X1 U3160 ( .B1(n2477), .B2(REG3_REG_8__SCAN_IN), .A(
        REG3_REG_9__SCAN_IN), .ZN(n2478) );
  OR2_X1 U3161 ( .A1(n2478), .A2(n2487), .ZN(n3654) );
  INV_X1 U3162 ( .A(n3654), .ZN(n3693) );
  NAND2_X1 U3163 ( .A1(n2422), .A2(n3693), .ZN(n2482) );
  NAND2_X1 U3164 ( .A1(n2732), .A2(REG0_REG_9__SCAN_IN), .ZN(n2481) );
  NAND2_X1 U3165 ( .A1(n2170), .A2(REG2_REG_9__SCAN_IN), .ZN(n2480) );
  INV_X1 U3166 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3744) );
  OR2_X1 U3167 ( .A1(n3146), .A2(n3744), .ZN(n2479) );
  NAND4_X1 U3168 ( .A1(n2482), .A2(n2481), .A3(n2480), .A4(n2479), .ZN(n3759)
         );
  NAND2_X1 U3169 ( .A1(n2484), .A2(IR_REG_31__SCAN_IN), .ZN(n2485) );
  MUX2_X1 U3170 ( .A(n4287), .B(DATAI_9_), .S(n2640), .Z(n3657) );
  AND2_X1 U3171 ( .A1(n3759), .A2(n3657), .ZN(n2486) );
  NAND2_X1 U3172 ( .A1(n2732), .A2(REG0_REG_10__SCAN_IN), .ZN(n2493) );
  OR2_X1 U3173 ( .A1(n2487), .A2(REG3_REG_10__SCAN_IN), .ZN(n2488) );
  AND2_X1 U3174 ( .A1(n2501), .A2(n2488), .ZN(n3730) );
  NAND2_X1 U3175 ( .A1(n2422), .A2(n3730), .ZN(n2492) );
  NAND2_X1 U3176 ( .A1(n2170), .A2(REG2_REG_10__SCAN_IN), .ZN(n2491) );
  INV_X1 U3177 ( .A(REG1_REG_10__SCAN_IN), .ZN(n2489) );
  OR2_X1 U3178 ( .A1(n3146), .A2(n2489), .ZN(n2490) );
  NAND4_X1 U3179 ( .A1(n2493), .A2(n2492), .A3(n2491), .A4(n2490), .ZN(n3801)
         );
  NAND2_X1 U3180 ( .A1(n2494), .A2(IR_REG_31__SCAN_IN), .ZN(n2495) );
  MUX2_X1 U3181 ( .A(IR_REG_31__SCAN_IN), .B(n2495), .S(IR_REG_10__SCAN_IN), 
        .Z(n2497) );
  NAND2_X1 U3182 ( .A1(n2497), .A2(n2335), .ZN(n4822) );
  MUX2_X1 U3183 ( .A(n4293), .B(DATAI_10_), .S(n2640), .Z(n3733) );
  NOR2_X1 U3184 ( .A1(n3801), .A2(n3733), .ZN(n2499) );
  NAND2_X1 U3185 ( .A1(n3801), .A2(n3733), .ZN(n2498) );
  OAI21_X1 U3186 ( .B1(n3726), .B2(n2499), .A(n2498), .ZN(n3704) );
  NAND2_X1 U3187 ( .A1(n2732), .A2(REG0_REG_11__SCAN_IN), .ZN(n2507) );
  NAND2_X1 U3188 ( .A1(n2501), .A2(n2500), .ZN(n2502) );
  AND2_X1 U3189 ( .A1(n2511), .A2(n2502), .ZN(n3754) );
  NAND2_X1 U3190 ( .A1(n2422), .A2(n3754), .ZN(n2506) );
  NAND2_X1 U3191 ( .A1(n2170), .A2(REG2_REG_11__SCAN_IN), .ZN(n2505) );
  INV_X1 U3192 ( .A(REG1_REG_11__SCAN_IN), .ZN(n2503) );
  OR2_X1 U3193 ( .A1(n3146), .A2(n2503), .ZN(n2504) );
  NAND4_X1 U3194 ( .A1(n2507), .A2(n2506), .A3(n2505), .A4(n2504), .ZN(n3724)
         );
  OR2_X1 U3195 ( .A1(n2496), .A2(n2663), .ZN(n2519) );
  XNOR2_X1 U3196 ( .A(n2519), .B(IR_REG_11__SCAN_IN), .ZN(n4285) );
  INV_X1 U3197 ( .A(DATAI_11_), .ZN(n2508) );
  MUX2_X1 U3198 ( .A(n4820), .B(n2508), .S(n2640), .Z(n3799) );
  OR2_X1 U3199 ( .A1(n3724), .A2(n3799), .ZN(n3770) );
  NAND2_X1 U3200 ( .A1(n3724), .A2(n3799), .ZN(n4102) );
  INV_X1 U3201 ( .A(n3799), .ZN(n3709) );
  OR2_X1 U3202 ( .A1(n3724), .A2(n3709), .ZN(n2509) );
  NAND2_X1 U3203 ( .A1(n2170), .A2(REG2_REG_12__SCAN_IN), .ZN(n2517) );
  AND2_X1 U3204 ( .A1(n2511), .A2(n2510), .ZN(n2512) );
  NOR2_X1 U3205 ( .A1(n2522), .A2(n2512), .ZN(n3791) );
  NAND2_X1 U3206 ( .A1(n2422), .A2(n3791), .ZN(n2516) );
  NAND2_X1 U3207 ( .A1(n2732), .A2(REG0_REG_12__SCAN_IN), .ZN(n2515) );
  INV_X1 U3208 ( .A(REG1_REG_12__SCAN_IN), .ZN(n2513) );
  OR2_X1 U3209 ( .A1(n3146), .A2(n2513), .ZN(n2514) );
  NAND4_X1 U32100 ( .A1(n2517), .A2(n2516), .A3(n2515), .A4(n2514), .ZN(n4232)
         );
  INV_X1 U32110 ( .A(IR_REG_11__SCAN_IN), .ZN(n2518) );
  NAND2_X1 U32120 ( .A1(n2519), .A2(n2518), .ZN(n2520) );
  NAND2_X1 U32130 ( .A1(n2520), .A2(IR_REG_31__SCAN_IN), .ZN(n2521) );
  XNOR2_X1 U32140 ( .A(n2521), .B(IR_REG_12__SCAN_IN), .ZN(n4709) );
  MUX2_X1 U32150 ( .A(n4709), .B(DATAI_12_), .S(n2640), .Z(n3794) );
  INV_X1 U32160 ( .A(n3811), .ZN(n2530) );
  NAND2_X1 U32170 ( .A1(n2170), .A2(REG2_REG_13__SCAN_IN), .ZN(n2527) );
  NOR2_X1 U32180 ( .A1(n2522), .A2(REG3_REG_13__SCAN_IN), .ZN(n2523) );
  OR2_X1 U32190 ( .A1(n2531), .A2(n2523), .ZN(n3823) );
  INV_X1 U32200 ( .A(n3823), .ZN(n3831) );
  NAND2_X1 U32210 ( .A1(n2422), .A2(n3831), .ZN(n2526) );
  NAND2_X1 U32220 ( .A1(n2732), .A2(REG0_REG_13__SCAN_IN), .ZN(n2525) );
  INV_X1 U32230 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4271) );
  OR2_X1 U32240 ( .A1(n3146), .A2(n4271), .ZN(n2524) );
  NAND4_X1 U32250 ( .A1(n2527), .A2(n2526), .A3(n2525), .A4(n2524), .ZN(n3843)
         );
  OR2_X1 U32260 ( .A1(n2528), .A2(n2663), .ZN(n2529) );
  XNOR2_X1 U32270 ( .A(n2529), .B(IR_REG_13__SCAN_IN), .ZN(n4299) );
  MUX2_X1 U32280 ( .A(n4299), .B(DATAI_13_), .S(n2640), .Z(n3817) );
  NAND2_X1 U32290 ( .A1(n2732), .A2(REG0_REG_14__SCAN_IN), .ZN(n2536) );
  OR2_X1 U32300 ( .A1(n2531), .A2(REG3_REG_14__SCAN_IN), .ZN(n2532) );
  AND2_X1 U32310 ( .A1(n2542), .A2(n2532), .ZN(n3900) );
  NAND2_X1 U32320 ( .A1(n2422), .A2(n3900), .ZN(n2535) );
  NAND2_X1 U32330 ( .A1(n2170), .A2(REG2_REG_14__SCAN_IN), .ZN(n2534) );
  INV_X1 U32340 ( .A(REG1_REG_14__SCAN_IN), .ZN(n3911) );
  OR2_X1 U32350 ( .A1(n3146), .A2(n3911), .ZN(n2533) );
  NAND4_X1 U32360 ( .A1(n2536), .A2(n2535), .A3(n2534), .A4(n2533), .ZN(n4058)
         );
  INV_X1 U32370 ( .A(n2568), .ZN(n2540) );
  NAND2_X1 U32380 ( .A1(n2537), .A2(IR_REG_31__SCAN_IN), .ZN(n2538) );
  MUX2_X1 U32390 ( .A(IR_REG_31__SCAN_IN), .B(n2538), .S(IR_REG_14__SCAN_IN), 
        .Z(n2539) );
  INV_X1 U32400 ( .A(DATAI_14_), .ZN(n4815) );
  MUX2_X1 U32410 ( .A(n4816), .B(n4815), .S(n2640), .Z(n3906) );
  OR2_X1 U32420 ( .A1(n4058), .A2(n3906), .ZN(n4107) );
  NAND2_X1 U32430 ( .A1(n4058), .A2(n3906), .ZN(n4087) );
  NAND2_X1 U32440 ( .A1(n4107), .A2(n4087), .ZN(n4146) );
  NAND2_X1 U32450 ( .A1(n2170), .A2(REG2_REG_15__SCAN_IN), .ZN(n2547) );
  NAND2_X1 U32460 ( .A1(n2542), .A2(n2541), .ZN(n2543) );
  AND2_X1 U32470 ( .A1(n2548), .A2(n2543), .ZN(n4052) );
  NAND2_X1 U32480 ( .A1(n2422), .A2(n4052), .ZN(n2546) );
  NAND2_X1 U32490 ( .A1(n2732), .A2(REG0_REG_15__SCAN_IN), .ZN(n2545) );
  INV_X1 U32500 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3889) );
  OR2_X1 U32510 ( .A1(n3146), .A2(n3889), .ZN(n2544) );
  NAND4_X1 U32520 ( .A1(n2547), .A2(n2546), .A3(n2545), .A4(n2544), .ZN(n4231)
         );
  XNOR2_X1 U32530 ( .A(n2555), .B(IR_REG_15__SCAN_IN), .ZN(n4303) );
  MUX2_X1 U32540 ( .A(n4303), .B(DATAI_15_), .S(n2640), .Z(n2882) );
  NAND2_X1 U32550 ( .A1(n2170), .A2(REG2_REG_16__SCAN_IN), .ZN(n2553) );
  NAND2_X1 U32560 ( .A1(n2548), .A2(n3458), .ZN(n2549) );
  AND2_X1 U32570 ( .A1(n2561), .A2(n2549), .ZN(n3979) );
  NAND2_X1 U32580 ( .A1(n2422), .A2(n3979), .ZN(n2552) );
  NAND2_X1 U32590 ( .A1(n2732), .A2(REG0_REG_16__SCAN_IN), .ZN(n2551) );
  INV_X1 U32600 ( .A(REG1_REG_16__SCAN_IN), .ZN(n3515) );
  OR2_X1 U32610 ( .A1(n3146), .A2(n3515), .ZN(n2550) );
  NAND4_X1 U32620 ( .A1(n2553), .A2(n2552), .A3(n2551), .A4(n2550), .ZN(n4230)
         );
  NAND2_X1 U32630 ( .A1(n2555), .A2(n2554), .ZN(n2556) );
  NAND2_X1 U32640 ( .A1(n2556), .A2(IR_REG_31__SCAN_IN), .ZN(n2557) );
  XNOR2_X1 U32650 ( .A(n2557), .B(IR_REG_16__SCAN_IN), .ZN(n4276) );
  INV_X1 U32660 ( .A(DATAI_16_), .ZN(n4811) );
  MUX2_X1 U32670 ( .A(n4812), .B(n4811), .S(n2640), .Z(n3879) );
  OR2_X1 U32680 ( .A1(n4230), .A2(n3879), .ZN(n4184) );
  NAND2_X1 U32690 ( .A1(n4230), .A2(n3879), .ZN(n4187) );
  NAND2_X1 U32700 ( .A1(n3874), .A2(n2558), .ZN(n3875) );
  NAND2_X1 U32710 ( .A1(n4230), .A2(n3982), .ZN(n2559) );
  NAND2_X1 U32720 ( .A1(n2732), .A2(REG0_REG_17__SCAN_IN), .ZN(n2566) );
  AND2_X1 U32730 ( .A1(n2561), .A2(n2560), .ZN(n2562) );
  NOR2_X1 U32740 ( .A1(n2572), .A2(n2562), .ZN(n3991) );
  NAND2_X1 U32750 ( .A1(n2422), .A2(n3991), .ZN(n2565) );
  NAND2_X1 U32760 ( .A1(n2170), .A2(REG2_REG_17__SCAN_IN), .ZN(n2564) );
  INV_X1 U32770 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4583) );
  OR2_X1 U32780 ( .A1(n3146), .A2(n4583), .ZN(n2563) );
  NAND4_X1 U32790 ( .A1(n2566), .A2(n2565), .A3(n2564), .A4(n2563), .ZN(n4507)
         );
  NOR2_X1 U32800 ( .A1(IR_REG_15__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2567) );
  NAND2_X1 U32810 ( .A1(n2568), .A2(n2567), .ZN(n2578) );
  NAND2_X1 U32820 ( .A1(n2578), .A2(IR_REG_31__SCAN_IN), .ZN(n2569) );
  XNOR2_X1 U32830 ( .A(n2569), .B(IR_REG_17__SCAN_IN), .ZN(n4306) );
  MUX2_X1 U32840 ( .A(n4306), .B(DATAI_17_), .S(n2640), .Z(n3926) );
  OR2_X1 U32850 ( .A1(n4507), .A2(n3926), .ZN(n2571) );
  AND2_X1 U32860 ( .A1(n4507), .A2(n3926), .ZN(n2570) );
  NAND2_X1 U32870 ( .A1(n2732), .A2(REG0_REG_18__SCAN_IN), .ZN(n2577) );
  OR2_X1 U32880 ( .A1(n2572), .A2(REG3_REG_18__SCAN_IN), .ZN(n2573) );
  AND2_X1 U32890 ( .A1(n2573), .A2(n2585), .ZN(n4500) );
  NAND2_X1 U32900 ( .A1(n2422), .A2(n4500), .ZN(n2576) );
  NAND2_X1 U32910 ( .A1(n2170), .A2(REG2_REG_18__SCAN_IN), .ZN(n2575) );
  INV_X1 U32920 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3546) );
  OR2_X1 U32930 ( .A1(n3146), .A2(n3546), .ZN(n2574) );
  NAND4_X1 U32940 ( .A1(n2577), .A2(n2576), .A3(n2575), .A4(n2574), .ZN(n4484)
         );
  NAND2_X1 U32950 ( .A1(n2591), .A2(IR_REG_31__SCAN_IN), .ZN(n2582) );
  INV_X1 U32960 ( .A(IR_REG_18__SCAN_IN), .ZN(n2581) );
  XNOR2_X1 U32970 ( .A(n2582), .B(n2581), .ZN(n4312) );
  INV_X1 U32980 ( .A(DATAI_18_), .ZN(n2583) );
  MUX2_X1 U32990 ( .A(n4312), .B(n2583), .S(n2640), .Z(n4512) );
  OR2_X1 U33000 ( .A1(n4484), .A2(n4512), .ZN(n4479) );
  NAND2_X1 U33010 ( .A1(n4484), .A2(n4512), .ZN(n4477) );
  INV_X1 U33020 ( .A(n4512), .ZN(n4034) );
  OR2_X1 U33030 ( .A1(n4034), .A2(n4484), .ZN(n4472) );
  NAND2_X1 U33040 ( .A1(n2170), .A2(REG2_REG_19__SCAN_IN), .ZN(n2590) );
  NAND2_X1 U33050 ( .A1(n2585), .A2(n2584), .ZN(n2586) );
  AND2_X1 U33060 ( .A1(n2596), .A2(n2586), .ZN(n4491) );
  NAND2_X1 U33070 ( .A1(n2422), .A2(n4491), .ZN(n2589) );
  NAND2_X1 U33080 ( .A1(n2732), .A2(REG0_REG_19__SCAN_IN), .ZN(n2588) );
  INV_X1 U33090 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4571) );
  OR2_X1 U33100 ( .A1(n3146), .A2(n4571), .ZN(n2587) );
  NAND4_X1 U33110 ( .A1(n2590), .A2(n2589), .A3(n2588), .A4(n2587), .ZN(n4509)
         );
  NAND2_X1 U33120 ( .A1(n2593), .A2(n2592), .ZN(n2683) );
  OR2_X1 U33130 ( .A1(n2593), .A2(n2592), .ZN(n2594) );
  MUX2_X1 U33140 ( .A(n4516), .B(DATAI_19_), .S(n2640), .Z(n3952) );
  OR2_X1 U33150 ( .A1(n4509), .A2(n3952), .ZN(n2595) );
  AND2_X1 U33160 ( .A1(n2596), .A2(n4011), .ZN(n2597) );
  NOR2_X1 U33170 ( .A1(n2603), .A2(n2597), .ZN(n4465) );
  NAND2_X1 U33180 ( .A1(n4465), .A2(n2422), .ZN(n2602) );
  NAND2_X1 U33190 ( .A1(n2423), .A2(REG2_REG_20__SCAN_IN), .ZN(n2601) );
  INV_X1 U33200 ( .A(REG1_REG_20__SCAN_IN), .ZN(n2598) );
  OR2_X1 U33210 ( .A1(n3146), .A2(n2598), .ZN(n2600) );
  NAND2_X1 U33220 ( .A1(n2732), .A2(REG0_REG_20__SCAN_IN), .ZN(n2599) );
  NAND4_X1 U33230 ( .A1(n2602), .A2(n2601), .A3(n2600), .A4(n2599), .ZN(n3961)
         );
  NAND2_X1 U33240 ( .A1(n3961), .A2(n4466), .ZN(n4132) );
  OR2_X1 U33250 ( .A1(n3961), .A2(n4466), .ZN(n4133) );
  NOR2_X1 U33260 ( .A1(n2603), .A2(REG3_REG_21__SCAN_IN), .ZN(n2604) );
  OR2_X1 U33270 ( .A1(n2611), .A2(n2604), .ZN(n4441) );
  NAND2_X1 U33280 ( .A1(n2170), .A2(REG2_REG_21__SCAN_IN), .ZN(n2606) );
  INV_X1 U33290 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4562) );
  OR2_X1 U33300 ( .A1(n3146), .A2(n4562), .ZN(n2605) );
  AND2_X1 U33310 ( .A1(n2606), .A2(n2605), .ZN(n2608) );
  NAND2_X1 U33320 ( .A1(n2413), .A2(REG0_REG_21__SCAN_IN), .ZN(n2607) );
  NAND2_X1 U33330 ( .A1(n2640), .A2(DATAI_21_), .ZN(n4557) );
  NAND2_X1 U33340 ( .A1(n4428), .A2(n4447), .ZN(n2610) );
  NOR2_X1 U33350 ( .A1(n4428), .A2(n4447), .ZN(n2609) );
  AOI21_X1 U33360 ( .B1(n4434), .B2(n2610), .A(n2609), .ZN(n4414) );
  OR2_X1 U33370 ( .A1(n2611), .A2(REG3_REG_22__SCAN_IN), .ZN(n2612) );
  NAND2_X1 U33380 ( .A1(n2616), .A2(n2612), .ZN(n4421) );
  INV_X1 U33390 ( .A(n3146), .ZN(n2613) );
  AOI22_X1 U33400 ( .A1(n2613), .A2(REG1_REG_22__SCAN_IN), .B1(n2170), .B2(
        REG2_REG_22__SCAN_IN), .ZN(n2615) );
  NAND2_X1 U33410 ( .A1(n2732), .A2(REG0_REG_22__SCAN_IN), .ZN(n2614) );
  XNOR2_X1 U33420 ( .A(n4403), .B(n4417), .ZN(n4425) );
  INV_X1 U33430 ( .A(n4417), .ZN(n4427) );
  NAND2_X1 U33440 ( .A1(n2616), .A2(n3941), .ZN(n2617) );
  AND2_X1 U33450 ( .A1(n2618), .A2(n2617), .ZN(n4409) );
  NAND2_X1 U33460 ( .A1(n4409), .A2(n2422), .ZN(n2621) );
  AOI22_X1 U33470 ( .A1(n2613), .A2(REG1_REG_23__SCAN_IN), .B1(n2732), .B2(
        REG0_REG_23__SCAN_IN), .ZN(n2620) );
  NAND2_X1 U33480 ( .A1(n2170), .A2(REG2_REG_23__SCAN_IN), .ZN(n2619) );
  INV_X1 U33490 ( .A(n4543), .ZN(n3138) );
  NOR2_X1 U33500 ( .A1(n3138), .A2(n4402), .ZN(n2622) );
  AOI21_X1 U33510 ( .B1(n4406), .B2(n4542), .A(n2623), .ZN(n4356) );
  NOR2_X1 U33520 ( .A1(n2624), .A2(REG3_REG_25__SCAN_IN), .ZN(n2625) );
  INV_X1 U3353 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4540) );
  NAND2_X1 U33540 ( .A1(n2423), .A2(REG2_REG_25__SCAN_IN), .ZN(n2627) );
  NAND2_X1 U3355 ( .A1(n2413), .A2(REG0_REG_25__SCAN_IN), .ZN(n2626) );
  OAI211_X1 U3356 ( .C1(n3146), .C2(n4540), .A(n2627), .B(n2626), .ZN(n2628)
         );
  INV_X1 U3357 ( .A(n2628), .ZN(n2629) );
  NAND2_X1 U3358 ( .A1(n4356), .A2(n2631), .ZN(n2632) );
  INV_X1 U3359 ( .A(n4343), .ZN(n4381) );
  OR2_X1 U3360 ( .A1(n2633), .A2(REG3_REG_26__SCAN_IN), .ZN(n2634) );
  NAND2_X1 U3361 ( .A1(n4351), .A2(n2422), .ZN(n2639) );
  INV_X1 U3362 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4536) );
  NAND2_X1 U3363 ( .A1(n2170), .A2(REG2_REG_26__SCAN_IN), .ZN(n2636) );
  NAND2_X1 U3364 ( .A1(n2413), .A2(REG0_REG_26__SCAN_IN), .ZN(n2635) );
  OAI211_X1 U3365 ( .C1(n3146), .C2(n4536), .A(n2636), .B(n2635), .ZN(n2637)
         );
  INV_X1 U3366 ( .A(n2637), .ZN(n2638) );
  NAND2_X1 U3367 ( .A1(n2640), .A2(DATAI_26_), .ZN(n4349) );
  NOR2_X1 U3368 ( .A1(n4528), .A2(n4349), .ZN(n2641) );
  XNOR2_X1 U3369 ( .A(n2648), .B(REG3_REG_27__SCAN_IN), .ZN(n4329) );
  NAND2_X1 U3370 ( .A1(n4329), .A2(n2422), .ZN(n2646) );
  INV_X1 U3371 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4532) );
  NAND2_X1 U3372 ( .A1(n2170), .A2(REG2_REG_27__SCAN_IN), .ZN(n2643) );
  NAND2_X1 U3373 ( .A1(n2732), .A2(REG0_REG_27__SCAN_IN), .ZN(n2642) );
  OAI211_X1 U3374 ( .C1(n3146), .C2(n4532), .A(n2643), .B(n2642), .ZN(n2644)
         );
  INV_X1 U3375 ( .A(n2644), .ZN(n2645) );
  INV_X1 U3376 ( .A(n4527), .ZN(n4330) );
  NOR2_X1 U3377 ( .A1(n4229), .A2(n4330), .ZN(n2647) );
  INV_X1 U3378 ( .A(n4229), .ZN(n4346) );
  INV_X1 U3379 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3001) );
  INV_X1 U3380 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2992) );
  OAI21_X1 U3381 ( .B1(n2648), .B2(n3001), .A(n2992), .ZN(n2649) );
  NAND2_X1 U3382 ( .A1(n4314), .A2(n2422), .ZN(n2655) );
  INV_X1 U3383 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2652) );
  NAND2_X1 U3384 ( .A1(n2170), .A2(REG2_REG_28__SCAN_IN), .ZN(n2651) );
  NAND2_X1 U3385 ( .A1(n2413), .A2(REG0_REG_28__SCAN_IN), .ZN(n2650) );
  OAI211_X1 U3386 ( .C1(n3146), .C2(n2652), .A(n2651), .B(n2650), .ZN(n2653)
         );
  INV_X1 U3387 ( .A(n2653), .ZN(n2654) );
  NAND2_X1 U3388 ( .A1(n4228), .A2(n2989), .ZN(n2726) );
  NAND2_X1 U3389 ( .A1(n4325), .A2(n2656), .ZN(n4123) );
  NAND2_X1 U3390 ( .A1(n2726), .A2(n4123), .ZN(n4131) );
  INV_X1 U3391 ( .A(n2740), .ZN(n2660) );
  NAND2_X1 U3392 ( .A1(n2423), .A2(REG2_REG_29__SCAN_IN), .ZN(n2658) );
  NAND2_X1 U3393 ( .A1(n2413), .A2(REG0_REG_29__SCAN_IN), .ZN(n2657) );
  OAI211_X1 U3394 ( .C1(n2767), .C2(n3146), .A(n2658), .B(n2657), .ZN(n2659)
         );
  AOI21_X1 U3395 ( .B1(n2660), .B2(n2422), .A(n2659), .ZN(n4125) );
  NAND2_X1 U3396 ( .A1(n2640), .A2(DATAI_29_), .ZN(n4065) );
  XNOR2_X1 U3397 ( .A(n4125), .B(n4065), .ZN(n4165) );
  XNOR2_X1 U3398 ( .A(n2661), .B(n4165), .ZN(n2766) );
  NAND2_X1 U3399 ( .A1(n2662), .A2(n2666), .ZN(n2667) );
  NAND2_X1 U3400 ( .A1(n2667), .A2(IR_REG_31__SCAN_IN), .ZN(n2668) );
  NAND2_X1 U3401 ( .A1(n2677), .A2(n3027), .ZN(n2669) );
  MUX2_X1 U3402 ( .A(n2677), .B(n2669), .S(B_REG_SCAN_IN), .Z(n2673) );
  NAND2_X1 U3403 ( .A1(n2662), .A2(n2670), .ZN(n2671) );
  INV_X1 U3404 ( .A(D_REG_0__SCAN_IN), .ZN(n3932) );
  NAND2_X1 U3405 ( .A1(n2700), .A2(n3932), .ZN(n2676) );
  INV_X1 U3406 ( .A(n2678), .ZN(n2674) );
  NAND2_X1 U3407 ( .A1(n2677), .A2(n2674), .ZN(n2675) );
  OAI22_X1 U3408 ( .A1(n3025), .A2(D_REG_1__SCAN_IN), .B1(n3015), .B2(n2678), 
        .ZN(n2751) );
  INV_X1 U3409 ( .A(n2751), .ZN(n2968) );
  INV_X1 U3410 ( .A(n2677), .ZN(n2679) );
  NAND2_X1 U3411 ( .A1(n2738), .A2(n4648), .ZN(n2970) );
  NAND2_X1 U3412 ( .A1(n2185), .A2(IR_REG_31__SCAN_IN), .ZN(n2686) );
  NAND2_X1 U3413 ( .A1(n2687), .A2(IR_REG_31__SCAN_IN), .ZN(n2688) );
  MUX2_X1 U3414 ( .A(IR_REG_31__SCAN_IN), .B(n2688), .S(IR_REG_21__SCAN_IN), 
        .Z(n2689) );
  NAND2_X1 U3415 ( .A1(n2689), .A2(n2185), .ZN(n2736) );
  NAND2_X1 U3416 ( .A1(n2970), .A2(n3029), .ZN(n2985) );
  NOR4_X1 U3417 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_22__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_18__SCAN_IN), .ZN(n2698) );
  NOR4_X1 U3418 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_5__SCAN_IN), .A3(
        D_REG_10__SCAN_IN), .A4(D_REG_27__SCAN_IN), .ZN(n2697) );
  INV_X1 U3419 ( .A(D_REG_17__SCAN_IN), .ZN(n4800) );
  INV_X1 U3420 ( .A(D_REG_3__SCAN_IN), .ZN(n4804) );
  INV_X1 U3421 ( .A(D_REG_19__SCAN_IN), .ZN(n4798) );
  INV_X1 U3422 ( .A(D_REG_28__SCAN_IN), .ZN(n4792) );
  NAND4_X1 U3423 ( .A1(n4800), .A2(n4804), .A3(n4798), .A4(n4792), .ZN(n2695)
         );
  NOR4_X1 U3424 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(D_REG_11__SCAN_IN), .ZN(n2693) );
  NOR4_X1 U3425 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_21__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_4__SCAN_IN), .ZN(n2692) );
  NOR4_X1 U3426 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_20__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_30__SCAN_IN), .ZN(n2691) );
  NOR4_X1 U3427 ( .A1(D_REG_12__SCAN_IN), .A2(D_REG_13__SCAN_IN), .A3(
        D_REG_14__SCAN_IN), .A4(D_REG_15__SCAN_IN), .ZN(n2690) );
  NAND4_X1 U3428 ( .A1(n2693), .A2(n2692), .A3(n2691), .A4(n2690), .ZN(n2694)
         );
  NOR4_X1 U3429 ( .A1(D_REG_25__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(n2695), 
        .A4(n2694), .ZN(n2696) );
  NAND3_X1 U3430 ( .A1(n2698), .A2(n2697), .A3(n2696), .ZN(n2699) );
  NAND2_X1 U3431 ( .A1(n2700), .A2(n2699), .ZN(n2966) );
  NAND4_X1 U3432 ( .A1(n2758), .A2(n2968), .A3(n3114), .A4(n2966), .ZN(n2702)
         );
  NAND2_X1 U3433 ( .A1(n2738), .A2(n4516), .ZN(n4783) );
  XNOR2_X1 U3434 ( .A(n2777), .B(n4631), .ZN(n2703) );
  NAND2_X1 U3435 ( .A1(n2703), .A2(n4648), .ZN(n3842) );
  OR2_X1 U3436 ( .A1(n2777), .A2(n4648), .ZN(n3253) );
  NAND2_X1 U3437 ( .A1(n3842), .A2(n3253), .ZN(n2704) );
  NAND2_X1 U3438 ( .A1(n3245), .A2(n2706), .ZN(n3213) );
  INV_X1 U3439 ( .A(n4145), .ZN(n3212) );
  NAND2_X1 U3440 ( .A1(n3213), .A2(n3212), .ZN(n2707) );
  NAND2_X1 U3441 ( .A1(n2707), .A2(n4069), .ZN(n3202) );
  INV_X2 U3442 ( .A(n3209), .ZN(n3203) );
  OR2_X1 U3443 ( .A1(n4234), .A2(n3203), .ZN(n4074) );
  NAND2_X1 U3444 ( .A1(n4234), .A2(n3203), .ZN(n4071) );
  AND2_X1 U3445 ( .A1(n4074), .A2(n4071), .ZN(n3200) );
  INV_X1 U3446 ( .A(n4075), .ZN(n2708) );
  INV_X1 U3447 ( .A(n3631), .ZN(n3298) );
  AND2_X1 U3448 ( .A1(n4233), .A2(n3298), .ZN(n3297) );
  OR2_X1 U3449 ( .A1(n4233), .A2(n3298), .ZN(n4090) );
  OAI21_X2 U3450 ( .B1(n3299), .B2(n3297), .A(n4090), .ZN(n3592) );
  NAND2_X1 U3451 ( .A1(n3665), .A2(n3595), .ZN(n4089) );
  OR2_X1 U3452 ( .A1(n3665), .A2(n3595), .ZN(n4080) );
  INV_X1 U3453 ( .A(n2709), .ZN(n2710) );
  INV_X1 U3454 ( .A(n3678), .ZN(n2711) );
  OR2_X1 U3455 ( .A1(n3695), .A2(n2711), .ZN(n4084) );
  NAND2_X1 U3456 ( .A1(n3638), .A2(n4084), .ZN(n2712) );
  NAND2_X1 U3457 ( .A1(n3695), .A2(n2711), .ZN(n4082) );
  INV_X1 U34580 ( .A(n3657), .ZN(n3739) );
  AND2_X1 U34590 ( .A1(n3759), .A2(n3739), .ZN(n4099) );
  OR2_X1 U3460 ( .A1(n3759), .A2(n3739), .ZN(n4085) );
  NAND2_X1 U3461 ( .A1(n3801), .A2(n3760), .ZN(n4101) );
  OR2_X1 U3462 ( .A1(n3801), .A2(n3760), .ZN(n4097) );
  NAND2_X1 U3463 ( .A1(n2713), .A2(n4097), .ZN(n3701) );
  INV_X1 U3464 ( .A(n3794), .ZN(n3777) );
  NAND2_X1 U3465 ( .A1(n4232), .A2(n3777), .ZN(n3813) );
  INV_X1 U3466 ( .A(n3817), .ZN(n3833) );
  NAND2_X1 U34670 ( .A1(n3843), .A2(n3833), .ZN(n2714) );
  NAND2_X1 U3468 ( .A1(n3813), .A2(n2714), .ZN(n2715) );
  INV_X1 U34690 ( .A(n2715), .ZN(n4103) );
  OR2_X1 U3470 ( .A1(n4232), .A2(n3777), .ZN(n3812) );
  NAND2_X1 U34710 ( .A1(n3770), .A2(n3812), .ZN(n2717) );
  NOR2_X1 U3472 ( .A1(n3843), .A2(n3833), .ZN(n2716) );
  AOI21_X1 U34730 ( .B1(n4103), .B2(n2717), .A(n2716), .ZN(n4105) );
  OR2_X1 U3474 ( .A1(n4231), .A2(n4055), .ZN(n4106) );
  NAND2_X1 U34750 ( .A1(n4231), .A2(n4055), .ZN(n4088) );
  NAND2_X1 U3476 ( .A1(n4106), .A2(n4088), .ZN(n4147) );
  INV_X1 U34770 ( .A(n4107), .ZN(n2718) );
  NOR2_X1 U3478 ( .A1(n4147), .A2(n2718), .ZN(n2719) );
  NAND2_X1 U34790 ( .A1(n3854), .A2(n2719), .ZN(n2720) );
  INV_X1 U3480 ( .A(n4187), .ZN(n4109) );
  INV_X1 U34810 ( .A(n3926), .ZN(n4576) );
  NAND2_X1 U3482 ( .A1(n4507), .A2(n4576), .ZN(n4186) );
  NAND2_X1 U34830 ( .A1(n4509), .A2(n4488), .ZN(n2721) );
  AND2_X1 U3484 ( .A1(n4477), .A2(n2721), .ZN(n4188) );
  OR2_X1 U34850 ( .A1(n4507), .A2(n4576), .ZN(n4474) );
  NAND2_X1 U3486 ( .A1(n4479), .A2(n4474), .ZN(n2723) );
  NOR2_X1 U34870 ( .A1(n4509), .A2(n4488), .ZN(n2722) );
  AOI21_X1 U3488 ( .B1(n4188), .B2(n2723), .A(n2722), .ZN(n4453) );
  INV_X1 U34890 ( .A(n4466), .ZN(n4457) );
  OR2_X1 U3490 ( .A1(n3961), .A2(n4457), .ZN(n2724) );
  AND2_X1 U34910 ( .A1(n3961), .A2(n4457), .ZN(n4190) );
  AOI21_X2 U3492 ( .B1(n4454), .B2(n4191), .A(n4190), .ZN(n4436) );
  OR2_X1 U34930 ( .A1(n4403), .A2(n4417), .ZN(n4398) );
  OR2_X1 U3494 ( .A1(n4428), .A2(n4557), .ZN(n4395) );
  NAND2_X1 U34950 ( .A1(n4398), .A2(n4395), .ZN(n4194) );
  AND2_X1 U3496 ( .A1(n4428), .A2(n4557), .ZN(n4140) );
  INV_X1 U34970 ( .A(n4403), .ZN(n4437) );
  OAI22_X1 U3498 ( .A1(n4543), .A2(n4402), .B1(n4437), .B2(n4427), .ZN(n4115)
         );
  AOI21_X1 U34990 ( .B1(n4140), .B2(n4398), .A(n4115), .ZN(n4193) );
  OAI21_X1 U3500 ( .B1(n4436), .B2(n4194), .A(n4193), .ZN(n4378) );
  NOR2_X1 U35010 ( .A1(n4363), .A2(n4542), .ZN(n4135) );
  NOR2_X1 U3502 ( .A1(n3138), .A2(n4408), .ZN(n4376) );
  NOR2_X1 U35030 ( .A1(n4135), .A2(n4376), .ZN(n4198) );
  NAND2_X1 U3504 ( .A1(n4343), .A2(n4367), .ZN(n4162) );
  NAND2_X1 U35050 ( .A1(n4363), .A2(n4542), .ZN(n4134) );
  NAND2_X1 U35060 ( .A1(n4162), .A2(n4134), .ZN(n4196) );
  OR2_X1 U35070 ( .A1(n4343), .A2(n4367), .ZN(n4163) );
  OAI21_X2 U35080 ( .B1(n4358), .B2(n4196), .A(n4163), .ZN(n4340) );
  NOR2_X1 U35090 ( .A1(n4332), .A2(n4349), .ZN(n4161) );
  NAND2_X1 U35100 ( .A1(n4332), .A2(n4349), .ZN(n4178) );
  OAI21_X1 U35110 ( .B1(n4340), .B2(n4161), .A(n4178), .ZN(n4324) );
  OR2_X1 U35120 ( .A1(n4229), .A2(n4527), .ZN(n4122) );
  NAND2_X1 U35130 ( .A1(n4229), .A2(n4527), .ZN(n4121) );
  NAND2_X1 U35140 ( .A1(n4122), .A2(n4121), .ZN(n4323) );
  NOR2_X2 U35150 ( .A1(n4324), .A2(n4323), .ZN(n4322) );
  INV_X1 U35160 ( .A(n4122), .ZN(n2725) );
  NOR2_X1 U35170 ( .A1(n4322), .A2(n2725), .ZN(n2747) );
  INV_X1 U35180 ( .A(n2726), .ZN(n4064) );
  INV_X1 U35190 ( .A(n2738), .ZN(n4632) );
  NAND2_X1 U35200 ( .A1(n4632), .A2(n4212), .ZN(n2728) );
  INV_X1 U35210 ( .A(n4631), .ZN(n2737) );
  OR2_X1 U35220 ( .A1(n4648), .A2(n2737), .ZN(n2727) );
  XNOR2_X1 U35230 ( .A(n2729), .B(IR_REG_27__SCAN_IN), .ZN(n4672) );
  NAND2_X1 U35240 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(
        n2730) );
  NAND2_X1 U35250 ( .A1(n2729), .A2(n2730), .ZN(n2731) );
  AOI21_X1 U35260 ( .B1(n4672), .B2(B_REG_SCAN_IN), .A(n4482), .ZN(n4523) );
  INV_X1 U35270 ( .A(REG1_REG_30__SCAN_IN), .ZN(n2735) );
  NAND2_X1 U35280 ( .A1(n2423), .A2(REG2_REG_30__SCAN_IN), .ZN(n2734) );
  NAND2_X1 U35290 ( .A1(n2732), .A2(REG0_REG_30__SCAN_IN), .ZN(n2733) );
  OAI211_X1 U35300 ( .C1(n2404), .C2(n2735), .A(n2734), .B(n2733), .ZN(n4226)
         );
  NAND2_X1 U35310 ( .A1(n2793), .A2(n3118), .ZN(n3257) );
  NAND2_X1 U35320 ( .A1(n3221), .A2(n3203), .ZN(n3207) );
  OR2_X2 U35330 ( .A1(n3207), .A2(n3193), .ZN(n3302) );
  NOR2_X4 U35340 ( .A1(n3302), .A2(n3631), .ZN(n3596) );
  AND2_X2 U35350 ( .A1(n3727), .A2(n3760), .ZN(n3729) );
  NAND2_X2 U35360 ( .A1(n4501), .A2(n4488), .ZN(n4490) );
  OAI21_X1 U35370 ( .B1(n2754), .B2(n4065), .A(n4522), .ZN(n2774) );
  AND2_X1 U35380 ( .A1(n4829), .A2(n4648), .ZN(n2739) );
  INV_X1 U35390 ( .A(n3029), .ZN(n2741) );
  NAND2_X1 U35400 ( .A1(n4517), .A2(n4506), .ZN(n4444) );
  INV_X1 U35410 ( .A(REG2_REG_29__SCAN_IN), .ZN(n2742) );
  OAI22_X1 U35420 ( .A1(n4325), .A2(n4444), .B1(n2742), .B2(n4517), .ZN(n2744)
         );
  INV_X1 U35430 ( .A(n4065), .ZN(n4124) );
  AND2_X1 U35440 ( .A1(n4446), .A2(n4124), .ZN(n2743) );
  XNOR2_X1 U35450 ( .A(n2747), .B(n4131), .ZN(n2750) );
  NOR2_X1 U35460 ( .A1(n4346), .A2(n4578), .ZN(n2749) );
  OAI22_X1 U35470 ( .A1(n4125), .A2(n4482), .B1(n4577), .B2(n2989), .ZN(n2748)
         );
  AOI211_X2 U35480 ( .C1(n2750), .C2(n4514), .A(n2749), .B(n2748), .ZN(n4313)
         );
  OAI21_X1 U35490 ( .B1(n4320), .B2(n4590), .A(n4313), .ZN(n2760) );
  INV_X1 U35500 ( .A(n2753), .ZN(n2757) );
  INV_X1 U35510 ( .A(n2754), .ZN(n2755) );
  OAI21_X1 U35520 ( .B1(n4327), .B2(n2989), .A(n2755), .ZN(n4316) );
  NAND2_X1 U35530 ( .A1(n2757), .A2(n2756), .ZN(U3546) );
  INV_X1 U35540 ( .A(n2761), .ZN(n2763) );
  NAND2_X1 U35550 ( .A1(n2763), .A2(n2762), .ZN(U3514) );
  AOI22_X1 U35560 ( .A1(n4228), .A2(n4506), .B1(n4124), .B2(n4658), .ZN(n2764)
         );
  NAND2_X1 U35570 ( .A1(n2773), .A2(n4867), .ZN(n2770) );
  NOR2_X1 U35580 ( .A1(n2774), .A2(n4585), .ZN(n2768) );
  NOR2_X1 U35590 ( .A1(n2768), .A2(n2349), .ZN(n2769) );
  OAI21_X1 U35600 ( .B1(n2773), .B2(n4858), .A(n2772), .ZN(n2775) );
  NAND2_X1 U35610 ( .A1(n2775), .A2(n2362), .ZN(U3515) );
  INV_X1 U35620 ( .A(n2777), .ZN(n2776) );
  NAND2_X2 U35630 ( .A1(n2776), .A2(n2172), .ZN(n2783) );
  NAND2_X1 U35640 ( .A1(n3229), .A2(n2804), .ZN(n2780) );
  NAND2_X1 U35650 ( .A1(n3193), .A2(n2789), .ZN(n2779) );
  NAND2_X1 U35660 ( .A1(n4648), .A2(n4631), .ZN(n2978) );
  AND2_X2 U35670 ( .A1(n2777), .A2(n2978), .ZN(n2956) );
  NAND2_X2 U35680 ( .A1(n2789), .A2(n2782), .ZN(n2866) );
  NOR2_X1 U35690 ( .A1(n3271), .A2(n2783), .ZN(n2784) );
  AOI21_X1 U35700 ( .B1(n3229), .B2(n2959), .A(n2784), .ZN(n2821) );
  NAND2_X1 U35710 ( .A1(n4234), .A2(n2919), .ZN(n2786) );
  NAND2_X1 U35720 ( .A1(n3209), .A2(n2789), .ZN(n2785) );
  INV_X1 U35730 ( .A(n2818), .ZN(n2788) );
  AOI22_X1 U35740 ( .A1(n4234), .A2(n2959), .B1(n3209), .B2(n2953), .ZN(n2817)
         );
  NAND2_X1 U35750 ( .A1(n2788), .A2(n2817), .ZN(n3190) );
  AND2_X1 U35760 ( .A1(n3189), .A2(n3190), .ZN(n2819) );
  XNOR2_X1 U35770 ( .A(n2792), .B(n2791), .ZN(n2801) );
  NOR2_X1 U35780 ( .A1(n2793), .A2(n2783), .ZN(n2794) );
  AOI21_X1 U35790 ( .B1(n2790), .B2(n2796), .A(n2794), .ZN(n2802) );
  XNOR2_X1 U35800 ( .A(n2801), .B(n2802), .ZN(n3119) );
  INV_X1 U35810 ( .A(IR_REG_0__SCAN_IN), .ZN(n4826) );
  AOI21_X1 U3582 ( .B1(n3247), .B2(n2796), .A(n2795), .ZN(n2797) );
  OAI21_X1 U3583 ( .B1(n3118), .B2(n2783), .A(n2797), .ZN(n3112) );
  NAND2_X1 U3584 ( .A1(n3247), .A2(n2804), .ZN(n2798) );
  NAND2_X1 U3585 ( .A1(n3255), .A2(n2789), .ZN(n2800) );
  OAI211_X1 U3586 ( .C1(n2172), .C2(n2799), .A(n2798), .B(n2800), .ZN(n3113)
         );
  AOI22_X1 U3587 ( .A1(n3112), .A2(n3113), .B1(n2956), .B2(n2800), .ZN(n3120)
         );
  OR2_X1 U3588 ( .A1(n2802), .A2(n2801), .ZN(n2803) );
  INV_X1 U3589 ( .A(n3124), .ZN(n2815) );
  NAND2_X1 U3590 ( .A1(n4236), .A2(n2804), .ZN(n2806) );
  NAND2_X1 U3591 ( .A1(n3222), .A2(n2789), .ZN(n2805) );
  NAND2_X1 U3592 ( .A1(n2806), .A2(n2805), .ZN(n2807) );
  NOR2_X1 U3593 ( .A1(n3214), .A2(n2783), .ZN(n2808) );
  AOI21_X1 U3594 ( .B1(n4236), .B2(n2959), .A(n2808), .ZN(n2810) );
  NAND2_X1 U3595 ( .A1(n2809), .A2(n2810), .ZN(n2816) );
  INV_X1 U3596 ( .A(n2809), .ZN(n2812) );
  NAND2_X1 U3597 ( .A1(n2812), .A2(n2811), .ZN(n2813) );
  NAND2_X1 U3598 ( .A1(n2816), .A2(n2813), .ZN(n3127) );
  INV_X1 U3599 ( .A(n3127), .ZN(n2814) );
  NAND2_X1 U3600 ( .A1(n2815), .A2(n2814), .ZN(n3125) );
  NAND2_X1 U3601 ( .A1(n3125), .A2(n2816), .ZN(n3180) );
  XNOR2_X1 U3602 ( .A(n2818), .B(n2817), .ZN(n3182) );
  NAND2_X1 U3603 ( .A1(n3180), .A2(n3182), .ZN(n3181) );
  NAND2_X1 U3604 ( .A1(n2819), .A2(n3181), .ZN(n3188) );
  INV_X1 U3605 ( .A(n2821), .ZN(n2822) );
  NAND2_X1 U3606 ( .A1(n2820), .A2(n2822), .ZN(n2823) );
  NAND2_X1 U3607 ( .A1(n3188), .A2(n2823), .ZN(n3226) );
  NAND2_X1 U3608 ( .A1(n4233), .A2(n2953), .ZN(n2825) );
  NAND2_X1 U3609 ( .A1(n3631), .A2(n2789), .ZN(n2824) );
  NAND2_X1 U3610 ( .A1(n2825), .A2(n2824), .ZN(n2826) );
  AOI22_X1 U3611 ( .A1(n4233), .A2(n2959), .B1(n2953), .B2(n3631), .ZN(n2828)
         );
  XNOR2_X1 U3612 ( .A(n2827), .B(n2828), .ZN(n3225) );
  INV_X1 U3613 ( .A(n2827), .ZN(n2829) );
  NOR2_X1 U3614 ( .A1(n2829), .A2(n2828), .ZN(n2830) );
  NAND2_X1 U3615 ( .A1(n3665), .A2(n2953), .ZN(n2832) );
  NAND2_X1 U3616 ( .A1(n3618), .A2(n2789), .ZN(n2831) );
  NAND2_X1 U3617 ( .A1(n2832), .A2(n2831), .ZN(n2833) );
  XNOR2_X1 U3618 ( .A(n2833), .B(n2956), .ZN(n2835) );
  AOI22_X1 U3619 ( .A1(n3665), .A2(n2959), .B1(n2953), .B2(n3618), .ZN(n2834)
         );
  OR2_X1 U3620 ( .A1(n2835), .A2(n2834), .ZN(n3235) );
  AND2_X1 U3621 ( .A1(n2835), .A2(n2834), .ZN(n3234) );
  AOI21_X1 U3622 ( .B1(n3233), .B2(n3235), .A(n3234), .ZN(n3308) );
  NAND2_X1 U3623 ( .A1(n3679), .A2(n2919), .ZN(n2837) );
  NAND2_X1 U3624 ( .A1(n3314), .A2(n2789), .ZN(n2836) );
  NAND2_X1 U3625 ( .A1(n2837), .A2(n2836), .ZN(n2838) );
  XNOR2_X1 U3626 ( .A(n2838), .B(n2791), .ZN(n2842) );
  NOR2_X1 U3627 ( .A1(n3668), .A2(n2783), .ZN(n2839) );
  AOI21_X1 U3628 ( .B1(n3679), .B2(n2959), .A(n2839), .ZN(n2840) );
  XNOR2_X1 U3629 ( .A(n2842), .B(n2840), .ZN(n3307) );
  INV_X1 U3630 ( .A(n2840), .ZN(n2841) );
  AOI22_X1 U3631 ( .A1(n3695), .A2(n2959), .B1(n2953), .B2(n3678), .ZN(n3605)
         );
  AOI22_X1 U3632 ( .A1(n3695), .A2(n2953), .B1(n2789), .B2(n3678), .ZN(n2843)
         );
  XNOR2_X1 U3633 ( .A(n2843), .B(n2791), .ZN(n3606) );
  INV_X1 U3634 ( .A(n3606), .ZN(n2845) );
  INV_X1 U3635 ( .A(n3605), .ZN(n2844) );
  AOI22_X1 U3636 ( .A1(n3759), .A2(n2959), .B1(n3657), .B2(n2953), .ZN(n2850)
         );
  AOI22_X1 U3637 ( .A1(n3759), .A2(n2953), .B1(n3657), .B2(n2789), .ZN(n2846)
         );
  XNOR2_X1 U3638 ( .A(n2846), .B(n2791), .ZN(n2851) );
  XOR2_X1 U3639 ( .A(n2850), .B(n2851), .Z(n3692) );
  NAND2_X1 U3640 ( .A1(n3801), .A2(n2919), .ZN(n2848) );
  NAND2_X1 U3641 ( .A1(n3733), .A2(n2789), .ZN(n2847) );
  NAND2_X1 U3642 ( .A1(n2848), .A2(n2847), .ZN(n2849) );
  XNOR2_X1 U3643 ( .A(n2849), .B(n2791), .ZN(n2852) );
  AOI22_X1 U3644 ( .A1(n3801), .A2(n2959), .B1(n2953), .B2(n3733), .ZN(n2853)
         );
  XNOR2_X1 U3645 ( .A(n2852), .B(n2853), .ZN(n3715) );
  NAND2_X1 U3646 ( .A1(n2851), .A2(n2850), .ZN(n3716) );
  NAND2_X1 U3647 ( .A1(n3714), .A2(n2855), .ZN(n3750) );
  NAND2_X1 U3648 ( .A1(n3724), .A2(n2919), .ZN(n2857) );
  NAND2_X1 U3649 ( .A1(n3709), .A2(n2789), .ZN(n2856) );
  NAND2_X1 U3650 ( .A1(n2857), .A2(n2856), .ZN(n2858) );
  XNOR2_X1 U3651 ( .A(n2858), .B(n2791), .ZN(n2863) );
  NAND2_X1 U3652 ( .A1(n3724), .A2(n2959), .ZN(n2860) );
  NAND2_X1 U3653 ( .A1(n3709), .A2(n2919), .ZN(n2859) );
  NAND2_X1 U3654 ( .A1(n2860), .A2(n2859), .ZN(n2862) );
  NOR2_X1 U3655 ( .A1(n2863), .A2(n2862), .ZN(n3752) );
  INV_X1 U3656 ( .A(n3752), .ZN(n2861) );
  NAND2_X1 U3657 ( .A1(n3750), .A2(n2861), .ZN(n2864) );
  NAND2_X1 U3658 ( .A1(n2863), .A2(n2862), .ZN(n3751) );
  AOI22_X1 U3659 ( .A1(n4232), .A2(n2953), .B1(n2789), .B2(n3794), .ZN(n2865)
         );
  XOR2_X1 U3660 ( .A(n2791), .B(n2865), .Z(n3787) );
  INV_X1 U3661 ( .A(n4232), .ZN(n3819) );
  OAI22_X1 U3662 ( .A1(n3819), .A2(n2963), .B1(n2783), .B2(n3777), .ZN(n3788)
         );
  NAND2_X1 U3663 ( .A1(n3843), .A2(n2919), .ZN(n2868) );
  NAND2_X1 U3664 ( .A1(n3817), .A2(n2789), .ZN(n2867) );
  NAND2_X1 U3665 ( .A1(n2868), .A2(n2867), .ZN(n2869) );
  XNOR2_X1 U3666 ( .A(n2869), .B(n2956), .ZN(n2871) );
  AOI22_X1 U3667 ( .A1(n3843), .A2(n2959), .B1(n2953), .B2(n3817), .ZN(n2870)
         );
  NOR2_X1 U3668 ( .A1(n2871), .A2(n2870), .ZN(n3828) );
  NAND2_X1 U3669 ( .A1(n4058), .A2(n2919), .ZN(n2873) );
  NAND2_X1 U3670 ( .A1(n3902), .A2(n2789), .ZN(n2872) );
  NAND2_X1 U3671 ( .A1(n2873), .A2(n2872), .ZN(n2874) );
  XNOR2_X1 U3672 ( .A(n2874), .B(n2791), .ZN(n2877) );
  NAND2_X1 U3673 ( .A1(n4058), .A2(n2959), .ZN(n2876) );
  NAND2_X1 U3674 ( .A1(n3902), .A2(n2919), .ZN(n2875) );
  NAND2_X1 U3675 ( .A1(n2876), .A2(n2875), .ZN(n2878) );
  NAND2_X1 U3676 ( .A1(n2877), .A2(n2878), .ZN(n3896) );
  NAND2_X1 U3677 ( .A1(n3895), .A2(n3896), .ZN(n3894) );
  INV_X1 U3678 ( .A(n2877), .ZN(n2880) );
  INV_X1 U3679 ( .A(n2878), .ZN(n2879) );
  NAND2_X1 U3680 ( .A1(n2880), .A2(n2879), .ZN(n3898) );
  NAND2_X1 U3681 ( .A1(n3894), .A2(n3898), .ZN(n2892) );
  AOI22_X1 U3682 ( .A1(n4231), .A2(n2953), .B1(n2789), .B2(n2882), .ZN(n2881)
         );
  XNOR2_X1 U3683 ( .A(n2881), .B(n2791), .ZN(n2893) );
  NAND2_X1 U3684 ( .A1(n4231), .A2(n2959), .ZN(n2884) );
  NAND2_X1 U3685 ( .A1(n2882), .A2(n2919), .ZN(n2883) );
  NAND2_X1 U3686 ( .A1(n2884), .A2(n2883), .ZN(n4051) );
  NAND2_X1 U3687 ( .A1(n4230), .A2(n2919), .ZN(n2886) );
  NAND2_X1 U3688 ( .A1(n3982), .A2(n2789), .ZN(n2885) );
  NAND2_X1 U3689 ( .A1(n2886), .A2(n2885), .ZN(n2887) );
  XNOR2_X1 U3690 ( .A(n2887), .B(n2791), .ZN(n2891) );
  NAND2_X1 U3691 ( .A1(n4230), .A2(n2959), .ZN(n2889) );
  NAND2_X1 U3692 ( .A1(n3982), .A2(n2953), .ZN(n2888) );
  NAND2_X1 U3693 ( .A1(n2889), .A2(n2888), .ZN(n2890) );
  NOR2_X1 U3694 ( .A1(n2891), .A2(n2890), .ZN(n2894) );
  AOI21_X1 U3695 ( .B1(n2891), .B2(n2890), .A(n2894), .ZN(n3978) );
  AOI22_X1 U3696 ( .A1(n4507), .A2(n2953), .B1(n2789), .B2(n3926), .ZN(n2895)
         );
  XOR2_X1 U3697 ( .A(n2791), .B(n2895), .Z(n2897) );
  INV_X1 U3698 ( .A(n4507), .ZN(n4032) );
  OAI22_X1 U3699 ( .A1(n4032), .A2(n2963), .B1(n2783), .B2(n4576), .ZN(n2896)
         );
  NAND2_X1 U3700 ( .A1(n2897), .A2(n2896), .ZN(n3988) );
  NOR2_X1 U3701 ( .A1(n2897), .A2(n2896), .ZN(n3987) );
  INV_X1 U3702 ( .A(n4484), .ZN(n3950) );
  OAI22_X1 U3703 ( .A1(n3950), .A2(n2963), .B1(n2783), .B2(n4512), .ZN(n4029)
         );
  AOI22_X1 U3704 ( .A1(n4484), .A2(n2953), .B1(n2789), .B2(n4034), .ZN(n2898)
         );
  XOR2_X1 U3705 ( .A(n2791), .B(n2898), .Z(n4028) );
  AOI22_X1 U3706 ( .A1(n4509), .A2(n2953), .B1(n2789), .B2(n3952), .ZN(n2899)
         );
  XNOR2_X1 U3707 ( .A(n2899), .B(n2791), .ZN(n2901) );
  AOI22_X1 U3708 ( .A1(n4509), .A2(n2959), .B1(n2953), .B2(n3952), .ZN(n2900)
         );
  NAND2_X1 U3709 ( .A1(n2901), .A2(n2900), .ZN(n2902) );
  OAI21_X1 U3710 ( .B1(n2901), .B2(n2900), .A(n2902), .ZN(n3949) );
  NAND2_X1 U3711 ( .A1(n3947), .A2(n2902), .ZN(n4006) );
  NAND2_X1 U3712 ( .A1(n3961), .A2(n2953), .ZN(n2904) );
  NAND2_X1 U3713 ( .A1(n4466), .A2(n2789), .ZN(n2903) );
  NAND2_X1 U3714 ( .A1(n2904), .A2(n2903), .ZN(n2905) );
  XNOR2_X1 U3715 ( .A(n2905), .B(n2791), .ZN(n2908) );
  NAND2_X1 U3716 ( .A1(n3961), .A2(n2959), .ZN(n2907) );
  NAND2_X1 U3717 ( .A1(n4466), .A2(n2953), .ZN(n2906) );
  NAND2_X1 U3718 ( .A1(n2907), .A2(n2906), .ZN(n2909) );
  NAND2_X1 U3719 ( .A1(n2908), .A2(n2909), .ZN(n4007) );
  INV_X1 U3720 ( .A(n2908), .ZN(n2911) );
  INV_X1 U3721 ( .A(n2909), .ZN(n2910) );
  NAND2_X1 U3722 ( .A1(n2911), .A2(n2910), .ZN(n4009) );
  NAND2_X1 U3723 ( .A1(n4428), .A2(n2953), .ZN(n2913) );
  NAND2_X1 U3724 ( .A1(n4447), .A2(n2789), .ZN(n2912) );
  NAND2_X1 U3725 ( .A1(n2913), .A2(n2912), .ZN(n2914) );
  XNOR2_X1 U3726 ( .A(n2914), .B(n2791), .ZN(n2918) );
  NAND2_X1 U3727 ( .A1(n4428), .A2(n2959), .ZN(n2916) );
  NAND2_X1 U3728 ( .A1(n4447), .A2(n2919), .ZN(n2915) );
  NAND2_X1 U3729 ( .A1(n2916), .A2(n2915), .ZN(n2917) );
  NOR2_X1 U3730 ( .A1(n2918), .A2(n2917), .ZN(n3956) );
  NAND2_X1 U3731 ( .A1(n2918), .A2(n2917), .ZN(n3957) );
  NAND2_X1 U3732 ( .A1(n4403), .A2(n2919), .ZN(n2921) );
  NAND2_X1 U3733 ( .A1(n4427), .A2(n2789), .ZN(n2920) );
  NAND2_X1 U3734 ( .A1(n2921), .A2(n2920), .ZN(n2922) );
  XNOR2_X1 U3735 ( .A(n2922), .B(n2791), .ZN(n2924) );
  OAI22_X1 U3736 ( .A1(n4437), .A2(n2963), .B1(n4417), .B2(n2783), .ZN(n2923)
         );
  XNOR2_X1 U3737 ( .A(n2924), .B(n2923), .ZN(n4020) );
  NAND2_X1 U3738 ( .A1(n4017), .A2(n2925), .ZN(n3937) );
  INV_X1 U3739 ( .A(n3937), .ZN(n2931) );
  OAI22_X1 U3740 ( .A1(n4543), .A2(n2783), .B1(n2926), .B2(n4408), .ZN(n2927)
         );
  XNOR2_X1 U3741 ( .A(n2927), .B(n2791), .ZN(n2933) );
  OR2_X1 U3742 ( .A1(n4543), .A2(n2963), .ZN(n2929) );
  NAND2_X1 U3743 ( .A1(n4402), .A2(n2953), .ZN(n2928) );
  NAND2_X1 U3744 ( .A1(n2929), .A2(n2928), .ZN(n2932) );
  XNOR2_X1 U3745 ( .A(n2933), .B(n2932), .ZN(n3938) );
  NAND2_X1 U3746 ( .A1(n2933), .A2(n2932), .ZN(n2934) );
  OAI22_X1 U3747 ( .A1(n4406), .A2(n2963), .B1(n2783), .B2(n4542), .ZN(n2936)
         );
  OAI22_X1 U3748 ( .A1(n4406), .A2(n2783), .B1(n2926), .B2(n4542), .ZN(n2935)
         );
  NAND2_X1 U3749 ( .A1(n3996), .A2(n3999), .ZN(n2938) );
  NAND2_X1 U3750 ( .A1(n2937), .A2(n2936), .ZN(n3997) );
  NAND2_X1 U3751 ( .A1(n2938), .A2(n3997), .ZN(n3967) );
  NAND2_X1 U3752 ( .A1(n4343), .A2(n2953), .ZN(n2940) );
  NAND2_X1 U3753 ( .A1(n4362), .A2(n2789), .ZN(n2939) );
  NAND2_X1 U3754 ( .A1(n2940), .A2(n2939), .ZN(n2941) );
  XNOR2_X1 U3755 ( .A(n2941), .B(n2956), .ZN(n3969) );
  NOR2_X1 U3756 ( .A1(n4367), .A2(n2783), .ZN(n2942) );
  AOI21_X1 U3757 ( .B1(n4343), .B2(n2959), .A(n2942), .ZN(n2943) );
  NAND2_X1 U3758 ( .A1(n3969), .A2(n2943), .ZN(n2945) );
  INV_X1 U3759 ( .A(n3969), .ZN(n2944) );
  INV_X1 U3760 ( .A(n2943), .ZN(n3968) );
  NAND2_X1 U3761 ( .A1(n4332), .A2(n2953), .ZN(n2947) );
  NAND2_X1 U3762 ( .A1(n4342), .A2(n2789), .ZN(n2946) );
  NAND2_X1 U3763 ( .A1(n2947), .A2(n2946), .ZN(n2948) );
  XNOR2_X1 U3764 ( .A(n2948), .B(n2791), .ZN(n2952) );
  NAND2_X1 U3765 ( .A1(n4332), .A2(n2959), .ZN(n2950) );
  NAND2_X1 U3766 ( .A1(n4342), .A2(n2953), .ZN(n2949) );
  NAND2_X1 U3767 ( .A1(n2950), .A2(n2949), .ZN(n2951) );
  NAND2_X1 U3768 ( .A1(n2952), .A2(n2951), .ZN(n4039) );
  NAND2_X1 U3769 ( .A1(n4229), .A2(n2953), .ZN(n2955) );
  NAND2_X1 U3770 ( .A1(n4330), .A2(n2789), .ZN(n2954) );
  NAND2_X1 U3771 ( .A1(n2955), .A2(n2954), .ZN(n2957) );
  XNOR2_X1 U3772 ( .A(n2957), .B(n2956), .ZN(n2961) );
  NOR2_X1 U3773 ( .A1(n4527), .A2(n2783), .ZN(n2958) );
  AOI21_X1 U3774 ( .B1(n4229), .B2(n2959), .A(n2958), .ZN(n2960) );
  NOR2_X1 U3775 ( .A1(n2961), .A2(n2960), .ZN(n2976) );
  AOI21_X1 U3776 ( .B1(n2961), .B2(n2960), .A(n2976), .ZN(n2999) );
  OAI22_X1 U3777 ( .A1(n4325), .A2(n2783), .B1(n2989), .B2(n2926), .ZN(n2962)
         );
  XNOR2_X1 U3778 ( .A(n2962), .B(n2791), .ZN(n2965) );
  OAI22_X1 U3779 ( .A1(n4325), .A2(n2963), .B1(n2989), .B2(n2783), .ZN(n2964)
         );
  XNOR2_X1 U3780 ( .A(n2965), .B(n2964), .ZN(n2977) );
  INV_X1 U3781 ( .A(n2977), .ZN(n2974) );
  INV_X1 U3782 ( .A(n2976), .ZN(n2972) );
  NAND3_X1 U3783 ( .A1(n2968), .A2(n2967), .A3(n2966), .ZN(n2984) );
  INV_X1 U3784 ( .A(n3031), .ZN(n2969) );
  AOI21_X1 U3785 ( .B1(n2970), .B2(n3098), .A(n3029), .ZN(n2971) );
  NAND2_X1 U3786 ( .A1(n2975), .A2(n2351), .ZN(n2998) );
  NAND3_X1 U3787 ( .A1(n3006), .A2(n3713), .A3(n2977), .ZN(n2997) );
  NAND3_X1 U3788 ( .A1(n2977), .A2(n3713), .A3(n2976), .ZN(n2996) );
  INV_X1 U3789 ( .A(n2984), .ZN(n2981) );
  NOR2_X1 U3790 ( .A1(n2777), .A2(n2978), .ZN(n2979) );
  AND2_X1 U3791 ( .A1(n3031), .A2(n2979), .ZN(n2980) );
  NAND2_X1 U3792 ( .A1(n2981), .A2(n2980), .ZN(n2991) );
  INV_X1 U3793 ( .A(n2991), .ZN(n2982) );
  INV_X1 U3794 ( .A(n4314), .ZN(n2990) );
  NAND2_X1 U3795 ( .A1(n2984), .A2(n2983), .ZN(n3115) );
  AND3_X1 U3796 ( .A1(n2985), .A2(n2172), .A3(n3030), .ZN(n2986) );
  NAND2_X1 U3797 ( .A1(n3115), .A2(n2986), .ZN(n2987) );
  OAI22_X1 U3798 ( .A1(n2990), .A2(n4021), .B1(n4056), .B2(n2989), .ZN(n2994)
         );
  OAI22_X1 U3799 ( .A1(n4125), .A2(n4022), .B1(STATE_REG_SCAN_IN), .B2(n2992), 
        .ZN(n2993) );
  AOI211_X1 U3800 ( .C1(n4059), .C2(n4229), .A(n2994), .B(n2993), .ZN(n2995)
         );
  NAND3_X1 U3801 ( .A1(n2998), .A2(n2997), .A3(n2357), .ZN(U3217) );
  OAI21_X1 U3802 ( .B1(n3000), .B2(n2999), .A(n3713), .ZN(n3007) );
  OAI22_X1 U3803 ( .A1(n4528), .A2(n4043), .B1(STATE_REG_SCAN_IN), .B2(n3001), 
        .ZN(n3004) );
  INV_X1 U3804 ( .A(n4329), .ZN(n3002) );
  OAI22_X1 U3805 ( .A1(n4325), .A2(n4022), .B1(n4021), .B2(n3002), .ZN(n3003)
         );
  AOI211_X1 U3806 ( .C1(n4330), .C2(n4041), .A(n3004), .B(n3003), .ZN(n3005)
         );
  INV_X1 U3807 ( .A(n4807), .ZN(n3026) );
  INV_X2 U3808 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  MUX2_X1 U3809 ( .A(n3008), .B(n3176), .S(STATE_REG_SCAN_IN), .Z(n3009) );
  INV_X1 U3810 ( .A(n3009), .ZN(U3348) );
  INV_X1 U3811 ( .A(DATAI_3_), .ZN(n3010) );
  INV_X1 U3812 ( .A(n3062), .ZN(n3051) );
  MUX2_X1 U3813 ( .A(n3010), .B(n3051), .S(STATE_REG_SCAN_IN), .Z(n3011) );
  INV_X1 U3814 ( .A(n3011), .ZN(U3349) );
  MUX2_X1 U3815 ( .A(n3460), .B(n3158), .S(STATE_REG_SCAN_IN), .Z(n3012) );
  INV_X1 U3816 ( .A(n3012), .ZN(U3345) );
  INV_X1 U3817 ( .A(DATAI_21_), .ZN(n3014) );
  NAND2_X1 U3818 ( .A1(n4212), .A2(STATE_REG_SCAN_IN), .ZN(n3013) );
  OAI21_X1 U3819 ( .B1(STATE_REG_SCAN_IN), .B2(n3014), .A(n3013), .ZN(U3331)
         );
  INV_X1 U3820 ( .A(DATAI_25_), .ZN(n3431) );
  NAND2_X1 U3821 ( .A1(n3015), .A2(STATE_REG_SCAN_IN), .ZN(n3016) );
  OAI21_X1 U3822 ( .B1(STATE_REG_SCAN_IN), .B2(n3431), .A(n3016), .ZN(U3327)
         );
  INV_X1 U3823 ( .A(DATAI_19_), .ZN(n3432) );
  MUX2_X1 U3824 ( .A(n4648), .B(n3432), .S(U3149), .Z(n3017) );
  INV_X1 U3825 ( .A(n3017), .ZN(U3333) );
  INV_X1 U3826 ( .A(DATAI_27_), .ZN(n3019) );
  NAND2_X1 U3827 ( .A1(n4672), .A2(STATE_REG_SCAN_IN), .ZN(n3018) );
  OAI21_X1 U3828 ( .B1(STATE_REG_SCAN_IN), .B2(n3019), .A(n3018), .ZN(U3325)
         );
  INV_X1 U3829 ( .A(DATAI_24_), .ZN(n3020) );
  MUX2_X1 U3830 ( .A(n2677), .B(n3020), .S(U3149), .Z(n3021) );
  INV_X1 U3831 ( .A(n3021), .ZN(U3328) );
  INV_X1 U3832 ( .A(DATAI_29_), .ZN(n3557) );
  NAND2_X1 U3833 ( .A1(n2382), .A2(STATE_REG_SCAN_IN), .ZN(n3022) );
  OAI21_X1 U3834 ( .B1(STATE_REG_SCAN_IN), .B2(n3557), .A(n3022), .ZN(U3323)
         );
  INV_X1 U3835 ( .A(DATAI_30_), .ZN(n3559) );
  NAND2_X1 U3836 ( .A1(n3023), .A2(STATE_REG_SCAN_IN), .ZN(n3024) );
  OAI21_X1 U3837 ( .B1(STATE_REG_SCAN_IN), .B2(n3559), .A(n3024), .ZN(U3322)
         );
  INV_X1 U3838 ( .A(D_REG_1__SCAN_IN), .ZN(n3028) );
  NOR2_X1 U3839 ( .A1(n3026), .A2(n2678), .ZN(n3931) );
  AOI22_X1 U3840 ( .A1(n4806), .A2(n3028), .B1(n3931), .B2(n3027), .ZN(U3459)
         );
  INV_X1 U3841 ( .A(n3042), .ZN(n3032) );
  OR2_X1 U3842 ( .A1(n3030), .A2(U3149), .ZN(n4224) );
  INV_X1 U3843 ( .A(n4224), .ZN(n4221) );
  NOR2_X1 U3844 ( .A1(n4768), .A2(U4043), .ZN(U3148) );
  INV_X1 U3845 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n3034) );
  NAND2_X1 U3846 ( .A1(n3961), .A2(U4043), .ZN(n3033) );
  OAI21_X1 U3847 ( .B1(U4043), .B2(n3034), .A(n3033), .ZN(U3570) );
  INV_X1 U3848 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n3036) );
  NAND2_X1 U3849 ( .A1(n3801), .A2(U4043), .ZN(n3035) );
  OAI21_X1 U3850 ( .B1(U4043), .B2(n3036), .A(n3035), .ZN(U3560) );
  INV_X1 U3851 ( .A(DATAO_REG_9__SCAN_IN), .ZN(n3038) );
  NAND2_X1 U3852 ( .A1(n3759), .A2(U4043), .ZN(n3037) );
  OAI21_X1 U3853 ( .B1(U4043), .B2(n3038), .A(n3037), .ZN(U3559) );
  INV_X1 U3854 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3040) );
  MUX2_X1 U3855 ( .A(n3040), .B(REG2_REG_2__SCAN_IN), .S(n4255), .Z(n4249) );
  XNOR2_X1 U3856 ( .A(n3047), .B(REG2_REG_1__SCAN_IN), .ZN(n4242) );
  AND2_X1 U3857 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n4241)
         );
  NAND2_X1 U3858 ( .A1(n4242), .A2(n4241), .ZN(n4240) );
  INV_X1 U3859 ( .A(n3047), .ZN(n4636) );
  NAND2_X1 U3860 ( .A1(n4636), .A2(REG2_REG_1__SCAN_IN), .ZN(n3039) );
  NAND2_X1 U3861 ( .A1(n4240), .A2(n3039), .ZN(n4248) );
  XNOR2_X1 U3862 ( .A(n3063), .B(REG2_REG_3__SCAN_IN), .ZN(n3055) );
  INV_X1 U3863 ( .A(n4672), .ZN(n3168) );
  NOR2_X1 U3864 ( .A1(n4654), .A2(n3168), .ZN(n3043) );
  INV_X1 U3865 ( .A(n4775), .ZN(n4256) );
  INV_X1 U3866 ( .A(n4768), .ZN(n3077) );
  INV_X1 U3867 ( .A(ADDR_REG_3__SCAN_IN), .ZN(n3045) );
  OAI22_X1 U3868 ( .A1(n3077), .A2(n3045), .B1(STATE_REG_SCAN_IN), .B2(n3044), 
        .ZN(n3046) );
  AOI21_X1 U3869 ( .B1(n3062), .B2(n4256), .A(n3046), .ZN(n3054) );
  XNOR2_X1 U3870 ( .A(n4255), .B(REG1_REG_2__SCAN_IN), .ZN(n4252) );
  XNOR2_X1 U3871 ( .A(n3047), .B(REG1_REG_1__SCAN_IN), .ZN(n4239) );
  AND2_X1 U3872 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n4238)
         );
  NAND2_X1 U3873 ( .A1(n4239), .A2(n4238), .ZN(n4237) );
  NAND2_X1 U3874 ( .A1(n4636), .A2(REG1_REG_1__SCAN_IN), .ZN(n3048) );
  NAND2_X1 U3875 ( .A1(n4237), .A2(n3048), .ZN(n4251) );
  NAND2_X1 U3876 ( .A1(n4252), .A2(n4251), .ZN(n4250) );
  OR2_X1 U3877 ( .A1(n4255), .A2(n3049), .ZN(n3050) );
  NAND2_X1 U3878 ( .A1(n4250), .A2(n3050), .ZN(n3056) );
  XNOR2_X1 U3879 ( .A(n3056), .B(n3051), .ZN(n3052) );
  NAND2_X1 U3880 ( .A1(n3052), .A2(REG1_REG_3__SCAN_IN), .ZN(n3058) );
  OAI211_X1 U3881 ( .C1(REG1_REG_3__SCAN_IN), .C2(n3052), .A(n4769), .B(n3058), 
        .ZN(n3053) );
  OAI211_X1 U3882 ( .C1(n3055), .C2(n4762), .A(n3054), .B(n3053), .ZN(U3243)
         );
  INV_X1 U3883 ( .A(n3176), .ZN(n3066) );
  NAND2_X1 U3884 ( .A1(n3056), .A2(n3062), .ZN(n3057) );
  NAND2_X1 U3885 ( .A1(n3058), .A2(n3057), .ZN(n3059) );
  XNOR2_X1 U3886 ( .A(n3059), .B(n3176), .ZN(n3172) );
  XNOR2_X1 U3887 ( .A(n4635), .B(REG1_REG_5__SCAN_IN), .ZN(n3060) );
  INV_X1 U3888 ( .A(n4769), .ZN(n3079) );
  AOI211_X1 U3889 ( .C1(n3061), .C2(n3060), .A(n3078), .B(n3079), .ZN(n3074)
         );
  XNOR2_X1 U3890 ( .A(n3064), .B(n3176), .ZN(n3170) );
  INV_X1 U3891 ( .A(n3170), .ZN(n3067) );
  INV_X1 U3892 ( .A(n3064), .ZN(n3065) );
  INV_X1 U3893 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3629) );
  MUX2_X1 U3894 ( .A(n3629), .B(REG2_REG_5__SCAN_IN), .S(n4635), .Z(n3068) );
  AOI211_X1 U3895 ( .C1(n3069), .C2(n3068), .A(n3075), .B(n4762), .ZN(n3073)
         );
  INV_X1 U3896 ( .A(n4635), .ZN(n3071) );
  AND2_X1 U3897 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3228) );
  AOI21_X1 U3898 ( .B1(n4768), .B2(ADDR_REG_5__SCAN_IN), .A(n3228), .ZN(n3070)
         );
  OAI21_X1 U3899 ( .B1(n3071), .B2(n4775), .A(n3070), .ZN(n3072) );
  OR3_X1 U3900 ( .A1(n3074), .A2(n3073), .A3(n3072), .ZN(U3245) );
  XNOR2_X1 U3901 ( .A(n3085), .B(REG2_REG_6__SCAN_IN), .ZN(n3084) );
  INV_X1 U3902 ( .A(ADDR_REG_6__SCAN_IN), .ZN(n3076) );
  NAND2_X1 U3903 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3238) );
  OAI21_X1 U3904 ( .B1(n3077), .B2(n3076), .A(n3238), .ZN(n3082) );
  AOI211_X1 U3905 ( .C1(n3080), .C2(n2450), .A(n3079), .B(n3089), .ZN(n3081)
         );
  AOI211_X1 U3906 ( .C1(n4256), .C2(n4634), .A(n3082), .B(n3081), .ZN(n3083)
         );
  OAI21_X1 U3907 ( .B1(n3084), .B2(n4762), .A(n3083), .ZN(U3246) );
  INV_X1 U3908 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3672) );
  MUX2_X1 U3909 ( .A(REG2_REG_7__SCAN_IN), .B(n3672), .S(n3158), .Z(n3086) );
  NOR2_X1 U3910 ( .A1(n3087), .A2(n3086), .ZN(n3153) );
  AOI211_X1 U3911 ( .C1(n3087), .C2(n3086), .A(n4762), .B(n3153), .ZN(n3096)
         );
  INV_X1 U3912 ( .A(n3088), .ZN(n3090) );
  INV_X1 U3913 ( .A(n3158), .ZN(n3154) );
  XNOR2_X1 U3914 ( .A(n3154), .B(REG1_REG_7__SCAN_IN), .ZN(n3092) );
  OAI21_X1 U3915 ( .B1(n3157), .B2(n3092), .A(n4769), .ZN(n3091) );
  AOI21_X1 U3916 ( .B1(n3157), .B2(n3092), .A(n3091), .ZN(n3095) );
  NAND2_X1 U3917 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3310) );
  NAND2_X1 U3918 ( .A1(n4768), .A2(ADDR_REG_7__SCAN_IN), .ZN(n3093) );
  OAI211_X1 U3919 ( .C1(n4775), .C2(n3158), .A(n3310), .B(n3093), .ZN(n3094)
         );
  OR3_X1 U3920 ( .A1(n3096), .A2(n3095), .A3(n3094), .ZN(U3247) );
  INV_X1 U3921 ( .A(n4831), .ZN(n4844) );
  NAND2_X1 U3922 ( .A1(n3247), .A2(n3118), .ZN(n4067) );
  AND2_X1 U3923 ( .A1(n3097), .A2(n4067), .ZN(n4169) );
  INV_X1 U3924 ( .A(n4169), .ZN(n4787) );
  AND2_X1 U3925 ( .A1(n3255), .A2(n3098), .ZN(n4784) );
  INV_X1 U3926 ( .A(n3842), .ZN(n4463) );
  NOR2_X1 U3927 ( .A1(n4463), .A2(n4514), .ZN(n3099) );
  OAI22_X1 U3928 ( .A1(n4169), .A2(n3099), .B1(n2397), .B2(n4482), .ZN(n4782)
         );
  AOI211_X1 U3929 ( .C1(n4844), .C2(n4787), .A(n4784), .B(n4782), .ZN(n4828)
         );
  NAND2_X1 U3930 ( .A1(n4865), .A2(REG1_REG_0__SCAN_IN), .ZN(n3100) );
  OAI21_X1 U3931 ( .B1(n4828), .B2(n4865), .A(n3100), .ZN(U3518) );
  INV_X1 U3932 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n3102) );
  NAND2_X1 U3933 ( .A1(n3843), .A2(U4043), .ZN(n3101) );
  OAI21_X1 U3934 ( .B1(U4043), .B2(n3102), .A(n3101), .ZN(U3563) );
  INV_X1 U3935 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n3104) );
  NAND2_X1 U3936 ( .A1(n4058), .A2(U4043), .ZN(n3103) );
  OAI21_X1 U3937 ( .B1(U4043), .B2(n3104), .A(n3103), .ZN(U3564) );
  INV_X1 U3938 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n3106) );
  NAND2_X1 U3939 ( .A1(n3695), .A2(U4043), .ZN(n3105) );
  OAI21_X1 U3940 ( .B1(U4043), .B2(n3106), .A(n3105), .ZN(U3558) );
  INV_X1 U3941 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n3549) );
  NAND2_X1 U3942 ( .A1(n3679), .A2(U4043), .ZN(n3107) );
  OAI21_X1 U3943 ( .B1(U4043), .B2(n3549), .A(n3107), .ZN(U3557) );
  INV_X1 U3944 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n3109) );
  NAND2_X1 U3945 ( .A1(n4507), .A2(U4043), .ZN(n3108) );
  OAI21_X1 U3946 ( .B1(U4043), .B2(n3109), .A(n3108), .ZN(U3567) );
  INV_X1 U3947 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n3111) );
  NAND2_X1 U3948 ( .A1(n3724), .A2(U4043), .ZN(n3110) );
  OAI21_X1 U3949 ( .B1(U4043), .B2(n3111), .A(n3110), .ZN(U3561) );
  XOR2_X1 U3950 ( .A(n3113), .B(n3112), .Z(n3166) );
  NAND2_X1 U3951 ( .A1(n3166), .A2(n3713), .ZN(n3117) );
  NAND2_X1 U3952 ( .A1(n3115), .A2(n3114), .ZN(n3128) );
  AOI22_X1 U3953 ( .A1(n4054), .A2(n2790), .B1(REG3_REG_0__SCAN_IN), .B2(n3128), .ZN(n3116) );
  OAI211_X1 U3954 ( .C1(n3118), .C2(n4056), .A(n3117), .B(n3116), .ZN(U3229)
         );
  XNOR2_X1 U3955 ( .A(n3120), .B(n3119), .ZN(n3123) );
  AOI22_X1 U3956 ( .A1(n4059), .A2(n3247), .B1(REG3_REG_1__SCAN_IN), .B2(n3128), .ZN(n3122) );
  AOI22_X1 U3957 ( .A1(n4041), .A2(n3256), .B1(n4054), .B2(n4236), .ZN(n3121)
         );
  OAI211_X1 U3958 ( .C1(n3123), .C2(n4062), .A(n3122), .B(n3121), .ZN(U3219)
         );
  INV_X1 U3959 ( .A(n3125), .ZN(n3126) );
  AOI21_X1 U3960 ( .B1(n3124), .B2(n3127), .A(n3126), .ZN(n3131) );
  AOI22_X1 U3961 ( .A1(n4059), .A2(n2790), .B1(REG3_REG_2__SCAN_IN), .B2(n3128), .ZN(n3130) );
  AOI22_X1 U3962 ( .A1(n4041), .A2(n3222), .B1(n4054), .B2(n4234), .ZN(n3129)
         );
  OAI211_X1 U3963 ( .C1(n3131), .C2(n4062), .A(n3130), .B(n3129), .ZN(U3234)
         );
  INV_X1 U3964 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n3133) );
  NAND2_X1 U3965 ( .A1(n3229), .A2(U4043), .ZN(n3132) );
  OAI21_X1 U3966 ( .B1(U4043), .B2(n3133), .A(n3132), .ZN(U3554) );
  INV_X1 U3967 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n3135) );
  NAND2_X1 U3968 ( .A1(n4509), .A2(U4043), .ZN(n3134) );
  OAI21_X1 U3969 ( .B1(U4043), .B2(n3135), .A(n3134), .ZN(U3569) );
  INV_X1 U3970 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n3137) );
  NAND2_X1 U3971 ( .A1(n3665), .A2(U4043), .ZN(n3136) );
  OAI21_X1 U3972 ( .B1(U4043), .B2(n3137), .A(n3136), .ZN(U3556) );
  INV_X1 U3973 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n3140) );
  NAND2_X1 U3974 ( .A1(n3138), .A2(U4043), .ZN(n3139) );
  OAI21_X1 U3975 ( .B1(U4043), .B2(n3140), .A(n3139), .ZN(U3573) );
  INV_X1 U3976 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n3142) );
  NAND2_X1 U3977 ( .A1(n4403), .A2(U4043), .ZN(n3141) );
  OAI21_X1 U3978 ( .B1(U4043), .B2(n3142), .A(n3141), .ZN(U3572) );
  INV_X1 U3979 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n3148) );
  INV_X1 U3980 ( .A(REG1_REG_31__SCAN_IN), .ZN(n3145) );
  NAND2_X1 U3981 ( .A1(n2423), .A2(REG2_REG_31__SCAN_IN), .ZN(n3144) );
  NAND2_X1 U3982 ( .A1(n2413), .A2(REG0_REG_31__SCAN_IN), .ZN(n3143) );
  OAI211_X1 U3983 ( .C1(n3146), .C2(n3145), .A(n3144), .B(n3143), .ZN(n4524)
         );
  NAND2_X1 U3984 ( .A1(n4524), .A2(U4043), .ZN(n3147) );
  OAI21_X1 U3985 ( .B1(U4043), .B2(n3148), .A(n3147), .ZN(U3581) );
  INV_X1 U3986 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n3150) );
  NAND2_X1 U3987 ( .A1(n3247), .A2(U4043), .ZN(n3149) );
  OAI21_X1 U3988 ( .B1(U4043), .B2(n3150), .A(n3149), .ZN(U3550) );
  INV_X1 U3989 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n3152) );
  NAND2_X1 U3990 ( .A1(n2790), .A2(U4043), .ZN(n3151) );
  OAI21_X1 U3991 ( .B1(U4043), .B2(n3152), .A(n3151), .ZN(U3551) );
  XNOR2_X1 U3992 ( .A(n4291), .B(n4633), .ZN(n4288) );
  XNOR2_X1 U3993 ( .A(n4288), .B(REG2_REG_8__SCAN_IN), .ZN(n3165) );
  NAND2_X1 U3994 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3608) );
  NOR2_X1 U3995 ( .A1(n3155), .A2(REG1_REG_7__SCAN_IN), .ZN(n3159) );
  OAI22_X1 U3996 ( .A1(n3159), .A2(n3158), .B1(n3157), .B2(n3156), .ZN(n4261)
         );
  XNOR2_X1 U3997 ( .A(n4261), .B(n4633), .ZN(n4264) );
  XNOR2_X1 U3998 ( .A(REG1_REG_8__SCAN_IN), .B(n4264), .ZN(n3160) );
  NAND2_X1 U3999 ( .A1(n4769), .A2(n3160), .ZN(n3161) );
  NAND2_X1 U4000 ( .A1(n3608), .A2(n3161), .ZN(n3162) );
  AOI21_X1 U4001 ( .B1(n4768), .B2(ADDR_REG_8__SCAN_IN), .A(n3162), .ZN(n3164)
         );
  NAND2_X1 U4002 ( .A1(n4256), .A2(n4633), .ZN(n3163) );
  OAI211_X1 U4003 ( .C1(n3165), .C2(n4762), .A(n3164), .B(n3163), .ZN(U3248)
         );
  INV_X1 U4004 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4789) );
  AOI21_X1 U4005 ( .B1(n4672), .B2(n4789), .A(n4654), .ZN(n4671) );
  NAND2_X1 U4006 ( .A1(n3166), .A2(n3168), .ZN(n3167) );
  OAI211_X1 U4007 ( .C1(n4241), .C2(n3168), .A(n3167), .B(n4218), .ZN(n3169)
         );
  OAI211_X1 U4008 ( .C1(IR_REG_0__SCAN_IN), .C2(n4671), .A(n3169), .B(U4043), 
        .ZN(n4260) );
  XNOR2_X1 U4009 ( .A(n3170), .B(REG2_REG_4__SCAN_IN), .ZN(n3178) );
  OAI211_X1 U4010 ( .C1(REG1_REG_4__SCAN_IN), .C2(n3172), .A(n4769), .B(n3171), 
        .ZN(n3175) );
  NAND2_X1 U4011 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3191) );
  INV_X1 U4012 ( .A(n3191), .ZN(n3173) );
  AOI21_X1 U4013 ( .B1(n4768), .B2(ADDR_REG_4__SCAN_IN), .A(n3173), .ZN(n3174)
         );
  OAI211_X1 U4014 ( .C1(n4775), .C2(n3176), .A(n3175), .B(n3174), .ZN(n3177)
         );
  AOI21_X1 U4015 ( .B1(n4711), .B2(n3178), .A(n3177), .ZN(n3179) );
  NAND2_X1 U4016 ( .A1(n4260), .A2(n3179), .ZN(U3244) );
  OAI21_X1 U4017 ( .B1(n3182), .B2(n3180), .A(n3181), .ZN(n3186) );
  AOI22_X1 U4018 ( .A1(n4054), .A2(n3229), .B1(n4059), .B2(n4236), .ZN(n3184)
         );
  MUX2_X1 U4019 ( .A(n4021), .B(STATE_REG_SCAN_IN), .S(REG3_REG_3__SCAN_IN), 
        .Z(n3183) );
  OAI211_X1 U4020 ( .C1(n3203), .C2(n4056), .A(n3184), .B(n3183), .ZN(n3185)
         );
  AOI21_X1 U4021 ( .B1(n3186), .B2(n3713), .A(n3185), .ZN(n3187) );
  INV_X1 U4022 ( .A(n3187), .ZN(U3215) );
  NAND2_X1 U4023 ( .A1(n3188), .A2(n3713), .ZN(n3197) );
  AOI21_X1 U4024 ( .B1(n3181), .B2(n3190), .A(n3189), .ZN(n3196) );
  AOI22_X1 U4025 ( .A1(n4054), .A2(n4233), .B1(n4053), .B2(n3285), .ZN(n3195)
         );
  OAI21_X1 U4026 ( .B1(n4043), .B2(n2431), .A(n3191), .ZN(n3192) );
  AOI21_X1 U4027 ( .B1(n3193), .B2(n4041), .A(n3192), .ZN(n3194) );
  OAI211_X1 U4028 ( .C1(n3197), .C2(n3196), .A(n3195), .B(n3194), .ZN(U3227)
         );
  NAND2_X1 U4029 ( .A1(n3198), .A2(n3199), .ZN(n3201) );
  INV_X1 U4030 ( .A(n3200), .ZN(n4141) );
  XNOR2_X1 U4031 ( .A(n3201), .B(n4141), .ZN(n3289) );
  XNOR2_X1 U4032 ( .A(n3202), .B(n4141), .ZN(n3206) );
  OAI22_X1 U4033 ( .A1(n2421), .A2(n4482), .B1(n4577), .B2(n3203), .ZN(n3204)
         );
  AOI21_X1 U4034 ( .B1(n4506), .B2(n4236), .A(n3204), .ZN(n3205) );
  OAI21_X1 U4035 ( .B1(n3206), .B2(n4486), .A(n3205), .ZN(n3290) );
  AOI21_X1 U4036 ( .B1(n4856), .B2(n3289), .A(n3290), .ZN(n3265) );
  INV_X1 U4037 ( .A(n3221), .ZN(n3208) );
  INV_X1 U4038 ( .A(n3207), .ZN(n3266) );
  AOI21_X1 U4039 ( .B1(n3209), .B2(n3208), .A(n3266), .ZN(n3292) );
  INV_X1 U4040 ( .A(n4585), .ZN(n4666) );
  AOI22_X1 U4041 ( .A1(n3292), .A2(n4666), .B1(REG1_REG_3__SCAN_IN), .B2(n4865), .ZN(n3210) );
  OAI21_X1 U4042 ( .B1(n3265), .B2(n4865), .A(n3210), .ZN(U3521) );
  OAI21_X1 U40430 ( .B1(n3211), .B2(n4145), .A(n3198), .ZN(n4777) );
  INV_X1 U4044 ( .A(n4777), .ZN(n3220) );
  XNOR2_X1 U4045 ( .A(n3213), .B(n3212), .ZN(n3219) );
  NAND2_X1 U4046 ( .A1(n4777), .A2(n4463), .ZN(n3217) );
  NOR2_X1 U4047 ( .A1(n3214), .A2(n4577), .ZN(n3215) );
  AOI21_X1 U4048 ( .B1(n2790), .B2(n4506), .A(n3215), .ZN(n3216) );
  OAI211_X1 U4049 ( .C1(n2431), .C2(n4482), .A(n3217), .B(n3216), .ZN(n3218)
         );
  AOI21_X1 U4050 ( .B1(n3219), .B2(n4514), .A(n3218), .ZN(n4780) );
  OAI21_X1 U4051 ( .B1(n3220), .B2(n4831), .A(n4780), .ZN(n4838) );
  INV_X1 U4052 ( .A(n4838), .ZN(n3224) );
  AOI21_X1 U4053 ( .B1(n3222), .B2(n3257), .A(n3221), .ZN(n4836) );
  AOI22_X1 U4054 ( .A1(n4836), .A2(n4666), .B1(REG1_REG_2__SCAN_IN), .B2(n4865), .ZN(n3223) );
  OAI21_X1 U4055 ( .B1(n3224), .B2(n4865), .A(n3223), .ZN(U3520) );
  XNOR2_X1 U4056 ( .A(n3226), .B(n3225), .ZN(n3232) );
  AOI22_X1 U4057 ( .A1(n4054), .A2(n3665), .B1(n4053), .B2(n3627), .ZN(n3231)
         );
  NOR2_X1 U4058 ( .A1(n4056), .A2(n3298), .ZN(n3227) );
  AOI211_X1 U4059 ( .C1(n4059), .C2(n3229), .A(n3228), .B(n3227), .ZN(n3230)
         );
  OAI211_X1 U4060 ( .C1(n3232), .C2(n4062), .A(n3231), .B(n3230), .ZN(U3224)
         );
  INV_X1 U4061 ( .A(n3234), .ZN(n3236) );
  NAND2_X1 U4062 ( .A1(n3236), .A2(n3235), .ZN(n3237) );
  XNOR2_X1 U4063 ( .A(n3233), .B(n3237), .ZN(n3242) );
  AOI22_X1 U4064 ( .A1(n4054), .A2(n3679), .B1(n4053), .B2(n3614), .ZN(n3241)
         );
  INV_X1 U4065 ( .A(n4233), .ZN(n3616) );
  OAI21_X1 U4066 ( .B1(n4043), .B2(n3616), .A(n3238), .ZN(n3239) );
  AOI21_X1 U4067 ( .B1(n3618), .B2(n4041), .A(n3239), .ZN(n3240) );
  OAI211_X1 U4068 ( .C1(n3242), .C2(n4062), .A(n3241), .B(n3240), .ZN(U3236)
         );
  OAI21_X1 U4069 ( .B1(n2705), .B2(n3244), .A(n3243), .ZN(n4832) );
  OAI21_X1 U4070 ( .B1(n3246), .B2(n4068), .A(n3245), .ZN(n3251) );
  AOI22_X1 U4071 ( .A1(n4236), .A2(n4508), .B1(n4658), .B2(n3256), .ZN(n3248)
         );
  OAI21_X1 U4072 ( .B1(n3249), .B2(n4578), .A(n3248), .ZN(n3250) );
  AOI21_X1 U4073 ( .B1(n3251), .B2(n4514), .A(n3250), .ZN(n3252) );
  OAI21_X1 U4074 ( .B1(n3842), .B2(n4832), .A(n3252), .ZN(n4834) );
  INV_X1 U4075 ( .A(n4834), .ZN(n3263) );
  INV_X1 U4076 ( .A(n4832), .ZN(n3261) );
  INV_X1 U4077 ( .A(n3253), .ZN(n3254) );
  NAND2_X1 U4078 ( .A1(n4517), .A2(n3254), .ZN(n4469) );
  INV_X1 U4079 ( .A(n4469), .ZN(n4786) );
  NAND2_X1 U4080 ( .A1(n3256), .A2(n3255), .ZN(n3258) );
  NAND2_X1 U4081 ( .A1(n3258), .A2(n3257), .ZN(n4830) );
  AOI22_X1 U4082 ( .A1(n4781), .A2(REG2_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(n4785), .ZN(n3259) );
  OAI21_X1 U4083 ( .B1(n4493), .B2(n4830), .A(n3259), .ZN(n3260) );
  AOI21_X1 U4084 ( .B1(n3261), .B2(n4786), .A(n3260), .ZN(n3262) );
  OAI21_X1 U4085 ( .B1(n3263), .B2(n4781), .A(n3262), .ZN(U3289) );
  INV_X1 U4086 ( .A(n4628), .ZN(n4837) );
  AOI22_X1 U4087 ( .A1(n3292), .A2(n4837), .B1(REG0_REG_3__SCAN_IN), .B2(n4858), .ZN(n3264) );
  OAI21_X1 U4088 ( .B1(n3265), .B2(n4858), .A(n3264), .ZN(U3473) );
  OAI211_X1 U4089 ( .C1(n3266), .C2(n3271), .A(n4829), .B(n3302), .ZN(n4841)
         );
  NOR2_X1 U4090 ( .A1(n4841), .A2(n4516), .ZN(n3284) );
  INV_X1 U4091 ( .A(n3267), .ZN(n3268) );
  XOR2_X1 U4092 ( .A(n3269), .B(n3268), .Z(n3283) );
  NAND2_X1 U4093 ( .A1(n4234), .A2(n4506), .ZN(n3270) );
  OAI21_X1 U4094 ( .B1(n4577), .B2(n3271), .A(n3270), .ZN(n3281) );
  AND2_X1 U4095 ( .A1(n3273), .A2(n3272), .ZN(n3279) );
  NAND2_X1 U4096 ( .A1(n3198), .A2(n3274), .ZN(n3276) );
  AND2_X1 U4097 ( .A1(n3276), .A2(n3275), .ZN(n3277) );
  NAND2_X1 U4098 ( .A1(n3277), .A2(n3268), .ZN(n3278) );
  NAND2_X1 U4099 ( .A1(n3279), .A2(n3278), .ZN(n3286) );
  NOR2_X1 U4100 ( .A1(n3286), .A2(n3842), .ZN(n3280) );
  AOI211_X1 U4101 ( .C1(n4508), .C2(n4233), .A(n3281), .B(n3280), .ZN(n3282)
         );
  OAI21_X1 U4102 ( .B1(n4486), .B2(n3283), .A(n3282), .ZN(n4842) );
  AOI211_X1 U4103 ( .C1(n4785), .C2(n3285), .A(n3284), .B(n4842), .ZN(n3288)
         );
  INV_X1 U4104 ( .A(n3286), .ZN(n4845) );
  AOI22_X1 U4105 ( .A1(n4845), .A2(n4786), .B1(REG2_REG_4__SCAN_IN), .B2(n4781), .ZN(n3287) );
  OAI21_X1 U4106 ( .B1(n3288), .B2(n4781), .A(n3287), .ZN(U3286) );
  INV_X1 U4107 ( .A(n3289), .ZN(n3295) );
  NAND2_X1 U4108 ( .A1(n3290), .A2(n4517), .ZN(n3294) );
  OAI22_X1 U4109 ( .A1(n4517), .A2(n3544), .B1(REG3_REG_3__SCAN_IN), .B2(n4420), .ZN(n3291) );
  AOI21_X1 U4110 ( .B1(n3292), .B2(n4776), .A(n3291), .ZN(n3293) );
  OAI211_X1 U4111 ( .C1(n4521), .C2(n3295), .A(n3294), .B(n3293), .ZN(U3287)
         );
  INV_X1 U4112 ( .A(n3297), .ZN(n4077) );
  AND2_X1 U4113 ( .A1(n4077), .A2(n4090), .ZN(n4144) );
  XNOR2_X1 U4114 ( .A(n3296), .B(n4144), .ZN(n3635) );
  OAI22_X1 U4115 ( .A1(n2421), .A2(n4578), .B1(n4577), .B2(n3298), .ZN(n3301)
         );
  XNOR2_X1 U4116 ( .A(n3299), .B(n4144), .ZN(n3300) );
  INV_X1 U4117 ( .A(n3665), .ZN(n3311) );
  OAI22_X1 U4118 ( .A1(n3300), .A2(n4486), .B1(n3311), .B2(n4482), .ZN(n3625)
         );
  AOI211_X1 U4119 ( .C1(n3635), .C2(n4856), .A(n3301), .B(n3625), .ZN(n3306)
         );
  AND2_X1 U4120 ( .A1(n3302), .A2(n3631), .ZN(n3303) );
  NOR2_X1 U4121 ( .A1(n3596), .A2(n3303), .ZN(n3626) );
  AOI22_X1 U4122 ( .A1(n3626), .A2(n4837), .B1(REG0_REG_5__SCAN_IN), .B2(n4858), .ZN(n3304) );
  OAI21_X1 U4123 ( .B1(n3306), .B2(n4858), .A(n3304), .ZN(U3477) );
  AOI22_X1 U4124 ( .A1(n3626), .A2(n4666), .B1(REG1_REG_5__SCAN_IN), .B2(n4865), .ZN(n3305) );
  OAI21_X1 U4125 ( .B1(n3306), .B2(n4865), .A(n3305), .ZN(U3523) );
  OAI21_X1 U4126 ( .B1(n3308), .B2(n3307), .A(n3713), .ZN(n3316) );
  INV_X1 U4127 ( .A(n3695), .ZN(n3740) );
  OAI22_X1 U4128 ( .A1(n3740), .A2(n4022), .B1(n4021), .B2(n3671), .ZN(n3313)
         );
  OAI21_X1 U4129 ( .B1(n4043), .B2(n3311), .A(n3310), .ZN(n3312) );
  AOI211_X1 U4130 ( .C1(n3314), .C2(n4041), .A(n3313), .B(n3312), .ZN(n3315)
         );
  OAI21_X1 U4131 ( .B1(n3316), .B2(n3309), .A(n3315), .ZN(n3590) );
  NOR2_X1 U4132 ( .A1(keyinput22), .A2(keyinput23), .ZN(n3317) );
  NAND3_X1 U4133 ( .A1(keyinput103), .A2(keyinput105), .A3(n3317), .ZN(n3332)
         );
  NAND4_X1 U4134 ( .A1(keyinput12), .A2(keyinput21), .A3(keyinput94), .A4(
        keyinput95), .ZN(n3331) );
  NOR2_X1 U4135 ( .A1(keyinput126), .A2(keyinput11), .ZN(n3318) );
  NAND3_X1 U4136 ( .A1(keyinput42), .A2(keyinput124), .A3(n3318), .ZN(n3319)
         );
  NOR3_X1 U4137 ( .A1(keyinput91), .A2(keyinput41), .A3(n3319), .ZN(n3320) );
  NAND3_X1 U4138 ( .A1(keyinput111), .A2(keyinput88), .A3(n3320), .ZN(n3330)
         );
  INV_X1 U4139 ( .A(keyinput78), .ZN(n3321) );
  NOR4_X1 U4140 ( .A1(keyinput65), .A2(keyinput7), .A3(keyinput10), .A4(n3321), 
        .ZN(n3328) );
  NAND2_X1 U4141 ( .A1(keyinput53), .A2(keyinput29), .ZN(n3322) );
  NOR3_X1 U4142 ( .A1(keyinput85), .A2(keyinput83), .A3(n3322), .ZN(n3327) );
  NAND2_X1 U4143 ( .A1(keyinput122), .A2(keyinput6), .ZN(n3323) );
  NOR3_X1 U4144 ( .A1(keyinput80), .A2(keyinput24), .A3(n3323), .ZN(n3326) );
  INV_X1 U4145 ( .A(keyinput27), .ZN(n3324) );
  NOR4_X1 U4146 ( .A1(keyinput62), .A2(keyinput108), .A3(keyinput84), .A4(
        n3324), .ZN(n3325) );
  NAND4_X1 U4147 ( .A1(n3328), .A2(n3327), .A3(n3326), .A4(n3325), .ZN(n3329)
         );
  NOR4_X1 U4148 ( .A1(n3332), .A2(n3331), .A3(n3330), .A4(n3329), .ZN(n3379)
         );
  NOR2_X1 U4149 ( .A1(keyinput60), .A2(keyinput3), .ZN(n3333) );
  NAND3_X1 U4150 ( .A1(keyinput52), .A2(keyinput90), .A3(n3333), .ZN(n3377) );
  INV_X1 U4151 ( .A(keyinput89), .ZN(n3571) );
  NAND4_X1 U4152 ( .A1(keyinput121), .A2(keyinput102), .A3(keyinput40), .A4(
        n3571), .ZN(n3376) );
  NAND2_X1 U4153 ( .A1(keyinput73), .A2(keyinput113), .ZN(n3334) );
  NOR3_X1 U4154 ( .A1(keyinput37), .A2(keyinput49), .A3(n3334), .ZN(n3342) );
  INV_X1 U4155 ( .A(keyinput31), .ZN(n3530) );
  INV_X1 U4156 ( .A(keyinput107), .ZN(n3531) );
  INV_X1 U4157 ( .A(keyinput92), .ZN(n3528) );
  AND4_X1 U4158 ( .A1(n3530), .A2(n3531), .A3(n3528), .A4(keyinput77), .ZN(
        n3341) );
  INV_X1 U4159 ( .A(keyinput72), .ZN(n3335) );
  NOR4_X1 U4160 ( .A1(keyinput48), .A2(keyinput25), .A3(keyinput112), .A4(
        n3335), .ZN(n3336) );
  NAND4_X1 U4161 ( .A1(keyinput34), .A2(keyinput35), .A3(keyinput8), .A4(n3336), .ZN(n3339) );
  NOR4_X1 U4162 ( .A1(keyinput39), .A2(keyinput51), .A3(keyinput98), .A4(
        keyinput17), .ZN(n3337) );
  NAND3_X1 U4163 ( .A1(keyinput63), .A2(keyinput70), .A3(n3337), .ZN(n3338) );
  NOR4_X1 U4164 ( .A1(keyinput30), .A2(keyinput32), .A3(n3339), .A4(n3338), 
        .ZN(n3340) );
  NAND3_X1 U4165 ( .A1(n3342), .A2(n3341), .A3(n3340), .ZN(n3375) );
  AND4_X1 U4166 ( .A1(keyinput1), .A2(keyinput15), .A3(keyinput119), .A4(
        keyinput13), .ZN(n3373) );
  NAND2_X1 U4167 ( .A1(keyinput100), .A2(keyinput96), .ZN(n3343) );
  NOR3_X1 U4168 ( .A1(keyinput86), .A2(keyinput55), .A3(n3343), .ZN(n3372) );
  NAND2_X1 U4169 ( .A1(keyinput82), .A2(keyinput28), .ZN(n3344) );
  NOR3_X1 U4170 ( .A1(keyinput81), .A2(keyinput93), .A3(n3344), .ZN(n3345) );
  NAND3_X1 U4171 ( .A1(keyinput110), .A2(keyinput123), .A3(n3345), .ZN(n3354)
         );
  NAND2_X1 U4172 ( .A1(keyinput75), .A2(keyinput99), .ZN(n3346) );
  NOR3_X1 U4173 ( .A1(keyinput45), .A2(keyinput56), .A3(n3346), .ZN(n3352) );
  NAND2_X1 U4174 ( .A1(keyinput87), .A2(keyinput61), .ZN(n3347) );
  NOR3_X1 U4175 ( .A1(keyinput127), .A2(keyinput57), .A3(n3347), .ZN(n3351) );
  NAND2_X1 U4176 ( .A1(keyinput69), .A2(keyinput54), .ZN(n3348) );
  NOR3_X1 U4177 ( .A1(keyinput14), .A2(keyinput64), .A3(n3348), .ZN(n3350) );
  NOR4_X1 U4178 ( .A1(keyinput101), .A2(keyinput106), .A3(keyinput74), .A4(
        keyinput44), .ZN(n3349) );
  NAND4_X1 U4179 ( .A1(n3352), .A2(n3351), .A3(n3350), .A4(n3349), .ZN(n3353)
         );
  NOR4_X1 U4180 ( .A1(keyinput0), .A2(keyinput120), .A3(n3354), .A4(n3353), 
        .ZN(n3371) );
  NAND2_X1 U4181 ( .A1(keyinput4), .A2(keyinput16), .ZN(n3355) );
  NOR3_X1 U4182 ( .A1(keyinput36), .A2(keyinput125), .A3(n3355), .ZN(n3356) );
  NAND3_X1 U4183 ( .A1(keyinput76), .A2(keyinput68), .A3(n3356), .ZN(n3369) );
  NOR2_X1 U4184 ( .A1(keyinput18), .A2(keyinput43), .ZN(n3357) );
  NAND3_X1 U4185 ( .A1(keyinput19), .A2(keyinput38), .A3(n3357), .ZN(n3358) );
  NOR3_X1 U4186 ( .A1(keyinput2), .A2(keyinput59), .A3(n3358), .ZN(n3367) );
  NOR2_X1 U4187 ( .A1(keyinput71), .A2(keyinput58), .ZN(n3359) );
  NAND3_X1 U4188 ( .A1(keyinput50), .A2(keyinput104), .A3(n3359), .ZN(n3365)
         );
  NOR2_X1 U4189 ( .A1(keyinput116), .A2(keyinput33), .ZN(n3360) );
  NAND3_X1 U4190 ( .A1(keyinput20), .A2(keyinput26), .A3(n3360), .ZN(n3364) );
  NAND4_X1 U4191 ( .A1(keyinput9), .A2(keyinput79), .A3(keyinput118), .A4(
        keyinput115), .ZN(n3363) );
  NOR3_X1 U4192 ( .A1(keyinput97), .A2(keyinput66), .A3(keyinput5), .ZN(n3361)
         );
  NAND2_X1 U4193 ( .A1(keyinput67), .A2(n3361), .ZN(n3362) );
  NOR4_X1 U4194 ( .A1(n3365), .A2(n3364), .A3(n3363), .A4(n3362), .ZN(n3366)
         );
  NAND4_X1 U4195 ( .A1(keyinput46), .A2(keyinput47), .A3(n3367), .A4(n3366), 
        .ZN(n3368) );
  NOR4_X1 U4196 ( .A1(keyinput117), .A2(keyinput109), .A3(n3369), .A4(n3368), 
        .ZN(n3370) );
  NAND4_X1 U4197 ( .A1(n3373), .A2(n3372), .A3(n3371), .A4(n3370), .ZN(n3374)
         );
  NOR4_X1 U4198 ( .A1(n3377), .A2(n3376), .A3(n3375), .A4(n3374), .ZN(n3378)
         );
  AOI21_X1 U4199 ( .B1(n3379), .B2(n3378), .A(keyinput114), .ZN(n3588) );
  INV_X1 U4200 ( .A(REG0_REG_21__SCAN_IN), .ZN(n3382) );
  INV_X1 U4201 ( .A(REG2_REG_21__SCAN_IN), .ZN(n3381) );
  AOI22_X1 U4202 ( .A1(n3382), .A2(keyinput96), .B1(keyinput1), .B2(n3381), 
        .ZN(n3380) );
  OAI221_X1 U4203 ( .B1(n3382), .B2(keyinput96), .C1(n3381), .C2(keyinput1), 
        .A(n3380), .ZN(n3393) );
  INV_X1 U4204 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4555) );
  INV_X1 U4205 ( .A(keyinput15), .ZN(n3384) );
  AOI22_X1 U4206 ( .A1(n4555), .A2(keyinput119), .B1(DATAO_REG_22__SCAN_IN), 
        .B2(n3384), .ZN(n3383) );
  OAI221_X1 U4207 ( .B1(n4555), .B2(keyinput119), .C1(n3384), .C2(
        DATAO_REG_22__SCAN_IN), .A(n3383), .ZN(n3392) );
  INV_X1 U4208 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4614) );
  INV_X1 U4209 ( .A(keyinput55), .ZN(n3386) );
  AOI22_X1 U4210 ( .A1(n4614), .A2(keyinput13), .B1(DATAO_REG_23__SCAN_IN), 
        .B2(n3386), .ZN(n3385) );
  OAI221_X1 U4211 ( .B1(n4614), .B2(keyinput13), .C1(n3386), .C2(
        DATAO_REG_23__SCAN_IN), .A(n3385), .ZN(n3391) );
  INV_X1 U4212 ( .A(REG1_REG_23__SCAN_IN), .ZN(n3389) );
  INV_X1 U4213 ( .A(REG0_REG_23__SCAN_IN), .ZN(n3388) );
  AOI22_X1 U4214 ( .A1(n3389), .A2(keyinput100), .B1(n3388), .B2(keyinput61), 
        .ZN(n3387) );
  OAI221_X1 U4215 ( .B1(n3389), .B2(keyinput100), .C1(n3388), .C2(keyinput61), 
        .A(n3387), .ZN(n3390) );
  NOR4_X1 U4216 ( .A1(n3393), .A2(n3392), .A3(n3391), .A4(n3390), .ZN(n3426)
         );
  INV_X1 U4217 ( .A(REG0_REG_25__SCAN_IN), .ZN(n3395) );
  AOI22_X1 U4218 ( .A1(n4547), .A2(keyinput127), .B1(n3395), .B2(keyinput87), 
        .ZN(n3394) );
  OAI221_X1 U4219 ( .B1(n4547), .B2(keyinput127), .C1(n3395), .C2(keyinput87), 
        .A(n3394), .ZN(n3403) );
  AOI22_X1 U4220 ( .A1(n4536), .A2(keyinput57), .B1(n4532), .B2(keyinput99), 
        .ZN(n3396) );
  OAI221_X1 U4221 ( .B1(n4536), .B2(keyinput57), .C1(n4532), .C2(keyinput99), 
        .A(n3396), .ZN(n3402) );
  AOI22_X1 U4222 ( .A1(n2767), .A2(keyinput56), .B1(keyinput45), .B2(n2771), 
        .ZN(n3397) );
  OAI221_X1 U4223 ( .B1(n2767), .B2(keyinput56), .C1(n2771), .C2(keyinput45), 
        .A(n3397), .ZN(n3401) );
  INV_X1 U4224 ( .A(keyinput75), .ZN(n3399) );
  AOI22_X1 U4225 ( .A1(n3145), .A2(keyinput101), .B1(DATAO_REG_31__SCAN_IN), 
        .B2(n3399), .ZN(n3398) );
  OAI221_X1 U4226 ( .B1(n3145), .B2(keyinput101), .C1(n3399), .C2(
        DATAO_REG_31__SCAN_IN), .A(n3398), .ZN(n3400) );
  NOR4_X1 U4227 ( .A1(n3403), .A2(n3402), .A3(n3401), .A4(n3400), .ZN(n3425)
         );
  INV_X1 U4228 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4827) );
  INV_X1 U4229 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4840) );
  AOI22_X1 U4230 ( .A1(n4827), .A2(keyinput106), .B1(n4840), .B2(keyinput74), 
        .ZN(n3404) );
  OAI221_X1 U4231 ( .B1(n4827), .B2(keyinput106), .C1(n4840), .C2(keyinput74), 
        .A(n3404), .ZN(n3414) );
  INV_X1 U4232 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4846) );
  INV_X1 U4233 ( .A(DATAI_6_), .ZN(n3406) );
  AOI22_X1 U4234 ( .A1(n4846), .A2(keyinput54), .B1(n3406), .B2(keyinput64), 
        .ZN(n3405) );
  OAI221_X1 U4235 ( .B1(n4846), .B2(keyinput54), .C1(n3406), .C2(keyinput64), 
        .A(n3405), .ZN(n3413) );
  XOR2_X1 U4236 ( .A(n3407), .B(keyinput44), .Z(n3411) );
  XNOR2_X1 U4237 ( .A(IR_REG_3__SCAN_IN), .B(keyinput14), .ZN(n3410) );
  XNOR2_X1 U4238 ( .A(REG3_REG_7__SCAN_IN), .B(keyinput28), .ZN(n3409) );
  XNOR2_X1 U4239 ( .A(IR_REG_28__SCAN_IN), .B(keyinput69), .ZN(n3408) );
  NAND4_X1 U4240 ( .A1(n3411), .A2(n3410), .A3(n3409), .A4(n3408), .ZN(n3412)
         );
  NOR3_X1 U4241 ( .A1(n3414), .A2(n3413), .A3(n3412), .ZN(n3424) );
  AOI22_X1 U4242 ( .A1(n4800), .A2(keyinput93), .B1(keyinput81), .B2(n4804), 
        .ZN(n3415) );
  OAI221_X1 U4243 ( .B1(n4800), .B2(keyinput93), .C1(n4804), .C2(keyinput81), 
        .A(n3415), .ZN(n3422) );
  AOI22_X1 U4244 ( .A1(n4798), .A2(keyinput82), .B1(keyinput110), .B2(n4792), 
        .ZN(n3416) );
  OAI221_X1 U4245 ( .B1(n4798), .B2(keyinput82), .C1(n4792), .C2(keyinput110), 
        .A(n3416), .ZN(n3421) );
  INV_X1 U4246 ( .A(D_REG_23__SCAN_IN), .ZN(n4795) );
  INV_X1 U4247 ( .A(D_REG_22__SCAN_IN), .ZN(n4796) );
  AOI22_X1 U4248 ( .A1(n4795), .A2(keyinput123), .B1(keyinput0), .B2(n4796), 
        .ZN(n3417) );
  OAI221_X1 U4249 ( .B1(n4795), .B2(keyinput123), .C1(n4796), .C2(keyinput0), 
        .A(n3417), .ZN(n3420) );
  INV_X1 U4250 ( .A(D_REG_9__SCAN_IN), .ZN(n4802) );
  INV_X1 U4251 ( .A(D_REG_18__SCAN_IN), .ZN(n4799) );
  AOI22_X1 U4252 ( .A1(n4802), .A2(keyinput120), .B1(keyinput116), .B2(n4799), 
        .ZN(n3418) );
  OAI221_X1 U4253 ( .B1(n4802), .B2(keyinput120), .C1(n4799), .C2(keyinput116), 
        .A(n3418), .ZN(n3419) );
  NOR4_X1 U4254 ( .A1(n3422), .A2(n3421), .A3(n3420), .A4(n3419), .ZN(n3423)
         );
  NAND4_X1 U4255 ( .A1(n3426), .A2(n3425), .A3(n3424), .A4(n3423), .ZN(n3586)
         );
  INV_X1 U4256 ( .A(D_REG_26__SCAN_IN), .ZN(n4794) );
  INV_X1 U4257 ( .A(D_REG_5__SCAN_IN), .ZN(n4803) );
  AOI22_X1 U4258 ( .A1(n4794), .A2(keyinput20), .B1(keyinput33), .B2(n4803), 
        .ZN(n3427) );
  OAI221_X1 U4259 ( .B1(n4794), .B2(keyinput20), .C1(n4803), .C2(keyinput33), 
        .A(n3427), .ZN(n3436) );
  INV_X1 U4260 ( .A(D_REG_10__SCAN_IN), .ZN(n4801) );
  INV_X1 U4261 ( .A(D_REG_27__SCAN_IN), .ZN(n4793) );
  AOI22_X1 U4262 ( .A1(n4801), .A2(keyinput26), .B1(keyinput50), .B2(n4793), 
        .ZN(n3428) );
  OAI221_X1 U4263 ( .B1(n4801), .B2(keyinput26), .C1(n4793), .C2(keyinput50), 
        .A(n3428), .ZN(n3435) );
  INV_X1 U4264 ( .A(D_REG_31__SCAN_IN), .ZN(n4791) );
  INV_X1 U4265 ( .A(D_REG_21__SCAN_IN), .ZN(n4797) );
  AOI22_X1 U4266 ( .A1(n4791), .A2(keyinput58), .B1(keyinput71), .B2(n4797), 
        .ZN(n3429) );
  OAI221_X1 U4267 ( .B1(n4791), .B2(keyinput58), .C1(n4797), .C2(keyinput71), 
        .A(n3429), .ZN(n3434) );
  AOI22_X1 U4268 ( .A1(n3432), .A2(keyinput104), .B1(n3431), .B2(keyinput76), 
        .ZN(n3430) );
  OAI221_X1 U4269 ( .B1(n3432), .B2(keyinput104), .C1(n3431), .C2(keyinput76), 
        .A(n3430), .ZN(n3433) );
  NOR4_X1 U4270 ( .A1(n3436), .A2(n3435), .A3(n3434), .A4(n3433), .ZN(n3471)
         );
  AOI22_X1 U4271 ( .A1(n2684), .A2(keyinput125), .B1(keyinput117), .B2(n3438), 
        .ZN(n3437) );
  OAI221_X1 U4272 ( .B1(n2684), .B2(keyinput125), .C1(n3438), .C2(keyinput117), 
        .A(n3437), .ZN(n3447) );
  INV_X1 U4273 ( .A(DATAI_23_), .ZN(n4808) );
  INV_X1 U4274 ( .A(ADDR_REG_18__SCAN_IN), .ZN(n3440) );
  AOI22_X1 U4275 ( .A1(n4808), .A2(keyinput16), .B1(keyinput4), .B2(n3440), 
        .ZN(n3439) );
  OAI221_X1 U4276 ( .B1(n4808), .B2(keyinput16), .C1(n3440), .C2(keyinput4), 
        .A(n3439), .ZN(n3446) );
  INV_X1 U4277 ( .A(DATAI_17_), .ZN(n4809) );
  XOR2_X1 U4278 ( .A(n4809), .B(keyinput36), .Z(n3444) );
  XNOR2_X1 U4279 ( .A(IR_REG_12__SCAN_IN), .B(keyinput68), .ZN(n3443) );
  XNOR2_X1 U4280 ( .A(DATAI_28_), .B(keyinput97), .ZN(n3442) );
  XNOR2_X1 U4281 ( .A(IR_REG_9__SCAN_IN), .B(keyinput109), .ZN(n3441) );
  NAND4_X1 U4282 ( .A1(n3444), .A2(n3443), .A3(n3442), .A4(n3441), .ZN(n3445)
         );
  NOR3_X1 U4283 ( .A1(n3447), .A2(n3446), .A3(n3445), .ZN(n3470) );
  INV_X1 U4284 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3832) );
  INV_X1 U4285 ( .A(IR_REG_30__SCAN_IN), .ZN(n3934) );
  AOI22_X1 U4286 ( .A1(n3832), .A2(keyinput79), .B1(n3934), .B2(keyinput67), 
        .ZN(n3448) );
  OAI221_X1 U4287 ( .B1(n3832), .B2(keyinput79), .C1(n3934), .C2(keyinput67), 
        .A(n3448), .ZN(n3456) );
  XNOR2_X1 U4288 ( .A(keyinput9), .B(n2369), .ZN(n3455) );
  XNOR2_X1 U4289 ( .A(keyinput46), .B(n3932), .ZN(n3454) );
  XNOR2_X1 U4290 ( .A(DATAI_26_), .B(keyinput118), .ZN(n3452) );
  XNOR2_X1 U4291 ( .A(IR_REG_16__SCAN_IN), .B(keyinput5), .ZN(n3451) );
  XNOR2_X1 U4292 ( .A(IR_REG_22__SCAN_IN), .B(keyinput115), .ZN(n3450) );
  XNOR2_X1 U4293 ( .A(IR_REG_4__SCAN_IN), .B(keyinput66), .ZN(n3449) );
  NAND4_X1 U4294 ( .A1(n3452), .A2(n3451), .A3(n3450), .A4(n3449), .ZN(n3453)
         );
  NOR4_X1 U4295 ( .A1(n3456), .A2(n3455), .A3(n3454), .A4(n3453), .ZN(n3469)
         );
  AOI22_X1 U4296 ( .A1(n3458), .A2(keyinput19), .B1(keyinput43), .B2(n2396), 
        .ZN(n3457) );
  OAI221_X1 U4297 ( .B1(n3458), .B2(keyinput19), .C1(n2396), .C2(keyinput43), 
        .A(n3457), .ZN(n3467) );
  INV_X1 U4298 ( .A(REG3_REG_10__SCAN_IN), .ZN(n3717) );
  AOI22_X1 U4299 ( .A1(n3460), .A2(keyinput34), .B1(n3717), .B2(keyinput38), 
        .ZN(n3459) );
  OAI221_X1 U4300 ( .B1(n3460), .B2(keyinput34), .C1(n3717), .C2(keyinput38), 
        .A(n3459), .ZN(n3466) );
  XNOR2_X1 U4301 ( .A(DATAI_22_), .B(keyinput47), .ZN(n3464) );
  XNOR2_X1 U4302 ( .A(IR_REG_25__SCAN_IN), .B(keyinput2), .ZN(n3463) );
  XNOR2_X1 U4303 ( .A(REG3_REG_6__SCAN_IN), .B(keyinput59), .ZN(n3462) );
  XNOR2_X1 U4304 ( .A(DATAI_14_), .B(keyinput18), .ZN(n3461) );
  NAND4_X1 U4305 ( .A1(n3464), .A2(n3463), .A3(n3462), .A4(n3461), .ZN(n3465)
         );
  NOR3_X1 U4306 ( .A1(n3467), .A2(n3466), .A3(n3465), .ZN(n3468) );
  NAND4_X1 U4307 ( .A1(n3471), .A2(n3470), .A3(n3469), .A4(n3468), .ZN(n3585)
         );
  INV_X1 U4308 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4721) );
  AOI22_X1 U4309 ( .A1(n4721), .A2(keyinput29), .B1(keyinput53), .B2(n4789), 
        .ZN(n3472) );
  OAI221_X1 U4310 ( .B1(n4721), .B2(keyinput29), .C1(n4789), .C2(keyinput53), 
        .A(n3472), .ZN(n3480) );
  INV_X1 U4311 ( .A(REG2_REG_11__SCAN_IN), .ZN(n4284) );
  AOI22_X1 U4312 ( .A1(n4284), .A2(keyinput7), .B1(keyinput65), .B2(n2436), 
        .ZN(n3473) );
  OAI221_X1 U4313 ( .B1(n4284), .B2(keyinput7), .C1(n2436), .C2(keyinput65), 
        .A(n3473), .ZN(n3479) );
  INV_X1 U4314 ( .A(REG2_REG_9__SCAN_IN), .ZN(n4286) );
  XOR2_X1 U4315 ( .A(n4286), .B(keyinput78), .Z(n3477) );
  XNOR2_X1 U4316 ( .A(REG2_REG_1__SCAN_IN), .B(keyinput83), .ZN(n3476) );
  XNOR2_X1 U4317 ( .A(IR_REG_15__SCAN_IN), .B(keyinput10), .ZN(n3475) );
  XNOR2_X1 U4318 ( .A(REG1_REG_14__SCAN_IN), .B(keyinput111), .ZN(n3474) );
  NAND4_X1 U4319 ( .A1(n3477), .A2(n3476), .A3(n3475), .A4(n3474), .ZN(n3478)
         );
  NOR3_X1 U4320 ( .A1(n3480), .A2(n3479), .A3(n3478), .ZN(n3525) );
  INV_X1 U4321 ( .A(keyinput103), .ZN(n3483) );
  INV_X1 U4322 ( .A(keyinput105), .ZN(n3482) );
  AOI22_X1 U4323 ( .A1(n3483), .A2(ADDR_REG_7__SCAN_IN), .B1(
        ADDR_REG_8__SCAN_IN), .B2(n3482), .ZN(n3481) );
  OAI221_X1 U4324 ( .B1(n3483), .B2(ADDR_REG_7__SCAN_IN), .C1(n3482), .C2(
        ADDR_REG_8__SCAN_IN), .A(n3481), .ZN(n3495) );
  INV_X1 U4325 ( .A(keyinput22), .ZN(n3485) );
  AOI22_X1 U4326 ( .A1(n4826), .A2(keyinput21), .B1(ADDR_REG_6__SCAN_IN), .B2(
        n3485), .ZN(n3484) );
  OAI221_X1 U4327 ( .B1(n4826), .B2(keyinput21), .C1(n3485), .C2(
        ADDR_REG_6__SCAN_IN), .A(n3484), .ZN(n3494) );
  INV_X1 U4328 ( .A(keyinput95), .ZN(n3488) );
  INV_X1 U4329 ( .A(keyinput85), .ZN(n3487) );
  AOI22_X1 U4330 ( .A1(n3488), .A2(ADDR_REG_13__SCAN_IN), .B1(
        ADDR_REG_15__SCAN_IN), .B2(n3487), .ZN(n3486) );
  OAI221_X1 U4331 ( .B1(n3488), .B2(ADDR_REG_13__SCAN_IN), .C1(n3487), .C2(
        ADDR_REG_15__SCAN_IN), .A(n3486), .ZN(n3493) );
  INV_X1 U4332 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3491) );
  INV_X1 U4333 ( .A(keyinput94), .ZN(n3490) );
  AOI22_X1 U4334 ( .A1(n3491), .A2(keyinput23), .B1(ADDR_REG_10__SCAN_IN), 
        .B2(n3490), .ZN(n3489) );
  OAI221_X1 U4335 ( .B1(n3491), .B2(keyinput23), .C1(n3490), .C2(
        ADDR_REG_10__SCAN_IN), .A(n3489), .ZN(n3492) );
  NOR4_X1 U4336 ( .A1(n3495), .A2(n3494), .A3(n3493), .A4(n3492), .ZN(n3524)
         );
  INV_X1 U4337 ( .A(REG0_REG_18__SCAN_IN), .ZN(n3498) );
  INV_X1 U4338 ( .A(keyinput80), .ZN(n3497) );
  AOI22_X1 U4339 ( .A1(n3498), .A2(keyinput84), .B1(DATAO_REG_19__SCAN_IN), 
        .B2(n3497), .ZN(n3496) );
  OAI221_X1 U4340 ( .B1(n3498), .B2(keyinput84), .C1(n3497), .C2(
        DATAO_REG_19__SCAN_IN), .A(n3496), .ZN(n3509) );
  INV_X1 U4341 ( .A(keyinput108), .ZN(n3500) );
  AOI22_X1 U4342 ( .A1(n2560), .A2(keyinput62), .B1(DATAO_REG_17__SCAN_IN), 
        .B2(n3500), .ZN(n3499) );
  OAI221_X1 U4343 ( .B1(n2560), .B2(keyinput62), .C1(n3500), .C2(
        DATAO_REG_17__SCAN_IN), .A(n3499), .ZN(n3508) );
  INV_X1 U4344 ( .A(keyinput122), .ZN(n3502) );
  AOI22_X1 U4345 ( .A1(n4562), .A2(keyinput86), .B1(DATAO_REG_21__SCAN_IN), 
        .B2(n3502), .ZN(n3501) );
  OAI221_X1 U4346 ( .B1(n4562), .B2(keyinput86), .C1(n3502), .C2(
        DATAO_REG_21__SCAN_IN), .A(n3501), .ZN(n3507) );
  INV_X1 U4347 ( .A(REG0_REG_19__SCAN_IN), .ZN(n3505) );
  INV_X1 U4348 ( .A(keyinput24), .ZN(n3504) );
  AOI22_X1 U4349 ( .A1(n3505), .A2(keyinput6), .B1(DATAO_REG_20__SCAN_IN), 
        .B2(n3504), .ZN(n3503) );
  OAI221_X1 U4350 ( .B1(n3505), .B2(keyinput6), .C1(n3504), .C2(
        DATAO_REG_20__SCAN_IN), .A(n3503), .ZN(n3506) );
  NOR4_X1 U4351 ( .A1(n3509), .A2(n3508), .A3(n3507), .A4(n3506), .ZN(n3523)
         );
  INV_X1 U4352 ( .A(DATAI_9_), .ZN(n4823) );
  AOI22_X1 U4353 ( .A1(n2513), .A2(keyinput42), .B1(keyinput91), .B2(n4823), 
        .ZN(n3510) );
  OAI221_X1 U4354 ( .B1(n2513), .B2(keyinput42), .C1(n4823), .C2(keyinput91), 
        .A(n3510), .ZN(n3521) );
  INV_X1 U4355 ( .A(DATAI_13_), .ZN(n4817) );
  INV_X1 U4356 ( .A(REG0_REG_15__SCAN_IN), .ZN(n3512) );
  AOI22_X1 U4357 ( .A1(n4817), .A2(keyinput41), .B1(n3512), .B2(keyinput11), 
        .ZN(n3511) );
  OAI221_X1 U4358 ( .B1(n4817), .B2(keyinput41), .C1(n3512), .C2(keyinput11), 
        .A(n3511), .ZN(n3520) );
  INV_X1 U4359 ( .A(REG0_REG_16__SCAN_IN), .ZN(n3514) );
  AOI22_X1 U4360 ( .A1(n3515), .A2(keyinput124), .B1(n3514), .B2(keyinput27), 
        .ZN(n3513) );
  OAI221_X1 U4361 ( .B1(n3515), .B2(keyinput124), .C1(n3514), .C2(keyinput27), 
        .A(n3513), .ZN(n3519) );
  XNOR2_X1 U4362 ( .A(REG0_REG_14__SCAN_IN), .B(keyinput88), .ZN(n3517) );
  XNOR2_X1 U4363 ( .A(IR_REG_11__SCAN_IN), .B(keyinput126), .ZN(n3516) );
  NAND2_X1 U4364 ( .A1(n3517), .A2(n3516), .ZN(n3518) );
  NOR4_X1 U4365 ( .A1(n3521), .A2(n3520), .A3(n3519), .A4(n3518), .ZN(n3522)
         );
  NAND4_X1 U4366 ( .A1(n3525), .A2(n3524), .A3(n3523), .A4(n3522), .ZN(n3584)
         );
  INV_X1 U4367 ( .A(keyinput37), .ZN(n3527) );
  AOI22_X1 U4368 ( .A1(n3528), .A2(DATAO_REG_10__SCAN_IN), .B1(
        DATAO_REG_8__SCAN_IN), .B2(n3527), .ZN(n3526) );
  OAI221_X1 U4369 ( .B1(n3528), .B2(DATAO_REG_10__SCAN_IN), .C1(n3527), .C2(
        DATAO_REG_8__SCAN_IN), .A(n3526), .ZN(n3541) );
  AOI22_X1 U4370 ( .A1(n3531), .A2(DATAO_REG_4__SCAN_IN), .B1(
        DATAO_REG_0__SCAN_IN), .B2(n3530), .ZN(n3529) );
  OAI221_X1 U4371 ( .B1(n3531), .B2(DATAO_REG_4__SCAN_IN), .C1(n3530), .C2(
        DATAO_REG_0__SCAN_IN), .A(n3529), .ZN(n3540) );
  INV_X1 U4372 ( .A(keyinput49), .ZN(n3534) );
  INV_X1 U4373 ( .A(keyinput102), .ZN(n3533) );
  AOI22_X1 U4374 ( .A1(n3534), .A2(DATAO_REG_11__SCAN_IN), .B1(
        DATAO_REG_13__SCAN_IN), .B2(n3533), .ZN(n3532) );
  OAI221_X1 U4375 ( .B1(n3534), .B2(DATAO_REG_11__SCAN_IN), .C1(n3533), .C2(
        DATAO_REG_13__SCAN_IN), .A(n3532), .ZN(n3539) );
  INV_X1 U4376 ( .A(keyinput113), .ZN(n3537) );
  INV_X1 U4377 ( .A(keyinput73), .ZN(n3536) );
  AOI22_X1 U4378 ( .A1(n3537), .A2(DATAO_REG_6__SCAN_IN), .B1(
        DATAO_REG_1__SCAN_IN), .B2(n3536), .ZN(n3535) );
  OAI221_X1 U4379 ( .B1(n3537), .B2(DATAO_REG_6__SCAN_IN), .C1(n3536), .C2(
        DATAO_REG_1__SCAN_IN), .A(n3535), .ZN(n3538) );
  NOR4_X1 U4380 ( .A1(n3541), .A2(n3540), .A3(n3539), .A4(n3538), .ZN(n3582)
         );
  INV_X1 U4381 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3544) );
  INV_X1 U4382 ( .A(keyinput48), .ZN(n3543) );
  AOI22_X1 U4383 ( .A1(n3544), .A2(keyinput8), .B1(ADDR_REG_3__SCAN_IN), .B2(
        n3543), .ZN(n3542) );
  OAI221_X1 U4384 ( .B1(n3544), .B2(keyinput8), .C1(n3543), .C2(
        ADDR_REG_3__SCAN_IN), .A(n3542), .ZN(n3555) );
  AOI22_X1 U4385 ( .A1(U3149), .A2(keyinput72), .B1(keyinput25), .B2(n3546), 
        .ZN(n3545) );
  OAI221_X1 U4386 ( .B1(U3149), .B2(keyinput72), .C1(n3546), .C2(keyinput25), 
        .A(n3545), .ZN(n3554) );
  INV_X1 U4387 ( .A(REG2_REG_17__SCAN_IN), .ZN(n3548) );
  NAND2_X1 U4388 ( .A1(n3548), .A2(keyinput35), .ZN(n3547) );
  OAI221_X1 U4389 ( .B1(n3549), .B2(keyinput114), .C1(n3548), .C2(keyinput35), 
        .A(n3547), .ZN(n3553) );
  INV_X1 U4390 ( .A(REG3_REG_0__SCAN_IN), .ZN(n4677) );
  XOR2_X1 U4391 ( .A(n4677), .B(keyinput77), .Z(n3551) );
  XNOR2_X1 U4392 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput112), .ZN(n3550) );
  NAND2_X1 U4393 ( .A1(n3551), .A2(n3550), .ZN(n3552) );
  NOR4_X1 U4394 ( .A1(n3555), .A2(n3554), .A3(n3553), .A4(n3552), .ZN(n3581)
         );
  INV_X1 U4395 ( .A(REG3_REG_9__SCAN_IN), .ZN(n3694) );
  AOI22_X1 U4396 ( .A1(n3557), .A2(keyinput51), .B1(n3694), .B2(keyinput98), 
        .ZN(n3556) );
  OAI221_X1 U4397 ( .B1(n3557), .B2(keyinput51), .C1(n3694), .C2(keyinput98), 
        .A(n3556), .ZN(n3568) );
  INV_X1 U4398 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4753) );
  AOI22_X1 U4399 ( .A1(n4753), .A2(keyinput30), .B1(keyinput39), .B2(n3559), 
        .ZN(n3558) );
  OAI221_X1 U4400 ( .B1(n4753), .B2(keyinput30), .C1(n3559), .C2(keyinput39), 
        .A(n3558), .ZN(n3567) );
  INV_X1 U4401 ( .A(REG2_REG_31__SCAN_IN), .ZN(n4661) );
  INV_X1 U4402 ( .A(REG2_REG_23__SCAN_IN), .ZN(n3561) );
  AOI22_X1 U4403 ( .A1(n4661), .A2(keyinput70), .B1(n3561), .B2(keyinput32), 
        .ZN(n3560) );
  OAI221_X1 U4404 ( .B1(n4661), .B2(keyinput70), .C1(n3561), .C2(keyinput32), 
        .A(n3560), .ZN(n3566) );
  INV_X1 U4405 ( .A(keyinput12), .ZN(n3562) );
  XOR2_X1 U4406 ( .A(ADDR_REG_1__SCAN_IN), .B(n3562), .Z(n3564) );
  XNOR2_X1 U4407 ( .A(REG1_REG_0__SCAN_IN), .B(keyinput17), .ZN(n3563) );
  NAND2_X1 U4408 ( .A1(n3564), .A2(n3563), .ZN(n3565) );
  NOR4_X1 U4409 ( .A1(n3568), .A2(n3567), .A3(n3566), .A4(n3565), .ZN(n3580)
         );
  INV_X1 U4410 ( .A(REG3_REG_26__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U4411 ( .A1(n2742), .A2(keyinput40), .B1(keyinput52), .B2(n4042), 
        .ZN(n3569) );
  OAI221_X1 U4412 ( .B1(n2742), .B2(keyinput40), .C1(n4042), .C2(keyinput52), 
        .A(n3569), .ZN(n3578) );
  INV_X1 U4413 ( .A(keyinput121), .ZN(n3572) );
  AOI22_X1 U4414 ( .A1(n3572), .A2(DATAO_REG_9__SCAN_IN), .B1(
        DATAO_REG_14__SCAN_IN), .B2(n3571), .ZN(n3570) );
  OAI221_X1 U4415 ( .B1(n3572), .B2(DATAO_REG_9__SCAN_IN), .C1(n3571), .C2(
        DATAO_REG_14__SCAN_IN), .A(n3570), .ZN(n3577) );
  INV_X1 U4416 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4023) );
  AOI22_X1 U4417 ( .A1(n4000), .A2(keyinput90), .B1(keyinput63), .B2(n4023), 
        .ZN(n3573) );
  OAI221_X1 U4418 ( .B1(n4000), .B2(keyinput90), .C1(n4023), .C2(keyinput63), 
        .A(n3573), .ZN(n3576) );
  AOI22_X1 U4419 ( .A1(n2992), .A2(keyinput3), .B1(keyinput60), .B2(n3941), 
        .ZN(n3574) );
  OAI221_X1 U4420 ( .B1(n2992), .B2(keyinput3), .C1(n3941), .C2(keyinput60), 
        .A(n3574), .ZN(n3575) );
  NOR4_X1 U4421 ( .A1(n3578), .A2(n3577), .A3(n3576), .A4(n3575), .ZN(n3579)
         );
  NAND4_X1 U4422 ( .A1(n3582), .A2(n3581), .A3(n3580), .A4(n3579), .ZN(n3583)
         );
  NOR4_X1 U4423 ( .A1(n3586), .A2(n3585), .A3(n3584), .A4(n3583), .ZN(n3587)
         );
  OAI21_X1 U4424 ( .B1(DATAO_REG_7__SCAN_IN), .B2(n3588), .A(n3587), .ZN(n3589) );
  XNOR2_X1 U4425 ( .A(n3590), .B(n3589), .ZN(U3210) );
  AND2_X1 U4426 ( .A1(n4080), .A2(n4089), .ZN(n4148) );
  XNOR2_X1 U4427 ( .A(n3591), .B(n4148), .ZN(n3622) );
  OAI22_X1 U4428 ( .A1(n3616), .A2(n4578), .B1(n3595), .B2(n4577), .ZN(n3594)
         );
  XOR2_X1 U4429 ( .A(n4148), .B(n3592), .Z(n3593) );
  INV_X1 U4430 ( .A(n3679), .ZN(n3643) );
  OAI22_X1 U4431 ( .A1(n3593), .A2(n4486), .B1(n3643), .B2(n4482), .ZN(n3613)
         );
  AOI211_X1 U4432 ( .C1(n3622), .C2(n4856), .A(n3594), .B(n3613), .ZN(n3603)
         );
  NOR2_X1 U4433 ( .A1(n3596), .A2(n3595), .ZN(n3597) );
  OR2_X1 U4434 ( .A1(n3663), .A2(n3597), .ZN(n3620) );
  OAI22_X1 U4435 ( .A1(n3620), .A2(n4585), .B1(n4867), .B2(n2450), .ZN(n3598)
         );
  INV_X1 U4436 ( .A(n3598), .ZN(n3599) );
  OAI21_X1 U4437 ( .B1(n3603), .B2(n4865), .A(n3599), .ZN(U3524) );
  INV_X1 U4438 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3600) );
  OAI22_X1 U4439 ( .A1(n3620), .A2(n4628), .B1(n4860), .B2(n3600), .ZN(n3601)
         );
  INV_X1 U4440 ( .A(n3601), .ZN(n3602) );
  OAI21_X1 U4441 ( .B1(n3603), .B2(n4858), .A(n3602), .ZN(U3479) );
  XNOR2_X1 U4442 ( .A(n3606), .B(n3605), .ZN(n3607) );
  XNOR2_X1 U4443 ( .A(n3604), .B(n3607), .ZN(n3612) );
  AOI22_X1 U4444 ( .A1(n4054), .A2(n3759), .B1(n4053), .B2(n3640), .ZN(n3611)
         );
  OAI21_X1 U4445 ( .B1(n4043), .B2(n3643), .A(n3608), .ZN(n3609) );
  AOI21_X1 U4446 ( .B1(n3678), .B2(n4041), .A(n3609), .ZN(n3610) );
  OAI211_X1 U4447 ( .C1(n3612), .C2(n4062), .A(n3611), .B(n3610), .ZN(U3218)
         );
  INV_X1 U4448 ( .A(n3613), .ZN(n3624) );
  INV_X1 U4449 ( .A(n4521), .ZN(n3783) );
  AOI22_X1 U4450 ( .A1(n4781), .A2(REG2_REG_6__SCAN_IN), .B1(n3614), .B2(n4785), .ZN(n3615) );
  OAI21_X1 U4451 ( .B1(n3616), .B2(n4444), .A(n3615), .ZN(n3617) );
  AOI21_X1 U4452 ( .B1(n3618), .B2(n4446), .A(n3617), .ZN(n3619) );
  OAI21_X1 U4453 ( .B1(n3620), .B2(n4493), .A(n3619), .ZN(n3621) );
  AOI21_X1 U4454 ( .B1(n3622), .B2(n3783), .A(n3621), .ZN(n3623) );
  OAI21_X1 U4455 ( .B1(n3624), .B2(n4781), .A(n3623), .ZN(U3284) );
  INV_X1 U4456 ( .A(n3625), .ZN(n3637) );
  NAND2_X1 U4457 ( .A1(n3626), .A2(n4776), .ZN(n3633) );
  INV_X1 U4458 ( .A(n3627), .ZN(n3628) );
  OAI22_X1 U4459 ( .A1(n4517), .A2(n3629), .B1(n3628), .B2(n4420), .ZN(n3630)
         );
  AOI21_X1 U4460 ( .B1(n3631), .B2(n4446), .A(n3630), .ZN(n3632) );
  OAI211_X1 U4461 ( .C1(n2421), .C2(n4444), .A(n3633), .B(n3632), .ZN(n3634)
         );
  AOI21_X1 U4462 ( .B1(n3635), .B2(n3783), .A(n3634), .ZN(n3636) );
  OAI21_X1 U4463 ( .B1(n3637), .B2(n4781), .A(n3636), .ZN(U3285) );
  AND2_X1 U4464 ( .A1(n4084), .A2(n4082), .ZN(n4156) );
  XOR2_X1 U4465 ( .A(n4156), .B(n3638), .Z(n3639) );
  AOI22_X1 U4466 ( .A1(n3639), .A2(n4514), .B1(n4508), .B2(n3759), .ZN(n3681)
         );
  INV_X1 U4467 ( .A(n2360), .ZN(n3653) );
  AOI21_X1 U4468 ( .B1(n3678), .B2(n3662), .A(n3653), .ZN(n3686) );
  AOI22_X1 U4469 ( .A1(n4781), .A2(REG2_REG_8__SCAN_IN), .B1(n3640), .B2(n4785), .ZN(n3642) );
  NAND2_X1 U4470 ( .A1(n4446), .A2(n3678), .ZN(n3641) );
  OAI211_X1 U4471 ( .C1(n3643), .C2(n4444), .A(n3642), .B(n3641), .ZN(n3646)
         );
  XOR2_X1 U4472 ( .A(n3644), .B(n4156), .Z(n3682) );
  NOR2_X1 U4473 ( .A1(n3682), .A2(n4521), .ZN(n3645) );
  AOI211_X1 U4474 ( .C1(n3686), .C2(n4776), .A(n3646), .B(n3645), .ZN(n3647)
         );
  OAI21_X1 U4475 ( .B1(n4781), .B2(n3681), .A(n3647), .ZN(U3282) );
  INV_X1 U4476 ( .A(n4099), .ZN(n3648) );
  AND2_X1 U4477 ( .A1(n3648), .A2(n4085), .ZN(n4159) );
  XNOR2_X1 U4478 ( .A(n3649), .B(n4159), .ZN(n3650) );
  INV_X1 U4479 ( .A(n3801), .ZN(n3707) );
  OAI22_X1 U4480 ( .A1(n3650), .A2(n4486), .B1(n3707), .B2(n4482), .ZN(n3741)
         );
  INV_X1 U4481 ( .A(n3741), .ZN(n3661) );
  XNOR2_X1 U4482 ( .A(n3651), .B(n4159), .ZN(n3743) );
  INV_X1 U4483 ( .A(n3727), .ZN(n3652) );
  OAI21_X1 U4484 ( .B1(n3653), .B2(n3739), .A(n3652), .ZN(n3749) );
  OAI22_X1 U4485 ( .A1(n3654), .A2(n4420), .B1(n4286), .B2(n4517), .ZN(n3656)
         );
  NOR2_X1 U4486 ( .A1(n4444), .A2(n3740), .ZN(n3655) );
  AOI211_X1 U4487 ( .C1(n4446), .C2(n3657), .A(n3656), .B(n3655), .ZN(n3658)
         );
  OAI21_X1 U4488 ( .B1(n3749), .B2(n4493), .A(n3658), .ZN(n3659) );
  AOI21_X1 U4489 ( .B1(n3743), .B2(n3783), .A(n3659), .ZN(n3660) );
  OAI21_X1 U4490 ( .B1(n3661), .B2(n4781), .A(n3660), .ZN(U3281) );
  OAI211_X1 U4491 ( .C1(n3663), .C2(n3668), .A(n4829), .B(n3662), .ZN(n4850)
         );
  XNOR2_X1 U4492 ( .A(n3664), .B(n4142), .ZN(n3670) );
  NAND2_X1 U4493 ( .A1(n3665), .A2(n4506), .ZN(n3667) );
  NAND2_X1 U4494 ( .A1(n3695), .A2(n4508), .ZN(n3666) );
  OAI211_X1 U4495 ( .C1(n4577), .C2(n3668), .A(n3667), .B(n3666), .ZN(n3669)
         );
  AOI21_X1 U4496 ( .B1(n3670), .B2(n4514), .A(n3669), .ZN(n4851) );
  OAI21_X1 U4497 ( .B1(n4516), .B2(n4850), .A(n4851), .ZN(n3676) );
  OAI22_X1 U4498 ( .A1(n4517), .A2(n3672), .B1(n3671), .B2(n4420), .ZN(n3675)
         );
  NAND2_X1 U4499 ( .A1(n3673), .A2(n4142), .ZN(n4847) );
  AND3_X1 U4500 ( .A1(n4848), .A2(n4847), .A3(n3783), .ZN(n3674) );
  AOI211_X1 U4501 ( .C1(n3676), .C2(n4517), .A(n3675), .B(n3674), .ZN(n3677)
         );
  INV_X1 U4502 ( .A(n3677), .ZN(U3283) );
  AOI22_X1 U4503 ( .A1(n3679), .A2(n4506), .B1(n4658), .B2(n3678), .ZN(n3680)
         );
  OAI211_X1 U4504 ( .C1(n3682), .C2(n4590), .A(n3681), .B(n3680), .ZN(n3685)
         );
  NAND2_X1 U4505 ( .A1(n3685), .A2(n4867), .ZN(n3684) );
  NAND2_X1 U4506 ( .A1(n3686), .A2(n4666), .ZN(n3683) );
  OAI211_X1 U4507 ( .C1(n4867), .C2(n4263), .A(n3684), .B(n3683), .ZN(U3526)
         );
  INV_X1 U4508 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3689) );
  NAND2_X1 U4509 ( .A1(n3685), .A2(n4860), .ZN(n3688) );
  NAND2_X1 U4510 ( .A1(n3686), .A2(n4837), .ZN(n3687) );
  OAI211_X1 U4511 ( .C1(n4860), .C2(n3689), .A(n3688), .B(n3687), .ZN(U3483)
         );
  OAI21_X1 U4512 ( .B1(n3692), .B2(n3691), .A(n3690), .ZN(n3699) );
  AOI22_X1 U4513 ( .A1(n4054), .A2(n3801), .B1(n4053), .B2(n3693), .ZN(n3697)
         );
  NOR2_X1 U4514 ( .A1(STATE_REG_SCAN_IN), .A2(n3694), .ZN(n4687) );
  AOI21_X1 U4515 ( .B1(n4059), .B2(n3695), .A(n4687), .ZN(n3696) );
  OAI211_X1 U4516 ( .C1(n4056), .C2(n3739), .A(n3697), .B(n3696), .ZN(n3698)
         );
  AOI21_X1 U4517 ( .B1(n3699), .B2(n3713), .A(n3698), .ZN(n3700) );
  INV_X1 U4518 ( .A(n3700), .ZN(U3228) );
  XNOR2_X1 U4519 ( .A(n3701), .B(n4143), .ZN(n3703) );
  AND2_X1 U4520 ( .A1(n4232), .A2(n4508), .ZN(n3702) );
  AOI21_X1 U4521 ( .B1(n3703), .B2(n4514), .A(n3702), .ZN(n3803) );
  NAND2_X1 U4522 ( .A1(n3704), .A2(n4143), .ZN(n3705) );
  NAND2_X1 U4523 ( .A1(n2356), .A2(n3705), .ZN(n3798) );
  OAI21_X1 U4524 ( .B1(n3729), .B2(n3799), .A(n3776), .ZN(n3810) );
  AOI22_X1 U4525 ( .A1(n4781), .A2(REG2_REG_11__SCAN_IN), .B1(n3754), .B2(
        n4785), .ZN(n3706) );
  OAI21_X1 U4526 ( .B1(n3707), .B2(n4444), .A(n3706), .ZN(n3708) );
  AOI21_X1 U4527 ( .B1(n3709), .B2(n4446), .A(n3708), .ZN(n3710) );
  OAI21_X1 U4528 ( .B1(n3810), .B2(n4493), .A(n3710), .ZN(n3711) );
  AOI21_X1 U4529 ( .B1(n3798), .B2(n3783), .A(n3711), .ZN(n3712) );
  OAI21_X1 U4530 ( .B1(n4781), .B2(n3803), .A(n3712), .ZN(U3279) );
  NAND2_X1 U4531 ( .A1(n3714), .A2(n3713), .ZN(n3722) );
  AOI21_X1 U4532 ( .B1(n3690), .B2(n3716), .A(n3715), .ZN(n3721) );
  AOI22_X1 U4533 ( .A1(n4054), .A2(n3724), .B1(n4053), .B2(n3730), .ZN(n3720)
         );
  NOR2_X1 U4534 ( .A1(STATE_REG_SCAN_IN), .A2(n3717), .ZN(n4696) );
  NOR2_X1 U4535 ( .A1(n4056), .A2(n3760), .ZN(n3718) );
  AOI211_X1 U4536 ( .C1(n4059), .C2(n3759), .A(n4696), .B(n3718), .ZN(n3719)
         );
  OAI211_X1 U4537 ( .C1(n3722), .C2(n3721), .A(n3720), .B(n3719), .ZN(U3214)
         );
  AND2_X1 U4538 ( .A1(n4097), .A2(n4101), .ZN(n4157) );
  XOR2_X1 U4539 ( .A(n4157), .B(n3723), .Z(n3725) );
  INV_X1 U4540 ( .A(n3724), .ZN(n3792) );
  OAI22_X1 U4541 ( .A1(n3725), .A2(n4486), .B1(n3792), .B2(n4482), .ZN(n3762)
         );
  INV_X1 U4542 ( .A(n3762), .ZN(n3738) );
  XOR2_X1 U4543 ( .A(n4157), .B(n3726), .Z(n3764) );
  NOR2_X1 U4544 ( .A1(n3727), .A2(n3760), .ZN(n3728) );
  OR2_X1 U4545 ( .A1(n3729), .A2(n3728), .ZN(n3769) );
  INV_X1 U4546 ( .A(n4444), .ZN(n4331) );
  INV_X1 U4547 ( .A(n3730), .ZN(n3731) );
  OAI22_X1 U4548 ( .A1(n4517), .A2(n3491), .B1(n3731), .B2(n4420), .ZN(n3732)
         );
  AOI21_X1 U4549 ( .B1(n4331), .B2(n3759), .A(n3732), .ZN(n3735) );
  NAND2_X1 U4550 ( .A1(n4446), .A2(n3733), .ZN(n3734) );
  OAI211_X1 U4551 ( .C1(n3769), .C2(n4493), .A(n3735), .B(n3734), .ZN(n3736)
         );
  AOI21_X1 U4552 ( .B1(n3764), .B2(n3783), .A(n3736), .ZN(n3737) );
  OAI21_X1 U4553 ( .B1(n3738), .B2(n4781), .A(n3737), .ZN(U3280) );
  OAI22_X1 U4554 ( .A1(n3740), .A2(n4578), .B1(n3739), .B2(n4577), .ZN(n3742)
         );
  AOI211_X1 U4555 ( .C1(n3743), .C2(n4856), .A(n3742), .B(n3741), .ZN(n3746)
         );
  MUX2_X1 U4556 ( .A(n3744), .B(n3746), .S(n4867), .Z(n3745) );
  OAI21_X1 U4557 ( .B1(n4585), .B2(n3749), .A(n3745), .ZN(U3527) );
  INV_X1 U4558 ( .A(REG0_REG_9__SCAN_IN), .ZN(n3747) );
  MUX2_X1 U4559 ( .A(n3747), .B(n3746), .S(n4860), .Z(n3748) );
  OAI21_X1 U4560 ( .B1(n3749), .B2(n4628), .A(n3748), .ZN(U3485) );
  NOR2_X1 U4561 ( .A1(n3752), .A2(n2307), .ZN(n3753) );
  XNOR2_X1 U4562 ( .A(n3750), .B(n3753), .ZN(n3758) );
  AOI22_X1 U4563 ( .A1(n4054), .A2(n4232), .B1(n4053), .B2(n3754), .ZN(n3757)
         );
  AND2_X1 U4564 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4707) );
  NOR2_X1 U4565 ( .A1(n4056), .A2(n3799), .ZN(n3755) );
  AOI211_X1 U4566 ( .C1(n4059), .C2(n3801), .A(n4707), .B(n3755), .ZN(n3756)
         );
  OAI211_X1 U4567 ( .C1(n3758), .C2(n4062), .A(n3757), .B(n3756), .ZN(U3233)
         );
  INV_X1 U4568 ( .A(n3759), .ZN(n3761) );
  OAI22_X1 U4569 ( .A1(n3761), .A2(n4578), .B1(n3760), .B2(n4577), .ZN(n3763)
         );
  AOI211_X1 U4570 ( .C1(n4856), .C2(n3764), .A(n3763), .B(n3762), .ZN(n3766)
         );
  MUX2_X1 U4571 ( .A(n2489), .B(n3766), .S(n4867), .Z(n3765) );
  OAI21_X1 U4572 ( .B1(n3769), .B2(n4585), .A(n3765), .ZN(U3528) );
  INV_X1 U4573 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3767) );
  MUX2_X1 U4574 ( .A(n3767), .B(n3766), .S(n4860), .Z(n3768) );
  OAI21_X1 U4575 ( .B1(n3769), .B2(n4628), .A(n3768), .ZN(U3487) );
  NAND2_X1 U4576 ( .A1(n3771), .A2(n3770), .ZN(n3815) );
  AND2_X1 U4577 ( .A1(n3812), .A2(n3813), .ZN(n4158) );
  XNOR2_X1 U4578 ( .A(n3815), .B(n4158), .ZN(n3772) );
  NAND2_X1 U4579 ( .A1(n3772), .A2(n4514), .ZN(n3774) );
  AOI22_X1 U4580 ( .A1(n3843), .A2(n4508), .B1(n4658), .B2(n3794), .ZN(n3773)
         );
  OAI211_X1 U4581 ( .C1(n3792), .C2(n4578), .A(n3774), .B(n3773), .ZN(n4854)
         );
  INV_X1 U4582 ( .A(n4854), .ZN(n3785) );
  XOR2_X1 U4583 ( .A(n4158), .B(n3775), .Z(n4857) );
  INV_X1 U4584 ( .A(n3776), .ZN(n3778) );
  NOR2_X1 U4585 ( .A1(n3778), .A2(n3777), .ZN(n4853) );
  NOR3_X1 U4586 ( .A1(n4853), .A2(n2227), .A3(n4493), .ZN(n3782) );
  INV_X1 U4587 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3780) );
  INV_X1 U4588 ( .A(n3791), .ZN(n3779) );
  OAI22_X1 U4589 ( .A1(n4517), .A2(n3780), .B1(n3779), .B2(n4420), .ZN(n3781)
         );
  AOI211_X1 U4590 ( .C1(n4857), .C2(n3783), .A(n3782), .B(n3781), .ZN(n3784)
         );
  OAI21_X1 U4591 ( .B1(n4781), .B2(n3785), .A(n3784), .ZN(U3278) );
  INV_X1 U4592 ( .A(n3787), .ZN(n3789) );
  XNOR2_X1 U4593 ( .A(n3789), .B(n3788), .ZN(n3790) );
  XNOR2_X1 U4594 ( .A(n3786), .B(n3790), .ZN(n3797) );
  AOI22_X1 U4595 ( .A1(n4054), .A2(n3843), .B1(n4053), .B2(n3791), .ZN(n3796)
         );
  NAND2_X1 U4596 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4713) );
  OAI21_X1 U4597 ( .B1(n4043), .B2(n3792), .A(n4713), .ZN(n3793) );
  AOI21_X1 U4598 ( .B1(n3794), .B2(n4041), .A(n3793), .ZN(n3795) );
  OAI211_X1 U4599 ( .C1(n3797), .C2(n4062), .A(n3796), .B(n3795), .ZN(U3221)
         );
  NAND2_X1 U4600 ( .A1(n3798), .A2(n4856), .ZN(n3804) );
  NOR2_X1 U4601 ( .A1(n3799), .A2(n4577), .ZN(n3800) );
  AOI21_X1 U4602 ( .B1(n3801), .B2(n4506), .A(n3800), .ZN(n3802) );
  NAND3_X1 U4603 ( .A1(n3804), .A2(n3803), .A3(n3802), .ZN(n3807) );
  MUX2_X1 U4604 ( .A(REG1_REG_11__SCAN_IN), .B(n3807), .S(n4867), .Z(n3805) );
  INV_X1 U4605 ( .A(n3805), .ZN(n3806) );
  OAI21_X1 U4606 ( .B1(n4585), .B2(n3810), .A(n3806), .ZN(U3529) );
  MUX2_X1 U4607 ( .A(REG0_REG_11__SCAN_IN), .B(n3807), .S(n4860), .Z(n3808) );
  INV_X1 U4608 ( .A(n3808), .ZN(n3809) );
  OAI21_X1 U4609 ( .B1(n3810), .B2(n4628), .A(n3809), .ZN(U3489) );
  XNOR2_X1 U4610 ( .A(n3843), .B(n3817), .ZN(n4149) );
  XNOR2_X1 U4611 ( .A(n3811), .B(n4149), .ZN(n3866) );
  INV_X1 U4612 ( .A(n3812), .ZN(n3814) );
  OAI21_X1 U4613 ( .B1(n3815), .B2(n3814), .A(n3813), .ZN(n3816) );
  XOR2_X1 U4614 ( .A(n4149), .B(n3816), .Z(n3821) );
  AOI22_X1 U4615 ( .A1(n4058), .A2(n4508), .B1(n4658), .B2(n3817), .ZN(n3818)
         );
  OAI21_X1 U4616 ( .B1(n3819), .B2(n4578), .A(n3818), .ZN(n3820) );
  AOI21_X1 U4617 ( .B1(n3821), .B2(n4514), .A(n3820), .ZN(n3822) );
  OAI21_X1 U4618 ( .B1(n3866), .B2(n3842), .A(n3822), .ZN(n3867) );
  NAND2_X1 U4619 ( .A1(n3867), .A2(n4517), .ZN(n3827) );
  OAI21_X1 U4620 ( .B1(n2227), .B2(n3833), .A(n3845), .ZN(n3873) );
  INV_X1 U4621 ( .A(n3873), .ZN(n3825) );
  OAI22_X1 U4622 ( .A1(n4517), .A2(n4721), .B1(n3823), .B2(n4420), .ZN(n3824)
         );
  AOI21_X1 U4623 ( .B1(n3825), .B2(n4776), .A(n3824), .ZN(n3826) );
  OAI211_X1 U4624 ( .C1(n3866), .C2(n4469), .A(n3827), .B(n3826), .ZN(U3277)
         );
  NOR2_X1 U4625 ( .A1(n3828), .A2(n2204), .ZN(n3829) );
  XNOR2_X1 U4626 ( .A(n3830), .B(n3829), .ZN(n3837) );
  AOI22_X1 U4627 ( .A1(n4054), .A2(n4058), .B1(n4053), .B2(n3831), .ZN(n3836)
         );
  NOR2_X1 U4628 ( .A1(STATE_REG_SCAN_IN), .A2(n3832), .ZN(n4726) );
  NOR2_X1 U4629 ( .A1(n4056), .A2(n3833), .ZN(n3834) );
  AOI211_X1 U4630 ( .C1(n4059), .C2(n4232), .A(n4726), .B(n3834), .ZN(n3835)
         );
  OAI211_X1 U4631 ( .C1(n3837), .C2(n4062), .A(n3836), .B(n3835), .ZN(U3231)
         );
  OAI21_X1 U4632 ( .B1(n3839), .B2(n4146), .A(n3838), .ZN(n3910) );
  INV_X1 U4633 ( .A(n3910), .ZN(n3852) );
  OAI21_X1 U4634 ( .B1(n2246), .B2(n4183), .A(n3854), .ZN(n3840) );
  AOI22_X1 U4635 ( .A1(n3840), .A2(n4514), .B1(n4508), .B2(n4231), .ZN(n3841)
         );
  OAI21_X1 U4636 ( .B1(n3852), .B2(n3842), .A(n3841), .ZN(n3908) );
  NAND2_X1 U4637 ( .A1(n3908), .A2(n4517), .ZN(n3851) );
  INV_X1 U4638 ( .A(n3843), .ZN(n3907) );
  AOI22_X1 U4639 ( .A1(n4781), .A2(REG2_REG_14__SCAN_IN), .B1(n3900), .B2(
        n4785), .ZN(n3844) );
  OAI21_X1 U4640 ( .B1(n3907), .B2(n4444), .A(n3844), .ZN(n3849) );
  INV_X1 U4641 ( .A(n3845), .ZN(n3847) );
  INV_X1 U4642 ( .A(n3859), .ZN(n3846) );
  OAI21_X1 U4643 ( .B1(n3847), .B2(n3906), .A(n3846), .ZN(n3916) );
  NOR2_X1 U4644 ( .A1(n3916), .A2(n4493), .ZN(n3848) );
  AOI211_X1 U4645 ( .C1(n4446), .C2(n3902), .A(n3849), .B(n3848), .ZN(n3850)
         );
  OAI211_X1 U4646 ( .C1(n3852), .C2(n4469), .A(n3851), .B(n3850), .ZN(U3276)
         );
  XNOR2_X1 U4647 ( .A(n3853), .B(n4147), .ZN(n3888) );
  INV_X1 U4648 ( .A(n3888), .ZN(n3865) );
  NAND2_X1 U4649 ( .A1(n3854), .A2(n4107), .ZN(n3855) );
  XNOR2_X1 U4650 ( .A(n3855), .B(n4147), .ZN(n3858) );
  INV_X1 U4651 ( .A(n4230), .ZN(n4579) );
  OAI22_X1 U4652 ( .A1(n4579), .A2(n4482), .B1(n4577), .B2(n4055), .ZN(n3856)
         );
  AOI21_X1 U4653 ( .B1(n4506), .B2(n4058), .A(n3856), .ZN(n3857) );
  OAI21_X1 U4654 ( .B1(n3858), .B2(n4486), .A(n3857), .ZN(n3887) );
  OAI21_X1 U4655 ( .B1(n3859), .B2(n4055), .A(n3882), .ZN(n3893) );
  NOR2_X1 U4656 ( .A1(n3893), .A2(n4493), .ZN(n3863) );
  INV_X1 U4657 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3861) );
  INV_X1 U4658 ( .A(n4052), .ZN(n3860) );
  OAI22_X1 U4659 ( .A1(n4517), .A2(n3861), .B1(n3860), .B2(n4420), .ZN(n3862)
         );
  AOI211_X1 U4660 ( .C1(n3887), .C2(n4517), .A(n3863), .B(n3862), .ZN(n3864)
         );
  OAI21_X1 U4661 ( .B1(n3865), .B2(n4521), .A(n3864), .ZN(U3275) );
  INV_X1 U4662 ( .A(n3866), .ZN(n3868) );
  AOI21_X1 U4663 ( .B1(n4844), .B2(n3868), .A(n3867), .ZN(n3870) );
  MUX2_X1 U4664 ( .A(n4271), .B(n3870), .S(n4867), .Z(n3869) );
  OAI21_X1 U4665 ( .B1(n4585), .B2(n3873), .A(n3869), .ZN(U3531) );
  INV_X1 U4666 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3871) );
  MUX2_X1 U4667 ( .A(n3871), .B(n3870), .S(n4860), .Z(n3872) );
  OAI21_X1 U4668 ( .B1(n3873), .B2(n4628), .A(n3872), .ZN(U3493) );
  OAI21_X1 U4669 ( .B1(n3874), .B2(n2558), .A(n3875), .ZN(n4591) );
  XNOR2_X1 U4670 ( .A(n3876), .B(n2558), .ZN(n3881) );
  NAND2_X1 U4671 ( .A1(n4231), .A2(n4506), .ZN(n3878) );
  NAND2_X1 U4672 ( .A1(n4507), .A2(n4508), .ZN(n3877) );
  OAI211_X1 U4673 ( .C1(n4577), .C2(n3879), .A(n3878), .B(n3877), .ZN(n3880)
         );
  AOI21_X1 U4674 ( .B1(n3881), .B2(n4514), .A(n3880), .ZN(n4589) );
  AOI22_X1 U4675 ( .A1(n4781), .A2(REG2_REG_16__SCAN_IN), .B1(n3979), .B2(
        n4785), .ZN(n3884) );
  NAND2_X1 U4676 ( .A1(n3882), .A2(n3982), .ZN(n4586) );
  NAND3_X1 U4677 ( .A1(n4587), .A2(n4776), .A3(n4586), .ZN(n3883) );
  OAI211_X1 U4678 ( .C1(n4589), .C2(n4781), .A(n3884), .B(n3883), .ZN(n3885)
         );
  INV_X1 U4679 ( .A(n3885), .ZN(n3886) );
  OAI21_X1 U4680 ( .B1(n4591), .B2(n4521), .A(n3886), .ZN(U3274) );
  AOI21_X1 U4681 ( .B1(n3888), .B2(n4856), .A(n3887), .ZN(n3891) );
  MUX2_X1 U4682 ( .A(n3891), .B(n3889), .S(n4865), .Z(n3890) );
  OAI21_X1 U4683 ( .B1(n4585), .B2(n3893), .A(n3890), .ZN(U3533) );
  MUX2_X1 U4684 ( .A(n3891), .B(n3512), .S(n4858), .Z(n3892) );
  OAI21_X1 U4685 ( .B1(n3893), .B2(n4628), .A(n3892), .ZN(U3497) );
  INV_X1 U4686 ( .A(n3894), .ZN(n3899) );
  AOI21_X1 U4687 ( .B1(n3898), .B2(n3896), .A(n3895), .ZN(n3897) );
  AOI21_X1 U4688 ( .B1(n3899), .B2(n3898), .A(n3897), .ZN(n3905) );
  AOI22_X1 U4689 ( .A1(n4054), .A2(n4231), .B1(n4053), .B2(n3900), .ZN(n3904)
         );
  INV_X1 U4690 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4732) );
  OAI22_X1 U4691 ( .A1(n4043), .A2(n3907), .B1(STATE_REG_SCAN_IN), .B2(n4732), 
        .ZN(n3901) );
  AOI21_X1 U4692 ( .B1(n3902), .B2(n4041), .A(n3901), .ZN(n3903) );
  OAI211_X1 U4693 ( .C1(n3905), .C2(n4062), .A(n3904), .B(n3903), .ZN(U3212)
         );
  OAI22_X1 U4694 ( .A1(n3907), .A2(n4578), .B1(n3906), .B2(n4577), .ZN(n3909)
         );
  AOI211_X1 U4695 ( .C1(n4844), .C2(n3910), .A(n3909), .B(n3908), .ZN(n3913)
         );
  MUX2_X1 U4696 ( .A(n3911), .B(n3913), .S(n4867), .Z(n3912) );
  OAI21_X1 U4697 ( .B1(n4585), .B2(n3916), .A(n3912), .ZN(U3532) );
  INV_X1 U4698 ( .A(REG0_REG_14__SCAN_IN), .ZN(n3914) );
  MUX2_X1 U4699 ( .A(n3914), .B(n3913), .S(n4860), .Z(n3915) );
  OAI21_X1 U4700 ( .B1(n3916), .B2(n4628), .A(n3915), .ZN(U3495) );
  AND2_X1 U4701 ( .A1(n4474), .A2(n4186), .ZN(n4136) );
  XNOR2_X1 U4702 ( .A(n3917), .B(n4136), .ZN(n4582) );
  INV_X1 U4703 ( .A(n4582), .ZN(n3930) );
  XNOR2_X1 U4704 ( .A(n3918), .B(n4136), .ZN(n3919) );
  NAND2_X1 U4705 ( .A1(n3919), .A2(n4514), .ZN(n3921) );
  NAND2_X1 U4706 ( .A1(n4484), .A2(n4508), .ZN(n3920) );
  NAND2_X1 U4707 ( .A1(n3921), .A2(n3920), .ZN(n4581) );
  INV_X1 U4708 ( .A(n4587), .ZN(n3923) );
  INV_X1 U4709 ( .A(n4503), .ZN(n3922) );
  OAI21_X1 U4710 ( .B1(n3923), .B2(n4576), .A(n3922), .ZN(n4629) );
  AOI22_X1 U4711 ( .A1(n4781), .A2(REG2_REG_17__SCAN_IN), .B1(n3991), .B2(
        n4785), .ZN(n3924) );
  OAI21_X1 U4712 ( .B1(n4579), .B2(n4444), .A(n3924), .ZN(n3925) );
  AOI21_X1 U4713 ( .B1(n3926), .B2(n4446), .A(n3925), .ZN(n3927) );
  OAI21_X1 U4714 ( .B1(n4629), .B2(n4493), .A(n3927), .ZN(n3928) );
  AOI21_X1 U4715 ( .B1(n4581), .B2(n4517), .A(n3928), .ZN(n3929) );
  OAI21_X1 U4716 ( .B1(n3930), .B2(n4521), .A(n3929), .ZN(U3273) );
  AOI22_X1 U4717 ( .A1(n4806), .A2(n3932), .B1(n3931), .B2(n2677), .ZN(U3458)
         );
  NAND3_X1 U4718 ( .A1(IR_REG_31__SCAN_IN), .A2(STATE_REG_SCAN_IN), .A3(n3934), 
        .ZN(n3936) );
  INV_X1 U4719 ( .A(DATAI_31_), .ZN(n3935) );
  OAI22_X1 U4720 ( .A1(n3933), .A2(n3936), .B1(STATE_REG_SCAN_IN), .B2(n3935), 
        .ZN(U3321) );
  AOI21_X1 U4721 ( .B1(n3937), .B2(n3938), .A(n4062), .ZN(n3940) );
  NAND2_X1 U4722 ( .A1(n3940), .A2(n3939), .ZN(n3945) );
  AOI22_X1 U4723 ( .A1(n4363), .A2(n4054), .B1(n4053), .B2(n4409), .ZN(n3944)
         );
  OAI22_X1 U4724 ( .A1(n4043), .A2(n4437), .B1(STATE_REG_SCAN_IN), .B2(n3941), 
        .ZN(n3942) );
  AOI21_X1 U4725 ( .B1(n4402), .B2(n4041), .A(n3942), .ZN(n3943) );
  NAND3_X1 U4726 ( .A1(n3945), .A2(n3944), .A3(n3943), .ZN(U3213) );
  INV_X1 U4727 ( .A(n3947), .ZN(n3948) );
  AOI21_X1 U4728 ( .B1(n3949), .B2(n3946), .A(n3948), .ZN(n3955) );
  AOI22_X1 U4729 ( .A1(n4054), .A2(n3961), .B1(n4053), .B2(n4491), .ZN(n3954)
         );
  NAND2_X1 U4730 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4647) );
  OAI21_X1 U4731 ( .B1(n4043), .B2(n3950), .A(n4647), .ZN(n3951) );
  AOI21_X1 U4732 ( .B1(n3952), .B2(n4041), .A(n3951), .ZN(n3953) );
  OAI211_X1 U4733 ( .C1(n3955), .C2(n4062), .A(n3954), .B(n3953), .ZN(U3216)
         );
  INV_X1 U4734 ( .A(n3956), .ZN(n3958) );
  NAND2_X1 U4735 ( .A1(n3958), .A2(n3957), .ZN(n3959) );
  XNOR2_X1 U4736 ( .A(n3960), .B(n3959), .ZN(n3966) );
  OAI22_X1 U4737 ( .A1(n4437), .A2(n4022), .B1(n4021), .B2(n4441), .ZN(n3964)
         );
  INV_X1 U4738 ( .A(n3961), .ZN(n4558) );
  INV_X1 U4739 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3962) );
  OAI22_X1 U4740 ( .A1(n4043), .A2(n4558), .B1(STATE_REG_SCAN_IN), .B2(n3962), 
        .ZN(n3963) );
  AOI211_X1 U4741 ( .C1(n4447), .C2(n4041), .A(n3964), .B(n3963), .ZN(n3965)
         );
  OAI21_X1 U4742 ( .B1(n3966), .B2(n4062), .A(n3965), .ZN(U3220) );
  XNOR2_X1 U4743 ( .A(n3969), .B(n3968), .ZN(n3970) );
  XNOR2_X1 U4744 ( .A(n3967), .B(n3970), .ZN(n3975) );
  INV_X1 U4745 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3971) );
  OAI22_X1 U4746 ( .A1(n4406), .A2(n4043), .B1(STATE_REG_SCAN_IN), .B2(n3971), 
        .ZN(n3973) );
  OAI22_X1 U4747 ( .A1(n4528), .A2(n4022), .B1(n4021), .B2(n4370), .ZN(n3972)
         );
  AOI211_X1 U4748 ( .C1(n4362), .C2(n4041), .A(n3973), .B(n3972), .ZN(n3974)
         );
  OAI21_X1 U4749 ( .B1(n3975), .B2(n4062), .A(n3974), .ZN(U3222) );
  INV_X1 U4750 ( .A(n4049), .ZN(n3976) );
  OAI21_X1 U4751 ( .B1(n3976), .B2(n4051), .A(n4048), .ZN(n3977) );
  XOR2_X1 U4752 ( .A(n3978), .B(n3977), .Z(n3985) );
  AOI22_X1 U4753 ( .A1(n4054), .A2(n4507), .B1(n4053), .B2(n3979), .ZN(n3984)
         );
  INV_X1 U4754 ( .A(n4231), .ZN(n3980) );
  NAND2_X1 U4755 ( .A1(REG3_REG_16__SCAN_IN), .A2(U3149), .ZN(n4752) );
  OAI21_X1 U4756 ( .B1(n4043), .B2(n3980), .A(n4752), .ZN(n3981) );
  AOI21_X1 U4757 ( .B1(n3982), .B2(n4041), .A(n3981), .ZN(n3983) );
  OAI211_X1 U4758 ( .C1(n3985), .C2(n4062), .A(n3984), .B(n3983), .ZN(U3223)
         );
  INV_X1 U4759 ( .A(n3987), .ZN(n3989) );
  NAND2_X1 U4760 ( .A1(n3989), .A2(n3988), .ZN(n3990) );
  XNOR2_X1 U4761 ( .A(n3986), .B(n3990), .ZN(n3995) );
  AOI22_X1 U4762 ( .A1(n4054), .A2(n4484), .B1(n4053), .B2(n3991), .ZN(n3994)
         );
  NOR2_X1 U4763 ( .A1(STATE_REG_SCAN_IN), .A2(n2560), .ZN(n4767) );
  NOR2_X1 U4764 ( .A1(n4056), .A2(n4576), .ZN(n3992) );
  AOI211_X1 U4765 ( .C1(n4059), .C2(n4230), .A(n4767), .B(n3992), .ZN(n3993)
         );
  OAI211_X1 U4766 ( .C1(n3995), .C2(n4062), .A(n3994), .B(n3993), .ZN(U3225)
         );
  NAND2_X1 U4767 ( .A1(n3996), .A2(n3997), .ZN(n3998) );
  XOR2_X1 U4768 ( .A(n3999), .B(n3998), .Z(n4004) );
  OAI22_X1 U4769 ( .A1(n4043), .A2(n4543), .B1(STATE_REG_SCAN_IN), .B2(n4000), 
        .ZN(n4002) );
  OAI22_X1 U4770 ( .A1(n4381), .A2(n4022), .B1(n4021), .B2(n4385), .ZN(n4001)
         );
  AOI211_X1 U4771 ( .C1(n4389), .C2(n4041), .A(n4002), .B(n4001), .ZN(n4003)
         );
  OAI21_X1 U4772 ( .B1(n4004), .B2(n4062), .A(n4003), .ZN(U3226) );
  INV_X1 U4773 ( .A(n4005), .ZN(n4010) );
  AOI21_X1 U4774 ( .B1(n4007), .B2(n4009), .A(n4006), .ZN(n4008) );
  AOI21_X1 U4775 ( .B1(n4010), .B2(n4009), .A(n4008), .ZN(n4016) );
  AOI22_X1 U4776 ( .A1(n4054), .A2(n4428), .B1(n4053), .B2(n4465), .ZN(n4015)
         );
  INV_X1 U4777 ( .A(n4509), .ZN(n4012) );
  OAI22_X1 U4778 ( .A1(n4043), .A2(n4012), .B1(STATE_REG_SCAN_IN), .B2(n4011), 
        .ZN(n4013) );
  AOI21_X1 U4779 ( .B1(n4466), .B2(n4041), .A(n4013), .ZN(n4014) );
  OAI211_X1 U4780 ( .C1(n4016), .C2(n4062), .A(n4015), .B(n4014), .ZN(U3230)
         );
  INV_X1 U4781 ( .A(n4017), .ZN(n4018) );
  AOI21_X1 U4782 ( .B1(n4020), .B2(n4019), .A(n4018), .ZN(n4027) );
  OAI22_X1 U4783 ( .A1(n4543), .A2(n4022), .B1(n4421), .B2(n4021), .ZN(n4025)
         );
  INV_X1 U4784 ( .A(n4428), .ZN(n4458) );
  OAI22_X1 U4785 ( .A1(n4043), .A2(n4458), .B1(STATE_REG_SCAN_IN), .B2(n4023), 
        .ZN(n4024) );
  AOI211_X1 U4786 ( .C1(n4427), .C2(n4041), .A(n4025), .B(n4024), .ZN(n4026)
         );
  OAI21_X1 U4787 ( .B1(n4027), .B2(n4062), .A(n4026), .ZN(U3232) );
  XOR2_X1 U4788 ( .A(n4029), .B(n4028), .Z(n4030) );
  XNOR2_X1 U4789 ( .A(n4031), .B(n4030), .ZN(n4037) );
  AOI22_X1 U4790 ( .A1(n4054), .A2(n4509), .B1(n4053), .B2(n4500), .ZN(n4036)
         );
  NAND2_X1 U4791 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4309) );
  OAI21_X1 U4792 ( .B1(n4043), .B2(n4032), .A(n4309), .ZN(n4033) );
  AOI21_X1 U4793 ( .B1(n4034), .B2(n4041), .A(n4033), .ZN(n4035) );
  OAI211_X1 U4794 ( .C1(n4037), .C2(n4062), .A(n4036), .B(n4035), .ZN(U3235)
         );
  NAND2_X1 U4795 ( .A1(n2196), .A2(n4039), .ZN(n4040) );
  XNOR2_X1 U4796 ( .A(n4038), .B(n4040), .ZN(n4047) );
  AOI22_X1 U4797 ( .A1(n4351), .A2(n4053), .B1(n4041), .B2(n4342), .ZN(n4046)
         );
  OAI22_X1 U4798 ( .A1(n4381), .A2(n4043), .B1(STATE_REG_SCAN_IN), .B2(n4042), 
        .ZN(n4044) );
  AOI21_X1 U4799 ( .B1(n4054), .B2(n4229), .A(n4044), .ZN(n4045) );
  OAI211_X1 U4800 ( .C1(n4047), .C2(n4062), .A(n4046), .B(n4045), .ZN(U3237)
         );
  NAND2_X1 U4801 ( .A1(n4049), .A2(n4048), .ZN(n4050) );
  XOR2_X1 U4802 ( .A(n4051), .B(n4050), .Z(n4063) );
  AOI22_X1 U4803 ( .A1(n4054), .A2(n4230), .B1(n4053), .B2(n4052), .ZN(n4061)
         );
  AND2_X1 U4804 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4746) );
  NOR2_X1 U4805 ( .A1(n4056), .A2(n4055), .ZN(n4057) );
  AOI211_X1 U4806 ( .C1(n4059), .C2(n4058), .A(n4746), .B(n4057), .ZN(n4060)
         );
  OAI211_X1 U4807 ( .C1(n4063), .C2(n4062), .A(n4061), .B(n4060), .ZN(U3238)
         );
  INV_X1 U4808 ( .A(n4125), .ZN(n4227) );
  AOI21_X1 U4809 ( .B1(n4227), .B2(n4065), .A(n4064), .ZN(n4180) );
  OAI211_X1 U4810 ( .C1(n4068), .C2(n4212), .A(n4067), .B(n4066), .ZN(n4070)
         );
  NAND3_X1 U4811 ( .A1(n4070), .A2(n4069), .A3(n2706), .ZN(n4073) );
  NAND3_X1 U4812 ( .A1(n4073), .A2(n4072), .A3(n4071), .ZN(n4076) );
  NAND3_X1 U4813 ( .A1(n4076), .A2(n4075), .A3(n4074), .ZN(n4078) );
  NAND4_X1 U4814 ( .A1(n4079), .A2(n4078), .A3(n4077), .A4(n4089), .ZN(n4081)
         );
  AND3_X1 U4815 ( .A1(n4081), .A2(n4142), .A3(n4080), .ZN(n4086) );
  NAND2_X1 U4816 ( .A1(n4083), .A2(n4082), .ZN(n4092) );
  OAI211_X1 U4817 ( .C1(n4086), .C2(n4092), .A(n4085), .B(n4084), .ZN(n4096)
         );
  NAND2_X1 U4818 ( .A1(n4088), .A2(n4087), .ZN(n4093) );
  INV_X1 U4819 ( .A(n4093), .ZN(n4095) );
  INV_X1 U4820 ( .A(n4089), .ZN(n4091) );
  NOR3_X1 U4821 ( .A1(n4092), .A2(n4091), .A3(n4090), .ZN(n4094) );
  NAND2_X1 U4822 ( .A1(n4093), .A2(n4106), .ZN(n4181) );
  AOI22_X1 U4823 ( .A1(n4096), .A2(n4095), .B1(n4094), .B2(n4181), .ZN(n4100)
         );
  INV_X1 U4824 ( .A(n4181), .ZN(n4098) );
  OAI22_X1 U4825 ( .A1(n4100), .A2(n4099), .B1(n4098), .B2(n4097), .ZN(n4104)
         );
  NAND4_X1 U4826 ( .A1(n4104), .A2(n4103), .A3(n4102), .A4(n4101), .ZN(n4111)
         );
  INV_X1 U4827 ( .A(n4105), .ZN(n4108) );
  NAND2_X1 U4828 ( .A1(n4107), .A2(n4106), .ZN(n4182) );
  OAI21_X1 U4829 ( .B1(n4108), .B2(n4182), .A(n4181), .ZN(n4110) );
  AOI21_X1 U4830 ( .B1(n4111), .B2(n4110), .A(n4109), .ZN(n4113) );
  INV_X1 U4831 ( .A(n4184), .ZN(n4112) );
  OAI211_X1 U4832 ( .C1(n4113), .C2(n4112), .A(n4188), .B(n4186), .ZN(n4114)
         );
  AOI211_X1 U4833 ( .C1(n4114), .C2(n4191), .A(n4190), .B(n4140), .ZN(n4117)
         );
  INV_X1 U4834 ( .A(n4115), .ZN(n4116) );
  OAI21_X1 U4835 ( .B1(n4117), .B2(n4194), .A(n4116), .ZN(n4119) );
  INV_X1 U4836 ( .A(n4163), .ZN(n4118) );
  NOR2_X1 U4837 ( .A1(n4161), .A2(n4118), .ZN(n4199) );
  OAI221_X1 U4838 ( .B1(n4196), .B2(n4198), .C1(n4196), .C2(n4119), .A(n4199), 
        .ZN(n4120) );
  NAND4_X1 U4839 ( .A1(n4180), .A2(n4178), .A3(n4121), .A4(n4120), .ZN(n4130)
         );
  NAND2_X1 U4840 ( .A1(n4123), .A2(n4122), .ZN(n4202) );
  NAND2_X1 U4841 ( .A1(n4125), .A2(n4124), .ZN(n4127) );
  NAND2_X1 U4842 ( .A1(n4524), .A2(n4656), .ZN(n4129) );
  OR2_X1 U4843 ( .A1(n4226), .A2(n4177), .ZN(n4126) );
  AND2_X1 U4844 ( .A1(n4129), .A2(n4126), .ZN(n4164) );
  NAND2_X1 U4845 ( .A1(n4127), .A2(n4164), .ZN(n4201) );
  AOI21_X1 U4846 ( .B1(n4202), .B2(n4180), .A(n4201), .ZN(n4206) );
  NAND2_X1 U4847 ( .A1(n4226), .A2(n4177), .ZN(n4209) );
  OR2_X1 U4848 ( .A1(n4524), .A2(n4656), .ZN(n4128) );
  NAND2_X1 U4849 ( .A1(n4209), .A2(n4128), .ZN(n4167) );
  AOI22_X1 U4850 ( .A1(n4130), .A2(n4206), .B1(n4129), .B2(n4167), .ZN(n4216)
         );
  INV_X1 U4851 ( .A(n4131), .ZN(n4176) );
  INV_X1 U4852 ( .A(n4323), .ZN(n4179) );
  AND2_X1 U4853 ( .A1(n4133), .A2(n4132), .ZN(n4455) );
  XNOR2_X1 U4854 ( .A(n4509), .B(n4488), .ZN(n4480) );
  INV_X1 U4855 ( .A(n4134), .ZN(n4357) );
  NOR2_X1 U4856 ( .A1(n4135), .A2(n4357), .ZN(n4380) );
  XNOR2_X1 U4857 ( .A(n4543), .B(n4402), .ZN(n4400) );
  INV_X1 U4858 ( .A(n4400), .ZN(n4137) );
  NAND4_X1 U4859 ( .A1(n4138), .A2(n4380), .A3(n4137), .A4(n4136), .ZN(n4139)
         );
  NOR3_X1 U4860 ( .A1(n4455), .A2(n4480), .A3(n4139), .ZN(n4175) );
  INV_X1 U4861 ( .A(n4140), .ZN(n4397) );
  NAND2_X1 U4862 ( .A1(n4397), .A2(n4395), .ZN(n4435) );
  NOR2_X1 U4863 ( .A1(n4435), .A2(n4141), .ZN(n4155) );
  AND4_X1 U4864 ( .A1(n4144), .A2(n4143), .A3(n4142), .A4(n3268), .ZN(n4154)
         );
  NOR2_X1 U4865 ( .A1(n4145), .A2(n2705), .ZN(n4153) );
  NOR2_X1 U4866 ( .A1(n4147), .A2(n4146), .ZN(n4151) );
  AND4_X1 U4867 ( .A1(n4151), .A2(n4150), .A3(n4149), .A4(n4148), .ZN(n4152)
         );
  NAND4_X1 U4868 ( .A1(n4155), .A2(n4154), .A3(n4153), .A4(n4152), .ZN(n4173)
         );
  INV_X1 U4869 ( .A(n4425), .ZN(n4171) );
  AND4_X1 U4870 ( .A1(n4159), .A2(n4158), .A3(n4157), .A4(n4156), .ZN(n4170)
         );
  INV_X1 U4871 ( .A(n4178), .ZN(n4160) );
  NOR2_X1 U4872 ( .A1(n4161), .A2(n4160), .ZN(n4339) );
  AND2_X1 U4873 ( .A1(n4163), .A2(n4162), .ZN(n4359) );
  NAND4_X1 U4874 ( .A1(n4165), .A2(n4339), .A3(n4359), .A4(n4164), .ZN(n4166)
         );
  NOR2_X1 U4875 ( .A1(n4167), .A2(n4166), .ZN(n4168) );
  NAND4_X1 U4876 ( .A1(n4171), .A2(n4170), .A3(n4169), .A4(n4168), .ZN(n4172)
         );
  NOR2_X1 U4877 ( .A1(n4173), .A2(n4172), .ZN(n4174) );
  AND4_X1 U4878 ( .A1(n4176), .A2(n4179), .A3(n4175), .A4(n4174), .ZN(n4214)
         );
  INV_X1 U4879 ( .A(n4524), .ZN(n4208) );
  NAND3_X1 U4880 ( .A1(n4180), .A2(n4179), .A3(n4178), .ZN(n4205) );
  OAI21_X1 U4881 ( .B1(n4183), .B2(n4182), .A(n4181), .ZN(n4185) );
  NAND2_X1 U4882 ( .A1(n4185), .A2(n4184), .ZN(n4189) );
  NAND4_X1 U4883 ( .A1(n4189), .A2(n4188), .A3(n4187), .A4(n4186), .ZN(n4192)
         );
  AOI21_X1 U4884 ( .B1(n4192), .B2(n4191), .A(n4190), .ZN(n4195) );
  OAI21_X1 U4885 ( .B1(n4195), .B2(n4194), .A(n4193), .ZN(n4197) );
  AOI21_X1 U4886 ( .B1(n4198), .B2(n4197), .A(n4196), .ZN(n4203) );
  INV_X1 U4887 ( .A(n4199), .ZN(n4200) );
  NOR4_X1 U4888 ( .A1(n4203), .A2(n4202), .A3(n4201), .A4(n4200), .ZN(n4204)
         );
  AOI21_X1 U4889 ( .B1(n4206), .B2(n4205), .A(n4204), .ZN(n4207) );
  AOI21_X1 U4890 ( .B1(n4525), .B2(n4208), .A(n4207), .ZN(n4211) );
  AOI21_X1 U4891 ( .B1(n4209), .B2(n4524), .A(n4656), .ZN(n4210) );
  NOR2_X1 U4892 ( .A1(n4211), .A2(n4210), .ZN(n4213) );
  MUX2_X1 U4893 ( .A(n4214), .B(n4213), .S(n4212), .Z(n4215) );
  MUX2_X1 U4894 ( .A(n4216), .B(n4215), .S(n4632), .Z(n4217) );
  XNOR2_X1 U4895 ( .A(n4217), .B(n4516), .ZN(n4225) );
  NAND4_X1 U4896 ( .A1(n4218), .A2(n4672), .A3(n4807), .A4(n4648), .ZN(n4219)
         );
  NOR2_X1 U4897 ( .A1(n4219), .A2(n2783), .ZN(n4220) );
  MUX2_X1 U4898 ( .A(n4221), .B(n4220), .S(n4631), .Z(n4223) );
  INV_X1 U4899 ( .A(B_REG_SCAN_IN), .ZN(n4222) );
  OAI22_X1 U4900 ( .A1(n4225), .A2(n4224), .B1(n4223), .B2(n4222), .ZN(U3239)
         );
  MUX2_X1 U4901 ( .A(n4226), .B(DATAO_REG_30__SCAN_IN), .S(n4235), .Z(U3580)
         );
  MUX2_X1 U4902 ( .A(DATAO_REG_29__SCAN_IN), .B(n4227), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4903 ( .A(DATAO_REG_28__SCAN_IN), .B(n4228), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4904 ( .A(DATAO_REG_27__SCAN_IN), .B(n4229), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4905 ( .A(n4332), .B(DATAO_REG_26__SCAN_IN), .S(n4235), .Z(U3576)
         );
  MUX2_X1 U4906 ( .A(n4343), .B(DATAO_REG_25__SCAN_IN), .S(n4235), .Z(U3575)
         );
  MUX2_X1 U4907 ( .A(n4363), .B(DATAO_REG_24__SCAN_IN), .S(n4235), .Z(U3574)
         );
  MUX2_X1 U4908 ( .A(n4428), .B(DATAO_REG_21__SCAN_IN), .S(n4235), .Z(U3571)
         );
  MUX2_X1 U4909 ( .A(n4484), .B(DATAO_REG_18__SCAN_IN), .S(n4235), .Z(U3568)
         );
  MUX2_X1 U4910 ( .A(n4230), .B(DATAO_REG_16__SCAN_IN), .S(n4235), .Z(U3566)
         );
  MUX2_X1 U4911 ( .A(n4231), .B(DATAO_REG_15__SCAN_IN), .S(n4235), .Z(U3565)
         );
  MUX2_X1 U4912 ( .A(n4232), .B(DATAO_REG_12__SCAN_IN), .S(n4235), .Z(U3562)
         );
  MUX2_X1 U4913 ( .A(n4233), .B(DATAO_REG_5__SCAN_IN), .S(n4235), .Z(U3555) );
  MUX2_X1 U4914 ( .A(n4234), .B(DATAO_REG_3__SCAN_IN), .S(n4235), .Z(U3553) );
  MUX2_X1 U4915 ( .A(n4236), .B(DATAO_REG_2__SCAN_IN), .S(n4235), .Z(U3552) );
  NAND2_X1 U4916 ( .A1(n4256), .A2(n4636), .ZN(n4246) );
  OAI211_X1 U4917 ( .C1(n4239), .C2(n4238), .A(n4769), .B(n4237), .ZN(n4245)
         );
  OAI211_X1 U4918 ( .C1(n4242), .C2(n4241), .A(n4711), .B(n4240), .ZN(n4244)
         );
  AOI22_X1 U4919 ( .A1(n4768), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4243) );
  NAND4_X1 U4920 ( .A1(n4246), .A2(n4245), .A3(n4244), .A4(n4243), .ZN(U3241)
         );
  AOI22_X1 U4921 ( .A1(n4768), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n4259) );
  OAI211_X1 U4922 ( .C1(n4249), .C2(n4248), .A(n4711), .B(n4247), .ZN(n4254)
         );
  OAI211_X1 U4923 ( .C1(n4252), .C2(n4251), .A(n4769), .B(n4250), .ZN(n4253)
         );
  AND2_X1 U4924 ( .A1(n4254), .A2(n4253), .ZN(n4258) );
  NAND2_X1 U4925 ( .A1(n4256), .A2(n2412), .ZN(n4257) );
  NAND4_X1 U4926 ( .A1(n4260), .A2(n4259), .A3(n4258), .A4(n4257), .ZN(U3242)
         );
  XNOR2_X1 U4927 ( .A(n4312), .B(REG1_REG_18__SCAN_IN), .ZN(n4642) );
  NOR2_X1 U4928 ( .A1(n4306), .A2(REG1_REG_17__SCAN_IN), .ZN(n4279) );
  NAND2_X1 U4929 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4303), .ZN(n4275) );
  INV_X1 U4930 ( .A(n4303), .ZN(n4814) );
  AOI22_X1 U4931 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4303), .B1(n4814), .B2(
        n3889), .ZN(n4749) );
  AOI22_X1 U4932 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4299), .B1(n4818), .B2(
        n4271), .ZN(n4729) );
  NAND2_X1 U4933 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4285), .ZN(n4268) );
  AOI22_X1 U4934 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4285), .B1(n4820), .B2(
        n2503), .ZN(n4700) );
  NAND2_X1 U4935 ( .A1(n4287), .A2(REG1_REG_9__SCAN_IN), .ZN(n4265) );
  INV_X1 U4936 ( .A(n4287), .ZN(n4824) );
  AOI22_X1 U4937 ( .A1(n4287), .A2(REG1_REG_9__SCAN_IN), .B1(n3744), .B2(n4824), .ZN(n4680) );
  INV_X1 U4938 ( .A(n4261), .ZN(n4262) );
  INV_X1 U4939 ( .A(n4633), .ZN(n4290) );
  NAND2_X1 U4940 ( .A1(n4293), .A2(n4266), .ZN(n4267) );
  NAND2_X1 U4941 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4690), .ZN(n4689) );
  NAND2_X1 U4942 ( .A1(n4709), .A2(n4269), .ZN(n4270) );
  NAND2_X1 U4943 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4717), .ZN(n4716) );
  NAND2_X1 U4944 ( .A1(n4272), .A2(n4273), .ZN(n4274) );
  NAND2_X1 U4945 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4739), .ZN(n4738) );
  NAND2_X1 U4946 ( .A1(n4274), .A2(n4738), .ZN(n4748) );
  NAND2_X1 U4947 ( .A1(n4749), .A2(n4748), .ZN(n4747) );
  NOR2_X1 U4948 ( .A1(n4276), .A2(n4277), .ZN(n4278) );
  INV_X1 U4949 ( .A(n4306), .ZN(n4810) );
  AOI22_X1 U4950 ( .A1(n4306), .A2(n4583), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4810), .ZN(n4770) );
  NOR2_X1 U4951 ( .A1(n4771), .A2(n4770), .ZN(n4772) );
  NOR2_X1 U4952 ( .A1(n4279), .A2(n4772), .ZN(n4643) );
  XOR2_X1 U4953 ( .A(n4642), .B(n4643), .Z(n4280) );
  NAND2_X1 U4954 ( .A1(n4280), .A2(n4769), .ZN(n4311) );
  INV_X1 U4955 ( .A(n4312), .ZN(n4641) );
  INV_X1 U4956 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4282) );
  NOR2_X1 U4957 ( .A1(n4641), .A2(n4282), .ZN(n4281) );
  AOI21_X1 U4958 ( .B1(n4641), .B2(n4282), .A(n4281), .ZN(n4308) );
  NOR2_X1 U4959 ( .A1(n4306), .A2(REG2_REG_17__SCAN_IN), .ZN(n4283) );
  AOI21_X1 U4960 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4306), .A(n4283), .ZN(n4765) );
  NOR2_X1 U4961 ( .A1(n4721), .A2(n4818), .ZN(n4720) );
  NAND2_X1 U4962 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4285), .ZN(n4296) );
  AOI22_X1 U4963 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4285), .B1(n4820), .B2(
        n4284), .ZN(n4703) );
  NAND2_X1 U4964 ( .A1(n4287), .A2(REG2_REG_9__SCAN_IN), .ZN(n4292) );
  AOI22_X1 U4965 ( .A1(n4287), .A2(REG2_REG_9__SCAN_IN), .B1(n4286), .B2(n4824), .ZN(n4683) );
  NAND2_X1 U4966 ( .A1(n4288), .A2(REG2_REG_8__SCAN_IN), .ZN(n4289) );
  OAI21_X1 U4967 ( .B1(n4291), .B2(n4290), .A(n4289), .ZN(n4682) );
  NAND2_X1 U4968 ( .A1(n4683), .A2(n4682), .ZN(n4681) );
  NAND2_X1 U4969 ( .A1(n4293), .A2(n4294), .ZN(n4295) );
  NAND2_X1 U4970 ( .A1(n4703), .A2(n4702), .ZN(n4701) );
  NAND2_X1 U4971 ( .A1(n4709), .A2(n4297), .ZN(n4298) );
  OAI22_X1 U4972 ( .A1(n4720), .A2(n4723), .B1(REG2_REG_13__SCAN_IN), .B2(
        n4299), .ZN(n4300) );
  NOR2_X1 U4973 ( .A1(n4816), .A2(n4300), .ZN(n4301) );
  INV_X1 U4974 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4735) );
  XNOR2_X1 U4975 ( .A(n4816), .B(n4300), .ZN(n4734) );
  NOR2_X1 U4976 ( .A1(n4735), .A2(n4734), .ZN(n4733) );
  NAND2_X1 U4977 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4303), .ZN(n4302) );
  OAI21_X1 U4978 ( .B1(REG2_REG_15__SCAN_IN), .B2(n4303), .A(n4302), .ZN(n4743) );
  NAND2_X1 U4979 ( .A1(n4304), .A2(n4812), .ZN(n4305) );
  NAND2_X1 U4980 ( .A1(n4765), .A2(n4763), .ZN(n4764) );
  OAI21_X1 U4981 ( .B1(n4306), .B2(REG2_REG_17__SCAN_IN), .A(n4764), .ZN(n4307) );
  NOR2_X1 U4982 ( .A1(n4307), .A2(n4308), .ZN(n4637) );
  OAI211_X1 U4983 ( .C1(n4775), .C2(n4312), .A(n4311), .B(n4310), .ZN(U3258)
         );
  INV_X1 U4984 ( .A(n4313), .ZN(n4318) );
  AOI22_X1 U4985 ( .A1(n4314), .A2(n4785), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4781), .ZN(n4315) );
  OAI21_X1 U4986 ( .B1(n4316), .B2(n4493), .A(n4315), .ZN(n4317) );
  AOI21_X1 U4987 ( .B1(n4318), .B2(n4517), .A(n4317), .ZN(n4319) );
  OAI21_X1 U4988 ( .B1(n4320), .B2(n4521), .A(n4319), .ZN(U3262) );
  XNOR2_X1 U4989 ( .A(n4321), .B(n4323), .ZN(n4531) );
  INV_X1 U4990 ( .A(n4531), .ZN(n4337) );
  AOI21_X1 U4991 ( .B1(n4324), .B2(n4323), .A(n4322), .ZN(n4326) );
  OAI22_X1 U4992 ( .A1(n4326), .A2(n4486), .B1(n4325), .B2(n4482), .ZN(n4530)
         );
  INV_X1 U4993 ( .A(n4327), .ZN(n4328) );
  OAI21_X1 U4994 ( .B1(n4347), .B2(n4527), .A(n4328), .ZN(n4598) );
  AOI22_X1 U4995 ( .A1(n4329), .A2(n4785), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4781), .ZN(n4334) );
  AOI22_X1 U4996 ( .A1(n4332), .A2(n4331), .B1(n4330), .B2(n4446), .ZN(n4333)
         );
  OAI211_X1 U4997 ( .C1(n4598), .C2(n4493), .A(n4334), .B(n4333), .ZN(n4335)
         );
  AOI21_X1 U4998 ( .B1(n4530), .B2(n4517), .A(n4335), .ZN(n4336) );
  OAI21_X1 U4999 ( .B1(n4337), .B2(n4521), .A(n4336), .ZN(U3263) );
  XNOR2_X1 U5000 ( .A(n4338), .B(n4339), .ZN(n4535) );
  INV_X1 U5001 ( .A(n4535), .ZN(n4355) );
  XNOR2_X1 U5002 ( .A(n4340), .B(n4339), .ZN(n4341) );
  NAND2_X1 U5003 ( .A1(n4341), .A2(n4514), .ZN(n4345) );
  AOI22_X1 U5004 ( .A1(n4343), .A2(n4506), .B1(n4342), .B2(n4658), .ZN(n4344)
         );
  OAI211_X1 U5005 ( .C1(n4346), .C2(n4482), .A(n4345), .B(n4344), .ZN(n4534)
         );
  INV_X1 U5006 ( .A(n4366), .ZN(n4350) );
  INV_X1 U5007 ( .A(n4347), .ZN(n4348) );
  OAI21_X1 U5008 ( .B1(n4350), .B2(n4349), .A(n4348), .ZN(n4602) );
  AOI22_X1 U5009 ( .A1(n4351), .A2(n4785), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4781), .ZN(n4352) );
  OAI21_X1 U5010 ( .B1(n4602), .B2(n4493), .A(n4352), .ZN(n4353) );
  AOI21_X1 U5011 ( .B1(n4534), .B2(n4517), .A(n4353), .ZN(n4354) );
  OAI21_X1 U5012 ( .B1(n4355), .B2(n4521), .A(n4354), .ZN(U3264) );
  XNOR2_X1 U5013 ( .A(n4356), .B(n4359), .ZN(n4539) );
  INV_X1 U5014 ( .A(n4539), .ZN(n4374) );
  NOR2_X1 U5015 ( .A1(n4358), .A2(n4357), .ZN(n4360) );
  XNOR2_X1 U5016 ( .A(n4360), .B(n4359), .ZN(n4361) );
  NAND2_X1 U5017 ( .A1(n4361), .A2(n4514), .ZN(n4365) );
  AOI22_X1 U5018 ( .A1(n4363), .A2(n4506), .B1(n4362), .B2(n4658), .ZN(n4364)
         );
  OAI211_X1 U5019 ( .C1(n4528), .C2(n4482), .A(n4365), .B(n4364), .ZN(n4538)
         );
  INV_X1 U5020 ( .A(n4383), .ZN(n4368) );
  OAI21_X1 U5021 ( .B1(n4368), .B2(n4367), .A(n4366), .ZN(n4605) );
  NOR2_X1 U5022 ( .A1(n4605), .A2(n4493), .ZN(n4372) );
  INV_X1 U5023 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4369) );
  OAI22_X1 U5024 ( .A1(n4370), .A2(n4420), .B1(n4369), .B2(n4517), .ZN(n4371)
         );
  AOI211_X1 U5025 ( .C1(n4538), .C2(n4517), .A(n4372), .B(n4371), .ZN(n4373)
         );
  OAI21_X1 U5026 ( .B1(n4374), .B2(n4521), .A(n4373), .ZN(U3265) );
  XNOR2_X1 U5027 ( .A(n4375), .B(n4380), .ZN(n4546) );
  INV_X1 U5028 ( .A(n4546), .ZN(n4393) );
  INV_X1 U5029 ( .A(n4376), .ZN(n4377) );
  NAND2_X1 U5030 ( .A1(n4378), .A2(n4377), .ZN(n4379) );
  XOR2_X1 U5031 ( .A(n4380), .B(n4379), .Z(n4382) );
  OAI22_X1 U5032 ( .A1(n4382), .A2(n4486), .B1(n4381), .B2(n4482), .ZN(n4545)
         );
  INV_X1 U5033 ( .A(n4407), .ZN(n4384) );
  OAI21_X1 U5034 ( .B1(n4384), .B2(n4542), .A(n4383), .ZN(n4609) );
  INV_X1 U5035 ( .A(n4385), .ZN(n4386) );
  AOI22_X1 U5036 ( .A1(n4386), .A2(n4785), .B1(REG2_REG_24__SCAN_IN), .B2(
        n4781), .ZN(n4387) );
  OAI21_X1 U5037 ( .B1(n4543), .B2(n4444), .A(n4387), .ZN(n4388) );
  AOI21_X1 U5038 ( .B1(n4389), .B2(n4446), .A(n4388), .ZN(n4390) );
  OAI21_X1 U5039 ( .B1(n4609), .B2(n4493), .A(n4390), .ZN(n4391) );
  AOI21_X1 U5040 ( .B1(n4545), .B2(n4517), .A(n4391), .ZN(n4392) );
  OAI21_X1 U5041 ( .B1(n4393), .B2(n4521), .A(n4392), .ZN(U3266) );
  XNOR2_X1 U5042 ( .A(n4394), .B(n4400), .ZN(n4550) );
  INV_X1 U5043 ( .A(n4550), .ZN(n4413) );
  INV_X1 U5044 ( .A(n4395), .ZN(n4396) );
  AOI21_X1 U5045 ( .B1(n4436), .B2(n4397), .A(n4396), .ZN(n4426) );
  OAI21_X1 U5046 ( .B1(n4426), .B2(n4425), .A(n4398), .ZN(n4399) );
  XOR2_X1 U5047 ( .A(n4400), .B(n4399), .Z(n4401) );
  NAND2_X1 U5048 ( .A1(n4401), .A2(n4514), .ZN(n4405) );
  AOI22_X1 U5049 ( .A1(n4403), .A2(n4506), .B1(n4658), .B2(n4402), .ZN(n4404)
         );
  OAI211_X1 U5050 ( .C1(n4406), .C2(n4482), .A(n4405), .B(n4404), .ZN(n4549)
         );
  OAI21_X1 U5051 ( .B1(n4419), .B2(n4408), .A(n4407), .ZN(n4612) );
  AOI22_X1 U5052 ( .A1(n4781), .A2(REG2_REG_23__SCAN_IN), .B1(n4409), .B2(
        n4785), .ZN(n4410) );
  OAI21_X1 U5053 ( .B1(n4612), .B2(n4493), .A(n4410), .ZN(n4411) );
  AOI21_X1 U5054 ( .B1(n4549), .B2(n4517), .A(n4411), .ZN(n4412) );
  OAI21_X1 U5055 ( .B1(n4413), .B2(n4521), .A(n4412), .ZN(U3267) );
  NOR2_X1 U5056 ( .A1(n4414), .A2(n4425), .ZN(n4415) );
  OR2_X1 U5057 ( .A1(n4416), .A2(n4415), .ZN(n4552) );
  NOR2_X1 U5058 ( .A1(n4439), .A2(n4417), .ZN(n4418) );
  OR2_X1 U5059 ( .A1(n4419), .A2(n4418), .ZN(n4616) );
  INV_X1 U5060 ( .A(n4616), .ZN(n4424) );
  INV_X1 U5061 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4422) );
  OAI22_X1 U5062 ( .A1(n4517), .A2(n4422), .B1(n4421), .B2(n4420), .ZN(n4423)
         );
  AOI21_X1 U5063 ( .B1(n4424), .B2(n4776), .A(n4423), .ZN(n4433) );
  XNOR2_X1 U5064 ( .A(n4426), .B(n4425), .ZN(n4431) );
  AOI22_X1 U5065 ( .A1(n4428), .A2(n4506), .B1(n4427), .B2(n4658), .ZN(n4429)
         );
  OAI21_X1 U5066 ( .B1(n4543), .B2(n4482), .A(n4429), .ZN(n4430) );
  AOI21_X1 U5067 ( .B1(n4431), .B2(n4514), .A(n4430), .ZN(n4553) );
  OR2_X1 U5068 ( .A1(n4553), .A2(n4781), .ZN(n4432) );
  OAI211_X1 U5069 ( .C1(n4552), .C2(n4521), .A(n4433), .B(n4432), .ZN(U3268)
         );
  XNOR2_X1 U5070 ( .A(n4434), .B(n4435), .ZN(n4561) );
  INV_X1 U5071 ( .A(n4561), .ZN(n4451) );
  XNOR2_X1 U5072 ( .A(n4436), .B(n4435), .ZN(n4438) );
  OAI22_X1 U5073 ( .A1(n4438), .A2(n4486), .B1(n4437), .B2(n4482), .ZN(n4560)
         );
  INV_X1 U5074 ( .A(n4439), .ZN(n4440) );
  OAI21_X1 U5075 ( .B1(n2228), .B2(n4557), .A(n4440), .ZN(n4619) );
  INV_X1 U5076 ( .A(n4441), .ZN(n4442) );
  AOI22_X1 U5077 ( .A1(n4781), .A2(REG2_REG_21__SCAN_IN), .B1(n4442), .B2(
        n4785), .ZN(n4443) );
  OAI21_X1 U5078 ( .B1(n4558), .B2(n4444), .A(n4443), .ZN(n4445) );
  AOI21_X1 U5079 ( .B1(n4447), .B2(n4446), .A(n4445), .ZN(n4448) );
  OAI21_X1 U5080 ( .B1(n4619), .B2(n4493), .A(n4448), .ZN(n4449) );
  AOI21_X1 U5081 ( .B1(n4560), .B2(n4517), .A(n4449), .ZN(n4450) );
  OAI21_X1 U5082 ( .B1(n4451), .B2(n4521), .A(n4450), .ZN(U3269) );
  XNOR2_X1 U5083 ( .A(n4452), .B(n4455), .ZN(n4464) );
  NAND2_X1 U5084 ( .A1(n4454), .A2(n4453), .ZN(n4456) );
  XNOR2_X1 U5085 ( .A(n4456), .B(n4455), .ZN(n4461) );
  OAI22_X1 U5086 ( .A1(n4458), .A2(n4482), .B1(n4457), .B2(n4577), .ZN(n4459)
         );
  AOI21_X1 U5087 ( .B1(n4506), .B2(n4509), .A(n4459), .ZN(n4460) );
  OAI21_X1 U5088 ( .B1(n4461), .B2(n4486), .A(n4460), .ZN(n4462) );
  AOI21_X1 U5089 ( .B1(n4464), .B2(n4463), .A(n4462), .ZN(n4567) );
  INV_X1 U5090 ( .A(n4464), .ZN(n4568) );
  AOI22_X1 U5091 ( .A1(n4781), .A2(REG2_REG_20__SCAN_IN), .B1(n4465), .B2(
        n4785), .ZN(n4468) );
  NAND2_X1 U5092 ( .A1(n4490), .A2(n4466), .ZN(n4564) );
  NAND3_X1 U5093 ( .A1(n4565), .A2(n4776), .A3(n4564), .ZN(n4467) );
  OAI211_X1 U5094 ( .C1(n4568), .C2(n4469), .A(n4468), .B(n4467), .ZN(n4470)
         );
  INV_X1 U5095 ( .A(n4470), .ZN(n4471) );
  OAI21_X1 U5096 ( .B1(n4781), .B2(n4567), .A(n4471), .ZN(U3270) );
  NAND2_X1 U5097 ( .A1(n4498), .A2(n4472), .ZN(n4473) );
  XNOR2_X1 U5098 ( .A(n4473), .B(n4480), .ZN(n4570) );
  INV_X1 U5099 ( .A(n4570), .ZN(n4496) );
  INV_X1 U5100 ( .A(n4474), .ZN(n4475) );
  NOR2_X1 U5101 ( .A1(n4476), .A2(n4475), .ZN(n4505) );
  INV_X1 U5102 ( .A(n4477), .ZN(n4478) );
  AOI21_X1 U5103 ( .B1(n4505), .B2(n4479), .A(n4478), .ZN(n4481) );
  XNOR2_X1 U5104 ( .A(n4481), .B(n4480), .ZN(n4487) );
  OAI22_X1 U5105 ( .A1(n4558), .A2(n4482), .B1(n4577), .B2(n4488), .ZN(n4483)
         );
  AOI21_X1 U5106 ( .B1(n4506), .B2(n4484), .A(n4483), .ZN(n4485) );
  OAI21_X1 U5107 ( .B1(n4487), .B2(n4486), .A(n4485), .ZN(n4569) );
  OR2_X1 U5108 ( .A1(n4501), .A2(n4488), .ZN(n4489) );
  NAND2_X1 U5109 ( .A1(n4490), .A2(n4489), .ZN(n4623) );
  AOI22_X1 U5110 ( .A1(n4781), .A2(REG2_REG_19__SCAN_IN), .B1(n4491), .B2(
        n4785), .ZN(n4492) );
  OAI21_X1 U5111 ( .B1(n4623), .B2(n4493), .A(n4492), .ZN(n4494) );
  AOI21_X1 U5112 ( .B1(n4569), .B2(n4517), .A(n4494), .ZN(n4495) );
  OAI21_X1 U5113 ( .B1(n4496), .B2(n4521), .A(n4495), .ZN(U3271) );
  OAI21_X1 U5114 ( .B1(n4497), .B2(n4504), .A(n4498), .ZN(n4499) );
  INV_X1 U5115 ( .A(n4499), .ZN(n4575) );
  AOI22_X1 U5116 ( .A1(n4781), .A2(REG2_REG_18__SCAN_IN), .B1(n4500), .B2(
        n4785), .ZN(n4520) );
  INV_X1 U5117 ( .A(n4501), .ZN(n4502) );
  OAI211_X1 U5118 ( .C1(n4503), .C2(n4512), .A(n4502), .B(n4829), .ZN(n4573)
         );
  XNOR2_X1 U5119 ( .A(n4505), .B(n4504), .ZN(n4515) );
  NAND2_X1 U5120 ( .A1(n4507), .A2(n4506), .ZN(n4511) );
  NAND2_X1 U5121 ( .A1(n4509), .A2(n4508), .ZN(n4510) );
  OAI211_X1 U5122 ( .C1(n4577), .C2(n4512), .A(n4511), .B(n4510), .ZN(n4513)
         );
  AOI21_X1 U5123 ( .B1(n4515), .B2(n4514), .A(n4513), .ZN(n4574) );
  OAI21_X1 U5124 ( .B1(n4516), .B2(n4573), .A(n4574), .ZN(n4518) );
  NAND2_X1 U5125 ( .A1(n4518), .A2(n4517), .ZN(n4519) );
  OAI211_X1 U5126 ( .C1(n4575), .C2(n4521), .A(n4520), .B(n4519), .ZN(U3272)
         );
  AOI21_X1 U5127 ( .B1(n4525), .B2(n4522), .A(n4655), .ZN(n4662) );
  INV_X1 U5128 ( .A(n4662), .ZN(n4594) );
  AND2_X1 U5129 ( .A1(n4524), .A2(n4523), .ZN(n4657) );
  AOI21_X1 U5130 ( .B1(n4525), .B2(n4658), .A(n4657), .ZN(n4664) );
  MUX2_X1 U5131 ( .A(n2735), .B(n4664), .S(n4867), .Z(n4526) );
  OAI21_X1 U5132 ( .B1(n4594), .B2(n4585), .A(n4526), .ZN(U3548) );
  OAI22_X1 U5133 ( .A1(n4528), .A2(n4578), .B1(n4527), .B2(n4577), .ZN(n4529)
         );
  AOI211_X1 U5134 ( .C1(n4531), .C2(n4856), .A(n4530), .B(n4529), .ZN(n4595)
         );
  MUX2_X1 U5135 ( .A(n4532), .B(n4595), .S(n4867), .Z(n4533) );
  OAI21_X1 U5136 ( .B1(n4585), .B2(n4598), .A(n4533), .ZN(U3545) );
  AOI21_X1 U5137 ( .B1(n4535), .B2(n4856), .A(n4534), .ZN(n4599) );
  MUX2_X1 U5138 ( .A(n4536), .B(n4599), .S(n4867), .Z(n4537) );
  OAI21_X1 U5139 ( .B1(n4585), .B2(n4602), .A(n4537), .ZN(U3544) );
  AOI21_X1 U5140 ( .B1(n4539), .B2(n4856), .A(n4538), .ZN(n4603) );
  MUX2_X1 U5141 ( .A(n4540), .B(n4603), .S(n4867), .Z(n4541) );
  OAI21_X1 U5142 ( .B1(n4585), .B2(n4605), .A(n4541), .ZN(U3543) );
  OAI22_X1 U5143 ( .A1(n4543), .A2(n4578), .B1(n4542), .B2(n4577), .ZN(n4544)
         );
  AOI211_X1 U5144 ( .C1(n4546), .C2(n4856), .A(n4545), .B(n4544), .ZN(n4606)
         );
  MUX2_X1 U5145 ( .A(n4547), .B(n4606), .S(n4867), .Z(n4548) );
  OAI21_X1 U5146 ( .B1(n4585), .B2(n4609), .A(n4548), .ZN(U3542) );
  AOI21_X1 U5147 ( .B1(n4550), .B2(n4856), .A(n4549), .ZN(n4610) );
  MUX2_X1 U5148 ( .A(n3389), .B(n4610), .S(n4867), .Z(n4551) );
  OAI21_X1 U5149 ( .B1(n4585), .B2(n4612), .A(n4551), .ZN(U3541) );
  OR2_X1 U5150 ( .A1(n4552), .A2(n4590), .ZN(n4554) );
  AND2_X1 U5151 ( .A1(n4554), .A2(n4553), .ZN(n4613) );
  MUX2_X1 U5152 ( .A(n4555), .B(n4613), .S(n4867), .Z(n4556) );
  OAI21_X1 U5153 ( .B1(n4585), .B2(n4616), .A(n4556), .ZN(U3540) );
  OAI22_X1 U5154 ( .A1(n4558), .A2(n4578), .B1(n4577), .B2(n4557), .ZN(n4559)
         );
  AOI211_X1 U5155 ( .C1(n4561), .C2(n4856), .A(n4560), .B(n4559), .ZN(n4617)
         );
  MUX2_X1 U5156 ( .A(n4562), .B(n4617), .S(n4867), .Z(n4563) );
  OAI21_X1 U5157 ( .B1(n4585), .B2(n4619), .A(n4563), .ZN(U3539) );
  NAND3_X1 U5158 ( .A1(n4565), .A2(n4829), .A3(n4564), .ZN(n4566) );
  OAI211_X1 U5159 ( .C1(n4568), .C2(n4831), .A(n4567), .B(n4566), .ZN(n4620)
         );
  MUX2_X1 U5160 ( .A(REG1_REG_20__SCAN_IN), .B(n4620), .S(n4867), .Z(U3538) );
  AOI21_X1 U5161 ( .B1(n4570), .B2(n4856), .A(n4569), .ZN(n4621) );
  MUX2_X1 U5162 ( .A(n4571), .B(n4621), .S(n4867), .Z(n4572) );
  OAI21_X1 U5163 ( .B1(n4585), .B2(n4623), .A(n4572), .ZN(U3537) );
  OAI211_X1 U5164 ( .C1(n4575), .C2(n4590), .A(n4574), .B(n4573), .ZN(n4624)
         );
  MUX2_X1 U5165 ( .A(REG1_REG_18__SCAN_IN), .B(n4624), .S(n4867), .Z(U3536) );
  OAI22_X1 U5166 ( .A1(n4579), .A2(n4578), .B1(n4577), .B2(n4576), .ZN(n4580)
         );
  AOI211_X1 U5167 ( .C1(n4582), .C2(n4856), .A(n4581), .B(n4580), .ZN(n4625)
         );
  MUX2_X1 U5168 ( .A(n4583), .B(n4625), .S(n4867), .Z(n4584) );
  OAI21_X1 U5169 ( .B1(n4585), .B2(n4629), .A(n4584), .ZN(U3535) );
  NAND3_X1 U5170 ( .A1(n4587), .A2(n4829), .A3(n4586), .ZN(n4588) );
  OAI211_X1 U5171 ( .C1(n4591), .C2(n4590), .A(n4589), .B(n4588), .ZN(n4630)
         );
  MUX2_X1 U5172 ( .A(REG1_REG_16__SCAN_IN), .B(n4630), .S(n4867), .Z(U3534) );
  INV_X1 U5173 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4592) );
  MUX2_X1 U5174 ( .A(n4592), .B(n4664), .S(n4860), .Z(n4593) );
  OAI21_X1 U5175 ( .B1(n4594), .B2(n4628), .A(n4593), .ZN(U3516) );
  INV_X1 U5176 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4596) );
  MUX2_X1 U5177 ( .A(n4596), .B(n4595), .S(n4860), .Z(n4597) );
  OAI21_X1 U5178 ( .B1(n4598), .B2(n4628), .A(n4597), .ZN(U3513) );
  INV_X1 U5179 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4600) );
  MUX2_X1 U5180 ( .A(n4600), .B(n4599), .S(n4860), .Z(n4601) );
  OAI21_X1 U5181 ( .B1(n4602), .B2(n4628), .A(n4601), .ZN(U3512) );
  MUX2_X1 U5182 ( .A(n3395), .B(n4603), .S(n4860), .Z(n4604) );
  OAI21_X1 U5183 ( .B1(n4605), .B2(n4628), .A(n4604), .ZN(U3511) );
  INV_X1 U5184 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4607) );
  MUX2_X1 U5185 ( .A(n4607), .B(n4606), .S(n4860), .Z(n4608) );
  OAI21_X1 U5186 ( .B1(n4609), .B2(n4628), .A(n4608), .ZN(U3510) );
  MUX2_X1 U5187 ( .A(n3388), .B(n4610), .S(n4860), .Z(n4611) );
  OAI21_X1 U5188 ( .B1(n4612), .B2(n4628), .A(n4611), .ZN(U3509) );
  MUX2_X1 U5189 ( .A(n4614), .B(n4613), .S(n4860), .Z(n4615) );
  OAI21_X1 U5190 ( .B1(n4616), .B2(n4628), .A(n4615), .ZN(U3508) );
  MUX2_X1 U5191 ( .A(n3382), .B(n4617), .S(n4860), .Z(n4618) );
  OAI21_X1 U5192 ( .B1(n4619), .B2(n4628), .A(n4618), .ZN(U3507) );
  MUX2_X1 U5193 ( .A(REG0_REG_20__SCAN_IN), .B(n4620), .S(n4860), .Z(U3506) );
  MUX2_X1 U5194 ( .A(n3505), .B(n4621), .S(n4860), .Z(n4622) );
  OAI21_X1 U5195 ( .B1(n4623), .B2(n4628), .A(n4622), .ZN(U3505) );
  MUX2_X1 U5196 ( .A(REG0_REG_18__SCAN_IN), .B(n4624), .S(n4860), .Z(U3503) );
  INV_X1 U5197 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4626) );
  MUX2_X1 U5198 ( .A(n4626), .B(n4625), .S(n4860), .Z(n4627) );
  OAI21_X1 U5199 ( .B1(n4629), .B2(n4628), .A(n4627), .ZN(U3501) );
  MUX2_X1 U5200 ( .A(REG0_REG_16__SCAN_IN), .B(n4630), .S(n4860), .Z(U3499) );
  MUX2_X1 U5201 ( .A(n2678), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5202 ( .A(DATAI_22_), .B(n4631), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U5203 ( .A(DATAI_20_), .B(n4632), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5204 ( .A(DATAI_18_), .B(n4641), .S(STATE_REG_SCAN_IN), .Z(U3334)
         );
  MUX2_X1 U5205 ( .A(DATAI_8_), .B(n4633), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U5206 ( .A(n4634), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5207 ( .A(n4635), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5208 ( .A(DATAI_2_), .B(n2412), .S(STATE_REG_SCAN_IN), .Z(U3350) );
  MUX2_X1 U5209 ( .A(n4636), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  AOI21_X1 U5210 ( .B1(n4641), .B2(REG2_REG_18__SCAN_IN), .A(n4637), .ZN(n4640) );
  INV_X1 U5211 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4638) );
  MUX2_X1 U5212 ( .A(REG2_REG_19__SCAN_IN), .B(n4638), .S(n4648), .Z(n4639) );
  XNOR2_X1 U5213 ( .A(n4640), .B(n4639), .ZN(n4652) );
  MUX2_X1 U5214 ( .A(REG1_REG_19__SCAN_IN), .B(n4571), .S(n4648), .Z(n4645) );
  AOI22_X1 U5215 ( .A1(n4643), .A2(n4642), .B1(REG1_REG_18__SCAN_IN), .B2(
        n4641), .ZN(n4644) );
  XOR2_X1 U5216 ( .A(n4645), .B(n4644), .Z(n4650) );
  NAND2_X1 U5217 ( .A1(n4768), .A2(ADDR_REG_19__SCAN_IN), .ZN(n4646) );
  OAI211_X1 U5218 ( .C1(n4775), .C2(n4648), .A(n4647), .B(n4646), .ZN(n4649)
         );
  AOI21_X1 U5219 ( .B1(n4650), .B2(n4769), .A(n4649), .ZN(n4651) );
  OAI21_X1 U5220 ( .B1(n4652), .B2(n4762), .A(n4651), .ZN(U3259) );
  INV_X1 U5221 ( .A(DATAI_28_), .ZN(n4653) );
  AOI22_X1 U5222 ( .A1(STATE_REG_SCAN_IN), .A2(n4654), .B1(n4653), .B2(U3149), 
        .ZN(U3324) );
  INV_X1 U5223 ( .A(n4656), .ZN(n4659) );
  AOI21_X1 U5224 ( .B1(n4659), .B2(n4658), .A(n4657), .ZN(n4670) );
  INV_X1 U5225 ( .A(n4670), .ZN(n4665) );
  AOI22_X1 U5226 ( .A1(n4668), .A2(n4776), .B1(n4517), .B2(n4665), .ZN(n4660)
         );
  OAI21_X1 U5227 ( .B1(n4517), .B2(n4661), .A(n4660), .ZN(U3260) );
  AOI22_X1 U5228 ( .A1(n4662), .A2(n4776), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4781), .ZN(n4663) );
  OAI21_X1 U5229 ( .B1(n4781), .B2(n4664), .A(n4663), .ZN(U3261) );
  AOI22_X1 U5230 ( .A1(n4668), .A2(n4666), .B1(n4867), .B2(n4665), .ZN(n4667)
         );
  OAI21_X1 U5231 ( .B1(n4867), .B2(n3145), .A(n4667), .ZN(U3549) );
  AOI22_X1 U5232 ( .A1(n4668), .A2(n4837), .B1(REG0_REG_31__SCAN_IN), .B2(
        n4858), .ZN(n4669) );
  OAI21_X1 U5233 ( .B1(n4670), .B2(n4858), .A(n4669), .ZN(U3517) );
  OAI21_X1 U5234 ( .B1(REG1_REG_0__SCAN_IN), .B2(n4672), .A(n4671), .ZN(n4673)
         );
  XNOR2_X1 U5235 ( .A(IR_REG_0__SCAN_IN), .B(n4673), .ZN(n4674) );
  AOI22_X1 U5236 ( .A1(n4675), .A2(n4674), .B1(n4768), .B2(ADDR_REG_0__SCAN_IN), .ZN(n4676) );
  OAI21_X1 U5237 ( .B1(STATE_REG_SCAN_IN), .B2(n4677), .A(n4676), .ZN(U3240)
         );
  OAI211_X1 U5238 ( .C1(n4680), .C2(n4679), .A(n4769), .B(n4678), .ZN(n4685)
         );
  OAI211_X1 U5239 ( .C1(n4683), .C2(n4682), .A(n4711), .B(n4681), .ZN(n4684)
         );
  OAI211_X1 U5240 ( .C1(n4775), .C2(n4824), .A(n4685), .B(n4684), .ZN(n4686)
         );
  AOI211_X1 U5241 ( .C1(n4768), .C2(ADDR_REG_9__SCAN_IN), .A(n4687), .B(n4686), 
        .ZN(n4688) );
  INV_X1 U5242 ( .A(n4688), .ZN(U3249) );
  OAI211_X1 U5243 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4690), .A(n4769), .B(n4689), .ZN(n4694) );
  OAI211_X1 U5244 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4692), .A(n4711), .B(n4691), .ZN(n4693) );
  OAI211_X1 U5245 ( .C1(n4775), .C2(n4822), .A(n4694), .B(n4693), .ZN(n4695)
         );
  AOI211_X1 U5246 ( .C1(n4768), .C2(ADDR_REG_10__SCAN_IN), .A(n4696), .B(n4695), .ZN(n4697) );
  INV_X1 U5247 ( .A(n4697), .ZN(U3250) );
  OAI211_X1 U5248 ( .C1(n4700), .C2(n4699), .A(n4769), .B(n4698), .ZN(n4705)
         );
  OAI211_X1 U5249 ( .C1(n4703), .C2(n4702), .A(n4711), .B(n4701), .ZN(n4704)
         );
  OAI211_X1 U5250 ( .C1(n4775), .C2(n4820), .A(n4705), .B(n4704), .ZN(n4706)
         );
  AOI211_X1 U5251 ( .C1(n4768), .C2(ADDR_REG_11__SCAN_IN), .A(n4707), .B(n4706), .ZN(n4708) );
  INV_X1 U5252 ( .A(n4708), .ZN(U3251) );
  OAI211_X1 U5253 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4712), .A(n4711), .B(n4710), .ZN(n4714) );
  NAND2_X1 U5254 ( .A1(n4714), .A2(n4713), .ZN(n4715) );
  AOI21_X1 U5255 ( .B1(n4768), .B2(ADDR_REG_12__SCAN_IN), .A(n4715), .ZN(n4719) );
  OAI211_X1 U5256 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4717), .A(n4769), .B(n4716), .ZN(n4718) );
  OAI211_X1 U5257 ( .C1(n4775), .C2(n2286), .A(n4719), .B(n4718), .ZN(U3252)
         );
  AOI21_X1 U5258 ( .B1(n4721), .B2(n4818), .A(n4720), .ZN(n4724) );
  NOR2_X1 U5259 ( .A1(n4724), .A2(n4723), .ZN(n4722) );
  AOI211_X1 U5260 ( .C1(n4724), .C2(n4723), .A(n4762), .B(n4722), .ZN(n4725)
         );
  AOI211_X1 U5261 ( .C1(n4768), .C2(ADDR_REG_13__SCAN_IN), .A(n4726), .B(n4725), .ZN(n4731) );
  OAI211_X1 U5262 ( .C1(n4729), .C2(n4728), .A(n4769), .B(n4727), .ZN(n4730)
         );
  OAI211_X1 U5263 ( .C1(n4775), .C2(n4818), .A(n4731), .B(n4730), .ZN(U3253)
         );
  NOR2_X1 U5264 ( .A1(STATE_REG_SCAN_IN), .A2(n4732), .ZN(n4737) );
  AOI211_X1 U5265 ( .C1(n4735), .C2(n4734), .A(n4733), .B(n4762), .ZN(n4736)
         );
  AOI211_X1 U5266 ( .C1(n4768), .C2(ADDR_REG_14__SCAN_IN), .A(n4737), .B(n4736), .ZN(n4741) );
  OAI211_X1 U5267 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4739), .A(n4769), .B(n4738), .ZN(n4740) );
  OAI211_X1 U5268 ( .C1(n4775), .C2(n4816), .A(n4741), .B(n4740), .ZN(U3254)
         );
  AOI211_X1 U5269 ( .C1(n4744), .C2(n4743), .A(n4742), .B(n4762), .ZN(n4745)
         );
  AOI211_X1 U5270 ( .C1(n4768), .C2(ADDR_REG_15__SCAN_IN), .A(n4746), .B(n4745), .ZN(n4751) );
  OAI211_X1 U5271 ( .C1(n4749), .C2(n4748), .A(n4769), .B(n4747), .ZN(n4750)
         );
  OAI211_X1 U5272 ( .C1(n4775), .C2(n4814), .A(n4751), .B(n4750), .ZN(U3255)
         );
  INV_X1 U5273 ( .A(n4752), .ZN(n4757) );
  AOI221_X1 U5274 ( .B1(n4755), .B2(n4754), .C1(n4753), .C2(n4754), .A(n4762), 
        .ZN(n4756) );
  AOI211_X1 U5275 ( .C1(n4768), .C2(ADDR_REG_16__SCAN_IN), .A(n4757), .B(n4756), .ZN(n4761) );
  OAI221_X1 U5276 ( .B1(n4759), .B2(REG1_REG_16__SCAN_IN), .C1(n4759), .C2(
        n4758), .A(n4769), .ZN(n4760) );
  OAI211_X1 U5277 ( .C1(n4775), .C2(n4812), .A(n4761), .B(n4760), .ZN(U3256)
         );
  AOI221_X1 U5278 ( .B1(n4765), .B2(n4764), .C1(n4763), .C2(n4764), .A(n4762), 
        .ZN(n4766) );
  AOI211_X1 U5279 ( .C1(n4768), .C2(ADDR_REG_17__SCAN_IN), .A(n4767), .B(n4766), .ZN(n4774) );
  OAI221_X1 U5280 ( .B1(n4772), .B2(n4771), .C1(n4772), .C2(n4770), .A(n4769), 
        .ZN(n4773) );
  OAI211_X1 U5281 ( .C1(n4775), .C2(n4810), .A(n4774), .B(n4773), .ZN(U3257)
         );
  AOI22_X1 U5282 ( .A1(REG2_REG_2__SCAN_IN), .A2(n4781), .B1(
        REG3_REG_2__SCAN_IN), .B2(n4785), .ZN(n4779) );
  AOI22_X1 U5283 ( .A1(n4777), .A2(n4786), .B1(n4776), .B2(n4836), .ZN(n4778)
         );
  OAI211_X1 U5284 ( .C1(n4781), .C2(n4780), .A(n4779), .B(n4778), .ZN(U3288)
         );
  AOI21_X1 U5285 ( .B1(n4784), .B2(n4783), .A(n4782), .ZN(n4790) );
  AOI22_X1 U5286 ( .A1(n4787), .A2(n4786), .B1(REG3_REG_0__SCAN_IN), .B2(n4785), .ZN(n4788) );
  OAI221_X1 U5287 ( .B1(n4781), .B2(n4790), .C1(n4517), .C2(n4789), .A(n4788), 
        .ZN(U3290) );
  NOR2_X1 U5288 ( .A1(n4805), .A2(n4791), .ZN(U3291) );
  AND2_X1 U5289 ( .A1(D_REG_30__SCAN_IN), .A2(n4806), .ZN(U3292) );
  AND2_X1 U5290 ( .A1(D_REG_29__SCAN_IN), .A2(n4806), .ZN(U3293) );
  NOR2_X1 U5291 ( .A1(n4805), .A2(n4792), .ZN(U3294) );
  NOR2_X1 U5292 ( .A1(n4805), .A2(n4793), .ZN(U3295) );
  NOR2_X1 U5293 ( .A1(n4805), .A2(n4794), .ZN(U3296) );
  AND2_X1 U5294 ( .A1(D_REG_25__SCAN_IN), .A2(n4806), .ZN(U3297) );
  AND2_X1 U5295 ( .A1(D_REG_24__SCAN_IN), .A2(n4806), .ZN(U3298) );
  NOR2_X1 U5296 ( .A1(n4805), .A2(n4795), .ZN(U3299) );
  NOR2_X1 U5297 ( .A1(n4805), .A2(n4796), .ZN(U3300) );
  NOR2_X1 U5298 ( .A1(n4805), .A2(n4797), .ZN(U3301) );
  AND2_X1 U5299 ( .A1(D_REG_20__SCAN_IN), .A2(n4806), .ZN(U3302) );
  NOR2_X1 U5300 ( .A1(n4805), .A2(n4798), .ZN(U3303) );
  NOR2_X1 U5301 ( .A1(n4805), .A2(n4799), .ZN(U3304) );
  NOR2_X1 U5302 ( .A1(n4805), .A2(n4800), .ZN(U3305) );
  AND2_X1 U5303 ( .A1(D_REG_16__SCAN_IN), .A2(n4806), .ZN(U3306) );
  AND2_X1 U5304 ( .A1(D_REG_15__SCAN_IN), .A2(n4806), .ZN(U3307) );
  AND2_X1 U5305 ( .A1(D_REG_14__SCAN_IN), .A2(n4806), .ZN(U3308) );
  AND2_X1 U5306 ( .A1(D_REG_13__SCAN_IN), .A2(n4806), .ZN(U3309) );
  AND2_X1 U5307 ( .A1(D_REG_12__SCAN_IN), .A2(n4806), .ZN(U3310) );
  AND2_X1 U5308 ( .A1(D_REG_11__SCAN_IN), .A2(n4806), .ZN(U3311) );
  NOR2_X1 U5309 ( .A1(n4805), .A2(n4801), .ZN(U3312) );
  NOR2_X1 U5310 ( .A1(n4805), .A2(n4802), .ZN(U3313) );
  AND2_X1 U5311 ( .A1(D_REG_8__SCAN_IN), .A2(n4806), .ZN(U3314) );
  AND2_X1 U5312 ( .A1(D_REG_7__SCAN_IN), .A2(n4806), .ZN(U3315) );
  AND2_X1 U5313 ( .A1(D_REG_6__SCAN_IN), .A2(n4806), .ZN(U3316) );
  NOR2_X1 U5314 ( .A1(n4805), .A2(n4803), .ZN(U3317) );
  AND2_X1 U5315 ( .A1(D_REG_4__SCAN_IN), .A2(n4806), .ZN(U3318) );
  NOR2_X1 U5316 ( .A1(n4805), .A2(n4804), .ZN(U3319) );
  AND2_X1 U5317 ( .A1(D_REG_2__SCAN_IN), .A2(n4806), .ZN(U3320) );
  AOI21_X1 U5318 ( .B1(U3149), .B2(n4808), .A(n4807), .ZN(U3329) );
  AOI22_X1 U5319 ( .A1(STATE_REG_SCAN_IN), .A2(n4810), .B1(n4809), .B2(U3149), 
        .ZN(U3335) );
  AOI22_X1 U5320 ( .A1(STATE_REG_SCAN_IN), .A2(n4812), .B1(n4811), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5321 ( .A(DATAI_15_), .ZN(n4813) );
  AOI22_X1 U5322 ( .A1(STATE_REG_SCAN_IN), .A2(n4814), .B1(n4813), .B2(U3149), 
        .ZN(U3337) );
  AOI22_X1 U5323 ( .A1(STATE_REG_SCAN_IN), .A2(n4816), .B1(n4815), .B2(U3149), 
        .ZN(U3338) );
  AOI22_X1 U5324 ( .A1(STATE_REG_SCAN_IN), .A2(n4818), .B1(n4817), .B2(U3149), 
        .ZN(U3339) );
  INV_X1 U5325 ( .A(DATAI_12_), .ZN(n4819) );
  AOI22_X1 U5326 ( .A1(STATE_REG_SCAN_IN), .A2(n2286), .B1(n4819), .B2(U3149), 
        .ZN(U3340) );
  AOI22_X1 U5327 ( .A1(STATE_REG_SCAN_IN), .A2(n4820), .B1(n2508), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5328 ( .A(DATAI_10_), .ZN(n4821) );
  AOI22_X1 U5329 ( .A1(STATE_REG_SCAN_IN), .A2(n4822), .B1(n4821), .B2(U3149), 
        .ZN(U3342) );
  AOI22_X1 U5330 ( .A1(STATE_REG_SCAN_IN), .A2(n4824), .B1(n4823), .B2(U3149), 
        .ZN(U3343) );
  INV_X1 U5331 ( .A(DATAI_0_), .ZN(n4825) );
  AOI22_X1 U5332 ( .A1(STATE_REG_SCAN_IN), .A2(n4826), .B1(n4825), .B2(U3149), 
        .ZN(U3352) );
  AOI22_X1 U5333 ( .A1(n4860), .A2(n4828), .B1(n4827), .B2(n4858), .ZN(U3467)
         );
  OAI22_X1 U5334 ( .A1(n4832), .A2(n4831), .B1(n2782), .B2(n4830), .ZN(n4833)
         );
  NOR2_X1 U5335 ( .A1(n4834), .A2(n4833), .ZN(n4862) );
  INV_X1 U5336 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4835) );
  AOI22_X1 U5337 ( .A1(n4860), .A2(n4862), .B1(n4835), .B2(n4858), .ZN(U3469)
         );
  AOI22_X1 U5338 ( .A1(n4838), .A2(n4860), .B1(n4837), .B2(n4836), .ZN(n4839)
         );
  OAI21_X1 U5339 ( .B1(n4860), .B2(n4840), .A(n4839), .ZN(U3471) );
  INV_X1 U5340 ( .A(n4841), .ZN(n4843) );
  AOI211_X1 U5341 ( .C1(n4845), .C2(n4844), .A(n4843), .B(n4842), .ZN(n4863)
         );
  AOI22_X1 U5342 ( .A1(n4860), .A2(n4863), .B1(n4846), .B2(n4858), .ZN(U3475)
         );
  NAND3_X1 U5343 ( .A1(n4848), .A2(n4847), .A3(n4856), .ZN(n4849) );
  AND3_X1 U5344 ( .A1(n4851), .A2(n4850), .A3(n4849), .ZN(n4864) );
  INV_X1 U5345 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4852) );
  AOI22_X1 U5346 ( .A1(n4860), .A2(n4864), .B1(n4852), .B2(n4858), .ZN(U3481)
         );
  NOR3_X1 U5347 ( .A1(n4853), .A2(n2227), .A3(n2782), .ZN(n4855) );
  AOI211_X1 U5348 ( .C1(n4857), .C2(n4856), .A(n4855), .B(n4854), .ZN(n4866)
         );
  INV_X1 U5349 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4859) );
  AOI22_X1 U5350 ( .A1(n4860), .A2(n4866), .B1(n4859), .B2(n4858), .ZN(U3491)
         );
  INV_X1 U5351 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4861) );
  AOI22_X1 U5352 ( .A1(n4867), .A2(n4862), .B1(n4861), .B2(n4865), .ZN(U3519)
         );
  AOI22_X1 U5353 ( .A1(n4867), .A2(n4863), .B1(n2414), .B2(n4865), .ZN(U3522)
         );
  AOI22_X1 U5354 ( .A1(n4867), .A2(n4864), .B1(n3156), .B2(n4865), .ZN(U3525)
         );
  AOI22_X1 U5355 ( .A1(n4867), .A2(n4866), .B1(n2513), .B2(n4865), .ZN(U3530)
         );
  INV_X2 U2436 ( .A(n2783), .ZN(n2804) );
  NOR2_X1 U2463 ( .A1(IR_REG_4__SCAN_IN), .A2(IR_REG_3__SCAN_IN), .ZN(n2224)
         );
  CLKBUF_X1 U2904 ( .A(n2404), .Z(n3146) );
endmodule

