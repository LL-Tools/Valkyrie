

module b22_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, 
        SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, 
        SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, 
        SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, 
        P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
         n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
         n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
         n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
         n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
         n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
         n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
         n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
         n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
         n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
         n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
         n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
         n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
         n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
         n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
         n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
         n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973,
         n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981,
         n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
         n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
         n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
         n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
         n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125,
         n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
         n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
         n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
         n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
         n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
         n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173,
         n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
         n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189,
         n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197,
         n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
         n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
         n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
         n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
         n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
         n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245,
         n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
         n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261,
         n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
         n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
         n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
         n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
         n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
         n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
         n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
         n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
         n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333,
         n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341,
         n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349,
         n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
         n16358, n16359, n16360, n16361, n16362;

  OR2_X1 U7516 ( .A1(n9131), .A2(n8933), .ZN(n8934) );
  INV_X1 U7517 ( .A(n14176), .ZN(n8307) );
  XNOR2_X1 U7519 ( .A(n8918), .B(n8917), .ZN(n13372) );
  AOI21_X1 U7520 ( .B1(n15436), .B2(n13359), .A(n13358), .ZN(n15424) );
  INV_X1 U7521 ( .A(n10312), .ZN(n12412) );
  BUF_X2 U7522 ( .A(n10327), .Z(n7425) );
  NAND2_X1 U7523 ( .A1(n11131), .A2(n10420), .ZN(n10322) );
  INV_X2 U7524 ( .A(n8952), .ZN(n8948) );
  CLKBUF_X2 U7525 ( .A(n8761), .Z(n8922) );
  NAND4_X1 U7526 ( .A1(n8742), .A2(n8741), .A3(n8740), .A4(n8739), .ZN(n15194)
         );
  INV_X1 U7527 ( .A(n8750), .ZN(n8926) );
  INV_X1 U7528 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n10646) );
  INV_X1 U7529 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n11221) );
  OAI21_X1 U7530 ( .B1(n9042), .B2(n8244), .A(n7651), .ZN(n7893) );
  NOR2_X1 U7531 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n10092) );
  AND3_X1 U7532 ( .A1(n7793), .A2(n10094), .A3(n10093), .ZN(n8077) );
  INV_X1 U7533 ( .A(n13594), .ZN(n13578) );
  NAND2_X1 U7534 ( .A1(n10872), .A2(n10877), .ZN(n8954) );
  INV_X1 U7535 ( .A(n13927), .ZN(n9276) );
  NAND2_X1 U7536 ( .A1(n14279), .A2(n7542), .ZN(n14278) );
  NAND2_X1 U7537 ( .A1(n14352), .A2(n14174), .ZN(n9932) );
  INV_X1 U7538 ( .A(n10129), .ZN(n10043) );
  BUF_X1 U7539 ( .A(n11125), .Z(n14525) );
  OR2_X1 U7540 ( .A1(n14975), .A2(n14845), .ZN(n14824) );
  CLKBUF_X3 U7541 ( .A(n10322), .Z(n13618) );
  INV_X1 U7542 ( .A(n15193), .ZN(n11297) );
  NAND2_X1 U7543 ( .A1(n15606), .A2(n15244), .ZN(n10877) );
  OR2_X1 U7544 ( .A1(n9571), .A2(n11438), .ZN(n9280) );
  NAND2_X1 U7545 ( .A1(n14212), .A2(n9671), .ZN(n14193) );
  INV_X1 U7546 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n9330) );
  OAI211_X1 U7547 ( .C1(n10312), .C2(n10465), .A(n8022), .B(n7959), .ZN(n13680) );
  OR2_X1 U7548 ( .A1(n15052), .A2(n10411), .ZN(n10268) );
  AND2_X1 U7550 ( .A1(n10294), .A2(n10295), .ZN(n10410) );
  INV_X1 U7551 ( .A(n8763), .ZN(n8750) );
  INV_X1 U7552 ( .A(n8750), .ZN(n8896) );
  INV_X1 U7553 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n7671) );
  NAND2_X1 U7554 ( .A1(n12259), .A2(n12258), .ZN(n12257) );
  CLKBUF_X3 U7555 ( .A(n9571), .Z(n9908) );
  NAND4_X1 U7556 ( .A1(n9282), .A2(n9281), .A3(n9280), .A4(n9279), .ZN(n9299)
         );
  OAI21_X1 U7557 ( .B1(n14349), .B2(n14341), .A(n7641), .ZN(n7640) );
  OR2_X1 U7558 ( .A1(n9273), .A2(n9330), .ZN(n9275) );
  NAND2_X1 U7559 ( .A1(n10327), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n10300) );
  NOR3_X1 U7560 ( .A1(n14785), .A2(n14944), .A3(n7968), .ZN(n14729) );
  NAND2_X1 U7561 ( .A1(n9695), .A2(n9694), .ZN(n14346) );
  INV_X1 U7562 ( .A(n16238), .ZN(n9764) );
  NAND4_X1 U7563 ( .A1(n11054), .A2(n11053), .A3(n11052), .A4(n11051), .ZN(
        n14687) );
  INV_X1 U7564 ( .A(n8847), .ZN(n15244) );
  XNOR2_X1 U7565 ( .A(n8518), .B(P1_IR_REG_19__SCAN_IN), .ZN(n8847) );
  AOI21_X2 U7566 ( .B1(n7997), .B2(n15973), .A(n7994), .ZN(n14154) );
  OAI21_X2 U7567 ( .B1(n12027), .B2(n8032), .A(n8029), .ZN(n12208) );
  NAND2_X2 U7568 ( .A1(n12025), .A2(n12024), .ZN(n12027) );
  OAI21_X2 U7569 ( .B1(n13838), .B2(n7805), .A(n7804), .ZN(n13843) );
  XNOR2_X2 U7570 ( .A(n10270), .B(P2_IR_REG_29__SCAN_IN), .ZN(n10272) );
  NAND2_X2 U7571 ( .A1(n10293), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10270) );
  NAND2_X2 U7572 ( .A1(n15082), .A2(n13274), .ZN(n13278) );
  NAND2_X2 U7573 ( .A1(n14980), .A2(n13541), .ZN(n14816) );
  NAND2_X2 U7574 ( .A1(n8162), .A2(n7531), .ZN(n14980) );
  NOR2_X2 U7575 ( .A1(n14065), .A2(n10124), .ZN(n10126) );
  NOR2_X2 U7576 ( .A1(n14067), .A2(n14066), .ZN(n14065) );
  XNOR2_X1 U7577 ( .A(n8771), .B(n8025), .ZN(n10465) );
  NAND2_X1 U7578 ( .A1(n11690), .A2(n11689), .ZN(n11692) );
  XNOR2_X2 U7579 ( .A(n15829), .B(n7925), .ZN(n15830) );
  NAND2_X2 U7580 ( .A1(n7926), .A2(n15820), .ZN(n15829) );
  XNOR2_X2 U7581 ( .A(n8473), .B(SI_24_), .ZN(n8877) );
  NAND2_X1 U7582 ( .A1(n11194), .A2(n7452), .ZN(n8081) );
  NOR2_X2 U7583 ( .A1(n11124), .A2(n11123), .ZN(n11194) );
  OAI222_X1 U7584 ( .A1(n10618), .A2(P1_U3086), .B1(n15604), .B2(n10465), .C1(
        n10464), .C2(n15597), .ZN(P1_U3354) );
  OAI222_X1 U7585 ( .A1(n15652), .A2(P2_U3088), .B1(n15061), .B2(n10465), .C1(
        n10452), .C2(n13255), .ZN(P2_U3326) );
  NOR2_X2 U7586 ( .A1(n7657), .A2(n7527), .ZN(n15339) );
  NOR2_X2 U7587 ( .A1(n15353), .A2(n15358), .ZN(n7657) );
  XNOR2_X2 U7588 ( .A(n9213), .B(n9212), .ZN(n13248) );
  NOR2_X2 U7589 ( .A1(n9379), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9392) );
  NAND2_X2 U7590 ( .A1(n10881), .A2(n12527), .ZN(n10878) );
  OR2_X2 U7591 ( .A1(n11090), .A2(n11438), .ZN(n11092) );
  NOR2_X2 U7592 ( .A1(n9448), .A2(n12155), .ZN(n12154) );
  XNOR2_X2 U7593 ( .A(n8526), .B(n8521), .ZN(n13616) );
  NAND2_X2 U7594 ( .A1(n8908), .A2(n8496), .ZN(n8526) );
  NOR2_X2 U7595 ( .A1(n14109), .A2(n14110), .ZN(n14115) );
  XNOR2_X1 U7596 ( .A(n10321), .B(n10320), .ZN(n14628) );
  NAND2_X2 U7597 ( .A1(n8015), .A2(n8012), .ZN(n15436) );
  OAI21_X4 U7598 ( .B1(n8660), .B2(n8441), .A(n8440), .ZN(n8442) );
  NOR2_X2 U7599 ( .A1(n16008), .A2(n9408), .ZN(n16007) );
  BUF_X2 U7600 ( .A(n9299), .Z(n16040) );
  XNOR2_X1 U7601 ( .A(n10291), .B(P2_IR_REG_19__SCAN_IN), .ZN(n10662) );
  OAI22_X2 U7602 ( .A1(n11670), .A2(n11669), .B1(n14649), .B2(n13631), .ZN(
        n11851) );
  XNOR2_X2 U7603 ( .A(n10117), .B(n16019), .ZN(n16008) );
  AND2_X2 U7604 ( .A1(n11375), .A2(n10116), .ZN(n10117) );
  XNOR2_X2 U7605 ( .A(n15192), .B(n8053), .ZN(n11488) );
  NAND4_X2 U7606 ( .A1(n8804), .A2(n8803), .A3(n8802), .A4(n8801), .ZN(n15192)
         );
  OAI21_X2 U7607 ( .B1(n8682), .B2(n8268), .A(n8265), .ZN(n8660) );
  OAI22_X2 U7608 ( .A1(n14532), .A2(n14533), .B1(n14511), .B2(n14510), .ZN(
        n14604) );
  XNOR2_X2 U7610 ( .A(n9218), .B(n9217), .ZN(n12383) );
  OAI21_X2 U7611 ( .B1(n9255), .B2(n8137), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n9218) );
  INV_X1 U7612 ( .A(n15516), .ZN(n7416) );
  INV_X1 U7613 ( .A(n7416), .ZN(n7417) );
  INV_X1 U7614 ( .A(n10170), .ZN(n10842) );
  NOR2_X2 U7615 ( .A1(n15798), .A2(n15799), .ZN(n15807) );
  NAND2_X2 U7616 ( .A1(n11546), .A2(n11545), .ZN(n13717) );
  AND2_X2 U7617 ( .A1(n15914), .A2(n15915), .ZN(n15917) );
  NAND2_X2 U7618 ( .A1(n8592), .A2(n8591), .ZN(n15528) );
  AOI21_X2 U7619 ( .B1(n7577), .B2(n7576), .A(n15789), .ZN(n15796) );
  AOI21_X1 U7620 ( .B1(n10054), .B2(n10076), .A(n10073), .ZN(n7732) );
  AOI21_X1 U7621 ( .B1(n7836), .B2(n14924), .A(n13528), .ZN(n14946) );
  OR2_X1 U7622 ( .A1(n14949), .A2(n14672), .ZN(n13512) );
  NOR2_X1 U7623 ( .A1(n8342), .A2(n7703), .ZN(n7702) );
  NAND2_X1 U7624 ( .A1(n7924), .A2(n15936), .ZN(n15943) );
  INV_X1 U7625 ( .A(n14949), .ZN(n7418) );
  NAND2_X1 U7626 ( .A1(n13375), .A2(n13374), .ZN(n14949) );
  OR3_X1 U7627 ( .A1(n13781), .A2(n8336), .A3(n13784), .ZN(n7809) );
  OR2_X1 U7628 ( .A1(n10126), .A2(n10125), .ZN(n10225) );
  NAND2_X1 U7629 ( .A1(n13449), .A2(n13448), .ZN(n14981) );
  OR2_X1 U7630 ( .A1(n11891), .A2(n13734), .ZN(n11892) );
  OAI22_X1 U7631 ( .A1(n8442), .A2(n7842), .B1(n7843), .B2(n7844), .ZN(n8449)
         );
  OR2_X1 U7632 ( .A1(n15992), .A2(n10114), .ZN(n7978) );
  NAND2_X1 U7633 ( .A1(n11205), .A2(n13625), .ZN(n11204) );
  CLKBUF_X2 U7634 ( .A(n9085), .Z(n7427) );
  INV_X2 U7635 ( .A(n11341), .ZN(n8053) );
  INV_X1 U7636 ( .A(n8948), .ZN(n9085) );
  INV_X1 U7637 ( .A(n13691), .ZN(n11389) );
  CLKBUF_X2 U7638 ( .A(n13677), .Z(n13870) );
  NAND2_X2 U7639 ( .A1(n13669), .A2(n11702), .ZN(n10767) );
  INV_X1 U7640 ( .A(n13695), .ZN(n11422) );
  INV_X1 U7641 ( .A(n14626), .ZN(n11367) );
  INV_X1 U7642 ( .A(n11727), .ZN(n7933) );
  INV_X1 U7643 ( .A(n13667), .ZN(n11702) );
  NAND2_X2 U7644 ( .A1(n10535), .A2(n10878), .ZN(n13594) );
  INV_X4 U7645 ( .A(n9587), .ZN(n9904) );
  INV_X1 U7646 ( .A(n8772), .ZN(n8814) );
  INV_X1 U7647 ( .A(n13902), .ZN(n7420) );
  NOR2_X1 U7648 ( .A1(n10504), .A2(n15600), .ZN(n9114) );
  NAND2_X2 U7649 ( .A1(n9715), .A2(n13248), .ZN(n10131) );
  INV_X2 U7650 ( .A(n10420), .ZN(n10431) );
  INV_X8 U7651 ( .A(n10420), .ZN(n10432) );
  NAND3_X1 U7652 ( .A1(n8188), .A2(n8603), .A3(n8187), .ZN(n8508) );
  AND2_X1 U7653 ( .A1(n8189), .A2(n8506), .ZN(n8378) );
  INV_X1 U7654 ( .A(n10720), .ZN(n10093) );
  INV_X1 U7655 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n10086) );
  INV_X1 U7656 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n10087) );
  INV_X2 U7657 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n7685) );
  AND2_X1 U7658 ( .A1(n7605), .A2(n7604), .ZN(n14957) );
  OR2_X1 U7659 ( .A1(n9745), .A2(n14163), .ZN(n8337) );
  OAI22_X1 U7660 ( .A1(n13860), .A2(n13859), .B1(n13875), .B2(n13874), .ZN(
        n13873) );
  AOI21_X1 U7661 ( .B1(n16330), .B2(n15286), .A(n15285), .ZN(n15490) );
  NAND2_X1 U7662 ( .A1(n13547), .A2(n13546), .ZN(n14750) );
  AND2_X1 U7663 ( .A1(n7587), .A2(n7586), .ZN(n14967) );
  NOR2_X1 U7664 ( .A1(n14757), .A2(n14758), .ZN(n7604) );
  AND2_X1 U7665 ( .A1(n7792), .A2(n7643), .ZN(n7642) );
  OR2_X1 U7666 ( .A1(n14219), .A2(n14218), .ZN(n14366) );
  OR2_X1 U7667 ( .A1(n15478), .A2(n16299), .ZN(n7643) );
  AOI211_X1 U7668 ( .C1(n14944), .C2(n7467), .A(n10363), .B(n14729), .ZN(
        n14943) );
  AND2_X1 U7669 ( .A1(n13345), .A2(n15258), .ZN(n15476) );
  AOI21_X1 U7670 ( .B1(n7702), .B2(n7700), .A(n7699), .ZN(n7698) );
  AND2_X1 U7671 ( .A1(n8184), .A2(n15076), .ZN(n8183) );
  XNOR2_X1 U7672 ( .A(n15943), .B(n7923), .ZN(n15942) );
  AND2_X1 U7673 ( .A1(n13620), .A2(n13619), .ZN(n14942) );
  AND2_X1 U7674 ( .A1(n8911), .A2(n8910), .ZN(n15474) );
  NAND2_X1 U7675 ( .A1(n13306), .A2(n13305), .ZN(n15147) );
  NAND2_X1 U7676 ( .A1(n14278), .A2(n9606), .ZN(n14264) );
  AOI21_X1 U7677 ( .B1(n8344), .B2(n9936), .A(n7449), .ZN(n8343) );
  NOR2_X1 U7678 ( .A1(n8345), .A2(n14204), .ZN(n8344) );
  XOR2_X1 U7679 ( .A(n13591), .B(n13590), .Z(n15076) );
  AND2_X1 U7680 ( .A1(n9739), .A2(n9940), .ZN(n14221) );
  AND2_X1 U7681 ( .A1(n15422), .A2(n13360), .ZN(n15403) );
  OR2_X1 U7682 ( .A1(n14227), .A2(n14208), .ZN(n9739) );
  NAND2_X1 U7683 ( .A1(n9647), .A2(n9646), .ZN(n14227) );
  NAND2_X1 U7684 ( .A1(n7904), .A2(n7903), .ZN(n14096) );
  NAND2_X1 U7685 ( .A1(n8562), .A2(n8561), .ZN(n15498) );
  NAND2_X1 U7686 ( .A1(n16319), .A2(n16320), .ZN(n16318) );
  OR2_X1 U7687 ( .A1(n14086), .A2(n10237), .ZN(n7904) );
  OAI21_X1 U7688 ( .B1(n9645), .B2(n13463), .A(n9189), .ZN(n9659) );
  OR2_X1 U7689 ( .A1(n9021), .A2(n7891), .ZN(n7888) );
  NAND2_X1 U7690 ( .A1(n13178), .A2(n9733), .ZN(n13175) );
  XNOR2_X1 U7691 ( .A(n14975), .B(n14837), .ZN(n14818) );
  NAND2_X1 U7692 ( .A1(n8895), .A2(n8894), .ZN(n15349) );
  OR2_X1 U7693 ( .A1(n12142), .A2(n12141), .ZN(n7981) );
  NAND2_X1 U7694 ( .A1(n12321), .A2(n12325), .ZN(n12320) );
  XOR2_X1 U7695 ( .A(n14496), .B(n14495), .Z(n14541) );
  NAND2_X1 U7696 ( .A1(n13420), .A2(n13419), .ZN(n14993) );
  NAND2_X2 U7697 ( .A1(n13408), .A2(n13407), .ZN(n15001) );
  OR2_X1 U7698 ( .A1(n9002), .A2(n9003), .ZN(n7882) );
  NAND2_X1 U7699 ( .A1(n8849), .A2(n8848), .ZN(n15534) );
  NAND2_X1 U7700 ( .A1(n8060), .A2(n16354), .ZN(n15451) );
  NAND2_X2 U7701 ( .A1(n13400), .A2(n13399), .ZN(n15005) );
  NAND2_X1 U7702 ( .A1(n7921), .A2(n15871), .ZN(n15878) );
  NAND2_X1 U7703 ( .A1(n8866), .A2(n8865), .ZN(n15542) );
  INV_X1 U7704 ( .A(n14346), .ZN(n14174) );
  NAND2_X1 U7705 ( .A1(n12536), .A2(n12535), .ZN(n15011) );
  NAND2_X1 U7706 ( .A1(n8607), .A2(n8606), .ZN(n15550) );
  NAND2_X1 U7707 ( .A1(n7573), .A2(n7465), .ZN(n7986) );
  NAND2_X1 U7708 ( .A1(n8633), .A2(n8632), .ZN(n13354) );
  NAND2_X1 U7709 ( .A1(n14644), .A2(n11602), .ZN(n11603) );
  NAND2_X1 U7710 ( .A1(n12213), .A2(n12212), .ZN(n13774) );
  OR2_X1 U7711 ( .A1(n14164), .A2(n9701), .ZN(n14172) );
  XNOR2_X1 U7712 ( .A(n10151), .B(n16019), .ZN(n16012) );
  NAND2_X2 U7713 ( .A1(n9656), .A2(n9655), .ZN(n14360) );
  AND2_X1 U7714 ( .A1(n11382), .A2(n10150), .ZN(n10151) );
  XNOR2_X1 U7715 ( .A(n15847), .B(n7929), .ZN(n15846) );
  NAND2_X1 U7716 ( .A1(n7930), .A2(n15839), .ZN(n15847) );
  NAND2_X1 U7717 ( .A1(n11862), .A2(n11861), .ZN(n13747) );
  NAND2_X1 U7718 ( .A1(n12103), .A2(n12102), .ZN(n13758) );
  NAND2_X1 U7719 ( .A1(n12185), .A2(n12184), .ZN(n13770) );
  NAND2_X1 U7720 ( .A1(n7978), .A2(n7977), .ZN(n11375) );
  NAND2_X1 U7721 ( .A1(n11857), .A2(n11856), .ZN(n13734) );
  NOR2_X1 U7722 ( .A1(n11781), .A2(n8046), .ZN(n8048) );
  AND2_X1 U7723 ( .A1(n7658), .A2(n7536), .ZN(n10952) );
  INV_X2 U7724 ( .A(n14843), .ZN(n14938) );
  INV_X2 U7725 ( .A(n16100), .ZN(n14341) );
  NOR2_X1 U7726 ( .A1(n15993), .A2(n9381), .ZN(n15992) );
  OR2_X1 U7727 ( .A1(n10674), .A2(n10673), .ZN(n7658) );
  INV_X2 U7728 ( .A(n16315), .ZN(n7419) );
  NAND2_X1 U7729 ( .A1(n8143), .A2(n11039), .ZN(n11203) );
  NOR2_X1 U7730 ( .A1(n10668), .A2(n10667), .ZN(n10674) );
  AND2_X1 U7731 ( .A1(n14562), .A2(n14563), .ZN(n14630) );
  AND2_X1 U7732 ( .A1(n9601), .A2(n12802), .ZN(n9611) );
  NAND2_X1 U7733 ( .A1(n8426), .A2(n8425), .ZN(n8427) );
  AND2_X1 U7734 ( .A1(n7709), .A2(n7708), .ZN(n10684) );
  NAND2_X1 U7735 ( .A1(n11134), .A2(n11133), .ZN(n13706) );
  NAND2_X1 U7736 ( .A1(n7873), .A2(n9768), .ZN(n9801) );
  INV_X1 U7737 ( .A(n16040), .ZN(n7579) );
  AND2_X1 U7738 ( .A1(n9958), .A2(n9953), .ZN(n10396) );
  INV_X1 U7739 ( .A(n13716), .ZN(n13676) );
  MUX2_X1 U7740 ( .A(n13258), .B(n10578), .S(n10577), .Z(n10580) );
  INV_X2 U7741 ( .A(n13677), .ZN(n13716) );
  INV_X1 U7742 ( .A(n14690), .ZN(n7422) );
  AND2_X1 U7743 ( .A1(n11890), .A2(n15711), .ZN(n10938) );
  AND2_X1 U7744 ( .A1(n7843), .A2(n7845), .ZN(n7842) );
  OAI211_X1 U7745 ( .C1(n10312), .C2(n10429), .A(n10325), .B(n10324), .ZN(
        n13695) );
  INV_X4 U7746 ( .A(n10669), .ZN(n13265) );
  NAND4_X1 U7747 ( .A1(n9297), .A2(n9296), .A3(n9295), .A4(n9294), .ZN(n14059)
         );
  AOI21_X1 U7748 ( .B1(n7610), .B2(n7609), .A(n15815), .ZN(n15823) );
  INV_X1 U7749 ( .A(n13680), .ZN(n7431) );
  AOI21_X1 U7750 ( .B1(n8269), .B2(n8267), .A(n8266), .ZN(n8265) );
  NOR2_X1 U7751 ( .A1(n10663), .A2(n8074), .ZN(n11890) );
  NAND4_X2 U7752 ( .A1(n9315), .A2(n9314), .A3(n9313), .A4(n9312), .ZN(n14057)
         );
  INV_X1 U7753 ( .A(n10876), .ZN(n11236) );
  AND2_X1 U7755 ( .A1(n8270), .A2(n8366), .ZN(n8269) );
  OR2_X1 U7756 ( .A1(n11151), .A2(n10176), .ZN(n11153) );
  NOR2_X1 U7757 ( .A1(n8249), .A2(n8248), .ZN(n7843) );
  CLKBUF_X3 U7758 ( .A(n8814), .Z(n7428) );
  CLKBUF_X1 U7759 ( .A(n12412), .Z(n13615) );
  CLKBUF_X3 U7760 ( .A(n9904), .Z(n9717) );
  INV_X2 U7761 ( .A(n8773), .ZN(n8758) );
  AND2_X1 U7762 ( .A1(n7726), .A2(n7725), .ZN(n10816) );
  OR2_X1 U7763 ( .A1(n9499), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9518) );
  BUF_X2 U7764 ( .A(n12110), .Z(n13522) );
  XNOR2_X1 U7765 ( .A(n15813), .B(n10860), .ZN(n15814) );
  INV_X1 U7766 ( .A(n10271), .ZN(n13329) );
  INV_X2 U7767 ( .A(n10455), .ZN(n8864) );
  NAND2_X1 U7768 ( .A1(n9254), .A2(n9253), .ZN(n11767) );
  INV_X1 U7769 ( .A(n13912), .ZN(n8074) );
  NOR2_X1 U7770 ( .A1(n8248), .A2(n7846), .ZN(n7844) );
  NAND2_X4 U7771 ( .A1(n15594), .A2(n13245), .ZN(n10455) );
  AND2_X1 U7772 ( .A1(n8247), .A2(n12974), .ZN(n7840) );
  NAND2_X4 U7773 ( .A1(n15064), .A2(n10370), .ZN(n11131) );
  INV_X1 U7774 ( .A(n8381), .ZN(n8540) );
  XNOR2_X1 U7775 ( .A(n9113), .B(P1_IR_REG_25__SCAN_IN), .ZN(n15602) );
  XNOR2_X1 U7776 ( .A(n10289), .B(P2_IR_REG_21__SCAN_IN), .ZN(n13662) );
  XNOR2_X1 U7777 ( .A(n9111), .B(n9110), .ZN(n15600) );
  XNOR2_X1 U7778 ( .A(n8429), .B(SI_10_), .ZN(n8246) );
  INV_X1 U7779 ( .A(n8704), .ZN(n8247) );
  INV_X2 U7780 ( .A(n15059), .ZN(n13255) );
  XNOR2_X1 U7781 ( .A(n9215), .B(n9211), .ZN(n9715) );
  NAND2_X1 U7782 ( .A1(n9112), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9113) );
  NAND2_X1 U7783 ( .A1(n10285), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10289) );
  XNOR2_X1 U7784 ( .A(n9259), .B(n9207), .ZN(n14145) );
  XNOR2_X1 U7785 ( .A(n8402), .B(n12761), .ZN(n8747) );
  NAND2_X2 U7786 ( .A1(n10432), .A2(P3_U3151), .ZN(n13926) );
  XNOR2_X1 U7787 ( .A(n8498), .B(n8497), .ZN(n13245) );
  NAND2_X1 U7788 ( .A1(n8499), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8501) );
  NAND2_X1 U7789 ( .A1(n9214), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9215) );
  NAND2_X1 U7790 ( .A1(n8517), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8518) );
  NAND2_X1 U7791 ( .A1(n8504), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8505) );
  NAND2_X1 U7792 ( .A1(n8079), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10291) );
  NAND2_X2 U7793 ( .A1(n10420), .A2(P1_U3086), .ZN(n15604) );
  INV_X1 U7794 ( .A(n8079), .ZN(n10286) );
  INV_X2 U7795 ( .A(n8767), .ZN(n10420) );
  INV_X1 U7796 ( .A(n8508), .ZN(n8225) );
  OR2_X1 U7797 ( .A1(n8510), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n8504) );
  AND2_X2 U7798 ( .A1(n8353), .A2(n8352), .ZN(n9208) );
  NAND2_X1 U7799 ( .A1(n8077), .A2(n7486), .ZN(n8079) );
  OAI211_X1 U7800 ( .C1(n9287), .C2(n7910), .A(n9288), .B(n7909), .ZN(n10475)
         );
  NAND4_X1 U7801 ( .A1(n7793), .A2(n10094), .A3(n10093), .A4(n10410), .ZN(
        n11769) );
  NAND2_X2 U7802 ( .A1(n7638), .A2(n7636), .ZN(n8767) );
  AND2_X1 U7803 ( .A1(n8355), .A2(n9207), .ZN(n8354) );
  AND4_X1 U7804 ( .A1(n10267), .A2(n10266), .A3(n10265), .A4(n10264), .ZN(
        n8365) );
  AND2_X2 U7805 ( .A1(n8372), .A2(n8190), .ZN(n8188) );
  NAND2_X1 U7806 ( .A1(n7608), .A2(n7607), .ZN(n7577) );
  AND2_X1 U7807 ( .A1(n8362), .A2(n9206), .ZN(n8352) );
  NOR2_X1 U7808 ( .A1(n10280), .A2(n10279), .ZN(n10281) );
  INV_X1 U7809 ( .A(n10719), .ZN(n10094) );
  AND2_X2 U7810 ( .A1(n8645), .A2(n8191), .ZN(n8187) );
  NAND3_X1 U7811 ( .A1(n7685), .A2(n7684), .A3(n7683), .ZN(n8116) );
  AND4_X1 U7812 ( .A1(n9205), .A2(n9204), .A3(n9203), .A4(n9202), .ZN(n8362)
         );
  NAND4_X1 U7813 ( .A1(n11221), .A2(n10088), .A3(n10087), .A4(n10086), .ZN(
        n11770) );
  INV_X1 U7814 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9100) );
  INV_X1 U7815 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n8862) );
  NOR2_X1 U7816 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n8191) );
  NOR2_X2 U7817 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n8774) );
  NOR2_X1 U7818 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n8370) );
  NOR2_X1 U7819 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n8371) );
  INV_X1 U7820 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n13154) );
  NOR2_X1 U7821 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n8377) );
  NOR2_X2 U7822 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n8645) );
  INV_X1 U7823 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n10263) );
  INV_X1 U7824 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n10261) );
  INV_X1 U7825 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8078) );
  NOR2_X1 U7826 ( .A1(P3_IR_REG_11__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n9202) );
  NOR2_X1 U7827 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_16__SCAN_IN), .ZN(
        n9203) );
  NOR2_X1 U7828 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_13__SCAN_IN), .ZN(
        n9204) );
  INV_X1 U7829 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9247) );
  INV_X1 U7830 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n9217) );
  INV_X1 U7831 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n10409) );
  INV_X1 U7832 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7683) );
  INV_X1 U7833 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7684) );
  INV_X1 U7834 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n9349) );
  NAND2_X4 U7835 ( .A1(n9278), .A2(n9276), .ZN(n9293) );
  NAND2_X1 U7836 ( .A1(n8487), .A2(n8486), .ZN(n8918) );
  NOR2_X2 U7837 ( .A1(n12430), .A2(n15025), .ZN(n7974) );
  INV_X1 U7838 ( .A(n8952), .ZN(n7421) );
  INV_X1 U7839 ( .A(n8952), .ZN(n8958) );
  NOR2_X2 U7840 ( .A1(n15833), .A2(n15956), .ZN(n15836) );
  NOR2_X2 U7841 ( .A1(n9687), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9700) );
  CLKBUF_X1 U7842 ( .A(n14690), .Z(n7423) );
  NAND4_X1 U7843 ( .A1(n10276), .A2(n10273), .A3(n10274), .A4(n10275), .ZN(
        n14690) );
  OR2_X2 U7844 ( .A1(n9093), .A2(n9094), .ZN(n7477) );
  AOI21_X2 U7845 ( .B1(n12533), .B2(n13643), .A(n12532), .ZN(n13403) );
  AOI21_X2 U7846 ( .B1(n12506), .B2(n13642), .A(n12505), .ZN(n12533) );
  NAND2_X2 U7847 ( .A1(n12420), .A2(n12419), .ZN(n12506) );
  INV_X1 U7848 ( .A(n9587), .ZN(n7424) );
  NAND2_X1 U7849 ( .A1(n9278), .A2(n13927), .ZN(n9587) );
  AOI22_X2 U7850 ( .A1(n14611), .A2(n14610), .B1(n14500), .B2(n14499), .ZN(
        n14569) );
  AND2_X2 U7851 ( .A1(n8602), .A2(n13154), .ZN(n8190) );
  NAND2_X2 U7852 ( .A1(n10535), .A2(n10532), .ZN(n10669) );
  OAI22_X2 U7853 ( .A1(n14193), .A2(n14199), .B1(n14351), .B2(n14356), .ZN(
        n14182) );
  XNOR2_X2 U7854 ( .A(n15883), .B(n15882), .ZN(n15884) );
  AND2_X2 U7855 ( .A1(n7611), .A2(n7585), .ZN(n15883) );
  AND3_X2 U7856 ( .A1(n13158), .A2(n8862), .A3(n12930), .ZN(n8372) );
  INV_X2 U7857 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n12930) );
  NAND2_X1 U7858 ( .A1(n10455), .A2(n10432), .ZN(n7426) );
  NOR2_X2 U7859 ( .A1(n9518), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9534) );
  XNOR2_X1 U7860 ( .A(n15194), .B(n11260), .ZN(n11104) );
  OAI21_X2 U7861 ( .B1(n8964), .B2(n11006), .A(n8963), .ZN(n8966) );
  NOR2_X2 U7863 ( .A1(n11892), .A2(n13747), .ZN(n12040) );
  CLKBUF_X1 U7864 ( .A(n8847), .Z(n7429) );
  OAI211_X1 U7865 ( .C1(n10455), .C2(n10972), .A(n8749), .B(n8748), .ZN(n11260) );
  AND2_X1 U7866 ( .A1(n15923), .A2(n15924), .ZN(n15928) );
  BUF_X4 U7867 ( .A(n10328), .Z(n13517) );
  NAND2_X1 U7868 ( .A1(n10455), .A2(n10432), .ZN(n8773) );
  AOI21_X2 U7869 ( .B1(n15897), .B2(n15896), .A(n15895), .ZN(n15910) );
  NOR2_X2 U7870 ( .A1(n14824), .A2(n14969), .ZN(n14802) );
  NOR2_X2 U7871 ( .A1(n11209), .A2(n13695), .ZN(n11211) );
  OR2_X1 U7872 ( .A1(n10773), .A2(n14626), .ZN(n11209) );
  NAND2_X1 U7874 ( .A1(n9856), .A2(n14197), .ZN(n7862) );
  AND2_X1 U7875 ( .A1(n10112), .A2(n10187), .ZN(n7993) );
  NOR2_X1 U7876 ( .A1(n8165), .A2(n13540), .ZN(n8164) );
  INV_X1 U7877 ( .A(n13539), .ZN(n8165) );
  AND2_X1 U7878 ( .A1(n8374), .A2(n8375), .ZN(n8506) );
  AOI21_X1 U7879 ( .B1(n14006), .B2(n14244), .A(n9848), .ZN(n13943) );
  INV_X1 U7880 ( .A(n9293), .ZN(n9718) );
  INV_X1 U7882 ( .A(n11742), .ZN(n8092) );
  AND2_X1 U7883 ( .A1(n8152), .A2(n12551), .ZN(n8149) );
  AND2_X1 U7884 ( .A1(n10539), .A2(n10371), .ZN(n14883) );
  NAND2_X1 U7885 ( .A1(n10539), .A2(n10370), .ZN(n14916) );
  NOR2_X1 U7886 ( .A1(n11924), .A2(n7787), .ZN(n7785) );
  NOR2_X1 U7887 ( .A1(n9019), .A2(n9016), .ZN(n8242) );
  INV_X1 U7888 ( .A(n9016), .ZN(n8241) );
  INV_X1 U7889 ( .A(n13819), .ZN(n7814) );
  OAI21_X1 U7890 ( .B1(n13813), .B2(n13812), .A(n7509), .ZN(n7813) );
  NAND2_X1 U7891 ( .A1(n8416), .A2(n8827), .ZN(n8414) );
  OR2_X1 U7892 ( .A1(n14356), .A2(n14186), .ZN(n9929) );
  OR2_X1 U7893 ( .A1(n14372), .A2(n14252), .ZN(n10039) );
  OR2_X1 U7894 ( .A1(n14389), .A2(n14268), .ZN(n10027) );
  NOR2_X1 U7895 ( .A1(n9470), .A2(n7947), .ZN(n7946) );
  INV_X1 U7896 ( .A(n9799), .ZN(n7947) );
  INV_X1 U7897 ( .A(n9278), .ZN(n9277) );
  OR2_X1 U7898 ( .A1(n9230), .A2(P3_D_REG_0__SCAN_IN), .ZN(n9229) );
  NAND2_X1 U7899 ( .A1(n12580), .A2(n12581), .ZN(n8115) );
  NAND2_X1 U7900 ( .A1(n7415), .A2(n13666), .ZN(n8071) );
  INV_X1 U7901 ( .A(n13475), .ZN(n7830) );
  INV_X1 U7902 ( .A(n7663), .ZN(n7662) );
  AOI21_X1 U7903 ( .B1(n7665), .B2(n7458), .A(n7664), .ZN(n7663) );
  INV_X1 U7904 ( .A(n15106), .ZN(n7664) );
  OR2_X1 U7905 ( .A1(n12486), .A2(n8369), .ZN(n8021) );
  XNOR2_X1 U7906 ( .A(n11074), .B(n10876), .ZN(n8003) );
  NAND2_X1 U7907 ( .A1(n12701), .A2(n12700), .ZN(n12703) );
  INV_X1 U7908 ( .A(n8269), .ZN(n8268) );
  INV_X1 U7909 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7928) );
  NAND2_X1 U7910 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n7607) );
  AND2_X1 U7911 ( .A1(n7856), .A2(n8127), .ZN(n7855) );
  NAND2_X1 U7912 ( .A1(n12257), .A2(n7483), .ZN(n12398) );
  INV_X1 U7913 ( .A(n9792), .ZN(n8129) );
  XNOR2_X1 U7914 ( .A(n9849), .B(n16049), .ZN(n9773) );
  NAND2_X1 U7915 ( .A1(n7872), .A2(n9783), .ZN(n11943) );
  OAI21_X1 U7916 ( .B1(n11413), .B2(n8132), .A(n8130), .ZN(n7872) );
  NAND2_X1 U7917 ( .A1(n7858), .A2(n7862), .ZN(n7857) );
  INV_X1 U7918 ( .A(n13967), .ZN(n7858) );
  NAND2_X1 U7919 ( .A1(n10475), .A2(n10136), .ZN(n7908) );
  NAND2_X1 U7920 ( .A1(n10111), .A2(n10850), .ZN(n10854) );
  NOR2_X1 U7921 ( .A1(n15996), .A2(n9378), .ZN(n15995) );
  NAND2_X1 U7922 ( .A1(n7912), .A2(n7911), .ZN(n11382) );
  INV_X1 U7923 ( .A(n11379), .ZN(n7911) );
  NOR2_X1 U7924 ( .A1(n16012), .A2(n9405), .ZN(n16011) );
  NOR2_X1 U7925 ( .A1(n14077), .A2(n10228), .ZN(n10232) );
  INV_X1 U7926 ( .A(n10238), .ZN(n7903) );
  AOI21_X1 U7927 ( .B1(n7649), .B2(n7951), .A(n7648), .ZN(n14220) );
  INV_X1 U7928 ( .A(n7949), .ZN(n7648) );
  AOI21_X1 U7929 ( .B1(n7951), .B2(n7950), .A(n7517), .ZN(n7949) );
  NAND2_X1 U7930 ( .A1(n9738), .A2(n7704), .ZN(n14235) );
  OR2_X1 U7931 ( .A1(n14385), .A2(n14281), .ZN(n10030) );
  NAND2_X1 U7932 ( .A1(n14270), .A2(n10031), .ZN(n8349) );
  NAND2_X1 U7933 ( .A1(n12286), .A2(n8348), .ZN(n12328) );
  NOR2_X1 U7934 ( .A1(n12325), .A2(n9978), .ZN(n8348) );
  INV_X1 U7935 ( .A(n9917), .ZN(n9686) );
  INV_X1 U7936 ( .A(n9562), .ZN(n9916) );
  INV_X1 U7937 ( .A(n7594), .ZN(n9581) );
  INV_X1 U7939 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n9206) );
  NOR2_X1 U7940 ( .A1(n7761), .A2(n7764), .ZN(n7760) );
  NOR2_X1 U7941 ( .A1(n9255), .A2(n9210), .ZN(n9219) );
  AOI21_X1 U7942 ( .B1(n7768), .B2(n7769), .A(n7767), .ZN(n7766) );
  INV_X1 U7943 ( .A(n9149), .ZN(n7767) );
  INV_X1 U7944 ( .A(n9145), .ZN(n7772) );
  AND2_X1 U7945 ( .A1(n9335), .A2(n9141), .ZN(n9353) );
  NAND2_X1 U7946 ( .A1(n7747), .A2(n7448), .ZN(n7746) );
  AND2_X1 U7947 ( .A1(n8091), .A2(n11741), .ZN(n8090) );
  AOI21_X1 U7948 ( .B1(n7592), .B2(n7591), .A(n13880), .ZN(n7590) );
  INV_X1 U7949 ( .A(n13858), .ZN(n7591) );
  AOI21_X1 U7950 ( .B1(n8148), .B2(n8146), .A(n7501), .ZN(n8145) );
  INV_X1 U7951 ( .A(n8148), .ZN(n8147) );
  AND2_X1 U7952 ( .A1(n14770), .A2(n13487), .ZN(n14794) );
  NAND2_X1 U7953 ( .A1(n14873), .A2(n8164), .ZN(n8162) );
  NOR2_X1 U7954 ( .A1(n13643), .A2(n8151), .ZN(n8150) );
  INV_X1 U7955 ( .A(n12521), .ZN(n8151) );
  NAND2_X1 U7956 ( .A1(n10660), .A2(n13861), .ZN(n14924) );
  INV_X1 U7957 ( .A(n10661), .ZN(n14902) );
  INV_X1 U7958 ( .A(n13871), .ZN(n14944) );
  NOR2_X1 U7959 ( .A1(n14734), .A2(n14737), .ZN(n7583) );
  INV_X1 U7960 ( .A(n13240), .ZN(n10352) );
  NAND2_X1 U7961 ( .A1(n8037), .A2(n8041), .ZN(n10292) );
  INV_X1 U7962 ( .A(n8042), .ZN(n8041) );
  OAI21_X1 U7963 ( .B1(n15076), .B2(n7680), .A(n7679), .ZN(n7678) );
  NOR2_X1 U7964 ( .A1(n15166), .A2(n8185), .ZN(n7680) );
  NAND2_X1 U7965 ( .A1(n15076), .A2(n13586), .ZN(n7679) );
  AND2_X1 U7966 ( .A1(n13557), .A2(n13554), .ZN(n8209) );
  OR2_X1 U7967 ( .A1(n15166), .A2(n8185), .ZN(n8184) );
  NAND2_X1 U7968 ( .A1(n10455), .A2(n10420), .ZN(n8772) );
  NAND2_X2 U7969 ( .A1(n9114), .A2(n15602), .ZN(n10535) );
  INV_X1 U7970 ( .A(n15282), .ZN(n15079) );
  NAND2_X1 U7971 ( .A1(n7619), .A2(n15474), .ZN(n15258) );
  NAND2_X1 U7972 ( .A1(n11489), .A2(n11485), .ZN(n8287) );
  AND2_X1 U7973 ( .A1(n11485), .A2(n11298), .ZN(n8285) );
  INV_X1 U7974 ( .A(n8506), .ZN(n8507) );
  OAI21_X1 U7975 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(n15868), .A(n15867), .ZN(
        n15874) );
  NAND2_X1 U7976 ( .A1(n12049), .A2(n12048), .ZN(n12047) );
  CLKBUF_X1 U7977 ( .A(n13943), .Z(n13989) );
  INV_X1 U7978 ( .A(n14186), .ZN(n14351) );
  OR2_X2 U7979 ( .A1(n10232), .A2(n10231), .ZN(n14107) );
  AND2_X1 U7980 ( .A1(n9628), .A2(n9627), .ZN(n14244) );
  NAND2_X1 U7981 ( .A1(n13435), .A2(n13434), .ZN(n14987) );
  INV_X1 U7982 ( .A(n14929), .ZN(n14840) );
  OAI21_X1 U7983 ( .B1(n15869), .B2(n15870), .A(P2_ADDR_REG_10__SCAN_IN), .ZN(
        n7921) );
  AOI22_X1 U7984 ( .A1(n13671), .A2(n13670), .B1(n13669), .B2(n13668), .ZN(
        n13672) );
  NAND2_X1 U7985 ( .A1(n13707), .A2(n13708), .ZN(n7795) );
  NAND2_X1 U7986 ( .A1(n7799), .A2(n7798), .ZN(n7797) );
  INV_X1 U7987 ( .A(n13708), .ZN(n7798) );
  INV_X1 U7988 ( .A(n7795), .ZN(n7794) );
  AND2_X1 U7989 ( .A1(n9003), .A2(n8220), .ZN(n8219) );
  OAI21_X1 U7990 ( .B1(n13750), .B2(n13749), .A(n7512), .ZN(n7808) );
  NAND2_X1 U7991 ( .A1(n7462), .A2(n7812), .ZN(n7811) );
  OR2_X1 U7992 ( .A1(n7554), .A2(n9029), .ZN(n7613) );
  AOI21_X1 U7993 ( .B1(n7886), .B2(n7891), .A(n7884), .ZN(n7883) );
  INV_X1 U7994 ( .A(n9045), .ZN(n7895) );
  NAND2_X1 U7995 ( .A1(n13788), .A2(n7479), .ZN(n8335) );
  NOR2_X1 U7996 ( .A1(n13788), .A2(n7479), .ZN(n8336) );
  NAND2_X1 U7997 ( .A1(n9047), .A2(n9045), .ZN(n7894) );
  NAND2_X1 U7998 ( .A1(n9062), .A2(n9064), .ZN(n7876) );
  INV_X1 U7999 ( .A(n13837), .ZN(n7806) );
  OAI211_X1 U8000 ( .C1(n9941), .C2(n8308), .A(n8305), .B(n8304), .ZN(n8303)
         );
  NAND2_X1 U8001 ( .A1(n8309), .A2(n10043), .ZN(n8308) );
  AND2_X1 U8002 ( .A1(n8307), .A2(n8306), .ZN(n8305) );
  NAND2_X1 U8003 ( .A1(n9938), .A2(n10129), .ZN(n8304) );
  NAND2_X1 U8004 ( .A1(n8329), .A2(n8326), .ZN(n8325) );
  NOR2_X1 U8005 ( .A1(n7806), .A2(n7482), .ZN(n7805) );
  AND2_X1 U8006 ( .A1(n13834), .A2(n8311), .ZN(n8310) );
  NAND2_X1 U8007 ( .A1(n7806), .A2(n7482), .ZN(n7804) );
  NAND2_X1 U8008 ( .A1(n8328), .A2(n8327), .ZN(n8326) );
  INV_X1 U8009 ( .A(n13841), .ZN(n8327) );
  INV_X1 U8010 ( .A(n13842), .ZN(n8328) );
  NAND2_X1 U8011 ( .A1(n7805), .A2(n7804), .ZN(n7801) );
  AND2_X1 U8012 ( .A1(n13841), .A2(n13842), .ZN(n8329) );
  NAND2_X1 U8013 ( .A1(n7833), .A2(n8454), .ZN(n8455) );
  NAND2_X1 U8014 ( .A1(n7832), .A2(n7494), .ZN(n7833) );
  INV_X1 U8015 ( .A(n8600), .ZN(n7831) );
  INV_X1 U8016 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n8602) );
  INV_X1 U8017 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n15788) );
  OAI21_X1 U8018 ( .B1(P3_ADDR_REG_15__SCAN_IN), .B2(n15922), .A(n15921), .ZN(
        n15929) );
  AND2_X1 U8019 ( .A1(n8126), .A2(n7537), .ZN(n8125) );
  NAND2_X1 U8020 ( .A1(n13928), .A2(n8128), .ZN(n8126) );
  NAND2_X1 U8021 ( .A1(n10144), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7920) );
  AND2_X1 U8022 ( .A1(n11623), .A2(n10153), .ZN(n10154) );
  NAND2_X1 U8023 ( .A1(n7981), .A2(n7980), .ZN(n7979) );
  INV_X1 U8024 ( .A(n10208), .ZN(n7980) );
  NAND2_X1 U8025 ( .A1(n7695), .A2(n7697), .ZN(n7693) );
  INV_X1 U8026 ( .A(n7696), .ZN(n7695) );
  OAI21_X1 U8027 ( .B1(n9576), .B2(n7697), .A(n14293), .ZN(n7696) );
  INV_X1 U8028 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n13158) );
  NAND2_X1 U8029 ( .A1(n9633), .A2(n9187), .ZN(n9188) );
  INV_X1 U8030 ( .A(n7756), .ZN(n7755) );
  OAI21_X1 U8031 ( .B1(n7758), .B2(n7757), .A(n9607), .ZN(n7756) );
  INV_X1 U8032 ( .A(n9179), .ZN(n7757) );
  NAND2_X1 U8033 ( .A1(n8140), .A2(n8138), .ZN(n9250) );
  AND2_X1 U8034 ( .A1(n9216), .A2(n9256), .ZN(n8141) );
  INV_X1 U8035 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n9216) );
  INV_X1 U8036 ( .A(n9255), .ZN(n8140) );
  NOR2_X1 U8037 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .ZN(
        n9199) );
  NAND2_X1 U8038 ( .A1(n9458), .A2(n9161), .ZN(n9162) );
  CLKBUF_X1 U8039 ( .A(n9329), .Z(n9350) );
  XNOR2_X1 U8040 ( .A(n11125), .B(n14626), .ZN(n10321) );
  NAND2_X1 U8041 ( .A1(n13912), .A2(n13662), .ZN(n13666) );
  NOR2_X1 U8042 ( .A1(n14954), .A2(n14959), .ZN(n7969) );
  NAND2_X1 U8043 ( .A1(n7827), .A2(n13475), .ZN(n7826) );
  NAND2_X1 U8044 ( .A1(n7826), .A2(n14794), .ZN(n7824) );
  AOI21_X1 U8045 ( .B1(n14818), .B2(n13542), .A(n14810), .ZN(n8148) );
  NOR2_X1 U8046 ( .A1(n13637), .A2(n8034), .ZN(n8033) );
  INV_X1 U8047 ( .A(n12026), .ZN(n8034) );
  OR2_X1 U8048 ( .A1(n11536), .A2(n11535), .ZN(n8049) );
  NAND2_X1 U8049 ( .A1(n7420), .A2(n8074), .ZN(n8073) );
  INV_X1 U8050 ( .A(n7972), .ZN(n14864) );
  NOR2_X2 U8051 ( .A1(n11770), .A2(n10090), .ZN(n7793) );
  INV_X1 U8052 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n10089) );
  OR2_X1 U8053 ( .A1(n11291), .A2(P2_IR_REG_15__SCAN_IN), .ZN(n11733) );
  INV_X1 U8054 ( .A(n11274), .ZN(n8199) );
  NOR2_X1 U8055 ( .A1(n11337), .A2(n8201), .ZN(n8200) );
  INV_X1 U8056 ( .A(n8256), .ZN(n8252) );
  OR2_X1 U8057 ( .A1(n15498), .A2(n15334), .ZN(n8058) );
  INV_X1 U8058 ( .A(n12702), .ZN(n8014) );
  INV_X1 U8059 ( .A(n13355), .ZN(n8016) );
  NOR2_X2 U8060 ( .A1(n12695), .A2(n13354), .ZN(n8060) );
  OR2_X1 U8061 ( .A1(n11920), .A2(n8274), .ZN(n8273) );
  INV_X1 U8062 ( .A(n15188), .ZN(n11931) );
  INV_X1 U8063 ( .A(n11642), .ZN(n8006) );
  NAND2_X1 U8064 ( .A1(n15450), .A2(n15461), .ZN(n8284) );
  OAI21_X1 U8065 ( .B1(n8918), .B2(n8917), .A(n8491), .ZN(n8905) );
  OAI21_X1 U8066 ( .B1(n8550), .B2(n8480), .A(n8483), .ZN(n8537) );
  OAI21_X1 U8067 ( .B1(n8560), .B2(n8559), .A(n8479), .ZN(n8550) );
  NAND2_X1 U8068 ( .A1(n8264), .A2(n8263), .ZN(n8261) );
  NOR2_X1 U8069 ( .A1(n8588), .A2(SI_20_), .ZN(n8264) );
  NAND2_X1 U8070 ( .A1(n8588), .A2(SI_20_), .ZN(n8263) );
  OR2_X1 U8071 ( .A1(n8449), .A2(n11069), .ZN(n8450) );
  NOR2_X1 U8072 ( .A1(n8246), .A2(n7840), .ZN(n7839) );
  OR2_X1 U8073 ( .A1(n8418), .A2(n8417), .ZN(n8419) );
  NAND2_X1 U8074 ( .A1(n8394), .A2(n7637), .ZN(n7636) );
  NOR2_X1 U8075 ( .A1(n15825), .A2(n15824), .ZN(n15835) );
  INV_X1 U8076 ( .A(n8125), .ZN(n8123) );
  OAI21_X1 U8077 ( .B1(n7436), .B2(n8122), .A(n8121), .ZN(n8120) );
  NOR2_X1 U8078 ( .A1(n7461), .A2(n8123), .ZN(n8122) );
  NAND2_X1 U8079 ( .A1(n7436), .A2(n8125), .ZN(n8121) );
  AND2_X1 U8080 ( .A1(n9796), .A2(n9795), .ZN(n7867) );
  AND4_X1 U8081 ( .A1(n9486), .A2(n9485), .A3(n9484), .A4(n9483), .ZN(n12601)
         );
  AND3_X1 U8082 ( .A1(n9326), .A2(n9327), .A3(n9325), .ZN(n7935) );
  NAND2_X1 U8083 ( .A1(n10143), .A2(n10142), .ZN(n10825) );
  NAND2_X1 U8084 ( .A1(n7990), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7987) );
  AOI21_X1 U8085 ( .B1(n10854), .B2(n10112), .A(n10187), .ZN(n7991) );
  OR2_X1 U8086 ( .A1(n15995), .A2(n10148), .ZN(n7912) );
  OR2_X1 U8087 ( .A1(n16011), .A2(n10152), .ZN(n7902) );
  NAND2_X1 U8088 ( .A1(n7902), .A2(n7901), .ZN(n11623) );
  INV_X1 U8089 ( .A(n11620), .ZN(n7901) );
  XNOR2_X1 U8090 ( .A(n7979), .B(n14072), .ZN(n14067) );
  AOI21_X1 U8091 ( .B1(n10242), .B2(n10729), .A(n10241), .ZN(n10243) );
  AOI22_X1 U8092 ( .A1(n12528), .A2(n9916), .B1(SI_27_), .B2(n9686), .ZN(n9860) );
  NOR2_X1 U8093 ( .A1(n14221), .A2(n9936), .ZN(n8345) );
  OAI21_X1 U8094 ( .B1(n9738), .B2(n7701), .A(n7698), .ZN(n14198) );
  INV_X1 U8095 ( .A(n7702), .ZN(n7701) );
  AND2_X1 U8096 ( .A1(n9929), .A2(n9931), .ZN(n14199) );
  NOR2_X1 U8097 ( .A1(n14227), .A2(n14360), .ZN(n7647) );
  NAND2_X1 U8098 ( .A1(n14235), .A2(n10039), .ZN(n14217) );
  AND2_X1 U8099 ( .A1(n14217), .A2(n14221), .ZN(n14219) );
  OAI21_X1 U8100 ( .B1(n14309), .B2(n7697), .A(n7695), .ZN(n14292) );
  AND2_X1 U8101 ( .A1(n9942), .A2(n9736), .ZN(n14293) );
  NAND2_X1 U8102 ( .A1(n14309), .A2(n9576), .ZN(n14308) );
  AND4_X1 U8103 ( .A1(n9575), .A2(n9574), .A3(n9573), .A4(n9572), .ZN(n14316)
         );
  NOR2_X1 U8104 ( .A1(n14333), .A2(n7937), .ZN(n7936) );
  INV_X1 U8105 ( .A(n9524), .ZN(n7937) );
  AOI21_X1 U8106 ( .B1(n7690), .B2(n9999), .A(n7688), .ZN(n7687) );
  INV_X1 U8107 ( .A(n10006), .ZN(n7688) );
  INV_X1 U8108 ( .A(n7691), .ZN(n7690) );
  OAI21_X1 U8109 ( .B1(n7439), .B2(n9999), .A(n13213), .ZN(n7691) );
  AOI21_X1 U8110 ( .B1(n7946), .B2(n7944), .A(n7560), .ZN(n7943) );
  OR2_X1 U8111 ( .A1(n16232), .A2(n14050), .ZN(n13177) );
  NAND2_X1 U8112 ( .A1(n12495), .A2(n9800), .ZN(n7948) );
  AND2_X1 U8113 ( .A1(n13177), .A2(n9993), .ZN(n12600) );
  NAND2_X1 U8114 ( .A1(n12320), .A2(n9440), .ZN(n12495) );
  NAND2_X1 U8115 ( .A1(n11959), .A2(n7469), .ZN(n12286) );
  INV_X1 U8116 ( .A(n11957), .ZN(n11960) );
  AND2_X1 U8117 ( .A1(n11804), .A2(n9339), .ZN(n7953) );
  NAND2_X1 U8118 ( .A1(n7706), .A2(n7485), .ZN(n16049) );
  INV_X1 U8119 ( .A(n7707), .ZN(n7706) );
  OR2_X1 U8120 ( .A1(n9917), .A2(n12989), .ZN(n9290) );
  AND2_X1 U8121 ( .A1(n9750), .A2(n9749), .ZN(n10393) );
  INV_X1 U8122 ( .A(n16103), .ZN(n14391) );
  OR2_X1 U8123 ( .A1(n9882), .A2(n10043), .ZN(n16054) );
  AND2_X1 U8124 ( .A1(n10105), .A2(n14467), .ZN(n10395) );
  INV_X1 U8125 ( .A(n12463), .ZN(n9227) );
  OR2_X1 U8126 ( .A1(n9895), .A2(n9894), .ZN(n9897) );
  INV_X1 U8127 ( .A(n9715), .ZN(n10164) );
  INV_X1 U8128 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n9222) );
  AND2_X1 U8129 ( .A1(n8141), .A2(n8139), .ZN(n8138) );
  INV_X1 U8130 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8139) );
  NOR2_X1 U8131 ( .A1(n9597), .A2(n7759), .ZN(n7758) );
  INV_X1 U8132 ( .A(n9176), .ZN(n7759) );
  NAND2_X1 U8133 ( .A1(n9561), .A2(n9174), .ZN(n9580) );
  NAND2_X1 U8134 ( .A1(n9162), .A2(n10727), .ZN(n9164) );
  OAI21_X1 U8135 ( .B1(n9163), .B2(n7735), .A(n7734), .ZN(n9490) );
  INV_X1 U8136 ( .A(n9164), .ZN(n7735) );
  AOI21_X1 U8137 ( .B1(n9164), .B2(n10725), .A(n8300), .ZN(n7734) );
  INV_X1 U8138 ( .A(n9487), .ZN(n8300) );
  NOR2_X1 U8139 ( .A1(n9492), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n9514) );
  NAND2_X1 U8140 ( .A1(n8301), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n9473) );
  INV_X1 U8141 ( .A(n9471), .ZN(n8301) );
  INV_X1 U8142 ( .A(n7741), .ZN(n7740) );
  OAI21_X1 U8143 ( .B1(n9154), .B2(n7742), .A(n9430), .ZN(n7741) );
  INV_X1 U8144 ( .A(n9155), .ZN(n7742) );
  NAND2_X1 U8145 ( .A1(n9414), .A2(n9154), .ZN(n7739) );
  XNOR2_X1 U8146 ( .A(n9401), .B(P3_IR_REG_8__SCAN_IN), .ZN(n10479) );
  AOI21_X1 U8147 ( .B1(n9352), .B2(n7771), .A(n7450), .ZN(n7769) );
  XNOR2_X1 U8148 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n9371) );
  NAND2_X1 U8149 ( .A1(n9144), .A2(n9143), .ZN(n9354) );
  NAND2_X1 U8150 ( .A1(n7746), .A2(n7745), .ZN(n9335) );
  AND2_X1 U8151 ( .A1(n7750), .A2(n9139), .ZN(n7745) );
  INV_X1 U8152 ( .A(n9332), .ZN(n7750) );
  NAND2_X1 U8153 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n7749), .ZN(n7748) );
  NAND3_X1 U8154 ( .A1(n9285), .A2(n7510), .A3(n9138), .ZN(n7747) );
  XNOR2_X1 U8155 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .ZN(n9137) );
  INV_X1 U8156 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7910) );
  OR2_X1 U8157 ( .A1(n12476), .A2(n8109), .ZN(n8103) );
  NAND2_X1 U8158 ( .A1(n7519), .A2(n8115), .ZN(n8110) );
  NAND2_X1 U8159 ( .A1(n12475), .A2(n12474), .ZN(n8114) );
  AND2_X1 U8160 ( .A1(n10941), .A2(n10308), .ZN(n14563) );
  OR2_X1 U8161 ( .A1(n13423), .A2(n13376), .ZN(n13436) );
  AOI21_X1 U8162 ( .B1(n8090), .B2(n11742), .A(n7464), .ZN(n8088) );
  INV_X1 U8163 ( .A(n8090), .ZN(n8089) );
  INV_X1 U8164 ( .A(n8110), .ZN(n8109) );
  AND2_X1 U8165 ( .A1(n12585), .A2(n8108), .ZN(n8107) );
  NAND2_X1 U8166 ( .A1(n8110), .A2(n8112), .ZN(n8108) );
  AND2_X1 U8167 ( .A1(n13662), .A2(n7420), .ZN(n10539) );
  INV_X1 U8168 ( .A(n13522), .ZN(n13504) );
  NAND4_X2 U8169 ( .A1(n10316), .A2(n10313), .A3(n10315), .A4(n10314), .ZN(
        n14691) );
  NAND2_X1 U8170 ( .A1(n10328), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n10313) );
  NOR2_X1 U8171 ( .A1(n14785), .A2(n7967), .ZN(n14759) );
  INV_X1 U8172 ( .A(n7969), .ZN(n7967) );
  NAND2_X1 U8173 ( .A1(n7972), .A2(n7971), .ZN(n14845) );
  INV_X1 U8174 ( .A(n13642), .ZN(n7633) );
  NAND2_X1 U8175 ( .A1(n12027), .A2(n8033), .ZN(n12119) );
  OAI21_X1 U8176 ( .B1(n11692), .B2(n8155), .A(n8153), .ZN(n11871) );
  AOI21_X1 U8177 ( .B1(n8156), .B2(n8154), .A(n7492), .ZN(n8153) );
  INV_X1 U8178 ( .A(n8156), .ZN(n8155) );
  INV_X1 U8179 ( .A(n11870), .ZN(n8154) );
  AND2_X1 U8180 ( .A1(n10658), .A2(n15647), .ZN(n14929) );
  INV_X1 U8181 ( .A(n13527), .ZN(n13528) );
  AOI21_X1 U8182 ( .B1(n14951), .B2(n14902), .A(n7655), .ZN(n14953) );
  INV_X1 U8183 ( .A(n10363), .ZN(n15027) );
  XNOR2_X1 U8184 ( .A(n10096), .B(n10261), .ZN(n13243) );
  NAND2_X1 U8185 ( .A1(n10099), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10102) );
  INV_X1 U8186 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n10411) );
  INV_X1 U8187 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n10303) );
  NAND2_X1 U8188 ( .A1(n8171), .A2(n8173), .ZN(n8170) );
  INV_X1 U8189 ( .A(n7666), .ZN(n7665) );
  OAI21_X1 U8190 ( .B1(n7458), .B2(n8171), .A(n7667), .ZN(n7666) );
  OR2_X1 U8191 ( .A1(n13293), .A2(n13292), .ZN(n7667) );
  INV_X1 U8192 ( .A(n8183), .ZN(n8178) );
  AOI21_X1 U8193 ( .B1(n8183), .B2(n8185), .A(n7514), .ZN(n8182) );
  AND2_X1 U8194 ( .A1(n13312), .A2(n13310), .ZN(n8210) );
  OAI21_X1 U8195 ( .B1(n7569), .B2(n8205), .A(n11468), .ZN(n8204) );
  AND2_X1 U8196 ( .A1(n8198), .A2(n11463), .ZN(n8194) );
  CLKBUF_X3 U8197 ( .A(n8762), .Z(n8921) );
  AND2_X1 U8198 ( .A1(n8380), .A2(n8381), .ZN(n8762) );
  AND2_X1 U8199 ( .A1(n8381), .A2(n8795), .ZN(n8761) );
  OR2_X1 U8200 ( .A1(n10782), .A2(n10781), .ZN(n7726) );
  OR2_X1 U8201 ( .A1(n10790), .A2(n10791), .ZN(n7709) );
  OR2_X1 U8202 ( .A1(n8683), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n8647) );
  NOR2_X1 U8203 ( .A1(n12618), .A2(n7719), .ZN(n12620) );
  AND2_X1 U8204 ( .A1(n12619), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7719) );
  NOR2_X1 U8205 ( .A1(n15205), .A2(n7714), .ZN(n15208) );
  AND2_X1 U8206 ( .A1(n15206), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n7714) );
  OR2_X1 U8207 ( .A1(n15208), .A2(n15207), .ZN(n7713) );
  XNOR2_X1 U8208 ( .A(n7711), .B(n15233), .ZN(n15217) );
  NAND2_X1 U8209 ( .A1(n7713), .A2(n7712), .ZN(n7711) );
  NAND2_X1 U8210 ( .A1(n15216), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n7712) );
  INV_X1 U8211 ( .A(n7619), .ZN(n15269) );
  NOR2_X1 U8212 ( .A1(n15334), .A2(n8259), .ZN(n8258) );
  NAND2_X1 U8213 ( .A1(n15321), .A2(n8257), .ZN(n8256) );
  INV_X1 U8214 ( .A(n8258), .ZN(n8257) );
  NOR2_X1 U8215 ( .A1(n15326), .A2(n15330), .ZN(n15325) );
  AOI21_X1 U8216 ( .B1(n7434), .B2(n15402), .A(n7516), .ZN(n7779) );
  INV_X1 U8217 ( .A(n7434), .ZN(n7780) );
  INV_X1 U8218 ( .A(n8276), .ZN(n15400) );
  OAI21_X1 U8219 ( .B1(n15450), .B2(n8279), .A(n8277), .ZN(n8276) );
  NAND2_X1 U8220 ( .A1(n8283), .A2(n13334), .ZN(n8279) );
  AOI21_X1 U8221 ( .B1(n8278), .B2(n13334), .A(n13333), .ZN(n8277) );
  AOI21_X1 U8222 ( .B1(n8283), .B2(n8281), .A(n7507), .ZN(n8280) );
  INV_X1 U8223 ( .A(n15461), .ZN(n8281) );
  NOR2_X1 U8224 ( .A1(n16301), .A2(n7789), .ZN(n12694) );
  AND2_X1 U8225 ( .A1(n15089), .A2(n16321), .ZN(n7789) );
  NAND2_X1 U8226 ( .A1(n7790), .A2(n8292), .ZN(n8289) );
  INV_X1 U8227 ( .A(n16244), .ZN(n7790) );
  AOI21_X1 U8228 ( .B1(n8021), .B2(n7466), .A(n8019), .ZN(n8018) );
  NOR2_X1 U8229 ( .A1(n12693), .A2(n15183), .ZN(n8019) );
  INV_X1 U8230 ( .A(n12650), .ZN(n12697) );
  INV_X1 U8231 ( .A(n15184), .ZN(n12687) );
  NAND3_X1 U8232 ( .A1(n16224), .A2(n8061), .A3(n16165), .ZN(n16246) );
  NOR2_X1 U8233 ( .A1(n16266), .A2(n8062), .ZN(n8061) );
  INV_X1 U8234 ( .A(n8063), .ZN(n8062) );
  NAND2_X1 U8235 ( .A1(n16249), .A2(n12687), .ZN(n8294) );
  OR2_X1 U8236 ( .A1(n12485), .A2(n8021), .ZN(n16250) );
  NAND2_X1 U8237 ( .A1(n8695), .A2(n8694), .ZN(n12272) );
  OR2_X1 U8238 ( .A1(n16156), .A2(n16157), .ZN(n16154) );
  AND2_X1 U8239 ( .A1(n13268), .A2(n10879), .ZN(n11295) );
  NOR2_X1 U8240 ( .A1(n11496), .A2(n16113), .ZN(n7787) );
  NAND2_X1 U8241 ( .A1(n11496), .A2(n16113), .ZN(n7788) );
  NAND2_X1 U8242 ( .A1(n11306), .A2(n11305), .ZN(n11490) );
  NAND2_X1 U8243 ( .A1(n7582), .A2(n7484), .ZN(n11306) );
  CLKBUF_X1 U8244 ( .A(n8003), .Z(n7599) );
  OR2_X1 U8245 ( .A1(n7599), .A2(n10874), .ZN(n11007) );
  AOI21_X1 U8246 ( .B1(n15476), .B2(n16247), .A(n15475), .ZN(n8008) );
  AND2_X1 U8247 ( .A1(n16254), .A2(n16135), .ZN(n16299) );
  OR2_X1 U8248 ( .A1(n8772), .A2(n10465), .ZN(n8778) );
  OR2_X1 U8249 ( .A1(n10455), .A2(n10618), .ZN(n8776) );
  NAND2_X1 U8250 ( .A1(n10528), .A2(n10533), .ZN(n16333) );
  OR2_X1 U8251 ( .A1(n10881), .A2(n15606), .ZN(n16031) );
  AND2_X1 U8252 ( .A1(n8497), .A2(n8500), .ZN(n8299) );
  INV_X1 U8253 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8497) );
  AND2_X2 U8254 ( .A1(n8371), .A2(n8370), .ZN(n8603) );
  NOR2_X1 U8255 ( .A1(n9105), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n8189) );
  AND2_X1 U8256 ( .A1(n7670), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n7669) );
  OR2_X1 U8257 ( .A1(n7672), .A2(n7671), .ZN(n7670) );
  NAND2_X1 U8258 ( .A1(n9103), .A2(n9100), .ZN(n9112) );
  XNOR2_X1 U8259 ( .A(n8520), .B(P1_IR_REG_23__SCAN_IN), .ZN(n10454) );
  INV_X1 U8260 ( .A(n7577), .ZN(n15790) );
  AOI21_X1 U8261 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n15854), .A(n15853), .ZN(
        n15858) );
  OAI21_X1 U8262 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n15890), .A(n15889), .ZN(
        n15900) );
  NAND2_X1 U8263 ( .A1(n11944), .A2(n9786), .ZN(n12049) );
  NAND2_X1 U8264 ( .A1(n13989), .A2(n7488), .ZN(n7850) );
  OAI21_X1 U8265 ( .B1(n7861), .B2(n7855), .A(n7848), .ZN(n7847) );
  NAND2_X1 U8266 ( .A1(n7849), .A2(n7855), .ZN(n7848) );
  NAND2_X1 U8267 ( .A1(n7853), .A2(n13928), .ZN(n7849) );
  NAND2_X1 U8268 ( .A1(n7852), .A2(n7861), .ZN(n7851) );
  INV_X1 U8269 ( .A(n7853), .ZN(n7852) );
  NAND2_X1 U8270 ( .A1(n12639), .A2(n8135), .ZN(n13194) );
  AND2_X1 U8271 ( .A1(n13196), .A2(n9808), .ZN(n8135) );
  NAND2_X1 U8272 ( .A1(n9776), .A2(n9775), .ZN(n11413) );
  AND2_X1 U8273 ( .A1(n9447), .A2(n9446), .ZN(n12712) );
  NAND2_X1 U8274 ( .A1(n7854), .A2(n7857), .ZN(n14022) );
  INV_X1 U8275 ( .A(n14017), .ZN(n16037) );
  OAI21_X1 U8276 ( .B1(n10081), .B2(n10080), .A(n7447), .ZN(n7705) );
  INV_X1 U8277 ( .A(n14244), .ZN(n14371) );
  INV_X1 U8278 ( .A(n14268), .ZN(n14383) );
  NAND2_X2 U8279 ( .A1(n9328), .A2(n7935), .ZN(n11806) );
  INV_X1 U8280 ( .A(n7904), .ZN(n10239) );
  NOR2_X1 U8281 ( .A1(n14115), .A2(n14116), .ZN(n14119) );
  OR2_X1 U8282 ( .A1(n14127), .A2(n7918), .ZN(n7917) );
  INV_X1 U8283 ( .A(n7914), .ZN(n7913) );
  AOI21_X1 U8284 ( .B1(n14132), .B2(n16017), .A(n14131), .ZN(n7914) );
  NAND2_X1 U8285 ( .A1(n7917), .A2(n7916), .ZN(n14136) );
  NAND2_X1 U8286 ( .A1(n7957), .A2(n7471), .ZN(n7956) );
  NAND2_X1 U8287 ( .A1(n9699), .A2(n9698), .ZN(n14347) );
  NAND2_X1 U8288 ( .A1(n14178), .A2(n14304), .ZN(n7626) );
  AND2_X1 U8289 ( .A1(n9683), .A2(n9682), .ZN(n14186) );
  INV_X1 U8290 ( .A(n9860), .ZN(n14352) );
  NAND2_X1 U8291 ( .A1(n9675), .A2(n9674), .ZN(n14356) );
  NAND2_X1 U8292 ( .A1(n9738), .A2(n10036), .ZN(n14233) );
  NAND2_X1 U8293 ( .A1(n9635), .A2(n9634), .ZN(n14372) );
  NAND2_X1 U8294 ( .A1(n9610), .A2(n9609), .ZN(n14385) );
  NAND2_X1 U8295 ( .A1(n9600), .A2(n9599), .ZN(n14389) );
  INV_X1 U8296 ( .A(n12075), .ZN(n12263) );
  NAND2_X1 U8297 ( .A1(n13477), .A2(n13476), .ZN(n14964) );
  NAND2_X1 U8298 ( .A1(n8084), .A2(n8083), .ZN(n8082) );
  INV_X1 U8299 ( .A(n11135), .ZN(n8083) );
  NOR2_X1 U8300 ( .A1(n14595), .A2(n14594), .ZN(n14593) );
  INV_X1 U8301 ( .A(n14811), .ZN(n14662) );
  AND2_X1 U8302 ( .A1(n10937), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14667) );
  INV_X1 U8303 ( .A(n14642), .ZN(n14658) );
  AND2_X1 U8304 ( .A1(n13889), .A2(n13888), .ZN(n13890) );
  AND2_X1 U8305 ( .A1(n13515), .A2(n13514), .ZN(n13871) );
  INV_X1 U8306 ( .A(n14946), .ZN(n8161) );
  XNOR2_X1 U8307 ( .A(n13550), .B(n7600), .ZN(n14947) );
  NAND2_X1 U8308 ( .A1(n14764), .A2(n14902), .ZN(n7605) );
  AOI22_X1 U8309 ( .A1(n14795), .A2(n14885), .B1(n14883), .B2(n14819), .ZN(
        n7587) );
  NAND2_X1 U8310 ( .A1(n14796), .A2(n14924), .ZN(n7586) );
  INV_X1 U8311 ( .A(n14851), .ZN(n8167) );
  NAND2_X1 U8312 ( .A1(n8162), .A2(n8163), .ZN(n14850) );
  NAND2_X1 U8313 ( .A1(n8166), .A2(n13539), .ZN(n14861) );
  OR2_X1 U8314 ( .A1(n14873), .A2(n13538), .ZN(n8166) );
  NAND2_X1 U8315 ( .A1(n14843), .A2(n11364), .ZN(n14932) );
  NAND2_X1 U8316 ( .A1(n14843), .A2(n11362), .ZN(n14933) );
  AND2_X1 U8317 ( .A1(n10354), .A2(n10353), .ZN(n15648) );
  NOR2_X1 U8318 ( .A1(n7444), .A2(n15175), .ZN(n7675) );
  NAND2_X1 U8319 ( .A1(n7678), .A2(n7681), .ZN(n7677) );
  NAND2_X1 U8320 ( .A1(n7682), .A2(n13586), .ZN(n7681) );
  INV_X1 U8321 ( .A(n15076), .ZN(n7682) );
  NAND2_X1 U8322 ( .A1(n13555), .A2(n13554), .ZN(n15095) );
  OR2_X1 U8323 ( .A1(n8772), .A2(n10421), .ZN(n8749) );
  NAND2_X1 U8324 ( .A1(n8798), .A2(n8797), .ZN(n15197) );
  NOR2_X1 U8325 ( .A1(n10968), .A2(n7727), .ZN(n10782) );
  AND2_X1 U8326 ( .A1(n10622), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7727) );
  NOR2_X1 U8327 ( .A1(n10816), .A2(n10815), .ZN(n10814) );
  NAND2_X1 U8328 ( .A1(n10679), .A2(n7710), .ZN(n10790) );
  OR2_X1 U8329 ( .A1(n10680), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n7710) );
  XNOR2_X1 U8330 ( .A(n12620), .B(n12627), .ZN(n15762) );
  NAND2_X1 U8331 ( .A1(n15762), .A2(n16340), .ZN(n15761) );
  OR2_X1 U8332 ( .A1(n15759), .A2(n15750), .ZN(n15240) );
  XNOR2_X1 U8333 ( .A(n13343), .B(n13342), .ZN(n15478) );
  NAND2_X1 U8334 ( .A1(n8920), .A2(n8919), .ZN(n15274) );
  NAND2_X1 U8335 ( .A1(n11508), .A2(n11487), .ZN(n11640) );
  INV_X1 U8336 ( .A(n15848), .ZN(n7929) );
  NAND2_X1 U8337 ( .A1(n7575), .A2(n7574), .ZN(n7585) );
  INV_X1 U8338 ( .A(n15879), .ZN(n7574) );
  INV_X1 U8339 ( .A(n8972), .ZN(n8235) );
  NOR2_X1 U8340 ( .A1(n8975), .A2(n8972), .ZN(n8236) );
  OAI21_X1 U8341 ( .B1(n13688), .B2(n13687), .A(n13686), .ZN(n13698) );
  INV_X1 U8342 ( .A(n8984), .ZN(n8237) );
  NOR2_X1 U8343 ( .A1(n8987), .A2(n8984), .ZN(n8238) );
  OAI211_X1 U8344 ( .C1(n13709), .C2(n7794), .A(n7797), .B(n7631), .ZN(n8312)
         );
  INV_X1 U8345 ( .A(n13713), .ZN(n7631) );
  NOR2_X1 U8346 ( .A1(n8996), .A2(n8999), .ZN(n8223) );
  NAND2_X1 U8347 ( .A1(n8999), .A2(n8996), .ZN(n8222) );
  NAND2_X1 U8348 ( .A1(n8223), .A2(n8222), .ZN(n8220) );
  NAND2_X1 U8349 ( .A1(n13731), .A2(n7451), .ZN(n7588) );
  NAND2_X1 U8350 ( .A1(n9005), .A2(n9007), .ZN(n7880) );
  NAND2_X1 U8351 ( .A1(n9020), .A2(n7890), .ZN(n7889) );
  NOR2_X1 U8352 ( .A1(n9026), .A2(n9023), .ZN(n8230) );
  NAND2_X1 U8353 ( .A1(n9026), .A2(n9023), .ZN(n8229) );
  NOR2_X1 U8354 ( .A1(n8230), .A2(n7887), .ZN(n7886) );
  INV_X1 U8355 ( .A(n7889), .ZN(n7887) );
  INV_X1 U8356 ( .A(n8229), .ZN(n7884) );
  AND2_X1 U8357 ( .A1(n9022), .A2(n7892), .ZN(n7891) );
  INV_X1 U8358 ( .A(n9020), .ZN(n7892) );
  NAND2_X1 U8359 ( .A1(n13777), .A2(n7481), .ZN(n8334) );
  NAND2_X1 U8360 ( .A1(n7612), .A2(n7874), .ZN(n9035) );
  NAND2_X1 U8361 ( .A1(n9031), .A2(n7875), .ZN(n7874) );
  NOR2_X1 U8362 ( .A1(n7503), .A2(n7652), .ZN(n7651) );
  NOR2_X1 U8363 ( .A1(n8243), .A2(n9043), .ZN(n7652) );
  INV_X1 U8364 ( .A(n9041), .ZN(n8243) );
  NOR2_X1 U8365 ( .A1(n9044), .A2(n9041), .ZN(n8244) );
  NAND2_X1 U8366 ( .A1(n7463), .A2(n8332), .ZN(n8330) );
  AND2_X1 U8367 ( .A1(n13337), .A2(n8232), .ZN(n8231) );
  NAND2_X1 U8368 ( .A1(n9055), .A2(n9057), .ZN(n8232) );
  NAND2_X1 U8369 ( .A1(n9063), .A2(n7879), .ZN(n7878) );
  NOR2_X1 U8370 ( .A1(n9068), .A2(n9065), .ZN(n8240) );
  INV_X1 U8371 ( .A(n9065), .ZN(n8239) );
  NAND2_X1 U8372 ( .A1(n9939), .A2(n10129), .ZN(n8306) );
  INV_X1 U8373 ( .A(n9939), .ZN(n8309) );
  INV_X1 U8374 ( .A(n14754), .ZN(n7819) );
  NAND2_X1 U8375 ( .A1(n8234), .A2(n9077), .ZN(n8233) );
  NOR2_X1 U8376 ( .A1(n8625), .A2(n8641), .ZN(n8249) );
  NAND2_X1 U8377 ( .A1(n8250), .A2(n7846), .ZN(n7845) );
  INV_X1 U8378 ( .A(n8625), .ZN(n8250) );
  INV_X1 U8379 ( .A(n8447), .ZN(n8248) );
  NAND2_X1 U8380 ( .A1(n8302), .A2(n7744), .ZN(n10049) );
  NAND2_X1 U8381 ( .A1(n8303), .A2(n7471), .ZN(n8302) );
  AND2_X1 U8382 ( .A1(n10046), .A2(n7532), .ZN(n7743) );
  NAND2_X1 U8383 ( .A1(n8325), .A2(n13850), .ZN(n8324) );
  AOI21_X1 U8384 ( .B1(n13838), .B2(n7802), .A(n7800), .ZN(n13852) );
  NOR2_X1 U8385 ( .A1(n8329), .A2(n7803), .ZN(n7802) );
  INV_X1 U8386 ( .A(n7804), .ZN(n7803) );
  INV_X1 U8387 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n10091) );
  NAND2_X1 U8388 ( .A1(n8457), .A2(n12956), .ZN(n8460) );
  NAND2_X1 U8389 ( .A1(n8681), .A2(n8433), .ZN(n8270) );
  INV_X1 U8390 ( .A(n8437), .ZN(n8266) );
  INV_X1 U8391 ( .A(n8433), .ZN(n8267) );
  NOR2_X1 U8392 ( .A1(n8247), .A2(n12974), .ZN(n7841) );
  INV_X1 U8393 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n8643) );
  OAI21_X1 U8394 ( .B1(n8767), .B2(n10425), .A(n7603), .ZN(n8412) );
  NAND2_X1 U8395 ( .A1(n8767), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7603) );
  INV_X1 U8396 ( .A(n7922), .ZN(n15813) );
  NOR2_X1 U8397 ( .A1(n11724), .A2(n8134), .ZN(n8133) );
  INV_X1 U8398 ( .A(n9778), .ZN(n8134) );
  INV_X1 U8399 ( .A(n9781), .ZN(n8132) );
  OAI21_X1 U8400 ( .B1(n8133), .B2(n8132), .A(n11832), .ZN(n8131) );
  OR2_X1 U8401 ( .A1(n10112), .A2(n10187), .ZN(n7990) );
  AND2_X1 U8402 ( .A1(n10235), .A2(n10234), .ZN(n10236) );
  INV_X1 U8403 ( .A(n8343), .ZN(n8342) );
  INV_X1 U8404 ( .A(n10039), .ZN(n7703) );
  INV_X1 U8405 ( .A(n8339), .ZN(n7699) );
  AOI21_X1 U8406 ( .B1(n8343), .B2(n8341), .A(n8340), .ZN(n8339) );
  INV_X1 U8407 ( .A(n14199), .ZN(n8340) );
  INV_X1 U8408 ( .A(n8344), .ZN(n8341) );
  INV_X1 U8409 ( .A(n7704), .ZN(n7700) );
  OR2_X1 U8410 ( .A1(n9676), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9687) );
  OR2_X1 U8411 ( .A1(n9636), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9637) );
  AND2_X1 U8412 ( .A1(n14236), .A2(n10036), .ZN(n7704) );
  NAND2_X1 U8413 ( .A1(n9611), .A2(n12787), .ZN(n9636) );
  NOR2_X1 U8414 ( .A1(n7945), .A2(n7942), .ZN(n7941) );
  INV_X1 U8415 ( .A(n9440), .ZN(n7942) );
  INV_X1 U8416 ( .A(n7946), .ZN(n7945) );
  INV_X1 U8417 ( .A(n9800), .ZN(n7944) );
  NOR2_X1 U8418 ( .A1(n9463), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9481) );
  INV_X1 U8419 ( .A(n11767), .ZN(n10400) );
  INV_X1 U8420 ( .A(n7763), .ZN(n7761) );
  INV_X1 U8421 ( .A(n9684), .ZN(n7764) );
  NOR2_X1 U8422 ( .A1(n7771), .A2(n9148), .ZN(n7768) );
  INV_X1 U8423 ( .A(n11125), .ZN(n14487) );
  NAND2_X1 U8424 ( .A1(n7418), .A2(n7969), .ZN(n7968) );
  INV_X1 U8425 ( .A(n13542), .ZN(n8146) );
  NOR2_X1 U8426 ( .A1(n14874), .A2(n14987), .ZN(n7972) );
  AOI21_X1 U8427 ( .B1(n14855), .B2(n13445), .A(n13444), .ZN(n14834) );
  NOR2_X1 U8428 ( .A1(n12555), .A2(n15011), .ZN(n13530) );
  OR2_X1 U8429 ( .A1(n12108), .A2(n12107), .ZN(n12190) );
  NOR2_X1 U8430 ( .A1(n12200), .A2(n13770), .ZN(n7976) );
  OR2_X1 U8431 ( .A1(n12123), .A2(n13758), .ZN(n12200) );
  INV_X1 U8432 ( .A(n8033), .ZN(n8031) );
  AND2_X1 U8433 ( .A1(n13634), .A2(n8157), .ZN(n8156) );
  NAND2_X1 U8434 ( .A1(n11691), .A2(n11870), .ZN(n8157) );
  OR2_X1 U8435 ( .A1(n11677), .A2(n11676), .ZN(n11864) );
  INV_X1 U8436 ( .A(n11538), .ZN(n8046) );
  OR2_X1 U8437 ( .A1(n13662), .A2(n13902), .ZN(n8075) );
  INV_X1 U8438 ( .A(n14912), .ZN(n14911) );
  INV_X1 U8439 ( .A(n14897), .ZN(n8027) );
  INV_X1 U8440 ( .A(n14896), .ZN(n8028) );
  AND2_X1 U8441 ( .A1(n13902), .A2(n10662), .ZN(n13665) );
  AND2_X1 U8442 ( .A1(n10094), .A2(n10093), .ZN(n8040) );
  AND2_X1 U8443 ( .A1(n10410), .A2(n8039), .ZN(n8038) );
  AND2_X1 U8444 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(n8322), .ZN(n8039) );
  OAI21_X1 U8445 ( .B1(P2_IR_REG_31__SCAN_IN), .B2(n8043), .A(n8044), .ZN(
        n8042) );
  NAND2_X1 U8446 ( .A1(n8043), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8044) );
  NOR2_X1 U8447 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n10095) );
  CLKBUF_X1 U8448 ( .A(n11769), .Z(n12233) );
  OR2_X1 U8449 ( .A1(n10419), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n10651) );
  INV_X1 U8450 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n10414) );
  AND2_X1 U8451 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n8880), .ZN(n8564) );
  NAND2_X1 U8452 ( .A1(n7774), .A2(n7476), .ZN(n8297) );
  OR2_X1 U8453 ( .A1(n15341), .A2(n15342), .ZN(n7774) );
  INV_X1 U8454 ( .A(n8280), .ZN(n8278) );
  AND2_X1 U8455 ( .A1(n15542), .A2(n15182), .ZN(n13333) );
  INV_X1 U8456 ( .A(n12487), .ZN(n8020) );
  NAND2_X1 U8457 ( .A1(n12488), .A2(n7473), .ZN(n16244) );
  NOR2_X1 U8458 ( .A1(n12010), .A2(n12272), .ZN(n8063) );
  NAND2_X1 U8459 ( .A1(n16165), .A2(n16197), .ZN(n12000) );
  INV_X1 U8460 ( .A(n11301), .ZN(n11112) );
  INV_X1 U8461 ( .A(n16031), .ZN(n10528) );
  NAND2_X1 U8462 ( .A1(n8537), .A2(n8535), .ZN(n8487) );
  AND2_X1 U8463 ( .A1(n9107), .A2(n7673), .ZN(n7672) );
  INV_X1 U8464 ( .A(n8858), .ZN(n8245) );
  OR2_X1 U8465 ( .A1(n8455), .A2(n12736), .ZN(n8456) );
  NAND2_X1 U8466 ( .A1(n8442), .A2(SI_14_), .ZN(n8443) );
  NAND2_X1 U8467 ( .A1(n8427), .A2(SI_9_), .ZN(n8428) );
  INV_X1 U8468 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n12914) );
  OAI21_X1 U8469 ( .B1(SI_9_), .B2(n8427), .A(n8428), .ZN(n8705) );
  NAND2_X1 U8470 ( .A1(n7821), .A2(n7597), .ZN(n8716) );
  INV_X1 U8471 ( .A(n7598), .ZN(n7597) );
  OAI21_X1 U8472 ( .B1(n8419), .B2(n8726), .A(n8422), .ZN(n7598) );
  INV_X1 U8473 ( .A(n9107), .ZN(n8829) );
  INV_X1 U8474 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n15795) );
  AOI22_X1 U8475 ( .A1(n15835), .A2(n15834), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n15989), .ZN(n15840) );
  AOI21_X1 U8476 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n15877), .A(n15876), .ZN(
        n15888) );
  NOR2_X1 U8477 ( .A1(n15932), .A2(n15931), .ZN(n15937) );
  AND2_X1 U8478 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n15930), .ZN(n15931) );
  NAND2_X1 U8479 ( .A1(n7518), .A2(n7864), .ZN(n7853) );
  INV_X1 U8480 ( .A(n9854), .ZN(n7864) );
  INV_X1 U8481 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n11376) );
  INV_X1 U8482 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n13020) );
  AND2_X1 U8483 ( .A1(n9534), .A2(n9533), .ZN(n9552) );
  NAND2_X1 U8484 ( .A1(n11413), .A2(n8133), .ZN(n11721) );
  OR2_X1 U8485 ( .A1(n12322), .A2(n12501), .ZN(n9987) );
  INV_X1 U8486 ( .A(n11247), .ZN(n9292) );
  OR2_X1 U8487 ( .A1(n9360), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9379) );
  OR2_X1 U8488 ( .A1(n13943), .A2(n9854), .ZN(n7863) );
  OR2_X1 U8489 ( .A1(n10073), .A2(n8367), .ZN(n9925) );
  NAND2_X1 U8490 ( .A1(n7440), .A2(n8142), .ZN(n7733) );
  OR2_X1 U8491 ( .A1(n9293), .A2(n10169), .ZN(n9306) );
  OR2_X1 U8492 ( .A1(n11087), .A2(n15961), .ZN(n10834) );
  NAND2_X1 U8493 ( .A1(n7622), .A2(n10851), .ZN(n11151) );
  OR2_X1 U8494 ( .A1(n10110), .A2(n10441), .ZN(n7622) );
  NAND2_X1 U8495 ( .A1(n10855), .A2(n7596), .ZN(n10859) );
  NAND2_X1 U8496 ( .A1(n7919), .A2(n10856), .ZN(n11157) );
  INV_X1 U8497 ( .A(n7920), .ZN(n7919) );
  NAND2_X1 U8498 ( .A1(n15970), .A2(n7992), .ZN(n11027) );
  OR2_X1 U8499 ( .A1(n11025), .A2(n9340), .ZN(n15978) );
  AND2_X1 U8500 ( .A1(n15984), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7621) );
  OR2_X1 U8501 ( .A1(n9400), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n9415) );
  NAND2_X1 U8502 ( .A1(n7986), .A2(n7985), .ZN(n11615) );
  INV_X1 U8503 ( .A(n11617), .ZN(n7985) );
  OAI22_X1 U8504 ( .A1(n16016), .A2(n16015), .B1(n10202), .B2(n10478), .ZN(
        n11628) );
  NAND2_X1 U8505 ( .A1(n12129), .A2(n10157), .ZN(n7906) );
  OR2_X1 U8506 ( .A1(n10156), .A2(n10207), .ZN(n7907) );
  INV_X1 U8507 ( .A(n7979), .ZN(n10123) );
  XNOR2_X1 U8508 ( .A(n10236), .B(n7905), .ZN(n14087) );
  NOR2_X1 U8509 ( .A1(n14087), .A2(n14416), .ZN(n14086) );
  OR2_X1 U8510 ( .A1(n14106), .A2(n7984), .ZN(n7983) );
  AOI21_X1 U8511 ( .B1(n14101), .B2(n14100), .A(n14099), .ZN(n14103) );
  NAND2_X1 U8512 ( .A1(n14096), .A2(n14095), .ZN(n14128) );
  AND2_X1 U8513 ( .A1(n7957), .A2(n7548), .ZN(n7955) );
  INV_X1 U8514 ( .A(n7958), .ZN(n7957) );
  OAI21_X1 U8515 ( .B1(n7471), .B2(n9707), .A(n9714), .ZN(n7958) );
  OAI21_X1 U8516 ( .B1(n14189), .B2(n7515), .A(n8350), .ZN(n9923) );
  AOI21_X1 U8517 ( .B1(n8307), .B2(n9740), .A(n8351), .ZN(n8350) );
  INV_X1 U8518 ( .A(n10047), .ZN(n8351) );
  NAND2_X1 U8519 ( .A1(n14361), .A2(n8346), .ZN(n9671) );
  NOR2_X1 U8520 ( .A1(n9648), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9663) );
  OR2_X1 U8521 ( .A1(n9637), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9648) );
  INV_X1 U8522 ( .A(n9629), .ZN(n7952) );
  NAND2_X1 U8523 ( .A1(n14249), .A2(n9629), .ZN(n14237) );
  NAND2_X1 U8524 ( .A1(n14251), .A2(n14250), .ZN(n14249) );
  AND2_X1 U8525 ( .A1(n10030), .A2(n10031), .ZN(n14269) );
  NAND2_X1 U8526 ( .A1(n7694), .A2(n7692), .ZN(n14276) );
  AND2_X1 U8527 ( .A1(n9737), .A2(n7693), .ZN(n7692) );
  OR2_X1 U8528 ( .A1(n9568), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9584) );
  NAND2_X1 U8529 ( .A1(n9552), .A2(n13020), .ZN(n9568) );
  OR2_X1 U8530 ( .A1(n9449), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9463) );
  OR2_X1 U8531 ( .A1(n9423), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9449) );
  AND2_X1 U8532 ( .A1(n9987), .A2(n9992), .ZN(n12498) );
  AND2_X1 U8533 ( .A1(n9392), .A2(n11376), .ZN(n9406) );
  AOI21_X1 U8534 ( .B1(n7646), .B2(n7433), .A(n7645), .ZN(n8368) );
  INV_X1 U8535 ( .A(n7938), .ZN(n7645) );
  AOI21_X1 U8536 ( .B1(n7433), .B2(n7939), .A(n7498), .ZN(n7938) );
  NAND2_X1 U8537 ( .A1(n11843), .A2(n11842), .ZN(n11841) );
  OR2_X1 U8538 ( .A1(n9293), .A2(n10175), .ZN(n9314) );
  INV_X1 U8539 ( .A(n9959), .ZN(n7934) );
  INV_X1 U8540 ( .A(n10396), .ZN(n9321) );
  INV_X1 U8541 ( .A(n9948), .ZN(n16050) );
  NOR2_X1 U8542 ( .A1(n14059), .A2(n11481), .ZN(n11243) );
  OR2_X1 U8543 ( .A1(n9244), .A2(n14466), .ZN(n9880) );
  INV_X1 U8544 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n9274) );
  AOI21_X1 U8545 ( .B1(n9697), .B2(n9197), .A(n9196), .ZN(n9895) );
  NAND2_X1 U8546 ( .A1(n9672), .A2(n7457), .ZN(n7763) );
  NAND2_X1 U8547 ( .A1(n9193), .A2(n7571), .ZN(n7762) );
  INV_X1 U8548 ( .A(n9214), .ZN(n7870) );
  OR2_X1 U8549 ( .A1(n9188), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n9189) );
  XNOR2_X1 U8550 ( .A(n9188), .B(P2_DATAO_REG_24__SCAN_IN), .ZN(n9645) );
  NAND2_X1 U8551 ( .A1(n9620), .A2(n9184), .ZN(n9631) );
  AND2_X1 U8552 ( .A1(n9187), .A2(n9186), .ZN(n9630) );
  NAND2_X1 U8553 ( .A1(n9631), .A2(n9630), .ZN(n9633) );
  XNOR2_X1 U8554 ( .A(n9248), .B(n9247), .ZN(n10128) );
  NAND2_X1 U8555 ( .A1(n7753), .A2(n7751), .ZN(n9618) );
  AOI21_X1 U8556 ( .B1(n7755), .B2(n7757), .A(n7752), .ZN(n7751) );
  INV_X1 U8557 ( .A(n9181), .ZN(n7752) );
  AND2_X1 U8558 ( .A1(n9184), .A2(n9183), .ZN(n9617) );
  NAND2_X1 U8559 ( .A1(n8140), .A2(n8141), .ZN(n9253) );
  INV_X1 U8560 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n9578) );
  AND2_X1 U8561 ( .A1(n9174), .A2(n9173), .ZN(n9558) );
  INV_X1 U8562 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n9198) );
  AND2_X1 U8563 ( .A1(n9172), .A2(n9171), .ZN(n9542) );
  AND2_X1 U8564 ( .A1(n9170), .A2(n9169), .ZN(n9526) );
  AND2_X1 U8565 ( .A1(n9168), .A2(n9167), .ZN(n9508) );
  INV_X1 U8566 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n9513) );
  NAND2_X1 U8567 ( .A1(n9163), .A2(n9164), .ZN(n9471) );
  INV_X1 U8568 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n9474) );
  AND2_X1 U8569 ( .A1(n9161), .A2(n9160), .ZN(n9455) );
  AOI21_X1 U8570 ( .B1(n7740), .B2(n7742), .A(n7738), .ZN(n7737) );
  INV_X1 U8571 ( .A(n9157), .ZN(n7738) );
  AND2_X1 U8572 ( .A1(n9159), .A2(n9158), .ZN(n9441) );
  INV_X1 U8573 ( .A(n8353), .ZN(n9435) );
  XNOR2_X1 U8574 ( .A(n9386), .B(P3_IR_REG_7__SCAN_IN), .ZN(n10466) );
  OR2_X1 U8575 ( .A1(n9350), .A2(n9330), .ZN(n9331) );
  INV_X1 U8576 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8001) );
  NOR2_X1 U8577 ( .A1(n10140), .A2(n9330), .ZN(n8002) );
  OR2_X1 U8578 ( .A1(n12059), .A2(n12058), .ZN(n12060) );
  XNOR2_X1 U8579 ( .A(n15001), .B(n14553), .ZN(n14495) );
  NAND2_X1 U8580 ( .A1(n8102), .A2(n8100), .ZN(n8099) );
  INV_X1 U8581 ( .A(n14594), .ZN(n8100) );
  INV_X1 U8582 ( .A(n14541), .ZN(n8097) );
  XNOR2_X1 U8583 ( .A(n15005), .B(n14553), .ZN(n14493) );
  AND2_X1 U8584 ( .A1(n8082), .A2(n7558), .ZN(n8080) );
  INV_X1 U8585 ( .A(n10326), .ZN(n12545) );
  AND2_X1 U8586 ( .A1(n13516), .A2(n13382), .ZN(n14743) );
  AOI21_X1 U8587 ( .B1(n7502), .B2(n7826), .A(n7828), .ZN(n7823) );
  INV_X1 U8588 ( .A(n14770), .ZN(n7828) );
  OAI21_X1 U8589 ( .B1(n14809), .B2(n7830), .A(n7829), .ZN(n14792) );
  INV_X1 U8590 ( .A(n7824), .ZN(n7829) );
  NAND2_X1 U8591 ( .A1(n14808), .A2(n13475), .ZN(n14793) );
  NAND2_X1 U8592 ( .A1(n14802), .A2(n14791), .ZN(n14785) );
  NAND2_X1 U8593 ( .A1(n14809), .A2(n14810), .ZN(n14808) );
  INV_X1 U8594 ( .A(n14810), .ZN(n7827) );
  AOI21_X1 U8595 ( .B1(n8164), .B2(n13538), .A(n7435), .ZN(n8163) );
  NAND2_X1 U8596 ( .A1(n14892), .A2(n14879), .ZN(n14874) );
  NAND2_X1 U8597 ( .A1(n13537), .A2(n13536), .ZN(n14873) );
  NAND2_X1 U8598 ( .A1(n14913), .A2(n14919), .ZN(n14912) );
  NAND2_X1 U8599 ( .A1(n7974), .A2(n7973), .ZN(n12555) );
  OR2_X1 U8600 ( .A1(n12215), .A2(n12214), .ZN(n12422) );
  NAND2_X1 U8601 ( .A1(n7976), .A2(n7975), .ZN(n12430) );
  INV_X1 U8602 ( .A(n7976), .ZN(n12227) );
  INV_X1 U8603 ( .A(n12118), .ZN(n8032) );
  AOI21_X1 U8604 ( .B1(n12118), .B2(n8031), .A(n8030), .ZN(n8029) );
  INV_X1 U8605 ( .A(n12186), .ZN(n8030) );
  NAND2_X1 U8606 ( .A1(n12027), .A2(n12026), .ZN(n12028) );
  AND2_X1 U8607 ( .A1(n11778), .A2(n16141), .ZN(n11685) );
  NAND2_X1 U8608 ( .A1(n8049), .A2(n11538), .ZN(n11782) );
  NAND2_X1 U8609 ( .A1(n8049), .A2(n8048), .ZN(n11784) );
  NAND2_X1 U8610 ( .A1(n7623), .A2(n11537), .ZN(n11777) );
  INV_X1 U8611 ( .A(n11399), .ZN(n7623) );
  NOR2_X1 U8612 ( .A1(n11777), .A2(n16122), .ZN(n11778) );
  NAND2_X1 U8613 ( .A1(n11391), .A2(n11390), .ZN(n11558) );
  NAND2_X1 U8614 ( .A1(n11211), .A2(n11389), .ZN(n11399) );
  NAND2_X1 U8615 ( .A1(n11040), .A2(n11059), .ZN(n11202) );
  OAI22_X1 U8616 ( .A1(n13622), .A2(n10736), .B1(n7580), .B2(n7432), .ZN(
        n11038) );
  INV_X1 U8617 ( .A(n13623), .ZN(n11037) );
  INV_X1 U8618 ( .A(n14916), .ZN(n14885) );
  NAND2_X1 U8619 ( .A1(n13664), .A2(n13622), .ZN(n10768) );
  NAND2_X1 U8620 ( .A1(n13489), .A2(n13488), .ZN(n14959) );
  NAND2_X1 U8621 ( .A1(n12023), .A2(n12022), .ZN(n13753) );
  INV_X1 U8622 ( .A(n13663), .ZN(n15031) );
  AND2_X1 U8623 ( .A1(n10661), .A2(n15031), .ZN(n14998) );
  AND2_X1 U8624 ( .A1(n8322), .A2(n8043), .ZN(n8321) );
  OAI21_X1 U8625 ( .B1(n10277), .B2(P2_IR_REG_23__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n10098) );
  INV_X1 U8626 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n10097) );
  AND2_X1 U8627 ( .A1(n10411), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n10280) );
  AND2_X1 U8628 ( .A1(n10278), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10279) );
  OR2_X1 U8629 ( .A1(n11771), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n11220) );
  AND2_X1 U8630 ( .A1(n10410), .A2(n10409), .ZN(n10722) );
  INV_X1 U8631 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n10295) );
  INV_X1 U8632 ( .A(n8881), .ZN(n8897) );
  AND2_X1 U8633 ( .A1(n8734), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8721) );
  AND2_X1 U8634 ( .A1(n10878), .A2(n10877), .ZN(n13258) );
  NAND2_X1 U8635 ( .A1(n11275), .A2(n11274), .ZN(n8197) );
  NOR2_X1 U8636 ( .A1(n11823), .A2(n8213), .ZN(n8212) );
  INV_X1 U8637 ( .A(n8358), .ZN(n8213) );
  AOI21_X1 U8638 ( .B1(n13286), .B2(n7665), .A(n7662), .ZN(n7661) );
  NOR2_X1 U8639 ( .A1(n12391), .A2(n8217), .ZN(n8216) );
  INV_X1 U8640 ( .A(n8356), .ZN(n8217) );
  OR2_X1 U8641 ( .A1(n11106), .A2(n13587), .ZN(n10672) );
  INV_X1 U8642 ( .A(n15130), .ZN(n8173) );
  AOI21_X1 U8643 ( .B1(n15130), .B2(n8172), .A(n7499), .ZN(n8171) );
  INV_X1 U8644 ( .A(n13285), .ZN(n8172) );
  AND3_X1 U8645 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n8834) );
  NAND2_X1 U8646 ( .A1(n8195), .A2(n8198), .ZN(n8206) );
  OR2_X1 U8647 ( .A1(n11275), .A2(n8200), .ZN(n8195) );
  NOR2_X1 U8648 ( .A1(n8668), .A2(n15086), .ZN(n8654) );
  INV_X1 U8649 ( .A(n13587), .ZN(n13572) );
  NAND2_X1 U8650 ( .A1(n9090), .A2(n9091), .ZN(n7617) );
  NAND2_X1 U8651 ( .A1(n9088), .A2(n9089), .ZN(n7618) );
  NAND2_X1 U8652 ( .A1(n8925), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n8742) );
  INV_X1 U8653 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10633) );
  NAND2_X1 U8654 ( .A1(n10608), .A2(n10609), .ZN(n10679) );
  NOR2_X1 U8655 ( .A1(n10755), .A2(n7724), .ZN(n10922) );
  AND2_X1 U8656 ( .A1(n10756), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7724) );
  NAND2_X1 U8657 ( .A1(n10922), .A2(n10921), .ZN(n10920) );
  NAND2_X1 U8658 ( .A1(n10920), .A2(n7723), .ZN(n10759) );
  OR2_X1 U8659 ( .A1(n10758), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7723) );
  NAND2_X1 U8660 ( .A1(n10759), .A2(n10760), .ZN(n11174) );
  NOR2_X1 U8661 ( .A1(n11318), .A2(n7718), .ZN(n11321) );
  AND2_X1 U8662 ( .A1(n11319), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7718) );
  NAND2_X1 U8663 ( .A1(n11321), .A2(n11320), .ZN(n11705) );
  NAND2_X1 U8664 ( .A1(n11705), .A2(n7715), .ZN(n11706) );
  NAND2_X1 U8665 ( .A1(n7717), .A2(n7716), .ZN(n7715) );
  XNOR2_X1 U8666 ( .A(n11706), .B(n15779), .ZN(n15775) );
  INV_X1 U8667 ( .A(n15474), .ZN(n13344) );
  AND2_X1 U8668 ( .A1(n8554), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8923) );
  NAND2_X1 U8669 ( .A1(n8057), .A2(n15485), .ZN(n8056) );
  INV_X1 U8670 ( .A(n8058), .ZN(n8057) );
  NAND2_X1 U8671 ( .A1(n15307), .A2(n13339), .ZN(n15303) );
  NOR3_X1 U8672 ( .A1(n15343), .A2(n8058), .A3(n15491), .ZN(n15297) );
  INV_X1 U8673 ( .A(n8254), .ZN(n8253) );
  OAI21_X1 U8674 ( .B1(n8256), .B2(n13338), .A(n8360), .ZN(n8254) );
  NOR2_X1 U8675 ( .A1(n15343), .A2(n8058), .ZN(n15309) );
  NOR2_X1 U8676 ( .A1(n15343), .A2(n15334), .ZN(n15331) );
  INV_X1 U8677 ( .A(n7774), .ZN(n15340) );
  AND2_X1 U8678 ( .A1(n7779), .A2(n15369), .ZN(n7777) );
  NOR2_X1 U8679 ( .A1(n8621), .A2(n8608), .ZN(n8867) );
  AND2_X1 U8680 ( .A1(n8867), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8869) );
  INV_X1 U8681 ( .A(n8059), .ZN(n15438) );
  AND2_X1 U8682 ( .A1(n8013), .A2(n7552), .ZN(n8012) );
  INV_X1 U8683 ( .A(n8060), .ZN(n15453) );
  OR2_X1 U8684 ( .A1(n16244), .A2(n16251), .ZN(n8295) );
  OR2_X1 U8685 ( .A1(n8698), .A2(n12392), .ZN(n8687) );
  OAI22_X1 U8686 ( .A1(n11921), .A2(n8271), .B1(n8272), .B2(n12166), .ZN(
        n12170) );
  NAND2_X1 U8687 ( .A1(n8275), .A2(n12011), .ZN(n8271) );
  AND2_X1 U8688 ( .A1(n12167), .A2(n8273), .ZN(n8272) );
  INV_X1 U8689 ( .A(n8005), .ZN(n8004) );
  OAI21_X1 U8690 ( .B1(n11494), .B2(n8006), .A(n11497), .ZN(n8005) );
  NAND2_X1 U8691 ( .A1(n8052), .A2(n8051), .ZN(n11647) );
  NAND2_X1 U8692 ( .A1(n11299), .A2(n11298), .ZN(n11300) );
  NAND2_X1 U8693 ( .A1(n11108), .A2(n11107), .ZN(n11304) );
  INV_X1 U8694 ( .A(n15455), .ZN(n15406) );
  XNOR2_X1 U8695 ( .A(n7599), .B(n11011), .ZN(n10884) );
  NAND2_X1 U8696 ( .A1(n8284), .A2(n8283), .ZN(n15554) );
  AND2_X1 U8697 ( .A1(n8284), .A2(n7470), .ZN(n15444) );
  NAND2_X1 U8698 ( .A1(n8664), .A2(n8663), .ZN(n16277) );
  NAND2_X1 U8699 ( .A1(n12012), .A2(n12011), .ZN(n12168) );
  NOR2_X2 U8700 ( .A1(n16031), .A2(n8224), .ZN(n16247) );
  INV_X1 U8701 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n8790) );
  NAND2_X1 U8702 ( .A1(n7581), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8379) );
  XNOR2_X1 U8703 ( .A(n8537), .B(n8536), .ZN(n15063) );
  XNOR2_X1 U8704 ( .A(n8550), .B(n8549), .ZN(n15067) );
  NAND2_X1 U8705 ( .A1(n8464), .A2(n8463), .ZN(n8887) );
  AND2_X1 U8706 ( .A1(n8261), .A2(n8461), .ZN(n8260) );
  XNOR2_X1 U8707 ( .A(n8887), .B(n9621), .ZN(n8890) );
  AND2_X1 U8708 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n8509) );
  INV_X1 U8709 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n7897) );
  NAND2_X1 U8710 ( .A1(n7832), .A2(n8450), .ZN(n8601) );
  NAND2_X1 U8711 ( .A1(n8812), .A2(n8413), .ZN(n7822) );
  NAND2_X1 U8712 ( .A1(n8404), .A2(n8403), .ZN(n8756) );
  NAND2_X1 U8713 ( .A1(n10431), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8026) );
  XNOR2_X1 U8714 ( .A(n15814), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n15819) );
  AOI21_X1 U8715 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n16028), .A(n15859), .ZN(
        n15866) );
  NAND2_X1 U8716 ( .A1(n12398), .A2(n9795), .ZN(n10254) );
  NAND2_X1 U8717 ( .A1(n11328), .A2(n9774), .ZN(n8117) );
  AND2_X1 U8718 ( .A1(n8120), .A2(n7526), .ZN(n8119) );
  NAND2_X1 U8719 ( .A1(n7436), .A2(n7461), .ZN(n8124) );
  NAND2_X1 U8720 ( .A1(n12047), .A2(n9789), .ZN(n12259) );
  AND2_X1 U8721 ( .A1(n12639), .A2(n9808), .ZN(n13195) );
  NAND2_X1 U8722 ( .A1(n12257), .A2(n9792), .ZN(n12400) );
  INV_X1 U8723 ( .A(n14032), .ZN(n16039) );
  NOR2_X1 U8724 ( .A1(n13225), .A2(n7866), .ZN(n7865) );
  INV_X1 U8725 ( .A(n9810), .ZN(n7866) );
  NAND2_X1 U8726 ( .A1(n13194), .A2(n9810), .ZN(n13226) );
  AND4_X1 U8727 ( .A1(n9469), .A2(n9468), .A3(n9467), .A4(n9466), .ZN(n13230)
         );
  NAND2_X1 U8728 ( .A1(n12641), .A2(n12640), .ZN(n12639) );
  XNOR2_X1 U8729 ( .A(n9773), .B(n14058), .ZN(n11330) );
  NAND2_X1 U8730 ( .A1(n7654), .A2(n7653), .ZN(n11944) );
  INV_X1 U8731 ( .A(n11942), .ZN(n7653) );
  OAI211_X1 U8732 ( .C1(n9908), .C2(n9593), .A(n9592), .B(n9591), .ZN(n14305)
         );
  INV_X1 U8733 ( .A(n14316), .ZN(n14290) );
  INV_X1 U8734 ( .A(n13230), .ZN(n14050) );
  INV_X1 U8735 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n15967) );
  NAND2_X1 U8736 ( .A1(n10856), .A2(n10144), .ZN(n11155) );
  INV_X1 U8737 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n15989) );
  INV_X1 U8738 ( .A(n7912), .ZN(n11380) );
  INV_X1 U8739 ( .A(n7902), .ZN(n11621) );
  INV_X1 U8740 ( .A(n7986), .ZN(n11618) );
  INV_X1 U8741 ( .A(n7981), .ZN(n12140) );
  NOR2_X1 U8742 ( .A1(n12154), .A2(n10156), .ZN(n12130) );
  NOR2_X1 U8743 ( .A1(n9479), .A2(n14061), .ZN(n14060) );
  NOR2_X1 U8744 ( .A1(n12134), .A2(n10209), .ZN(n14064) );
  XNOR2_X1 U8745 ( .A(n14128), .B(n14129), .ZN(n14097) );
  INV_X1 U8746 ( .A(n14130), .ZN(n7916) );
  XNOR2_X1 U8747 ( .A(n7998), .B(n14149), .ZN(n7997) );
  NAND2_X1 U8748 ( .A1(n8000), .A2(n7999), .ZN(n7998) );
  NAND2_X1 U8749 ( .A1(n14148), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n7999) );
  NAND2_X1 U8750 ( .A1(n14153), .A2(n16017), .ZN(n7996) );
  NAND2_X1 U8751 ( .A1(n14150), .A2(n14151), .ZN(n7995) );
  XNOR2_X1 U8752 ( .A(n9923), .B(n7471), .ZN(n14168) );
  NAND2_X1 U8753 ( .A1(n8338), .A2(n8343), .ZN(n14200) );
  NAND2_X1 U8754 ( .A1(n14217), .A2(n8344), .ZN(n8338) );
  NOR2_X1 U8755 ( .A1(n14219), .A2(n9936), .ZN(n14205) );
  NAND2_X1 U8756 ( .A1(n8349), .A2(n10030), .ZN(n14248) );
  NAND2_X1 U8757 ( .A1(n9623), .A2(n9622), .ZN(n14377) );
  AND3_X1 U8758 ( .A1(n9605), .A2(n9604), .A3(n9603), .ZN(n14268) );
  NAND2_X1 U8759 ( .A1(n14308), .A2(n10020), .ZN(n14294) );
  NAND2_X1 U8760 ( .A1(n9525), .A2(n9524), .ZN(n14328) );
  OAI21_X1 U8761 ( .B1(n13175), .B2(n9999), .A(n7690), .ZN(n13212) );
  NAND2_X1 U8762 ( .A1(n7689), .A2(n9998), .ZN(n13214) );
  NAND2_X1 U8763 ( .A1(n13175), .A2(n7439), .ZN(n7689) );
  NAND2_X1 U8764 ( .A1(n13175), .A2(n9989), .ZN(n13189) );
  NAND2_X1 U8765 ( .A1(n7948), .A2(n9799), .ZN(n12599) );
  NAND2_X1 U8766 ( .A1(n12286), .A2(n9977), .ZN(n12326) );
  NAND2_X1 U8767 ( .A1(n11959), .A2(n9730), .ZN(n12284) );
  AND2_X1 U8768 ( .A1(n11573), .A2(n9339), .ZN(n11805) );
  INV_X1 U8769 ( .A(n16094), .ZN(n16059) );
  OR3_X1 U8770 ( .A1(n10401), .A2(n16061), .A3(n16231), .ZN(n14337) );
  AND2_X1 U8771 ( .A1(n10395), .A2(n10394), .ZN(n16094) );
  AND3_X1 U8772 ( .A1(n9419), .A2(n9418), .A3(n9417), .ZN(n12440) );
  INV_X1 U8773 ( .A(n9924), .ZN(n14428) );
  OR2_X1 U8774 ( .A1(n14376), .A2(n14375), .ZN(n14437) );
  NAND2_X1 U8775 ( .A1(n9550), .A2(n9549), .ZN(n14455) );
  NAND2_X1 U8776 ( .A1(n9517), .A2(n9516), .ZN(n14463) );
  INV_X1 U8777 ( .A(n12440), .ZN(n12444) );
  AND3_X1 U8778 ( .A1(n9404), .A2(n9403), .A3(n9402), .ZN(n12075) );
  INV_X1 U8779 ( .A(n16038), .ZN(n11481) );
  NAND2_X1 U8780 ( .A1(n16242), .A2(n16102), .ZN(n14464) );
  AND2_X1 U8781 ( .A1(n10128), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14467) );
  INV_X1 U8782 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n14470) );
  NAND2_X1 U8783 ( .A1(n7871), .A2(n7868), .ZN(n12463) );
  NOR2_X1 U8784 ( .A1(n7870), .A2(n7869), .ZN(n7868) );
  NAND2_X1 U8785 ( .A1(n9225), .A2(n7500), .ZN(n7871) );
  NOR2_X1 U8786 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_26__SCAN_IN), .ZN(
        n7869) );
  NAND2_X1 U8787 ( .A1(n9223), .A2(n9225), .ZN(n12378) );
  MUX2_X1 U8788 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9221), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n9223) );
  NAND2_X1 U8789 ( .A1(n8138), .A2(n9247), .ZN(n8137) );
  NAND2_X1 U8790 ( .A1(n7754), .A2(n9179), .ZN(n9608) );
  NAND2_X1 U8791 ( .A1(n9177), .A2(n7758), .ZN(n7754) );
  XNOR2_X1 U8792 ( .A(n9257), .B(n9256), .ZN(n11614) );
  NAND2_X1 U8793 ( .A1(n9177), .A2(n9176), .ZN(n9598) );
  INV_X1 U8794 ( .A(SI_19_), .ZN(n12956) );
  INV_X1 U8795 ( .A(SI_18_), .ZN(n12736) );
  INV_X1 U8796 ( .A(SI_16_), .ZN(n11069) );
  INV_X1 U8797 ( .A(SI_15_), .ZN(n10936) );
  NAND2_X1 U8798 ( .A1(n9473), .A2(n9164), .ZN(n9488) );
  NAND2_X1 U8799 ( .A1(n9495), .A2(n9494), .ZN(n10729) );
  INV_X1 U8800 ( .A(SI_11_), .ZN(n12973) );
  INV_X1 U8801 ( .A(n10155), .ZN(n12153) );
  OAI21_X1 U8802 ( .B1(n9414), .B2(n7742), .A(n7740), .ZN(n9433) );
  NAND2_X1 U8803 ( .A1(n7739), .A2(n9155), .ZN(n9431) );
  OAI21_X1 U8804 ( .B1(n9144), .B2(n7770), .A(n7769), .ZN(n9388) );
  NAND2_X1 U8805 ( .A1(n9354), .A2(n9145), .ZN(n9372) );
  NAND2_X1 U8806 ( .A1(n7746), .A2(n9139), .ZN(n9333) );
  NAND2_X1 U8807 ( .A1(n7747), .A2(n7748), .ZN(n9318) );
  INV_X1 U8808 ( .A(n9137), .ZN(n9284) );
  INV_X1 U8809 ( .A(n10140), .ZN(n9288) );
  NAND2_X1 U8810 ( .A1(n7910), .A2(n9330), .ZN(n7909) );
  AND2_X1 U8811 ( .A1(n13243), .A2(n10103), .ZN(n10538) );
  NOR2_X1 U8812 ( .A1(n11603), .A2(n11604), .ZN(n11743) );
  NAND2_X1 U8813 ( .A1(n8106), .A2(n8110), .ZN(n12584) );
  NAND2_X1 U8814 ( .A1(n8103), .A2(n8107), .ZN(n12611) );
  NAND2_X1 U8815 ( .A1(n12476), .A2(n8111), .ZN(n8106) );
  NAND2_X1 U8816 ( .A1(n8069), .A2(n10320), .ZN(n8068) );
  OAI21_X1 U8817 ( .B1(n14595), .B2(n8099), .A(n8098), .ZN(n14542) );
  NAND2_X1 U8818 ( .A1(n11603), .A2(n8092), .ZN(n8087) );
  NAND2_X1 U8819 ( .A1(n11194), .A2(n11193), .ZN(n11192) );
  INV_X1 U8820 ( .A(n14684), .ZN(n11911) );
  OAI21_X1 U8821 ( .B1(n11603), .B2(n8089), .A(n8088), .ZN(n11907) );
  NAND2_X1 U8822 ( .A1(n8113), .A2(n12474), .ZN(n12583) );
  OR2_X1 U8823 ( .A1(n12476), .A2(n12475), .ZN(n8113) );
  NOR2_X1 U8824 ( .A1(n10373), .A2(n14916), .ZN(n14627) );
  NOR2_X1 U8825 ( .A1(n14593), .A2(n14491), .ZN(n14636) );
  AND2_X1 U8826 ( .A1(n8080), .A2(n8081), .ZN(n14646) );
  AND2_X1 U8827 ( .A1(n13501), .A2(n13491), .ZN(n14777) );
  AOI21_X1 U8828 ( .B1(n10364), .B2(n11364), .A(n14929), .ZN(n14670) );
  INV_X1 U8829 ( .A(n14677), .ZN(n13776) );
  NAND2_X1 U8830 ( .A1(n10372), .A2(n14883), .ZN(n14661) );
  INV_X1 U8831 ( .A(n14667), .ZN(n14638) );
  AOI21_X1 U8832 ( .B1(n8107), .B2(n8109), .A(n12610), .ZN(n8104) );
  INV_X1 U8833 ( .A(n14670), .ZN(n14651) );
  OR2_X1 U8834 ( .A1(n10360), .A2(n10359), .ZN(n14642) );
  INV_X1 U8835 ( .A(n13869), .ZN(n14740) );
  INV_X1 U8836 ( .A(n14752), .ZN(n14672) );
  NAND2_X1 U8837 ( .A1(n13510), .A2(n13509), .ZN(n14774) );
  OR2_X1 U8838 ( .A1(n14760), .A2(n13504), .ZN(n13510) );
  NAND2_X1 U8839 ( .A1(n13486), .A2(n13485), .ZN(n14811) );
  OR2_X1 U8840 ( .A1(n14788), .A2(n13504), .ZN(n13486) );
  NAND2_X1 U8841 ( .A1(n13473), .A2(n13472), .ZN(n14819) );
  NAND2_X1 U8842 ( .A1(n13397), .A2(n13396), .ZN(n14837) );
  NAND2_X1 U8843 ( .A1(n13458), .A2(n13457), .ZN(n14858) );
  NAND2_X1 U8844 ( .A1(n13430), .A2(n13429), .ZN(n14857) );
  CLKBUF_X1 U8845 ( .A(n14691), .Z(n7580) );
  INV_X1 U8846 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8393) );
  NAND2_X1 U8847 ( .A1(n7965), .A2(n15027), .ZN(n14939) );
  XNOR2_X1 U8848 ( .A(n14728), .B(n7966), .ZN(n7965) );
  NAND2_X1 U8849 ( .A1(n7629), .A2(n12551), .ZN(n12552) );
  NAND2_X1 U8851 ( .A1(n12522), .A2(n12521), .ZN(n12523) );
  NAND2_X1 U8852 ( .A1(n12416), .A2(n12415), .ZN(n15025) );
  NAND2_X1 U8853 ( .A1(n12119), .A2(n12118), .ZN(n12187) );
  NAND2_X1 U8854 ( .A1(n16188), .A2(n11870), .ZN(n11889) );
  NAND2_X1 U8855 ( .A1(n8158), .A2(n13633), .ZN(n16188) );
  INV_X1 U8856 ( .A(n11692), .ZN(n8158) );
  NAND2_X1 U8857 ( .A1(n14939), .A2(n7963), .ZN(n15034) );
  INV_X1 U8858 ( .A(n7964), .ZN(n7963) );
  OAI21_X1 U8859 ( .B1(n7966), .B2(n16307), .A(n14940), .ZN(n7964) );
  OAI211_X1 U8860 ( .C1(n15031), .C2(n14958), .A(n14957), .B(n14956), .ZN(
        n15038) );
  OR3_X1 U8861 ( .A1(n14985), .A2(n14984), .A3(n14983), .ZN(n15043) );
  OR2_X1 U8862 ( .A1(n14992), .A2(n14991), .ZN(n15044) );
  INV_X1 U8863 ( .A(n8365), .ZN(n7970) );
  XNOR2_X1 U8864 ( .A(n10101), .B(P2_IR_REG_26__SCAN_IN), .ZN(n15066) );
  NAND2_X1 U8865 ( .A1(n10100), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10101) );
  XNOR2_X1 U8866 ( .A(n10102), .B(P2_IR_REG_25__SCAN_IN), .ZN(n15071) );
  XNOR2_X1 U8867 ( .A(n10098), .B(n10097), .ZN(n13240) );
  XNOR2_X1 U8868 ( .A(n8890), .B(n8889), .ZN(n13446) );
  INV_X1 U8869 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n10288) );
  INV_X1 U8870 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n10287) );
  INV_X1 U8871 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11775) );
  INV_X1 U8872 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11294) );
  INV_X1 U8873 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10653) );
  INV_X1 U8874 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10501) );
  INV_X1 U8875 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10461) );
  INV_X1 U8876 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10449) );
  INV_X1 U8877 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10418) );
  INV_X1 U8878 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n11044) );
  INV_X1 U8879 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10408) );
  NAND2_X1 U8880 ( .A1(n13264), .A2(n8359), .ZN(n15084) );
  NAND2_X1 U8881 ( .A1(n8652), .A2(n8651), .ZN(n15089) );
  INV_X1 U8882 ( .A(n15185), .ZN(n12489) );
  OAI21_X1 U8883 ( .B1(n13286), .B2(n7458), .A(n7665), .ZN(n15105) );
  NAND2_X1 U8884 ( .A1(n8186), .A2(n8182), .ZN(n8175) );
  NAND2_X1 U8885 ( .A1(n8182), .A2(n8178), .ZN(n8177) );
  NAND2_X1 U8886 ( .A1(n11821), .A2(n8358), .ZN(n11822) );
  NOR2_X1 U8887 ( .A1(n10579), .A2(n10580), .ZN(n10668) );
  NAND2_X1 U8888 ( .A1(n15147), .A2(n13310), .ZN(n15114) );
  NAND2_X1 U8889 ( .A1(n8218), .A2(n8215), .ZN(n12678) );
  AND2_X1 U8890 ( .A1(n12570), .A2(n7443), .ZN(n8215) );
  AND2_X1 U8891 ( .A1(n8218), .A2(n7443), .ZN(n12571) );
  NAND2_X1 U8892 ( .A1(n16318), .A2(n7659), .ZN(n16347) );
  NAND2_X1 U8893 ( .A1(n13278), .A2(n7660), .ZN(n7659) );
  INV_X1 U8894 ( .A(n13279), .ZN(n7660) );
  NAND2_X1 U8895 ( .A1(n8214), .A2(n8211), .ZN(n12268) );
  AND2_X1 U8896 ( .A1(n11983), .A2(n7442), .ZN(n8211) );
  AND2_X1 U8897 ( .A1(n8214), .A2(n7442), .ZN(n11984) );
  NAND2_X1 U8898 ( .A1(n12686), .A2(n12685), .ZN(n13264) );
  NAND2_X1 U8899 ( .A1(n15607), .A2(n10455), .ZN(n15516) );
  NAND2_X1 U8900 ( .A1(n15112), .A2(n7490), .ZN(n13555) );
  NAND2_X1 U8901 ( .A1(n15112), .A2(n13315), .ZN(n13317) );
  NAND2_X1 U8902 ( .A1(n12389), .A2(n8356), .ZN(n12390) );
  INV_X1 U8903 ( .A(n7658), .ZN(n10949) );
  OAI21_X1 U8904 ( .B1(n13286), .B2(n8173), .A(n8171), .ZN(n15156) );
  NAND2_X1 U8905 ( .A1(n8193), .A2(n8192), .ZN(n11656) );
  AND2_X1 U8906 ( .A1(n8196), .A2(n8203), .ZN(n8192) );
  INV_X1 U8907 ( .A(n8204), .ZN(n8203) );
  NAND2_X1 U8908 ( .A1(n8202), .A2(n11463), .ZN(n11469) );
  NAND2_X1 U8909 ( .A1(n8206), .A2(n7569), .ZN(n8202) );
  XNOR2_X1 U8910 ( .A(n13278), .B(n13279), .ZN(n16319) );
  OAI21_X1 U8911 ( .B1(n15390), .B2(n8872), .A(n8599), .ZN(n15375) );
  OAI21_X1 U8912 ( .B1(n15410), .B2(n8872), .A(n8857), .ZN(n15421) );
  OR2_X1 U8913 ( .A1(n10454), .A2(P1_U3086), .ZN(n10104) );
  INV_X1 U8914 ( .A(n7726), .ZN(n10780) );
  NAND2_X1 U8915 ( .A1(n10623), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7725) );
  INV_X1 U8916 ( .A(n7709), .ZN(n10789) );
  NAND2_X1 U8917 ( .A1(n10687), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7708) );
  AND2_X1 U8918 ( .A1(n11709), .A2(n11708), .ZN(n12080) );
  NAND2_X1 U8919 ( .A1(n15761), .A2(n7468), .ZN(n12623) );
  INV_X1 U8920 ( .A(n7713), .ZN(n15215) );
  INV_X1 U8921 ( .A(n7711), .ZN(n15228) );
  INV_X1 U8922 ( .A(n15257), .ZN(n15472) );
  NAND2_X1 U8923 ( .A1(n8007), .A2(n8009), .ZN(n15477) );
  OR2_X1 U8924 ( .A1(n15325), .A2(n8256), .ZN(n15320) );
  NAND2_X1 U8925 ( .A1(n7778), .A2(n7779), .ZN(n15370) );
  OR2_X1 U8926 ( .A1(n15400), .A2(n7780), .ZN(n7778) );
  NAND2_X1 U8927 ( .A1(n7781), .A2(n7434), .ZN(n15395) );
  AND2_X1 U8928 ( .A1(n7781), .A2(n7783), .ZN(n15394) );
  NAND2_X1 U8929 ( .A1(n15400), .A2(n13335), .ZN(n7781) );
  OAI21_X1 U8930 ( .B1(n15450), .B2(n8282), .A(n8280), .ZN(n15420) );
  NAND2_X1 U8931 ( .A1(n13356), .A2(n13355), .ZN(n15460) );
  AND2_X1 U8932 ( .A1(n8289), .A2(n8288), .ZN(n16301) );
  NOR2_X1 U8933 ( .A1(n8291), .A2(n12697), .ZN(n8288) );
  NAND2_X1 U8934 ( .A1(n8289), .A2(n8290), .ZN(n12660) );
  NAND2_X1 U8935 ( .A1(n16250), .A2(n12487), .ZN(n12649) );
  NAND2_X1 U8936 ( .A1(n8676), .A2(n8675), .ZN(n16266) );
  NAND2_X1 U8937 ( .A1(n16154), .A2(n11929), .ZN(n12005) );
  NAND2_X1 U8938 ( .A1(n8296), .A2(n11918), .ZN(n16150) );
  OR2_X1 U8939 ( .A1(n16275), .A2(n11296), .ZN(n15466) );
  INV_X1 U8940 ( .A(n7787), .ZN(n7784) );
  NAND2_X1 U8941 ( .A1(n11495), .A2(n11494), .ZN(n11641) );
  INV_X1 U8942 ( .A(n15466), .ZN(n15366) );
  NAND2_X1 U8943 ( .A1(n7599), .A2(n10874), .ZN(n10875) );
  OR2_X1 U8944 ( .A1(n16275), .A2(n11079), .ZN(n15416) );
  NAND2_X1 U8945 ( .A1(n10524), .A2(n10523), .ZN(n16110) );
  INV_X1 U8946 ( .A(n16114), .ZN(n16265) );
  INV_X1 U8947 ( .A(n15416), .ZN(n16073) );
  AND2_X1 U8948 ( .A1(n8008), .A2(n8009), .ZN(n7792) );
  AOI21_X1 U8949 ( .B1(n15482), .B2(n16337), .A(n15481), .ZN(n15484) );
  NAND2_X1 U8950 ( .A1(n7441), .A2(n7474), .ZN(n15588) );
  INV_X1 U8951 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7791) );
  AND3_X1 U8952 ( .A1(n8187), .A2(n8603), .A3(n8500), .ZN(n8054) );
  AND2_X1 U8953 ( .A1(n8378), .A2(n9107), .ZN(n7632) );
  INV_X1 U8954 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9110) );
  NAND2_X1 U8955 ( .A1(n9102), .A2(n9101), .ZN(n9104) );
  NAND2_X1 U8956 ( .A1(n9100), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9101) );
  AND2_X1 U8957 ( .A1(n10432), .A2(P1_U3086), .ZN(n15601) );
  XNOR2_X1 U8958 ( .A(n8570), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15607) );
  NAND2_X1 U8959 ( .A1(n8890), .A2(n10420), .ZN(n8570) );
  INV_X1 U8960 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n13252) );
  INV_X1 U8961 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n11737) );
  INV_X1 U8962 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n11289) );
  INV_X1 U8963 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n11226) );
  INV_X1 U8964 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10727) );
  INV_X1 U8965 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10503) );
  INV_X1 U8966 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10496) );
  INV_X1 U8967 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10483) );
  INV_X1 U8968 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10463) );
  INV_X1 U8969 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10451) );
  INV_X1 U8970 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10423) );
  INV_X1 U8971 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10428) );
  NAND2_X1 U8972 ( .A1(n8775), .A2(n7720), .ZN(n10618) );
  INV_X1 U8973 ( .A(n7721), .ZN(n7720) );
  OAI21_X1 U8974 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(P1_IR_REG_1__SCAN_IN), .A(
        n7722), .ZN(n7721) );
  INV_X1 U8975 ( .A(P1_RD_REG_SCAN_IN), .ZN(n16030) );
  INV_X1 U8976 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7624) );
  XNOR2_X1 U8977 ( .A(n15819), .B(n7927), .ZN(n15818) );
  NOR2_X1 U8978 ( .A1(n15832), .A2(n15831), .ZN(n15955) );
  XNOR2_X1 U8979 ( .A(n15836), .B(n7931), .ZN(n15838) );
  NAND2_X1 U8980 ( .A1(n15850), .A2(n15849), .ZN(n15860) );
  NAND2_X1 U8981 ( .A1(n15862), .A2(n7584), .ZN(n15869) );
  OAI21_X1 U8982 ( .B1(n15860), .B2(n15861), .A(P2_ADDR_REG_9__SCAN_IN), .ZN(
        n7584) );
  NOR2_X1 U8983 ( .A1(n15927), .A2(n15928), .ZN(n15935) );
  INV_X1 U8984 ( .A(n15944), .ZN(n7923) );
  OAI211_X1 U8985 ( .C1(n13989), .C2(n7851), .A(n7850), .B(n7847), .ZN(n13933)
         );
  NAND2_X1 U8986 ( .A1(n11413), .A2(n9778), .ZN(n11723) );
  OAI21_X1 U8987 ( .B1(n7595), .B2(n14041), .A(n14027), .ZN(P3_U3180) );
  XNOR2_X1 U8988 ( .A(n14022), .B(n7559), .ZN(n7595) );
  NAND2_X1 U8989 ( .A1(n7705), .A2(n10127), .ZN(n7728) );
  OR4_X1 U8990 ( .A1(n10251), .A2(n10250), .A3(n10249), .A4(n10248), .ZN(
        P3_U3198) );
  OAI21_X1 U8991 ( .B1(n7917), .B2(n7916), .A(n14136), .ZN(n7915) );
  INV_X1 U8992 ( .A(n7640), .ZN(n14181) );
  AOI21_X1 U8993 ( .B1(n14347), .B2(n16096), .A(n14180), .ZN(n7641) );
  NAND2_X1 U8994 ( .A1(n8337), .A2(n16238), .ZN(n9765) );
  AND2_X1 U8995 ( .A1(n9270), .A2(n9269), .ZN(n9747) );
  NAND2_X1 U8996 ( .A1(n8337), .A2(n16242), .ZN(n9746) );
  NAND2_X1 U8997 ( .A1(n8081), .A2(n8082), .ZN(n11596) );
  INV_X1 U8998 ( .A(n13919), .ZN(n8316) );
  OAI211_X1 U8999 ( .C1(n14947), .C2(n14891), .A(n8160), .B(n8159), .ZN(
        P2_U3236) );
  AOI21_X1 U9000 ( .B1(n14943), .B2(n14832), .A(n13551), .ZN(n8159) );
  NAND2_X1 U9001 ( .A1(n8161), .A2(n14843), .ZN(n8160) );
  OR2_X1 U9002 ( .A1(n14749), .A2(n14933), .ZN(n7635) );
  NOR2_X1 U9003 ( .A1(n14967), .A2(n14938), .ZN(n14797) );
  MUX2_X1 U9004 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n15036), .S(n16293), .Z(
        P2_U3528) );
  INV_X1 U9005 ( .A(n7960), .ZN(P2_U3498) );
  AOI21_X1 U9006 ( .B1(n15034), .B2(n7419), .A(n7961), .ZN(n7960) );
  NOR2_X1 U9007 ( .A1(n7419), .A2(n7962), .ZN(n7961) );
  INV_X1 U9008 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n7962) );
  NAND2_X1 U9009 ( .A1(n16315), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n7834) );
  NAND2_X1 U9010 ( .A1(n7677), .A2(n16356), .ZN(n7676) );
  INV_X1 U9011 ( .A(n7585), .ZN(n15880) );
  AND2_X1 U9012 ( .A1(n11957), .A2(n9391), .ZN(n7433) );
  NOR2_X2 U9013 ( .A1(n13336), .A2(n7782), .ZN(n7434) );
  AND2_X1 U9014 ( .A1(n8169), .A2(n8168), .ZN(n7435) );
  NAND2_X1 U9015 ( .A1(n8879), .A2(n8878), .ZN(n15334) );
  XOR2_X1 U9016 ( .A(n14176), .B(n9863), .Z(n7436) );
  OR3_X2 U9017 ( .A1(n15343), .A2(n15491), .A3(n8056), .ZN(n7437) );
  OR2_X1 U9018 ( .A1(n15385), .A2(n15396), .ZN(n7438) );
  AND2_X1 U9019 ( .A1(n9734), .A2(n9989), .ZN(n7439) );
  CLKBUF_X3 U9020 ( .A(n13716), .Z(n13857) );
  NAND2_X1 U9021 ( .A1(n13663), .A2(n13662), .ZN(n13677) );
  XOR2_X1 U9022 ( .A(n10077), .B(n14145), .Z(n7440) );
  INV_X1 U9023 ( .A(n14250), .ZN(n7950) );
  INV_X1 U9024 ( .A(n11842), .ZN(n7939) );
  AND4_X1 U9025 ( .A1(n8378), .A2(n9107), .A3(n8188), .A4(n7791), .ZN(n7441)
         );
  NAND2_X1 U9026 ( .A1(n11977), .A2(n11976), .ZN(n7442) );
  NAND2_X1 U9027 ( .A1(n12566), .A2(n12565), .ZN(n7443) );
  NAND2_X1 U9028 ( .A1(n9661), .A2(n9660), .ZN(n14361) );
  INV_X1 U9029 ( .A(n14361), .ZN(n8347) );
  INV_X1 U9030 ( .A(n9022), .ZN(n7890) );
  AND2_X1 U9031 ( .A1(n7678), .A2(n7496), .ZN(n7444) );
  AND2_X1 U9032 ( .A1(n13762), .A2(n13761), .ZN(n7445) );
  OR2_X1 U9033 ( .A1(n15334), .A2(n15311), .ZN(n7446) );
  AND3_X1 U9034 ( .A1(n7729), .A2(n7731), .A3(n7733), .ZN(n7447) );
  AND2_X1 U9035 ( .A1(n7748), .A2(n7495), .ZN(n7448) );
  AND2_X1 U9036 ( .A1(n8347), .A2(n8346), .ZN(n7449) );
  AND2_X1 U9037 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n7773), .ZN(n7450) );
  AND2_X1 U9038 ( .A1(n13728), .A2(n13727), .ZN(n7451) );
  AND2_X1 U9039 ( .A1(n8084), .A2(n11193), .ZN(n7452) );
  INV_X1 U9040 ( .A(n12527), .ZN(n8224) );
  NAND2_X1 U9041 ( .A1(n8386), .A2(n8504), .ZN(n12527) );
  AND2_X1 U9042 ( .A1(n7520), .A2(n10095), .ZN(n7453) );
  INV_X1 U9043 ( .A(n9029), .ZN(n8227) );
  NAND2_X1 U9044 ( .A1(n8120), .A2(n8124), .ZN(n7454) );
  INV_X1 U9045 ( .A(n15311), .ZN(n8259) );
  INV_X1 U9046 ( .A(n14987), .ZN(n8169) );
  NAND2_X1 U9047 ( .A1(n11841), .A2(n7433), .ZN(n11956) );
  AND2_X1 U9048 ( .A1(n11275), .A2(n8207), .ZN(n7455) );
  AND2_X1 U9049 ( .A1(n14106), .A2(n7984), .ZN(n7456) );
  INV_X1 U9050 ( .A(n11587), .ZN(n8051) );
  NAND2_X1 U9051 ( .A1(n15598), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n7457) );
  NAND2_X1 U9052 ( .A1(n15157), .A2(n8170), .ZN(n7458) );
  NOR2_X1 U9053 ( .A1(n15461), .A2(n8016), .ZN(n7459) );
  INV_X2 U9054 ( .A(n9801), .ZN(n9849) );
  NOR2_X1 U9055 ( .A1(n9406), .A2(n9393), .ZN(n7460) );
  INV_X1 U9056 ( .A(n13928), .ZN(n7861) );
  INV_X1 U9057 ( .A(n13653), .ZN(n7600) );
  AND3_X1 U9058 ( .A1(n9099), .A2(n8516), .A3(n8515), .ZN(n15606) );
  AND2_X1 U9059 ( .A1(n7559), .A2(n13928), .ZN(n7461) );
  XNOR2_X1 U9060 ( .A(n14954), .B(n14774), .ZN(n14753) );
  INV_X1 U9061 ( .A(n15186), .ZN(n12271) );
  AND2_X1 U9062 ( .A1(n13769), .A2(n13768), .ZN(n7462) );
  AND2_X1 U9063 ( .A1(n13796), .A2(n13795), .ZN(n7463) );
  NOR2_X1 U9064 ( .A1(n11906), .A2(n11905), .ZN(n7464) );
  OR2_X1 U9065 ( .A1(n16019), .A2(n10117), .ZN(n7465) );
  INV_X1 U9066 ( .A(n15652), .ZN(n8023) );
  NOR2_X1 U9067 ( .A1(n12648), .A2(n8020), .ZN(n7466) );
  OR2_X1 U9068 ( .A1(n14785), .A2(n7968), .ZN(n7467) );
  NAND2_X1 U9069 ( .A1(n13286), .A2(n13285), .ZN(n15129) );
  OR2_X1 U9070 ( .A1(n12621), .A2(n12627), .ZN(n7468) );
  INV_X1 U9071 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n9211) );
  NAND2_X1 U9072 ( .A1(n13608), .A2(n13607), .ZN(n14725) );
  INV_X1 U9073 ( .A(n14725), .ZN(n7966) );
  INV_X1 U9074 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8322) );
  NAND2_X1 U9075 ( .A1(n8616), .A2(n8615), .ZN(n15454) );
  INV_X1 U9076 ( .A(n15454), .ZN(n16354) );
  AND2_X1 U9077 ( .A1(n10063), .A2(n9730), .ZN(n7469) );
  NAND4_X1 U9078 ( .A1(n8188), .A2(n8187), .A3(n7896), .A4(n9107), .ZN(n8510)
         );
  INV_X1 U9079 ( .A(n11463), .ZN(n8205) );
  INV_X1 U9080 ( .A(n9032), .ZN(n7875) );
  NAND2_X1 U9081 ( .A1(n16354), .A2(n13357), .ZN(n7470) );
  AND2_X1 U9082 ( .A1(n10046), .A2(n10044), .ZN(n7471) );
  AND2_X1 U9083 ( .A1(n16122), .A2(n11556), .ZN(n7472) );
  INV_X1 U9084 ( .A(n13598), .ZN(n8186) );
  NOR2_X1 U9085 ( .A1(n14236), .A2(n7952), .ZN(n7951) );
  OR2_X1 U9086 ( .A1(n16224), .A2(n12489), .ZN(n7473) );
  AND3_X1 U9087 ( .A1(n8187), .A2(n8299), .A3(n8603), .ZN(n7474) );
  OR2_X1 U9088 ( .A1(n15511), .A2(n15180), .ZN(n7475) );
  NOR2_X1 U9089 ( .A1(n13338), .A2(n8298), .ZN(n7476) );
  AND2_X1 U9090 ( .A1(n10044), .A2(n9940), .ZN(n7478) );
  INV_X1 U9091 ( .A(n12010), .ZN(n16197) );
  NAND2_X1 U9092 ( .A1(n8710), .A2(n8709), .ZN(n12010) );
  AND2_X1 U9093 ( .A1(n13786), .A2(n13785), .ZN(n7479) );
  AND3_X1 U9094 ( .A1(n7478), .A2(n9941), .A3(n10046), .ZN(n7480) );
  AND2_X1 U9095 ( .A1(n13773), .A2(n13772), .ZN(n7481) );
  AND2_X1 U9096 ( .A1(n13836), .A2(n13835), .ZN(n7482) );
  NOR2_X1 U9097 ( .A1(n12401), .A2(n8129), .ZN(n7483) );
  OR2_X1 U9098 ( .A1(n15193), .A2(n16077), .ZN(n7484) );
  OR2_X1 U9099 ( .A1(n9917), .A2(SI_2_), .ZN(n7485) );
  XNOR2_X1 U9100 ( .A(n13344), .B(n15179), .ZN(n13368) );
  INV_X1 U9101 ( .A(n7771), .ZN(n7770) );
  NOR2_X1 U9102 ( .A1(n9146), .A2(n7772), .ZN(n7771) );
  AND2_X1 U9103 ( .A1(n10410), .A2(n8078), .ZN(n7486) );
  AND2_X1 U9104 ( .A1(n9049), .A2(n9048), .ZN(n7487) );
  INV_X1 U9105 ( .A(n8208), .ZN(n8207) );
  INV_X1 U9106 ( .A(n9078), .ZN(n8234) );
  AND2_X1 U9107 ( .A1(n7855), .A2(n13928), .ZN(n7488) );
  AND2_X1 U9108 ( .A1(n14107), .A2(n14106), .ZN(n7489) );
  AND2_X1 U9109 ( .A1(n13319), .A2(n13315), .ZN(n7490) );
  AND4_X1 U9110 ( .A1(n8603), .A2(n8190), .A3(n8299), .A4(n8372), .ZN(n7491)
         );
  INV_X1 U9111 ( .A(n12011), .ZN(n8274) );
  AND2_X1 U9112 ( .A1(n13734), .A2(n14682), .ZN(n7492) );
  INV_X1 U9113 ( .A(n8291), .ZN(n8290) );
  OAI21_X1 U9114 ( .B1(n12659), .B2(n8294), .A(n8293), .ZN(n8291) );
  AND2_X1 U9115 ( .A1(n12010), .A2(n12006), .ZN(n7493) );
  AND2_X1 U9116 ( .A1(n9149), .A2(n9147), .ZN(n9387) );
  AND2_X1 U9117 ( .A1(n8450), .A2(n7831), .ZN(n7494) );
  INV_X1 U9118 ( .A(n8128), .ZN(n8127) );
  NOR2_X1 U9119 ( .A1(n9859), .A2(n14351), .ZN(n8128) );
  OR2_X1 U9120 ( .A1(n10408), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7495) );
  NAND2_X1 U9121 ( .A1(n15076), .A2(n15166), .ZN(n7496) );
  NOR2_X1 U9122 ( .A1(n15340), .A2(n8298), .ZN(n7497) );
  INV_X1 U9123 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n9212) );
  NOR2_X1 U9124 ( .A1(n12659), .A2(n16251), .ZN(n8292) );
  NOR2_X1 U9125 ( .A1(n14053), .A2(n12263), .ZN(n7498) );
  INV_X1 U9126 ( .A(n8112), .ZN(n8111) );
  NAND2_X1 U9127 ( .A1(n8115), .A2(n12474), .ZN(n8112) );
  NOR2_X1 U9128 ( .A1(n13291), .A2(n13290), .ZN(n7499) );
  AND2_X1 U9129 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_26__SCAN_IN), .ZN(
        n7500) );
  NOR2_X1 U9130 ( .A1(n14969), .A2(n14819), .ZN(n7501) );
  AND2_X1 U9131 ( .A1(n14794), .A2(n7830), .ZN(n7502) );
  AND2_X1 U9132 ( .A1(n9046), .A2(n7895), .ZN(n7503) );
  OR2_X1 U9133 ( .A1(n13777), .A2(n7481), .ZN(n7504) );
  OR2_X1 U9134 ( .A1(n15485), .A2(n15295), .ZN(n7505) );
  OR2_X1 U9135 ( .A1(n9255), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n7506) );
  INV_X1 U9136 ( .A(n8641), .ZN(n8251) );
  INV_X1 U9137 ( .A(n12166), .ZN(n8275) );
  NOR2_X1 U9138 ( .A1(n12272), .A2(n15186), .ZN(n12166) );
  NOR2_X1 U9139 ( .A1(n13332), .A2(n15158), .ZN(n7507) );
  OR2_X1 U9140 ( .A1(n11493), .A2(n11587), .ZN(n7508) );
  OR2_X1 U9141 ( .A1(n13819), .A2(n13821), .ZN(n7509) );
  NAND2_X1 U9142 ( .A1(n10407), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7510) );
  OR2_X1 U9143 ( .A1(n14785), .A2(n14959), .ZN(n7511) );
  INV_X1 U9144 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10464) );
  NAND2_X1 U9145 ( .A1(n13754), .A2(n13755), .ZN(n7512) );
  AND2_X1 U9146 ( .A1(n16157), .A2(n11918), .ZN(n7513) );
  AND2_X1 U9147 ( .A1(n13593), .A2(n13592), .ZN(n7514) );
  OAI21_X1 U9148 ( .B1(n8329), .B2(n7801), .A(n8326), .ZN(n7800) );
  NAND2_X1 U9149 ( .A1(n8307), .A2(n9935), .ZN(n7515) );
  NOR2_X1 U9150 ( .A1(n15393), .A2(n15409), .ZN(n7516) );
  INV_X1 U9151 ( .A(n8283), .ZN(n8282) );
  AND2_X1 U9152 ( .A1(n15443), .A2(n7470), .ZN(n8283) );
  AND2_X1 U9153 ( .A1(n14372), .A2(n14223), .ZN(n7517) );
  AND2_X1 U9154 ( .A1(n7559), .A2(n7857), .ZN(n7518) );
  NAND2_X1 U9155 ( .A1(n12582), .A2(n8114), .ZN(n7519) );
  NOR2_X1 U9156 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n7520) );
  INV_X1 U9157 ( .A(n9062), .ZN(n7879) );
  INV_X1 U9158 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10425) );
  NAND2_X1 U9159 ( .A1(n9932), .A2(n9933), .ZN(n14188) );
  INV_X1 U9160 ( .A(n14188), .ZN(n9935) );
  INV_X1 U9161 ( .A(n12486), .ZN(n16251) );
  AND2_X1 U9162 ( .A1(n7769), .A2(n9387), .ZN(n7521) );
  INV_X1 U9163 ( .A(n9080), .ZN(n7899) );
  OR2_X1 U9164 ( .A1(P3_IR_REG_26__SCAN_IN), .A2(P3_IR_REG_25__SCAN_IN), .ZN(
        n7522) );
  OR2_X1 U9165 ( .A1(n15807), .A2(n15806), .ZN(n7523) );
  AND2_X1 U9166 ( .A1(n14249), .A2(n7951), .ZN(n7524) );
  INV_X1 U9167 ( .A(n13338), .ZN(n15330) );
  NOR2_X1 U9168 ( .A1(n14975), .A2(n14620), .ZN(n7525) );
  OR2_X1 U9169 ( .A1(n7436), .A2(n8123), .ZN(n7526) );
  AND2_X1 U9170 ( .A1(n15362), .A2(n15097), .ZN(n7527) );
  NOR2_X1 U9171 ( .A1(n15325), .A2(n8258), .ZN(n7528) );
  AND2_X1 U9172 ( .A1(n8429), .A2(SI_10_), .ZN(n7529) );
  AND2_X1 U9173 ( .A1(n7950), .A2(n10030), .ZN(n7530) );
  NAND2_X1 U9174 ( .A1(n7928), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n7625) );
  INV_X1 U9175 ( .A(n7625), .ZN(n7576) );
  AND2_X1 U9176 ( .A1(n8167), .A2(n8163), .ZN(n7531) );
  AND2_X1 U9177 ( .A1(n10042), .A2(n10041), .ZN(n7532) );
  AND2_X1 U9178 ( .A1(n8365), .A2(n8321), .ZN(n7533) );
  AND2_X1 U9179 ( .A1(n11487), .A2(n7788), .ZN(n7534) );
  AND2_X1 U9180 ( .A1(n7795), .A2(n13713), .ZN(n7535) );
  NAND2_X1 U9181 ( .A1(n10948), .A2(n10947), .ZN(n7536) );
  NAND2_X1 U9182 ( .A1(n9862), .A2(n14174), .ZN(n7537) );
  NOR2_X1 U9183 ( .A1(n15525), .A2(n15181), .ZN(n7538) );
  AND2_X1 U9184 ( .A1(n8297), .A2(n7446), .ZN(n7539) );
  AND2_X1 U9185 ( .A1(n15308), .A2(n7446), .ZN(n7540) );
  OR2_X1 U9186 ( .A1(n7463), .A2(n8332), .ZN(n7541) );
  INV_X1 U9187 ( .A(n14236), .ZN(n14232) );
  AND2_X1 U9188 ( .A1(n10039), .A2(n10040), .ZN(n14236) );
  NAND2_X1 U9189 ( .A1(n10027), .A2(n10028), .ZN(n7542) );
  OR2_X1 U9190 ( .A1(n8234), .A2(n9077), .ZN(n7543) );
  OR2_X1 U9191 ( .A1(n9057), .A2(n9055), .ZN(n7544) );
  OR2_X1 U9192 ( .A1(n9007), .A2(n9005), .ZN(n7545) );
  OR2_X1 U9193 ( .A1(n7462), .A2(n7812), .ZN(n7546) );
  AND2_X1 U9194 ( .A1(n13270), .A2(n8359), .ZN(n7547) );
  NAND2_X1 U9195 ( .A1(n7471), .A2(n9707), .ZN(n7548) );
  AND2_X1 U9196 ( .A1(n13341), .A2(n13340), .ZN(n7549) );
  OR2_X1 U9197 ( .A1(n7875), .A2(n9031), .ZN(n7550) );
  OR2_X1 U9198 ( .A1(n13731), .A2(n7451), .ZN(n7551) );
  NAND2_X1 U9199 ( .A1(n15454), .A2(n13357), .ZN(n7552) );
  AND2_X1 U9200 ( .A1(n7878), .A2(n9060), .ZN(n7553) );
  NAND2_X1 U9201 ( .A1(n7885), .A2(n7883), .ZN(n7554) );
  AND2_X1 U9202 ( .A1(n7504), .A2(n7811), .ZN(n7555) );
  AND2_X1 U9203 ( .A1(n8028), .A2(n8027), .ZN(n7556) );
  AND2_X1 U9204 ( .A1(n9211), .A2(n9212), .ZN(n7557) );
  NAND2_X1 U9205 ( .A1(n11598), .A2(n11597), .ZN(n7558) );
  INV_X1 U9206 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8500) );
  INV_X1 U9207 ( .A(n13336), .ZN(n15396) );
  INV_X1 U9208 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8043) );
  INV_X1 U9209 ( .A(n7860), .ZN(n7859) );
  NAND2_X1 U9210 ( .A1(n7862), .A2(n9853), .ZN(n7860) );
  INV_X1 U9211 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n7673) );
  MUX2_X2 U9212 ( .A(n12527), .B(n10881), .S(n8954), .Z(n8952) );
  XOR2_X1 U9213 ( .A(n9858), .B(n14186), .Z(n7559) );
  AND2_X1 U9214 ( .A1(n9670), .A2(n9669), .ZN(n14197) );
  INV_X1 U9215 ( .A(n14197), .ZN(n8346) );
  OR2_X1 U9216 ( .A1(n12703), .A2(n12702), .ZN(n13356) );
  AOI21_X1 U9217 ( .B1(n14172), .B2(n9708), .A(n9705), .ZN(n14044) );
  INV_X1 U9218 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n7749) );
  INV_X1 U9219 ( .A(n13645), .ZN(n8152) );
  INV_X1 U9220 ( .A(n10020), .ZN(n7697) );
  INV_X1 U9221 ( .A(n14981), .ZN(n7971) );
  NAND2_X1 U9222 ( .A1(n13443), .A2(n13442), .ZN(n14886) );
  INV_X1 U9223 ( .A(n14886), .ZN(n8168) );
  AND2_X1 U9224 ( .A1(n16232), .A2(n13230), .ZN(n7560) );
  NAND2_X1 U9225 ( .A1(n8353), .A2(n8362), .ZN(n9563) );
  NOR2_X1 U9226 ( .A1(n12130), .A2(n12129), .ZN(n7561) );
  INV_X1 U9227 ( .A(n7974), .ZN(n12554) );
  NOR2_X1 U9228 ( .A1(n12485), .A2(n8369), .ZN(n7562) );
  AND2_X1 U9229 ( .A1(n13356), .A2(n7459), .ZN(n7563) );
  INV_X1 U9230 ( .A(n7783), .ZN(n7782) );
  NAND2_X1 U9231 ( .A1(n15412), .A2(n13361), .ZN(n7783) );
  OR2_X1 U9232 ( .A1(n15079), .A2(n15406), .ZN(n8009) );
  NAND2_X1 U9233 ( .A1(n13349), .A2(n16110), .ZN(n16179) );
  NAND2_X1 U9234 ( .A1(n11894), .A2(n14840), .ZN(n14843) );
  NAND2_X1 U9235 ( .A1(n10978), .A2(n10977), .ZN(n16315) );
  INV_X1 U9236 ( .A(n13637), .ZN(n8035) );
  INV_X1 U9237 ( .A(n13774), .ZN(n7975) );
  INV_X1 U9238 ( .A(n14085), .ZN(n7905) );
  INV_X1 U9239 ( .A(SI_20_), .ZN(n11612) );
  INV_X1 U9240 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7716) );
  AND2_X1 U9241 ( .A1(n16165), .A2(n8063), .ZN(n7564) );
  NAND2_X1 U9242 ( .A1(n9104), .A2(n9112), .ZN(n10504) );
  NAND2_X1 U9243 ( .A1(n12510), .A2(n12509), .ZN(n15017) );
  INV_X1 U9244 ( .A(n15017), .ZN(n7973) );
  NAND2_X1 U9245 ( .A1(n11721), .A2(n9781), .ZN(n11831) );
  AND2_X1 U9246 ( .A1(n7786), .A2(n7784), .ZN(n11917) );
  AND2_X1 U9247 ( .A1(n11797), .A2(n10400), .ZN(n10129) );
  NAND2_X1 U9248 ( .A1(n9229), .A2(n9228), .ZN(n9767) );
  NAND2_X1 U9249 ( .A1(n12170), .A2(n12169), .ZN(n12488) );
  NAND2_X1 U9250 ( .A1(n11921), .A2(n11920), .ZN(n12012) );
  INV_X1 U9251 ( .A(n8050), .ZN(n11646) );
  OR2_X1 U9252 ( .A1(n11647), .A2(n11648), .ZN(n8050) );
  AND2_X1 U9253 ( .A1(n8087), .A2(n8090), .ZN(n7565) );
  AND2_X1 U9254 ( .A1(n8197), .A2(n8201), .ZN(n7566) );
  INV_X1 U9255 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10725) );
  AND2_X1 U9256 ( .A1(n8295), .A2(n8294), .ZN(n7567) );
  AND2_X1 U9257 ( .A1(n11841), .A2(n9391), .ZN(n7568) );
  AND2_X1 U9258 ( .A1(n12131), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n10207) );
  INV_X1 U9259 ( .A(n14129), .ZN(n7984) );
  NAND2_X1 U9260 ( .A1(n8070), .A2(n15711), .ZN(n10661) );
  INV_X1 U9261 ( .A(n15175), .ZN(n16356) );
  NAND2_X1 U9262 ( .A1(n10162), .A2(n14141), .ZN(n16013) );
  OR2_X1 U9263 ( .A1(n11282), .A2(n11281), .ZN(n7569) );
  NAND2_X1 U9264 ( .A1(n10531), .A2(n10530), .ZN(n15175) );
  INV_X1 U9265 ( .A(n7991), .ZN(n15970) );
  AND2_X1 U9266 ( .A1(n8064), .A2(n14628), .ZN(n7570) );
  AND2_X1 U9267 ( .A1(n7457), .A2(n9192), .ZN(n7571) );
  NAND2_X1 U9268 ( .A1(n11112), .A2(n8053), .ZN(n11509) );
  INV_X1 U9269 ( .A(n11509), .ZN(n8052) );
  NOR2_X1 U9270 ( .A1(n14152), .A2(n7995), .ZN(n7572) );
  AND2_X1 U9271 ( .A1(n9866), .A2(n10395), .ZN(n16041) );
  INV_X1 U9272 ( .A(n16041), .ZN(n14041) );
  INV_X2 U9273 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U9274 ( .A(n11711), .ZN(n7717) );
  INV_X1 U9275 ( .A(n10078), .ZN(n8142) );
  INV_X1 U9276 ( .A(n11374), .ZN(n7977) );
  INV_X1 U9277 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n7609) );
  INV_X1 U9278 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7773) );
  INV_X1 U9279 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7927) );
  INV_X1 U9280 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7931) );
  INV_X1 U9281 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7637) );
  NOR2_X2 U9282 ( .A1(n10616), .A2(n13245), .ZN(n15780) );
  OR2_X2 U9283 ( .A1(n10535), .A2(n10104), .ZN(n15196) );
  INV_X1 U9284 ( .A(n16007), .ZN(n7573) );
  NAND2_X1 U9285 ( .A1(n7989), .A2(n7992), .ZN(n15972) );
  NOR2_X1 U9286 ( .A1(n15975), .A2(n7621), .ZN(n10113) );
  INV_X1 U9287 ( .A(n15878), .ZN(n7575) );
  NOR2_X1 U9288 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n15884), .ZN(n15885) );
  NOR2_X1 U9289 ( .A1(n15894), .A2(n15893), .ZN(n15895) );
  NOR2_X2 U9290 ( .A1(n15923), .A2(n15924), .ZN(n15926) );
  AOI22_X2 U9291 ( .A1(n14182), .A2(n14188), .B1(n14174), .B2(n9860), .ZN(
        n14175) );
  AOI21_X2 U9292 ( .B1(n14220), .B2(n9657), .A(n7647), .ZN(n14209) );
  NAND2_X2 U9293 ( .A1(n10131), .A2(n10420), .ZN(n9562) );
  OAI21_X2 U9294 ( .B1(n13172), .B2(n9812), .A(n9811), .ZN(n13186) );
  AND2_X2 U9295 ( .A1(n9596), .A2(n9595), .ZN(n14279) );
  NAND2_X1 U9296 ( .A1(n13208), .A2(n13209), .ZN(n9525) );
  NAND2_X1 U9297 ( .A1(n14301), .A2(n9577), .ZN(n14289) );
  NAND2_X1 U9298 ( .A1(n9376), .A2(n9375), .ZN(n11757) );
  NAND2_X1 U9299 ( .A1(n9311), .A2(n9310), .ZN(n10383) );
  NAND2_X1 U9300 ( .A1(n7578), .A2(n9321), .ZN(n10385) );
  INV_X1 U9301 ( .A(n10383), .ZN(n7578) );
  NAND2_X1 U9302 ( .A1(n7579), .A2(n11247), .ZN(n9300) );
  AND3_X2 U9303 ( .A1(n9290), .A2(n9291), .A3(n9289), .ZN(n11247) );
  NAND2_X1 U9304 ( .A1(n14177), .A2(n8307), .ZN(n7628) );
  NAND2_X1 U9305 ( .A1(n12062), .A2(n12063), .ZN(n12295) );
  AOI21_X2 U9306 ( .B1(n14577), .B2(n14576), .A(n14520), .ZN(n14656) );
  OAI22_X1 U9307 ( .A1(n14569), .A2(n14568), .B1(n14503), .B2(n14502), .ZN(
        n14504) );
  NOR2_X2 U9308 ( .A1(n14584), .A2(n14585), .ZN(n14583) );
  NAND2_X1 U9309 ( .A1(n11393), .A2(n11392), .ZN(n11536) );
  OR3_X2 U9310 ( .A1(n14739), .A2(n14821), .A3(n14738), .ZN(n14742) );
  AOI21_X1 U9311 ( .B1(n14817), .B2(n14818), .A(n7525), .ZN(n8036) );
  NAND2_X1 U9312 ( .A1(n13498), .A2(n14768), .ZN(n14773) );
  NAND2_X1 U9313 ( .A1(n13598), .A2(n8177), .ZN(n8176) );
  NAND2_X1 U9314 ( .A1(n8176), .A2(n8175), .ZN(n8174) );
  NAND2_X1 U9315 ( .A1(n15403), .A2(n15402), .ZN(n15401) );
  OAI21_X2 U9316 ( .B1(n11495), .B2(n8006), .A(n8004), .ZN(n11925) );
  OAI21_X2 U9317 ( .B1(n15278), .B2(n15280), .A(n7505), .ZN(n15262) );
  INV_X1 U9318 ( .A(n11304), .ZN(n7582) );
  NAND2_X1 U9319 ( .A1(n8003), .A2(n11011), .ZN(n11013) );
  NAND2_X1 U9320 ( .A1(n12165), .A2(n12164), .ZN(n12483) );
  NAND4_X1 U9321 ( .A1(n7491), .A2(n8378), .A3(n8187), .A4(n9107), .ZN(n7581)
         );
  NAND2_X1 U9322 ( .A1(n11492), .A2(n11491), .ZN(n11511) );
  NAND2_X1 U9323 ( .A1(n15371), .A2(n13365), .ZN(n15353) );
  NAND2_X1 U9324 ( .A1(n15372), .A2(n15373), .ZN(n15371) );
  NAND2_X1 U9325 ( .A1(n8905), .A2(n8495), .ZN(n8908) );
  NAND2_X1 U9326 ( .A1(n9092), .A2(n7477), .ZN(n9135) );
  NAND2_X1 U9327 ( .A1(n13860), .A2(n13859), .ZN(n7592) );
  OAI21_X1 U9328 ( .B1(n13794), .B2(n13793), .A(n7541), .ZN(n8331) );
  NAND2_X1 U9329 ( .A1(n7593), .A2(n7590), .ZN(n8319) );
  OR2_X1 U9330 ( .A1(n13828), .A2(n13827), .ZN(n13833) );
  OAI22_X1 U9331 ( .A1(n13833), .A2(n8310), .B1(n13834), .B2(n8311), .ZN(
        n13838) );
  OAI21_X1 U9332 ( .B1(n7445), .B2(n7810), .A(n7555), .ZN(n8333) );
  OAI22_X1 U9333 ( .A1(n7813), .A2(n13814), .B1(n13820), .B2(n7814), .ZN(
        n13826) );
  NAND4_X4 U9334 ( .A1(n10302), .A2(n10301), .A3(n10300), .A4(n10299), .ZN(
        n13669) );
  OR2_X1 U9335 ( .A1(n13694), .A2(n13699), .ZN(n13703) );
  NAND2_X1 U9336 ( .A1(n7589), .A2(n7588), .ZN(n13739) );
  INV_X1 U9337 ( .A(n13873), .ZN(n7593) );
  OAI21_X1 U9338 ( .B1(n13792), .B2(n8331), .A(n8330), .ZN(n13803) );
  INV_X1 U9339 ( .A(n7583), .ZN(n14735) );
  OAI21_X2 U9340 ( .B1(n14918), .B2(n14919), .A(n13535), .ZN(n14893) );
  AOI21_X1 U9341 ( .B1(n14756), .B2(n13511), .A(n13651), .ZN(n14738) );
  OAI22_X2 U9342 ( .A1(n14482), .A2(n14481), .B1(n14480), .B2(n14479), .ZN(
        n14584) );
  NAND2_X1 U9343 ( .A1(n11859), .A2(n11858), .ZN(n12025) );
  NAND2_X1 U9344 ( .A1(n13461), .A2(n13460), .ZN(n14817) );
  NAND2_X1 U9345 ( .A1(n12366), .A2(n12365), .ZN(n12476) );
  NAND3_X1 U9346 ( .A1(n8086), .A2(n11908), .A3(n8085), .ZN(n12061) );
  NOR2_X1 U9347 ( .A1(n15926), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n15927) );
  NOR2_X1 U9348 ( .A1(n15910), .A2(n15909), .ZN(n15911) );
  NOR2_X1 U9349 ( .A1(n15915), .A2(n15914), .ZN(n15918) );
  OAI22_X1 U9350 ( .A1(n14551), .A2(n14550), .B1(n14549), .B2(n14548), .ZN(
        n14556) );
  NAND3_X1 U9351 ( .A1(n13726), .A2(n13725), .A3(n7551), .ZN(n7589) );
  AOI22_X1 U9352 ( .A1(n13406), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n13405), 
        .B2(n11132), .ZN(n11133) );
  XNOR2_X2 U9353 ( .A(n8144), .B(n8322), .ZN(n15064) );
  NAND2_X1 U9354 ( .A1(n11329), .A2(n11330), .ZN(n11328) );
  INV_X1 U9355 ( .A(n11943), .ZN(n7654) );
  NAND2_X1 U9356 ( .A1(n9830), .A2(n9829), .ZN(n14013) );
  NAND2_X1 U9357 ( .A1(n13934), .A2(n9819), .ZN(n14030) );
  NAND2_X1 U9358 ( .A1(n13227), .A2(n9817), .ZN(n13936) );
  NAND2_X1 U9359 ( .A1(n8136), .A2(n9841), .ZN(n13960) );
  NAND2_X1 U9360 ( .A1(n7920), .A2(n10856), .ZN(n7596) );
  NAND2_X1 U9361 ( .A1(n10139), .A2(n7908), .ZN(n11088) );
  NAND2_X1 U9362 ( .A1(n14635), .A2(n14490), .ZN(n8101) );
  NAND2_X1 U9363 ( .A1(n8098), .A2(n8099), .ZN(n8096) );
  NAND2_X1 U9364 ( .A1(n7620), .A2(n7508), .ZN(n11495) );
  AOI22_X1 U9365 ( .A1(n15294), .A2(n15293), .B1(n15125), .B2(n15491), .ZN(
        n15278) );
  NAND2_X1 U9366 ( .A1(n7438), .A2(n13363), .ZN(n15372) );
  NAND2_X1 U9367 ( .A1(n12008), .A2(n12007), .ZN(n12163) );
  NOR2_X2 U9368 ( .A1(n12483), .A2(n12482), .ZN(n12485) );
  NAND2_X2 U9369 ( .A1(n15588), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8783) );
  NAND2_X1 U9370 ( .A1(n11928), .A2(n11927), .ZN(n16156) );
  NAND2_X1 U9371 ( .A1(n8255), .A2(n8253), .ZN(n15294) );
  NAND2_X1 U9372 ( .A1(n15401), .A2(n13362), .ZN(n15385) );
  INV_X1 U9373 ( .A(n11511), .ZN(n7620) );
  XNOR2_X1 U9374 ( .A(n13369), .B(n13342), .ZN(n7644) );
  NAND2_X1 U9375 ( .A1(n7644), .A2(n16330), .ZN(n8007) );
  AOI21_X1 U9376 ( .B1(n7839), .B2(n7841), .A(n7529), .ZN(n7837) );
  NAND2_X1 U9377 ( .A1(n8297), .A2(n7540), .ZN(n15307) );
  INV_X1 U9378 ( .A(n13586), .ZN(n8185) );
  AOI22_X1 U9379 ( .A1(n15303), .A2(n15302), .B1(n15312), .B2(n15491), .ZN(
        n15281) );
  NAND2_X1 U9380 ( .A1(n15279), .A2(n7549), .ZN(n15268) );
  NAND2_X1 U9381 ( .A1(n13598), .A2(n8182), .ZN(n8181) );
  NAND2_X1 U9382 ( .A1(n7776), .A2(n7775), .ZN(n15359) );
  XNOR2_X1 U9383 ( .A(n7601), .B(n7600), .ZN(n7836) );
  NAND2_X1 U9384 ( .A1(n7656), .A2(n7602), .ZN(n7601) );
  NAND2_X1 U9385 ( .A1(n7418), .A2(n14672), .ZN(n7602) );
  OAI21_X1 U9386 ( .B1(n14773), .B2(n7820), .A(n7816), .ZN(n7656) );
  OAI211_X1 U9387 ( .C1(n14947), .C2(n14998), .A(n14945), .B(n14946), .ZN(
        n15036) );
  OR2_X2 U9388 ( .A1(n8613), .A2(n8448), .ZN(n7832) );
  OAI21_X1 U9389 ( .B1(n14750), .B2(n14753), .A(n13548), .ZN(n14734) );
  NAND2_X1 U9390 ( .A1(n12522), .A2(n8150), .ZN(n15020) );
  NAND2_X1 U9391 ( .A1(n11042), .A2(n11041), .ZN(n11388) );
  INV_X1 U9392 ( .A(n11202), .ZN(n13625) );
  NAND2_X1 U9393 ( .A1(n7634), .A2(n7633), .ZN(n12522) );
  NAND2_X1 U9394 ( .A1(n15020), .A2(n8149), .ZN(n13534) );
  NAND2_X1 U9395 ( .A1(n12411), .A2(n12410), .ZN(n12520) );
  NAND2_X1 U9396 ( .A1(n11037), .A2(n11038), .ZN(n8143) );
  NAND2_X1 U9397 ( .A1(n10327), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10314) );
  NAND2_X1 U9398 ( .A1(n14734), .A2(n14737), .ZN(n14736) );
  NAND2_X1 U9399 ( .A1(n13545), .A2(n13544), .ZN(n14769) );
  NAND2_X1 U9400 ( .A1(n15869), .A2(n15870), .ZN(n15871) );
  NAND2_X1 U9401 ( .A1(n7606), .A2(n15881), .ZN(n7611) );
  NAND2_X1 U9402 ( .A1(n15878), .A2(n15879), .ZN(n7606) );
  AOI21_X2 U9403 ( .B1(n15913), .B2(n15912), .A(n15911), .ZN(n15914) );
  NOR2_X2 U9404 ( .A1(n15886), .A2(n15885), .ZN(n15893) );
  INV_X1 U9405 ( .A(n15828), .ZN(n7925) );
  NAND2_X1 U9406 ( .A1(n15788), .A2(n10633), .ZN(n7608) );
  INV_X1 U9407 ( .A(n15814), .ZN(n7610) );
  XNOR2_X1 U9408 ( .A(n15807), .B(n15806), .ZN(n15805) );
  XNOR2_X1 U9409 ( .A(n15796), .B(n15795), .ZN(n15797) );
  NAND2_X1 U9410 ( .A1(n9086), .A2(n9087), .ZN(n7616) );
  NAND3_X1 U9411 ( .A1(n9030), .A2(n7550), .A3(n7613), .ZN(n7612) );
  NOR2_X1 U9412 ( .A1(n15797), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n15798) );
  NAND2_X1 U9413 ( .A1(n9098), .A2(n8847), .ZN(n10872) );
  OAI22_X2 U9414 ( .A1(n9017), .A2(n8242), .B1(n9018), .B2(n8241), .ZN(n9021)
         );
  OAI22_X1 U9415 ( .A1(n9066), .A2(n8240), .B1(n9067), .B2(n8239), .ZN(n9071)
         );
  OAI22_X2 U9416 ( .A1(n8985), .A2(n8238), .B1(n8986), .B2(n8237), .ZN(n8990)
         );
  OAI22_X2 U9417 ( .A1(n8973), .A2(n8236), .B1(n8974), .B2(n8235), .ZN(n8978)
         );
  NAND2_X1 U9418 ( .A1(n7615), .A2(n7614), .ZN(n8970) );
  OAI21_X1 U9419 ( .B1(n9085), .B2(n15193), .A(n11114), .ZN(n7614) );
  NAND2_X1 U9420 ( .A1(n8969), .A2(n16077), .ZN(n7615) );
  AOI21_X1 U9421 ( .B1(n7777), .B2(n7780), .A(n7538), .ZN(n7775) );
  NAND2_X1 U9422 ( .A1(n7881), .A2(n7880), .ZN(n9010) );
  NAND2_X1 U9423 ( .A1(n7900), .A2(n8233), .ZN(n9082) );
  AND3_X2 U9424 ( .A1(n7618), .A2(n7617), .A3(n7616), .ZN(n9093) );
  NAND2_X1 U9425 ( .A1(n9061), .A2(n7553), .ZN(n7877) );
  AND3_X2 U9426 ( .A1(n8778), .A2(n8777), .A3(n8776), .ZN(n10876) );
  OR2_X2 U9427 ( .A1(n15089), .A2(n12651), .ZN(n12695) );
  NAND2_X1 U9428 ( .A1(n8059), .A2(n15428), .ZN(n15404) );
  NOR2_X2 U9429 ( .A1(n15525), .A2(n15388), .ZN(n15378) );
  NOR2_X2 U9430 ( .A1(n7437), .A2(n15274), .ZN(n7619) );
  INV_X1 U9431 ( .A(n7656), .ZN(n14739) );
  XNOR2_X2 U9432 ( .A(n14691), .B(n7432), .ZN(n13622) );
  AND2_X1 U9433 ( .A1(n8762), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n8364) );
  AND3_X2 U9434 ( .A1(n8764), .A2(n8766), .A3(n8765), .ZN(n11074) );
  NOR2_X2 U9435 ( .A1(n14079), .A2(n14078), .ZN(n14077) );
  NOR2_X2 U9436 ( .A1(n12147), .A2(n10121), .ZN(n12142) );
  NOR2_X2 U9437 ( .A1(n12148), .A2(n12500), .ZN(n12147) );
  AOI21_X2 U9438 ( .B1(n15972), .B2(n15970), .A(n15971), .ZN(n15975) );
  NAND2_X1 U9439 ( .A1(n10110), .A2(n10441), .ZN(n10851) );
  AND2_X2 U9440 ( .A1(n8072), .A2(n8071), .ZN(n11125) );
  NOR2_X2 U9441 ( .A1(n14583), .A2(n14486), .ZN(n14595) );
  NAND2_X1 U9442 ( .A1(n13530), .A2(n13529), .ZN(n14925) );
  NAND2_X1 U9443 ( .A1(n15036), .A2(n7419), .ZN(n7835) );
  XNOR2_X1 U9444 ( .A(n15791), .B(n7624), .ZN(n15959) );
  XNOR2_X1 U9445 ( .A(n15790), .B(n7625), .ZN(n15791) );
  NAND3_X1 U9446 ( .A1(n8393), .A2(n16030), .A3(n8392), .ZN(n7639) );
  XNOR2_X1 U9447 ( .A(n8449), .B(n11069), .ZN(n8613) );
  NAND2_X2 U9448 ( .A1(n7838), .A2(n7837), .ZN(n8682) );
  INV_X1 U9449 ( .A(P2_RD_REG_SCAN_IN), .ZN(n8391) );
  NOR2_X1 U9450 ( .A1(n7522), .A2(n9210), .ZN(n8355) );
  NAND2_X1 U9451 ( .A1(n11572), .A2(n11574), .ZN(n11573) );
  NAND2_X1 U9452 ( .A1(n9301), .A2(n9300), .ZN(n16051) );
  AND3_X2 U9453 ( .A1(n9208), .A2(n7557), .A3(n8354), .ZN(n9273) );
  AND2_X2 U9454 ( .A1(n7627), .A2(n7626), .ZN(n14349) );
  NAND3_X1 U9455 ( .A1(n7628), .A2(n14179), .A3(n9714), .ZN(n7627) );
  NAND2_X2 U9456 ( .A1(n14326), .A2(n10008), .ZN(n14314) );
  NAND2_X1 U9457 ( .A1(n7639), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n7638) );
  INV_X1 U9458 ( .A(n12520), .ZN(n7634) );
  NAND2_X1 U9459 ( .A1(n7996), .A2(n7572), .ZN(n7994) );
  NOR2_X1 U9460 ( .A1(n14138), .A2(n7630), .ZN(n14144) );
  AND2_X1 U9461 ( .A1(n14140), .A2(n14139), .ZN(n7630) );
  INV_X1 U9462 ( .A(n11136), .ZN(n8084) );
  NOR2_X2 U9463 ( .A1(n13669), .A2(n13667), .ZN(n13664) );
  NAND2_X1 U9464 ( .A1(n13854), .A2(n13853), .ZN(n13860) );
  NAND2_X1 U9465 ( .A1(n7809), .A2(n8335), .ZN(n13794) );
  AOI21_X1 U9466 ( .B1(n13750), .B2(n13749), .A(n13748), .ZN(n7807) );
  NAND2_X1 U9467 ( .A1(n8225), .A2(n7632), .ZN(n8499) );
  NAND2_X1 U9468 ( .A1(n13744), .A2(n13743), .ZN(n13750) );
  NAND2_X1 U9469 ( .A1(n13808), .A2(n13807), .ZN(n13813) );
  OAI22_X1 U9470 ( .A1(n7808), .A2(n7807), .B1(n13754), .B2(n13755), .ZN(
        n13763) );
  AOI21_X1 U9471 ( .B1(n13843), .B2(n8326), .A(n8324), .ZN(n8323) );
  INV_X2 U9472 ( .A(n11195), .ZN(n14689) );
  NAND2_X1 U9473 ( .A1(n11195), .A2(n13695), .ZN(n11059) );
  AND4_X2 U9474 ( .A1(n10329), .A2(n10330), .A3(n10332), .A4(n10331), .ZN(
        n11195) );
  NAND2_X1 U9475 ( .A1(n14912), .A2(n7556), .ZN(n14899) );
  NAND2_X1 U9476 ( .A1(n12210), .A2(n12209), .ZN(n12418) );
  AND2_X2 U9477 ( .A1(n14899), .A2(n13416), .ZN(n14882) );
  NAND3_X1 U9478 ( .A1(n14748), .A2(n14747), .A3(n7635), .ZN(P2_U3237) );
  NAND3_X1 U9479 ( .A1(n8812), .A2(n8413), .A3(n8420), .ZN(n7821) );
  OAI22_X1 U9480 ( .A1(n14541), .A2(n8096), .B1(n14496), .B2(n14497), .ZN(
        n8095) );
  INV_X1 U9481 ( .A(n8095), .ZN(n8094) );
  OAI21_X2 U9482 ( .B1(n14314), .B2(n14319), .A(n8357), .ZN(n14301) );
  NAND2_X1 U9483 ( .A1(n9946), .A2(n9945), .ZN(n10057) );
  NAND2_X1 U9484 ( .A1(n8368), .A2(n9420), .ZN(n12287) );
  INV_X1 U9485 ( .A(n11843), .ZN(n7646) );
  NAND2_X1 U9486 ( .A1(n7835), .A2(n7834), .ZN(P2_U3496) );
  NAND2_X1 U9487 ( .A1(n8007), .A2(n7642), .ZN(n15568) );
  INV_X1 U9488 ( .A(n14251), .ZN(n7649) );
  NAND2_X1 U9489 ( .A1(n15838), .A2(n15837), .ZN(n7930) );
  AND2_X2 U9490 ( .A1(n9201), .A2(n9329), .ZN(n8353) );
  NAND2_X1 U9491 ( .A1(n15935), .A2(n15934), .ZN(n7924) );
  NAND2_X1 U9492 ( .A1(n11803), .A2(n9358), .ZN(n11755) );
  OAI21_X1 U9493 ( .B1(n15917), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7932), .ZN(
        n15923) );
  AOI21_X1 U9494 ( .B1(n8048), .B2(n11535), .A(n7472), .ZN(n8047) );
  NAND2_X1 U9495 ( .A1(n14742), .A2(n14741), .ZN(n7655) );
  OAI21_X1 U9496 ( .B1(n7487), .B2(n7650), .A(n8231), .ZN(n9061) );
  NAND2_X1 U9497 ( .A1(n9054), .A2(n7544), .ZN(n7650) );
  NAND2_X1 U9498 ( .A1(n9035), .A2(n9036), .ZN(n9034) );
  NAND2_X1 U9499 ( .A1(n7877), .A2(n7876), .ZN(n9066) );
  NAND2_X1 U9500 ( .A1(n9082), .A2(n7899), .ZN(n7898) );
  NAND2_X1 U9501 ( .A1(n7898), .A2(n9079), .ZN(n9081) );
  NAND2_X1 U9502 ( .A1(n7888), .A2(n7889), .ZN(n9024) );
  AOI21_X1 U9503 ( .B1(n7988), .B2(n11024), .A(n7987), .ZN(n7989) );
  INV_X1 U9504 ( .A(n14147), .ZN(n8000) );
  XNOR2_X1 U9505 ( .A(n10113), .B(n10466), .ZN(n15993) );
  NAND2_X1 U9506 ( .A1(n7822), .A2(n8419), .ZN(n8727) );
  NAND2_X1 U9507 ( .A1(n12061), .A2(n12060), .ZN(n12062) );
  NAND2_X1 U9508 ( .A1(n14516), .A2(n14515), .ZN(n14577) );
  NAND2_X1 U9509 ( .A1(n8088), .A2(n8089), .ZN(n8085) );
  NAND2_X1 U9510 ( .A1(n8105), .A2(n8104), .ZN(n14482) );
  NAND2_X1 U9511 ( .A1(n11604), .A2(n8092), .ZN(n8091) );
  INV_X1 U9512 ( .A(n15918), .ZN(n7932) );
  NAND2_X1 U9513 ( .A1(n15818), .A2(n15817), .ZN(n7926) );
  OAI21_X1 U9514 ( .B1(n13960), .B2(n13958), .A(n13956), .ZN(n9847) );
  NOR2_X2 U9515 ( .A1(n8116), .A2(P3_IR_REG_3__SCAN_IN), .ZN(n9329) );
  NAND2_X1 U9516 ( .A1(n14000), .A2(n13999), .ZN(n8136) );
  INV_X1 U9517 ( .A(n9208), .ZN(n9258) );
  NAND2_X2 U9518 ( .A1(n9208), .A2(n9207), .ZN(n9255) );
  INV_X1 U9519 ( .A(n8131), .ZN(n8130) );
  OAI21_X2 U9520 ( .B1(n14816), .B2(n8147), .A(n8145), .ZN(n14784) );
  OAI21_X1 U9521 ( .B1(n7825), .B2(n7824), .A(n7823), .ZN(n13498) );
  AOI21_X1 U9522 ( .B1(n13403), .B2(n13402), .A(n13401), .ZN(n14913) );
  NOR2_X2 U9523 ( .A1(n10269), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n15052) );
  NAND2_X1 U9524 ( .A1(n8320), .A2(n7533), .ZN(n10269) );
  NAND2_X1 U9525 ( .A1(n15326), .A2(n8252), .ZN(n8255) );
  NAND2_X1 U9526 ( .A1(n12703), .A2(n7459), .ZN(n8015) );
  NAND2_X1 U9527 ( .A1(n11925), .A2(n11924), .ZN(n11928) );
  NAND2_X2 U9528 ( .A1(n10952), .A2(n10951), .ZN(n11275) );
  NAND2_X1 U9529 ( .A1(n13555), .A2(n8209), .ZN(n15093) );
  INV_X1 U9530 ( .A(n7661), .ZN(n13300) );
  OR2_X1 U9531 ( .A1(n9108), .A2(n7671), .ZN(n7668) );
  AND2_X1 U9532 ( .A1(n9108), .A2(n7672), .ZN(n9103) );
  NAND2_X1 U9533 ( .A1(n7668), .A2(n7669), .ZN(n9102) );
  NAND2_X1 U9534 ( .A1(n9108), .A2(n9107), .ZN(n9099) );
  NAND2_X1 U9535 ( .A1(n15165), .A2(n7675), .ZN(n7674) );
  OAI211_X1 U9536 ( .C1(n15165), .C2(n7676), .A(n7674), .B(n15081), .ZN(
        P1_U3214) );
  NAND2_X1 U9537 ( .A1(n13175), .A2(n7690), .ZN(n7686) );
  NAND2_X1 U9538 ( .A1(n7686), .A2(n7687), .ZN(n14334) );
  NAND2_X1 U9539 ( .A1(n14309), .A2(n7695), .ZN(n7694) );
  XNOR2_X1 U9540 ( .A(n14058), .B(n16049), .ZN(n9948) );
  NAND2_X4 U9541 ( .A1(n10131), .A2(n10432), .ZN(n9917) );
  OAI22_X1 U9542 ( .A1(n9562), .A2(n10472), .B1(n10131), .B2(n10170), .ZN(
        n7707) );
  NAND3_X1 U9543 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .A3(
        P1_IR_REG_0__SCAN_IN), .ZN(n7722) );
  NAND2_X1 U9544 ( .A1(n7728), .A2(n10085), .ZN(P3_U3296) );
  NAND2_X1 U9545 ( .A1(n7730), .A2(n16061), .ZN(n7729) );
  INV_X1 U9546 ( .A(n7732), .ZN(n7730) );
  NAND2_X1 U9547 ( .A1(n7732), .A2(n10079), .ZN(n7731) );
  NAND2_X1 U9548 ( .A1(n9414), .A2(n7740), .ZN(n7736) );
  NAND2_X1 U9549 ( .A1(n7736), .A2(n7737), .ZN(n9442) );
  NAND3_X1 U9550 ( .A1(n7478), .A2(n9941), .A3(n7743), .ZN(n7744) );
  NAND2_X1 U9551 ( .A1(n9285), .A2(n9138), .ZN(n9309) );
  NAND2_X1 U9552 ( .A1(n9177), .A2(n7755), .ZN(n7753) );
  NAND2_X1 U9553 ( .A1(n7762), .A2(n7763), .ZN(n9685) );
  NAND2_X1 U9554 ( .A1(n7762), .A2(n7760), .ZN(n9195) );
  NAND2_X1 U9555 ( .A1(n9193), .A2(n9192), .ZN(n9673) );
  NAND2_X1 U9556 ( .A1(n9144), .A2(n7521), .ZN(n7765) );
  NAND2_X1 U9557 ( .A1(n7765), .A2(n7766), .ZN(n9399) );
  NAND2_X1 U9558 ( .A1(n15400), .A2(n7777), .ZN(n7776) );
  NAND2_X1 U9559 ( .A1(n11508), .A2(n7534), .ZN(n7786) );
  NAND2_X1 U9560 ( .A1(n7786), .A2(n7785), .ZN(n8296) );
  NAND4_X1 U9561 ( .A1(n11109), .A2(n7599), .A3(n11104), .A4(n16033), .ZN(
        n8811) );
  NAND4_X1 U9562 ( .A1(n7793), .A2(n8038), .A3(n8040), .A4(n8365), .ZN(n8037)
         );
  NAND2_X1 U9563 ( .A1(n7796), .A2(n7535), .ZN(n8315) );
  NAND2_X1 U9564 ( .A1(n13709), .A2(n7797), .ZN(n7796) );
  INV_X1 U9565 ( .A(n13707), .ZN(n7799) );
  NAND2_X1 U9566 ( .A1(n10286), .A2(n7453), .ZN(n10277) );
  NAND2_X1 U9567 ( .A1(n10286), .A2(n10095), .ZN(n10285) );
  INV_X1 U9568 ( .A(n10277), .ZN(n10282) );
  NAND2_X1 U9569 ( .A1(n13767), .A2(n7546), .ZN(n7810) );
  INV_X1 U9570 ( .A(n13771), .ZN(n7812) );
  NAND2_X1 U9571 ( .A1(n14773), .A2(n14754), .ZN(n7815) );
  NAND2_X1 U9572 ( .A1(n7815), .A2(n14753), .ZN(n14756) );
  NOR2_X1 U9573 ( .A1(n14737), .A2(n7817), .ZN(n7816) );
  NAND2_X1 U9574 ( .A1(n13511), .A2(n7818), .ZN(n7817) );
  NAND2_X1 U9575 ( .A1(n14753), .A2(n7819), .ZN(n7818) );
  INV_X1 U9576 ( .A(n14753), .ZN(n7820) );
  INV_X1 U9577 ( .A(n8036), .ZN(n7825) );
  XNOR2_X2 U9578 ( .A(n8455), .B(n12736), .ZN(n8859) );
  NAND2_X1 U9579 ( .A1(n8427), .A2(n7839), .ZN(n7838) );
  INV_X1 U9580 ( .A(SI_14_), .ZN(n7846) );
  OAI21_X1 U9581 ( .B1(SI_14_), .B2(n8442), .A(n8443), .ZN(n8642) );
  NAND2_X1 U9582 ( .A1(n7863), .A2(n7859), .ZN(n7854) );
  NAND2_X1 U9583 ( .A1(n7863), .A2(n9853), .ZN(n13966) );
  NAND3_X1 U9584 ( .A1(n7860), .A2(n7857), .A3(n7559), .ZN(n7856) );
  NAND2_X1 U9585 ( .A1(n13194), .A2(n7865), .ZN(n13227) );
  NAND2_X1 U9586 ( .A1(n12398), .A2(n7867), .ZN(n10252) );
  NAND3_X1 U9587 ( .A1(n9229), .A2(n8142), .A3(n9228), .ZN(n7873) );
  NAND3_X1 U9588 ( .A1(n9004), .A2(n7882), .A3(n7545), .ZN(n7881) );
  NAND2_X1 U9589 ( .A1(n9021), .A2(n7886), .ZN(n7885) );
  INV_X1 U9590 ( .A(n9050), .ZN(n9053) );
  NAND2_X1 U9591 ( .A1(n7893), .A2(n7894), .ZN(n9050) );
  AND2_X1 U9592 ( .A1(n8603), .A2(n7897), .ZN(n7896) );
  NAND2_X1 U9593 ( .A1(n8225), .A2(n9107), .ZN(n8517) );
  NAND3_X1 U9594 ( .A1(n9076), .A2(n9075), .A3(n7543), .ZN(n7900) );
  XNOR2_X2 U9595 ( .A(n8505), .B(P1_IR_REG_21__SCAN_IN), .ZN(n10881) );
  OAI21_X1 U9596 ( .B1(n12154), .B2(n7907), .A(n7906), .ZN(n10158) );
  XNOR2_X1 U9597 ( .A(n10158), .B(n10210), .ZN(n14061) );
  AOI21_X1 U9598 ( .B1(n7915), .B2(n15979), .A(n7913), .ZN(n14133) );
  AND2_X1 U9599 ( .A1(n14128), .A2(n14129), .ZN(n7918) );
  OAI21_X1 U9600 ( .B1(n15805), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n7523), .ZN(
        n7922) );
  NAND3_X1 U9601 ( .A1(n9328), .A2(n7935), .A3(n7933), .ZN(n9959) );
  NOR2_X2 U9602 ( .A1(n9338), .A2(n7934), .ZN(n11578) );
  NAND2_X1 U9603 ( .A1(n9525), .A2(n7936), .ZN(n14326) );
  NAND2_X1 U9604 ( .A1(n12320), .A2(n7941), .ZN(n7940) );
  NAND2_X1 U9605 ( .A1(n7940), .A2(n7943), .ZN(n13172) );
  INV_X1 U9606 ( .A(n11755), .ZN(n9376) );
  NAND2_X1 U9607 ( .A1(n11573), .A2(n7953), .ZN(n11803) );
  NAND2_X1 U9608 ( .A1(n14179), .A2(n7955), .ZN(n7954) );
  OAI211_X1 U9609 ( .C1(n14179), .C2(n7956), .A(n9725), .B(n7954), .ZN(n14163)
         );
  NAND3_X1 U9610 ( .A1(n9208), .A2(n9211), .A3(n8354), .ZN(n9271) );
  NAND2_X1 U9611 ( .A1(n9208), .A2(n8354), .ZN(n9214) );
  OR2_X1 U9612 ( .A1(n10322), .A2(n10452), .ZN(n7959) );
  OAI21_X2 U9613 ( .B1(n11769), .B2(n7970), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8144) );
  NOR2_X2 U9614 ( .A1(n14925), .A2(n15001), .ZN(n14892) );
  NAND2_X1 U9615 ( .A1(n14107), .A2(n7456), .ZN(n7982) );
  OAI211_X1 U9616 ( .C1(n14107), .C2(n7984), .A(n7982), .B(n7983), .ZN(n14109)
         );
  INV_X1 U9617 ( .A(n10854), .ZN(n7988) );
  NAND2_X1 U9618 ( .A1(n10854), .A2(n7993), .ZN(n7992) );
  XNOR2_X2 U9619 ( .A(n8002), .B(n8001), .ZN(n10170) );
  AND2_X2 U9620 ( .A1(n7685), .A2(n7910), .ZN(n10140) );
  NAND2_X1 U9621 ( .A1(n16156), .A2(n11929), .ZN(n8010) );
  NAND2_X1 U9622 ( .A1(n8010), .A2(n8011), .ZN(n12008) );
  AOI21_X1 U9623 ( .B1(n16157), .B2(n11929), .A(n7493), .ZN(n8011) );
  OR3_X1 U9624 ( .A1(n15461), .A2(n8016), .A3(n8014), .ZN(n8013) );
  NAND2_X1 U9625 ( .A1(n12485), .A2(n7466), .ZN(n8017) );
  NAND2_X1 U9626 ( .A1(n8017), .A2(n8018), .ZN(n12698) );
  OAI21_X2 U9627 ( .B1(n15339), .B2(n13366), .A(n7475), .ZN(n15326) );
  OAI22_X1 U9628 ( .A1(n15262), .A2(n13367), .B1(n15079), .B2(n15274), .ZN(
        n13369) );
  NAND2_X1 U9629 ( .A1(n8024), .A2(n8023), .ZN(n8022) );
  INV_X1 U9630 ( .A(n11131), .ZN(n8024) );
  OAI21_X1 U9632 ( .B1(n10431), .B2(n10464), .A(n8026), .ZN(n8025) );
  NAND2_X1 U9633 ( .A1(n11536), .A2(n8048), .ZN(n8045) );
  NAND2_X1 U9634 ( .A1(n8045), .A2(n8047), .ZN(n11670) );
  NOR2_X2 U9635 ( .A1(n8050), .A2(n16132), .ZN(n16163) );
  NAND4_X1 U9636 ( .A1(n8378), .A2(n8054), .A3(n8188), .A4(n9107), .ZN(n8055)
         );
  NAND2_X1 U9637 ( .A1(n8055), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8498) );
  NOR2_X2 U9638 ( .A1(n15451), .A2(n15550), .ZN(n8059) );
  NAND3_X1 U9639 ( .A1(n16224), .A2(n16165), .A3(n8063), .ZN(n16245) );
  NAND2_X1 U9640 ( .A1(n14628), .A2(n14629), .ZN(n8066) );
  OR2_X1 U9641 ( .A1(n14630), .A2(n14629), .ZN(n8064) );
  NAND2_X1 U9642 ( .A1(n8067), .A2(n8065), .ZN(n10362) );
  AND2_X1 U9643 ( .A1(n8066), .A2(n8068), .ZN(n8065) );
  NAND2_X1 U9644 ( .A1(n14630), .A2(n14628), .ZN(n8067) );
  INV_X1 U9645 ( .A(n10321), .ZN(n8069) );
  XNOR2_X1 U9646 ( .A(n10318), .B(n10317), .ZN(n14562) );
  NAND3_X1 U9647 ( .A1(n8073), .A2(n8075), .A3(n8076), .ZN(n8070) );
  NAND4_X1 U9648 ( .A1(n8073), .A2(n13666), .A3(n8075), .A4(n8076), .ZN(n8072)
         );
  NAND3_X1 U9649 ( .A1(n13912), .A2(n13902), .A3(n13662), .ZN(n8076) );
  NAND3_X1 U9650 ( .A1(n8080), .A2(n14645), .A3(n8081), .ZN(n14644) );
  NAND2_X1 U9651 ( .A1(n11603), .A2(n8088), .ZN(n8086) );
  NAND2_X1 U9652 ( .A1(n8093), .A2(n8094), .ZN(n14611) );
  NAND3_X1 U9653 ( .A1(n14595), .A2(n8097), .A3(n8098), .ZN(n8093) );
  NAND2_X1 U9654 ( .A1(n8101), .A2(n8102), .ZN(n8098) );
  NAND2_X1 U9655 ( .A1(n14493), .A2(n14494), .ZN(n8102) );
  NAND2_X1 U9656 ( .A1(n12476), .A2(n8107), .ZN(n8105) );
  NAND2_X1 U9657 ( .A1(n8116), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9316) );
  INV_X1 U9658 ( .A(n8117), .ZN(n9776) );
  AOI21_X1 U9659 ( .B1(n8117), .B2(n11412), .A(n14041), .ZN(n11414) );
  NAND2_X1 U9660 ( .A1(n14022), .A2(n8119), .ZN(n8118) );
  OAI211_X1 U9661 ( .C1(n14022), .C2(n7454), .A(n8118), .B(n16041), .ZN(n9892)
         );
  OAI21_X1 U9662 ( .B1(n14816), .B2(n14818), .A(n13542), .ZN(n14800) );
  INV_X2 U9663 ( .A(n11080), .ZN(n16032) );
  MUX2_X1 U9664 ( .A(P1_IR_REG_0__SCAN_IN), .B(n15608), .S(n10455), .Z(n11080)
         );
  XNOR2_X2 U9665 ( .A(n8501), .B(n8500), .ZN(n15594) );
  OR2_X1 U9666 ( .A1(n15165), .A2(n8181), .ZN(n8180) );
  NAND3_X1 U9667 ( .A1(n8180), .A2(n8179), .A3(n8174), .ZN(n13603) );
  NAND3_X1 U9668 ( .A1(n15165), .A2(n8183), .A3(n8186), .ZN(n8179) );
  NAND2_X1 U9669 ( .A1(n13264), .A2(n7547), .ZN(n15082) );
  NAND2_X1 U9670 ( .A1(n8194), .A2(n11275), .ZN(n8193) );
  NAND3_X1 U9671 ( .A1(n8198), .A2(n8200), .A3(n11463), .ZN(n8196) );
  AOI22_X1 U9672 ( .A1(n11337), .A2(n8208), .B1(n8201), .B2(n8199), .ZN(n8198)
         );
  INV_X1 U9673 ( .A(n11273), .ZN(n8201) );
  INV_X1 U9674 ( .A(n8206), .ZN(n11464) );
  NAND2_X1 U9675 ( .A1(n11274), .A2(n11273), .ZN(n8208) );
  NAND2_X1 U9676 ( .A1(n15147), .A2(n8210), .ZN(n15112) );
  NAND2_X1 U9677 ( .A1(n11821), .A2(n8212), .ZN(n8214) );
  INV_X1 U9678 ( .A(n8214), .ZN(n11978) );
  NAND2_X1 U9679 ( .A1(n12389), .A2(n8216), .ZN(n8218) );
  INV_X1 U9680 ( .A(n8218), .ZN(n12567) );
  OAI21_X1 U9681 ( .B1(n8997), .B2(n8223), .A(n8222), .ZN(n9002) );
  NAND2_X1 U9682 ( .A1(n8221), .A2(n8219), .ZN(n9001) );
  NAND2_X1 U9683 ( .A1(n8997), .A2(n8222), .ZN(n8221) );
  AND3_X4 U9684 ( .A1(n8774), .A2(n8376), .A3(n8377), .ZN(n9107) );
  NAND2_X1 U9685 ( .A1(n8228), .A2(n8226), .ZN(n9028) );
  AOI21_X1 U9686 ( .B1(n8230), .B2(n8229), .A(n8227), .ZN(n8226) );
  NAND2_X1 U9687 ( .A1(n9024), .A2(n8229), .ZN(n8228) );
  NAND2_X1 U9688 ( .A1(n8978), .A2(n8979), .ZN(n8977) );
  NAND2_X1 U9689 ( .A1(n8990), .A2(n8991), .ZN(n8989) );
  NAND2_X1 U9690 ( .A1(n9071), .A2(n9072), .ZN(n9070) );
  NAND2_X1 U9691 ( .A1(n9010), .A2(n9011), .ZN(n9009) );
  OAI21_X2 U9692 ( .B1(n8859), .B2(n8245), .A(n8456), .ZN(n8846) );
  OAI21_X1 U9693 ( .B1(n8705), .B2(n8247), .A(n8428), .ZN(n8692) );
  OAI21_X1 U9694 ( .B1(n8642), .B2(n8251), .A(n8443), .ZN(n8626) );
  OAI21_X1 U9695 ( .B1(n8590), .B2(n8264), .A(n8263), .ZN(n8577) );
  NAND2_X1 U9696 ( .A1(n8262), .A2(n8260), .ZN(n8464) );
  NAND2_X1 U9697 ( .A1(n8590), .A2(n8263), .ZN(n8262) );
  OAI21_X1 U9698 ( .B1(n8682), .B2(n8681), .A(n8433), .ZN(n8673) );
  NAND2_X1 U9699 ( .A1(n11299), .A2(n8285), .ZN(n8286) );
  NAND3_X1 U9700 ( .A1(n8287), .A2(n11505), .A3(n8286), .ZN(n11508) );
  NAND2_X1 U9701 ( .A1(n11486), .A2(n11485), .ZN(n11506) );
  NAND2_X1 U9702 ( .A1(n11300), .A2(n11488), .ZN(n11486) );
  INV_X1 U9703 ( .A(n8295), .ZN(n16243) );
  OR2_X1 U9704 ( .A1(n16277), .A2(n15183), .ZN(n8293) );
  NAND2_X1 U9705 ( .A1(n15281), .A2(n15280), .ZN(n15279) );
  NAND2_X1 U9706 ( .A1(n15279), .A2(n13340), .ZN(n15266) );
  NAND2_X1 U9707 ( .A1(n8296), .A2(n7513), .ZN(n16152) );
  AND2_X1 U9708 ( .A1(n15349), .A2(n15180), .ZN(n8298) );
  INV_X1 U9709 ( .A(n13832), .ZN(n8311) );
  NAND2_X1 U9710 ( .A1(n8313), .A2(n8312), .ZN(n13721) );
  NAND2_X1 U9711 ( .A1(n8315), .A2(n8314), .ZN(n8313) );
  INV_X1 U9712 ( .A(n13712), .ZN(n8314) );
  OAI211_X1 U9713 ( .C1(n8318), .C2(n13921), .A(n8317), .B(n8316), .ZN(
        P2_U3328) );
  NAND2_X1 U9714 ( .A1(n8318), .A2(n13920), .ZN(n8317) );
  NAND2_X1 U9715 ( .A1(n8319), .A2(n13890), .ZN(n8318) );
  INV_X1 U9716 ( .A(n11769), .ZN(n8320) );
  INV_X1 U9717 ( .A(n8323), .ZN(n13849) );
  NAND2_X1 U9718 ( .A1(n13739), .A2(n13740), .ZN(n13738) );
  INV_X1 U9719 ( .A(n13797), .ZN(n8332) );
  NAND2_X1 U9720 ( .A1(n8333), .A2(n8334), .ZN(n13783) );
  NAND2_X1 U9721 ( .A1(n13763), .A2(n13764), .ZN(n13762) );
  OR2_X2 U9722 ( .A1(n9299), .A2(n11247), .ZN(n9946) );
  INV_X1 U9723 ( .A(n11251), .ZN(n9726) );
  NAND2_X1 U9724 ( .A1(n8349), .A2(n7530), .ZN(n9738) );
  NOR2_X1 U9725 ( .A1(n14189), .A2(n14188), .ZN(n14187) );
  NOR2_X1 U9726 ( .A1(n14187), .A2(n9740), .ZN(n14171) );
  NAND2_X1 U9727 ( .A1(n10535), .A2(n9115), .ZN(n10954) );
  AND2_X1 U9728 ( .A1(n10574), .A2(n10573), .ZN(n10575) );
  NAND2_X1 U9729 ( .A1(n9251), .A2(n9250), .ZN(n9755) );
  NAND2_X1 U9730 ( .A1(n9250), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9248) );
  NAND2_X1 U9731 ( .A1(n11228), .A2(n11229), .ZN(n11227) );
  OAI21_X1 U9732 ( .B1(n15602), .B2(n10507), .A(n10506), .ZN(n15582) );
  INV_X1 U9733 ( .A(n13245), .ZN(n10804) );
  AND2_X1 U9734 ( .A1(n15268), .A2(n15267), .ZN(n15482) );
  AND2_X1 U9735 ( .A1(n16152), .A2(n16151), .ZN(n16178) );
  INV_X1 U9736 ( .A(n8795), .ZN(n8380) );
  INV_X1 U9737 ( .A(n13721), .ZN(n13724) );
  CLKBUF_X1 U9738 ( .A(n10057), .Z(n11251) );
  XNOR2_X1 U9739 ( .A(n9292), .B(n9801), .ZN(n9770) );
  INV_X1 U9740 ( .A(n12272), .ZN(n16216) );
  INV_X2 U9741 ( .A(n16239), .ZN(n16242) );
  NAND2_X1 U9742 ( .A1(n16238), .A2(n16102), .ZN(n14418) );
  AND2_X2 U9743 ( .A1(n10393), .A2(n9761), .ZN(n16238) );
  OR2_X1 U9744 ( .A1(n12388), .A2(n12387), .ZN(n8356) );
  NOR2_X1 U9745 ( .A1(n9576), .A2(n14300), .ZN(n8357) );
  OR2_X1 U9746 ( .A1(n11820), .A2(n11819), .ZN(n8358) );
  OR2_X1 U9747 ( .A1(n13263), .A2(n13262), .ZN(n8359) );
  OR2_X1 U9748 ( .A1(n15318), .A2(n15329), .ZN(n8360) );
  AND2_X1 U9749 ( .A1(n15829), .A2(n15828), .ZN(n8361) );
  INV_X1 U9750 ( .A(n11890), .ZN(n10363) );
  INV_X1 U9751 ( .A(n15485), .ZN(n15288) );
  NOR2_X1 U9752 ( .A1(n14314), .A2(n14319), .ZN(n8363) );
  INV_X1 U9753 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n8732) );
  AND2_X1 U9754 ( .A1(n10432), .A2(P2_U3088), .ZN(n13242) );
  INV_X4 U9755 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  AND2_X1 U9756 ( .A1(n8437), .A2(n8436), .ZN(n8366) );
  INV_X1 U9757 ( .A(n14145), .ZN(n9927) );
  AND2_X1 U9758 ( .A1(n10072), .A2(n14156), .ZN(n8367) );
  INV_X2 U9759 ( .A(P2_U3947), .ZN(n14683) );
  INV_X1 U9760 ( .A(n14166), .ZN(n9268) );
  INV_X1 U9761 ( .A(n16053), .ZN(n9714) );
  AND2_X1 U9762 ( .A1(n12484), .A2(n12489), .ZN(n8369) );
  INV_X1 U9763 ( .A(n11920), .ZN(n11930) );
  CLKBUF_X3 U9764 ( .A(n10669), .Z(n13588) );
  INV_X1 U9765 ( .A(n15171), .ZN(n15295) );
  AND4_X1 U9766 ( .A1(n8548), .A2(n8547), .A3(n8546), .A4(n8545), .ZN(n15171)
         );
  AND2_X1 U9767 ( .A1(n13716), .A2(n13667), .ZN(n13668) );
  NAND2_X1 U9768 ( .A1(n14626), .A2(n13870), .ZN(n13678) );
  INV_X1 U9769 ( .A(n13722), .ZN(n13723) );
  INV_X1 U9770 ( .A(n14044), .ZN(n9706) );
  INV_X1 U9771 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n10088) );
  NAND2_X1 U9772 ( .A1(n14347), .A2(n9706), .ZN(n9707) );
  INV_X1 U9773 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n8373) );
  INV_X1 U9774 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n9480) );
  INV_X1 U9775 ( .A(n9960), .ZN(n9338) );
  INV_X1 U9776 ( .A(n10063), .ZN(n9420) );
  INV_X1 U9777 ( .A(n12540), .ZN(n12539) );
  INV_X1 U9778 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n11863) );
  INV_X1 U9779 ( .A(n12422), .ZN(n12421) );
  OR2_X1 U9780 ( .A1(n11074), .A2(n13587), .ZN(n10574) );
  OR2_X1 U9781 ( .A1(n13273), .A2(n13272), .ZN(n13274) );
  NAND2_X1 U9782 ( .A1(n15485), .A2(n15171), .ZN(n13340) );
  INV_X1 U9783 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n13147) );
  INV_X1 U9784 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n8392) );
  INV_X1 U9785 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n9533) );
  OAI22_X1 U9786 ( .A1(n14044), .A2(n16054), .B1(n14157), .B2(n11792), .ZN(
        n9724) );
  INV_X1 U9787 ( .A(n12325), .ZN(n9731) );
  OR4_X1 U9788 ( .A1(n12929), .A2(n12928), .A3(n12927), .A4(n12926), .ZN(
        n12933) );
  INV_X1 U9789 ( .A(n11754), .ZN(n9375) );
  AND2_X1 U9790 ( .A1(n10129), .A2(n10079), .ZN(n11083) );
  INV_X1 U9791 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13373) );
  INV_X1 U9792 ( .A(n9219), .ZN(n9220) );
  INV_X1 U9793 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n9207) );
  OR2_X1 U9794 ( .A1(n9491), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n9492) );
  AND4_X1 U9795 ( .A1(n9200), .A2(n9199), .A3(n9349), .A4(n9198), .ZN(n9201)
         );
  CLKBUF_X3 U9796 ( .A(n13857), .Z(n13891) );
  OR2_X1 U9797 ( .A1(n13503), .A2(n13381), .ZN(n13516) );
  OR2_X1 U9798 ( .A1(n13452), .A2(n14534), .ZN(n13466) );
  NAND2_X1 U9799 ( .A1(n12539), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13423) );
  OR2_X1 U9800 ( .A1(n11864), .A2(n11863), .ZN(n11875) );
  INV_X1 U9801 ( .A(n13651), .ZN(n14737) );
  OR2_X1 U9802 ( .A1(n13450), .A2(n14619), .ZN(n13452) );
  INV_X1 U9803 ( .A(n15005), .ZN(n13529) );
  NAND2_X1 U9804 ( .A1(n12421), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n12512) );
  INV_X1 U9805 ( .A(n11131), .ZN(n13405) );
  NAND2_X1 U9806 ( .A1(n11131), .A2(n15074), .ZN(n10307) );
  INV_X1 U9807 ( .A(n15085), .ZN(n13270) );
  AND2_X1 U9808 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n8541) );
  INV_X1 U9809 ( .A(n8898), .ZN(n8571) );
  OR2_X1 U9810 ( .A1(n13298), .A2(n13297), .ZN(n13299) );
  AND2_X1 U9811 ( .A1(n8564), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8554) );
  INV_X1 U9812 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8608) );
  INV_X1 U9813 ( .A(n13258), .ZN(n13268) );
  OR2_X1 U9814 ( .A1(n12010), .A2(n15187), .ZN(n12011) );
  AND2_X1 U9815 ( .A1(n9116), .A2(n10533), .ZN(n10953) );
  NOR2_X1 U9816 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n8376) );
  NAND3_X1 U9817 ( .A1(n8391), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n8394) );
  INV_X1 U9818 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n15806) );
  INV_X1 U9819 ( .A(n11412), .ZN(n9775) );
  AND2_X1 U9820 ( .A1(n9700), .A2(n9885), .ZN(n14164) );
  INV_X1 U9821 ( .A(n9551), .ZN(n9708) );
  INV_X1 U9822 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n15868) );
  INV_X1 U9823 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n15890) );
  INV_X1 U9824 ( .A(n9724), .ZN(n9725) );
  INV_X1 U9825 ( .A(n14360), .ZN(n14208) );
  AND2_X1 U9826 ( .A1(n10019), .A2(n9943), .ZN(n14319) );
  INV_X1 U9827 ( .A(n12712), .ZN(n12501) );
  INV_X1 U9828 ( .A(n16061), .ZN(n11435) );
  AND2_X1 U9829 ( .A1(n9748), .A2(n10395), .ZN(n9749) );
  AND2_X1 U9830 ( .A1(n14168), .A2(n16103), .ZN(n9745) );
  NAND2_X1 U9831 ( .A1(n12596), .A2(n12600), .ZN(n13178) );
  AND2_X1 U9832 ( .A1(n9753), .A2(n10080), .ZN(n16053) );
  NAND2_X1 U9833 ( .A1(n9882), .A2(n10129), .ZN(n16056) );
  AND2_X1 U9834 ( .A1(n9181), .A2(n9180), .ZN(n9607) );
  AND2_X1 U9835 ( .A1(n9166), .A2(n9165), .ZN(n9487) );
  AND2_X1 U9836 ( .A1(n9157), .A2(n9156), .ZN(n9430) );
  INV_X1 U9837 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n14534) );
  CLKBUF_X3 U9838 ( .A(n11125), .Z(n14553) );
  OR2_X1 U9839 ( .A1(n12364), .A2(n12363), .ZN(n12365) );
  INV_X1 U9840 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n14619) );
  NAND2_X1 U9841 ( .A1(n12298), .A2(n12299), .ZN(n12366) );
  INV_X1 U9842 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n14660) );
  OR2_X1 U9843 ( .A1(n13490), .A2(n14660), .ZN(n13501) );
  NAND2_X1 U9844 ( .A1(n13887), .A2(n13886), .ZN(n13888) );
  OR2_X1 U9845 ( .A1(n12512), .A2(n12511), .ZN(n12540) );
  AND2_X1 U9846 ( .A1(n10545), .A2(n15058), .ZN(n10554) );
  INV_X1 U9847 ( .A(n14678), .ZN(n12587) );
  INV_X1 U9848 ( .A(n13629), .ZN(n11781) );
  AND2_X1 U9849 ( .A1(n10357), .A2(n13904), .ZN(n15026) );
  INV_X1 U9850 ( .A(n14924), .ZN(n14821) );
  AND2_X1 U9851 ( .A1(n15066), .A2(n10336), .ZN(n15643) );
  OR2_X1 U9852 ( .A1(n15066), .A2(n10352), .ZN(n10353) );
  NAND2_X1 U9853 ( .A1(n11653), .A2(n11654), .ZN(n11655) );
  INV_X1 U9854 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n15086) );
  INV_X1 U9855 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8619) );
  AND2_X1 U9856 ( .A1(n8897), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8880) );
  INV_X1 U9857 ( .A(n13258), .ZN(n11815) );
  OR2_X1 U9858 ( .A1(n8687), .A2(n8542), .ZN(n8668) );
  OR2_X1 U9859 ( .A1(n10526), .A2(n15583), .ZN(n10527) );
  AND2_X1 U9860 ( .A1(n8851), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n8594) );
  AND2_X1 U9861 ( .A1(n8869), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8851) );
  INV_X1 U9862 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n12392) );
  INV_X1 U9863 ( .A(n15274), .ZN(n15480) );
  XNOR2_X1 U9864 ( .A(n15288), .B(n15171), .ZN(n15280) );
  INV_X1 U9865 ( .A(n16321), .ZN(n12699) );
  INV_X1 U9866 ( .A(n12484), .ZN(n16224) );
  INV_X1 U9867 ( .A(n16333), .ZN(n16278) );
  INV_X1 U9868 ( .A(n16247), .ZN(n16198) );
  AND3_X1 U9869 ( .A1(n10870), .A2(n10869), .A3(n10868), .ZN(n10871) );
  NAND2_X1 U9870 ( .A1(n8475), .A2(n8474), .ZN(n8560) );
  AOI21_X1 U9871 ( .B1(n15830), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n8361), .ZN(
        n15832) );
  OR2_X1 U9872 ( .A1(n10395), .A2(n10127), .ZN(n10217) );
  NAND2_X1 U9873 ( .A1(n9884), .A2(n9883), .ZN(n14015) );
  NAND2_X1 U9874 ( .A1(n9827), .A2(n9826), .ZN(n13982) );
  NAND2_X1 U9875 ( .A1(n9838), .A2(n9837), .ZN(n14000) );
  NAND2_X1 U9876 ( .A1(n10252), .A2(n9798), .ZN(n12641) );
  NAND2_X1 U9877 ( .A1(n9879), .A2(n9878), .ZN(n14023) );
  AND2_X1 U9878 ( .A1(n9912), .A2(n9911), .ZN(n14158) );
  AND2_X1 U9879 ( .A1(n9644), .A2(n9643), .ZN(n14252) );
  INV_X1 U9880 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n12403) );
  INV_X1 U9881 ( .A(n15997), .ZN(n16020) );
  AND2_X1 U9882 ( .A1(P3_U3897), .A2(n13248), .ZN(n16017) );
  INV_X1 U9883 ( .A(n16056), .ZN(n14304) );
  INV_X1 U9884 ( .A(n14337), .ZN(n16096) );
  AND2_X1 U9885 ( .A1(n16100), .A2(n16088), .ZN(n14339) );
  AND2_X1 U9886 ( .A1(n11614), .A2(n9927), .ZN(n16061) );
  INV_X1 U9887 ( .A(n14418), .ZN(n12441) );
  NAND2_X1 U9888 ( .A1(n9755), .A2(n11767), .ZN(n16231) );
  INV_X1 U9889 ( .A(n16054), .ZN(n14384) );
  NAND2_X1 U9890 ( .A1(n14256), .A2(n14365), .ZN(n16103) );
  INV_X1 U9891 ( .A(n16231), .ZN(n16102) );
  INV_X1 U9892 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n9256) );
  AND2_X1 U9893 ( .A1(n9151), .A2(n9150), .ZN(n9398) );
  AND2_X1 U9894 ( .A1(n10542), .A2(n10541), .ZN(n10544) );
  NOR2_X1 U9895 ( .A1(n10369), .A2(n15649), .ZN(n10364) );
  AND3_X1 U9896 ( .A1(n13526), .A2(n13525), .A3(n13524), .ZN(n13866) );
  INV_X1 U9897 ( .A(n7425), .ZN(n13612) );
  INV_X1 U9898 ( .A(n15724), .ZN(n15741) );
  AND2_X1 U9899 ( .A1(n10554), .A2(n13906), .ZN(n15718) );
  AND2_X1 U9900 ( .A1(n10554), .A2(n15064), .ZN(n15743) );
  INV_X1 U9901 ( .A(n7415), .ZN(n15711) );
  AND2_X1 U9902 ( .A1(n12182), .A2(n12106), .ZN(n12352) );
  INV_X1 U9903 ( .A(n14936), .ZN(n14846) );
  INV_X1 U9904 ( .A(n14891), .ZN(n14870) );
  INV_X1 U9905 ( .A(n14933), .ZN(n14908) );
  INV_X1 U9906 ( .A(n15026), .ZN(n16307) );
  INV_X1 U9907 ( .A(n14998), .ZN(n16310) );
  AND2_X1 U9908 ( .A1(n13243), .A2(n10356), .ZN(n15647) );
  AND2_X1 U9909 ( .A1(n10724), .A2(n11220), .ZN(n15717) );
  NOR2_X1 U9910 ( .A1(n10431), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15059) );
  OR2_X1 U9911 ( .A1(n8635), .A2(n8619), .ZN(n8621) );
  INV_X1 U9912 ( .A(n16361), .ZN(n15167) );
  OAI21_X2 U9913 ( .B1(n10527), .B2(n16174), .A(n16110), .ZN(n15173) );
  AND3_X1 U9914 ( .A1(n8384), .A2(n8383), .A3(n8382), .ZN(n15252) );
  AND4_X1 U9915 ( .A1(n8575), .A2(n8574), .A3(n8573), .A4(n8572), .ZN(n15097)
         );
  INV_X1 U9916 ( .A(n8925), .ZN(n8872) );
  INV_X1 U9917 ( .A(n15240), .ZN(n15776) );
  INV_X1 U9918 ( .A(n15778), .ZN(n15765) );
  AND2_X1 U9919 ( .A1(n9116), .A2(n10804), .ZN(n15455) );
  INV_X1 U9920 ( .A(n15408), .ZN(n15457) );
  INV_X1 U9921 ( .A(n12648), .ZN(n12659) );
  INV_X1 U9922 ( .A(n16181), .ZN(n16269) );
  INV_X1 U9923 ( .A(n15435), .ZN(n16270) );
  AND2_X1 U9924 ( .A1(n10522), .A2(n15586), .ZN(n10891) );
  AND2_X1 U9925 ( .A1(n10883), .A2(n10882), .ZN(n16280) );
  INV_X1 U9926 ( .A(n16280), .ZN(n16330) );
  INV_X1 U9927 ( .A(n16299), .ZN(n16337) );
  INV_X1 U9928 ( .A(n16135), .ZN(n16257) );
  OR2_X1 U9929 ( .A1(n10954), .A2(P1_U3086), .ZN(n15583) );
  AND2_X1 U9930 ( .A1(n10454), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13236) );
  NOR2_X1 U9931 ( .A1(n8631), .A2(n8630), .ZN(n12627) );
  AND2_X1 U9932 ( .A1(n8708), .A2(n8707), .ZN(n11175) );
  AND2_X1 U9933 ( .A1(n10217), .A2(n10216), .ZN(n15646) );
  INV_X1 U9934 ( .A(n9890), .ZN(n9891) );
  NAND2_X1 U9935 ( .A1(n9868), .A2(n9867), .ZN(n14017) );
  INV_X1 U9936 ( .A(n14023), .ZN(n14036) );
  AND2_X1 U9937 ( .A1(n9912), .A2(n9723), .ZN(n11792) );
  INV_X1 U9938 ( .A(n14252), .ZN(n14223) );
  INV_X1 U9939 ( .A(n12601), .ZN(n14049) );
  INV_X1 U9940 ( .A(P3_U3897), .ZN(n14055) );
  MUX2_X1 U9941 ( .A(n10215), .B(n14055), .S(n10214), .Z(n15997) );
  NAND2_X1 U9942 ( .A1(n10162), .A2(n10134), .ZN(n16009) );
  NAND2_X1 U9943 ( .A1(n10401), .A2(n16059), .ZN(n16100) );
  INV_X1 U9944 ( .A(n14339), .ZN(n14288) );
  AND2_X1 U9945 ( .A1(n9763), .A2(n9762), .ZN(n9766) );
  INV_X1 U9946 ( .A(n14227), .ZN(n14436) );
  AND2_X1 U9947 ( .A1(n9266), .A2(n9265), .ZN(n16239) );
  NAND2_X1 U9948 ( .A1(n9230), .A2(n14467), .ZN(n10645) );
  AND2_X1 U9949 ( .A1(n9243), .A2(n9242), .ZN(n14466) );
  INV_X1 U9950 ( .A(n10164), .ZN(n14141) );
  NOR2_X1 U9951 ( .A1(n10431), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14474) );
  INV_X1 U9952 ( .A(SI_17_), .ZN(n12737) );
  INV_X1 U9953 ( .A(SI_12_), .ZN(n12970) );
  INV_X1 U9954 ( .A(n10187), .ZN(n11024) );
  AND2_X1 U9955 ( .A1(n10544), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15683) );
  INV_X1 U9956 ( .A(n14627), .ZN(n14663) );
  INV_X1 U9957 ( .A(n15718), .ZN(n15736) );
  INV_X1 U9958 ( .A(n15743), .ZN(n15728) );
  INV_X1 U9959 ( .A(n16293), .ZN(n16314) );
  AND2_X2 U9960 ( .A1(n10978), .A2(n15648), .ZN(n16293) );
  OR3_X1 U9961 ( .A1(n15016), .A2(n15015), .A3(n15014), .ZN(n15048) );
  NAND2_X1 U9962 ( .A1(n15647), .A2(n15644), .ZN(n15645) );
  INV_X1 U9963 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13617) );
  INV_X1 U9964 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n13388) );
  INV_X1 U9965 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n11735) );
  INV_X1 U9966 ( .A(n16266), .ZN(n16249) );
  INV_X1 U9967 ( .A(n15334), .ZN(n15503) );
  INV_X1 U9968 ( .A(n16277), .ZN(n12693) );
  INV_X1 U9969 ( .A(n15173), .ZN(n16353) );
  INV_X1 U9970 ( .A(n13599), .ZN(n15179) );
  INV_X1 U9971 ( .A(n15097), .ZN(n15374) );
  OR2_X1 U9972 ( .A1(n8624), .A2(n8623), .ZN(n16322) );
  INV_X1 U9973 ( .A(n11074), .ZN(n15195) );
  INV_X1 U9974 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15922) );
  OR2_X1 U9975 ( .A1(n16275), .A2(n16174), .ZN(n16114) );
  OR2_X1 U9976 ( .A1(n16264), .A2(n16280), .ZN(n15462) );
  INV_X1 U9977 ( .A(n16179), .ZN(n16275) );
  AND2_X1 U9978 ( .A1(n10880), .A2(n8799), .ZN(n16033) );
  INV_X1 U9979 ( .A(n16341), .ZN(n16339) );
  AND4_X1 U9980 ( .A1(n16186), .A2(n16167), .A3(n16182), .A4(n16166), .ZN(
        n16169) );
  INV_X1 U9981 ( .A(n16345), .ZN(n16342) );
  NOR2_X1 U9982 ( .A1(n15584), .A2(n15583), .ZN(n15625) );
  CLKBUF_X1 U9983 ( .A(n15625), .Z(n15640) );
  INV_X1 U9984 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n13246) );
  INV_X1 U9985 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n11768) );
  INV_X1 U9986 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10655) );
  AND2_X2 U9987 ( .A1(n10106), .A2(n14467), .ZN(P3_U3897) );
  OR4_X1 U9988 ( .A1(n10223), .A2(n10222), .A3(n10221), .A4(n10220), .ZN(
        P3_U3196) );
  AND2_X1 U9989 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10538), .ZN(P2_U3947) );
  INV_X1 U9990 ( .A(n15196), .ZN(P1_U4016) );
  NAND3_X1 U9991 ( .A1(n7673), .A2(n9100), .A3(n8373), .ZN(n9105) );
  NOR2_X1 U9992 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n8375) );
  NOR2_X1 U9993 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n8374) );
  XNOR2_X2 U9994 ( .A(n8783), .B(n8790), .ZN(n8381) );
  XNOR2_X2 U9995 ( .A(n8379), .B(P1_IR_REG_29__SCAN_IN), .ZN(n8795) );
  NAND2_X1 U9996 ( .A1(n8922), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n8384) );
  AND2_X2 U9997 ( .A1(n8540), .A2(n8380), .ZN(n8763) );
  NAND2_X1 U9998 ( .A1(n8926), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n8383) );
  NAND2_X1 U9999 ( .A1(n8921), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8382) );
  INV_X1 U10000 ( .A(n15252), .ZN(n15177) );
  NAND2_X1 U10001 ( .A1(n8510), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8385) );
  MUX2_X1 U10002 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8385), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n8386) );
  INV_X1 U10003 ( .A(n8922), .ZN(n8855) );
  INV_X1 U10004 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8389) );
  NAND2_X1 U10005 ( .A1(n8926), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8388) );
  NAND2_X1 U10006 ( .A1(n8921), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8387) );
  OAI211_X1 U10007 ( .C1(n8855), .C2(n8389), .A(n8388), .B(n8387), .ZN(n15178)
         );
  OAI21_X1 U10008 ( .B1(n15177), .B2(n12527), .A(n15178), .ZN(n8390) );
  INV_X1 U10009 ( .A(n8390), .ZN(n8519) );
  INV_X1 U10010 ( .A(SI_1_), .ZN(n12989) );
  NAND2_X1 U10011 ( .A1(n10464), .A2(n12989), .ZN(n8395) );
  AND2_X1 U10012 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n8768) );
  AOI22_X1 U10013 ( .A1(n8395), .A2(n8768), .B1(P2_DATAO_REG_1__SCAN_IN), .B2(
        SI_1_), .ZN(n8401) );
  NOR2_X1 U10014 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8398) );
  AND2_X1 U10015 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8769) );
  INV_X1 U10016 ( .A(n8769), .ZN(n8397) );
  NAND2_X1 U10017 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8396) );
  OAI21_X1 U10018 ( .B1(n8398), .B2(n8397), .A(n8396), .ZN(n8399) );
  NAND2_X1 U10019 ( .A1(n8767), .A2(n8399), .ZN(n8400) );
  OAI21_X2 U10020 ( .B1(n8767), .B2(n8401), .A(n8400), .ZN(n8402) );
  INV_X1 U10021 ( .A(SI_2_), .ZN(n12761) );
  MUX2_X1 U10022 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n8767), .Z(n8746) );
  NAND2_X1 U10023 ( .A1(n8747), .A2(n8746), .ZN(n8404) );
  NAND2_X1 U10024 ( .A1(n8402), .A2(SI_2_), .ZN(n8403) );
  MUX2_X1 U10025 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n8767), .Z(n8405) );
  INV_X1 U10026 ( .A(SI_3_), .ZN(n10440) );
  XNOR2_X1 U10027 ( .A(n8405), .B(n10440), .ZN(n8755) );
  NAND2_X1 U10028 ( .A1(n8756), .A2(n8755), .ZN(n8407) );
  NAND2_X1 U10029 ( .A1(n8405), .A2(SI_3_), .ZN(n8406) );
  NAND2_X1 U10030 ( .A1(n8407), .A2(n8406), .ZN(n8806) );
  MUX2_X1 U10031 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n8767), .Z(n8409) );
  XNOR2_X1 U10032 ( .A(n8409), .B(SI_4_), .ZN(n8805) );
  INV_X1 U10033 ( .A(n8805), .ZN(n8408) );
  NAND2_X1 U10034 ( .A1(n8806), .A2(n8408), .ZN(n8411) );
  NAND2_X1 U10035 ( .A1(n8409), .A2(SI_4_), .ZN(n8410) );
  NAND2_X2 U10036 ( .A1(n8411), .A2(n8410), .ZN(n8812) );
  MUX2_X1 U10037 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n8767), .Z(n8415) );
  XNOR2_X1 U10038 ( .A(n8415), .B(SI_5_), .ZN(n8813) );
  INV_X1 U10039 ( .A(n8813), .ZN(n8824) );
  NAND2_X1 U10040 ( .A1(n8412), .A2(SI_6_), .ZN(n8416) );
  XNOR2_X1 U10041 ( .A(n8412), .B(SI_6_), .ZN(n8827) );
  AND2_X1 U10042 ( .A1(n8414), .A2(n8824), .ZN(n8413) );
  INV_X1 U10043 ( .A(n8414), .ZN(n8418) );
  NAND2_X1 U10044 ( .A1(n8415), .A2(SI_5_), .ZN(n8825) );
  AND2_X1 U10045 ( .A1(n8825), .A2(n8416), .ZN(n8417) );
  MUX2_X1 U10046 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n8767), .Z(n8421) );
  XNOR2_X1 U10047 ( .A(n8421), .B(SI_7_), .ZN(n8726) );
  INV_X1 U10048 ( .A(n8726), .ZN(n8420) );
  NAND2_X1 U10049 ( .A1(n8421), .A2(SI_7_), .ZN(n8422) );
  MUX2_X1 U10050 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n10431), .Z(n8424) );
  XNOR2_X1 U10051 ( .A(n8424), .B(SI_8_), .ZN(n8715) );
  INV_X1 U10052 ( .A(n8715), .ZN(n8423) );
  NAND2_X1 U10053 ( .A1(n8716), .A2(n8423), .ZN(n8426) );
  NAND2_X1 U10054 ( .A1(n8424), .A2(SI_8_), .ZN(n8425) );
  MUX2_X1 U10055 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n10432), .Z(n8704) );
  MUX2_X1 U10056 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n10432), .Z(n8429) );
  MUX2_X1 U10057 ( .A(n10503), .B(n10501), .S(n10431), .Z(n8430) );
  NAND2_X1 U10058 ( .A1(n8430), .A2(n12973), .ZN(n8433) );
  INV_X1 U10059 ( .A(n8430), .ZN(n8431) );
  NAND2_X1 U10060 ( .A1(n8431), .A2(SI_11_), .ZN(n8432) );
  NAND2_X1 U10061 ( .A1(n8433), .A2(n8432), .ZN(n8681) );
  MUX2_X1 U10062 ( .A(n10655), .B(n10653), .S(n10432), .Z(n8434) );
  NAND2_X1 U10063 ( .A1(n8434), .A2(n12970), .ZN(n8437) );
  INV_X1 U10064 ( .A(n8434), .ZN(n8435) );
  NAND2_X1 U10065 ( .A1(n8435), .A2(SI_12_), .ZN(n8436) );
  MUX2_X1 U10066 ( .A(n10727), .B(n10725), .S(n10431), .Z(n8438) );
  XNOR2_X1 U10067 ( .A(n8438), .B(SI_13_), .ZN(n8659) );
  INV_X1 U10068 ( .A(n8659), .ZN(n8441) );
  INV_X1 U10069 ( .A(n8438), .ZN(n8439) );
  NAND2_X1 U10070 ( .A1(n8439), .A2(SI_13_), .ZN(n8440) );
  MUX2_X1 U10071 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n10431), .Z(n8641) );
  MUX2_X1 U10072 ( .A(n11289), .B(n11294), .S(n10432), .Z(n8444) );
  NAND2_X1 U10073 ( .A1(n8444), .A2(n10936), .ZN(n8447) );
  INV_X1 U10074 ( .A(n8444), .ZN(n8445) );
  NAND2_X1 U10075 ( .A1(n8445), .A2(SI_15_), .ZN(n8446) );
  NAND2_X1 U10076 ( .A1(n8447), .A2(n8446), .ZN(n8625) );
  MUX2_X1 U10077 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(P1_DATAO_REG_16__SCAN_IN), 
        .S(n10432), .Z(n8612) );
  INV_X1 U10078 ( .A(n8612), .ZN(n8448) );
  MUX2_X1 U10079 ( .A(n11768), .B(n11775), .S(n10432), .Z(n8451) );
  NAND2_X1 U10080 ( .A1(n8451), .A2(n12737), .ZN(n8454) );
  INV_X1 U10081 ( .A(n8451), .ZN(n8452) );
  NAND2_X1 U10082 ( .A1(n8452), .A2(SI_17_), .ZN(n8453) );
  NAND2_X1 U10083 ( .A1(n8454), .A2(n8453), .ZN(n8600) );
  MUX2_X1 U10084 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n10432), .Z(n8858) );
  MUX2_X1 U10085 ( .A(n13252), .B(n9578), .S(n10431), .Z(n8457) );
  INV_X1 U10086 ( .A(n8457), .ZN(n8458) );
  NAND2_X1 U10087 ( .A1(n8458), .A2(SI_19_), .ZN(n8459) );
  NAND2_X1 U10088 ( .A1(n8460), .A2(n8459), .ZN(n8845) );
  OAI21_X2 U10089 ( .B1(n8846), .B2(n8845), .A(n8460), .ZN(n8590) );
  MUX2_X1 U10090 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n10432), .Z(n8588) );
  MUX2_X1 U10091 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n10431), .Z(n8462) );
  XNOR2_X1 U10092 ( .A(n8462), .B(SI_21_), .ZN(n8576) );
  INV_X1 U10093 ( .A(n8576), .ZN(n8461) );
  NAND2_X1 U10094 ( .A1(n8462), .A2(SI_21_), .ZN(n8463) );
  MUX2_X1 U10095 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n10432), .Z(n13253) );
  MUX2_X1 U10096 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n10432), .Z(n8891) );
  INV_X1 U10097 ( .A(n8891), .ZN(n8465) );
  INV_X1 U10098 ( .A(SI_23_), .ZN(n11955) );
  NAND2_X1 U10099 ( .A1(n8465), .A2(n11955), .ZN(n8468) );
  OAI21_X1 U10100 ( .B1(SI_22_), .B2(n13253), .A(n8468), .ZN(n8466) );
  INV_X1 U10101 ( .A(n8466), .ZN(n8467) );
  NAND2_X1 U10102 ( .A1(n8887), .A2(n8467), .ZN(n8471) );
  INV_X1 U10103 ( .A(n13253), .ZN(n8889) );
  INV_X1 U10104 ( .A(SI_22_), .ZN(n9621) );
  NOR2_X1 U10105 ( .A1(n8889), .A2(n9621), .ZN(n8469) );
  AOI22_X1 U10106 ( .A1(n8469), .A2(n8468), .B1(n8891), .B2(SI_23_), .ZN(n8470) );
  NAND2_X1 U10107 ( .A1(n8471), .A2(n8470), .ZN(n8473) );
  INV_X1 U10108 ( .A(n8877), .ZN(n8472) );
  MUX2_X1 U10109 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n10431), .Z(n8876) );
  NAND2_X1 U10110 ( .A1(n8472), .A2(n8876), .ZN(n8475) );
  NAND2_X1 U10111 ( .A1(n8473), .A2(SI_24_), .ZN(n8474) );
  INV_X1 U10112 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n9191) );
  INV_X1 U10113 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n15073) );
  MUX2_X1 U10114 ( .A(n9191), .B(n15073), .S(n10432), .Z(n8476) );
  INV_X1 U10115 ( .A(SI_25_), .ZN(n12724) );
  NAND2_X1 U10116 ( .A1(n8476), .A2(n12724), .ZN(n8479) );
  INV_X1 U10117 ( .A(n8476), .ZN(n8477) );
  NAND2_X1 U10118 ( .A1(n8477), .A2(SI_25_), .ZN(n8478) );
  NAND2_X1 U10119 ( .A1(n8479), .A2(n8478), .ZN(n8559) );
  INV_X1 U10120 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n15598) );
  INV_X1 U10121 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n15068) );
  MUX2_X1 U10122 ( .A(n15598), .B(n15068), .S(n10431), .Z(n8481) );
  XNOR2_X1 U10123 ( .A(n8481), .B(SI_26_), .ZN(n8549) );
  INV_X1 U10124 ( .A(n8549), .ZN(n8480) );
  INV_X1 U10125 ( .A(n8481), .ZN(n8482) );
  NAND2_X1 U10126 ( .A1(n8482), .A2(SI_26_), .ZN(n8483) );
  INV_X1 U10127 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n15596) );
  INV_X1 U10128 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n15065) );
  MUX2_X1 U10129 ( .A(n15596), .B(n15065), .S(n10432), .Z(n8484) );
  XNOR2_X1 U10130 ( .A(n8484), .B(SI_27_), .ZN(n8535) );
  INV_X1 U10131 ( .A(n8484), .ZN(n8485) );
  NAND2_X1 U10132 ( .A1(n8485), .A2(SI_27_), .ZN(n8486) );
  MUX2_X1 U10133 ( .A(n13246), .B(n13373), .S(n10432), .Z(n8488) );
  INV_X1 U10134 ( .A(SI_28_), .ZN(n13249) );
  NAND2_X1 U10135 ( .A1(n8488), .A2(n13249), .ZN(n8491) );
  INV_X1 U10136 ( .A(n8488), .ZN(n8489) );
  NAND2_X1 U10137 ( .A1(n8489), .A2(SI_28_), .ZN(n8490) );
  NAND2_X1 U10138 ( .A1(n8491), .A2(n8490), .ZN(n8917) );
  INV_X1 U10139 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n15593) );
  INV_X1 U10140 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n15057) );
  MUX2_X1 U10141 ( .A(n15593), .B(n15057), .S(n10431), .Z(n8492) );
  INV_X1 U10142 ( .A(SI_29_), .ZN(n13925) );
  NAND2_X1 U10143 ( .A1(n8492), .A2(n13925), .ZN(n8496) );
  INV_X1 U10144 ( .A(n8492), .ZN(n8493) );
  NAND2_X1 U10145 ( .A1(n8493), .A2(SI_29_), .ZN(n8494) );
  NAND2_X1 U10146 ( .A1(n8496), .A2(n8494), .ZN(n8906) );
  INV_X1 U10147 ( .A(n8906), .ZN(n8495) );
  INV_X1 U10148 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n13604) );
  MUX2_X1 U10149 ( .A(n13604), .B(n13617), .S(n10432), .Z(n8522) );
  XNOR2_X1 U10150 ( .A(n8522), .B(SI_30_), .ZN(n8521) );
  NAND2_X1 U10151 ( .A1(n13616), .A2(n7428), .ZN(n8503) );
  NAND2_X1 U10152 ( .A1(n8758), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8502) );
  NAND2_X2 U10153 ( .A1(n8503), .A2(n8502), .ZN(n15257) );
  NOR2_X2 U10154 ( .A1(n8508), .A2(n8507), .ZN(n9108) );
  NAND2_X1 U10155 ( .A1(n8510), .A2(n8509), .ZN(n8516) );
  INV_X1 U10156 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8512) );
  INV_X1 U10157 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8511) );
  NAND3_X1 U10158 ( .A1(n8512), .A2(n8511), .A3(P1_IR_REG_22__SCAN_IN), .ZN(
        n8514) );
  XNOR2_X1 U10159 ( .A(P1_IR_REG_22__SCAN_IN), .B(P1_IR_REG_31__SCAN_IN), .ZN(
        n8513) );
  NAND2_X1 U10160 ( .A1(n8514), .A2(n8513), .ZN(n8515) );
  INV_X1 U10161 ( .A(n15606), .ZN(n9098) );
  MUX2_X1 U10162 ( .A(n8519), .B(n15257), .S(n8948), .Z(n9121) );
  NAND2_X1 U10163 ( .A1(n9099), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8520) );
  NAND2_X1 U10164 ( .A1(n9121), .A2(n13236), .ZN(n9118) );
  INV_X1 U10165 ( .A(n8521), .ZN(n8525) );
  INV_X1 U10166 ( .A(n8522), .ZN(n8523) );
  NAND2_X1 U10167 ( .A1(n8523), .A2(SI_30_), .ZN(n8524) );
  OAI21_X1 U10168 ( .B1(n8526), .B2(n8525), .A(n8524), .ZN(n8529) );
  MUX2_X1 U10169 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n10432), .Z(n8527) );
  XNOR2_X1 U10170 ( .A(n8527), .B(SI_31_), .ZN(n8528) );
  XNOR2_X1 U10171 ( .A(n8529), .B(n8528), .ZN(n15051) );
  NAND2_X1 U10172 ( .A1(n15051), .A2(n7428), .ZN(n8531) );
  NAND2_X1 U10173 ( .A1(n8758), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8530) );
  NAND2_X2 U10174 ( .A1(n8531), .A2(n8530), .ZN(n15253) );
  NAND2_X1 U10175 ( .A1(n15177), .A2(n7427), .ZN(n8936) );
  OR2_X1 U10176 ( .A1(n10878), .A2(n15244), .ZN(n16170) );
  NAND2_X1 U10177 ( .A1(n10881), .A2(n15606), .ZN(n10529) );
  OAI21_X1 U10178 ( .B1(n15606), .B2(n8224), .A(n10529), .ZN(n8532) );
  NAND2_X1 U10179 ( .A1(n16170), .A2(n8532), .ZN(n9095) );
  INV_X1 U10180 ( .A(n10881), .ZN(n12593) );
  NAND2_X1 U10181 ( .A1(n12593), .A2(n8224), .ZN(n8939) );
  AND2_X1 U10182 ( .A1(n9095), .A2(n8939), .ZN(n9128) );
  OR2_X1 U10183 ( .A1(n15177), .A2(n7427), .ZN(n8937) );
  INV_X1 U10184 ( .A(n8937), .ZN(n8533) );
  NAND2_X1 U10185 ( .A1(n15253), .A2(n8533), .ZN(n8534) );
  OAI211_X1 U10186 ( .C1(n15253), .C2(n8936), .A(n9128), .B(n8534), .ZN(n9119)
         );
  XNOR2_X1 U10187 ( .A(n15253), .B(n15252), .ZN(n9131) );
  XNOR2_X1 U10188 ( .A(n15257), .B(n15178), .ZN(n8932) );
  INV_X1 U10189 ( .A(n8535), .ZN(n8536) );
  NAND2_X1 U10190 ( .A1(n15063), .A2(n7428), .ZN(n8539) );
  NAND2_X1 U10191 ( .A1(n8758), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8538) );
  AND2_X2 U10192 ( .A1(n8539), .A2(n8538), .ZN(n15485) );
  NAND2_X1 U10193 ( .A1(n8921), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8548) );
  NAND2_X1 U10194 ( .A1(n8922), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n8547) );
  AND2_X4 U10195 ( .A1(n8795), .A2(n8540), .ZN(n8925) );
  NAND2_X1 U10196 ( .A1(n8834), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8833) );
  NOR2_X1 U10197 ( .A1(n8833), .A2(n8732), .ZN(n8734) );
  NAND2_X1 U10198 ( .A1(n8721), .A2(n8541), .ZN(n8698) );
  NAND2_X1 U10199 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .ZN(n8542) );
  NAND2_X1 U10200 ( .A1(n8654), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8635) );
  NAND2_X1 U10201 ( .A1(n8594), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8580) );
  INV_X1 U10202 ( .A(n8580), .ZN(n8543) );
  NAND2_X1 U10203 ( .A1(n8543), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8898) );
  NAND2_X1 U10204 ( .A1(n8571), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8881) );
  NOR2_X1 U10205 ( .A1(n8554), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8544) );
  NOR2_X1 U10206 ( .A1(n8923), .A2(n8544), .ZN(n15287) );
  NAND2_X1 U10207 ( .A1(n8925), .A2(n15287), .ZN(n8546) );
  NAND2_X1 U10208 ( .A1(n8896), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8545) );
  NAND2_X1 U10209 ( .A1(n15067), .A2(n7428), .ZN(n8552) );
  NAND2_X1 U10210 ( .A1(n8758), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8551) );
  NAND2_X2 U10211 ( .A1(n8552), .A2(n8551), .ZN(n15491) );
  NAND2_X1 U10212 ( .A1(n8921), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8558) );
  NAND2_X1 U10213 ( .A1(n8922), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8557) );
  NOR2_X1 U10214 ( .A1(n8564), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8553) );
  NOR2_X1 U10215 ( .A1(n8554), .A2(n8553), .ZN(n15299) );
  NAND2_X1 U10216 ( .A1(n8925), .A2(n15299), .ZN(n8556) );
  NAND2_X1 U10217 ( .A1(n8926), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8555) );
  NAND4_X1 U10218 ( .A1(n8558), .A2(n8557), .A3(n8556), .A4(n8555), .ZN(n15312) );
  XNOR2_X1 U10219 ( .A(n15491), .B(n15312), .ZN(n15293) );
  XNOR2_X1 U10220 ( .A(n8560), .B(n8559), .ZN(n15070) );
  NAND2_X1 U10221 ( .A1(n15070), .A2(n7428), .ZN(n8562) );
  NAND2_X1 U10222 ( .A1(n8758), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8561) );
  NAND2_X1 U10223 ( .A1(n8922), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8568) );
  NAND2_X1 U10224 ( .A1(n8896), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8567) );
  NOR2_X1 U10225 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n8880), .ZN(n8563) );
  NOR2_X1 U10226 ( .A1(n8564), .A2(n8563), .ZN(n15315) );
  NAND2_X1 U10227 ( .A1(n8925), .A2(n15315), .ZN(n8566) );
  NAND2_X1 U10228 ( .A1(n8921), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8565) );
  NAND4_X1 U10229 ( .A1(n8568), .A2(n8567), .A3(n8566), .A4(n8565), .ZN(n15329) );
  NAND2_X1 U10230 ( .A1(n15498), .A2(n15329), .ZN(n13339) );
  OR2_X1 U10231 ( .A1(n15498), .A2(n15329), .ZN(n8569) );
  NAND2_X1 U10232 ( .A1(n13339), .A2(n8569), .ZN(n15321) );
  NAND2_X1 U10233 ( .A1(n8921), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8575) );
  NAND2_X1 U10234 ( .A1(n8922), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n8574) );
  INV_X1 U10235 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13321) );
  AOI21_X1 U10236 ( .B1(n13321), .B2(n8580), .A(n8571), .ZN(n15361) );
  NAND2_X1 U10237 ( .A1(n8925), .A2(n15361), .ZN(n8573) );
  NAND2_X1 U10238 ( .A1(n8896), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8572) );
  XNOR2_X1 U10239 ( .A(n15516), .B(n15097), .ZN(n13337) );
  XNOR2_X1 U10240 ( .A(n8577), .B(n8576), .ZN(n13432) );
  NAND2_X1 U10241 ( .A1(n13432), .A2(n7428), .ZN(n8579) );
  NAND2_X1 U10242 ( .A1(n8758), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8578) );
  NAND2_X2 U10243 ( .A1(n8579), .A2(n8578), .ZN(n15525) );
  OR2_X1 U10244 ( .A1(n8594), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8581) );
  AND2_X1 U10245 ( .A1(n8581), .A2(n8580), .ZN(n15380) );
  NAND2_X1 U10246 ( .A1(n15380), .A2(n8925), .ZN(n8587) );
  INV_X1 U10247 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n8584) );
  NAND2_X1 U10248 ( .A1(n8921), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8583) );
  NAND2_X1 U10249 ( .A1(n8926), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8582) );
  OAI211_X1 U10250 ( .C1(n8855), .C2(n8584), .A(n8583), .B(n8582), .ZN(n8585)
         );
  INV_X1 U10251 ( .A(n8585), .ZN(n8586) );
  NAND2_X1 U10252 ( .A1(n8587), .A2(n8586), .ZN(n15181) );
  INV_X1 U10253 ( .A(n15181), .ZN(n13364) );
  XNOR2_X1 U10254 ( .A(n15525), .B(n13364), .ZN(n15369) );
  XNOR2_X1 U10255 ( .A(n8588), .B(n11612), .ZN(n8589) );
  XNOR2_X1 U10256 ( .A(n8590), .B(n8589), .ZN(n13417) );
  NAND2_X1 U10257 ( .A1(n13417), .A2(n7428), .ZN(n8592) );
  NAND2_X1 U10258 ( .A1(n8758), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8591) );
  NOR2_X1 U10259 ( .A1(n8851), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n8593) );
  OR2_X1 U10260 ( .A1(n8594), .A2(n8593), .ZN(n15390) );
  INV_X1 U10261 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n8597) );
  NAND2_X1 U10262 ( .A1(n8896), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8596) );
  NAND2_X1 U10263 ( .A1(n8921), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n8595) );
  OAI211_X1 U10264 ( .C1(n8855), .C2(n8597), .A(n8596), .B(n8595), .ZN(n8598)
         );
  INV_X1 U10265 ( .A(n8598), .ZN(n8599) );
  XNOR2_X1 U10266 ( .A(n15528), .B(n15375), .ZN(n13336) );
  XNOR2_X1 U10267 ( .A(n8601), .B(n8600), .ZN(n12534) );
  NAND2_X1 U10268 ( .A1(n12534), .A2(n7428), .ZN(n8607) );
  OR2_X1 U10269 ( .A1(n8829), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n8728) );
  NAND4_X1 U10270 ( .A1(n8603), .A2(n8645), .A3(n8602), .A4(n8643), .ZN(n8604)
         );
  NOR2_X1 U10271 ( .A1(n8728), .A2(n8604), .ZN(n8627) );
  NAND2_X1 U10272 ( .A1(n8627), .A2(n13154), .ZN(n8629) );
  OR2_X1 U10273 ( .A1(n8629), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n8605) );
  NAND2_X1 U10274 ( .A1(n8605), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8861) );
  XNOR2_X1 U10275 ( .A(n8861), .B(P1_IR_REG_17__SCAN_IN), .ZN(n15216) );
  AOI22_X1 U10276 ( .A1(n8758), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n8864), 
        .B2(n15216), .ZN(n8606) );
  AND2_X1 U10277 ( .A1(n8621), .A2(n8608), .ZN(n8609) );
  OR2_X1 U10278 ( .A1(n8609), .A2(n8867), .ZN(n15439) );
  AOI22_X1 U10279 ( .A1(n8922), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n8921), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n8611) );
  NAND2_X1 U10280 ( .A1(n8926), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8610) );
  OAI211_X1 U10281 ( .C1(n15439), .C2(n8872), .A(n8611), .B(n8610), .ZN(n16350) );
  INV_X1 U10282 ( .A(n16350), .ZN(n15158) );
  XNOR2_X1 U10283 ( .A(n15550), .B(n15158), .ZN(n15443) );
  XNOR2_X1 U10284 ( .A(n8613), .B(n8612), .ZN(n12507) );
  NAND2_X1 U10285 ( .A1(n12507), .A2(n7428), .ZN(n8616) );
  NAND2_X1 U10286 ( .A1(n8629), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8614) );
  XNOR2_X1 U10287 ( .A(n8614), .B(P1_IR_REG_16__SCAN_IN), .ZN(n15206) );
  AOI22_X1 U10288 ( .A1(n8758), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n8864), 
        .B2(n15206), .ZN(n8615) );
  INV_X1 U10289 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n8618) );
  NAND2_X1 U10290 ( .A1(n8921), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n8617) );
  OAI21_X1 U10291 ( .B1(n8618), .B2(n8750), .A(n8617), .ZN(n8624) );
  NAND2_X1 U10292 ( .A1(n8635), .A2(n8619), .ZN(n8620) );
  NAND2_X1 U10293 ( .A1(n8621), .A2(n8620), .ZN(n16360) );
  INV_X1 U10294 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n8622) );
  OAI22_X1 U10295 ( .A1(n16360), .A2(n8872), .B1(n8855), .B2(n8622), .ZN(n8623) );
  INV_X1 U10296 ( .A(n16322), .ZN(n13357) );
  XNOR2_X1 U10297 ( .A(n15454), .B(n13357), .ZN(n15461) );
  XNOR2_X1 U10298 ( .A(n8626), .B(n8625), .ZN(n12413) );
  NAND2_X1 U10299 ( .A1(n12413), .A2(n7428), .ZN(n8633) );
  NOR2_X1 U10300 ( .A1(n8627), .A2(n7671), .ZN(n8628) );
  MUX2_X1 U10301 ( .A(n7671), .B(n8628), .S(P1_IR_REG_15__SCAN_IN), .Z(n8631)
         );
  INV_X1 U10302 ( .A(n8629), .ZN(n8630) );
  AOI22_X1 U10303 ( .A1(n8758), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n8864), 
        .B2(n12627), .ZN(n8632) );
  NAND2_X1 U10304 ( .A1(n8922), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n8640) );
  OR2_X1 U10305 ( .A1(n8654), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8634) );
  NAND2_X1 U10306 ( .A1(n8635), .A2(n8634), .ZN(n16328) );
  INV_X1 U10307 ( .A(n16328), .ZN(n8636) );
  NAND2_X1 U10308 ( .A1(n8925), .A2(n8636), .ZN(n8639) );
  NAND2_X1 U10309 ( .A1(n8896), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n8638) );
  NAND2_X1 U10310 ( .A1(n8921), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n8637) );
  NAND4_X1 U10311 ( .A1(n8640), .A2(n8639), .A3(n8638), .A4(n8637), .ZN(n16348) );
  INV_X1 U10312 ( .A(n16348), .ZN(n13353) );
  XNOR2_X1 U10313 ( .A(n13354), .B(n13353), .ZN(n12702) );
  XNOR2_X1 U10314 ( .A(n8642), .B(n8641), .ZN(n12211) );
  NAND2_X1 U10315 ( .A1(n12211), .A2(n7428), .ZN(n8652) );
  OAI21_X1 U10316 ( .B1(n8728), .B2(P1_IR_REG_7__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8717) );
  NAND2_X1 U10317 ( .A1(n8717), .A2(n8643), .ZN(n8644) );
  NAND2_X1 U10318 ( .A1(n8644), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8706) );
  OR2_X1 U10319 ( .A1(n8645), .A2(n7671), .ZN(n8646) );
  NAND2_X1 U10320 ( .A1(n8706), .A2(n8646), .ZN(n8683) );
  NAND2_X1 U10321 ( .A1(n8647), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8674) );
  NAND2_X1 U10322 ( .A1(n8674), .A2(n13147), .ZN(n8648) );
  NAND2_X1 U10323 ( .A1(n8648), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8661) );
  INV_X1 U10324 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n13148) );
  NAND2_X1 U10325 ( .A1(n8661), .A2(n13148), .ZN(n8649) );
  NAND2_X1 U10326 ( .A1(n8649), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8650) );
  XNOR2_X1 U10327 ( .A(n8650), .B(P1_IR_REG_14__SCAN_IN), .ZN(n12619) );
  AOI22_X1 U10328 ( .A1(n12619), .A2(n8864), .B1(n8758), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n8651) );
  NAND2_X1 U10329 ( .A1(n8922), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n8658) );
  NAND2_X1 U10330 ( .A1(n8921), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n8657) );
  AND2_X1 U10331 ( .A1(n8668), .A2(n15086), .ZN(n8653) );
  NOR2_X1 U10332 ( .A1(n8654), .A2(n8653), .ZN(n15088) );
  NAND2_X1 U10333 ( .A1(n8925), .A2(n15088), .ZN(n8656) );
  NAND2_X1 U10334 ( .A1(n8896), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n8655) );
  NAND4_X1 U10335 ( .A1(n8658), .A2(n8657), .A3(n8656), .A4(n8655), .ZN(n16321) );
  XNOR2_X1 U10336 ( .A(n15089), .B(n12699), .ZN(n12650) );
  XNOR2_X1 U10337 ( .A(n8660), .B(n8659), .ZN(n12183) );
  NAND2_X1 U10338 ( .A1(n12183), .A2(n7428), .ZN(n8664) );
  XNOR2_X1 U10339 ( .A(n8661), .B(P1_IR_REG_13__SCAN_IN), .ZN(n12081) );
  NOR2_X1 U10340 ( .A1(n8773), .A2(n10727), .ZN(n8662) );
  AOI21_X1 U10341 ( .B1(n12081), .B2(n8864), .A(n8662), .ZN(n8663) );
  NAND2_X1 U10342 ( .A1(n8922), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8672) );
  NAND2_X1 U10343 ( .A1(n8926), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n8671) );
  INV_X1 U10344 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n8666) );
  INV_X1 U10345 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8665) );
  OAI21_X1 U10346 ( .B1(n8687), .B2(n8666), .A(n8665), .ZN(n8667) );
  AND2_X1 U10347 ( .A1(n8668), .A2(n8667), .ZN(n12690) );
  NAND2_X1 U10348 ( .A1(n8925), .A2(n12690), .ZN(n8670) );
  NAND2_X1 U10349 ( .A1(n8921), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n8669) );
  NAND4_X1 U10350 ( .A1(n8672), .A2(n8671), .A3(n8670), .A4(n8669), .ZN(n15183) );
  INV_X1 U10351 ( .A(n15183), .ZN(n12681) );
  XNOR2_X1 U10352 ( .A(n16277), .B(n12681), .ZN(n12648) );
  XNOR2_X1 U10353 ( .A(n8673), .B(n8366), .ZN(n12101) );
  NAND2_X1 U10354 ( .A1(n12101), .A2(n7428), .ZN(n8676) );
  XNOR2_X1 U10355 ( .A(n8674), .B(P1_IR_REG_12__SCAN_IN), .ZN(n15779) );
  AOI22_X1 U10356 ( .A1(n8864), .A2(n15779), .B1(n8758), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n8675) );
  NAND2_X1 U10357 ( .A1(n8921), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n8680) );
  NAND2_X1 U10358 ( .A1(n8922), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n8679) );
  XNOR2_X1 U10359 ( .A(n8687), .B(P1_REG3_REG_12__SCAN_IN), .ZN(n16263) );
  NAND2_X1 U10360 ( .A1(n8925), .A2(n16263), .ZN(n8678) );
  NAND2_X1 U10361 ( .A1(n8926), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n8677) );
  NAND4_X1 U10362 ( .A1(n8680), .A2(n8679), .A3(n8678), .A4(n8677), .ZN(n15184) );
  XNOR2_X1 U10363 ( .A(n16266), .B(n12687), .ZN(n12486) );
  XNOR2_X1 U10364 ( .A(n8682), .B(n8681), .ZN(n12020) );
  NAND2_X1 U10365 ( .A1(n12020), .A2(n7428), .ZN(n8685) );
  INV_X1 U10366 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n12923) );
  XNOR2_X1 U10367 ( .A(n8683), .B(n12923), .ZN(n11711) );
  AOI22_X1 U10368 ( .A1(n8758), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n8864), 
        .B2(n11711), .ZN(n8684) );
  NAND2_X1 U10369 ( .A1(n8685), .A2(n8684), .ZN(n12484) );
  NAND2_X1 U10370 ( .A1(n8921), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n8691) );
  NAND2_X1 U10371 ( .A1(n8922), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n8690) );
  NAND2_X1 U10372 ( .A1(n8698), .A2(n12392), .ZN(n8686) );
  AND2_X1 U10373 ( .A1(n8687), .A2(n8686), .ZN(n12395) );
  NAND2_X1 U10374 ( .A1(n8925), .A2(n12395), .ZN(n8689) );
  NAND2_X1 U10375 ( .A1(n8896), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n8688) );
  NAND4_X1 U10376 ( .A1(n8691), .A2(n8690), .A3(n8689), .A4(n8688), .ZN(n15185) );
  XNOR2_X1 U10377 ( .A(n12484), .B(n12489), .ZN(n12169) );
  XNOR2_X1 U10378 ( .A(n8692), .B(n8246), .ZN(n11860) );
  NAND2_X1 U10379 ( .A1(n11860), .A2(n7428), .ZN(n8695) );
  NAND2_X1 U10380 ( .A1(n8706), .A2(n12914), .ZN(n8708) );
  NAND2_X1 U10381 ( .A1(n8708), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8693) );
  XNOR2_X1 U10382 ( .A(n8693), .B(P1_IR_REG_10__SCAN_IN), .ZN(n11319) );
  AOI22_X1 U10383 ( .A1(n8758), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n11319), 
        .B2(n8864), .ZN(n8694) );
  NAND2_X1 U10384 ( .A1(n8922), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8703) );
  NAND2_X1 U10385 ( .A1(n8896), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n8702) );
  NAND2_X1 U10386 ( .A1(n8721), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n8697) );
  INV_X1 U10387 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n8696) );
  NAND2_X1 U10388 ( .A1(n8697), .A2(n8696), .ZN(n8699) );
  AND2_X1 U10389 ( .A1(n8699), .A2(n8698), .ZN(n12281) );
  NAND2_X1 U10390 ( .A1(n8925), .A2(n12281), .ZN(n8701) );
  NAND2_X1 U10391 ( .A1(n8921), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n8700) );
  NAND4_X1 U10392 ( .A1(n8703), .A2(n8702), .A3(n8701), .A4(n8700), .ZN(n15186) );
  XNOR2_X1 U10393 ( .A(n12272), .B(n12271), .ZN(n12167) );
  XNOR2_X1 U10394 ( .A(n8705), .B(n8704), .ZN(n11854) );
  NAND2_X1 U10395 ( .A1(n11854), .A2(n7428), .ZN(n8710) );
  OR2_X1 U10396 ( .A1(n8706), .A2(n12914), .ZN(n8707) );
  AOI22_X1 U10397 ( .A1(n8758), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n8864), .B2(
        n11175), .ZN(n8709) );
  NAND2_X1 U10398 ( .A1(n8921), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n8714) );
  NAND2_X1 U10399 ( .A1(n8922), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n8713) );
  XNOR2_X1 U10400 ( .A(n8721), .B(n11986), .ZN(n11935) );
  NAND2_X1 U10401 ( .A1(n8925), .A2(n11935), .ZN(n8712) );
  NAND2_X1 U10402 ( .A1(n8926), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n8711) );
  NAND4_X1 U10403 ( .A1(n8714), .A2(n8713), .A3(n8712), .A4(n8711), .ZN(n15187) );
  INV_X1 U10404 ( .A(n15187), .ZN(n12006) );
  XNOR2_X1 U10405 ( .A(n12010), .B(n12006), .ZN(n11920) );
  XNOR2_X1 U10406 ( .A(n8716), .B(n8715), .ZN(n11671) );
  NAND2_X1 U10407 ( .A1(n11671), .A2(n7428), .ZN(n8719) );
  XNOR2_X1 U10408 ( .A(n8717), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10758) );
  AOI22_X1 U10409 ( .A1(n8758), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n8864), .B2(
        n10758), .ZN(n8718) );
  NAND2_X1 U10410 ( .A1(n8719), .A2(n8718), .ZN(n16162) );
  NAND2_X1 U10411 ( .A1(n8922), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n8725) );
  NAND2_X1 U10412 ( .A1(n8921), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n8724) );
  NOR2_X1 U10413 ( .A1(n8734), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8720) );
  OR2_X1 U10414 ( .A1(n8721), .A2(n8720), .ZN(n11827) );
  INV_X1 U10415 ( .A(n11827), .ZN(n16172) );
  NAND2_X1 U10416 ( .A1(n8925), .A2(n16172), .ZN(n8723) );
  NAND2_X1 U10417 ( .A1(n8926), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n8722) );
  NAND4_X1 U10418 ( .A1(n8725), .A2(n8724), .A3(n8723), .A4(n8722), .ZN(n15188) );
  XNOR2_X1 U10419 ( .A(n16162), .B(n11931), .ZN(n16157) );
  XNOR2_X1 U10420 ( .A(n8727), .B(n8726), .ZN(n11543) );
  NAND2_X1 U10421 ( .A1(n11543), .A2(n7428), .ZN(n8731) );
  NAND2_X1 U10422 ( .A1(n8728), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8729) );
  XNOR2_X1 U10423 ( .A(n8729), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10756) );
  AOI22_X1 U10424 ( .A1(n8758), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n8864), .B2(
        n10756), .ZN(n8730) );
  NAND2_X1 U10425 ( .A1(n8731), .A2(n8730), .ZN(n16132) );
  NAND2_X1 U10426 ( .A1(n8922), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n8738) );
  NAND2_X1 U10427 ( .A1(n8896), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n8737) );
  AND2_X1 U10428 ( .A1(n8833), .A2(n8732), .ZN(n8733) );
  NOR2_X1 U10429 ( .A1(n8734), .A2(n8733), .ZN(n11665) );
  NAND2_X1 U10430 ( .A1(n8925), .A2(n11665), .ZN(n8736) );
  NAND2_X1 U10431 ( .A1(n8921), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n8735) );
  NAND4_X1 U10432 ( .A1(n8738), .A2(n8737), .A3(n8736), .A4(n8735), .ZN(n15189) );
  XNOR2_X1 U10433 ( .A(n16132), .B(n15189), .ZN(n11924) );
  NAND2_X1 U10434 ( .A1(n8762), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n8741) );
  NAND2_X1 U10435 ( .A1(n8763), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n8740) );
  NAND2_X1 U10436 ( .A1(n8761), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n8739) );
  NOR2_X1 U10437 ( .A1(n8774), .A2(n7671), .ZN(n8743) );
  MUX2_X1 U10438 ( .A(n7671), .B(n8743), .S(P1_IR_REG_2__SCAN_IN), .Z(n8744)
         );
  INV_X1 U10439 ( .A(n8744), .ZN(n8745) );
  INV_X1 U10440 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n13132) );
  NAND2_X1 U10441 ( .A1(n8774), .A2(n13132), .ZN(n8807) );
  NAND2_X1 U10442 ( .A1(n8745), .A2(n8807), .ZN(n10972) );
  XNOR2_X1 U10443 ( .A(n8747), .B(n8746), .ZN(n10421) );
  OR2_X1 U10444 ( .A1(n7426), .A2(n7749), .ZN(n8748) );
  NAND2_X1 U10445 ( .A1(n8761), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n8754) );
  INV_X1 U10446 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n10958) );
  NAND2_X1 U10447 ( .A1(n8925), .A2(n10958), .ZN(n8753) );
  NAND2_X1 U10448 ( .A1(n8926), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n8752) );
  NAND2_X1 U10449 ( .A1(n8921), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n8751) );
  NAND4_X2 U10450 ( .A1(n8754), .A2(n8753), .A3(n8752), .A4(n8751), .ZN(n15193) );
  XNOR2_X1 U10451 ( .A(n8756), .B(n8755), .ZN(n10429) );
  NAND2_X1 U10452 ( .A1(n8807), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8757) );
  XNOR2_X1 U10453 ( .A(n8757), .B(P1_IR_REG_3__SCAN_IN), .ZN(n10623) );
  NAND2_X1 U10454 ( .A1(n8864), .A2(n10623), .ZN(n8760) );
  NAND2_X1 U10455 ( .A1(n8758), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8759) );
  OAI211_X1 U10456 ( .C1(n8772), .C2(n10429), .A(n8760), .B(n8759), .ZN(n11114) );
  XNOR2_X1 U10457 ( .A(n15193), .B(n11114), .ZN(n11109) );
  NAND2_X1 U10458 ( .A1(n8925), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n8766) );
  NAND2_X1 U10459 ( .A1(n8761), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8765) );
  AOI21_X1 U10460 ( .B1(P1_REG2_REG_1__SCAN_IN), .B2(n8763), .A(n8364), .ZN(
        n8764) );
  NAND2_X1 U10461 ( .A1(n10420), .A2(n8768), .ZN(n8782) );
  NAND2_X1 U10462 ( .A1(n8767), .A2(n8769), .ZN(n10305) );
  NAND2_X1 U10463 ( .A1(n8782), .A2(n10305), .ZN(n8770) );
  XNOR2_X1 U10464 ( .A(n8770), .B(n12989), .ZN(n8771) );
  OR2_X1 U10465 ( .A1(n7426), .A2(n10464), .ZN(n8777) );
  INV_X1 U10466 ( .A(n8774), .ZN(n8775) );
  INV_X1 U10467 ( .A(SI_0_), .ZN(n8780) );
  INV_X1 U10468 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8779) );
  OAI21_X1 U10469 ( .B1(n10432), .B2(n8780), .A(n8779), .ZN(n8781) );
  AND2_X1 U10470 ( .A1(n8782), .A2(n8781), .ZN(n15608) );
  AOI22_X1 U10471 ( .A1(n8790), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_IR_REG_30__SCAN_IN), .B2(P1_REG0_REG_0__SCAN_IN), .ZN(n8788) );
  INV_X1 U10472 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n8785) );
  NAND2_X1 U10473 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(P1_IR_REG_30__SCAN_IN), 
        .ZN(n8784) );
  OAI21_X1 U10474 ( .B1(n8785), .B2(P1_IR_REG_30__SCAN_IN), .A(n8784), .ZN(
        n8786) );
  NAND2_X1 U10475 ( .A1(n8783), .A2(n8786), .ZN(n8787) );
  OAI21_X1 U10476 ( .B1(n8783), .B2(n8788), .A(n8787), .ZN(n8789) );
  NAND2_X1 U10477 ( .A1(n8789), .A2(n8380), .ZN(n8798) );
  AOI22_X1 U10478 ( .A1(n8790), .A2(P1_REG3_REG_0__SCAN_IN), .B1(
        P1_REG1_REG_0__SCAN_IN), .B2(P1_IR_REG_30__SCAN_IN), .ZN(n8794) );
  INV_X1 U10479 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n15751) );
  NAND2_X1 U10480 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(P1_REG3_REG_0__SCAN_IN), 
        .ZN(n8791) );
  OAI21_X1 U10481 ( .B1(n15751), .B2(P1_IR_REG_30__SCAN_IN), .A(n8791), .ZN(
        n8792) );
  NAND2_X1 U10482 ( .A1(n8783), .A2(n8792), .ZN(n8793) );
  OAI21_X1 U10483 ( .B1(n8783), .B2(n8794), .A(n8793), .ZN(n8796) );
  NAND2_X1 U10484 ( .A1(n8796), .A2(n8795), .ZN(n8797) );
  INV_X1 U10485 ( .A(n15197), .ZN(n10534) );
  NAND2_X1 U10486 ( .A1(n11080), .A2(n10534), .ZN(n10880) );
  NAND2_X1 U10487 ( .A1(n16032), .A2(n15197), .ZN(n8799) );
  NAND2_X1 U10488 ( .A1(n8922), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n8804) );
  NAND2_X1 U10489 ( .A1(n8926), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n8803) );
  INV_X1 U10490 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n8800) );
  XNOR2_X1 U10491 ( .A(n8800), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n11342) );
  NAND2_X1 U10492 ( .A1(n8925), .A2(n11342), .ZN(n8802) );
  NAND2_X1 U10493 ( .A1(n8921), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n8801) );
  XNOR2_X1 U10494 ( .A(n8806), .B(n8805), .ZN(n11043) );
  NAND2_X1 U10495 ( .A1(n11043), .A2(n8814), .ZN(n8810) );
  OR2_X1 U10496 ( .A1(n8807), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n8815) );
  NAND2_X1 U10497 ( .A1(n8815), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8808) );
  XNOR2_X1 U10498 ( .A(n8808), .B(P1_IR_REG_4__SCAN_IN), .ZN(n10817) );
  AOI22_X1 U10499 ( .A1(n8758), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n8864), .B2(
        n10817), .ZN(n8809) );
  NAND2_X1 U10500 ( .A1(n8810), .A2(n8809), .ZN(n11341) );
  NOR2_X1 U10501 ( .A1(n8811), .A2(n11488), .ZN(n8840) );
  XNOR2_X1 U10502 ( .A(n8812), .B(n8813), .ZN(n11130) );
  NAND2_X1 U10503 ( .A1(n11130), .A2(n7428), .ZN(n8818) );
  OAI21_X1 U10504 ( .B1(n8815), .B2(P1_IR_REG_4__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8816) );
  XNOR2_X1 U10505 ( .A(n8816), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10680) );
  AOI22_X1 U10506 ( .A1(n8758), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n8864), .B2(
        n10680), .ZN(n8817) );
  NAND2_X1 U10507 ( .A1(n8818), .A2(n8817), .ZN(n11587) );
  NAND2_X1 U10508 ( .A1(n8921), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n8823) );
  NAND2_X1 U10509 ( .A1(n8922), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n8822) );
  AOI21_X1 U10510 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n8819) );
  NOR2_X1 U10511 ( .A1(n8819), .A2(n8834), .ZN(n11586) );
  NAND2_X1 U10512 ( .A1(n8925), .A2(n11586), .ZN(n8821) );
  NAND2_X1 U10513 ( .A1(n8896), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n8820) );
  NAND4_X1 U10514 ( .A1(n8823), .A2(n8822), .A3(n8821), .A4(n8820), .ZN(n15191) );
  XNOR2_X1 U10515 ( .A(n11587), .B(n15191), .ZN(n11510) );
  NAND2_X1 U10516 ( .A1(n8812), .A2(n8824), .ZN(n8826) );
  NAND2_X1 U10517 ( .A1(n8826), .A2(n8825), .ZN(n8828) );
  XNOR2_X1 U10518 ( .A(n8828), .B(n8827), .ZN(n11539) );
  NAND2_X1 U10519 ( .A1(n11539), .A2(n7428), .ZN(n8832) );
  NAND2_X1 U10520 ( .A1(n8829), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8830) );
  XNOR2_X1 U10521 ( .A(n8830), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10687) );
  AOI22_X1 U10522 ( .A1(n8758), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n8864), .B2(
        n10687), .ZN(n8831) );
  NAND2_X1 U10523 ( .A1(n8832), .A2(n8831), .ZN(n11648) );
  NAND2_X1 U10524 ( .A1(n8921), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n8839) );
  NAND2_X1 U10525 ( .A1(n8922), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n8838) );
  OAI21_X1 U10526 ( .B1(n8834), .B2(P1_REG3_REG_6__SCAN_IN), .A(n8833), .ZN(
        n16109) );
  INV_X1 U10527 ( .A(n16109), .ZN(n8835) );
  NAND2_X1 U10528 ( .A1(n8925), .A2(n8835), .ZN(n8837) );
  NAND2_X1 U10529 ( .A1(n8896), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n8836) );
  NAND4_X1 U10530 ( .A1(n8839), .A2(n8838), .A3(n8837), .A4(n8836), .ZN(n15190) );
  XNOR2_X1 U10531 ( .A(n11648), .B(n15190), .ZN(n11642) );
  NAND4_X1 U10532 ( .A1(n11924), .A2(n8840), .A3(n11510), .A4(n11642), .ZN(
        n8841) );
  OR4_X1 U10533 ( .A1(n12167), .A2(n11920), .A3(n16157), .A4(n8841), .ZN(n8842) );
  OR4_X1 U10534 ( .A1(n12648), .A2(n12486), .A3(n12169), .A4(n8842), .ZN(n8843) );
  OR4_X1 U10535 ( .A1(n15461), .A2(n12702), .A3(n12650), .A4(n8843), .ZN(n8844) );
  NOR2_X1 U10536 ( .A1(n15443), .A2(n8844), .ZN(n8873) );
  XNOR2_X1 U10537 ( .A(n8846), .B(n8845), .ZN(n13404) );
  NAND2_X1 U10538 ( .A1(n13404), .A2(n7428), .ZN(n8849) );
  AOI22_X1 U10539 ( .A1(n8758), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n8864), 
        .B2(n7429), .ZN(n8848) );
  NOR2_X1 U10540 ( .A1(n8869), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8850) );
  OR2_X1 U10541 ( .A1(n8851), .A2(n8850), .ZN(n15410) );
  INV_X1 U10542 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n8854) );
  NAND2_X1 U10543 ( .A1(n8921), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8853) );
  NAND2_X1 U10544 ( .A1(n8926), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n8852) );
  OAI211_X1 U10545 ( .C1(n8855), .C2(n8854), .A(n8853), .B(n8852), .ZN(n8856)
         );
  INV_X1 U10546 ( .A(n8856), .ZN(n8857) );
  XNOR2_X1 U10547 ( .A(n15534), .B(n15421), .ZN(n15402) );
  XNOR2_X1 U10548 ( .A(n8859), .B(n8858), .ZN(n13398) );
  NAND2_X1 U10549 ( .A1(n13398), .A2(n7428), .ZN(n8866) );
  NAND2_X1 U10550 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n8860) );
  NAND2_X1 U10551 ( .A1(n8861), .A2(n8860), .ZN(n8863) );
  XNOR2_X1 U10552 ( .A(n8863), .B(n8862), .ZN(n15233) );
  AOI22_X1 U10553 ( .A1(n8758), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n15233), 
        .B2(n8864), .ZN(n8865) );
  NOR2_X1 U10554 ( .A1(n8867), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8868) );
  OR2_X1 U10555 ( .A1(n8869), .A2(n8868), .ZN(n15429) );
  AOI22_X1 U10556 ( .A1(n8922), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n8896), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n8871) );
  NAND2_X1 U10557 ( .A1(n8921), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n8870) );
  OAI211_X1 U10558 ( .C1(n15429), .C2(n8872), .A(n8871), .B(n8870), .ZN(n15182) );
  XNOR2_X1 U10559 ( .A(n15542), .B(n15182), .ZN(n15423) );
  NAND4_X1 U10560 ( .A1(n13336), .A2(n8873), .A3(n15402), .A4(n15423), .ZN(
        n8874) );
  NOR2_X1 U10561 ( .A1(n15369), .A2(n8874), .ZN(n8875) );
  AND3_X1 U10562 ( .A1(n15321), .A2(n13337), .A3(n8875), .ZN(n8903) );
  XNOR2_X1 U10563 ( .A(n8877), .B(n8876), .ZN(n13462) );
  NAND2_X1 U10564 ( .A1(n13462), .A2(n7428), .ZN(n8879) );
  NAND2_X1 U10565 ( .A1(n8758), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8878) );
  NAND2_X1 U10566 ( .A1(n8921), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n8886) );
  NAND2_X1 U10567 ( .A1(n8922), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8885) );
  INV_X1 U10568 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8882) );
  AOI21_X1 U10569 ( .B1(n8882), .B2(n8881), .A(n8880), .ZN(n15333) );
  NAND2_X1 U10570 ( .A1(n8925), .A2(n15333), .ZN(n8884) );
  NAND2_X1 U10571 ( .A1(n8896), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8883) );
  NAND4_X1 U10572 ( .A1(n8886), .A2(n8885), .A3(n8884), .A4(n8883), .ZN(n15311) );
  XNOR2_X1 U10573 ( .A(n15334), .B(n15311), .ZN(n13338) );
  NOR2_X1 U10574 ( .A1(n8887), .A2(SI_22_), .ZN(n8888) );
  AOI21_X1 U10575 ( .B1(n8890), .B2(n8889), .A(n8888), .ZN(n8893) );
  XNOR2_X1 U10576 ( .A(n8891), .B(SI_23_), .ZN(n8892) );
  XNOR2_X1 U10577 ( .A(n8893), .B(n8892), .ZN(n13387) );
  NAND2_X1 U10578 ( .A1(n13387), .A2(n7428), .ZN(n8895) );
  NAND2_X1 U10579 ( .A1(n8758), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8894) );
  NAND2_X1 U10580 ( .A1(n8922), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n8902) );
  NAND2_X1 U10581 ( .A1(n8896), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n8901) );
  INV_X1 U10582 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n15100) );
  AOI21_X1 U10583 ( .B1(n15100), .B2(n8898), .A(n8897), .ZN(n15345) );
  NAND2_X1 U10584 ( .A1(n8925), .A2(n15345), .ZN(n8900) );
  NAND2_X1 U10585 ( .A1(n8921), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8899) );
  NAND4_X1 U10586 ( .A1(n8902), .A2(n8901), .A3(n8900), .A4(n8899), .ZN(n15180) );
  XNOR2_X1 U10587 ( .A(n15349), .B(n15180), .ZN(n15342) );
  NAND4_X1 U10588 ( .A1(n15293), .A2(n8903), .A3(n13338), .A4(n15342), .ZN(
        n8904) );
  NOR2_X1 U10589 ( .A1(n15280), .A2(n8904), .ZN(n8931) );
  INV_X1 U10590 ( .A(n8905), .ZN(n8907) );
  NAND2_X1 U10591 ( .A1(n8907), .A2(n8906), .ZN(n8909) );
  NAND2_X1 U10592 ( .A1(n8909), .A2(n8908), .ZN(n13513) );
  NAND2_X1 U10593 ( .A1(n13513), .A2(n7428), .ZN(n8911) );
  NAND2_X1 U10594 ( .A1(n8758), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8910) );
  NAND2_X1 U10595 ( .A1(n8923), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n13348) );
  INV_X1 U10596 ( .A(n13348), .ZN(n8912) );
  NAND2_X1 U10597 ( .A1(n8925), .A2(n8912), .ZN(n8916) );
  NAND2_X1 U10598 ( .A1(n8922), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8915) );
  NAND2_X1 U10599 ( .A1(n8926), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8914) );
  NAND2_X1 U10600 ( .A1(n8921), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8913) );
  AND4_X1 U10601 ( .A1(n8916), .A2(n8915), .A3(n8914), .A4(n8913), .ZN(n13599)
         );
  NAND2_X1 U10602 ( .A1(n13372), .A2(n7428), .ZN(n8920) );
  NAND2_X1 U10603 ( .A1(n8758), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8919) );
  NAND2_X1 U10604 ( .A1(n8921), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8930) );
  NAND2_X1 U10605 ( .A1(n8922), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n8929) );
  OAI21_X1 U10606 ( .B1(n8923), .B2(P1_REG3_REG_28__SCAN_IN), .A(n13348), .ZN(
        n15272) );
  INV_X1 U10607 ( .A(n15272), .ZN(n8924) );
  NAND2_X1 U10608 ( .A1(n8925), .A2(n8924), .ZN(n8928) );
  NAND2_X1 U10609 ( .A1(n8926), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n8927) );
  NAND4_X1 U10610 ( .A1(n8930), .A2(n8929), .A3(n8928), .A4(n8927), .ZN(n15282) );
  XNOR2_X1 U10611 ( .A(n15274), .B(n15282), .ZN(n15265) );
  NAND4_X1 U10612 ( .A1(n8932), .A2(n8931), .A3(n13368), .A4(n15265), .ZN(
        n8933) );
  XNOR2_X1 U10613 ( .A(n8934), .B(n15244), .ZN(n8945) );
  INV_X1 U10614 ( .A(n8939), .ZN(n8944) );
  INV_X1 U10615 ( .A(n9095), .ZN(n8935) );
  XNOR2_X1 U10616 ( .A(n8936), .B(n8935), .ZN(n8941) );
  XNOR2_X1 U10617 ( .A(n8937), .B(n9095), .ZN(n8938) );
  NAND2_X1 U10618 ( .A1(n15253), .A2(n8938), .ZN(n8940) );
  OAI211_X1 U10619 ( .C1(n15253), .C2(n8941), .A(n8940), .B(n8939), .ZN(n8942)
         );
  INV_X1 U10620 ( .A(n8942), .ZN(n8943) );
  AOI21_X2 U10621 ( .B1(n8945), .B2(n8944), .A(n8943), .ZN(n9129) );
  OAI21_X1 U10622 ( .B1(n15177), .B2(n8954), .A(n15178), .ZN(n8946) );
  MUX2_X1 U10623 ( .A(n8946), .B(n15472), .S(n7427), .Z(n9122) );
  NAND3_X1 U10624 ( .A1(n9129), .A2(n13236), .A3(n9122), .ZN(n8947) );
  OAI21_X1 U10625 ( .B1(n9118), .B2(n9119), .A(n8947), .ZN(n9092) );
  MUX2_X1 U10626 ( .A(n15282), .B(n15274), .S(n7427), .Z(n9089) );
  MUX2_X1 U10627 ( .A(n15171), .B(n15485), .S(n7427), .Z(n9080) );
  NAND2_X1 U10628 ( .A1(n15194), .A2(n8958), .ZN(n8950) );
  INV_X1 U10629 ( .A(n15194), .ZN(n11106) );
  NAND2_X1 U10630 ( .A1(n11106), .A2(n8952), .ZN(n8949) );
  MUX2_X1 U10631 ( .A(n8950), .B(n8949), .S(n7430), .Z(n8951) );
  OAI21_X1 U10632 ( .B1(n7421), .B2(n15197), .A(n10878), .ZN(n8953) );
  NAND2_X1 U10633 ( .A1(n8953), .A2(n11080), .ZN(n8962) );
  OR2_X1 U10634 ( .A1(n8954), .A2(n12593), .ZN(n8956) );
  INV_X1 U10635 ( .A(n8954), .ZN(n8955) );
  OAI22_X1 U10636 ( .A1(n15197), .A2(n8956), .B1(n8955), .B2(n10881), .ZN(
        n8957) );
  NAND2_X1 U10637 ( .A1(n8957), .A2(n16032), .ZN(n8961) );
  INV_X1 U10638 ( .A(n10878), .ZN(n10532) );
  NAND2_X1 U10639 ( .A1(n15197), .A2(n8952), .ZN(n8959) );
  OAI21_X1 U10640 ( .B1(n15197), .B2(n10532), .A(n8959), .ZN(n8960) );
  OR2_X1 U10641 ( .A1(n15195), .A2(n11236), .ZN(n11006) );
  MUX2_X1 U10642 ( .A(n11074), .B(n10876), .S(n8952), .Z(n8963) );
  NAND3_X1 U10643 ( .A1(n8964), .A2(n15195), .A3(n11236), .ZN(n8965) );
  NAND3_X1 U10644 ( .A1(n8966), .A2(n8965), .A3(n11104), .ZN(n8968) );
  INV_X1 U10645 ( .A(n11109), .ZN(n8967) );
  NAND3_X1 U10646 ( .A1(n8951), .A2(n8968), .A3(n11109), .ZN(n8971) );
  NAND2_X1 U10647 ( .A1(n15193), .A2(n8952), .ZN(n8969) );
  INV_X2 U10648 ( .A(n11114), .ZN(n16077) );
  NAND2_X1 U10649 ( .A1(n8971), .A2(n8970), .ZN(n8973) );
  MUX2_X1 U10650 ( .A(n11341), .B(n15192), .S(n8952), .Z(n8974) );
  MUX2_X1 U10651 ( .A(n15192), .B(n11341), .S(n8952), .Z(n8972) );
  INV_X1 U10652 ( .A(n8974), .ZN(n8975) );
  MUX2_X1 U10653 ( .A(n15191), .B(n11587), .S(n8952), .Z(n8979) );
  MUX2_X1 U10654 ( .A(n15191), .B(n11587), .S(n8948), .Z(n8976) );
  NAND2_X1 U10655 ( .A1(n8977), .A2(n8976), .ZN(n8983) );
  INV_X1 U10656 ( .A(n8978), .ZN(n8981) );
  INV_X1 U10657 ( .A(n8979), .ZN(n8980) );
  NAND2_X1 U10658 ( .A1(n8981), .A2(n8980), .ZN(n8982) );
  NAND2_X1 U10659 ( .A1(n8983), .A2(n8982), .ZN(n8985) );
  MUX2_X1 U10660 ( .A(n15190), .B(n11648), .S(n8948), .Z(n8986) );
  MUX2_X1 U10661 ( .A(n15190), .B(n11648), .S(n9085), .Z(n8984) );
  INV_X1 U10662 ( .A(n8986), .ZN(n8987) );
  MUX2_X1 U10663 ( .A(n15189), .B(n16132), .S(n7427), .Z(n8991) );
  MUX2_X1 U10664 ( .A(n15189), .B(n16132), .S(n8948), .Z(n8988) );
  NAND2_X1 U10665 ( .A1(n8989), .A2(n8988), .ZN(n8995) );
  INV_X1 U10666 ( .A(n8990), .ZN(n8993) );
  INV_X1 U10667 ( .A(n8991), .ZN(n8992) );
  NAND2_X1 U10668 ( .A1(n8993), .A2(n8992), .ZN(n8994) );
  NAND2_X1 U10669 ( .A1(n8995), .A2(n8994), .ZN(n8997) );
  MUX2_X1 U10670 ( .A(n15188), .B(n16162), .S(n8948), .Z(n8998) );
  MUX2_X1 U10671 ( .A(n15188), .B(n16162), .S(n7427), .Z(n8996) );
  INV_X1 U10672 ( .A(n8998), .ZN(n8999) );
  MUX2_X1 U10673 ( .A(n15187), .B(n12010), .S(n7427), .Z(n9003) );
  MUX2_X1 U10674 ( .A(n15187), .B(n12010), .S(n8948), .Z(n9000) );
  NAND2_X1 U10675 ( .A1(n9001), .A2(n9000), .ZN(n9004) );
  MUX2_X1 U10676 ( .A(n15186), .B(n12272), .S(n8948), .Z(n9006) );
  MUX2_X1 U10677 ( .A(n15186), .B(n12272), .S(n7427), .Z(n9005) );
  INV_X1 U10678 ( .A(n9006), .ZN(n9007) );
  MUX2_X1 U10679 ( .A(n15185), .B(n12484), .S(n7427), .Z(n9011) );
  MUX2_X1 U10680 ( .A(n15185), .B(n12484), .S(n8948), .Z(n9008) );
  NAND2_X1 U10681 ( .A1(n9009), .A2(n9008), .ZN(n9015) );
  INV_X1 U10682 ( .A(n9010), .ZN(n9013) );
  INV_X1 U10683 ( .A(n9011), .ZN(n9012) );
  NAND2_X1 U10684 ( .A1(n9013), .A2(n9012), .ZN(n9014) );
  NAND2_X1 U10685 ( .A1(n9015), .A2(n9014), .ZN(n9017) );
  MUX2_X1 U10686 ( .A(n15184), .B(n16266), .S(n8948), .Z(n9018) );
  MUX2_X1 U10687 ( .A(n15184), .B(n16266), .S(n7427), .Z(n9016) );
  INV_X1 U10688 ( .A(n9018), .ZN(n9019) );
  MUX2_X1 U10689 ( .A(n15183), .B(n16277), .S(n7427), .Z(n9022) );
  MUX2_X1 U10690 ( .A(n15183), .B(n16277), .S(n8948), .Z(n9020) );
  MUX2_X1 U10691 ( .A(n16321), .B(n15089), .S(n8948), .Z(n9025) );
  MUX2_X1 U10692 ( .A(n16321), .B(n15089), .S(n7427), .Z(n9023) );
  INV_X1 U10693 ( .A(n9025), .ZN(n9026) );
  MUX2_X1 U10694 ( .A(n16348), .B(n13354), .S(n7427), .Z(n9029) );
  MUX2_X1 U10695 ( .A(n16348), .B(n13354), .S(n8948), .Z(n9027) );
  NAND2_X1 U10696 ( .A1(n9028), .A2(n9027), .ZN(n9030) );
  MUX2_X1 U10697 ( .A(n16322), .B(n15454), .S(n8948), .Z(n9032) );
  MUX2_X1 U10698 ( .A(n16322), .B(n15454), .S(n7427), .Z(n9031) );
  MUX2_X1 U10699 ( .A(n16350), .B(n15550), .S(n7427), .Z(n9036) );
  MUX2_X1 U10700 ( .A(n16350), .B(n15550), .S(n8948), .Z(n9033) );
  NAND2_X1 U10701 ( .A1(n9034), .A2(n9033), .ZN(n9040) );
  INV_X1 U10702 ( .A(n9035), .ZN(n9038) );
  INV_X1 U10703 ( .A(n9036), .ZN(n9037) );
  NAND2_X1 U10704 ( .A1(n9038), .A2(n9037), .ZN(n9039) );
  NAND2_X1 U10705 ( .A1(n9040), .A2(n9039), .ZN(n9042) );
  MUX2_X1 U10706 ( .A(n15542), .B(n15182), .S(n7427), .Z(n9043) );
  MUX2_X1 U10707 ( .A(n15182), .B(n15542), .S(n7427), .Z(n9041) );
  INV_X1 U10708 ( .A(n9043), .ZN(n9044) );
  MUX2_X1 U10709 ( .A(n15421), .B(n15534), .S(n7427), .Z(n9046) );
  MUX2_X1 U10710 ( .A(n15421), .B(n15534), .S(n8948), .Z(n9045) );
  INV_X1 U10711 ( .A(n9046), .ZN(n9047) );
  MUX2_X1 U10712 ( .A(n15375), .B(n15528), .S(n8948), .Z(n9051) );
  NAND2_X1 U10713 ( .A1(n9050), .A2(n9051), .ZN(n9049) );
  MUX2_X1 U10714 ( .A(n15375), .B(n15528), .S(n7427), .Z(n9048) );
  INV_X1 U10715 ( .A(n9051), .ZN(n9052) );
  NAND2_X1 U10716 ( .A1(n9053), .A2(n9052), .ZN(n9054) );
  MUX2_X1 U10717 ( .A(n15181), .B(n15525), .S(n7427), .Z(n9056) );
  MUX2_X1 U10718 ( .A(n15181), .B(n15525), .S(n8948), .Z(n9055) );
  INV_X1 U10719 ( .A(n9056), .ZN(n9057) );
  NOR2_X1 U10720 ( .A1(n15374), .A2(n8948), .ZN(n9059) );
  OAI21_X1 U10721 ( .B1(n15097), .B2(n7427), .A(n7417), .ZN(n9058) );
  OAI21_X1 U10722 ( .B1(n9059), .B2(n7417), .A(n9058), .ZN(n9060) );
  MUX2_X1 U10723 ( .A(n15180), .B(n15349), .S(n7427), .Z(n9063) );
  MUX2_X1 U10724 ( .A(n15180), .B(n15349), .S(n8948), .Z(n9062) );
  INV_X1 U10725 ( .A(n9063), .ZN(n9064) );
  MUX2_X1 U10726 ( .A(n15311), .B(n15334), .S(n8948), .Z(n9067) );
  MUX2_X1 U10727 ( .A(n15311), .B(n15334), .S(n7427), .Z(n9065) );
  INV_X1 U10728 ( .A(n9067), .ZN(n9068) );
  MUX2_X1 U10729 ( .A(n15329), .B(n15498), .S(n7427), .Z(n9072) );
  MUX2_X1 U10730 ( .A(n15329), .B(n15498), .S(n8948), .Z(n9069) );
  NAND2_X1 U10731 ( .A1(n9070), .A2(n9069), .ZN(n9076) );
  INV_X1 U10732 ( .A(n9071), .ZN(n9074) );
  INV_X1 U10733 ( .A(n9072), .ZN(n9073) );
  NAND2_X1 U10734 ( .A1(n9074), .A2(n9073), .ZN(n9075) );
  MUX2_X1 U10735 ( .A(n15312), .B(n15491), .S(n8948), .Z(n9078) );
  MUX2_X1 U10736 ( .A(n15312), .B(n15491), .S(n7427), .Z(n9077) );
  MUX2_X1 U10737 ( .A(n15288), .B(n15295), .S(n7427), .Z(n9079) );
  OAI21_X1 U10738 ( .B1(n7899), .B2(n9082), .A(n9081), .ZN(n9084) );
  MUX2_X1 U10739 ( .A(n15274), .B(n15282), .S(n7427), .Z(n9083) );
  NAND2_X1 U10740 ( .A1(n9084), .A2(n9083), .ZN(n9088) );
  INV_X1 U10741 ( .A(n9083), .ZN(n9087) );
  INV_X1 U10742 ( .A(n9084), .ZN(n9086) );
  MUX2_X1 U10743 ( .A(n15179), .B(n13344), .S(n7427), .Z(n9090) );
  MUX2_X1 U10744 ( .A(n15474), .B(n13599), .S(n7427), .Z(n9091) );
  NOR2_X1 U10745 ( .A1(n9091), .A2(n9090), .ZN(n9094) );
  INV_X1 U10746 ( .A(n9093), .ZN(n9097) );
  INV_X1 U10747 ( .A(n13236), .ZN(n10453) );
  AOI211_X1 U10748 ( .C1(n9121), .C2(n9122), .A(n10453), .B(n9094), .ZN(n9096)
         );
  NOR2_X1 U10749 ( .A1(n9131), .A2(n9095), .ZN(n9120) );
  NAND3_X1 U10750 ( .A1(n9097), .A2(n9096), .A3(n9120), .ZN(n9134) );
  INV_X1 U10751 ( .A(P1_B_REG_SCAN_IN), .ZN(n13346) );
  AOI21_X1 U10752 ( .B1(n13236), .B2(n9098), .A(n13346), .ZN(n9127) );
  INV_X1 U10753 ( .A(n9105), .ZN(n9106) );
  NAND3_X1 U10754 ( .A1(n9108), .A2(n9107), .A3(n9106), .ZN(n9109) );
  NAND2_X1 U10755 ( .A1(n9109), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9111) );
  INV_X1 U10756 ( .A(n10454), .ZN(n9115) );
  INV_X1 U10757 ( .A(n10529), .ZN(n9116) );
  NAND2_X1 U10758 ( .A1(n12527), .A2(n15244), .ZN(n10533) );
  NOR2_X1 U10759 ( .A1(n15583), .A2(n10953), .ZN(n11071) );
  INV_X1 U10760 ( .A(n15594), .ZN(n15750) );
  NAND3_X1 U10761 ( .A1(n11071), .A2(n15750), .A3(n15455), .ZN(n9126) );
  INV_X1 U10762 ( .A(n9122), .ZN(n9117) );
  NOR3_X1 U10763 ( .A1(n9119), .A2(n9118), .A3(n9117), .ZN(n9125) );
  INV_X1 U10764 ( .A(n9120), .ZN(n9123) );
  NOR4_X1 U10765 ( .A1(n9123), .A2(n9122), .A3(n9121), .A4(n10453), .ZN(n9124)
         );
  AOI211_X1 U10766 ( .C1(n9127), .C2(n9126), .A(n9125), .B(n9124), .ZN(n9133)
         );
  INV_X1 U10767 ( .A(n9128), .ZN(n9130) );
  OAI211_X1 U10768 ( .C1(n9131), .C2(n9130), .A(n9129), .B(n13236), .ZN(n9132)
         );
  NAND4_X1 U10769 ( .A1(n9135), .A2(n9134), .A3(n9133), .A4(n9132), .ZN(
        P1_U3242) );
  NAND2_X1 U10770 ( .A1(n10303), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n9283) );
  INV_X1 U10771 ( .A(n9283), .ZN(n9136) );
  NAND2_X1 U10772 ( .A1(n9137), .A2(n9136), .ZN(n9285) );
  INV_X1 U10773 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10452) );
  NAND2_X1 U10774 ( .A1(n10452), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9138) );
  INV_X1 U10775 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10407) );
  NAND2_X1 U10776 ( .A1(n10408), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n9139) );
  NAND2_X1 U10777 ( .A1(n10428), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n9141) );
  NAND2_X1 U10778 ( .A1(n11044), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n9140) );
  NAND2_X1 U10779 ( .A1(n9141), .A2(n9140), .ZN(n9332) );
  INV_X1 U10780 ( .A(n9353), .ZN(n9144) );
  NAND2_X1 U10781 ( .A1(n10423), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n9145) );
  NAND2_X1 U10782 ( .A1(n10418), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n9142) );
  NAND2_X1 U10783 ( .A1(n9145), .A2(n9142), .ZN(n9352) );
  INV_X1 U10784 ( .A(n9352), .ZN(n9143) );
  INV_X1 U10785 ( .A(n9371), .ZN(n9146) );
  NAND2_X1 U10786 ( .A1(n10451), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n9149) );
  NAND2_X1 U10787 ( .A1(n10449), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n9147) );
  INV_X1 U10788 ( .A(n9387), .ZN(n9148) );
  NAND2_X1 U10789 ( .A1(n10463), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n9151) );
  NAND2_X1 U10790 ( .A1(n10461), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n9150) );
  NAND2_X1 U10791 ( .A1(n9399), .A2(n9398), .ZN(n9152) );
  NAND2_X1 U10792 ( .A1(n9152), .A2(n9151), .ZN(n9414) );
  NAND2_X1 U10793 ( .A1(n10483), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n9155) );
  INV_X1 U10794 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10488) );
  NAND2_X1 U10795 ( .A1(n10488), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n9153) );
  NAND2_X1 U10796 ( .A1(n9155), .A2(n9153), .ZN(n9413) );
  INV_X1 U10797 ( .A(n9413), .ZN(n9154) );
  NAND2_X1 U10798 ( .A1(n10496), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n9157) );
  INV_X1 U10799 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10494) );
  NAND2_X1 U10800 ( .A1(n10494), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n9156) );
  NAND2_X1 U10801 ( .A1(n10503), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n9159) );
  NAND2_X1 U10802 ( .A1(n10501), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n9158) );
  NAND2_X1 U10803 ( .A1(n9442), .A2(n9441), .ZN(n9444) );
  NAND2_X1 U10804 ( .A1(n9444), .A2(n9159), .ZN(n9456) );
  NAND2_X1 U10805 ( .A1(n10655), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n9161) );
  NAND2_X1 U10806 ( .A1(n10653), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n9160) );
  NAND2_X1 U10807 ( .A1(n9456), .A2(n9455), .ZN(n9458) );
  OR2_X1 U10808 ( .A1(n9162), .A2(n10727), .ZN(n9163) );
  NAND2_X1 U10809 ( .A1(n11226), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n9166) );
  INV_X1 U10810 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n11224) );
  NAND2_X1 U10811 ( .A1(n11224), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n9165) );
  NAND2_X1 U10812 ( .A1(n9490), .A2(n9166), .ZN(n9509) );
  NAND2_X1 U10813 ( .A1(n11289), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n9168) );
  NAND2_X1 U10814 ( .A1(n11294), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n9167) );
  NAND2_X1 U10815 ( .A1(n9509), .A2(n9508), .ZN(n9511) );
  NAND2_X1 U10816 ( .A1(n9511), .A2(n9168), .ZN(n9527) );
  NAND2_X1 U10817 ( .A1(n11737), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n9170) );
  NAND2_X1 U10818 ( .A1(n11735), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n9169) );
  NAND2_X1 U10819 ( .A1(n9527), .A2(n9526), .ZN(n9529) );
  NAND2_X1 U10820 ( .A1(n9529), .A2(n9170), .ZN(n9543) );
  NAND2_X1 U10821 ( .A1(n11768), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n9172) );
  NAND2_X1 U10822 ( .A1(n11775), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n9171) );
  NAND2_X1 U10823 ( .A1(n9543), .A2(n9542), .ZN(n9545) );
  NAND2_X1 U10824 ( .A1(n9545), .A2(n9172), .ZN(n9559) );
  INV_X1 U10825 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n12237) );
  NAND2_X1 U10826 ( .A1(n12237), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n9174) );
  INV_X1 U10827 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n12235) );
  NAND2_X1 U10828 ( .A1(n12235), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n9173) );
  NAND2_X1 U10829 ( .A1(n9559), .A2(n9558), .ZN(n9561) );
  NAND2_X1 U10830 ( .A1(n9578), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n9175) );
  NAND2_X1 U10831 ( .A1(n9580), .A2(n9175), .ZN(n9177) );
  NAND2_X1 U10832 ( .A1(n13252), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n9176) );
  INV_X1 U10833 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n13418) );
  NAND2_X1 U10834 ( .A1(n13418), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9179) );
  INV_X1 U10835 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n12526) );
  NAND2_X1 U10836 ( .A1(n12526), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9178) );
  NAND2_X1 U10837 ( .A1(n9179), .A2(n9178), .ZN(n9597) );
  INV_X1 U10838 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n13433) );
  NAND2_X1 U10839 ( .A1(n13433), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9181) );
  INV_X1 U10840 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n12594) );
  NAND2_X1 U10841 ( .A1(n12594), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9180) );
  INV_X1 U10842 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n13447) );
  NAND2_X1 U10843 ( .A1(n13447), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n9184) );
  INV_X1 U10844 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9182) );
  NAND2_X1 U10845 ( .A1(n9182), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n9183) );
  NAND2_X1 U10846 ( .A1(n9618), .A2(n9617), .ZN(n9620) );
  NAND2_X1 U10847 ( .A1(n13388), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9187) );
  INV_X1 U10848 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n9185) );
  NAND2_X1 U10849 ( .A1(n9185), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n9186) );
  XNOR2_X1 U10850 ( .A(n15073), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n9658) );
  INV_X1 U10851 ( .A(n9658), .ZN(n9190) );
  NAND2_X1 U10852 ( .A1(n9659), .A2(n9190), .ZN(n9193) );
  NAND2_X1 U10853 ( .A1(n9191), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9192) );
  XNOR2_X1 U10854 ( .A(n15068), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n9672) );
  XNOR2_X1 U10855 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n9684) );
  NAND2_X1 U10856 ( .A1(n15596), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9194) );
  NAND2_X1 U10857 ( .A1(n9195), .A2(n9194), .ZN(n9697) );
  XNOR2_X1 U10858 ( .A(n13373), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n9696) );
  INV_X1 U10859 ( .A(n9696), .ZN(n9197) );
  AND2_X1 U10860 ( .A1(n13246), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9196) );
  XNOR2_X1 U10861 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n9893) );
  XNOR2_X1 U10862 ( .A(n9895), .B(n9893), .ZN(n13922) );
  NOR2_X1 U10863 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_5__SCAN_IN), .ZN(
        n9200) );
  NOR2_X1 U10864 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), 
        .ZN(n9205) );
  NOR2_X1 U10865 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), 
        .ZN(n9209) );
  NAND4_X1 U10866 ( .A1(n9209), .A2(n9256), .A3(n9247), .A4(n9217), .ZN(n9210)
         );
  NAND2_X1 U10867 ( .A1(n9271), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9213) );
  AOI22_X1 U10868 ( .A1(n13922), .A2(n9916), .B1(SI_29_), .B2(n9686), .ZN(
        n14166) );
  XNOR2_X1 U10869 ( .A(n12383), .B(P3_B_REG_SCAN_IN), .ZN(n9224) );
  NAND2_X1 U10870 ( .A1(n9220), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9221) );
  NAND2_X1 U10871 ( .A1(n9219), .A2(n9222), .ZN(n9225) );
  NAND2_X1 U10872 ( .A1(n9224), .A2(n12378), .ZN(n9226) );
  NAND2_X1 U10873 ( .A1(n9226), .A2(n9227), .ZN(n9230) );
  NAND2_X1 U10874 ( .A1(n12383), .A2(n12463), .ZN(n9228) );
  NOR2_X1 U10875 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .ZN(
        n9234) );
  NOR4_X1 U10876 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n9233) );
  NOR4_X1 U10877 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n9232) );
  NOR4_X1 U10878 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n9231) );
  NAND4_X1 U10879 ( .A1(n9234), .A2(n9233), .A3(n9232), .A4(n9231), .ZN(n9240)
         );
  NOR4_X1 U10880 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n9238) );
  NOR4_X1 U10881 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n9237) );
  NOR4_X1 U10882 ( .A1(P3_D_REG_7__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_2__SCAN_IN), .ZN(n9236) );
  NOR4_X1 U10883 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_8__SCAN_IN), .ZN(n9235) );
  NAND4_X1 U10884 ( .A1(n9238), .A2(n9237), .A3(n9236), .A4(n9235), .ZN(n9239)
         );
  NOR2_X1 U10885 ( .A1(n9240), .A2(n9239), .ZN(n9241) );
  OR2_X1 U10886 ( .A1(n9230), .A2(n9241), .ZN(n9748) );
  NAND2_X1 U10887 ( .A1(n9767), .A2(n9748), .ZN(n9244) );
  OR2_X1 U10888 ( .A1(n9230), .A2(P3_D_REG_1__SCAN_IN), .ZN(n9243) );
  NAND2_X1 U10889 ( .A1(n12463), .A2(n12378), .ZN(n9242) );
  INV_X1 U10890 ( .A(n12383), .ZN(n9246) );
  NOR2_X1 U10891 ( .A1(n12463), .A2(n12378), .ZN(n9245) );
  NAND2_X1 U10892 ( .A1(n9246), .A2(n9245), .ZN(n10105) );
  NAND2_X1 U10893 ( .A1(n9253), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9249) );
  MUX2_X1 U10894 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9249), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n9251) );
  INV_X1 U10895 ( .A(n9755), .ZN(n11797) );
  NAND2_X1 U10896 ( .A1(n7506), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9252) );
  MUX2_X1 U10897 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9252), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n9254) );
  NAND2_X1 U10898 ( .A1(n9255), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9257) );
  NAND2_X1 U10899 ( .A1(n11767), .A2(n11614), .ZN(n9754) );
  XNOR2_X1 U10900 ( .A(n11797), .B(n9754), .ZN(n9261) );
  NAND2_X1 U10901 ( .A1(n9258), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9259) );
  NAND2_X1 U10902 ( .A1(n11767), .A2(n14145), .ZN(n9260) );
  NAND2_X1 U10903 ( .A1(n9261), .A2(n9260), .ZN(n9869) );
  NAND2_X1 U10904 ( .A1(n10395), .A2(n9869), .ZN(n9262) );
  OR2_X1 U10905 ( .A1(n9880), .A2(n9262), .ZN(n9266) );
  INV_X1 U10906 ( .A(n9767), .ZN(n14468) );
  NAND3_X1 U10907 ( .A1(n14468), .A2(n14466), .A3(n9748), .ZN(n9870) );
  NAND2_X1 U10908 ( .A1(n11614), .A2(n14145), .ZN(n9752) );
  INV_X1 U10909 ( .A(n9752), .ZN(n10079) );
  NAND2_X1 U10910 ( .A1(n10395), .A2(n11083), .ZN(n10082) );
  OR2_X1 U10911 ( .A1(n9755), .A2(n14145), .ZN(n9753) );
  INV_X1 U10912 ( .A(n11614), .ZN(n9742) );
  NAND2_X1 U10913 ( .A1(n11767), .A2(n9742), .ZN(n10078) );
  NOR2_X1 U10914 ( .A1(n9753), .A2(n10078), .ZN(n9872) );
  NAND2_X1 U10915 ( .A1(n10395), .A2(n9872), .ZN(n9263) );
  AND2_X1 U10916 ( .A1(n10082), .A2(n9263), .ZN(n9264) );
  OR2_X1 U10917 ( .A1(n9870), .A2(n9264), .ZN(n9265) );
  INV_X1 U10918 ( .A(n14464), .ZN(n9267) );
  NAND2_X1 U10919 ( .A1(n9268), .A2(n9267), .ZN(n9270) );
  NAND2_X1 U10920 ( .A1(n16239), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9269) );
  NAND2_X1 U10921 ( .A1(n9273), .A2(n9274), .ZN(n14469) );
  XNOR2_X2 U10922 ( .A(n9272), .B(n14470), .ZN(n9278) );
  XNOR2_X2 U10923 ( .A(n9275), .B(n9274), .ZN(n13927) );
  NAND2_X2 U10924 ( .A1(n9277), .A2(n9276), .ZN(n9537) );
  INV_X1 U10925 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n11234) );
  OR2_X1 U10926 ( .A1(n9537), .A2(n11234), .ZN(n9282) );
  INV_X1 U10927 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n11256) );
  OR2_X1 U10928 ( .A1(n9293), .A2(n11256), .ZN(n9281) );
  NAND2_X4 U10929 ( .A1(n13927), .A2(n9277), .ZN(n9571) );
  INV_X1 U10930 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n11438) );
  NAND2_X1 U10931 ( .A1(n7424), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n9279) );
  NAND2_X1 U10932 ( .A1(n9284), .A2(n9283), .ZN(n9286) );
  AND2_X1 U10933 ( .A1(n9286), .A2(n9285), .ZN(n10474) );
  OR2_X1 U10934 ( .A1(n9562), .A2(n10474), .ZN(n9291) );
  NAND2_X1 U10935 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n9287) );
  INV_X1 U10936 ( .A(n10475), .ZN(n11096) );
  OR2_X1 U10937 ( .A1(n10131), .A2(n10475), .ZN(n9289) );
  NAND2_X1 U10938 ( .A1(n9299), .A2(n11247), .ZN(n9945) );
  NAND2_X1 U10939 ( .A1(n9904), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n9297) );
  INV_X1 U10940 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10168) );
  OR2_X1 U10941 ( .A1(n9293), .A2(n10168), .ZN(n9296) );
  INV_X1 U10942 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n16044) );
  OR2_X1 U10943 ( .A1(n9537), .A2(n16044), .ZN(n9295) );
  INV_X1 U10944 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11477) );
  OR2_X1 U10945 ( .A1(n9571), .A2(n11477), .ZN(n9294) );
  XNOR2_X1 U10946 ( .A(n10303), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9298) );
  MUX2_X1 U10947 ( .A(n9298), .B(SI_0_), .S(n10431), .Z(n14477) );
  MUX2_X1 U10948 ( .A(P3_IR_REG_0__SCAN_IN), .B(n14477), .S(n7594), .Z(n16038)
         );
  NAND2_X1 U10949 ( .A1(n14059), .A2(n16038), .ZN(n11250) );
  NAND2_X1 U10950 ( .A1(n10057), .A2(n11250), .ZN(n9301) );
  INV_X1 U10951 ( .A(n9571), .ZN(n9302) );
  NAND2_X1 U10952 ( .A1(n9302), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n9307) );
  INV_X1 U10953 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10169) );
  INV_X1 U10954 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n16060) );
  OR2_X1 U10955 ( .A1(n9537), .A2(n16060), .ZN(n9305) );
  INV_X1 U10956 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n9303) );
  OR2_X1 U10957 ( .A1(n9587), .A2(n9303), .ZN(n9304) );
  NAND4_X2 U10958 ( .A1(n9307), .A2(n9306), .A3(n9305), .A4(n9304), .ZN(n14058) );
  XNOR2_X1 U10959 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n9308) );
  XNOR2_X1 U10960 ( .A(n9309), .B(n9308), .ZN(n10472) );
  NAND2_X1 U10961 ( .A1(n16051), .A2(n9948), .ZN(n9311) );
  INV_X1 U10962 ( .A(n16049), .ZN(n9772) );
  OR2_X1 U10963 ( .A1(n14058), .A2(n9772), .ZN(n9310) );
  NAND2_X1 U10964 ( .A1(n9904), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n9315) );
  INV_X1 U10965 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10175) );
  OR2_X1 U10966 ( .A1(n9537), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n9313) );
  INV_X1 U10967 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10176) );
  OR2_X1 U10968 ( .A1(n9571), .A2(n10176), .ZN(n9312) );
  XNOR2_X1 U10969 ( .A(n9316), .B(P3_IR_REG_3__SCAN_IN), .ZN(n11171) );
  XNOR2_X1 U10970 ( .A(n10408), .B(P2_DATAO_REG_3__SCAN_IN), .ZN(n9317) );
  XNOR2_X1 U10971 ( .A(n9318), .B(n9317), .ZN(n10438) );
  OR2_X1 U10972 ( .A1(n9562), .A2(n10438), .ZN(n9320) );
  OR2_X1 U10973 ( .A1(n9917), .A2(SI_3_), .ZN(n9319) );
  OAI211_X1 U10974 ( .C1(n11171), .C2(n10131), .A(n9320), .B(n9319), .ZN(
        n11522) );
  OR2_X1 U10975 ( .A1(n14057), .A2(n11522), .ZN(n9958) );
  NAND2_X1 U10976 ( .A1(n14057), .A2(n11522), .ZN(n9953) );
  INV_X1 U10977 ( .A(n11522), .ZN(n11431) );
  NAND2_X1 U10978 ( .A1(n14057), .A2(n11431), .ZN(n9322) );
  NAND2_X1 U10979 ( .A1(n10385), .A2(n9322), .ZN(n11572) );
  NAND2_X1 U10980 ( .A1(n9717), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n9328) );
  INV_X1 U10981 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n9323) );
  OR2_X1 U10982 ( .A1(n9293), .A2(n9323), .ZN(n9327) );
  NOR2_X1 U10983 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n9342) );
  AND2_X1 U10984 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n9324) );
  NOR2_X1 U10985 ( .A1(n9342), .A2(n9324), .ZN(n11725) );
  OR2_X1 U10986 ( .A1(n9551), .A2(n11725), .ZN(n9326) );
  INV_X1 U10987 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11634) );
  OR2_X1 U10988 ( .A1(n9571), .A2(n11634), .ZN(n9325) );
  XNOR2_X1 U10989 ( .A(n9331), .B(P3_IR_REG_4__SCAN_IN), .ZN(n10183) );
  NAND2_X1 U10990 ( .A1(n9333), .A2(n9332), .ZN(n9334) );
  AND2_X1 U10991 ( .A1(n9335), .A2(n9334), .ZN(n10442) );
  OR2_X1 U10992 ( .A1(n9562), .A2(n10442), .ZN(n9337) );
  OR2_X1 U10993 ( .A1(n9917), .A2(SI_4_), .ZN(n9336) );
  OAI211_X1 U10994 ( .C1(n10183), .C2(n10131), .A(n9337), .B(n9336), .ZN(
        n11727) );
  NAND2_X1 U10995 ( .A1(n11806), .A2(n11727), .ZN(n9960) );
  INV_X1 U10996 ( .A(n11578), .ZN(n11574) );
  NAND2_X1 U10997 ( .A1(n11806), .A2(n7933), .ZN(n9339) );
  NAND2_X1 U10998 ( .A1(n9717), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n9348) );
  INV_X1 U10999 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n9340) );
  OR2_X1 U11000 ( .A1(n9293), .A2(n9340), .ZN(n9347) );
  INV_X1 U11001 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n9341) );
  NAND2_X1 U11002 ( .A1(n9342), .A2(n9341), .ZN(n9360) );
  OR2_X1 U11003 ( .A1(n9342), .A2(n9341), .ZN(n9343) );
  AND2_X1 U11004 ( .A1(n9360), .A2(n9343), .ZN(n16093) );
  OR2_X1 U11005 ( .A1(n9537), .A2(n16093), .ZN(n9346) );
  INV_X1 U11006 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n9344) );
  OR2_X1 U11007 ( .A1(n9908), .A2(n9344), .ZN(n9345) );
  NAND4_X1 U11008 ( .A1(n9348), .A2(n9347), .A3(n9346), .A4(n9345), .ZN(n11575) );
  NAND2_X1 U11009 ( .A1(n9350), .A2(n9349), .ZN(n9366) );
  NAND2_X1 U11010 ( .A1(n9366), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9351) );
  XNOR2_X1 U11011 ( .A(n9351), .B(P3_IR_REG_5__SCAN_IN), .ZN(n10187) );
  NAND2_X1 U11012 ( .A1(n9353), .A2(n9352), .ZN(n9355) );
  AND2_X1 U11013 ( .A1(n9355), .A2(n9354), .ZN(n10435) );
  OR2_X1 U11014 ( .A1(n9562), .A2(n10435), .ZN(n9357) );
  OR2_X1 U11015 ( .A1(n9917), .A2(SI_5_), .ZN(n9356) );
  OAI211_X1 U11016 ( .C1(n10187), .C2(n7594), .A(n9357), .B(n9356), .ZN(n11810) );
  OR2_X1 U11017 ( .A1(n11575), .A2(n11810), .ZN(n9963) );
  NAND2_X1 U11018 ( .A1(n11575), .A2(n11810), .ZN(n9964) );
  NAND2_X1 U11019 ( .A1(n9963), .A2(n9964), .ZN(n11804) );
  INV_X1 U11020 ( .A(n11810), .ZN(n16097) );
  OR2_X1 U11021 ( .A1(n11575), .A2(n16097), .ZN(n9358) );
  NAND2_X1 U11022 ( .A1(n9718), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n9365) );
  INV_X1 U11023 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n9359) );
  OR2_X1 U11024 ( .A1(n9587), .A2(n9359), .ZN(n9364) );
  NAND2_X1 U11025 ( .A1(n9360), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9361) );
  AND2_X1 U11026 ( .A1(n9379), .A2(n9361), .ZN(n11951) );
  OR2_X1 U11027 ( .A1(n9537), .A2(n11951), .ZN(n9363) );
  INV_X1 U11028 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11759) );
  OR2_X1 U11029 ( .A1(n9571), .A2(n11759), .ZN(n9362) );
  NAND4_X1 U11030 ( .A1(n9365), .A2(n9364), .A3(n9363), .A4(n9362), .ZN(n14056) );
  NOR2_X1 U11031 ( .A1(n9366), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n9369) );
  OR2_X1 U11032 ( .A1(n9369), .A2(n9330), .ZN(n9367) );
  MUX2_X1 U11033 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9367), .S(
        P3_IR_REG_6__SCAN_IN), .Z(n9370) );
  INV_X1 U11034 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n9368) );
  NAND2_X1 U11035 ( .A1(n9369), .A2(n9368), .ZN(n9400) );
  NAND2_X1 U11036 ( .A1(n9370), .A2(n9400), .ZN(n15984) );
  INV_X1 U11037 ( .A(SI_6_), .ZN(n10433) );
  OR2_X1 U11038 ( .A1(n9917), .A2(n10433), .ZN(n9374) );
  XNOR2_X1 U11039 ( .A(n9372), .B(n9371), .ZN(n10434) );
  OR2_X1 U11040 ( .A1(n9562), .A2(n10434), .ZN(n9373) );
  OAI211_X1 U11041 ( .C1(n7594), .C2(n15984), .A(n9374), .B(n9373), .ZN(n16101) );
  XNOR2_X1 U11042 ( .A(n14056), .B(n16101), .ZN(n11754) );
  NAND2_X1 U11043 ( .A1(n14056), .A2(n16101), .ZN(n9377) );
  NAND2_X1 U11044 ( .A1(n11757), .A2(n9377), .ZN(n11843) );
  NAND2_X1 U11045 ( .A1(n9717), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n9385) );
  INV_X1 U11046 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n9378) );
  OR2_X1 U11047 ( .A1(n9293), .A2(n9378), .ZN(n9384) );
  AND2_X1 U11048 ( .A1(n9379), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9380) );
  NOR2_X1 U11049 ( .A1(n9392), .A2(n9380), .ZN(n12056) );
  OR2_X1 U11050 ( .A1(n9551), .A2(n12056), .ZN(n9383) );
  INV_X1 U11051 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n9381) );
  OR2_X1 U11052 ( .A1(n9908), .A2(n9381), .ZN(n9382) );
  NAND4_X1 U11053 ( .A1(n9385), .A2(n9384), .A3(n9383), .A4(n9382), .ZN(n14054) );
  NAND2_X1 U11054 ( .A1(n9400), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9386) );
  XNOR2_X1 U11055 ( .A(n9388), .B(n9387), .ZN(n10467) );
  OR2_X1 U11056 ( .A1(n9562), .A2(n10467), .ZN(n9390) );
  OR2_X1 U11057 ( .A1(n9917), .A2(SI_7_), .ZN(n9389) );
  OAI211_X1 U11058 ( .C1(n10466), .C2(n7594), .A(n9390), .B(n9389), .ZN(n11995) );
  OR2_X1 U11059 ( .A1(n14054), .A2(n11995), .ZN(n9970) );
  NAND2_X1 U11060 ( .A1(n14054), .A2(n11995), .ZN(n9971) );
  NAND2_X1 U11061 ( .A1(n9970), .A2(n9971), .ZN(n11842) );
  INV_X1 U11062 ( .A(n11995), .ZN(n12053) );
  NAND2_X1 U11063 ( .A1(n14054), .A2(n12053), .ZN(n9391) );
  NAND2_X1 U11064 ( .A1(n9717), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n9397) );
  INV_X1 U11065 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n10149) );
  OR2_X1 U11066 ( .A1(n9293), .A2(n10149), .ZN(n9396) );
  NOR2_X1 U11067 ( .A1(n9392), .A2(n11376), .ZN(n9393) );
  OR2_X1 U11068 ( .A1(n9551), .A2(n7460), .ZN(n9395) );
  INV_X1 U11069 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n10115) );
  OR2_X1 U11070 ( .A1(n9571), .A2(n10115), .ZN(n9394) );
  NAND4_X1 U11071 ( .A1(n9397), .A2(n9396), .A3(n9395), .A4(n9394), .ZN(n14053) );
  XNOR2_X1 U11072 ( .A(n9399), .B(n9398), .ZN(n10481) );
  OR2_X1 U11073 ( .A1(n9562), .A2(n10481), .ZN(n9404) );
  INV_X1 U11074 ( .A(SI_8_), .ZN(n10480) );
  OR2_X1 U11075 ( .A1(n9917), .A2(n10480), .ZN(n9403) );
  NAND2_X1 U11076 ( .A1(n9415), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9401) );
  NAND2_X1 U11077 ( .A1(n9581), .A2(n10479), .ZN(n9402) );
  XNOR2_X1 U11078 ( .A(n14053), .B(n12075), .ZN(n11957) );
  NAND2_X1 U11079 ( .A1(n9717), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n9412) );
  INV_X1 U11080 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n9405) );
  OR2_X1 U11081 ( .A1(n9293), .A2(n9405), .ZN(n9411) );
  NAND2_X1 U11082 ( .A1(n9406), .A2(n12403), .ZN(n9423) );
  OR2_X1 U11083 ( .A1(n9406), .A2(n12403), .ZN(n9407) );
  AND2_X1 U11084 ( .A1(n9423), .A2(n9407), .ZN(n12402) );
  OR2_X1 U11085 ( .A1(n9537), .A2(n12402), .ZN(n9410) );
  INV_X1 U11086 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n9408) );
  OR2_X1 U11087 ( .A1(n9908), .A2(n9408), .ZN(n9409) );
  NAND4_X1 U11088 ( .A1(n9412), .A2(n9411), .A3(n9410), .A4(n9409), .ZN(n14052) );
  XNOR2_X1 U11089 ( .A(n9414), .B(n9413), .ZN(n10476) );
  OR2_X1 U11090 ( .A1(n9562), .A2(n10476), .ZN(n9419) );
  OR2_X1 U11091 ( .A1(n9917), .A2(SI_9_), .ZN(n9418) );
  OAI21_X1 U11092 ( .B1(n9415), .B2(P3_IR_REG_8__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9416) );
  XNOR2_X1 U11093 ( .A(n9416), .B(P3_IR_REG_9__SCAN_IN), .ZN(n16019) );
  INV_X1 U11094 ( .A(n16019), .ZN(n10478) );
  NAND2_X1 U11095 ( .A1(n9581), .A2(n10478), .ZN(n9417) );
  XNOR2_X1 U11096 ( .A(n14052), .B(n12440), .ZN(n10063) );
  NAND2_X1 U11097 ( .A1(n14052), .A2(n12440), .ZN(n9421) );
  NAND2_X1 U11098 ( .A1(n12287), .A2(n9421), .ZN(n12321) );
  NAND2_X1 U11099 ( .A1(n9718), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n9429) );
  INV_X1 U11100 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n9422) );
  OR2_X1 U11101 ( .A1(n9571), .A2(n9422), .ZN(n9428) );
  NAND2_X1 U11102 ( .A1(n9423), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9424) );
  AND2_X1 U11103 ( .A1(n9449), .A2(n9424), .ZN(n12329) );
  OR2_X1 U11104 ( .A1(n9551), .A2(n12329), .ZN(n9427) );
  INV_X1 U11105 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n9425) );
  OR2_X1 U11106 ( .A1(n9587), .A2(n9425), .ZN(n9426) );
  NAND4_X1 U11107 ( .A1(n9429), .A2(n9428), .A3(n9427), .A4(n9426), .ZN(n14051) );
  OR2_X1 U11108 ( .A1(n9431), .A2(n9430), .ZN(n9432) );
  NAND2_X1 U11109 ( .A1(n9433), .A2(n9432), .ZN(n10470) );
  NAND2_X1 U11110 ( .A1(n10470), .A2(n9916), .ZN(n9438) );
  NAND2_X1 U11111 ( .A1(n9435), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9434) );
  MUX2_X1 U11112 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9434), .S(
        P3_IR_REG_10__SCAN_IN), .Z(n9436) );
  OR2_X1 U11113 ( .A1(n9435), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n9459) );
  NAND2_X1 U11114 ( .A1(n9436), .A2(n9459), .ZN(n10471) );
  NAND2_X1 U11115 ( .A1(n9581), .A2(n10471), .ZN(n9437) );
  OAI211_X1 U11116 ( .C1(SI_10_), .C2(n9917), .A(n9438), .B(n9437), .ZN(n12473) );
  OR2_X1 U11117 ( .A1(n14051), .A2(n12473), .ZN(n9983) );
  NAND2_X1 U11118 ( .A1(n14051), .A2(n12473), .ZN(n9984) );
  NAND2_X1 U11119 ( .A1(n9983), .A2(n9984), .ZN(n12325) );
  INV_X1 U11120 ( .A(n12473), .ZN(n9439) );
  NAND2_X1 U11121 ( .A1(n14051), .A2(n9439), .ZN(n9440) );
  OR2_X1 U11122 ( .A1(n9442), .A2(n9441), .ZN(n9443) );
  NAND2_X1 U11123 ( .A1(n9444), .A2(n9443), .ZN(n10482) );
  NAND2_X1 U11124 ( .A1(n10482), .A2(n9916), .ZN(n9447) );
  NAND2_X1 U11125 ( .A1(n9459), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9445) );
  XNOR2_X1 U11126 ( .A(n9445), .B(P3_IR_REG_11__SCAN_IN), .ZN(n10155) );
  AOI22_X1 U11127 ( .A1(n9686), .A2(n12973), .B1(n9581), .B2(n12153), .ZN(
        n9446) );
  NAND2_X1 U11128 ( .A1(n9717), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n9454) );
  INV_X1 U11129 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n9448) );
  OR2_X1 U11130 ( .A1(n9293), .A2(n9448), .ZN(n9453) );
  NAND2_X1 U11131 ( .A1(n9449), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9450) );
  AND2_X1 U11132 ( .A1(n9463), .A2(n9450), .ZN(n12647) );
  OR2_X1 U11133 ( .A1(n9537), .A2(n12647), .ZN(n9452) );
  INV_X1 U11134 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n12500) );
  OR2_X1 U11135 ( .A1(n9908), .A2(n12500), .ZN(n9451) );
  NAND4_X1 U11136 ( .A1(n9454), .A2(n9453), .A3(n9452), .A4(n9451), .ZN(n12322) );
  OR2_X1 U11137 ( .A1(n12712), .A2(n12322), .ZN(n9800) );
  NAND2_X1 U11138 ( .A1(n12712), .A2(n12322), .ZN(n9799) );
  OR2_X1 U11139 ( .A1(n9456), .A2(n9455), .ZN(n9457) );
  NAND2_X1 U11140 ( .A1(n9458), .A2(n9457), .ZN(n10489) );
  NAND2_X1 U11141 ( .A1(n10489), .A2(n9916), .ZN(n9462) );
  NOR2_X1 U11142 ( .A1(n9459), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n9475) );
  OR2_X1 U11143 ( .A1(n9475), .A2(n9330), .ZN(n9460) );
  XNOR2_X1 U11144 ( .A(n9460), .B(n9474), .ZN(n12131) );
  AOI22_X1 U11145 ( .A1(n9686), .A2(n12970), .B1(n9581), .B2(n12131), .ZN(
        n9461) );
  NAND2_X1 U11146 ( .A1(n9462), .A2(n9461), .ZN(n16232) );
  NAND2_X1 U11147 ( .A1(n9717), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n9469) );
  INV_X1 U11148 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n16237) );
  OR2_X1 U11149 ( .A1(n9293), .A2(n16237), .ZN(n9468) );
  AND2_X1 U11150 ( .A1(n9463), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9464) );
  NOR2_X1 U11151 ( .A1(n9481), .A2(n9464), .ZN(n13198) );
  OR2_X1 U11152 ( .A1(n9551), .A2(n13198), .ZN(n9467) );
  INV_X1 U11153 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n9465) );
  OR2_X1 U11154 ( .A1(n9571), .A2(n9465), .ZN(n9466) );
  NOR2_X1 U11155 ( .A1(n16232), .A2(n13230), .ZN(n9470) );
  NAND2_X1 U11156 ( .A1(n9471), .A2(n10725), .ZN(n9472) );
  NAND2_X1 U11157 ( .A1(n9473), .A2(n9472), .ZN(n10600) );
  NAND2_X1 U11158 ( .A1(n10600), .A2(n9916), .ZN(n9478) );
  INV_X1 U11159 ( .A(SI_13_), .ZN(n12971) );
  NAND2_X1 U11160 ( .A1(n9475), .A2(n9474), .ZN(n9491) );
  NAND2_X1 U11161 ( .A1(n9491), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9476) );
  XNOR2_X1 U11162 ( .A(n9476), .B(P3_IR_REG_13__SCAN_IN), .ZN(n10210) );
  INV_X1 U11163 ( .A(n10210), .ZN(n14072) );
  AOI22_X1 U11164 ( .A1(n9686), .A2(n12971), .B1(n9581), .B2(n14072), .ZN(
        n9477) );
  NAND2_X1 U11165 ( .A1(n9478), .A2(n9477), .ZN(n13235) );
  NAND2_X1 U11166 ( .A1(n9717), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n9486) );
  INV_X1 U11167 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n9479) );
  OR2_X1 U11168 ( .A1(n9293), .A2(n9479), .ZN(n9485) );
  INV_X1 U11169 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n14066) );
  OR2_X1 U11170 ( .A1(n9908), .A2(n14066), .ZN(n9484) );
  OR2_X1 U11171 ( .A1(n9481), .A2(n9480), .ZN(n9482) );
  NAND2_X1 U11172 ( .A1(n9481), .A2(n9480), .ZN(n9499) );
  AND2_X1 U11173 ( .A1(n9482), .A2(n9499), .ZN(n13181) );
  OR2_X1 U11174 ( .A1(n9537), .A2(n13181), .ZN(n9483) );
  AND2_X1 U11175 ( .A1(n13235), .A2(n12601), .ZN(n9812) );
  OR2_X1 U11176 ( .A1(n13235), .A2(n12601), .ZN(n9811) );
  OR2_X1 U11177 ( .A1(n9488), .A2(n9487), .ZN(n9489) );
  NAND2_X1 U11178 ( .A1(n9490), .A2(n9489), .ZN(n10728) );
  NAND2_X1 U11179 ( .A1(n10728), .A2(n9916), .ZN(n9497) );
  INV_X1 U11180 ( .A(n9514), .ZN(n9495) );
  NAND2_X1 U11181 ( .A1(n9492), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9493) );
  MUX2_X1 U11182 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9493), .S(
        P3_IR_REG_14__SCAN_IN), .Z(n9494) );
  AOI22_X1 U11183 ( .A1(n9686), .A2(n7846), .B1(n9581), .B2(n10729), .ZN(n9496) );
  NAND2_X1 U11184 ( .A1(n9497), .A2(n9496), .ZN(n14422) );
  NAND2_X1 U11185 ( .A1(n9718), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n9505) );
  INV_X1 U11186 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n9498) );
  OR2_X1 U11187 ( .A1(n9587), .A2(n9498), .ZN(n9504) );
  NAND2_X1 U11188 ( .A1(n9499), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9500) );
  AND2_X1 U11189 ( .A1(n9518), .A2(n9500), .ZN(n13190) );
  OR2_X1 U11190 ( .A1(n9551), .A2(n13190), .ZN(n9503) );
  INV_X1 U11191 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n9501) );
  OR2_X1 U11192 ( .A1(n9571), .A2(n9501), .ZN(n9502) );
  NAND4_X1 U11193 ( .A1(n9505), .A2(n9504), .A3(n9503), .A4(n9502), .ZN(n14048) );
  OR2_X1 U11194 ( .A1(n14422), .A2(n14048), .ZN(n9998) );
  NAND2_X1 U11195 ( .A1(n14422), .A2(n14048), .ZN(n10002) );
  NAND2_X1 U11196 ( .A1(n9998), .A2(n10002), .ZN(n13188) );
  NAND2_X1 U11197 ( .A1(n13186), .A2(n13188), .ZN(n9507) );
  INV_X1 U11198 ( .A(n14048), .ZN(n13211) );
  OR2_X1 U11199 ( .A1(n14422), .A2(n13211), .ZN(n9506) );
  NAND2_X1 U11200 ( .A1(n9507), .A2(n9506), .ZN(n13208) );
  OR2_X1 U11201 ( .A1(n9509), .A2(n9508), .ZN(n9510) );
  NAND2_X1 U11202 ( .A1(n9511), .A2(n9510), .ZN(n10935) );
  NAND2_X1 U11203 ( .A1(n10935), .A2(n9916), .ZN(n9517) );
  OR2_X1 U11204 ( .A1(n9514), .A2(n9330), .ZN(n9512) );
  MUX2_X1 U11205 ( .A(n9512), .B(P3_IR_REG_31__SCAN_IN), .S(n9513), .Z(n9515)
         );
  NAND2_X1 U11206 ( .A1(n9514), .A2(n9513), .ZN(n9546) );
  NAND2_X1 U11207 ( .A1(n9515), .A2(n9546), .ZN(n14085) );
  AOI22_X1 U11208 ( .A1(n9686), .A2(n10936), .B1(n9581), .B2(n14085), .ZN(
        n9516) );
  NAND2_X1 U11209 ( .A1(n9717), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n9523) );
  INV_X1 U11210 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n14416) );
  OR2_X1 U11211 ( .A1(n9293), .A2(n14416), .ZN(n9522) );
  AND2_X1 U11212 ( .A1(n9518), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9519) );
  NOR2_X1 U11213 ( .A1(n9534), .A2(n9519), .ZN(n14037) );
  OR2_X1 U11214 ( .A1(n9537), .A2(n14037), .ZN(n9521) );
  INV_X1 U11215 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n14078) );
  OR2_X1 U11216 ( .A1(n9908), .A2(n14078), .ZN(n9520) );
  NAND4_X1 U11217 ( .A1(n9523), .A2(n9522), .A3(n9521), .A4(n9520), .ZN(n14047) );
  OR2_X1 U11218 ( .A1(n14463), .A2(n14047), .ZN(n10006) );
  NAND2_X1 U11219 ( .A1(n14463), .A2(n14047), .ZN(n10007) );
  NAND2_X1 U11220 ( .A1(n10006), .A2(n10007), .ZN(n13209) );
  INV_X1 U11221 ( .A(n14047), .ZN(n14331) );
  OR2_X1 U11222 ( .A1(n14463), .A2(n14331), .ZN(n9524) );
  OR2_X1 U11223 ( .A1(n9527), .A2(n9526), .ZN(n9528) );
  NAND2_X1 U11224 ( .A1(n9529), .A2(n9528), .ZN(n11068) );
  OR2_X1 U11225 ( .A1(n11068), .A2(n9562), .ZN(n9532) );
  NAND2_X1 U11226 ( .A1(n9546), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9530) );
  XNOR2_X1 U11227 ( .A(n9530), .B(P3_IR_REG_16__SCAN_IN), .ZN(n14094) );
  AOI22_X1 U11228 ( .A1(n9686), .A2(SI_16_), .B1(n9581), .B2(n14094), .ZN(
        n9531) );
  NAND2_X1 U11229 ( .A1(n9532), .A2(n9531), .ZN(n9944) );
  NAND2_X1 U11230 ( .A1(n9717), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n9541) );
  INV_X1 U11231 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n14412) );
  OR2_X1 U11232 ( .A1(n9293), .A2(n14412), .ZN(n9540) );
  INV_X1 U11233 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n10229) );
  OR2_X1 U11234 ( .A1(n9908), .A2(n10229), .ZN(n9539) );
  NOR2_X1 U11235 ( .A1(n9534), .A2(n9533), .ZN(n9535) );
  OR2_X1 U11236 ( .A1(n9552), .A2(n9535), .ZN(n14335) );
  INV_X1 U11237 ( .A(n14335), .ZN(n9536) );
  OR2_X1 U11238 ( .A1(n9537), .A2(n9536), .ZN(n9538) );
  NAND4_X1 U11239 ( .A1(n9541), .A2(n9540), .A3(n9539), .A4(n9538), .ZN(n14046) );
  OR2_X1 U11240 ( .A1(n9944), .A2(n14046), .ZN(n10008) );
  NAND2_X1 U11241 ( .A1(n9944), .A2(n14046), .ZN(n10014) );
  NAND2_X1 U11242 ( .A1(n10008), .A2(n10014), .ZN(n14333) );
  OR2_X1 U11243 ( .A1(n9543), .A2(n9542), .ZN(n9544) );
  NAND2_X1 U11244 ( .A1(n9545), .A2(n9544), .ZN(n11258) );
  NAND2_X1 U11245 ( .A1(n11258), .A2(n9916), .ZN(n9550) );
  OAI21_X1 U11246 ( .B1(n9546), .B2(P3_IR_REG_16__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9548) );
  INV_X1 U11247 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n9547) );
  XNOR2_X1 U11248 ( .A(n9548), .B(n9547), .ZN(n14129) );
  AOI22_X1 U11249 ( .A1(n9686), .A2(n12737), .B1(n9581), .B2(n14129), .ZN(
        n9549) );
  OR2_X1 U11250 ( .A1(n9552), .A2(n13020), .ZN(n9553) );
  NAND2_X1 U11251 ( .A1(n9568), .A2(n9553), .ZN(n14321) );
  NAND2_X1 U11252 ( .A1(n9708), .A2(n14321), .ZN(n9557) );
  INV_X1 U11253 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n14453) );
  OR2_X1 U11254 ( .A1(n9587), .A2(n14453), .ZN(n9556) );
  INV_X1 U11255 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n14408) );
  OR2_X1 U11256 ( .A1(n9293), .A2(n14408), .ZN(n9555) );
  INV_X1 U11257 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14110) );
  OR2_X1 U11258 ( .A1(n9908), .A2(n14110), .ZN(n9554) );
  NAND4_X1 U11259 ( .A1(n9557), .A2(n9556), .A3(n9555), .A4(n9554), .ZN(n14306) );
  OR2_X1 U11260 ( .A1(n14455), .A2(n14306), .ZN(n10019) );
  NAND2_X1 U11261 ( .A1(n14455), .A2(n14306), .ZN(n9943) );
  OR2_X1 U11262 ( .A1(n9559), .A2(n9558), .ZN(n9560) );
  NAND2_X1 U11263 ( .A1(n9561), .A2(n9560), .ZN(n11336) );
  OR2_X1 U11264 ( .A1(n11336), .A2(n9562), .ZN(n9567) );
  NAND2_X1 U11265 ( .A1(n9563), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9564) );
  MUX2_X1 U11266 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9564), .S(
        P3_IR_REG_18__SCAN_IN), .Z(n9565) );
  NAND2_X1 U11267 ( .A1(n9565), .A2(n9258), .ZN(n14148) );
  INV_X1 U11268 ( .A(n14148), .ZN(n14139) );
  AOI22_X1 U11269 ( .A1(n9686), .A2(SI_18_), .B1(n9581), .B2(n14139), .ZN(
        n9566) );
  NAND2_X1 U11270 ( .A1(n9567), .A2(n9566), .ZN(n14016) );
  NAND2_X1 U11271 ( .A1(n9568), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9569) );
  NAND2_X1 U11272 ( .A1(n9584), .A2(n9569), .ZN(n14310) );
  NAND2_X1 U11273 ( .A1(n9708), .A2(n14310), .ZN(n9575) );
  INV_X1 U11274 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n14449) );
  OR2_X1 U11275 ( .A1(n9587), .A2(n14449), .ZN(n9574) );
  INV_X1 U11276 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n14404) );
  OR2_X1 U11277 ( .A1(n9293), .A2(n14404), .ZN(n9573) );
  INV_X1 U11278 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n9570) );
  OR2_X1 U11279 ( .A1(n9571), .A2(n9570), .ZN(n9572) );
  OR2_X1 U11280 ( .A1(n14016), .A2(n14316), .ZN(n10022) );
  NAND2_X1 U11281 ( .A1(n14016), .A2(n14316), .ZN(n10020) );
  NAND2_X1 U11282 ( .A1(n10022), .A2(n10020), .ZN(n14302) );
  INV_X1 U11283 ( .A(n14302), .ZN(n9576) );
  INV_X1 U11284 ( .A(n14306), .ZN(n14330) );
  NOR2_X1 U11285 ( .A1(n14455), .A2(n14330), .ZN(n14300) );
  OR2_X1 U11286 ( .A1(n14016), .A2(n14290), .ZN(n9577) );
  XNOR2_X1 U11287 ( .A(n9578), .B(P2_DATAO_REG_19__SCAN_IN), .ZN(n9579) );
  XNOR2_X1 U11288 ( .A(n9580), .B(n9579), .ZN(n11482) );
  NAND2_X1 U11289 ( .A1(n11482), .A2(n9916), .ZN(n9583) );
  AOI22_X1 U11290 ( .A1(n9686), .A2(SI_19_), .B1(n9581), .B2(n9927), .ZN(n9582) );
  NAND2_X1 U11291 ( .A1(n9583), .A2(n9582), .ZN(n14397) );
  INV_X1 U11292 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n9593) );
  AND2_X1 U11293 ( .A1(n9584), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9585) );
  NOR2_X2 U11294 ( .A1(n9584), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9601) );
  OR2_X1 U11295 ( .A1(n9585), .A2(n9601), .ZN(n14295) );
  NAND2_X1 U11296 ( .A1(n14295), .A2(n9708), .ZN(n9592) );
  INV_X1 U11297 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n9586) );
  OR2_X1 U11298 ( .A1(n9587), .A2(n9586), .ZN(n9590) );
  INV_X1 U11299 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n9588) );
  OR2_X1 U11300 ( .A1(n9293), .A2(n9588), .ZN(n9589) );
  AND2_X1 U11301 ( .A1(n9590), .A2(n9589), .ZN(n9591) );
  NAND2_X1 U11302 ( .A1(n14397), .A2(n14305), .ZN(n9594) );
  NAND2_X1 U11303 ( .A1(n14289), .A2(n9594), .ZN(n9596) );
  OR2_X1 U11304 ( .A1(n14397), .A2(n14305), .ZN(n9595) );
  XNOR2_X1 U11305 ( .A(n9598), .B(n9597), .ZN(n11611) );
  NAND2_X1 U11306 ( .A1(n11611), .A2(n9916), .ZN(n9600) );
  OR2_X1 U11307 ( .A1(n9917), .A2(n11612), .ZN(n9599) );
  INV_X1 U11308 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n12802) );
  NOR2_X1 U11309 ( .A1(n9601), .A2(n12802), .ZN(n9602) );
  OR2_X1 U11310 ( .A1(n9611), .A2(n9602), .ZN(n14282) );
  NAND2_X1 U11311 ( .A1(n14282), .A2(n9708), .ZN(n9605) );
  AOI22_X1 U11312 ( .A1(n9717), .A2(P3_REG0_REG_20__SCAN_IN), .B1(n9718), .B2(
        P3_REG1_REG_20__SCAN_IN), .ZN(n9604) );
  NAND2_X1 U11313 ( .A1(n9302), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n9603) );
  NAND2_X1 U11314 ( .A1(n14389), .A2(n14268), .ZN(n10028) );
  NAND2_X1 U11315 ( .A1(n14389), .A2(n14383), .ZN(n9606) );
  XNOR2_X1 U11316 ( .A(n9608), .B(n9607), .ZN(n11764) );
  NAND2_X1 U11317 ( .A1(n11764), .A2(n9916), .ZN(n9610) );
  INV_X1 U11318 ( .A(SI_21_), .ZN(n11766) );
  OR2_X1 U11319 ( .A1(n9917), .A2(n11766), .ZN(n9609) );
  INV_X1 U11320 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n9615) );
  INV_X1 U11321 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n12787) );
  OR2_X1 U11322 ( .A1(n9611), .A2(n12787), .ZN(n9612) );
  NAND2_X1 U11323 ( .A1(n9636), .A2(n9612), .ZN(n14266) );
  NAND2_X1 U11324 ( .A1(n14266), .A2(n9708), .ZN(n9614) );
  AOI22_X1 U11325 ( .A1(n9717), .A2(P3_REG0_REG_21__SCAN_IN), .B1(n9718), .B2(
        P3_REG1_REG_21__SCAN_IN), .ZN(n9613) );
  OAI211_X1 U11326 ( .C1(n9908), .C2(n9615), .A(n9614), .B(n9613), .ZN(n14045)
         );
  OR2_X1 U11327 ( .A1(n14385), .A2(n14045), .ZN(n9616) );
  AND2_X1 U11328 ( .A1(n14385), .A2(n14045), .ZN(n9843) );
  AOI21_X2 U11329 ( .B1(n14264), .B2(n9616), .A(n9843), .ZN(n14251) );
  OR2_X1 U11330 ( .A1(n9618), .A2(n9617), .ZN(n9619) );
  NAND2_X1 U11331 ( .A1(n9620), .A2(n9619), .ZN(n11796) );
  NAND2_X1 U11332 ( .A1(n11796), .A2(n9916), .ZN(n9623) );
  OR2_X1 U11333 ( .A1(n9917), .A2(n9621), .ZN(n9622) );
  XNOR2_X1 U11334 ( .A(n9636), .B(P3_REG3_REG_22__SCAN_IN), .ZN(n14257) );
  NAND2_X1 U11335 ( .A1(n14257), .A2(n9708), .ZN(n9628) );
  INV_X1 U11336 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n14259) );
  NAND2_X1 U11337 ( .A1(n9717), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n9625) );
  NAND2_X1 U11338 ( .A1(n9718), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n9624) );
  OAI211_X1 U11339 ( .C1(n14259), .C2(n9908), .A(n9625), .B(n9624), .ZN(n9626)
         );
  INV_X1 U11340 ( .A(n9626), .ZN(n9627) );
  OR2_X1 U11341 ( .A1(n14377), .A2(n14244), .ZN(n10035) );
  NAND2_X1 U11342 ( .A1(n14377), .A2(n14244), .ZN(n10036) );
  NAND2_X1 U11343 ( .A1(n10035), .A2(n10036), .ZN(n14250) );
  OR2_X1 U11344 ( .A1(n14377), .A2(n14371), .ZN(n9629) );
  OR2_X1 U11345 ( .A1(n9631), .A2(n9630), .ZN(n9632) );
  NAND2_X1 U11346 ( .A1(n9633), .A2(n9632), .ZN(n11952) );
  NAND2_X1 U11347 ( .A1(n11952), .A2(n9916), .ZN(n9635) );
  OR2_X1 U11348 ( .A1(n9917), .A2(n11955), .ZN(n9634) );
  NAND2_X1 U11349 ( .A1(n9637), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9638) );
  NAND2_X1 U11350 ( .A1(n9648), .A2(n9638), .ZN(n14242) );
  NAND2_X1 U11351 ( .A1(n14242), .A2(n9708), .ZN(n9644) );
  INV_X1 U11352 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n9641) );
  NAND2_X1 U11353 ( .A1(n9717), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n9640) );
  NAND2_X1 U11354 ( .A1(n9718), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n9639) );
  OAI211_X1 U11355 ( .C1(n9641), .C2(n9908), .A(n9640), .B(n9639), .ZN(n9642)
         );
  INV_X1 U11356 ( .A(n9642), .ZN(n9643) );
  NAND2_X1 U11357 ( .A1(n14372), .A2(n14252), .ZN(n10040) );
  XNOR2_X1 U11358 ( .A(n9645), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n12380) );
  NAND2_X1 U11359 ( .A1(n12380), .A2(n9916), .ZN(n9647) );
  INV_X1 U11360 ( .A(SI_24_), .ZN(n12381) );
  OR2_X1 U11361 ( .A1(n9917), .A2(n12381), .ZN(n9646) );
  INV_X1 U11362 ( .A(n9663), .ZN(n9650) );
  NAND2_X1 U11363 ( .A1(n9648), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9649) );
  NAND2_X1 U11364 ( .A1(n9650), .A2(n9649), .ZN(n14226) );
  NAND2_X1 U11365 ( .A1(n14226), .A2(n9708), .ZN(n9656) );
  INV_X1 U11366 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n9653) );
  NAND2_X1 U11367 ( .A1(n9718), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n9652) );
  NAND2_X1 U11368 ( .A1(n9717), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n9651) );
  OAI211_X1 U11369 ( .C1(n9908), .C2(n9653), .A(n9652), .B(n9651), .ZN(n9654)
         );
  INV_X1 U11370 ( .A(n9654), .ZN(n9655) );
  NAND2_X1 U11371 ( .A1(n14227), .A2(n14360), .ZN(n9657) );
  XNOR2_X1 U11372 ( .A(n9659), .B(n9658), .ZN(n12377) );
  NAND2_X1 U11373 ( .A1(n12377), .A2(n9916), .ZN(n9661) );
  OR2_X1 U11374 ( .A1(n9917), .A2(n12724), .ZN(n9660) );
  INV_X1 U11375 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n9662) );
  NAND2_X1 U11376 ( .A1(n9663), .A2(n9662), .ZN(n9676) );
  OR2_X1 U11377 ( .A1(n9663), .A2(n9662), .ZN(n9664) );
  NAND2_X1 U11378 ( .A1(n9676), .A2(n9664), .ZN(n14206) );
  NAND2_X1 U11379 ( .A1(n14206), .A2(n9708), .ZN(n9670) );
  INV_X1 U11380 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n9667) );
  NAND2_X1 U11381 ( .A1(n9904), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n9666) );
  NAND2_X1 U11382 ( .A1(n9718), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n9665) );
  OAI211_X1 U11383 ( .C1(n9667), .C2(n9908), .A(n9666), .B(n9665), .ZN(n9668)
         );
  INV_X1 U11384 ( .A(n9668), .ZN(n9669) );
  XNOR2_X1 U11385 ( .A(n14361), .B(n14197), .ZN(n14204) );
  NAND2_X1 U11386 ( .A1(n14209), .A2(n14204), .ZN(n14212) );
  XNOR2_X1 U11387 ( .A(n9673), .B(n9672), .ZN(n12462) );
  NAND2_X1 U11388 ( .A1(n12462), .A2(n9916), .ZN(n9675) );
  INV_X1 U11389 ( .A(SI_26_), .ZN(n12464) );
  OR2_X1 U11390 ( .A1(n9917), .A2(n12464), .ZN(n9674) );
  NAND2_X1 U11391 ( .A1(n9676), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9677) );
  NAND2_X1 U11392 ( .A1(n9687), .A2(n9677), .ZN(n14195) );
  NAND2_X1 U11393 ( .A1(n14195), .A2(n9708), .ZN(n9683) );
  INV_X1 U11394 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n9680) );
  NAND2_X1 U11395 ( .A1(n9718), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n9679) );
  NAND2_X1 U11396 ( .A1(n9904), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n9678) );
  OAI211_X1 U11397 ( .C1(n9908), .C2(n9680), .A(n9679), .B(n9678), .ZN(n9681)
         );
  INV_X1 U11398 ( .A(n9681), .ZN(n9682) );
  NAND2_X1 U11399 ( .A1(n14356), .A2(n14186), .ZN(n9931) );
  XNOR2_X1 U11400 ( .A(n9685), .B(n9684), .ZN(n12528) );
  INV_X1 U11401 ( .A(n9700), .ZN(n9689) );
  NAND2_X1 U11402 ( .A1(n9687), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9688) );
  NAND2_X1 U11403 ( .A1(n9689), .A2(n9688), .ZN(n14184) );
  NAND2_X1 U11404 ( .A1(n14184), .A2(n9708), .ZN(n9695) );
  INV_X1 U11405 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n9692) );
  NAND2_X1 U11406 ( .A1(n9904), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n9691) );
  NAND2_X1 U11407 ( .A1(n9718), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n9690) );
  OAI211_X1 U11408 ( .C1(n9692), .C2(n9908), .A(n9691), .B(n9690), .ZN(n9693)
         );
  INV_X1 U11409 ( .A(n9693), .ZN(n9694) );
  NAND2_X1 U11410 ( .A1(n9860), .A2(n14346), .ZN(n9933) );
  XNOR2_X1 U11411 ( .A(n9697), .B(n9696), .ZN(n13247) );
  NAND2_X1 U11412 ( .A1(n13247), .A2(n9916), .ZN(n9699) );
  OR2_X1 U11413 ( .A1(n9917), .A2(n13249), .ZN(n9698) );
  INV_X1 U11414 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n9885) );
  NOR2_X1 U11415 ( .A1(n9700), .A2(n9885), .ZN(n9701) );
  INV_X1 U11416 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n9704) );
  NAND2_X1 U11417 ( .A1(n9904), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n9703) );
  NAND2_X1 U11418 ( .A1(n9718), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n9702) );
  OAI211_X1 U11419 ( .C1(n9704), .C2(n9908), .A(n9703), .B(n9702), .ZN(n9705)
         );
  OR2_X1 U11420 ( .A1(n14347), .A2(n14044), .ZN(n10048) );
  NAND2_X1 U11421 ( .A1(n14347), .A2(n14044), .ZN(n10047) );
  NAND2_X1 U11422 ( .A1(n14175), .A2(n14176), .ZN(n14179) );
  INV_X1 U11423 ( .A(n14347), .ZN(n9889) );
  NAND2_X1 U11424 ( .A1(n14164), .A2(n9708), .ZN(n9912) );
  INV_X1 U11425 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n9711) );
  NAND2_X1 U11426 ( .A1(n9718), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n9710) );
  NAND2_X1 U11427 ( .A1(n9904), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9709) );
  OAI211_X1 U11428 ( .C1(n9908), .C2(n9711), .A(n9710), .B(n9709), .ZN(n9712)
         );
  INV_X1 U11429 ( .A(n9712), .ZN(n9713) );
  NAND2_X1 U11430 ( .A1(n9912), .A2(n9713), .ZN(n14178) );
  NAND2_X1 U11431 ( .A1(n14166), .A2(n14178), .ZN(n10044) );
  INV_X1 U11432 ( .A(n14178), .ZN(n9881) );
  NAND2_X1 U11433 ( .A1(n9268), .A2(n9881), .ZN(n10046) );
  NAND2_X1 U11434 ( .A1(n10400), .A2(n9742), .ZN(n10080) );
  INV_X1 U11435 ( .A(n13248), .ZN(n10214) );
  NAND2_X1 U11436 ( .A1(n10214), .A2(n10164), .ZN(n10133) );
  NAND2_X1 U11437 ( .A1(n7594), .A2(n10133), .ZN(n9882) );
  AND2_X1 U11438 ( .A1(n10214), .A2(P3_B_REG_SCAN_IN), .ZN(n9716) );
  OR2_X1 U11439 ( .A1(n16056), .A2(n9716), .ZN(n14157) );
  INV_X1 U11440 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n9721) );
  NAND2_X1 U11441 ( .A1(n9904), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9720) );
  NAND2_X1 U11442 ( .A1(n9718), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n9719) );
  OAI211_X1 U11443 ( .C1(n9721), .C2(n9908), .A(n9720), .B(n9719), .ZN(n9722)
         );
  INV_X1 U11444 ( .A(n9722), .ZN(n9723) );
  NAND2_X1 U11445 ( .A1(n9726), .A2(n11243), .ZN(n11245) );
  NAND2_X1 U11446 ( .A1(n11245), .A2(n9946), .ZN(n16048) );
  NAND2_X1 U11447 ( .A1(n16048), .A2(n16050), .ZN(n9728) );
  OR2_X1 U11448 ( .A1(n14058), .A2(n16049), .ZN(n9727) );
  NAND2_X1 U11449 ( .A1(n9728), .A2(n9727), .ZN(n10397) );
  NAND2_X1 U11450 ( .A1(n10397), .A2(n10396), .ZN(n10399) );
  NAND2_X1 U11451 ( .A1(n10399), .A2(n9958), .ZN(n11579) );
  NAND2_X1 U11452 ( .A1(n11579), .A2(n11578), .ZN(n11581) );
  NAND2_X1 U11453 ( .A1(n11581), .A2(n9959), .ZN(n11802) );
  INV_X1 U11454 ( .A(n11804), .ZN(n11801) );
  NAND2_X1 U11455 ( .A1(n11802), .A2(n11801), .ZN(n11800) );
  NAND2_X1 U11456 ( .A1(n11800), .A2(n9963), .ZN(n11753) );
  NAND2_X1 U11457 ( .A1(n11753), .A2(n11754), .ZN(n11752) );
  INV_X1 U11458 ( .A(n16101), .ZN(n9784) );
  OR2_X1 U11459 ( .A1(n14056), .A2(n9784), .ZN(n9729) );
  NAND2_X1 U11460 ( .A1(n11752), .A2(n9729), .ZN(n11840) );
  NAND2_X1 U11461 ( .A1(n11840), .A2(n7939), .ZN(n11839) );
  NAND2_X1 U11462 ( .A1(n11839), .A2(n9970), .ZN(n11961) );
  NAND2_X1 U11463 ( .A1(n11961), .A2(n11960), .ZN(n11959) );
  OR2_X1 U11464 ( .A1(n14053), .A2(n12075), .ZN(n9730) );
  NAND2_X1 U11465 ( .A1(n14052), .A2(n12444), .ZN(n9977) );
  NAND2_X1 U11466 ( .A1(n12328), .A2(n9983), .ZN(n12499) );
  NAND2_X1 U11467 ( .A1(n12322), .A2(n12501), .ZN(n9992) );
  NAND2_X1 U11468 ( .A1(n12499), .A2(n12498), .ZN(n12497) );
  NAND2_X1 U11469 ( .A1(n12497), .A2(n9987), .ZN(n12596) );
  NAND2_X1 U11470 ( .A1(n16232), .A2(n14050), .ZN(n9993) );
  OR2_X1 U11471 ( .A1(n13235), .A2(n14049), .ZN(n9997) );
  NAND2_X1 U11472 ( .A1(n13235), .A2(n14049), .ZN(n9989) );
  NAND2_X1 U11473 ( .A1(n9997), .A2(n9989), .ZN(n10066) );
  INV_X1 U11474 ( .A(n13177), .ZN(n9732) );
  NOR2_X1 U11475 ( .A1(n10066), .A2(n9732), .ZN(n9733) );
  INV_X1 U11476 ( .A(n13188), .ZN(n9734) );
  INV_X1 U11477 ( .A(n13209), .ZN(n13213) );
  NAND2_X1 U11478 ( .A1(n14334), .A2(n14333), .ZN(n14332) );
  INV_X1 U11479 ( .A(n14046), .ZN(n14317) );
  NAND2_X1 U11480 ( .A1(n9944), .A2(n14317), .ZN(n9735) );
  NAND2_X1 U11481 ( .A1(n14332), .A2(n9735), .ZN(n14320) );
  NAND2_X1 U11482 ( .A1(n14320), .A2(n14319), .ZN(n14318) );
  NAND2_X1 U11483 ( .A1(n14318), .A2(n10019), .ZN(n14309) );
  INV_X1 U11484 ( .A(n14305), .ZN(n14390) );
  OR2_X1 U11485 ( .A1(n14397), .A2(n14390), .ZN(n9942) );
  NAND2_X1 U11486 ( .A1(n14397), .A2(n14390), .ZN(n9736) );
  INV_X1 U11487 ( .A(n9736), .ZN(n14274) );
  NOR2_X1 U11488 ( .A1(n7542), .A2(n14274), .ZN(n9737) );
  NAND2_X1 U11489 ( .A1(n14276), .A2(n10027), .ZN(n14270) );
  INV_X1 U11490 ( .A(n14045), .ZN(n14281) );
  NAND2_X1 U11491 ( .A1(n14385), .A2(n14281), .ZN(n10031) );
  NAND2_X1 U11492 ( .A1(n14227), .A2(n14208), .ZN(n9940) );
  INV_X1 U11493 ( .A(n9739), .ZN(n9936) );
  NAND2_X1 U11494 ( .A1(n14198), .A2(n9929), .ZN(n14189) );
  INV_X1 U11495 ( .A(n9932), .ZN(n9740) );
  AND2_X1 U11496 ( .A1(n16231), .A2(n10079), .ZN(n9741) );
  NAND2_X1 U11497 ( .A1(n9869), .A2(n9741), .ZN(n9744) );
  NAND2_X1 U11498 ( .A1(n9742), .A2(n14145), .ZN(n9743) );
  OR2_X1 U11499 ( .A1(n9755), .A2(n9743), .ZN(n9751) );
  AND2_X1 U11500 ( .A1(n9744), .A2(n9751), .ZN(n14256) );
  NAND2_X1 U11501 ( .A1(n9755), .A2(n16061), .ZN(n14365) );
  NAND2_X1 U11502 ( .A1(n9747), .A2(n9746), .ZN(P3_U3456) );
  XNOR2_X1 U11503 ( .A(n9767), .B(n14466), .ZN(n9750) );
  INV_X1 U11504 ( .A(n14466), .ZN(n9759) );
  NAND2_X1 U11505 ( .A1(n10129), .A2(n9752), .ZN(n9871) );
  NAND2_X1 U11506 ( .A1(n10043), .A2(n9751), .ZN(n10388) );
  AND2_X1 U11507 ( .A1(n9871), .A2(n10388), .ZN(n10390) );
  NAND2_X1 U11508 ( .A1(n9753), .A2(n9752), .ZN(n9756) );
  AOI22_X1 U11509 ( .A1(n9756), .A2(n11767), .B1(n9755), .B2(n9754), .ZN(n9757) );
  NAND2_X1 U11510 ( .A1(n9759), .A2(n9757), .ZN(n9758) );
  OAI21_X1 U11511 ( .B1(n9759), .B2(n10390), .A(n9758), .ZN(n9760) );
  INV_X1 U11512 ( .A(n9760), .ZN(n9761) );
  NAND2_X1 U11513 ( .A1(n9268), .A2(n12441), .ZN(n9763) );
  NAND2_X1 U11514 ( .A1(n9764), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n9762) );
  NAND2_X1 U11515 ( .A1(n9766), .A2(n9765), .ZN(P3_U3488) );
  OAI21_X1 U11516 ( .B1(n10400), .B2(n14145), .A(n11614), .ZN(n9768) );
  XNOR2_X1 U11517 ( .A(n9770), .B(n16040), .ZN(n11228) );
  NAND2_X1 U11518 ( .A1(n9801), .A2(n11481), .ZN(n9769) );
  AND2_X1 U11519 ( .A1(n9769), .A2(n11250), .ZN(n11229) );
  NAND2_X1 U11520 ( .A1(n9770), .A2(n7579), .ZN(n9771) );
  NAND2_X1 U11521 ( .A1(n11227), .A2(n9771), .ZN(n11329) );
  INV_X1 U11522 ( .A(n14058), .ZN(n11427) );
  NAND2_X1 U11523 ( .A1(n9773), .A2(n11427), .ZN(n9774) );
  INV_X2 U11524 ( .A(n9849), .ZN(n9857) );
  XNOR2_X1 U11525 ( .A(n9857), .B(n11522), .ZN(n9777) );
  XNOR2_X1 U11526 ( .A(n9777), .B(n14057), .ZN(n11412) );
  NAND2_X1 U11527 ( .A1(n9777), .A2(n14057), .ZN(n9778) );
  XNOR2_X1 U11528 ( .A(n9801), .B(n11727), .ZN(n9779) );
  XNOR2_X1 U11529 ( .A(n9779), .B(n11806), .ZN(n11724) );
  INV_X1 U11530 ( .A(n9779), .ZN(n9780) );
  INV_X1 U11531 ( .A(n11806), .ZN(n11834) );
  NAND2_X1 U11532 ( .A1(n9780), .A2(n11834), .ZN(n9781) );
  INV_X2 U11533 ( .A(n9849), .ZN(n9863) );
  XNOR2_X1 U11534 ( .A(n9863), .B(n16097), .ZN(n9782) );
  XNOR2_X1 U11535 ( .A(n9782), .B(n11575), .ZN(n11832) );
  INV_X1 U11536 ( .A(n11575), .ZN(n11946) );
  NAND2_X1 U11537 ( .A1(n9782), .A2(n11946), .ZN(n9783) );
  XNOR2_X1 U11538 ( .A(n9863), .B(n9784), .ZN(n9785) );
  XNOR2_X1 U11539 ( .A(n9785), .B(n14056), .ZN(n11942) );
  NAND2_X1 U11540 ( .A1(n9785), .A2(n14056), .ZN(n9786) );
  XNOR2_X1 U11541 ( .A(n9863), .B(n12053), .ZN(n9787) );
  XNOR2_X1 U11542 ( .A(n9787), .B(n14054), .ZN(n12048) );
  INV_X1 U11543 ( .A(n9787), .ZN(n9788) );
  NAND2_X1 U11544 ( .A1(n9788), .A2(n14054), .ZN(n9789) );
  XNOR2_X1 U11545 ( .A(n9863), .B(n12263), .ZN(n9790) );
  XNOR2_X1 U11546 ( .A(n9790), .B(n14053), .ZN(n12258) );
  INV_X1 U11547 ( .A(n9790), .ZN(n9791) );
  NAND2_X1 U11548 ( .A1(n9791), .A2(n14053), .ZN(n9792) );
  XNOR2_X1 U11549 ( .A(n9863), .B(n12444), .ZN(n9793) );
  XNOR2_X1 U11550 ( .A(n9793), .B(n14052), .ZN(n12401) );
  INV_X1 U11551 ( .A(n9793), .ZN(n9794) );
  INV_X1 U11552 ( .A(n14052), .ZN(n12332) );
  NAND2_X1 U11553 ( .A1(n9794), .A2(n12332), .ZN(n9795) );
  XNOR2_X1 U11554 ( .A(n9863), .B(n12473), .ZN(n9797) );
  XNOR2_X1 U11555 ( .A(n9797), .B(n14051), .ZN(n10255) );
  INV_X1 U11556 ( .A(n10255), .ZN(n9796) );
  NAND2_X1 U11557 ( .A1(n9797), .A2(n14051), .ZN(n9798) );
  AND2_X1 U11558 ( .A1(n9799), .A2(n9849), .ZN(n9804) );
  NAND2_X1 U11559 ( .A1(n9804), .A2(n9800), .ZN(n9803) );
  AND2_X1 U11560 ( .A1(n9992), .A2(n9801), .ZN(n9805) );
  NAND2_X1 U11561 ( .A1(n9805), .A2(n9987), .ZN(n9802) );
  NAND2_X1 U11562 ( .A1(n9803), .A2(n9802), .ZN(n12640) );
  INV_X1 U11563 ( .A(n9804), .ZN(n9807) );
  INV_X1 U11564 ( .A(n9805), .ZN(n9806) );
  NAND2_X1 U11565 ( .A1(n9807), .A2(n9806), .ZN(n9808) );
  XNOR2_X1 U11566 ( .A(n12600), .B(n9863), .ZN(n13196) );
  INV_X1 U11567 ( .A(n13196), .ZN(n9809) );
  NAND2_X1 U11568 ( .A1(n9809), .A2(n13230), .ZN(n9810) );
  OR2_X1 U11569 ( .A1(n10066), .A2(n9849), .ZN(n9814) );
  NAND2_X1 U11570 ( .A1(n9811), .A2(n9849), .ZN(n9816) );
  OR2_X1 U11571 ( .A1(n9816), .A2(n9812), .ZN(n9813) );
  AND2_X1 U11572 ( .A1(n9814), .A2(n9813), .ZN(n13225) );
  NAND2_X1 U11573 ( .A1(n9989), .A2(n9863), .ZN(n9815) );
  NAND2_X1 U11574 ( .A1(n9816), .A2(n9815), .ZN(n9817) );
  XNOR2_X1 U11575 ( .A(n14422), .B(n9863), .ZN(n9818) );
  XNOR2_X1 U11576 ( .A(n9818), .B(n13211), .ZN(n13935) );
  NAND2_X1 U11577 ( .A1(n13936), .A2(n13935), .ZN(n13934) );
  NAND2_X1 U11578 ( .A1(n9818), .A2(n14048), .ZN(n9819) );
  XNOR2_X1 U11579 ( .A(n14463), .B(n9849), .ZN(n14028) );
  NAND2_X1 U11580 ( .A1(n14028), .A2(n14331), .ZN(n9820) );
  NAND2_X1 U11581 ( .A1(n14030), .A2(n9820), .ZN(n9823) );
  INV_X1 U11582 ( .A(n14028), .ZN(n9821) );
  NAND2_X1 U11583 ( .A1(n9821), .A2(n14047), .ZN(n9822) );
  NAND2_X1 U11584 ( .A1(n9823), .A2(n9822), .ZN(n13974) );
  XNOR2_X1 U11585 ( .A(n9944), .B(n9863), .ZN(n9824) );
  XNOR2_X1 U11586 ( .A(n9824), .B(n14046), .ZN(n13973) );
  NAND2_X1 U11587 ( .A1(n13974), .A2(n13973), .ZN(n9827) );
  INV_X1 U11588 ( .A(n9824), .ZN(n9825) );
  NAND2_X1 U11589 ( .A1(n9825), .A2(n14046), .ZN(n9826) );
  XNOR2_X1 U11590 ( .A(n14455), .B(n9863), .ZN(n9828) );
  XNOR2_X1 U11591 ( .A(n9828), .B(n14330), .ZN(n13981) );
  NAND2_X1 U11592 ( .A1(n13982), .A2(n13981), .ZN(n9830) );
  NAND2_X1 U11593 ( .A1(n9828), .A2(n14306), .ZN(n9829) );
  XNOR2_X1 U11594 ( .A(n14016), .B(n9857), .ZN(n9831) );
  XNOR2_X1 U11595 ( .A(n9831), .B(n14290), .ZN(n14012) );
  NAND2_X1 U11596 ( .A1(n14013), .A2(n14012), .ZN(n9834) );
  INV_X1 U11597 ( .A(n9831), .ZN(n9832) );
  NAND2_X1 U11598 ( .A1(n9832), .A2(n14290), .ZN(n9833) );
  NAND2_X1 U11599 ( .A1(n9834), .A2(n9833), .ZN(n13950) );
  XNOR2_X1 U11600 ( .A(n14397), .B(n9857), .ZN(n9835) );
  XNOR2_X1 U11601 ( .A(n9835), .B(n14305), .ZN(n13949) );
  NAND2_X1 U11602 ( .A1(n13950), .A2(n13949), .ZN(n9838) );
  INV_X1 U11603 ( .A(n9835), .ZN(n9836) );
  NAND2_X1 U11604 ( .A1(n9836), .A2(n14305), .ZN(n9837) );
  XNOR2_X1 U11605 ( .A(n14389), .B(n9857), .ZN(n9839) );
  XNOR2_X1 U11606 ( .A(n9839), .B(n14383), .ZN(n13999) );
  INV_X1 U11607 ( .A(n9839), .ZN(n9840) );
  NAND2_X1 U11608 ( .A1(n9840), .A2(n14383), .ZN(n9841) );
  INV_X1 U11609 ( .A(n10030), .ZN(n9842) );
  MUX2_X1 U11610 ( .A(n9843), .B(n9842), .S(n9863), .Z(n13958) );
  XNOR2_X1 U11611 ( .A(n14385), .B(n9857), .ZN(n9844) );
  NAND2_X1 U11612 ( .A1(n9844), .A2(n14281), .ZN(n13956) );
  XNOR2_X1 U11613 ( .A(n14377), .B(n9849), .ZN(n9845) );
  XNOR2_X1 U11614 ( .A(n9847), .B(n9845), .ZN(n14006) );
  INV_X1 U11615 ( .A(n9845), .ZN(n9846) );
  AND2_X1 U11616 ( .A1(n9847), .A2(n9846), .ZN(n9848) );
  XNOR2_X1 U11617 ( .A(n14227), .B(n9857), .ZN(n13991) );
  XNOR2_X1 U11618 ( .A(n14372), .B(n9849), .ZN(n13988) );
  INV_X1 U11619 ( .A(n13988), .ZN(n9850) );
  OAI22_X1 U11620 ( .A1(n13991), .A2(n14208), .B1(n14252), .B2(n9850), .ZN(
        n9854) );
  OAI21_X1 U11621 ( .B1(n13988), .B2(n14223), .A(n14360), .ZN(n9852) );
  NOR2_X1 U11622 ( .A1(n14360), .A2(n14223), .ZN(n9851) );
  AOI22_X1 U11623 ( .A1(n13991), .A2(n9852), .B1(n9851), .B2(n9850), .ZN(n9853) );
  XNOR2_X1 U11624 ( .A(n8347), .B(n9857), .ZN(n9855) );
  XNOR2_X1 U11625 ( .A(n9855), .B(n14197), .ZN(n13967) );
  INV_X1 U11626 ( .A(n9855), .ZN(n9856) );
  XNOR2_X1 U11627 ( .A(n14356), .B(n9857), .ZN(n9858) );
  INV_X1 U11628 ( .A(n9858), .ZN(n9859) );
  XNOR2_X1 U11629 ( .A(n9860), .B(n9863), .ZN(n9861) );
  XNOR2_X1 U11630 ( .A(n9861), .B(n14174), .ZN(n13928) );
  INV_X1 U11631 ( .A(n9861), .ZN(n9862) );
  NAND2_X1 U11632 ( .A1(n9869), .A2(n16231), .ZN(n9865) );
  INV_X1 U11633 ( .A(n9872), .ZN(n9864) );
  OAI22_X1 U11634 ( .A1(n9870), .A2(n9865), .B1(n9880), .B2(n9864), .ZN(n9866)
         );
  NAND2_X1 U11635 ( .A1(n9870), .A2(n11435), .ZN(n9868) );
  AND2_X1 U11636 ( .A1(n10395), .A2(n16102), .ZN(n9867) );
  NAND2_X1 U11637 ( .A1(n9870), .A2(n9869), .ZN(n9875) );
  AND3_X1 U11638 ( .A1(n9871), .A2(n10105), .A3(n10128), .ZN(n9874) );
  NAND2_X1 U11639 ( .A1(n9880), .A2(n9872), .ZN(n9873) );
  NAND3_X1 U11640 ( .A1(n9875), .A2(n9874), .A3(n9873), .ZN(n9876) );
  NAND2_X1 U11641 ( .A1(n9876), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9879) );
  INV_X1 U11642 ( .A(n10082), .ZN(n9877) );
  NAND2_X1 U11643 ( .A1(n9880), .A2(n9877), .ZN(n9878) );
  NOR2_X1 U11644 ( .A1(n9880), .A2(n10082), .ZN(n9884) );
  NAND2_X1 U11645 ( .A1(n9884), .A2(n9882), .ZN(n14032) );
  NOR2_X1 U11646 ( .A1(n9881), .A2(n14032), .ZN(n9887) );
  INV_X1 U11647 ( .A(n9882), .ZN(n9883) );
  OAI22_X1 U11648 ( .A1(n14174), .A2(n14015), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n9885), .ZN(n9886) );
  AOI211_X1 U11649 ( .C1(n14172), .C2(n14023), .A(n9887), .B(n9886), .ZN(n9888) );
  OAI21_X1 U11650 ( .B1(n9889), .B2(n14017), .A(n9888), .ZN(n9890) );
  NAND2_X1 U11651 ( .A1(n9892), .A2(n9891), .ZN(P3_U3160) );
  INV_X4 U11652 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U11653 ( .A(n9893), .ZN(n9894) );
  NAND2_X1 U11654 ( .A1(n15593), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n9896) );
  NAND2_X1 U11655 ( .A1(n9897), .A2(n9896), .ZN(n9915) );
  XNOR2_X1 U11656 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .ZN(n9913) );
  NAND2_X1 U11657 ( .A1(n9915), .A2(n9913), .ZN(n9899) );
  NAND2_X1 U11658 ( .A1(n13604), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n9898) );
  NAND2_X1 U11659 ( .A1(n9899), .A2(n9898), .ZN(n9901) );
  INV_X1 U11660 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n13606) );
  XNOR2_X1 U11661 ( .A(n13606), .B(P2_DATAO_REG_31__SCAN_IN), .ZN(n9900) );
  XNOR2_X1 U11662 ( .A(n9901), .B(n9900), .ZN(n14475) );
  NAND2_X1 U11663 ( .A1(n14475), .A2(n9916), .ZN(n9903) );
  INV_X1 U11664 ( .A(SI_31_), .ZN(n14471) );
  OR2_X1 U11665 ( .A1(n9917), .A2(n14471), .ZN(n9902) );
  NAND2_X1 U11666 ( .A1(n9903), .A2(n9902), .ZN(n14156) );
  INV_X1 U11667 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n9909) );
  NAND2_X1 U11668 ( .A1(n9904), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n9907) );
  INV_X1 U11669 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n9905) );
  OR2_X1 U11670 ( .A1(n9293), .A2(n9905), .ZN(n9906) );
  OAI211_X1 U11671 ( .C1(n9909), .C2(n9908), .A(n9907), .B(n9906), .ZN(n9910)
         );
  INV_X1 U11672 ( .A(n9910), .ZN(n9911) );
  OR2_X1 U11673 ( .A1(n14156), .A2(n14158), .ZN(n9921) );
  INV_X1 U11674 ( .A(n9913), .ZN(n9914) );
  XNOR2_X1 U11675 ( .A(n9915), .B(n9914), .ZN(n13326) );
  NAND2_X1 U11676 ( .A1(n13326), .A2(n9916), .ZN(n9919) );
  INV_X1 U11677 ( .A(SI_30_), .ZN(n13328) );
  OR2_X1 U11678 ( .A1(n9917), .A2(n13328), .ZN(n9918) );
  NAND2_X1 U11679 ( .A1(n9919), .A2(n9918), .ZN(n9924) );
  NAND2_X1 U11680 ( .A1(n9924), .A2(n11792), .ZN(n9920) );
  NAND2_X1 U11681 ( .A1(n9921), .A2(n9920), .ZN(n10053) );
  INV_X1 U11682 ( .A(n14158), .ZN(n14043) );
  OAI21_X1 U11683 ( .B1(n14428), .B2(n14043), .A(n10046), .ZN(n9922) );
  AOI211_X1 U11684 ( .C1(n9923), .C2(n10044), .A(n10053), .B(n9922), .ZN(n9926) );
  AND2_X1 U11685 ( .A1(n14156), .A2(n14158), .ZN(n10073) );
  NOR2_X1 U11686 ( .A1(n9924), .A2(n11792), .ZN(n10072) );
  NOR2_X1 U11687 ( .A1(n9926), .A2(n9925), .ZN(n9928) );
  XNOR2_X1 U11688 ( .A(n9928), .B(n9927), .ZN(n10081) );
  NAND3_X1 U11689 ( .A1(n9929), .A2(n14197), .A3(n14361), .ZN(n9930) );
  NAND3_X1 U11690 ( .A1(n9932), .A2(n9931), .A3(n9930), .ZN(n9934) );
  AND2_X1 U11691 ( .A1(n9934), .A2(n9933), .ZN(n9939) );
  INV_X1 U11692 ( .A(n14204), .ZN(n14210) );
  NAND3_X1 U11693 ( .A1(n9935), .A2(n14199), .A3(n14210), .ZN(n9937) );
  NOR2_X1 U11694 ( .A1(n9937), .A2(n9940), .ZN(n9938) );
  NOR2_X1 U11695 ( .A1(n9937), .A2(n9936), .ZN(n9941) );
  OAI211_X1 U11696 ( .C1(n7697), .C2(n9943), .A(n9942), .B(n10022), .ZN(n10018) );
  INV_X1 U11697 ( .A(n9944), .ZN(n14459) );
  MUX2_X1 U11698 ( .A(n14317), .B(n14459), .S(n10043), .Z(n10009) );
  INV_X1 U11699 ( .A(n10009), .ZN(n10013) );
  MUX2_X1 U11700 ( .A(n10043), .B(n14056), .S(n16101), .Z(n9969) );
  NOR2_X1 U11701 ( .A1(n14056), .A2(n10043), .ZN(n9968) );
  NAND2_X1 U11702 ( .A1(n14059), .A2(n11481), .ZN(n10055) );
  NAND2_X1 U11703 ( .A1(n9945), .A2(n10055), .ZN(n9947) );
  NAND3_X1 U11704 ( .A1(n16050), .A2(n9946), .A3(n9947), .ZN(n9952) );
  INV_X1 U11705 ( .A(n9958), .ZN(n9950) );
  NOR3_X1 U11706 ( .A1(n9948), .A2(n9947), .A3(n11767), .ZN(n9949) );
  NOR3_X1 U11707 ( .A1(n10397), .A2(n9950), .A3(n9949), .ZN(n9951) );
  MUX2_X1 U11708 ( .A(n9952), .B(n9951), .S(n10043), .Z(n9956) );
  INV_X1 U11709 ( .A(n9953), .ZN(n9955) );
  AOI21_X1 U11710 ( .B1(n14058), .B2(n16049), .A(n9955), .ZN(n9954) );
  OAI22_X1 U11711 ( .A1(n9956), .A2(n9955), .B1(n9954), .B2(n10043), .ZN(n9957) );
  OAI211_X1 U11712 ( .C1(n9958), .C2(n10043), .A(n9957), .B(n11578), .ZN(n9962) );
  MUX2_X1 U11713 ( .A(n9960), .B(n9959), .S(n10043), .Z(n9961) );
  NAND3_X1 U11714 ( .A1(n9962), .A2(n11801), .A3(n9961), .ZN(n9966) );
  MUX2_X1 U11715 ( .A(n9964), .B(n9963), .S(n10129), .Z(n9965) );
  NAND3_X1 U11716 ( .A1(n9966), .A2(n11754), .A3(n9965), .ZN(n9967) );
  OAI211_X1 U11717 ( .C1(n9969), .C2(n9968), .A(n9967), .B(n7939), .ZN(n9973)
         );
  MUX2_X1 U11718 ( .A(n9971), .B(n9970), .S(n10129), .Z(n9972) );
  NAND3_X1 U11719 ( .A1(n9973), .A2(n11960), .A3(n9972), .ZN(n9982) );
  NOR2_X1 U11720 ( .A1(n12075), .A2(n10129), .ZN(n9975) );
  NOR2_X1 U11721 ( .A1(n12263), .A2(n10043), .ZN(n9974) );
  MUX2_X1 U11722 ( .A(n9975), .B(n9974), .S(n14053), .Z(n9976) );
  NOR2_X1 U11723 ( .A1(n9420), .A2(n9976), .ZN(n9981) );
  NOR2_X1 U11724 ( .A1(n14052), .A2(n12444), .ZN(n9979) );
  INV_X1 U11725 ( .A(n9977), .ZN(n9978) );
  MUX2_X1 U11726 ( .A(n9979), .B(n9978), .S(n10043), .Z(n9980) );
  AOI21_X1 U11727 ( .B1(n9982), .B2(n9981), .A(n9980), .ZN(n9986) );
  MUX2_X1 U11728 ( .A(n9984), .B(n9983), .S(n10129), .Z(n9985) );
  OAI211_X1 U11729 ( .C1(n9986), .C2(n12325), .A(n12498), .B(n9985), .ZN(n9994) );
  NAND3_X1 U11730 ( .A1(n9994), .A2(n13177), .A3(n9987), .ZN(n9988) );
  NAND3_X1 U11731 ( .A1(n9988), .A2(n9993), .A3(n10043), .ZN(n9991) );
  INV_X1 U11732 ( .A(n10066), .ZN(n13176) );
  INV_X1 U11733 ( .A(n9989), .ZN(n9990) );
  AOI22_X1 U11734 ( .A1(n9991), .A2(n13176), .B1(n9990), .B2(n10043), .ZN(
        n10005) );
  NAND3_X1 U11735 ( .A1(n9994), .A2(n9993), .A3(n9992), .ZN(n9995) );
  NAND3_X1 U11736 ( .A1(n9995), .A2(n10129), .A3(n13177), .ZN(n9996) );
  NAND2_X1 U11737 ( .A1(n9996), .A2(n9734), .ZN(n10004) );
  INV_X1 U11738 ( .A(n9997), .ZN(n10000) );
  INV_X1 U11739 ( .A(n9998), .ZN(n9999) );
  AOI21_X1 U11740 ( .B1(n10000), .B2(n10002), .A(n9999), .ZN(n10001) );
  MUX2_X1 U11741 ( .A(n10002), .B(n10001), .S(n10129), .Z(n10003) );
  OAI211_X1 U11742 ( .C1(n10005), .C2(n10004), .A(n13213), .B(n10003), .ZN(
        n10011) );
  MUX2_X1 U11743 ( .A(n10007), .B(n10006), .S(n10043), .Z(n10010) );
  AOI22_X1 U11744 ( .A1(n10011), .A2(n10010), .B1(n10009), .B2(n10008), .ZN(
        n10012) );
  AOI21_X1 U11745 ( .B1(n10014), .B2(n10013), .A(n10012), .ZN(n10016) );
  INV_X1 U11746 ( .A(n14319), .ZN(n10015) );
  NOR3_X1 U11747 ( .A1(n10016), .A2(n14302), .A3(n10015), .ZN(n10017) );
  AOI21_X1 U11748 ( .B1(n10129), .B2(n10018), .A(n10017), .ZN(n10024) );
  NAND2_X1 U11749 ( .A1(n10020), .A2(n10019), .ZN(n10021) );
  AOI21_X1 U11750 ( .B1(n10022), .B2(n10021), .A(n14274), .ZN(n10023) );
  OAI22_X1 U11751 ( .A1(n10024), .A2(n14274), .B1(n10129), .B2(n10023), .ZN(
        n10026) );
  INV_X1 U11752 ( .A(n14397), .ZN(n14297) );
  NAND3_X1 U11753 ( .A1(n14297), .A2(n14305), .A3(n10043), .ZN(n10025) );
  AOI21_X1 U11754 ( .B1(n10026), .B2(n10025), .A(n7542), .ZN(n10034) );
  MUX2_X1 U11755 ( .A(n10028), .B(n10027), .S(n10043), .Z(n10029) );
  NAND2_X1 U11756 ( .A1(n14269), .A2(n10029), .ZN(n10033) );
  MUX2_X1 U11757 ( .A(n10031), .B(n10030), .S(n10129), .Z(n10032) );
  OAI211_X1 U11758 ( .C1(n10034), .C2(n10033), .A(n7950), .B(n10032), .ZN(
        n10038) );
  MUX2_X1 U11759 ( .A(n10036), .B(n10035), .S(n10043), .Z(n10037) );
  NAND3_X1 U11760 ( .A1(n10038), .A2(n14236), .A3(n10037), .ZN(n10042) );
  MUX2_X1 U11761 ( .A(n10040), .B(n10039), .S(n10129), .Z(n10041) );
  NAND2_X1 U11762 ( .A1(n10044), .A2(n10043), .ZN(n10045) );
  AOI22_X1 U11763 ( .A1(n10049), .A2(n10047), .B1(n10046), .B2(n10045), .ZN(
        n10052) );
  AND3_X1 U11764 ( .A1(n10049), .A2(n10129), .A3(n10048), .ZN(n10051) );
  INV_X1 U11765 ( .A(n10072), .ZN(n10050) );
  OAI21_X1 U11766 ( .B1(n10052), .B2(n10051), .A(n10050), .ZN(n10054) );
  INV_X1 U11767 ( .A(n10053), .ZN(n10076) );
  INV_X1 U11768 ( .A(n14269), .ZN(n10070) );
  AND2_X1 U11769 ( .A1(n7939), .A2(n10396), .ZN(n10060) );
  INV_X1 U11770 ( .A(n10055), .ZN(n10056) );
  OR2_X1 U11771 ( .A1(n11243), .A2(n10056), .ZN(n16042) );
  NOR2_X1 U11772 ( .A1(n16042), .A2(n11251), .ZN(n10059) );
  NOR2_X1 U11773 ( .A1(n11574), .A2(n11804), .ZN(n10058) );
  NAND4_X1 U11774 ( .A1(n10060), .A2(n10059), .A3(n9731), .A4(n10058), .ZN(
        n10062) );
  NAND3_X1 U11775 ( .A1(n16050), .A2(n11960), .A3(n11754), .ZN(n10061) );
  NOR2_X1 U11776 ( .A1(n10062), .A2(n10061), .ZN(n10064) );
  NAND4_X1 U11777 ( .A1(n10064), .A2(n12600), .A3(n10063), .A4(n12498), .ZN(
        n10065) );
  NOR2_X1 U11778 ( .A1(n10066), .A2(n10065), .ZN(n10067) );
  AND4_X1 U11779 ( .A1(n14333), .A2(n9734), .A3(n13213), .A4(n10067), .ZN(
        n10068) );
  NAND4_X1 U11780 ( .A1(n14293), .A2(n14319), .A3(n9576), .A4(n10068), .ZN(
        n10069) );
  OR4_X1 U11781 ( .A1(n14250), .A2(n7542), .A3(n10070), .A4(n10069), .ZN(
        n10071) );
  NOR4_X1 U11782 ( .A1(n10072), .A2(n14232), .A3(n14176), .A4(n10071), .ZN(
        n10075) );
  INV_X1 U11783 ( .A(n10073), .ZN(n10074) );
  NAND4_X1 U11784 ( .A1(n7480), .A2(n10076), .A3(n10075), .A4(n10074), .ZN(
        n10077) );
  OR2_X1 U11785 ( .A1(n10128), .A2(P3_U3151), .ZN(n11953) );
  INV_X1 U11786 ( .A(n11953), .ZN(n10127) );
  NOR3_X1 U11787 ( .A1(n10082), .A2(n10164), .A3(n13248), .ZN(n10084) );
  OAI21_X1 U11788 ( .B1(n11953), .B2(n11797), .A(P3_B_REG_SCAN_IN), .ZN(n10083) );
  OR2_X1 U11789 ( .A1(n10084), .A2(n10083), .ZN(n10085) );
  NAND2_X1 U11790 ( .A1(n10409), .A2(n10089), .ZN(n10090) );
  NAND4_X1 U11791 ( .A1(n10092), .A2(n10091), .A3(n10414), .A4(n10646), .ZN(
        n10719) );
  NOR2_X2 U11792 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n10648) );
  NOR2_X2 U11793 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n10649) );
  NAND2_X1 U11794 ( .A1(n10648), .A2(n10649), .ZN(n10720) );
  NOR2_X2 U11795 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n10294) );
  NAND2_X1 U11796 ( .A1(n10277), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10096) );
  NAND2_X1 U11797 ( .A1(n10098), .A2(n10097), .ZN(n10099) );
  NAND2_X1 U11798 ( .A1(n10102), .A2(n10263), .ZN(n10100) );
  NAND3_X1 U11799 ( .A1(n10352), .A2(n15066), .A3(n15071), .ZN(n10366) );
  INV_X1 U11800 ( .A(n10366), .ZN(n10103) );
  INV_X1 U11801 ( .A(n10105), .ZN(n10106) );
  AND2_X1 U11802 ( .A1(n12131), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n10208) );
  INV_X1 U11803 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n16067) );
  MUX2_X1 U11804 ( .A(n16067), .B(P3_REG2_REG_2__SCAN_IN), .S(n10170), .Z(
        n10824) );
  INV_X1 U11805 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10137) );
  AND2_X1 U11806 ( .A1(P3_REG2_REG_0__SCAN_IN), .A2(n10137), .ZN(n10107) );
  NAND2_X1 U11807 ( .A1(n10140), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10108) );
  OAI21_X1 U11808 ( .B1(n10475), .B2(n10107), .A(n10108), .ZN(n11090) );
  NAND2_X1 U11809 ( .A1(n11092), .A2(n10108), .ZN(n10823) );
  NAND2_X1 U11810 ( .A1(n10824), .A2(n10823), .ZN(n10822) );
  NAND2_X1 U11811 ( .A1(n10842), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10109) );
  NAND2_X1 U11812 ( .A1(n10822), .A2(n10109), .ZN(n10110) );
  INV_X1 U11813 ( .A(n11171), .ZN(n10441) );
  NAND2_X1 U11814 ( .A1(n11153), .A2(n10851), .ZN(n10111) );
  XNOR2_X1 U11815 ( .A(n10183), .B(P3_REG2_REG_4__SCAN_IN), .ZN(n10850) );
  INV_X1 U11816 ( .A(n10183), .ZN(n10867) );
  NAND2_X1 U11817 ( .A1(n10867), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n10112) );
  XNOR2_X1 U11818 ( .A(n15984), .B(P3_REG2_REG_6__SCAN_IN), .ZN(n15971) );
  NOR2_X1 U11819 ( .A1(n10466), .A2(n10113), .ZN(n10114) );
  MUX2_X1 U11820 ( .A(P3_REG2_REG_8__SCAN_IN), .B(n10115), .S(n10479), .Z(
        n11374) );
  OR2_X1 U11821 ( .A1(n10479), .A2(n10115), .ZN(n10116) );
  NAND2_X1 U11822 ( .A1(n10471), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n10118) );
  OAI21_X1 U11823 ( .B1(n10471), .B2(P3_REG2_REG_10__SCAN_IN), .A(n10118), 
        .ZN(n11617) );
  NAND2_X1 U11824 ( .A1(n11615), .A2(n10118), .ZN(n10120) );
  INV_X1 U11825 ( .A(n10120), .ZN(n10119) );
  NOR2_X1 U11826 ( .A1(n10155), .A2(n10119), .ZN(n10121) );
  XNOR2_X1 U11827 ( .A(n10120), .B(n12153), .ZN(n12148) );
  NOR2_X1 U11828 ( .A1(n12131), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n10122) );
  OR2_X1 U11829 ( .A1(n10208), .A2(n10122), .ZN(n12141) );
  NOR2_X1 U11830 ( .A1(n10210), .A2(n10123), .ZN(n10124) );
  NAND2_X1 U11831 ( .A1(n10729), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n10224) );
  OAI21_X1 U11832 ( .B1(n10729), .B2(P3_REG2_REG_14__SCAN_IN), .A(n10224), 
        .ZN(n10125) );
  NAND2_X1 U11833 ( .A1(n10126), .A2(n10125), .ZN(n10135) );
  NAND2_X1 U11834 ( .A1(n10129), .A2(n10128), .ZN(n10130) );
  NAND2_X1 U11835 ( .A1(n7594), .A2(n10130), .ZN(n10216) );
  INV_X1 U11836 ( .A(n10216), .ZN(n10132) );
  NAND2_X1 U11837 ( .A1(n10217), .A2(n10132), .ZN(n10215) );
  INV_X1 U11838 ( .A(n10215), .ZN(n10162) );
  INV_X1 U11839 ( .A(n10133), .ZN(n10134) );
  AOI21_X1 U11840 ( .B1(n10225), .B2(n10135), .A(n16009), .ZN(n10223) );
  NAND2_X1 U11841 ( .A1(n10140), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n10136) );
  NAND2_X1 U11842 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n10137), .ZN(n10138) );
  OR2_X1 U11843 ( .A1(n10138), .A2(n10140), .ZN(n10139) );
  AND2_X1 U11844 ( .A1(n10140), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n10141) );
  AOI21_X1 U11845 ( .B1(n11088), .B2(P3_REG1_REG_1__SCAN_IN), .A(n10141), .ZN(
        n10829) );
  NAND2_X1 U11846 ( .A1(n10842), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10826) );
  NAND2_X1 U11847 ( .A1(n10829), .A2(n10826), .ZN(n10143) );
  NAND2_X1 U11848 ( .A1(n10170), .A2(n10169), .ZN(n10142) );
  OR2_X1 U11849 ( .A1(n10825), .A2(n11171), .ZN(n10856) );
  NAND2_X1 U11850 ( .A1(n10825), .A2(n11171), .ZN(n10144) );
  XNOR2_X1 U11851 ( .A(n10183), .B(P3_REG1_REG_4__SCAN_IN), .ZN(n10855) );
  NAND2_X1 U11852 ( .A1(n10867), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n10145) );
  NAND2_X1 U11853 ( .A1(n10859), .A2(n10145), .ZN(n10146) );
  NAND2_X1 U11854 ( .A1(n10146), .A2(n11024), .ZN(n15976) );
  OAI21_X1 U11855 ( .B1(n10146), .B2(n11024), .A(n15976), .ZN(n11025) );
  XNOR2_X1 U11856 ( .A(n15984), .B(P3_REG1_REG_6__SCAN_IN), .ZN(n15977) );
  AOI21_X1 U11857 ( .B1(n15978), .B2(n15976), .A(n15977), .ZN(n15981) );
  AOI21_X1 U11858 ( .B1(P3_REG1_REG_6__SCAN_IN), .B2(n15984), .A(n15981), .ZN(
        n10147) );
  NOR2_X1 U11859 ( .A1(n10466), .A2(n10147), .ZN(n10148) );
  XNOR2_X1 U11860 ( .A(n10466), .B(n10147), .ZN(n15996) );
  MUX2_X1 U11861 ( .A(P3_REG1_REG_8__SCAN_IN), .B(n10149), .S(n10479), .Z(
        n11379) );
  OR2_X1 U11862 ( .A1(n10479), .A2(n10149), .ZN(n10150) );
  NOR2_X1 U11863 ( .A1(n16019), .A2(n10151), .ZN(n10152) );
  NAND2_X1 U11864 ( .A1(n10471), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n10153) );
  OAI21_X1 U11865 ( .B1(n10471), .B2(P3_REG1_REG_10__SCAN_IN), .A(n10153), 
        .ZN(n11620) );
  NOR2_X1 U11866 ( .A1(n10155), .A2(n10154), .ZN(n10156) );
  XNOR2_X1 U11867 ( .A(n10155), .B(n10154), .ZN(n12155) );
  INV_X1 U11868 ( .A(n10207), .ZN(n10157) );
  OAI21_X1 U11869 ( .B1(P3_REG1_REG_12__SCAN_IN), .B2(n12131), .A(n10157), 
        .ZN(n12129) );
  NOR2_X1 U11870 ( .A1(n10210), .A2(n10158), .ZN(n10159) );
  NOR2_X1 U11871 ( .A1(n10159), .A2(n14060), .ZN(n10161) );
  NAND2_X1 U11872 ( .A1(n10729), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n10234) );
  OAI21_X1 U11873 ( .B1(n10729), .B2(P3_REG1_REG_14__SCAN_IN), .A(n10234), 
        .ZN(n10160) );
  OR2_X1 U11874 ( .A1(n10161), .A2(n10160), .ZN(n10235) );
  NAND2_X1 U11875 ( .A1(n10161), .A2(n10160), .ZN(n10163) );
  AOI21_X1 U11876 ( .B1(n10235), .B2(n10163), .A(n16013), .ZN(n10222) );
  INV_X2 U11877 ( .A(n10164), .ZN(n10205) );
  MUX2_X1 U11878 ( .A(P3_REG2_REG_14__SCAN_IN), .B(P3_REG1_REG_14__SCAN_IN), 
        .S(n10205), .Z(n10242) );
  XNOR2_X1 U11879 ( .A(n10242), .B(n10729), .ZN(n10213) );
  MUX2_X1 U11880 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n14141), .Z(n10211) );
  MUX2_X1 U11881 ( .A(n11438), .B(n11256), .S(n9715), .Z(n10165) );
  NAND2_X1 U11882 ( .A1(n10165), .A2(n11096), .ZN(n10835) );
  INV_X1 U11883 ( .A(n10165), .ZN(n10166) );
  NAND2_X1 U11884 ( .A1(n10166), .A2(n10475), .ZN(n10167) );
  NAND2_X1 U11885 ( .A1(n10835), .A2(n10167), .ZN(n11087) );
  MUX2_X1 U11886 ( .A(n11477), .B(n10168), .S(n10205), .Z(n15962) );
  NAND2_X1 U11887 ( .A1(n15962), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n15961) );
  NAND2_X1 U11888 ( .A1(n10834), .A2(n10835), .ZN(n10174) );
  MUX2_X1 U11889 ( .A(n16067), .B(n10169), .S(n10205), .Z(n10171) );
  NAND2_X1 U11890 ( .A1(n10171), .A2(n10170), .ZN(n11165) );
  INV_X1 U11891 ( .A(n10171), .ZN(n10172) );
  NAND2_X1 U11892 ( .A1(n10172), .A2(n10842), .ZN(n10173) );
  AND2_X1 U11893 ( .A1(n11165), .A2(n10173), .ZN(n10836) );
  NAND2_X1 U11894 ( .A1(n10174), .A2(n10836), .ZN(n11166) );
  NAND2_X1 U11895 ( .A1(n11166), .A2(n11165), .ZN(n10180) );
  MUX2_X1 U11896 ( .A(n10176), .B(n10175), .S(n10205), .Z(n10177) );
  NAND2_X1 U11897 ( .A1(n10177), .A2(n11171), .ZN(n10843) );
  INV_X1 U11898 ( .A(n10177), .ZN(n10178) );
  NAND2_X1 U11899 ( .A1(n10178), .A2(n10441), .ZN(n10179) );
  AND2_X1 U11900 ( .A1(n10843), .A2(n10179), .ZN(n11163) );
  NAND2_X1 U11901 ( .A1(n10180), .A2(n11163), .ZN(n11168) );
  NAND2_X1 U11902 ( .A1(n11168), .A2(n10843), .ZN(n10181) );
  MUX2_X1 U11903 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n10205), .Z(n10182) );
  XNOR2_X1 U11904 ( .A(n10182), .B(n10183), .ZN(n10844) );
  NAND2_X1 U11905 ( .A1(n10181), .A2(n10844), .ZN(n10847) );
  INV_X1 U11906 ( .A(n10182), .ZN(n10184) );
  NAND2_X1 U11907 ( .A1(n10184), .A2(n10183), .ZN(n10185) );
  NAND2_X1 U11908 ( .A1(n10847), .A2(n10185), .ZN(n11022) );
  MUX2_X1 U11909 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n10205), .Z(n10186) );
  NAND2_X1 U11910 ( .A1(n10186), .A2(n11024), .ZN(n11021) );
  NAND2_X1 U11911 ( .A1(n11022), .A2(n11021), .ZN(n10189) );
  INV_X1 U11912 ( .A(n10186), .ZN(n10188) );
  NAND2_X1 U11913 ( .A1(n10188), .A2(n10187), .ZN(n11020) );
  NAND2_X1 U11914 ( .A1(n10189), .A2(n11020), .ZN(n15969) );
  MUX2_X1 U11915 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n10205), .Z(n10190) );
  INV_X1 U11916 ( .A(n15984), .ZN(n10191) );
  XNOR2_X1 U11917 ( .A(n10190), .B(n10191), .ZN(n15968) );
  NAND2_X1 U11918 ( .A1(n15969), .A2(n15968), .ZN(n10194) );
  INV_X1 U11919 ( .A(n10190), .ZN(n10192) );
  NAND2_X1 U11920 ( .A1(n10192), .A2(n10191), .ZN(n10193) );
  NAND2_X1 U11921 ( .A1(n10194), .A2(n10193), .ZN(n15991) );
  MUX2_X1 U11922 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n10205), .Z(n10195) );
  XNOR2_X1 U11923 ( .A(n10195), .B(n10466), .ZN(n15990) );
  NAND2_X1 U11924 ( .A1(n15991), .A2(n15990), .ZN(n10198) );
  INV_X1 U11925 ( .A(n10195), .ZN(n10196) );
  NAND2_X1 U11926 ( .A1(n10196), .A2(n10466), .ZN(n10197) );
  NAND2_X1 U11927 ( .A1(n10198), .A2(n10197), .ZN(n11372) );
  MUX2_X1 U11928 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n10205), .Z(n10199) );
  XNOR2_X1 U11929 ( .A(n10199), .B(n10479), .ZN(n11373) );
  INV_X1 U11930 ( .A(n10199), .ZN(n10200) );
  AND2_X1 U11931 ( .A1(n10200), .A2(n10479), .ZN(n10201) );
  AOI21_X1 U11932 ( .B1(n11372), .B2(n11373), .A(n10201), .ZN(n16016) );
  MUX2_X1 U11933 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n10205), .Z(n10202) );
  XNOR2_X1 U11934 ( .A(n10202), .B(n10478), .ZN(n16015) );
  MUX2_X1 U11935 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n10205), .Z(n10203) );
  XOR2_X1 U11936 ( .A(n10471), .B(n10203), .Z(n11627) );
  INV_X1 U11937 ( .A(n10471), .ZN(n11626) );
  INV_X1 U11938 ( .A(n10203), .ZN(n10204) );
  AOI22_X1 U11939 ( .A1(n11628), .A2(n11627), .B1(n11626), .B2(n10204), .ZN(
        n12150) );
  MUX2_X1 U11940 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n10205), .Z(n10206) );
  XNOR2_X1 U11941 ( .A(n10206), .B(n12153), .ZN(n12149) );
  OAI22_X1 U11942 ( .A1(n12150), .A2(n12149), .B1(n10206), .B2(n12153), .ZN(
        n12135) );
  MUX2_X1 U11943 ( .A(n12141), .B(n12129), .S(n14141), .Z(n12136) );
  NOR2_X1 U11944 ( .A1(n12135), .A2(n12136), .ZN(n12134) );
  MUX2_X1 U11945 ( .A(n10208), .B(n10207), .S(n14141), .Z(n10209) );
  XNOR2_X1 U11946 ( .A(n10211), .B(n10210), .ZN(n14063) );
  NAND2_X1 U11947 ( .A1(n14064), .A2(n14063), .ZN(n14062) );
  OAI21_X1 U11948 ( .B1(n10211), .B2(n14072), .A(n14062), .ZN(n10212) );
  INV_X1 U11949 ( .A(n16017), .ZN(n15960) );
  NOR2_X1 U11950 ( .A1(n10212), .A2(n10213), .ZN(n10241) );
  AOI211_X1 U11951 ( .C1(n10213), .C2(n10212), .A(n15960), .B(n10241), .ZN(
        n10221) );
  INV_X1 U11952 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n10218) );
  NOR2_X1 U11953 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10218), .ZN(n13937) );
  AOI21_X1 U11954 ( .B1(n15646), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n13937), 
        .ZN(n10219) );
  OAI21_X1 U11955 ( .B1(n15997), .B2(n10729), .A(n10219), .ZN(n10220) );
  NAND2_X1 U11956 ( .A1(n10225), .A2(n10224), .ZN(n10227) );
  INV_X1 U11957 ( .A(n10227), .ZN(n10226) );
  NOR2_X1 U11958 ( .A1(n7905), .A2(n10226), .ZN(n10228) );
  XNOR2_X1 U11959 ( .A(n10227), .B(n14085), .ZN(n14079) );
  OR2_X1 U11960 ( .A1(n14094), .A2(n10229), .ZN(n14106) );
  NAND2_X1 U11961 ( .A1(n14094), .A2(n10229), .ZN(n10230) );
  NAND2_X1 U11962 ( .A1(n14106), .A2(n10230), .ZN(n10231) );
  NAND2_X1 U11963 ( .A1(n10232), .A2(n10231), .ZN(n10233) );
  AOI21_X1 U11964 ( .B1(n14107), .B2(n10233), .A(n16009), .ZN(n10251) );
  NOR2_X1 U11965 ( .A1(n7905), .A2(n10236), .ZN(n10237) );
  XNOR2_X1 U11966 ( .A(n14094), .B(n14412), .ZN(n10238) );
  NAND2_X1 U11967 ( .A1(n10239), .A2(n10238), .ZN(n10240) );
  AOI21_X1 U11968 ( .B1(n14096), .B2(n10240), .A(n16013), .ZN(n10250) );
  MUX2_X1 U11969 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n14141), .Z(n14101) );
  XOR2_X1 U11970 ( .A(n14094), .B(n14101), .Z(n10246) );
  INV_X1 U11971 ( .A(n10243), .ZN(n10244) );
  XNOR2_X1 U11972 ( .A(n10243), .B(n14085), .ZN(n14082) );
  MUX2_X1 U11973 ( .A(n14078), .B(n14416), .S(n14141), .Z(n14081) );
  NAND2_X1 U11974 ( .A1(n14082), .A2(n14081), .ZN(n14080) );
  OAI21_X1 U11975 ( .B1(n10244), .B2(n14085), .A(n14080), .ZN(n10245) );
  NOR2_X1 U11976 ( .A1(n10245), .A2(n10246), .ZN(n14099) );
  AOI211_X1 U11977 ( .C1(n10246), .C2(n10245), .A(n15960), .B(n14099), .ZN(
        n10249) );
  INV_X1 U11978 ( .A(n14094), .ZN(n14100) );
  NAND2_X1 U11979 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(P3_U3151), .ZN(n13975)
         );
  NAND2_X1 U11980 ( .A1(n15646), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n10247) );
  OAI211_X1 U11981 ( .C1(n15997), .C2(n14100), .A(n13975), .B(n10247), .ZN(
        n10248) );
  INV_X1 U11982 ( .A(n10252), .ZN(n10253) );
  AOI211_X1 U11983 ( .C1(n10255), .C2(n10254), .A(n14041), .B(n10253), .ZN(
        n10260) );
  NOR2_X1 U11984 ( .A1(n14036), .A2(n12329), .ZN(n10259) );
  INV_X1 U11985 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n10256) );
  OR2_X1 U11986 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10256), .ZN(n11619) );
  OAI21_X1 U11987 ( .B1(n14017), .B2(n12473), .A(n11619), .ZN(n10258) );
  INV_X1 U11988 ( .A(n12322), .ZN(n13200) );
  OAI22_X1 U11989 ( .A1(n12332), .A2(n14015), .B1(n14032), .B2(n13200), .ZN(
        n10257) );
  OR4_X1 U11990 ( .A1(n10260), .A2(n10259), .A3(n10258), .A4(n10257), .ZN(
        P3_U3157) );
  INV_X1 U11991 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n10262) );
  AND3_X1 U11992 ( .A1(n10263), .A2(n10262), .A3(n10261), .ZN(n10267) );
  NOR2_X1 U11993 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), 
        .ZN(n10266) );
  NOR2_X1 U11994 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), 
        .ZN(n10265) );
  NOR2_X1 U11995 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), 
        .ZN(n10264) );
  XNOR2_X2 U11996 ( .A(n10268), .B(P2_IR_REG_30__SCAN_IN), .ZN(n10271) );
  BUF_X2 U11997 ( .A(n10269), .Z(n10293) );
  AND2_X2 U11998 ( .A1(n10271), .A2(n10272), .ZN(n12110) );
  NAND2_X1 U11999 ( .A1(n12110), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n10276) );
  INV_X1 U12000 ( .A(n10272), .ZN(n15056) );
  AND2_X2 U12001 ( .A1(n10271), .A2(n15056), .ZN(n10326) );
  NAND2_X1 U12002 ( .A1(n10326), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n10275) );
  AND2_X2 U12003 ( .A1(n13329), .A2(n10272), .ZN(n10327) );
  NAND2_X1 U12004 ( .A1(n10327), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10274) );
  AND2_X2 U12005 ( .A1(n13329), .A2(n15056), .ZN(n10328) );
  NAND2_X1 U12006 ( .A1(n10328), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n10273) );
  NAND2_X1 U12007 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), 
        .ZN(n10278) );
  NOR2_X1 U12008 ( .A1(n10282), .A2(n10281), .ZN(n10284) );
  NAND3_X1 U12009 ( .A1(n10285), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_IR_REG_22__SCAN_IN), .ZN(n10283) );
  NAND2_X2 U12010 ( .A1(n10283), .A2(n10284), .ZN(n13902) );
  OR2_X2 U12011 ( .A1(n7420), .A2(n13662), .ZN(n10663) );
  AOI21_X1 U12012 ( .B1(n10291), .B2(n10287), .A(n10411), .ZN(n10290) );
  MUX2_X2 U12013 ( .A(n10290), .B(n10289), .S(n10288), .Z(n13912) );
  INV_X2 U12014 ( .A(n10938), .ZN(n11126) );
  NAND2_X1 U12015 ( .A1(n7423), .A2(n11126), .ZN(n10320) );
  NAND2_X2 U12016 ( .A1(n10293), .A2(n10292), .ZN(n10370) );
  OR2_X1 U12017 ( .A1(n10294), .A2(n10411), .ZN(n10296) );
  XNOR2_X1 U12018 ( .A(n10296), .B(n10295), .ZN(n14698) );
  OR2_X1 U12019 ( .A1(n10322), .A2(n10407), .ZN(n10298) );
  OR2_X1 U12020 ( .A1(n10312), .A2(n10421), .ZN(n10297) );
  OAI211_X2 U12021 ( .C1(n11131), .C2(n14698), .A(n10298), .B(n10297), .ZN(
        n14626) );
  NAND2_X1 U12022 ( .A1(n12110), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n10302) );
  NAND2_X1 U12023 ( .A1(n10328), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n10301) );
  NAND2_X1 U12024 ( .A1(n10326), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n10299) );
  INV_X1 U12025 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n15659) );
  NAND2_X1 U12026 ( .A1(n10432), .A2(SI_0_), .ZN(n10304) );
  NAND2_X1 U12027 ( .A1(n10304), .A2(n10303), .ZN(n10306) );
  NAND2_X1 U12028 ( .A1(n10306), .A2(n10305), .ZN(n15074) );
  OAI21_X2 U12029 ( .B1(n11131), .B2(P2_IR_REG_0__SCAN_IN), .A(n10307), .ZN(
        n13667) );
  OR2_X1 U12030 ( .A1(n10767), .A2(n10938), .ZN(n10941) );
  NAND2_X1 U12031 ( .A1(n14487), .A2(n13667), .ZN(n10308) );
  NAND2_X1 U12032 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n10309) );
  MUX2_X1 U12033 ( .A(P2_IR_REG_31__SCAN_IN), .B(n10309), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n10311) );
  INV_X1 U12034 ( .A(n10294), .ZN(n10310) );
  NAND2_X1 U12035 ( .A1(n10311), .A2(n10310), .ZN(n15652) );
  XNOR2_X1 U12036 ( .A(n11125), .B(n7432), .ZN(n10318) );
  NAND2_X1 U12037 ( .A1(n12110), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n10316) );
  NAND2_X1 U12038 ( .A1(n10326), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10315) );
  NAND2_X1 U12039 ( .A1(n14691), .A2(n11126), .ZN(n10317) );
  INV_X1 U12040 ( .A(n10317), .ZN(n10319) );
  NOR2_X1 U12041 ( .A1(n10319), .A2(n10318), .ZN(n14629) );
  OR2_X1 U12042 ( .A1(n13618), .A2(n10408), .ZN(n10325) );
  OR2_X1 U12043 ( .A1(n10410), .A2(n10411), .ZN(n10323) );
  XNOR2_X1 U12044 ( .A(n10323), .B(n10409), .ZN(n14714) );
  OR2_X1 U12045 ( .A1(n11131), .A2(n14714), .ZN(n10324) );
  XNOR2_X1 U12046 ( .A(n14525), .B(n13695), .ZN(n10334) );
  INV_X1 U12047 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n14706) );
  NAND2_X1 U12048 ( .A1(n13522), .A2(n14706), .ZN(n10332) );
  NAND2_X1 U12049 ( .A1(n10326), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10331) );
  NAND2_X1 U12050 ( .A1(n7425), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10330) );
  NAND2_X1 U12051 ( .A1(n13517), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n10329) );
  AND2_X1 U12052 ( .A1(n14689), .A2(n11126), .ZN(n10333) );
  NAND2_X1 U12053 ( .A1(n10334), .A2(n10333), .ZN(n11122) );
  OAI21_X1 U12054 ( .B1(n10334), .B2(n10333), .A(n11122), .ZN(n10361) );
  INV_X1 U12055 ( .A(P2_B_REG_SCAN_IN), .ZN(n13901) );
  AOI22_X1 U12056 ( .A1(P2_B_REG_SCAN_IN), .A2(n13240), .B1(n10352), .B2(
        n13901), .ZN(n10335) );
  OR2_X1 U12057 ( .A1(n15071), .A2(n10335), .ZN(n10336) );
  INV_X1 U12058 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10337) );
  NAND2_X1 U12059 ( .A1(n15643), .A2(n10337), .ZN(n10339) );
  OR2_X1 U12060 ( .A1(n15066), .A2(n15071), .ZN(n10338) );
  NAND2_X1 U12061 ( .A1(n10339), .A2(n10338), .ZN(n11359) );
  NOR4_X1 U12062 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n10343) );
  NOR4_X1 U12063 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n10342) );
  NOR4_X1 U12064 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n10341) );
  NOR4_X1 U12065 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n10340) );
  NAND4_X1 U12066 ( .A1(n10343), .A2(n10342), .A3(n10341), .A4(n10340), .ZN(
        n10349) );
  NOR2_X1 U12067 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n10347) );
  NOR4_X1 U12068 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n10346) );
  NOR4_X1 U12069 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n10345) );
  NOR4_X1 U12070 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n10344) );
  NAND4_X1 U12071 ( .A1(n10347), .A2(n10346), .A3(n10345), .A4(n10344), .ZN(
        n10348) );
  OAI21_X1 U12072 ( .B1(n10349), .B2(n10348), .A(n15643), .ZN(n10657) );
  INV_X1 U12073 ( .A(n10657), .ZN(n10350) );
  NOR2_X1 U12074 ( .A1(n11359), .A2(n10350), .ZN(n10355) );
  INV_X1 U12075 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10351) );
  NAND2_X1 U12076 ( .A1(n15643), .A2(n10351), .ZN(n10354) );
  NAND2_X1 U12077 ( .A1(n10355), .A2(n15648), .ZN(n10369) );
  AND2_X1 U12078 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10366), .ZN(n10356) );
  INV_X1 U12079 ( .A(n15647), .ZN(n15649) );
  INV_X1 U12080 ( .A(n10364), .ZN(n10360) );
  INV_X1 U12081 ( .A(n10663), .ZN(n10357) );
  NAND2_X1 U12082 ( .A1(n13912), .A2(n15711), .ZN(n13904) );
  INV_X1 U12083 ( .A(n10539), .ZN(n10358) );
  NAND2_X1 U12084 ( .A1(n16307), .A2(n10358), .ZN(n10359) );
  NOR2_X1 U12085 ( .A1(n10362), .A2(n10361), .ZN(n11124) );
  AOI211_X1 U12086 ( .C1(n10362), .C2(n10361), .A(n14642), .B(n11124), .ZN(
        n10382) );
  INV_X1 U12087 ( .A(n13662), .ZN(n13899) );
  NAND2_X1 U12088 ( .A1(n8074), .A2(n13899), .ZN(n13894) );
  NOR2_X1 U12089 ( .A1(n13894), .A2(n7420), .ZN(n11364) );
  AND2_X1 U12090 ( .A1(n15027), .A2(n7415), .ZN(n10658) );
  NOR2_X1 U12091 ( .A1(n14670), .A2(n11422), .ZN(n10381) );
  INV_X1 U12092 ( .A(n10658), .ZN(n10365) );
  NAND2_X1 U12093 ( .A1(n10369), .A2(n10365), .ZN(n10368) );
  AND2_X1 U12094 ( .A1(n13904), .A2(n13662), .ZN(n13862) );
  NAND2_X1 U12095 ( .A1(n13862), .A2(n7420), .ZN(n10656) );
  AND3_X1 U12096 ( .A1(n10656), .A2(n10366), .A3(n13243), .ZN(n10367) );
  NAND2_X1 U12097 ( .A1(n10368), .A2(n10367), .ZN(n10937) );
  OR3_X1 U12098 ( .A1(n10369), .A2(n15649), .A3(n13904), .ZN(n10373) );
  INV_X1 U12099 ( .A(n10373), .ZN(n10372) );
  INV_X1 U12100 ( .A(n10370), .ZN(n10371) );
  OAI22_X1 U12101 ( .A1(n14638), .A2(P2_REG3_REG_3__SCAN_IN), .B1(n7422), .B2(
        n14661), .ZN(n10380) );
  NAND2_X1 U12102 ( .A1(n13523), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n10378) );
  NAND2_X1 U12103 ( .A1(n7425), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10377) );
  INV_X1 U12104 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10374) );
  XNOR2_X1 U12105 ( .A(n10374), .B(P2_REG3_REG_3__SCAN_IN), .ZN(n11456) );
  NAND2_X1 U12106 ( .A1(n13522), .A2(n11456), .ZN(n10376) );
  NAND2_X1 U12107 ( .A1(n13517), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n10375) );
  NAND4_X1 U12108 ( .A1(n10378), .A2(n10377), .A3(n10376), .A4(n10375), .ZN(
        n14688) );
  INV_X1 U12109 ( .A(n14688), .ZN(n11394) );
  OAI22_X1 U12110 ( .A1(n14663), .A2(n11394), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14706), .ZN(n10379) );
  OR4_X1 U12111 ( .A1(n10382), .A2(n10381), .A3(n10380), .A4(n10379), .ZN(
        P2_U3190) );
  NAND2_X1 U12112 ( .A1(n10383), .A2(n10396), .ZN(n10384) );
  NAND3_X1 U12113 ( .A1(n10385), .A2(n9714), .A3(n10384), .ZN(n10387) );
  NAND2_X1 U12114 ( .A1(n11806), .A2(n14304), .ZN(n10386) );
  NAND2_X1 U12115 ( .A1(n10387), .A2(n10386), .ZN(n11428) );
  NAND2_X1 U12116 ( .A1(n14466), .A2(n10388), .ZN(n10389) );
  OAI21_X1 U12117 ( .B1(n14466), .B2(n10390), .A(n10389), .ZN(n10391) );
  INV_X1 U12118 ( .A(n10391), .ZN(n10392) );
  NAND2_X1 U12119 ( .A1(n10393), .A2(n10392), .ZN(n10401) );
  NOR2_X1 U12120 ( .A1(n16231), .A2(n11435), .ZN(n10394) );
  MUX2_X1 U12121 ( .A(n11428), .B(P3_REG2_REG_3__SCAN_IN), .S(n14341), .Z(
        n10406) );
  OR2_X1 U12122 ( .A1(n10397), .A2(n10396), .ZN(n10398) );
  NAND2_X1 U12123 ( .A1(n10399), .A2(n10398), .ZN(n11430) );
  NAND2_X1 U12124 ( .A1(n10400), .A2(n16061), .ZN(n12597) );
  NAND2_X1 U12125 ( .A1(n14256), .A2(n12597), .ZN(n16088) );
  NAND2_X1 U12126 ( .A1(n11430), .A2(n14339), .ZN(n10404) );
  NAND2_X1 U12127 ( .A1(n16100), .A2(n14384), .ZN(n14284) );
  INV_X1 U12128 ( .A(n14284), .ZN(n12291) );
  OAI22_X1 U12129 ( .A1(n14337), .A2(n11522), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(n16059), .ZN(n10402) );
  AOI21_X1 U12130 ( .B1(n12291), .B2(n14058), .A(n10402), .ZN(n10403) );
  NAND2_X1 U12131 ( .A1(n10404), .A2(n10403), .ZN(n10405) );
  OR2_X1 U12132 ( .A1(n10406), .A2(n10405), .ZN(P3_U3230) );
  INV_X2 U12133 ( .A(n13242), .ZN(n15061) );
  OAI222_X1 U12134 ( .A1(n13255), .A2(n10407), .B1(n15061), .B2(n10421), .C1(
        P2_U3088), .C2(n14698), .ZN(P2_U3325) );
  OAI222_X1 U12135 ( .A1(n13255), .A2(n10408), .B1(n15061), .B2(n10429), .C1(
        P2_U3088), .C2(n14714), .ZN(P2_U3324) );
  INV_X1 U12136 ( .A(n11043), .ZN(n10427) );
  NOR2_X1 U12137 ( .A1(n10722), .A2(n10411), .ZN(n10412) );
  MUX2_X1 U12138 ( .A(n10411), .B(n10412), .S(P2_IR_REG_4__SCAN_IN), .Z(n10413) );
  INV_X1 U12139 ( .A(n10413), .ZN(n10415) );
  NAND2_X1 U12140 ( .A1(n10722), .A2(n10414), .ZN(n10419) );
  NAND2_X1 U12141 ( .A1(n10415), .A2(n10419), .ZN(n11047) );
  OAI222_X1 U12142 ( .A1(n13255), .A2(n11044), .B1(n15061), .B2(n10427), .C1(
        P2_U3088), .C2(n11047), .ZN(P2_U3323) );
  INV_X1 U12143 ( .A(n11130), .ZN(n10422) );
  NAND2_X1 U12144 ( .A1(n10419), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10416) );
  XNOR2_X1 U12145 ( .A(n10416), .B(P2_IR_REG_5__SCAN_IN), .ZN(n11132) );
  INV_X1 U12146 ( .A(n11132), .ZN(n10417) );
  OAI222_X1 U12147 ( .A1(n13255), .A2(n10418), .B1(n15061), .B2(n10422), .C1(
        P2_U3088), .C2(n10417), .ZN(P2_U3322) );
  INV_X1 U12148 ( .A(n11539), .ZN(n10424) );
  NAND2_X1 U12149 ( .A1(n10651), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10446) );
  XNOR2_X1 U12150 ( .A(n10446), .B(P2_IR_REG_6__SCAN_IN), .ZN(n11540) );
  INV_X1 U12151 ( .A(n11540), .ZN(n15667) );
  OAI222_X1 U12152 ( .A1(n13255), .A2(n7773), .B1(n15061), .B2(n10424), .C1(
        P2_U3088), .C2(n15667), .ZN(P2_U3321) );
  INV_X2 U12153 ( .A(n15601), .ZN(n15597) );
  OAI222_X1 U12154 ( .A1(n15597), .A2(n7749), .B1(n15604), .B2(n10421), .C1(
        P1_U3086), .C2(n10972), .ZN(P1_U3353) );
  INV_X1 U12155 ( .A(n10680), .ZN(n10685) );
  OAI222_X1 U12156 ( .A1(n15597), .A2(n10423), .B1(n15604), .B2(n10422), .C1(
        P1_U3086), .C2(n10685), .ZN(P1_U3350) );
  INV_X1 U12157 ( .A(n10687), .ZN(n10799) );
  OAI222_X1 U12158 ( .A1(n15597), .A2(n10425), .B1(n15604), .B2(n10424), .C1(
        P1_U3086), .C2(n10799), .ZN(P1_U3349) );
  INV_X1 U12159 ( .A(n10817), .ZN(n10426) );
  OAI222_X1 U12160 ( .A1(n15597), .A2(n10428), .B1(n15604), .B2(n10427), .C1(
        P1_U3086), .C2(n10426), .ZN(P1_U3351) );
  INV_X1 U12161 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10430) );
  INV_X1 U12162 ( .A(n10623), .ZN(n10785) );
  OAI222_X1 U12163 ( .A1(n15597), .A2(n10430), .B1(n15604), .B2(n10429), .C1(
        P1_U3086), .C2(n10785), .ZN(P1_U3352) );
  INV_X2 U12164 ( .A(n14474), .ZN(n13924) );
  OAI222_X1 U12165 ( .A1(n13924), .A2(n10434), .B1(n13926), .B2(n10433), .C1(
        P3_U3151), .C2(n15984), .ZN(P3_U3289) );
  INV_X1 U12166 ( .A(SI_5_), .ZN(n10437) );
  INV_X1 U12167 ( .A(n10435), .ZN(n10436) );
  OAI222_X1 U12168 ( .A1(P3_U3151), .A2(n11024), .B1(n13926), .B2(n10437), 
        .C1(n13924), .C2(n10436), .ZN(P3_U3290) );
  INV_X1 U12169 ( .A(n10438), .ZN(n10439) );
  OAI222_X1 U12170 ( .A1(P3_U3151), .A2(n10441), .B1(n13926), .B2(n10440), 
        .C1(n13924), .C2(n10439), .ZN(P3_U3292) );
  INV_X1 U12171 ( .A(SI_4_), .ZN(n10444) );
  INV_X1 U12172 ( .A(n10442), .ZN(n10443) );
  OAI222_X1 U12173 ( .A1(P3_U3151), .A2(n10867), .B1(n13926), .B2(n10444), 
        .C1(n13924), .C2(n10443), .ZN(P3_U3291) );
  INV_X1 U12174 ( .A(n11543), .ZN(n10450) );
  INV_X1 U12175 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n10445) );
  NAND2_X1 U12176 ( .A1(n10446), .A2(n10445), .ZN(n10447) );
  NAND2_X1 U12177 ( .A1(n10447), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10458) );
  XNOR2_X1 U12178 ( .A(n10458), .B(P2_IR_REG_7__SCAN_IN), .ZN(n11544) );
  INV_X1 U12179 ( .A(n11544), .ZN(n10448) );
  OAI222_X1 U12180 ( .A1(n13255), .A2(n10449), .B1(n15061), .B2(n10450), .C1(
        P2_U3088), .C2(n10448), .ZN(P2_U3320) );
  INV_X1 U12181 ( .A(n10756), .ZN(n10750) );
  OAI222_X1 U12182 ( .A1(n15597), .A2(n10451), .B1(n15604), .B2(n10450), .C1(
        P1_U3086), .C2(n10750), .ZN(P1_U3348) );
  NAND2_X1 U12183 ( .A1(n15583), .A2(n10453), .ZN(n10611) );
  OR2_X1 U12184 ( .A1(n10529), .A2(n10454), .ZN(n10456) );
  AND2_X1 U12185 ( .A1(n10456), .A2(n10455), .ZN(n10610) );
  INV_X1 U12186 ( .A(n10610), .ZN(n10457) );
  AND2_X1 U12187 ( .A1(n10611), .A2(n10457), .ZN(n15757) );
  NOR2_X1 U12188 ( .A1(n15757), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U12189 ( .A(n11671), .ZN(n10462) );
  NAND2_X1 U12190 ( .A1(n10458), .A2(n10646), .ZN(n10459) );
  NAND2_X1 U12191 ( .A1(n10459), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10485) );
  XNOR2_X1 U12192 ( .A(n10485), .B(P2_IR_REG_8__SCAN_IN), .ZN(n11672) );
  INV_X1 U12193 ( .A(n11672), .ZN(n10460) );
  OAI222_X1 U12194 ( .A1(n13255), .A2(n10461), .B1(n15061), .B2(n10462), .C1(
        P2_U3088), .C2(n10460), .ZN(P2_U3319) );
  INV_X1 U12195 ( .A(n10758), .ZN(n10930) );
  OAI222_X1 U12196 ( .A1(n15597), .A2(n10463), .B1(n15604), .B2(n10462), .C1(
        P1_U3086), .C2(n10930), .ZN(P1_U3347) );
  INV_X1 U12197 ( .A(n10466), .ZN(n15998) );
  INV_X1 U12198 ( .A(SI_7_), .ZN(n10469) );
  INV_X1 U12199 ( .A(n10467), .ZN(n10468) );
  OAI222_X1 U12200 ( .A1(P3_U3151), .A2(n15998), .B1(n13926), .B2(n10469), 
        .C1(n13924), .C2(n10468), .ZN(P3_U3288) );
  INV_X1 U12201 ( .A(SI_10_), .ZN(n12745) );
  OAI222_X1 U12202 ( .A1(P3_U3151), .A2(n10471), .B1(n13926), .B2(n12745), 
        .C1(n13924), .C2(n10470), .ZN(P3_U3285) );
  INV_X1 U12203 ( .A(n10472), .ZN(n10473) );
  OAI222_X1 U12204 ( .A1(n10842), .A2(P3_U3151), .B1(n13924), .B2(n10473), 
        .C1(n12761), .C2(n13926), .ZN(P3_U3293) );
  OAI222_X1 U12205 ( .A1(n10475), .A2(P3_U3151), .B1(n13924), .B2(n10474), 
        .C1(n12989), .C2(n13926), .ZN(P3_U3294) );
  INV_X1 U12206 ( .A(n10476), .ZN(n10477) );
  INV_X1 U12207 ( .A(SI_9_), .ZN(n12974) );
  OAI222_X1 U12208 ( .A1(n10478), .A2(P3_U3151), .B1(n13924), .B2(n10477), 
        .C1(n12974), .C2(n13926), .ZN(P3_U3286) );
  INV_X1 U12209 ( .A(n10479), .ZN(n11378) );
  OAI222_X1 U12210 ( .A1(n11378), .A2(P3_U3151), .B1(n13924), .B2(n10481), 
        .C1(n10480), .C2(n13926), .ZN(P3_U3287) );
  OAI222_X1 U12211 ( .A1(P3_U3151), .A2(n12153), .B1(n13926), .B2(n12973), 
        .C1(n13924), .C2(n10482), .ZN(P3_U3284) );
  INV_X1 U12212 ( .A(n11854), .ZN(n10487) );
  INV_X1 U12213 ( .A(n11175), .ZN(n11179) );
  OAI222_X1 U12214 ( .A1(n15597), .A2(n10483), .B1(n15604), .B2(n10487), .C1(
        P1_U3086), .C2(n11179), .ZN(P1_U3346) );
  INV_X1 U12215 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n10484) );
  NAND2_X1 U12216 ( .A1(n10485), .A2(n10484), .ZN(n10486) );
  NAND2_X1 U12217 ( .A1(n10486), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10491) );
  XNOR2_X1 U12218 ( .A(n10491), .B(P2_IR_REG_9__SCAN_IN), .ZN(n11855) );
  INV_X1 U12219 ( .A(n11855), .ZN(n10986) );
  OAI222_X1 U12220 ( .A1(n13255), .A2(n10488), .B1(n15061), .B2(n10487), .C1(
        P2_U3088), .C2(n10986), .ZN(P2_U3318) );
  OAI222_X1 U12221 ( .A1(P3_U3151), .A2(n12131), .B1(n13926), .B2(n12970), 
        .C1(n13924), .C2(n10489), .ZN(P3_U3283) );
  AND2_X1 U12222 ( .A1(n10645), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U12223 ( .A1(n10645), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U12224 ( .A1(n10645), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U12225 ( .A1(n10645), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U12226 ( .A1(n10645), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U12227 ( .A1(n10645), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U12228 ( .A1(n10645), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U12229 ( .A1(n10645), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U12230 ( .A1(n10645), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U12231 ( .A1(n10645), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U12232 ( .A1(n10645), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U12233 ( .A1(n10645), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U12234 ( .A1(n10645), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U12235 ( .A1(n10645), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U12236 ( .A1(n10645), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U12237 ( .A1(n10645), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  INV_X1 U12238 ( .A(n11860), .ZN(n10495) );
  INV_X1 U12239 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n10490) );
  NAND2_X1 U12240 ( .A1(n10491), .A2(n10490), .ZN(n10492) );
  NAND2_X1 U12241 ( .A1(n10492), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10498) );
  XNOR2_X1 U12242 ( .A(n10498), .B(P2_IR_REG_10__SCAN_IN), .ZN(n15742) );
  INV_X1 U12243 ( .A(n15742), .ZN(n10493) );
  OAI222_X1 U12244 ( .A1(n13255), .A2(n10494), .B1(n15061), .B2(n10495), .C1(
        P2_U3088), .C2(n10493), .ZN(P2_U3317) );
  INV_X1 U12245 ( .A(n11319), .ZN(n11189) );
  OAI222_X1 U12246 ( .A1(n15597), .A2(n10496), .B1(n15604), .B2(n10495), .C1(
        P1_U3086), .C2(n11189), .ZN(P1_U3345) );
  INV_X1 U12247 ( .A(n12020), .ZN(n10502) );
  INV_X1 U12248 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n10497) );
  NAND2_X1 U12249 ( .A1(n10498), .A2(n10497), .ZN(n10499) );
  NAND2_X1 U12250 ( .A1(n10499), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10500) );
  XNOR2_X1 U12251 ( .A(n10500), .B(P2_IR_REG_11__SCAN_IN), .ZN(n12021) );
  INV_X1 U12252 ( .A(n12021), .ZN(n11348) );
  OAI222_X1 U12253 ( .A1(n13255), .A2(n10501), .B1(n15061), .B2(n10502), .C1(
        P2_U3088), .C2(n11348), .ZN(P2_U3316) );
  OAI222_X1 U12254 ( .A1(n10503), .A2(n15597), .B1(P1_U3086), .B2(n7717), .C1(
        n15604), .C2(n10502), .ZN(P1_U3344) );
  NAND2_X1 U12255 ( .A1(n10504), .A2(P1_B_REG_SCAN_IN), .ZN(n10507) );
  INV_X1 U12256 ( .A(n15600), .ZN(n10519) );
  OAI21_X1 U12257 ( .B1(n10504), .B2(P1_B_REG_SCAN_IN), .A(n10519), .ZN(n10505) );
  INV_X1 U12258 ( .A(n10505), .ZN(n10506) );
  NOR4_X1 U12259 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n10511) );
  NOR4_X1 U12260 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n10510) );
  NOR4_X1 U12261 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n10509) );
  NOR4_X1 U12262 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n10508) );
  NAND4_X1 U12263 ( .A1(n10511), .A2(n10510), .A3(n10509), .A4(n10508), .ZN(
        n10517) );
  NOR2_X1 U12264 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .ZN(
        n10515) );
  NOR4_X1 U12265 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n10514) );
  NOR4_X1 U12266 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n10513) );
  NOR4_X1 U12267 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n10512) );
  NAND4_X1 U12268 ( .A1(n10515), .A2(n10514), .A3(n10513), .A4(n10512), .ZN(
        n10516) );
  NOR2_X1 U12269 ( .A1(n10517), .A2(n10516), .ZN(n10518) );
  OR2_X1 U12270 ( .A1(n15582), .A2(n10518), .ZN(n10868) );
  INV_X1 U12271 ( .A(n10868), .ZN(n10521) );
  OR2_X1 U12272 ( .A1(n15582), .A2(P1_D_REG_1__SCAN_IN), .ZN(n10520) );
  OR2_X1 U12273 ( .A1(n15602), .A2(n10519), .ZN(n15585) );
  NAND2_X1 U12274 ( .A1(n10520), .A2(n15585), .ZN(n10870) );
  NOR2_X1 U12275 ( .A1(n10521), .A2(n10870), .ZN(n11072) );
  OR2_X1 U12276 ( .A1(n15582), .A2(P1_D_REG_0__SCAN_IN), .ZN(n10522) );
  NAND2_X1 U12277 ( .A1(n10504), .A2(n15600), .ZN(n15586) );
  NAND2_X1 U12278 ( .A1(n11072), .A2(n10891), .ZN(n10526) );
  NAND2_X1 U12279 ( .A1(n10528), .A2(n8224), .ZN(n16174) );
  INV_X1 U12280 ( .A(n15583), .ZN(n10524) );
  NAND2_X1 U12281 ( .A1(n16247), .A2(n7429), .ZN(n10869) );
  INV_X1 U12282 ( .A(n10869), .ZN(n10523) );
  INV_X1 U12283 ( .A(n11071), .ZN(n10525) );
  OR2_X1 U12284 ( .A1(n10526), .A2(n10525), .ZN(n15132) );
  INV_X1 U12285 ( .A(n15132), .ZN(n15153) );
  OR2_X1 U12286 ( .A1(n10529), .A2(n10804), .ZN(n15408) );
  NAND2_X1 U12287 ( .A1(n15153), .A2(n15457), .ZN(n15170) );
  INV_X1 U12288 ( .A(n15170), .ZN(n16351) );
  NAND2_X1 U12289 ( .A1(n10526), .A2(n10869), .ZN(n10956) );
  NAND2_X1 U12290 ( .A1(n10956), .A2(n11071), .ZN(n10675) );
  AOI22_X1 U12291 ( .A1(n16351), .A2(n15195), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n10675), .ZN(n10537) );
  INV_X1 U12292 ( .A(n10527), .ZN(n10531) );
  AND2_X1 U12293 ( .A1(n16333), .A2(n10529), .ZN(n10530) );
  NOR2_X1 U12294 ( .A1(n16031), .A2(n10533), .ZN(n11078) );
  OR2_X4 U12295 ( .A1(n13594), .A2(n11078), .ZN(n13587) );
  INV_X1 U12296 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10606) );
  OAI222_X1 U12297 ( .A1(n13588), .A2(n16032), .B1(n13587), .B2(n10534), .C1(
        n10606), .C2(n10535), .ZN(n10578) );
  OAI222_X1 U12298 ( .A1(n10535), .A2(n15751), .B1(n10669), .B2(n10534), .C1(
        n16032), .C2(n13594), .ZN(n10577) );
  XOR2_X1 U12299 ( .A(n10578), .B(n10577), .Z(n10805) );
  NAND2_X1 U12300 ( .A1(n16356), .A2(n10805), .ZN(n10536) );
  OAI211_X1 U12301 ( .C1(n16353), .C2(n16032), .A(n10537), .B(n10536), .ZN(
        P1_U3232) );
  INV_X1 U12302 ( .A(n10538), .ZN(n10542) );
  NAND2_X1 U12303 ( .A1(n10539), .A2(n13243), .ZN(n10540) );
  NAND2_X1 U12304 ( .A1(n10540), .A2(n11131), .ZN(n10541) );
  INV_X1 U12305 ( .A(n15683), .ZN(n15749) );
  NAND2_X1 U12306 ( .A1(n10370), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10543) );
  OR2_X1 U12307 ( .A1(n10544), .A2(n10543), .ZN(n15724) );
  INV_X1 U12308 ( .A(n11047), .ZN(n10585) );
  NAND2_X1 U12309 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n11197) );
  INV_X1 U12310 ( .A(n10544), .ZN(n10545) );
  NOR2_X1 U12311 ( .A1(n10370), .A2(P2_U3088), .ZN(n15058) );
  INV_X1 U12312 ( .A(n14714), .ZN(n10562) );
  INV_X1 U12313 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10776) );
  MUX2_X1 U12314 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n10776), .S(n15652), .Z(
        n15658) );
  INV_X1 U12315 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10546) );
  NOR3_X1 U12316 ( .A1(n15658), .A2(n10546), .A3(n15659), .ZN(n15657) );
  NOR2_X1 U12317 ( .A1(n15652), .A2(n10776), .ZN(n14694) );
  INV_X1 U12318 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10547) );
  MUX2_X1 U12319 ( .A(n10547), .B(P2_REG1_REG_2__SCAN_IN), .S(n14698), .Z(
        n10548) );
  OAI21_X1 U12320 ( .B1(n15657), .B2(n14694), .A(n10548), .ZN(n14711) );
  INV_X1 U12321 ( .A(n14698), .ZN(n10558) );
  NAND2_X1 U12322 ( .A1(n10558), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n14710) );
  INV_X1 U12323 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n11215) );
  MUX2_X1 U12324 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n11215), .S(n14714), .Z(
        n14709) );
  AOI21_X1 U12325 ( .B1(n14711), .B2(n14710), .A(n14709), .ZN(n14708) );
  AOI21_X1 U12326 ( .B1(P2_REG1_REG_3__SCAN_IN), .B2(n10562), .A(n14708), .ZN(
        n10550) );
  INV_X1 U12327 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10584) );
  MUX2_X1 U12328 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n10584), .S(n11047), .Z(
        n10549) );
  OR2_X1 U12329 ( .A1(n10550), .A2(n10549), .ZN(n10588) );
  NAND2_X1 U12330 ( .A1(n10550), .A2(n10549), .ZN(n10551) );
  NAND3_X1 U12331 ( .A1(n15743), .A2(n10588), .A3(n10551), .ZN(n10552) );
  NAND2_X1 U12332 ( .A1(n11197), .A2(n10552), .ZN(n10553) );
  AOI21_X1 U12333 ( .B1(n15741), .B2(n10585), .A(n10553), .ZN(n10569) );
  INV_X1 U12334 ( .A(n15064), .ZN(n13906) );
  INV_X1 U12335 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10555) );
  MUX2_X1 U12336 ( .A(n10555), .B(P2_REG2_REG_1__SCAN_IN), .S(n15652), .Z(
        n15655) );
  AND2_X1 U12337 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n15656) );
  NAND2_X1 U12338 ( .A1(n15655), .A2(n15656), .ZN(n15654) );
  NAND2_X1 U12339 ( .A1(n8023), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n14701) );
  NAND2_X1 U12340 ( .A1(n15654), .A2(n14701), .ZN(n10557) );
  INV_X1 U12341 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n14699) );
  MUX2_X1 U12342 ( .A(n14699), .B(P2_REG2_REG_2__SCAN_IN), .S(n14698), .Z(
        n10556) );
  NAND2_X1 U12343 ( .A1(n10557), .A2(n10556), .ZN(n14717) );
  NAND2_X1 U12344 ( .A1(n10558), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n14716) );
  NAND2_X1 U12345 ( .A1(n14717), .A2(n14716), .ZN(n10561) );
  INV_X1 U12346 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10559) );
  MUX2_X1 U12347 ( .A(n10559), .B(P2_REG2_REG_3__SCAN_IN), .S(n14714), .Z(
        n10560) );
  NAND2_X1 U12348 ( .A1(n10561), .A2(n10560), .ZN(n14719) );
  NAND2_X1 U12349 ( .A1(n10562), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10565) );
  NAND2_X1 U12350 ( .A1(n14719), .A2(n10565), .ZN(n10564) );
  INV_X1 U12351 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11455) );
  MUX2_X1 U12352 ( .A(n11455), .B(P2_REG2_REG_4__SCAN_IN), .S(n11047), .Z(
        n10563) );
  NAND2_X1 U12353 ( .A1(n10564), .A2(n10563), .ZN(n10592) );
  MUX2_X1 U12354 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n11455), .S(n11047), .Z(
        n10566) );
  NAND3_X1 U12355 ( .A1(n10566), .A2(n14719), .A3(n10565), .ZN(n10567) );
  NAND3_X1 U12356 ( .A1(n15718), .A2(n10592), .A3(n10567), .ZN(n10568) );
  OAI211_X1 U12357 ( .C1(n15749), .C2(n7927), .A(n10569), .B(n10568), .ZN(
        P2_U3218) );
  INV_X1 U12358 ( .A(P3_DATAO_REG_4__SCAN_IN), .ZN(n10571) );
  NAND2_X1 U12359 ( .A1(n11806), .A2(P3_U3897), .ZN(n10570) );
  OAI21_X1 U12360 ( .B1(P3_U3897), .B2(n10571), .A(n10570), .ZN(P3_U3495) );
  OAI22_X1 U12361 ( .A1(n11074), .A2(n10669), .B1(n10876), .B2(n13594), .ZN(
        n10572) );
  XNOR2_X1 U12362 ( .A(n10572), .B(n13258), .ZN(n10576) );
  NAND2_X1 U12363 ( .A1(n11236), .A2(n13265), .ZN(n10573) );
  NAND2_X1 U12364 ( .A1(n10576), .A2(n10575), .ZN(n10666) );
  OAI21_X1 U12365 ( .B1(n10576), .B2(n10575), .A(n10666), .ZN(n10579) );
  AOI21_X1 U12366 ( .B1(n10579), .B2(n10580), .A(n10668), .ZN(n10583) );
  AOI22_X1 U12367 ( .A1(n16351), .A2(n15194), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n10675), .ZN(n10582) );
  NOR2_X1 U12368 ( .A1(n15132), .A2(n15406), .ZN(n16349) );
  AOI22_X1 U12369 ( .A1(n11236), .A2(n15173), .B1(n16349), .B2(n15197), .ZN(
        n10581) );
  OAI211_X1 U12370 ( .C1(n10583), .C2(n15175), .A(n10582), .B(n10581), .ZN(
        P1_U3222) );
  INV_X1 U12371 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10599) );
  NAND2_X1 U12372 ( .A1(n10585), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10587) );
  INV_X1 U12373 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n11402) );
  MUX2_X1 U12374 ( .A(n11402), .B(P2_REG1_REG_5__SCAN_IN), .S(n11132), .Z(
        n10586) );
  AOI21_X1 U12375 ( .B1(n10588), .B2(n10587), .A(n10586), .ZN(n10711) );
  INV_X1 U12376 ( .A(n10711), .ZN(n10590) );
  NAND3_X1 U12377 ( .A1(n10588), .A2(n10587), .A3(n10586), .ZN(n10589) );
  NAND3_X1 U12378 ( .A1(n10590), .A2(n15743), .A3(n10589), .ZN(n10598) );
  NAND2_X1 U12379 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n11146) );
  OR2_X1 U12380 ( .A1(n11047), .A2(n11455), .ZN(n10591) );
  NAND2_X1 U12381 ( .A1(n10592), .A2(n10591), .ZN(n10594) );
  INV_X1 U12382 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11445) );
  MUX2_X1 U12383 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n11445), .S(n11132), .Z(
        n10593) );
  NAND2_X1 U12384 ( .A1(n10594), .A2(n10593), .ZN(n10698) );
  OAI211_X1 U12385 ( .C1(n10594), .C2(n10593), .A(n15718), .B(n10698), .ZN(
        n10595) );
  NAND2_X1 U12386 ( .A1(n11146), .A2(n10595), .ZN(n10596) );
  AOI21_X1 U12387 ( .B1(n15741), .B2(n11132), .A(n10596), .ZN(n10597) );
  OAI211_X1 U12388 ( .C1(n15749), .C2(n10599), .A(n10598), .B(n10597), .ZN(
        P2_U3219) );
  OAI222_X1 U12389 ( .A1(P3_U3151), .A2(n14072), .B1(n13926), .B2(n12971), 
        .C1(n13924), .C2(n10600), .ZN(P3_U3282) );
  INV_X1 U12390 ( .A(P3_DATAO_REG_11__SCAN_IN), .ZN(n10602) );
  NAND2_X1 U12391 ( .A1(n12322), .A2(P3_U3897), .ZN(n10601) );
  OAI21_X1 U12392 ( .B1(P3_U3897), .B2(n10602), .A(n10601), .ZN(P3_U3502) );
  INV_X1 U12393 ( .A(P3_DATAO_REG_5__SCAN_IN), .ZN(n10604) );
  NAND2_X1 U12394 ( .A1(n11575), .A2(P3_U3897), .ZN(n10603) );
  OAI21_X1 U12395 ( .B1(P3_U3897), .B2(n10604), .A(n10603), .ZN(P3_U3496) );
  XOR2_X1 U12396 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10680), .Z(n10609) );
  INV_X1 U12397 ( .A(n10972), .ZN(n10622) );
  INV_X1 U12398 ( .A(n10618), .ZN(n10639) );
  INV_X1 U12399 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10605) );
  XNOR2_X1 U12400 ( .A(n10618), .B(n10605), .ZN(n10635) );
  NOR3_X1 U12401 ( .A1(n10635), .A2(n15751), .A3(n10606), .ZN(n10634) );
  AOI21_X1 U12402 ( .B1(n10639), .B2(P1_REG1_REG_1__SCAN_IN), .A(n10634), .ZN(
        n10970) );
  XOR2_X1 U12403 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10972), .Z(n10969) );
  NOR2_X1 U12404 ( .A1(n10970), .A2(n10969), .ZN(n10968) );
  XNOR2_X1 U12405 ( .A(n10623), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n10781) );
  INV_X1 U12406 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10607) );
  MUX2_X1 U12407 ( .A(n10607), .B(P1_REG1_REG_4__SCAN_IN), .S(n10817), .Z(
        n10815) );
  AOI21_X1 U12408 ( .B1(n10817), .B2(P1_REG1_REG_4__SCAN_IN), .A(n10814), .ZN(
        n10608) );
  OAI21_X1 U12409 ( .B1(n10609), .B2(n10608), .A(n10679), .ZN(n10615) );
  NAND2_X1 U12410 ( .A1(n10611), .A2(n10610), .ZN(n15759) );
  NOR2_X1 U12411 ( .A1(n15759), .A2(n10804), .ZN(n15778) );
  AND2_X1 U12412 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10612) );
  AOI21_X1 U12413 ( .B1(n15757), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n10612), .ZN(
        n10613) );
  OAI21_X1 U12414 ( .B1(n15765), .B2(n10685), .A(n10613), .ZN(n10614) );
  AOI21_X1 U12415 ( .B1(n10615), .B2(n15776), .A(n10614), .ZN(n10631) );
  NOR2_X1 U12416 ( .A1(n15759), .A2(n15594), .ZN(n15237) );
  INV_X1 U12417 ( .A(n15237), .ZN(n10616) );
  INV_X1 U12418 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10617) );
  MUX2_X1 U12419 ( .A(n10617), .B(P1_REG2_REG_2__SCAN_IN), .S(n10972), .Z(
        n10621) );
  INV_X1 U12420 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10619) );
  MUX2_X1 U12421 ( .A(n10619), .B(P1_REG2_REG_1__SCAN_IN), .S(n10618), .Z(
        n10641) );
  AND2_X1 U12422 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n10642) );
  NAND2_X1 U12423 ( .A1(n10641), .A2(n10642), .ZN(n10640) );
  NAND2_X1 U12424 ( .A1(n10639), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10620) );
  NAND2_X1 U12425 ( .A1(n10640), .A2(n10620), .ZN(n10963) );
  NAND2_X1 U12426 ( .A1(n10621), .A2(n10963), .ZN(n10964) );
  NAND2_X1 U12427 ( .A1(n10622), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n10778) );
  INV_X1 U12428 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n16074) );
  MUX2_X1 U12429 ( .A(n16074), .B(P1_REG2_REG_3__SCAN_IN), .S(n10623), .Z(
        n10777) );
  AOI21_X1 U12430 ( .B1(n10964), .B2(n10778), .A(n10777), .ZN(n10811) );
  NOR2_X1 U12431 ( .A1(n10785), .A2(n16074), .ZN(n10810) );
  INV_X1 U12432 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10624) );
  MUX2_X1 U12433 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10624), .S(n10817), .Z(
        n10809) );
  OAI21_X1 U12434 ( .B1(n10811), .B2(n10810), .A(n10809), .ZN(n10808) );
  NAND2_X1 U12435 ( .A1(n10817), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10627) );
  INV_X1 U12436 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10625) );
  MUX2_X1 U12437 ( .A(n10625), .B(P1_REG2_REG_5__SCAN_IN), .S(n10680), .Z(
        n10626) );
  AOI21_X1 U12438 ( .B1(n10808), .B2(n10627), .A(n10626), .ZN(n10795) );
  INV_X1 U12439 ( .A(n10795), .ZN(n10629) );
  NAND3_X1 U12440 ( .A1(n10808), .A2(n10627), .A3(n10626), .ZN(n10628) );
  NAND3_X1 U12441 ( .A1(n15780), .A2(n10629), .A3(n10628), .ZN(n10630) );
  NAND2_X1 U12442 ( .A1(n10631), .A2(n10630), .ZN(P1_U3248) );
  INV_X1 U12443 ( .A(n15757), .ZN(n15784) );
  INV_X1 U12444 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10632) );
  OAI22_X1 U12445 ( .A1(n15784), .A2(n10633), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10632), .ZN(n10638) );
  NAND2_X1 U12446 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n10636) );
  AOI211_X1 U12447 ( .C1(n10636), .C2(n10635), .A(n10634), .B(n15240), .ZN(
        n10637) );
  AOI211_X1 U12448 ( .C1(n15778), .C2(n10639), .A(n10638), .B(n10637), .ZN(
        n10644) );
  OAI211_X1 U12449 ( .C1(n10642), .C2(n10641), .A(n15780), .B(n10640), .ZN(
        n10643) );
  NAND2_X1 U12450 ( .A1(n10644), .A2(n10643), .ZN(P1_U3244) );
  AND2_X1 U12451 ( .A1(n10645), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U12452 ( .A1(n10645), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U12453 ( .A1(n10645), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U12454 ( .A1(n10645), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U12455 ( .A1(n10645), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U12456 ( .A1(n10645), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U12457 ( .A1(n10645), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U12458 ( .A1(n10645), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U12459 ( .A1(n10645), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U12460 ( .A1(n10645), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U12461 ( .A1(n10645), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U12462 ( .A1(n10645), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U12463 ( .A1(n10645), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U12464 ( .A1(n10645), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  INV_X1 U12465 ( .A(n12101), .ZN(n10654) );
  INV_X1 U12466 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n10647) );
  NAND4_X1 U12467 ( .A1(n10649), .A2(n10648), .A3(n10647), .A4(n10646), .ZN(
        n10650) );
  OAI21_X1 U12468 ( .B1(n10651), .B2(n10650), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n10652) );
  XNOR2_X1 U12469 ( .A(n10652), .B(P2_IR_REG_12__SCAN_IN), .ZN(n12243) );
  INV_X1 U12470 ( .A(n12243), .ZN(n11354) );
  OAI222_X1 U12471 ( .A1(n13255), .A2(n10653), .B1(n15061), .B2(n10654), .C1(
        n11354), .C2(P2_U3088), .ZN(P2_U3315) );
  INV_X1 U12472 ( .A(n15779), .ZN(n11707) );
  OAI222_X1 U12473 ( .A1(n15597), .A2(n10655), .B1(n15604), .B2(n10654), .C1(
        n11707), .C2(P1_U3086), .ZN(P1_U3343) );
  AND2_X1 U12474 ( .A1(n10657), .A2(n10656), .ZN(n11361) );
  NAND2_X1 U12475 ( .A1(n11359), .A2(n15647), .ZN(n15641) );
  NOR2_X1 U12476 ( .A1(n15641), .A2(n10658), .ZN(n10659) );
  AND2_X1 U12477 ( .A1(n11361), .A2(n10659), .ZN(n10978) );
  OAI21_X1 U12478 ( .B1(n13669), .B2(n11702), .A(n10767), .ZN(n13621) );
  NAND2_X1 U12479 ( .A1(n8074), .A2(n13662), .ZN(n10660) );
  NAND2_X1 U12480 ( .A1(n7420), .A2(n7415), .ZN(n13861) );
  INV_X1 U12481 ( .A(n14691), .ZN(n10944) );
  OAI22_X1 U12482 ( .A1(n13621), .A2(n14821), .B1(n10944), .B2(n14916), .ZN(
        n11697) );
  AND2_X2 U12483 ( .A1(n13665), .A2(n13912), .ZN(n13663) );
  OAI22_X1 U12484 ( .A1(n13621), .A2(n14998), .B1(n10663), .B2(n13667), .ZN(
        n10664) );
  OR2_X1 U12485 ( .A1(n11697), .A2(n10664), .ZN(n10979) );
  NAND2_X1 U12486 ( .A1(n16293), .A2(n10979), .ZN(n10665) );
  OAI21_X1 U12487 ( .B1(n16293), .B2(n10546), .A(n10665), .ZN(P2_U3499) );
  INV_X1 U12488 ( .A(n10666), .ZN(n10667) );
  INV_X1 U12489 ( .A(n7430), .ZN(n11100) );
  OAI22_X1 U12490 ( .A1(n11106), .A2(n13588), .B1(n11100), .B2(n13594), .ZN(
        n10670) );
  XNOR2_X1 U12491 ( .A(n10670), .B(n11815), .ZN(n10946) );
  NAND2_X1 U12492 ( .A1(n13265), .A2(n7430), .ZN(n10671) );
  NAND2_X1 U12493 ( .A1(n10672), .A2(n10671), .ZN(n10945) );
  XNOR2_X1 U12494 ( .A(n10946), .B(n10945), .ZN(n10673) );
  AOI21_X1 U12495 ( .B1(n10674), .B2(n10673), .A(n10949), .ZN(n10678) );
  AOI22_X1 U12496 ( .A1(n16351), .A2(n15193), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n10675), .ZN(n10677) );
  AOI22_X1 U12497 ( .A1(n7430), .A2(n15173), .B1(n16349), .B2(n15195), .ZN(
        n10676) );
  OAI211_X1 U12498 ( .C1(n10678), .C2(n15175), .A(n10677), .B(n10676), .ZN(
        P1_U3237) );
  INV_X1 U12499 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10681) );
  MUX2_X1 U12500 ( .A(n10681), .B(P1_REG1_REG_6__SCAN_IN), .S(n10687), .Z(
        n10791) );
  INV_X1 U12501 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10682) );
  MUX2_X1 U12502 ( .A(n10682), .B(P1_REG1_REG_7__SCAN_IN), .S(n10756), .Z(
        n10683) );
  NOR2_X1 U12503 ( .A1(n10684), .A2(n10683), .ZN(n10755) );
  AOI211_X1 U12504 ( .C1(n10684), .C2(n10683), .A(n15240), .B(n10755), .ZN(
        n10696) );
  NOR2_X1 U12505 ( .A1(n10685), .A2(n10625), .ZN(n10794) );
  INV_X1 U12506 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10686) );
  MUX2_X1 U12507 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10686), .S(n10687), .Z(
        n10793) );
  OAI21_X1 U12508 ( .B1(n10795), .B2(n10794), .A(n10793), .ZN(n10792) );
  NAND2_X1 U12509 ( .A1(n10687), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10689) );
  INV_X1 U12510 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10749) );
  MUX2_X1 U12511 ( .A(n10749), .B(P1_REG2_REG_7__SCAN_IN), .S(n10756), .Z(
        n10688) );
  AOI21_X1 U12512 ( .B1(n10792), .B2(n10689), .A(n10688), .ZN(n10926) );
  INV_X1 U12513 ( .A(n10926), .ZN(n10691) );
  NAND3_X1 U12514 ( .A1(n10792), .A2(n10689), .A3(n10688), .ZN(n10690) );
  NAND3_X1 U12515 ( .A1(n10691), .A2(n15780), .A3(n10690), .ZN(n10694) );
  NOR2_X1 U12516 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8732), .ZN(n10692) );
  AOI21_X1 U12517 ( .B1(n15757), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n10692), .ZN(
        n10693) );
  OAI211_X1 U12518 ( .C1(n15765), .C2(n10750), .A(n10694), .B(n10693), .ZN(
        n10695) );
  OR2_X1 U12519 ( .A1(n10696), .A2(n10695), .ZN(P1_U3250) );
  NAND2_X1 U12520 ( .A1(n11132), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10697) );
  NAND2_X1 U12521 ( .A1(n10698), .A2(n10697), .ZN(n15671) );
  INV_X1 U12522 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10699) );
  MUX2_X1 U12523 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10699), .S(n11540), .Z(
        n15670) );
  NAND2_X1 U12524 ( .A1(n15671), .A2(n15670), .ZN(n15669) );
  NAND2_X1 U12525 ( .A1(n11540), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n10902) );
  NAND2_X1 U12526 ( .A1(n15669), .A2(n10902), .ZN(n10702) );
  INV_X1 U12527 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10700) );
  MUX2_X1 U12528 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10700), .S(n11544), .Z(
        n10701) );
  NAND2_X1 U12529 ( .A1(n10702), .A2(n10701), .ZN(n10908) );
  NAND2_X1 U12530 ( .A1(n11544), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10907) );
  NAND2_X1 U12531 ( .A1(n10908), .A2(n10907), .ZN(n10705) );
  INV_X1 U12532 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10703) );
  MUX2_X1 U12533 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10703), .S(n11672), .Z(
        n10704) );
  NAND2_X1 U12534 ( .A1(n10705), .A2(n10704), .ZN(n10910) );
  NAND2_X1 U12535 ( .A1(n11672), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10706) );
  NAND2_X1 U12536 ( .A1(n10910), .A2(n10706), .ZN(n10710) );
  INV_X1 U12537 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10707) );
  MUX2_X1 U12538 ( .A(n10707), .B(P2_REG2_REG_9__SCAN_IN), .S(n11855), .Z(
        n10709) );
  OR2_X1 U12539 ( .A1(n10710), .A2(n10709), .ZN(n10993) );
  INV_X1 U12540 ( .A(n10993), .ZN(n10708) );
  AOI21_X1 U12541 ( .B1(n10710), .B2(n10709), .A(n10708), .ZN(n10718) );
  AOI21_X1 U12542 ( .B1(P2_REG1_REG_5__SCAN_IN), .B2(n11132), .A(n10711), .ZN(
        n15674) );
  INV_X1 U12543 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n16128) );
  MUX2_X1 U12544 ( .A(n16128), .B(P2_REG1_REG_6__SCAN_IN), .S(n11540), .Z(
        n15673) );
  NOR2_X1 U12545 ( .A1(n15674), .A2(n15673), .ZN(n15672) );
  AOI21_X1 U12546 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n11540), .A(n15672), .ZN(
        n10897) );
  INV_X1 U12547 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n16146) );
  MUX2_X1 U12548 ( .A(n16146), .B(P2_REG1_REG_7__SCAN_IN), .S(n11544), .Z(
        n10896) );
  NOR2_X1 U12549 ( .A1(n10897), .A2(n10896), .ZN(n10895) );
  AOI21_X1 U12550 ( .B1(n11544), .B2(P2_REG1_REG_7__SCAN_IN), .A(n10895), .ZN(
        n10913) );
  INV_X1 U12551 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n16194) );
  MUX2_X1 U12552 ( .A(n16194), .B(P2_REG1_REG_8__SCAN_IN), .S(n11672), .Z(
        n10912) );
  NOR2_X1 U12553 ( .A1(n10913), .A2(n10912), .ZN(n10911) );
  AOI21_X1 U12554 ( .B1(n11672), .B2(P2_REG1_REG_8__SCAN_IN), .A(n10911), .ZN(
        n10713) );
  INV_X1 U12555 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n16211) );
  MUX2_X1 U12556 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n16211), .S(n11855), .Z(
        n10712) );
  NOR2_X1 U12557 ( .A1(n10713), .A2(n10712), .ZN(n10714) );
  AND2_X1 U12558 ( .A1(n10713), .A2(n10712), .ZN(n10985) );
  OAI21_X1 U12559 ( .B1(n10714), .B2(n10985), .A(n15743), .ZN(n10717) );
  AND2_X1 U12560 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n11914) );
  INV_X1 U12561 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n15863) );
  NOR2_X1 U12562 ( .A1(n15749), .A2(n15863), .ZN(n10715) );
  AOI211_X1 U12563 ( .C1(n11855), .C2(n15741), .A(n11914), .B(n10715), .ZN(
        n10716) );
  OAI211_X1 U12564 ( .C1(n10718), .C2(n15736), .A(n10717), .B(n10716), .ZN(
        P2_U3223) );
  INV_X1 U12565 ( .A(n12183), .ZN(n10726) );
  NOR2_X1 U12566 ( .A1(n10720), .A2(n10719), .ZN(n10721) );
  NAND2_X1 U12567 ( .A1(n10722), .A2(n10721), .ZN(n11771) );
  NAND2_X1 U12568 ( .A1(n11771), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10723) );
  MUX2_X1 U12569 ( .A(P2_IR_REG_31__SCAN_IN), .B(n10723), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n10724) );
  INV_X1 U12570 ( .A(n15717), .ZN(n15725) );
  OAI222_X1 U12571 ( .A1(n13255), .A2(n10725), .B1(n15061), .B2(n10726), .C1(
        n15725), .C2(P2_U3088), .ZN(P2_U3314) );
  INV_X1 U12572 ( .A(n12081), .ZN(n12086) );
  OAI222_X1 U12573 ( .A1(n15597), .A2(n10727), .B1(n15604), .B2(n10726), .C1(
        n12086), .C2(P1_U3086), .ZN(P1_U3342) );
  OAI222_X1 U12574 ( .A1(P3_U3151), .A2(n10729), .B1(n13926), .B2(n7846), .C1(
        n13924), .C2(n10728), .ZN(P3_U3281) );
  AOI22_X1 U12575 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n15718), .B1(n15743), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n10733) );
  INV_X1 U12576 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10731) );
  NOR2_X1 U12577 ( .A1(n15728), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n10730) );
  AOI211_X1 U12578 ( .C1(n15718), .C2(n10731), .A(n15741), .B(n10730), .ZN(
        n10732) );
  MUX2_X1 U12579 ( .A(n10733), .B(n10732), .S(P2_IR_REG_0__SCAN_IN), .Z(n10735) );
  AOI22_X1 U12580 ( .A1(n15683), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n10734) );
  NAND2_X1 U12581 ( .A1(n10735), .A2(n10734), .ZN(P2_U3214) );
  INV_X1 U12582 ( .A(n10767), .ZN(n10736) );
  NAND2_X1 U12583 ( .A1(n7422), .A2(n14626), .ZN(n11055) );
  NAND2_X1 U12584 ( .A1(n7423), .A2(n11367), .ZN(n10737) );
  AND2_X1 U12585 ( .A1(n11055), .A2(n10737), .ZN(n13623) );
  XNOR2_X1 U12586 ( .A(n11038), .B(n11037), .ZN(n11370) );
  INV_X1 U12587 ( .A(n11370), .ZN(n10747) );
  NAND2_X1 U12588 ( .A1(n10944), .A2(n7432), .ZN(n10739) );
  NAND2_X1 U12589 ( .A1(n10768), .A2(n10739), .ZN(n10738) );
  NAND2_X1 U12590 ( .A1(n10738), .A2(n13623), .ZN(n11056) );
  NAND3_X1 U12591 ( .A1(n11037), .A2(n10768), .A3(n10739), .ZN(n10740) );
  AND2_X1 U12592 ( .A1(n11056), .A2(n10740), .ZN(n10743) );
  NAND2_X1 U12593 ( .A1(n11370), .A2(n14902), .ZN(n10742) );
  AOI22_X1 U12594 ( .A1(n14883), .A2(n7580), .B1(n14689), .B2(n14885), .ZN(
        n10741) );
  OAI211_X1 U12595 ( .C1(n14821), .C2(n10743), .A(n10742), .B(n10741), .ZN(
        n11363) );
  INV_X1 U12596 ( .A(n11363), .ZN(n10746) );
  NAND2_X1 U12597 ( .A1(n7431), .A2(n13667), .ZN(n10773) );
  NAND2_X1 U12598 ( .A1(n10773), .A2(n14626), .ZN(n10744) );
  AND2_X1 U12599 ( .A1(n11209), .A2(n10744), .ZN(n11365) );
  AOI22_X1 U12600 ( .A1(n11365), .A2(n15027), .B1(n15026), .B2(n14626), .ZN(
        n10745) );
  OAI211_X1 U12601 ( .C1(n10747), .C2(n15031), .A(n10746), .B(n10745), .ZN(
        n10982) );
  NAND2_X1 U12602 ( .A1(n10982), .A2(n16293), .ZN(n10748) );
  OAI21_X1 U12603 ( .B1(n16293), .B2(n10547), .A(n10748), .ZN(P2_U3501) );
  NOR2_X1 U12604 ( .A1(n10750), .A2(n10749), .ZN(n10925) );
  INV_X1 U12605 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n16180) );
  MUX2_X1 U12606 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n16180), .S(n10758), .Z(
        n10924) );
  OAI21_X1 U12607 ( .B1(n10926), .B2(n10925), .A(n10924), .ZN(n10923) );
  NAND2_X1 U12608 ( .A1(n10758), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10752) );
  INV_X1 U12609 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n11936) );
  MUX2_X1 U12610 ( .A(n11936), .B(P1_REG2_REG_9__SCAN_IN), .S(n11175), .Z(
        n10751) );
  AOI21_X1 U12611 ( .B1(n10923), .B2(n10752), .A(n10751), .ZN(n11185) );
  NAND3_X1 U12612 ( .A1(n10923), .A2(n10752), .A3(n10751), .ZN(n10753) );
  NAND2_X1 U12613 ( .A1(n10753), .A2(n15780), .ZN(n10766) );
  INV_X1 U12614 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10754) );
  MUX2_X1 U12615 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10754), .S(n11175), .Z(
        n10760) );
  INV_X1 U12616 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10757) );
  MUX2_X1 U12617 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10757), .S(n10758), .Z(
        n10921) );
  OAI21_X1 U12618 ( .B1(n10760), .B2(n10759), .A(n11174), .ZN(n10761) );
  NAND2_X1 U12619 ( .A1(n10761), .A2(n15776), .ZN(n10765) );
  INV_X1 U12620 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n11986) );
  NOR2_X1 U12621 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11986), .ZN(n10763) );
  NOR2_X1 U12622 ( .A1(n15765), .A2(n11179), .ZN(n10762) );
  AOI211_X1 U12623 ( .C1(n15757), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n10763), .B(
        n10762), .ZN(n10764) );
  OAI211_X1 U12624 ( .C1(n11185), .C2(n10766), .A(n10765), .B(n10764), .ZN(
        P1_U3252) );
  XNOR2_X1 U12625 ( .A(n13622), .B(n10767), .ZN(n11406) );
  OAI21_X1 U12626 ( .B1(n13664), .B2(n13622), .A(n10768), .ZN(n10771) );
  INV_X1 U12627 ( .A(n13669), .ZN(n10939) );
  INV_X1 U12628 ( .A(n14883), .ZN(n14914) );
  OAI22_X1 U12629 ( .A1(n10939), .A2(n14914), .B1(n7422), .B2(n14916), .ZN(
        n10770) );
  NOR2_X1 U12630 ( .A1(n11406), .A2(n10661), .ZN(n10769) );
  AOI211_X1 U12631 ( .C1(n14924), .C2(n10771), .A(n10770), .B(n10769), .ZN(
        n11411) );
  NAND2_X1 U12632 ( .A1(n11702), .A2(n7432), .ZN(n10772) );
  AND2_X1 U12633 ( .A1(n10773), .A2(n10772), .ZN(n11409) );
  AOI22_X1 U12634 ( .A1(n11409), .A2(n15027), .B1(n15026), .B2(n7432), .ZN(
        n10774) );
  OAI211_X1 U12635 ( .C1(n15031), .C2(n11406), .A(n11411), .B(n10774), .ZN(
        n11003) );
  NAND2_X1 U12636 ( .A1(n11003), .A2(n16293), .ZN(n10775) );
  OAI21_X1 U12637 ( .B1(n16293), .B2(n10776), .A(n10775), .ZN(P2_U3500) );
  INV_X1 U12638 ( .A(n15780), .ZN(n15767) );
  AND3_X1 U12639 ( .A1(n10964), .A2(n10778), .A3(n10777), .ZN(n10779) );
  NOR3_X1 U12640 ( .A1(n15767), .A2(n10811), .A3(n10779), .ZN(n10788) );
  AOI211_X1 U12641 ( .C1(n10782), .C2(n10781), .A(n10780), .B(n15240), .ZN(
        n10787) );
  NOR2_X1 U12642 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10958), .ZN(n10783) );
  AOI21_X1 U12643 ( .B1(n15757), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n10783), .ZN(
        n10784) );
  OAI21_X1 U12644 ( .B1(n15765), .B2(n10785), .A(n10784), .ZN(n10786) );
  OR3_X1 U12645 ( .A1(n10788), .A2(n10787), .A3(n10786), .ZN(P1_U3246) );
  AOI211_X1 U12646 ( .C1(n10791), .C2(n10790), .A(n15240), .B(n10789), .ZN(
        n10802) );
  INV_X1 U12647 ( .A(n10792), .ZN(n10797) );
  NOR3_X1 U12648 ( .A1(n10795), .A2(n10794), .A3(n10793), .ZN(n10796) );
  NOR3_X1 U12649 ( .A1(n15767), .A2(n10797), .A3(n10796), .ZN(n10801) );
  NAND2_X1 U12650 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n11473) );
  NAND2_X1 U12651 ( .A1(n15757), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n10798) );
  OAI211_X1 U12652 ( .C1(n15765), .C2(n10799), .A(n11473), .B(n10798), .ZN(
        n10800) );
  OR3_X1 U12653 ( .A1(n10802), .A2(n10801), .A3(n10800), .ZN(P1_U3249) );
  INV_X1 U12654 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n11076) );
  NAND2_X1 U12655 ( .A1(n15750), .A2(n11076), .ZN(n10803) );
  NAND2_X1 U12656 ( .A1(n10804), .A2(n10803), .ZN(n15752) );
  NOR3_X1 U12657 ( .A1(n10805), .A2(n15750), .A3(n15752), .ZN(n10807) );
  NOR2_X1 U12658 ( .A1(n15752), .A2(n15594), .ZN(n10806) );
  MUX2_X1 U12659 ( .A(n15752), .B(n10806), .S(P1_IR_REG_0__SCAN_IN), .Z(n15756) );
  NOR3_X1 U12660 ( .A1(n10807), .A2(n15196), .A3(n15756), .ZN(n10976) );
  INV_X1 U12661 ( .A(n10808), .ZN(n10813) );
  NOR3_X1 U12662 ( .A1(n10811), .A2(n10810), .A3(n10809), .ZN(n10812) );
  NOR3_X1 U12663 ( .A1(n15767), .A2(n10813), .A3(n10812), .ZN(n10821) );
  AOI211_X1 U12664 ( .C1(n10816), .C2(n10815), .A(n15240), .B(n10814), .ZN(
        n10820) );
  NAND2_X1 U12665 ( .A1(n15778), .A2(n10817), .ZN(n10818) );
  NAND2_X1 U12666 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n11339) );
  OAI211_X1 U12667 ( .C1(n7609), .C2(n15784), .A(n10818), .B(n11339), .ZN(
        n10819) );
  OR4_X1 U12668 ( .A1(n10976), .A2(n10821), .A3(n10820), .A4(n10819), .ZN(
        P1_U3247) );
  INV_X1 U12669 ( .A(n16009), .ZN(n15973) );
  OAI21_X1 U12670 ( .B1(n10824), .B2(n10823), .A(n10822), .ZN(n10833) );
  OAI21_X1 U12671 ( .B1(P3_REG1_REG_2__SCAN_IN), .B2(n10842), .A(n10825), .ZN(
        n10828) );
  INV_X1 U12672 ( .A(n10825), .ZN(n10827) );
  AOI22_X1 U12673 ( .A1(n10829), .A2(n10828), .B1(n10827), .B2(n10826), .ZN(
        n10831) );
  AOI22_X1 U12674 ( .A1(n15646), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10830) );
  OAI21_X1 U12675 ( .B1(n10831), .B2(n16013), .A(n10830), .ZN(n10832) );
  AOI21_X1 U12676 ( .B1(n15973), .B2(n10833), .A(n10832), .ZN(n10841) );
  INV_X1 U12677 ( .A(n10834), .ZN(n11086) );
  INV_X1 U12678 ( .A(n10835), .ZN(n10837) );
  NOR3_X1 U12679 ( .A1(n11086), .A2(n10837), .A3(n10836), .ZN(n10839) );
  INV_X1 U12680 ( .A(n11166), .ZN(n10838) );
  OAI21_X1 U12681 ( .B1(n10839), .B2(n10838), .A(n16017), .ZN(n10840) );
  OAI211_X1 U12682 ( .C1(n15997), .C2(n10842), .A(n10841), .B(n10840), .ZN(
        P3_U3184) );
  INV_X1 U12683 ( .A(n11168), .ZN(n10846) );
  INV_X1 U12684 ( .A(n10843), .ZN(n10845) );
  NOR3_X1 U12685 ( .A1(n10846), .A2(n10845), .A3(n10844), .ZN(n10849) );
  INV_X1 U12686 ( .A(n10847), .ZN(n10848) );
  OAI21_X1 U12687 ( .B1(n10849), .B2(n10848), .A(n16017), .ZN(n10866) );
  INV_X1 U12688 ( .A(n10850), .ZN(n10852) );
  NAND3_X1 U12689 ( .A1(n11153), .A2(n10852), .A3(n10851), .ZN(n10853) );
  AOI21_X1 U12690 ( .B1(n10854), .B2(n10853), .A(n16009), .ZN(n10864) );
  INV_X1 U12691 ( .A(n10855), .ZN(n10857) );
  NAND3_X1 U12692 ( .A1(n11157), .A2(n10857), .A3(n10856), .ZN(n10858) );
  AOI21_X1 U12693 ( .B1(n10859), .B2(n10858), .A(n16013), .ZN(n10863) );
  INV_X1 U12694 ( .A(n15646), .ZN(n16027) );
  INV_X1 U12695 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n10860) );
  NOR2_X1 U12696 ( .A1(n16027), .A2(n10860), .ZN(n10862) );
  NAND2_X1 U12697 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_U3151), .ZN(n11726) );
  INV_X1 U12698 ( .A(n11726), .ZN(n10861) );
  NOR4_X1 U12699 ( .A1(n10864), .A2(n10863), .A3(n10862), .A4(n10861), .ZN(
        n10865) );
  OAI211_X1 U12700 ( .C1(n15997), .C2(n10867), .A(n10866), .B(n10865), .ZN(
        P3_U3186) );
  AND2_X1 U12701 ( .A1(n10871), .A2(n11071), .ZN(n10892) );
  INV_X1 U12702 ( .A(n10891), .ZN(n11070) );
  AND2_X2 U12703 ( .A1(n10892), .A2(n11070), .ZN(n16345) );
  INV_X1 U12704 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10890) );
  INV_X1 U12705 ( .A(n10872), .ZN(n10873) );
  NAND2_X1 U12706 ( .A1(n10873), .A2(n12527), .ZN(n16135) );
  AND2_X1 U12707 ( .A1(n11080), .A2(n15197), .ZN(n10874) );
  NAND2_X1 U12708 ( .A1(n11007), .A2(n10875), .ZN(n11241) );
  NAND2_X1 U12709 ( .A1(n16032), .A2(n10876), .ZN(n11009) );
  OAI21_X1 U12710 ( .B1(n16032), .B2(n10876), .A(n11009), .ZN(n11238) );
  OAI22_X1 U12711 ( .A1(n11238), .A2(n16198), .B1(n10876), .B2(n16333), .ZN(
        n10888) );
  OR2_X1 U12712 ( .A1(n10878), .A2(n10877), .ZN(n10879) );
  NAND2_X1 U12713 ( .A1(n11295), .A2(n15244), .ZN(n16254) );
  INV_X1 U12714 ( .A(n16254), .ZN(n16160) );
  NAND2_X1 U12715 ( .A1(n11241), .A2(n16160), .ZN(n10887) );
  INV_X1 U12716 ( .A(n10880), .ZN(n11011) );
  NAND2_X1 U12717 ( .A1(n10881), .A2(n8224), .ZN(n10883) );
  NAND2_X1 U12718 ( .A1(n7429), .A2(n15606), .ZN(n10882) );
  NAND2_X1 U12719 ( .A1(n10884), .A2(n16330), .ZN(n10886) );
  AOI22_X1 U12720 ( .A1(n15194), .A2(n15457), .B1(n15455), .B2(n15197), .ZN(
        n10885) );
  NAND3_X1 U12721 ( .A1(n10887), .A2(n10886), .A3(n10885), .ZN(n11235) );
  AOI211_X1 U12722 ( .C1(n16257), .C2(n11241), .A(n10888), .B(n11235), .ZN(
        n10893) );
  OR2_X1 U12723 ( .A1(n10893), .A2(n16342), .ZN(n10889) );
  OAI21_X1 U12724 ( .B1(n16345), .B2(n10890), .A(n10889), .ZN(P1_U3462) );
  AND2_X2 U12725 ( .A1(n10892), .A2(n10891), .ZN(n16341) );
  OR2_X1 U12726 ( .A1(n10893), .A2(n16339), .ZN(n10894) );
  OAI21_X1 U12727 ( .B1(n16341), .B2(n10605), .A(n10894), .ZN(P1_U3529) );
  NAND2_X1 U12728 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n11606) );
  AOI211_X1 U12729 ( .C1(n10897), .C2(n10896), .A(n10895), .B(n15728), .ZN(
        n10898) );
  INV_X1 U12730 ( .A(n10898), .ZN(n10899) );
  NAND2_X1 U12731 ( .A1(n11606), .A2(n10899), .ZN(n10900) );
  AOI21_X1 U12732 ( .B1(n15741), .B2(n11544), .A(n10900), .ZN(n10905) );
  MUX2_X1 U12733 ( .A(n10700), .B(P2_REG2_REG_7__SCAN_IN), .S(n11544), .Z(
        n10901) );
  NAND3_X1 U12734 ( .A1(n15669), .A2(n10902), .A3(n10901), .ZN(n10903) );
  NAND3_X1 U12735 ( .A1(n15718), .A2(n10908), .A3(n10903), .ZN(n10904) );
  OAI211_X1 U12736 ( .C1(n15749), .C2(n7931), .A(n10905), .B(n10904), .ZN(
        P2_U3221) );
  INV_X1 U12737 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10919) );
  MUX2_X1 U12738 ( .A(n10703), .B(P2_REG2_REG_8__SCAN_IN), .S(n11672), .Z(
        n10906) );
  NAND3_X1 U12739 ( .A1(n10908), .A2(n10907), .A3(n10906), .ZN(n10909) );
  NAND3_X1 U12740 ( .A1(n10910), .A2(n15718), .A3(n10909), .ZN(n10918) );
  NAND2_X1 U12741 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n11745) );
  AOI211_X1 U12742 ( .C1(n10913), .C2(n10912), .A(n10911), .B(n15728), .ZN(
        n10914) );
  INV_X1 U12743 ( .A(n10914), .ZN(n10915) );
  NAND2_X1 U12744 ( .A1(n11745), .A2(n10915), .ZN(n10916) );
  AOI21_X1 U12745 ( .B1(n15741), .B2(n11672), .A(n10916), .ZN(n10917) );
  OAI211_X1 U12746 ( .C1(n15749), .C2(n10919), .A(n10918), .B(n10917), .ZN(
        P2_U3222) );
  OAI21_X1 U12747 ( .B1(n10922), .B2(n10921), .A(n10920), .ZN(n10933) );
  INV_X1 U12748 ( .A(n10923), .ZN(n10928) );
  NOR3_X1 U12749 ( .A1(n10926), .A2(n10925), .A3(n10924), .ZN(n10927) );
  NOR3_X1 U12750 ( .A1(n10928), .A2(n10927), .A3(n15767), .ZN(n10932) );
  NAND2_X1 U12751 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n11826) );
  NAND2_X1 U12752 ( .A1(n15757), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n10929) );
  OAI211_X1 U12753 ( .C1(n15765), .C2(n10930), .A(n11826), .B(n10929), .ZN(
        n10931) );
  AOI211_X1 U12754 ( .C1(n10933), .C2(n15776), .A(n10932), .B(n10931), .ZN(
        n10934) );
  INV_X1 U12755 ( .A(n10934), .ZN(P1_U3251) );
  OAI222_X1 U12756 ( .A1(P3_U3151), .A2(n14085), .B1(n13926), .B2(n10936), 
        .C1(n13924), .C2(n10935), .ZN(P3_U3280) );
  OR2_X1 U12757 ( .A1(n10937), .A2(P2_U3088), .ZN(n14625) );
  AOI22_X1 U12758 ( .A1(n14651), .A2(n11702), .B1(n14625), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n10943) );
  OAI21_X1 U12759 ( .B1(n10939), .B2(n10938), .A(n13667), .ZN(n10940) );
  NAND3_X1 U12760 ( .A1(n14658), .A2(n10941), .A3(n10940), .ZN(n10942) );
  OAI211_X1 U12761 ( .C1(n10944), .C2(n14663), .A(n10943), .B(n10942), .ZN(
        P2_U3204) );
  INV_X1 U12762 ( .A(n10945), .ZN(n10948) );
  INV_X1 U12763 ( .A(n10946), .ZN(n10947) );
  OAI22_X1 U12764 ( .A1(n11297), .A2(n13587), .B1(n16077), .B2(n13588), .ZN(
        n11270) );
  OAI22_X1 U12765 ( .A1(n11297), .A2(n13588), .B1(n16077), .B2(n13594), .ZN(
        n10950) );
  XNOR2_X1 U12766 ( .A(n10950), .B(n11815), .ZN(n11271) );
  XOR2_X1 U12767 ( .A(n11270), .B(n11271), .Z(n10951) );
  OAI211_X1 U12768 ( .C1(n10952), .C2(n10951), .A(n11275), .B(n16356), .ZN(
        n10962) );
  NOR2_X1 U12769 ( .A1(n10954), .A2(n10953), .ZN(n10955) );
  NAND2_X1 U12770 ( .A1(n10956), .A2(n10955), .ZN(n10957) );
  NAND2_X1 U12771 ( .A1(n10957), .A2(P1_STATE_REG_SCAN_IN), .ZN(n16361) );
  INV_X1 U12772 ( .A(n15192), .ZN(n11484) );
  OAI22_X1 U12773 ( .A1(n15170), .A2(n11484), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10958), .ZN(n10960) );
  INV_X1 U12774 ( .A(n16349), .ZN(n15159) );
  OAI22_X1 U12775 ( .A1(n16077), .A2(n16353), .B1(n15159), .B2(n11106), .ZN(
        n10959) );
  AOI211_X1 U12776 ( .C1(n15167), .C2(n10958), .A(n10960), .B(n10959), .ZN(
        n10961) );
  NAND2_X1 U12777 ( .A1(n10962), .A2(n10961), .ZN(P1_U3218) );
  INV_X1 U12778 ( .A(n10963), .ZN(n10967) );
  MUX2_X1 U12779 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10617), .S(n10972), .Z(
        n10966) );
  INV_X1 U12780 ( .A(n10964), .ZN(n10965) );
  AOI211_X1 U12781 ( .C1(n10967), .C2(n10966), .A(n10965), .B(n15767), .ZN(
        n10975) );
  AOI211_X1 U12782 ( .C1(n10970), .C2(n10969), .A(n10968), .B(n15240), .ZN(
        n10974) );
  AOI22_X1 U12783 ( .A1(n15757), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n10971) );
  OAI21_X1 U12784 ( .B1(n15765), .B2(n10972), .A(n10971), .ZN(n10973) );
  OR4_X1 U12785 ( .A1(n10976), .A2(n10975), .A3(n10974), .A4(n10973), .ZN(
        P1_U3245) );
  INV_X1 U12786 ( .A(n15648), .ZN(n10977) );
  INV_X1 U12787 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10981) );
  NAND2_X1 U12788 ( .A1(n7419), .A2(n10979), .ZN(n10980) );
  OAI21_X1 U12789 ( .B1(n7419), .B2(n10981), .A(n10980), .ZN(P2_U3430) );
  INV_X1 U12790 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10984) );
  NAND2_X1 U12791 ( .A1(n10982), .A2(n7419), .ZN(n10983) );
  OAI21_X1 U12792 ( .B1(n7419), .B2(n10984), .A(n10983), .ZN(P2_U3436) );
  AOI21_X1 U12793 ( .B1(n16211), .B2(n10986), .A(n10985), .ZN(n15746) );
  INV_X1 U12794 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10987) );
  MUX2_X1 U12795 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n10987), .S(n15742), .Z(
        n15745) );
  NAND2_X1 U12796 ( .A1(n15746), .A2(n15745), .ZN(n15744) );
  NAND2_X1 U12797 ( .A1(n15742), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10989) );
  INV_X1 U12798 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n12316) );
  MUX2_X1 U12799 ( .A(n12316), .B(P2_REG1_REG_11__SCAN_IN), .S(n12021), .Z(
        n10988) );
  AOI21_X1 U12800 ( .B1(n15744), .B2(n10989), .A(n10988), .ZN(n11350) );
  NAND3_X1 U12801 ( .A1(n15744), .A2(n10989), .A3(n10988), .ZN(n10990) );
  NAND2_X1 U12802 ( .A1(n10990), .A2(n15743), .ZN(n11002) );
  INV_X1 U12803 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n15881) );
  NAND2_X1 U12804 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n12301)
         );
  OAI21_X1 U12805 ( .B1(n15749), .B2(n15881), .A(n12301), .ZN(n10991) );
  AOI21_X1 U12806 ( .B1(n12021), .B2(n15741), .A(n10991), .ZN(n11001) );
  OR2_X1 U12807 ( .A1(n11855), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n10992) );
  NAND2_X1 U12808 ( .A1(n10993), .A2(n10992), .ZN(n15738) );
  INV_X1 U12809 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10994) );
  MUX2_X1 U12810 ( .A(n10994), .B(P2_REG2_REG_10__SCAN_IN), .S(n15742), .Z(
        n15737) );
  OR2_X1 U12811 ( .A1(n15738), .A2(n15737), .ZN(n15734) );
  NAND2_X1 U12812 ( .A1(n15742), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10995) );
  AND2_X1 U12813 ( .A1(n15734), .A2(n10995), .ZN(n10998) );
  INV_X1 U12814 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10996) );
  MUX2_X1 U12815 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n10996), .S(n12021), .Z(
        n10997) );
  NAND2_X1 U12816 ( .A1(n10998), .A2(n10997), .ZN(n11346) );
  OAI21_X1 U12817 ( .B1(n10998), .B2(n10997), .A(n11346), .ZN(n10999) );
  NAND2_X1 U12818 ( .A1(n10999), .A2(n15718), .ZN(n11000) );
  OAI211_X1 U12819 ( .C1(n11350), .C2(n11002), .A(n11001), .B(n11000), .ZN(
        P2_U3225) );
  INV_X1 U12820 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n11005) );
  NAND2_X1 U12821 ( .A1(n11003), .A2(n7419), .ZN(n11004) );
  OAI21_X1 U12822 ( .B1(n7419), .B2(n11005), .A(n11004), .ZN(P2_U3433) );
  NAND2_X1 U12823 ( .A1(n11007), .A2(n11006), .ZN(n11008) );
  INV_X1 U12824 ( .A(n11104), .ZN(n11014) );
  NAND2_X1 U12825 ( .A1(n11008), .A2(n11014), .ZN(n11102) );
  OAI21_X1 U12826 ( .B1(n11008), .B2(n11014), .A(n11102), .ZN(n11265) );
  INV_X1 U12827 ( .A(n11009), .ZN(n11010) );
  NOR2_X1 U12828 ( .A1(n11009), .A2(n7430), .ZN(n11111) );
  INV_X1 U12829 ( .A(n11111), .ZN(n11113) );
  OAI21_X1 U12830 ( .B1(n11100), .B2(n11010), .A(n11113), .ZN(n11263) );
  OAI22_X1 U12831 ( .A1(n11263), .A2(n16198), .B1(n11100), .B2(n16333), .ZN(
        n11018) );
  NAND2_X1 U12832 ( .A1(n11074), .A2(n11236), .ZN(n11012) );
  NAND2_X1 U12833 ( .A1(n11013), .A2(n11012), .ZN(n11105) );
  XNOR2_X1 U12834 ( .A(n11105), .B(n11014), .ZN(n11017) );
  OAI22_X1 U12835 ( .A1(n11297), .A2(n15408), .B1(n11074), .B2(n15406), .ZN(
        n11015) );
  AOI21_X1 U12836 ( .B1(n11265), .B2(n16160), .A(n11015), .ZN(n11016) );
  OAI21_X1 U12837 ( .B1(n16280), .B2(n11017), .A(n11016), .ZN(n11259) );
  AOI211_X1 U12838 ( .C1(n16257), .C2(n11265), .A(n11018), .B(n11259), .ZN(
        n16069) );
  NAND2_X1 U12839 ( .A1(n16339), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n11019) );
  OAI21_X1 U12840 ( .B1(n16069), .B2(n16339), .A(n11019), .ZN(P1_U3530) );
  NAND2_X1 U12841 ( .A1(n11021), .A2(n11020), .ZN(n11023) );
  XOR2_X1 U12842 ( .A(n11023), .B(n11022), .Z(n11035) );
  NOR2_X1 U12843 ( .A1(n15997), .A2(n11024), .ZN(n11034) );
  NAND2_X1 U12844 ( .A1(n11025), .A2(n9340), .ZN(n11026) );
  AND2_X1 U12845 ( .A1(n15978), .A2(n11026), .ZN(n11032) );
  NAND2_X1 U12846 ( .A1(n11027), .A2(n9344), .ZN(n11028) );
  NAND2_X1 U12847 ( .A1(n15972), .A2(n11028), .ZN(n11029) );
  NAND2_X1 U12848 ( .A1(n15973), .A2(n11029), .ZN(n11031) );
  AND2_X1 U12849 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n11836) );
  AOI21_X1 U12850 ( .B1(n15646), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n11836), .ZN(
        n11030) );
  OAI211_X1 U12851 ( .C1(n11032), .C2(n16013), .A(n11031), .B(n11030), .ZN(
        n11033) );
  AOI211_X1 U12852 ( .C1(n11035), .C2(n16017), .A(n11034), .B(n11033), .ZN(
        n11036) );
  INV_X1 U12853 ( .A(n11036), .ZN(P3_U3187) );
  INV_X1 U12854 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n11067) );
  NAND2_X1 U12855 ( .A1(n7422), .A2(n11367), .ZN(n11039) );
  NAND2_X1 U12856 ( .A1(n14689), .A2(n11422), .ZN(n11040) );
  NAND2_X1 U12857 ( .A1(n11203), .A2(n11202), .ZN(n11042) );
  NAND2_X1 U12858 ( .A1(n11195), .A2(n11422), .ZN(n11041) );
  NAND2_X1 U12859 ( .A1(n11043), .A2(n12412), .ZN(n11046) );
  OR2_X1 U12860 ( .A1(n13618), .A2(n11044), .ZN(n11045) );
  OAI211_X1 U12861 ( .C1(n11131), .C2(n11047), .A(n11046), .B(n11045), .ZN(
        n13691) );
  XNOR2_X1 U12862 ( .A(n14688), .B(n11389), .ZN(n13626) );
  XNOR2_X1 U12863 ( .A(n11388), .B(n13626), .ZN(n11063) );
  INV_X1 U12864 ( .A(n11063), .ZN(n11462) );
  NAND3_X1 U12865 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_5__SCAN_IN), 
        .A3(P2_REG3_REG_3__SCAN_IN), .ZN(n11140) );
  INV_X1 U12866 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n11049) );
  NAND2_X1 U12867 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n11048) );
  NAND2_X1 U12868 ( .A1(n11049), .A2(n11048), .ZN(n11050) );
  AND2_X1 U12869 ( .A1(n11140), .A2(n11050), .ZN(n11447) );
  NAND2_X1 U12870 ( .A1(n13522), .A2(n11447), .ZN(n11054) );
  NAND2_X1 U12871 ( .A1(n13523), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n11053) );
  NAND2_X1 U12872 ( .A1(n7425), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n11052) );
  NAND2_X1 U12873 ( .A1(n13517), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n11051) );
  INV_X1 U12874 ( .A(n14687), .ZN(n11534) );
  OAI22_X1 U12875 ( .A1(n11195), .A2(n14914), .B1(n11534), .B2(n14916), .ZN(
        n11062) );
  NAND2_X1 U12876 ( .A1(n11056), .A2(n11055), .ZN(n11205) );
  NAND2_X1 U12877 ( .A1(n11204), .A2(n11059), .ZN(n11058) );
  INV_X1 U12878 ( .A(n13626), .ZN(n11057) );
  NAND2_X1 U12879 ( .A1(n11058), .A2(n11057), .ZN(n11393) );
  NAND3_X1 U12880 ( .A1(n11204), .A2(n13626), .A3(n11059), .ZN(n11060) );
  AOI21_X1 U12881 ( .B1(n11393), .B2(n11060), .A(n14821), .ZN(n11061) );
  AOI211_X1 U12882 ( .C1(n11063), .C2(n14902), .A(n11062), .B(n11061), .ZN(
        n11454) );
  OAI21_X1 U12883 ( .B1(n11211), .B2(n11389), .A(n11399), .ZN(n11458) );
  INV_X1 U12884 ( .A(n11458), .ZN(n11064) );
  AOI22_X1 U12885 ( .A1(n11064), .A2(n15027), .B1(n15026), .B2(n13691), .ZN(
        n11065) );
  OAI211_X1 U12886 ( .C1(n15031), .C2(n11462), .A(n11454), .B(n11065), .ZN(
        n15033) );
  NAND2_X1 U12887 ( .A1(n15033), .A2(n7419), .ZN(n11066) );
  OAI21_X1 U12888 ( .B1(n7419), .B2(n11067), .A(n11066), .ZN(P2_U3442) );
  OAI222_X1 U12889 ( .A1(P3_U3151), .A2(n14100), .B1(n13926), .B2(n11069), 
        .C1(n13924), .C2(n11068), .ZN(P3_U3279) );
  NAND3_X1 U12890 ( .A1(n11072), .A2(n11071), .A3(n11070), .ZN(n13349) );
  OR2_X1 U12891 ( .A1(n16275), .A2(n16170), .ZN(n15435) );
  NOR2_X1 U12892 ( .A1(n16160), .A2(n16330), .ZN(n11073) );
  OAI22_X1 U12893 ( .A1(n11074), .A2(n15408), .B1(n11073), .B2(n16033), .ZN(
        n16035) );
  INV_X1 U12894 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n11075) );
  OAI22_X1 U12895 ( .A1(n16179), .A2(n11076), .B1(n11075), .B2(n16110), .ZN(
        n11077) );
  AOI21_X1 U12896 ( .B1(n16179), .B2(n16035), .A(n11077), .ZN(n11082) );
  INV_X1 U12897 ( .A(n11078), .ZN(n11079) );
  OAI21_X1 U12898 ( .B1(n16073), .B2(n16265), .A(n11080), .ZN(n11081) );
  OAI211_X1 U12899 ( .C1(n16033), .C2(n15435), .A(n11082), .B(n11081), .ZN(
        P1_U3293) );
  NOR2_X1 U12900 ( .A1(n11083), .A2(n16102), .ZN(n11084) );
  AOI22_X1 U12901 ( .A1(n16042), .A2(n11084), .B1(n14304), .B2(n16040), .ZN(
        n11478) );
  MUX2_X1 U12902 ( .A(n10168), .B(n11478), .S(n16238), .Z(n11085) );
  OAI21_X1 U12903 ( .B1(n11481), .B2(n14418), .A(n11085), .ZN(P3_U3459) );
  AOI21_X1 U12904 ( .B1(n11087), .B2(n15961), .A(n11086), .ZN(n11099) );
  INV_X1 U12905 ( .A(n16013), .ZN(n15979) );
  XNOR2_X1 U12906 ( .A(n11088), .B(P3_REG1_REG_1__SCAN_IN), .ZN(n11095) );
  NAND2_X1 U12907 ( .A1(n15646), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n11089) );
  OAI21_X1 U12908 ( .B1(P3_STATE_REG_SCAN_IN), .B2(n11234), .A(n11089), .ZN(
        n11094) );
  NAND2_X1 U12909 ( .A1(n11090), .A2(n11438), .ZN(n11091) );
  AOI21_X1 U12910 ( .B1(n11092), .B2(n11091), .A(n16009), .ZN(n11093) );
  AOI211_X1 U12911 ( .C1(n15979), .C2(n11095), .A(n11094), .B(n11093), .ZN(
        n11098) );
  NAND2_X1 U12912 ( .A1(n16020), .A2(n11096), .ZN(n11097) );
  OAI211_X1 U12913 ( .C1(n11099), .C2(n15960), .A(n11098), .B(n11097), .ZN(
        P3_U3183) );
  INV_X1 U12914 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n11118) );
  NAND2_X1 U12915 ( .A1(n11106), .A2(n11100), .ZN(n11101) );
  NAND2_X1 U12916 ( .A1(n11102), .A2(n11101), .ZN(n11103) );
  NAND2_X1 U12917 ( .A1(n11103), .A2(n8967), .ZN(n11299) );
  OAI21_X1 U12918 ( .B1(n11103), .B2(n8967), .A(n11299), .ZN(n16079) );
  INV_X1 U12919 ( .A(n16079), .ZN(n11116) );
  NAND2_X1 U12920 ( .A1(n11105), .A2(n11104), .ZN(n11108) );
  NAND2_X1 U12921 ( .A1(n11106), .A2(n7430), .ZN(n11107) );
  XNOR2_X1 U12922 ( .A(n11304), .B(n11109), .ZN(n11110) );
  AOI222_X1 U12923 ( .A1(n16330), .A2(n11110), .B1(n15192), .B2(n15457), .C1(
        n15194), .C2(n15455), .ZN(n16070) );
  NAND2_X1 U12924 ( .A1(n11111), .A2(n16077), .ZN(n11301) );
  AOI21_X1 U12925 ( .B1(n11114), .B2(n11113), .A(n11112), .ZN(n16072) );
  AOI22_X1 U12926 ( .A1(n16072), .A2(n16247), .B1(n16278), .B2(n11114), .ZN(
        n11115) );
  OAI211_X1 U12927 ( .C1(n16299), .C2(n11116), .A(n16070), .B(n11115), .ZN(
        n11119) );
  NAND2_X1 U12928 ( .A1(n11119), .A2(n16345), .ZN(n11117) );
  OAI21_X1 U12929 ( .B1(n16345), .B2(n11118), .A(n11117), .ZN(P1_U3468) );
  INV_X1 U12930 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n11121) );
  NAND2_X1 U12931 ( .A1(n11119), .A2(n16341), .ZN(n11120) );
  OAI21_X1 U12932 ( .B1(n16341), .B2(n11121), .A(n11120), .ZN(P1_U3531) );
  INV_X1 U12933 ( .A(n11122), .ZN(n11123) );
  XNOR2_X1 U12934 ( .A(n13691), .B(n14553), .ZN(n11127) );
  BUF_X2 U12935 ( .A(n11126), .Z(n14552) );
  NAND2_X1 U12936 ( .A1(n14688), .A2(n14552), .ZN(n11128) );
  XNOR2_X1 U12937 ( .A(n11127), .B(n11128), .ZN(n11193) );
  INV_X1 U12938 ( .A(n11127), .ZN(n11129) );
  NAND2_X1 U12939 ( .A1(n11129), .A2(n11128), .ZN(n11135) );
  NAND2_X1 U12940 ( .A1(n14687), .A2(n14552), .ZN(n11597) );
  NAND2_X1 U12941 ( .A1(n11130), .A2(n12412), .ZN(n11134) );
  INV_X2 U12942 ( .A(n13618), .ZN(n13406) );
  XNOR2_X1 U12943 ( .A(n13706), .B(n14553), .ZN(n11595) );
  XOR2_X1 U12944 ( .A(n11597), .B(n11595), .Z(n11136) );
  AND3_X1 U12945 ( .A1(n11192), .A2(n11136), .A3(n11135), .ZN(n11137) );
  OAI21_X1 U12946 ( .B1(n11596), .B2(n11137), .A(n14658), .ZN(n11150) );
  INV_X4 U12947 ( .A(n12545), .ZN(n13523) );
  NAND2_X1 U12948 ( .A1(n13523), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n11145) );
  NAND2_X1 U12949 ( .A1(n7425), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n11144) );
  INV_X1 U12950 ( .A(n11140), .ZN(n11138) );
  NAND2_X1 U12951 ( .A1(n11138), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n11548) );
  INV_X1 U12952 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n11139) );
  NAND2_X1 U12953 ( .A1(n11140), .A2(n11139), .ZN(n11141) );
  AND2_X1 U12954 ( .A1(n11548), .A2(n11141), .ZN(n14647) );
  NAND2_X1 U12955 ( .A1(n13522), .A2(n14647), .ZN(n11143) );
  NAND2_X1 U12956 ( .A1(n13517), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n11142) );
  NAND4_X1 U12957 ( .A1(n11145), .A2(n11144), .A3(n11143), .A4(n11142), .ZN(
        n14686) );
  INV_X1 U12958 ( .A(n14686), .ZN(n11556) );
  OAI21_X1 U12959 ( .B1(n14663), .B2(n11556), .A(n11146), .ZN(n11148) );
  INV_X1 U12960 ( .A(n13706), .ZN(n11537) );
  OAI22_X1 U12961 ( .A1(n14670), .A2(n11537), .B1(n11394), .B2(n14661), .ZN(
        n11147) );
  AOI211_X1 U12962 ( .C1(n11447), .C2(n14667), .A(n11148), .B(n11147), .ZN(
        n11149) );
  NAND2_X1 U12963 ( .A1(n11150), .A2(n11149), .ZN(P2_U3199) );
  NAND2_X1 U12964 ( .A1(n11151), .A2(n10176), .ZN(n11152) );
  NAND2_X1 U12965 ( .A1(n11153), .A2(n11152), .ZN(n11154) );
  NAND2_X1 U12966 ( .A1(n15973), .A2(n11154), .ZN(n11162) );
  NAND2_X1 U12967 ( .A1(n11155), .A2(n10175), .ZN(n11156) );
  NAND2_X1 U12968 ( .A1(n11157), .A2(n11156), .ZN(n11158) );
  NAND2_X1 U12969 ( .A1(n15979), .A2(n11158), .ZN(n11161) );
  INV_X1 U12970 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n11159) );
  NOR2_X1 U12971 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11159), .ZN(n11416) );
  AOI21_X1 U12972 ( .B1(n15646), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n11416), .ZN(
        n11160) );
  NAND3_X1 U12973 ( .A1(n11162), .A2(n11161), .A3(n11160), .ZN(n11170) );
  INV_X1 U12974 ( .A(n11163), .ZN(n11164) );
  NAND3_X1 U12975 ( .A1(n11166), .A2(n11165), .A3(n11164), .ZN(n11167) );
  AOI21_X1 U12976 ( .B1(n11168), .B2(n11167), .A(n15960), .ZN(n11169) );
  AOI211_X1 U12977 ( .C1(n16020), .C2(n11171), .A(n11170), .B(n11169), .ZN(
        n11172) );
  INV_X1 U12978 ( .A(n11172), .ZN(P3_U3185) );
  INV_X1 U12979 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n11173) );
  MUX2_X1 U12980 ( .A(n11173), .B(P1_REG1_REG_10__SCAN_IN), .S(n11319), .Z(
        n11177) );
  OAI21_X1 U12981 ( .B1(n11175), .B2(P1_REG1_REG_9__SCAN_IN), .A(n11174), .ZN(
        n11176) );
  NOR2_X1 U12982 ( .A1(n11176), .A2(n11177), .ZN(n11318) );
  AOI211_X1 U12983 ( .C1(n11177), .C2(n11176), .A(n15240), .B(n11318), .ZN(
        n11191) );
  INV_X1 U12984 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n11178) );
  MUX2_X1 U12985 ( .A(n11178), .B(P1_REG2_REG_10__SCAN_IN), .S(n11319), .Z(
        n11181) );
  NOR2_X1 U12986 ( .A1(n11179), .A2(n11936), .ZN(n11183) );
  INV_X1 U12987 ( .A(n11183), .ZN(n11180) );
  NAND2_X1 U12988 ( .A1(n11181), .A2(n11180), .ZN(n11184) );
  MUX2_X1 U12989 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n11178), .S(n11319), .Z(
        n11182) );
  OAI21_X1 U12990 ( .B1(n11185), .B2(n11183), .A(n11182), .ZN(n11316) );
  OAI211_X1 U12991 ( .C1(n11185), .C2(n11184), .A(n11316), .B(n15780), .ZN(
        n11188) );
  NAND2_X1 U12992 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n12278)
         );
  INV_X1 U12993 ( .A(n12278), .ZN(n11186) );
  AOI21_X1 U12994 ( .B1(n15757), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n11186), 
        .ZN(n11187) );
  OAI211_X1 U12995 ( .C1(n15765), .C2(n11189), .A(n11188), .B(n11187), .ZN(
        n11190) );
  OR2_X1 U12996 ( .A1(n11191), .A2(n11190), .ZN(P1_U3253) );
  OAI21_X1 U12997 ( .B1(n11194), .B2(n11193), .A(n11192), .ZN(n11200) );
  OAI22_X1 U12998 ( .A1(n14670), .A2(n11389), .B1(n11195), .B2(n14661), .ZN(
        n11199) );
  NAND2_X1 U12999 ( .A1(n14667), .A2(n11456), .ZN(n11196) );
  OAI211_X1 U13000 ( .C1(n14663), .C2(n11534), .A(n11197), .B(n11196), .ZN(
        n11198) );
  AOI211_X1 U13001 ( .C1(n11200), .C2(n14658), .A(n11199), .B(n11198), .ZN(
        n11201) );
  INV_X1 U13002 ( .A(n11201), .ZN(P2_U3202) );
  XNOR2_X1 U13003 ( .A(n11202), .B(n11203), .ZN(n11424) );
  INV_X1 U13004 ( .A(n11424), .ZN(n11213) );
  OAI21_X1 U13005 ( .B1(n13625), .B2(n11205), .A(n11204), .ZN(n11208) );
  OAI22_X1 U13006 ( .A1(n7422), .A2(n14914), .B1(n11394), .B2(n14916), .ZN(
        n11207) );
  NOR2_X1 U13007 ( .A1(n11213), .A2(n10661), .ZN(n11206) );
  AOI211_X1 U13008 ( .C1(n14924), .C2(n11208), .A(n11207), .B(n11206), .ZN(
        n11426) );
  AND2_X1 U13009 ( .A1(n11209), .A2(n13695), .ZN(n11210) );
  NOR2_X1 U13010 ( .A1(n11211), .A2(n11210), .ZN(n11420) );
  AOI22_X1 U13011 ( .A1(n11420), .A2(n15027), .B1(n15026), .B2(n13695), .ZN(
        n11212) );
  OAI211_X1 U13012 ( .C1(n11213), .C2(n15031), .A(n11426), .B(n11212), .ZN(
        n11216) );
  NAND2_X1 U13013 ( .A1(n11216), .A2(n16293), .ZN(n11214) );
  OAI21_X1 U13014 ( .B1(n16293), .B2(n11215), .A(n11214), .ZN(P2_U3502) );
  INV_X1 U13015 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n11218) );
  NAND2_X1 U13016 ( .A1(n11216), .A2(n7419), .ZN(n11217) );
  OAI21_X1 U13017 ( .B1(n7419), .B2(n11218), .A(n11217), .ZN(P2_U3439) );
  INV_X1 U13018 ( .A(n12211), .ZN(n11225) );
  NAND2_X1 U13019 ( .A1(n11220), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n11219) );
  MUX2_X1 U13020 ( .A(P2_IR_REG_31__SCAN_IN), .B(n11219), .S(
        P2_IR_REG_14__SCAN_IN), .Z(n11223) );
  INV_X1 U13021 ( .A(n11220), .ZN(n11222) );
  NAND2_X1 U13022 ( .A1(n11222), .A2(n11221), .ZN(n11291) );
  NAND2_X1 U13023 ( .A1(n11223), .A2(n11291), .ZN(n15680) );
  OAI222_X1 U13024 ( .A1(n13255), .A2(n11224), .B1(n15061), .B2(n11225), .C1(
        P2_U3088), .C2(n15680), .ZN(P2_U3313) );
  INV_X1 U13025 ( .A(n12619), .ZN(n12625) );
  OAI222_X1 U13026 ( .A1(n15597), .A2(n11226), .B1(n15604), .B2(n11225), .C1(
        P1_U3086), .C2(n12625), .ZN(P1_U3341) );
  NOR2_X1 U13027 ( .A1(n14023), .A2(P3_U3151), .ZN(n16045) );
  OAI21_X1 U13028 ( .B1(n11229), .B2(n11228), .A(n11227), .ZN(n11230) );
  NAND2_X1 U13029 ( .A1(n11230), .A2(n16041), .ZN(n11233) );
  INV_X1 U13030 ( .A(n14015), .ZN(n14034) );
  OAI22_X1 U13031 ( .A1(n14032), .A2(n11427), .B1(n14017), .B2(n11247), .ZN(
        n11231) );
  AOI21_X1 U13032 ( .B1(n14034), .B2(n14059), .A(n11231), .ZN(n11232) );
  OAI211_X1 U13033 ( .C1(n16045), .C2(n11234), .A(n11233), .B(n11232), .ZN(
        P3_U3162) );
  MUX2_X1 U13034 ( .A(n11235), .B(P1_REG2_REG_1__SCAN_IN), .S(n16264), .Z(
        n11240) );
  INV_X1 U13035 ( .A(n16110), .ZN(n16262) );
  AOI22_X1 U13036 ( .A1(n16265), .A2(n11236), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n16262), .ZN(n11237) );
  OAI21_X1 U13037 ( .B1(n15416), .B2(n11238), .A(n11237), .ZN(n11239) );
  AOI211_X1 U13038 ( .C1(n16270), .C2(n11241), .A(n11240), .B(n11239), .ZN(
        n11242) );
  INV_X1 U13039 ( .A(n11242), .ZN(P1_U3292) );
  INV_X1 U13040 ( .A(n11243), .ZN(n11244) );
  NAND2_X1 U13041 ( .A1(n11244), .A2(n11251), .ZN(n11246) );
  NAND2_X1 U13042 ( .A1(n11246), .A2(n11245), .ZN(n11439) );
  NOR2_X1 U13043 ( .A1(n11247), .A2(n16231), .ZN(n11436) );
  AOI21_X1 U13044 ( .B1(n11439), .B2(n16103), .A(n11436), .ZN(n11255) );
  NAND2_X1 U13045 ( .A1(n16038), .A2(n9714), .ZN(n11248) );
  OAI21_X1 U13046 ( .B1(n11251), .B2(n11248), .A(n16054), .ZN(n11249) );
  NAND2_X1 U13047 ( .A1(n11249), .A2(n14059), .ZN(n11254) );
  AND2_X1 U13048 ( .A1(n11250), .A2(n9714), .ZN(n11252) );
  AOI22_X1 U13049 ( .A1(n11252), .A2(n11251), .B1(n14304), .B2(n14058), .ZN(
        n11253) );
  AND2_X1 U13050 ( .A1(n11254), .A2(n11253), .ZN(n11433) );
  AND2_X1 U13051 ( .A1(n11255), .A2(n11433), .ZN(n16047) );
  MUX2_X1 U13052 ( .A(n16047), .B(n11256), .S(n9764), .Z(n11257) );
  INV_X1 U13053 ( .A(n11257), .ZN(P3_U3460) );
  OAI222_X1 U13054 ( .A1(P3_U3151), .A2(n14129), .B1(n13926), .B2(n12737), 
        .C1(n13924), .C2(n11258), .ZN(P3_U3278) );
  INV_X1 U13055 ( .A(n11259), .ZN(n11267) );
  INV_X2 U13056 ( .A(n16179), .ZN(n16264) );
  NAND2_X1 U13057 ( .A1(n16265), .A2(n7430), .ZN(n11262) );
  AOI22_X1 U13058 ( .A1(n16264), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n16262), .ZN(n11261) );
  OAI211_X1 U13059 ( .C1(n11263), .C2(n15416), .A(n11262), .B(n11261), .ZN(
        n11264) );
  AOI21_X1 U13060 ( .B1(n16270), .B2(n11265), .A(n11264), .ZN(n11266) );
  OAI21_X1 U13061 ( .B1(n11267), .B2(n16264), .A(n11266), .ZN(P1_U3291) );
  NAND2_X1 U13062 ( .A1(n15192), .A2(n13572), .ZN(n11269) );
  NAND2_X1 U13063 ( .A1(n11341), .A2(n13265), .ZN(n11268) );
  AND2_X1 U13064 ( .A1(n11269), .A2(n11268), .ZN(n11273) );
  NAND2_X1 U13065 ( .A1(n11271), .A2(n11270), .ZN(n11274) );
  OAI22_X1 U13066 ( .A1(n11484), .A2(n13588), .B1(n8053), .B2(n13594), .ZN(
        n11272) );
  XNOR2_X1 U13067 ( .A(n11272), .B(n11815), .ZN(n11337) );
  NAND2_X1 U13068 ( .A1(n11587), .A2(n13578), .ZN(n11277) );
  NAND2_X1 U13069 ( .A1(n15191), .A2(n13265), .ZN(n11276) );
  NAND2_X1 U13070 ( .A1(n11277), .A2(n11276), .ZN(n11278) );
  XNOR2_X1 U13071 ( .A(n11278), .B(n11815), .ZN(n11282) );
  NAND2_X1 U13072 ( .A1(n11587), .A2(n13265), .ZN(n11280) );
  NAND2_X1 U13073 ( .A1(n15191), .A2(n13572), .ZN(n11279) );
  NAND2_X1 U13074 ( .A1(n11280), .A2(n11279), .ZN(n11281) );
  NAND2_X1 U13075 ( .A1(n11282), .A2(n11281), .ZN(n11463) );
  NAND2_X1 U13076 ( .A1(n7569), .A2(n11463), .ZN(n11283) );
  XNOR2_X1 U13077 ( .A(n11464), .B(n11283), .ZN(n11288) );
  AOI22_X1 U13078 ( .A1(n16351), .A2(n15190), .B1(P1_REG3_REG_5__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11285) );
  NAND2_X1 U13079 ( .A1(n15167), .A2(n11586), .ZN(n11284) );
  OAI211_X1 U13080 ( .C1(n11484), .C2(n15159), .A(n11285), .B(n11284), .ZN(
        n11286) );
  AOI21_X1 U13081 ( .B1(n11587), .B2(n15173), .A(n11286), .ZN(n11287) );
  OAI21_X1 U13082 ( .B1(n11288), .B2(n15175), .A(n11287), .ZN(P1_U3227) );
  INV_X1 U13083 ( .A(n12413), .ZN(n11293) );
  INV_X1 U13084 ( .A(n12627), .ZN(n15766) );
  OAI222_X1 U13085 ( .A1(n15597), .A2(n11289), .B1(n15604), .B2(n11293), .C1(
        P1_U3086), .C2(n15766), .ZN(P1_U3340) );
  NAND2_X1 U13086 ( .A1(n11291), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n11290) );
  MUX2_X1 U13087 ( .A(P2_IR_REG_31__SCAN_IN), .B(n11290), .S(
        P2_IR_REG_15__SCAN_IN), .Z(n11292) );
  AND2_X1 U13088 ( .A1(n11292), .A2(n11733), .ZN(n12414) );
  INV_X1 U13089 ( .A(n12414), .ZN(n12337) );
  OAI222_X1 U13090 ( .A1(n13255), .A2(n11294), .B1(n15061), .B2(n11293), .C1(
        P2_U3088), .C2(n12337), .ZN(P2_U3312) );
  INV_X1 U13091 ( .A(n11295), .ZN(n11296) );
  NAND2_X1 U13092 ( .A1(n11297), .A2(n16077), .ZN(n11298) );
  OAI21_X1 U13093 ( .B1(n11300), .B2(n11488), .A(n11486), .ZN(n16085) );
  NAND2_X1 U13094 ( .A1(n11301), .A2(n11341), .ZN(n11302) );
  NAND2_X1 U13095 ( .A1(n11509), .A2(n11302), .ZN(n16082) );
  AOI22_X1 U13096 ( .A1(n16265), .A2(n11341), .B1(n11342), .B2(n16262), .ZN(
        n11303) );
  OAI21_X1 U13097 ( .B1(n15416), .B2(n16082), .A(n11303), .ZN(n11311) );
  NAND2_X1 U13098 ( .A1(n15193), .A2(n16077), .ZN(n11305) );
  XNOR2_X1 U13099 ( .A(n11490), .B(n11488), .ZN(n11307) );
  NAND2_X1 U13100 ( .A1(n11307), .A2(n16330), .ZN(n11309) );
  AOI22_X1 U13101 ( .A1(n15455), .A2(n15193), .B1(n15191), .B2(n15457), .ZN(
        n11308) );
  NAND2_X1 U13102 ( .A1(n11309), .A2(n11308), .ZN(n16083) );
  MUX2_X1 U13103 ( .A(n16083), .B(P1_REG2_REG_4__SCAN_IN), .S(n16264), .Z(
        n11310) );
  AOI211_X1 U13104 ( .C1(n15366), .C2(n16085), .A(n11311), .B(n11310), .ZN(
        n11312) );
  INV_X1 U13105 ( .A(n11312), .ZN(P1_U3289) );
  NAND2_X1 U13106 ( .A1(n11319), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n11315) );
  INV_X1 U13107 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11313) );
  MUX2_X1 U13108 ( .A(n11313), .B(P1_REG2_REG_11__SCAN_IN), .S(n11711), .Z(
        n11314) );
  AOI21_X1 U13109 ( .B1(n11316), .B2(n11315), .A(n11314), .ZN(n11710) );
  NAND3_X1 U13110 ( .A1(n11316), .A2(n11315), .A3(n11314), .ZN(n11317) );
  NAND2_X1 U13111 ( .A1(n11317), .A2(n15780), .ZN(n11327) );
  MUX2_X1 U13112 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n7716), .S(n11711), .Z(
        n11320) );
  OAI21_X1 U13113 ( .B1(n11321), .B2(n11320), .A(n11705), .ZN(n11322) );
  NAND2_X1 U13114 ( .A1(n11322), .A2(n15776), .ZN(n11326) );
  NOR2_X1 U13115 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n12392), .ZN(n11324) );
  NOR2_X1 U13116 ( .A1(n15765), .A2(n7717), .ZN(n11323) );
  AOI211_X1 U13117 ( .C1(n15757), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n11324), 
        .B(n11323), .ZN(n11325) );
  OAI211_X1 U13118 ( .C1(n11710), .C2(n11327), .A(n11326), .B(n11325), .ZN(
        P1_U3254) );
  OAI21_X1 U13119 ( .B1(n11330), .B2(n11329), .A(n11328), .ZN(n11331) );
  NAND2_X1 U13120 ( .A1(n11331), .A2(n16041), .ZN(n11335) );
  INV_X1 U13121 ( .A(n14057), .ZN(n16055) );
  OAI22_X1 U13122 ( .A1(n14032), .A2(n16055), .B1(n14017), .B2(n16049), .ZN(
        n11333) );
  NOR2_X1 U13123 ( .A1(n14015), .A2(n7579), .ZN(n11332) );
  NOR2_X1 U13124 ( .A1(n11333), .A2(n11332), .ZN(n11334) );
  OAI211_X1 U13125 ( .C1(n16045), .C2(n16060), .A(n11335), .B(n11334), .ZN(
        P3_U3177) );
  OAI222_X1 U13126 ( .A1(P3_U3151), .A2(n14148), .B1(n13926), .B2(n12736), 
        .C1(n13924), .C2(n11336), .ZN(P3_U3277) );
  NOR2_X1 U13127 ( .A1(n7455), .A2(n7566), .ZN(n11338) );
  XNOR2_X1 U13128 ( .A(n11338), .B(n11337), .ZN(n11345) );
  INV_X1 U13129 ( .A(n15191), .ZN(n11493) );
  OAI21_X1 U13130 ( .B1(n15170), .B2(n11493), .A(n11339), .ZN(n11340) );
  AOI21_X1 U13131 ( .B1(n16349), .B2(n15193), .A(n11340), .ZN(n11344) );
  AOI22_X1 U13132 ( .A1(n11342), .A2(n15167), .B1(n15173), .B2(n11341), .ZN(
        n11343) );
  OAI211_X1 U13133 ( .C1(n11345), .C2(n15175), .A(n11344), .B(n11343), .ZN(
        P1_U3230) );
  INV_X1 U13134 ( .A(n11346), .ZN(n11347) );
  AOI21_X1 U13135 ( .B1(n11348), .B2(n10996), .A(n11347), .ZN(n12242) );
  XOR2_X1 U13136 ( .A(n11354), .B(n12242), .Z(n11349) );
  NOR2_X1 U13137 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n11349), .ZN(n12244) );
  AOI21_X1 U13138 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n11349), .A(n12244), 
        .ZN(n11358) );
  AOI21_X1 U13139 ( .B1(n12021), .B2(P2_REG1_REG_11__SCAN_IN), .A(n11350), 
        .ZN(n11352) );
  INV_X1 U13140 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n12358) );
  MUX2_X1 U13141 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n12358), .S(n12243), .Z(
        n11351) );
  NAND2_X1 U13142 ( .A1(n11352), .A2(n11351), .ZN(n12238) );
  OAI21_X1 U13143 ( .B1(n11352), .B2(n11351), .A(n12238), .ZN(n11356) );
  NAND2_X1 U13144 ( .A1(n15683), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n11353) );
  NAND2_X1 U13145 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n12372)
         );
  OAI211_X1 U13146 ( .C1(n11354), .C2(n15724), .A(n11353), .B(n12372), .ZN(
        n11355) );
  AOI21_X1 U13147 ( .B1(n11356), .B2(n15743), .A(n11355), .ZN(n11357) );
  OAI21_X1 U13148 ( .B1(n11358), .B2(n15736), .A(n11357), .ZN(P2_U3226) );
  NOR3_X1 U13149 ( .A1(n15648), .A2(n11359), .A3(n15649), .ZN(n11360) );
  NAND2_X1 U13150 ( .A1(n11361), .A2(n11360), .ZN(n11894) );
  INV_X1 U13151 ( .A(n13666), .ZN(n13895) );
  NAND2_X1 U13152 ( .A1(n13895), .A2(n7415), .ZN(n11563) );
  INV_X1 U13153 ( .A(n11563), .ZN(n11362) );
  MUX2_X1 U13154 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n11363), .S(n14843), .Z(
        n11369) );
  NOR2_X2 U13155 ( .A1(n11894), .A2(n14552), .ZN(n14936) );
  AOI22_X1 U13156 ( .A1(n14936), .A2(n11365), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n14929), .ZN(n11366) );
  OAI21_X1 U13157 ( .B1(n11367), .B2(n14932), .A(n11366), .ZN(n11368) );
  AOI211_X1 U13158 ( .C1(n14908), .C2(n11370), .A(n11369), .B(n11368), .ZN(
        n11371) );
  INV_X1 U13159 ( .A(n11371), .ZN(P2_U3263) );
  XOR2_X1 U13160 ( .A(n11373), .B(n11372), .Z(n11387) );
  OAI21_X1 U13161 ( .B1(n7978), .B2(n7977), .A(n11375), .ZN(n11385) );
  NOR2_X1 U13162 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11376), .ZN(n12262) );
  AOI21_X1 U13163 ( .B1(n15646), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n12262), .ZN(
        n11377) );
  OAI21_X1 U13164 ( .B1(n15997), .B2(n11378), .A(n11377), .ZN(n11384) );
  NAND2_X1 U13165 ( .A1(n11380), .A2(n11379), .ZN(n11381) );
  AOI21_X1 U13166 ( .B1(n11382), .B2(n11381), .A(n16013), .ZN(n11383) );
  AOI211_X1 U13167 ( .C1(n15973), .C2(n11385), .A(n11384), .B(n11383), .ZN(
        n11386) );
  OAI21_X1 U13168 ( .B1(n11387), .B2(n15960), .A(n11386), .ZN(P3_U3190) );
  NAND2_X1 U13169 ( .A1(n11388), .A2(n13626), .ZN(n11391) );
  NAND2_X1 U13170 ( .A1(n11394), .A2(n11389), .ZN(n11390) );
  XNOR2_X1 U13171 ( .A(n13706), .B(n14687), .ZN(n13628) );
  XNOR2_X1 U13172 ( .A(n11558), .B(n13628), .ZN(n11453) );
  NAND2_X1 U13173 ( .A1(n11394), .A2(n13691), .ZN(n11392) );
  XNOR2_X1 U13174 ( .A(n11536), .B(n13628), .ZN(n11397) );
  OAI22_X1 U13175 ( .A1(n11394), .A2(n14914), .B1(n11556), .B2(n14916), .ZN(
        n11396) );
  NOR2_X1 U13176 ( .A1(n11453), .A2(n10661), .ZN(n11395) );
  AOI211_X1 U13177 ( .C1(n14924), .C2(n11397), .A(n11396), .B(n11395), .ZN(
        n11444) );
  INV_X1 U13178 ( .A(n11777), .ZN(n11398) );
  AOI21_X1 U13179 ( .B1(n13706), .B2(n11399), .A(n11398), .ZN(n11446) );
  AOI22_X1 U13180 ( .A1(n11446), .A2(n15027), .B1(n15026), .B2(n13706), .ZN(
        n11400) );
  OAI211_X1 U13181 ( .C1(n15031), .C2(n11453), .A(n11444), .B(n11400), .ZN(
        n11403) );
  NAND2_X1 U13182 ( .A1(n11403), .A2(n16293), .ZN(n11401) );
  OAI21_X1 U13183 ( .B1(n16293), .B2(n11402), .A(n11401), .ZN(P2_U3504) );
  INV_X1 U13184 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n11405) );
  NAND2_X1 U13185 ( .A1(n11403), .A2(n7419), .ZN(n11404) );
  OAI21_X1 U13186 ( .B1(n7419), .B2(n11405), .A(n11404), .ZN(P2_U3445) );
  INV_X1 U13187 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n15651) );
  OAI22_X1 U13188 ( .A1(n14843), .A2(n10555), .B1(n15651), .B2(n14840), .ZN(
        n11408) );
  OAI22_X1 U13189 ( .A1(n7431), .A2(n14932), .B1(n14933), .B2(n11406), .ZN(
        n11407) );
  AOI211_X1 U13190 ( .C1(n14936), .C2(n11409), .A(n11408), .B(n11407), .ZN(
        n11410) );
  OAI21_X1 U13191 ( .B1(n14938), .B2(n11411), .A(n11410), .ZN(P2_U3264) );
  NAND2_X1 U13192 ( .A1(n11414), .A2(n11413), .ZN(n11418) );
  OAI22_X1 U13193 ( .A1(n11427), .A2(n14015), .B1(n14032), .B2(n11834), .ZN(
        n11415) );
  AOI211_X1 U13194 ( .C1(n16037), .C2(n11431), .A(n11416), .B(n11415), .ZN(
        n11417) );
  OAI211_X1 U13195 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n14036), .A(n11418), .B(
        n11417), .ZN(P3_U3158) );
  OAI22_X1 U13196 ( .A1(n14843), .A2(n10559), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n14840), .ZN(n11419) );
  AOI21_X1 U13197 ( .B1(n14936), .B2(n11420), .A(n11419), .ZN(n11421) );
  OAI21_X1 U13198 ( .B1(n11422), .B2(n14932), .A(n11421), .ZN(n11423) );
  AOI21_X1 U13199 ( .B1(n14908), .B2(n11424), .A(n11423), .ZN(n11425) );
  OAI21_X1 U13200 ( .B1(n11426), .B2(n14938), .A(n11425), .ZN(P2_U3262) );
  NOR2_X1 U13201 ( .A1(n11427), .A2(n16054), .ZN(n11429) );
  AOI211_X1 U13202 ( .C1(n16103), .C2(n11430), .A(n11429), .B(n11428), .ZN(
        n11525) );
  AOI22_X1 U13203 ( .A1(n12441), .A2(n11431), .B1(n9764), .B2(
        P3_REG1_REG_3__SCAN_IN), .ZN(n11432) );
  OAI21_X1 U13204 ( .B1(n11525), .B2(n9764), .A(n11432), .ZN(P3_U3462) );
  INV_X1 U13205 ( .A(n11433), .ZN(n11434) );
  AOI21_X1 U13206 ( .B1(n11436), .B2(n11435), .A(n11434), .ZN(n11437) );
  MUX2_X1 U13207 ( .A(n11438), .B(n11437), .S(n16100), .Z(n11441) );
  AOI22_X1 U13208 ( .A1(n14339), .A2(n11439), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n16094), .ZN(n11440) );
  NAND2_X1 U13209 ( .A1(n11441), .A2(n11440), .ZN(P3_U3232) );
  INV_X1 U13210 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n11442) );
  MUX2_X1 U13211 ( .A(n11478), .B(n11442), .S(n16239), .Z(n11443) );
  OAI21_X1 U13212 ( .B1(n11481), .B2(n14464), .A(n11443), .ZN(P3_U3390) );
  MUX2_X1 U13213 ( .A(n11445), .B(n11444), .S(n14843), .Z(n11452) );
  INV_X1 U13214 ( .A(n14932), .ZN(n14849) );
  INV_X1 U13215 ( .A(n11446), .ZN(n11449) );
  INV_X1 U13216 ( .A(n11447), .ZN(n11448) );
  OAI22_X1 U13217 ( .A1(n14846), .A2(n11449), .B1(n11448), .B2(n14840), .ZN(
        n11450) );
  AOI21_X1 U13218 ( .B1(n14849), .B2(n13706), .A(n11450), .ZN(n11451) );
  OAI211_X1 U13219 ( .C1(n11453), .C2(n14933), .A(n11452), .B(n11451), .ZN(
        P2_U3260) );
  MUX2_X1 U13220 ( .A(n11455), .B(n11454), .S(n14843), .Z(n11461) );
  INV_X1 U13221 ( .A(n11456), .ZN(n11457) );
  OAI22_X1 U13222 ( .A1(n14846), .A2(n11458), .B1(n11457), .B2(n14840), .ZN(
        n11459) );
  AOI21_X1 U13223 ( .B1(n14849), .B2(n13691), .A(n11459), .ZN(n11460) );
  OAI211_X1 U13224 ( .C1(n11462), .C2(n14933), .A(n11461), .B(n11460), .ZN(
        P2_U3261) );
  INV_X1 U13225 ( .A(n11648), .ZN(n16113) );
  INV_X1 U13226 ( .A(n15190), .ZN(n11496) );
  OAI22_X1 U13227 ( .A1(n16113), .A2(n13588), .B1(n11496), .B2(n13587), .ZN(
        n11654) );
  NAND2_X1 U13228 ( .A1(n11648), .A2(n13578), .ZN(n11466) );
  NAND2_X1 U13229 ( .A1(n15190), .A2(n13265), .ZN(n11465) );
  NAND2_X1 U13230 ( .A1(n11466), .A2(n11465), .ZN(n11467) );
  XNOR2_X1 U13231 ( .A(n11467), .B(n11815), .ZN(n11653) );
  XOR2_X1 U13232 ( .A(n11654), .B(n11653), .Z(n11468) );
  OAI211_X1 U13233 ( .C1(n11469), .C2(n11468), .A(n11656), .B(n16356), .ZN(
        n11476) );
  NAND2_X1 U13234 ( .A1(n15189), .A2(n15457), .ZN(n11471) );
  NAND2_X1 U13235 ( .A1(n15191), .A2(n15455), .ZN(n11470) );
  NAND2_X1 U13236 ( .A1(n11471), .A2(n11470), .ZN(n11645) );
  NAND2_X1 U13237 ( .A1(n15153), .A2(n11645), .ZN(n11472) );
  OAI211_X1 U13238 ( .C1(n16361), .C2(n16109), .A(n11473), .B(n11472), .ZN(
        n11474) );
  INV_X1 U13239 ( .A(n11474), .ZN(n11475) );
  OAI211_X1 U13240 ( .C1(n16113), .C2(n16353), .A(n11476), .B(n11475), .ZN(
        P1_U3239) );
  MUX2_X1 U13241 ( .A(n11478), .B(n11477), .S(n14341), .Z(n11480) );
  NAND2_X1 U13242 ( .A1(n16094), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n11479) );
  OAI211_X1 U13243 ( .C1(n11481), .C2(n14337), .A(n11480), .B(n11479), .ZN(
        P3_U3233) );
  INV_X1 U13244 ( .A(n11482), .ZN(n11483) );
  OAI222_X1 U13245 ( .A1(n13924), .A2(n11483), .B1(n13926), .B2(n12956), .C1(
        P3_U3151), .C2(n14145), .ZN(P3_U3276) );
  NAND2_X1 U13246 ( .A1(n11484), .A2(n8053), .ZN(n11485) );
  INV_X1 U13247 ( .A(n11510), .ZN(n11505) );
  OR2_X1 U13248 ( .A1(n15191), .A2(n11587), .ZN(n11487) );
  XNOR2_X1 U13249 ( .A(n11917), .B(n11924), .ZN(n16136) );
  INV_X1 U13250 ( .A(n11488), .ZN(n11489) );
  NAND2_X1 U13251 ( .A1(n11490), .A2(n11489), .ZN(n11492) );
  NAND2_X1 U13252 ( .A1(n15192), .A2(n8053), .ZN(n11491) );
  NAND2_X1 U13253 ( .A1(n11493), .A2(n11587), .ZN(n11494) );
  NAND2_X1 U13254 ( .A1(n11648), .A2(n11496), .ZN(n11497) );
  XNOR2_X1 U13255 ( .A(n11925), .B(n11924), .ZN(n11500) );
  NAND2_X1 U13256 ( .A1(n15188), .A2(n15457), .ZN(n11499) );
  NAND2_X1 U13257 ( .A1(n15190), .A2(n15455), .ZN(n11498) );
  NAND2_X1 U13258 ( .A1(n11499), .A2(n11498), .ZN(n11662) );
  AOI21_X1 U13259 ( .B1(n11500), .B2(n16330), .A(n11662), .ZN(n16134) );
  MUX2_X1 U13260 ( .A(n16134), .B(n10749), .S(n16264), .Z(n11504) );
  INV_X1 U13261 ( .A(n16132), .ZN(n11668) );
  AOI211_X1 U13262 ( .C1(n16132), .C2(n8050), .A(n16198), .B(n16163), .ZN(
        n16131) );
  OR2_X1 U13263 ( .A1(n13349), .A2(n7429), .ZN(n16181) );
  INV_X1 U13264 ( .A(n11665), .ZN(n11501) );
  OAI22_X1 U13265 ( .A1(n16114), .A2(n11668), .B1(n11501), .B2(n16110), .ZN(
        n11502) );
  AOI21_X1 U13266 ( .B1(n16131), .B2(n16269), .A(n11502), .ZN(n11503) );
  OAI211_X1 U13267 ( .C1(n15466), .C2(n16136), .A(n11504), .B(n11503), .ZN(
        P1_U3286) );
  INV_X1 U13268 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n11517) );
  OR2_X1 U13269 ( .A1(n11506), .A2(n11505), .ZN(n11507) );
  NAND2_X1 U13270 ( .A1(n11508), .A2(n11507), .ZN(n11593) );
  OAI21_X1 U13271 ( .B1(n8051), .B2(n8052), .A(n11647), .ZN(n11589) );
  OAI22_X1 U13272 ( .A1(n11589), .A2(n16198), .B1(n8051), .B2(n16333), .ZN(
        n11515) );
  XNOR2_X1 U13273 ( .A(n11511), .B(n11510), .ZN(n11514) );
  NAND2_X1 U13274 ( .A1(n11593), .A2(n16160), .ZN(n11513) );
  AOI22_X1 U13275 ( .A1(n15455), .A2(n15192), .B1(n15190), .B2(n15457), .ZN(
        n11512) );
  OAI211_X1 U13276 ( .C1(n16280), .C2(n11514), .A(n11513), .B(n11512), .ZN(
        n11590) );
  AOI211_X1 U13277 ( .C1(n16257), .C2(n11593), .A(n11515), .B(n11590), .ZN(
        n11518) );
  OR2_X1 U13278 ( .A1(n11518), .A2(n16342), .ZN(n11516) );
  OAI21_X1 U13279 ( .B1(n16345), .B2(n11517), .A(n11516), .ZN(P1_U3474) );
  INV_X1 U13280 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n11520) );
  OR2_X1 U13281 ( .A1(n11518), .A2(n16339), .ZN(n11519) );
  OAI21_X1 U13282 ( .B1(n16341), .B2(n11520), .A(n11519), .ZN(P1_U3533) );
  INV_X1 U13283 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n11521) );
  OAI22_X1 U13284 ( .A1(n14464), .A2(n11522), .B1(n11521), .B2(n16242), .ZN(
        n11523) );
  INV_X1 U13285 ( .A(n11523), .ZN(n11524) );
  OAI21_X1 U13286 ( .B1(n11525), .B2(n16239), .A(n11524), .ZN(P3_U3399) );
  NAND2_X1 U13287 ( .A1(n13523), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n11533) );
  NAND2_X1 U13288 ( .A1(n7425), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n11532) );
  INV_X1 U13289 ( .A(n11548), .ZN(n11526) );
  NAND2_X1 U13290 ( .A1(n11526), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n11550) );
  INV_X1 U13291 ( .A(n11550), .ZN(n11527) );
  NAND2_X1 U13292 ( .A1(n11527), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n11677) );
  INV_X1 U13293 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n11528) );
  NAND2_X1 U13294 ( .A1(n11550), .A2(n11528), .ZN(n11529) );
  AND2_X1 U13295 ( .A1(n11677), .A2(n11529), .ZN(n11746) );
  NAND2_X1 U13296 ( .A1(n13522), .A2(n11746), .ZN(n11531) );
  NAND2_X1 U13297 ( .A1(n13517), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n11530) );
  NAND4_X1 U13298 ( .A1(n11533), .A2(n11532), .A3(n11531), .A4(n11530), .ZN(
        n14684) );
  AND2_X1 U13299 ( .A1(n11534), .A2(n13706), .ZN(n11535) );
  NAND2_X1 U13300 ( .A1(n11537), .A2(n14687), .ZN(n11538) );
  NAND2_X1 U13301 ( .A1(n11539), .A2(n12412), .ZN(n11542) );
  AOI22_X1 U13302 ( .A1(n13406), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n13405), 
        .B2(n11540), .ZN(n11541) );
  NAND2_X1 U13303 ( .A1(n11542), .A2(n11541), .ZN(n16122) );
  XNOR2_X1 U13304 ( .A(n16122), .B(n14686), .ZN(n13629) );
  NAND2_X1 U13305 ( .A1(n11543), .A2(n12412), .ZN(n11546) );
  AOI22_X1 U13306 ( .A1(n13406), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n13405), 
        .B2(n11544), .ZN(n11545) );
  NAND2_X1 U13307 ( .A1(n13517), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n11554) );
  NAND2_X1 U13308 ( .A1(n13523), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n11553) );
  INV_X1 U13309 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n11547) );
  NAND2_X1 U13310 ( .A1(n11548), .A2(n11547), .ZN(n11549) );
  AND2_X1 U13311 ( .A1(n11550), .A2(n11549), .ZN(n11605) );
  NAND2_X1 U13312 ( .A1(n12110), .A2(n11605), .ZN(n11552) );
  NAND2_X1 U13313 ( .A1(n7425), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n11551) );
  NAND4_X1 U13314 ( .A1(n11554), .A2(n11553), .A3(n11552), .A4(n11551), .ZN(
        n14685) );
  XNOR2_X1 U13315 ( .A(n13717), .B(n14685), .ZN(n13631) );
  INV_X1 U13316 ( .A(n13631), .ZN(n11687) );
  XNOR2_X1 U13317 ( .A(n11670), .B(n11687), .ZN(n11555) );
  OAI222_X1 U13318 ( .A1(n14914), .A2(n11556), .B1(n14916), .B2(n11911), .C1(
        n14821), .C2(n11555), .ZN(n16143) );
  INV_X1 U13319 ( .A(n16143), .ZN(n11571) );
  NAND2_X1 U13320 ( .A1(n13706), .A2(n14687), .ZN(n11557) );
  NAND2_X1 U13321 ( .A1(n11558), .A2(n11557), .ZN(n11560) );
  OR2_X1 U13322 ( .A1(n14687), .A2(n13706), .ZN(n11559) );
  NAND2_X1 U13323 ( .A1(n11560), .A2(n11559), .ZN(n11776) );
  NAND2_X1 U13324 ( .A1(n11776), .A2(n11781), .ZN(n11562) );
  OR2_X1 U13325 ( .A1(n16122), .A2(n14686), .ZN(n11561) );
  NAND2_X1 U13326 ( .A1(n11562), .A2(n11561), .ZN(n11688) );
  XNOR2_X1 U13327 ( .A(n11688), .B(n11687), .ZN(n16145) );
  NAND2_X1 U13328 ( .A1(n10661), .A2(n11563), .ZN(n11564) );
  NAND2_X1 U13329 ( .A1(n14843), .A2(n11564), .ZN(n14891) );
  INV_X1 U13330 ( .A(n13717), .ZN(n16141) );
  INV_X1 U13331 ( .A(n11685), .ZN(n11565) );
  OAI21_X1 U13332 ( .B1(n16141), .B2(n11778), .A(n11565), .ZN(n16142) );
  INV_X1 U13333 ( .A(n11605), .ZN(n11566) );
  OAI22_X1 U13334 ( .A1(n14843), .A2(n10700), .B1(n11566), .B2(n14840), .ZN(
        n11567) );
  AOI21_X1 U13335 ( .B1(n14849), .B2(n13717), .A(n11567), .ZN(n11568) );
  OAI21_X1 U13336 ( .B1(n14846), .B2(n16142), .A(n11568), .ZN(n11569) );
  AOI21_X1 U13337 ( .B1(n16145), .B2(n14870), .A(n11569), .ZN(n11570) );
  OAI21_X1 U13338 ( .B1(n11571), .B2(n14938), .A(n11570), .ZN(P2_U3258) );
  OAI211_X1 U13339 ( .C1(n11572), .C2(n11574), .A(n11573), .B(n9714), .ZN(
        n11577) );
  NAND2_X1 U13340 ( .A1(n11575), .A2(n14304), .ZN(n11576) );
  AND2_X1 U13341 ( .A1(n11577), .A2(n11576), .ZN(n11635) );
  OR2_X1 U13342 ( .A1(n11579), .A2(n11578), .ZN(n11580) );
  NAND2_X1 U13343 ( .A1(n11581), .A2(n11580), .ZN(n11633) );
  NAND2_X1 U13344 ( .A1(n11633), .A2(n16103), .ZN(n11582) );
  OAI211_X1 U13345 ( .C1(n16055), .C2(n16054), .A(n11635), .B(n11582), .ZN(
        n11793) );
  INV_X1 U13346 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n11583) );
  OAI22_X1 U13347 ( .A1(n14464), .A2(n11727), .B1(n11583), .B2(n16242), .ZN(
        n11584) );
  AOI21_X1 U13348 ( .B1(n11793), .B2(n16242), .A(n11584), .ZN(n11585) );
  INV_X1 U13349 ( .A(n11585), .ZN(P3_U3402) );
  AOI22_X1 U13350 ( .A1(n16265), .A2(n11587), .B1(n11586), .B2(n16262), .ZN(
        n11588) );
  OAI21_X1 U13351 ( .B1(n15416), .B2(n11589), .A(n11588), .ZN(n11592) );
  MUX2_X1 U13352 ( .A(n11590), .B(P1_REG2_REG_5__SCAN_IN), .S(n16264), .Z(
        n11591) );
  AOI211_X1 U13353 ( .C1(n16270), .C2(n11593), .A(n11592), .B(n11591), .ZN(
        n11594) );
  INV_X1 U13354 ( .A(n11594), .ZN(P1_U3288) );
  NAND2_X1 U13355 ( .A1(n14685), .A2(n14552), .ZN(n11738) );
  XNOR2_X1 U13356 ( .A(n13717), .B(n14525), .ZN(n11740) );
  XOR2_X1 U13357 ( .A(n11738), .B(n11740), .Z(n11604) );
  INV_X1 U13358 ( .A(n11595), .ZN(n11598) );
  XNOR2_X1 U13359 ( .A(n16122), .B(n14487), .ZN(n11600) );
  NAND2_X1 U13360 ( .A1(n14686), .A2(n14552), .ZN(n11599) );
  NOR2_X1 U13361 ( .A1(n11600), .A2(n11599), .ZN(n11601) );
  AOI21_X1 U13362 ( .B1(n11600), .B2(n11599), .A(n11601), .ZN(n14645) );
  INV_X1 U13363 ( .A(n11601), .ZN(n11602) );
  AOI21_X1 U13364 ( .B1(n11604), .B2(n11603), .A(n11743), .ZN(n11610) );
  INV_X1 U13365 ( .A(n14661), .ZN(n14648) );
  AOI22_X1 U13366 ( .A1(n14648), .A2(n14686), .B1(n14667), .B2(n11605), .ZN(
        n11607) );
  OAI211_X1 U13367 ( .C1(n11911), .C2(n14663), .A(n11607), .B(n11606), .ZN(
        n11608) );
  AOI21_X1 U13368 ( .B1(n13717), .B2(n14651), .A(n11608), .ZN(n11609) );
  OAI21_X1 U13369 ( .B1(n11610), .B2(n14642), .A(n11609), .ZN(P2_U3185) );
  INV_X1 U13370 ( .A(n11611), .ZN(n11613) );
  OAI222_X1 U13371 ( .A1(P3_U3151), .A2(n11614), .B1(n13924), .B2(n11613), 
        .C1(n11612), .C2(n13926), .ZN(P3_U3275) );
  INV_X1 U13372 ( .A(n11615), .ZN(n11616) );
  AOI21_X1 U13373 ( .B1(n11618), .B2(n11617), .A(n11616), .ZN(n11632) );
  OAI21_X1 U13374 ( .B1(n16027), .B2(n15868), .A(n11619), .ZN(n11625) );
  NAND2_X1 U13375 ( .A1(n11621), .A2(n11620), .ZN(n11622) );
  AOI21_X1 U13376 ( .B1(n11623), .B2(n11622), .A(n16013), .ZN(n11624) );
  AOI211_X1 U13377 ( .C1(n16020), .C2(n11626), .A(n11625), .B(n11624), .ZN(
        n11631) );
  XNOR2_X1 U13378 ( .A(n11628), .B(n11627), .ZN(n11629) );
  NAND2_X1 U13379 ( .A1(n11629), .A2(n16017), .ZN(n11630) );
  OAI211_X1 U13380 ( .C1(n11632), .C2(n16009), .A(n11631), .B(n11630), .ZN(
        P3_U3192) );
  INV_X1 U13381 ( .A(n11633), .ZN(n11639) );
  MUX2_X1 U13382 ( .A(n11635), .B(n11634), .S(n14341), .Z(n11638) );
  OAI22_X1 U13383 ( .A1(n14337), .A2(n11727), .B1(n11725), .B2(n16059), .ZN(
        n11636) );
  AOI21_X1 U13384 ( .B1(n12291), .B2(n14057), .A(n11636), .ZN(n11637) );
  OAI211_X1 U13385 ( .C1(n14288), .C2(n11639), .A(n11638), .B(n11637), .ZN(
        P3_U3229) );
  INV_X1 U13386 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n11652) );
  XOR2_X1 U13387 ( .A(n11642), .B(n11640), .Z(n16117) );
  INV_X1 U13388 ( .A(n16117), .ZN(n11650) );
  XOR2_X1 U13389 ( .A(n11642), .B(n11641), .Z(n11643) );
  NOR2_X1 U13390 ( .A1(n11643), .A2(n16280), .ZN(n11644) );
  AOI211_X1 U13391 ( .C1(n16117), .C2(n16160), .A(n11645), .B(n11644), .ZN(
        n16120) );
  AOI211_X1 U13392 ( .C1(n11648), .C2(n11647), .A(n16198), .B(n11646), .ZN(
        n16116) );
  AOI21_X1 U13393 ( .B1(n16278), .B2(n11648), .A(n16116), .ZN(n11649) );
  OAI211_X1 U13394 ( .C1(n16135), .C2(n11650), .A(n16120), .B(n11649), .ZN(
        n15565) );
  NAND2_X1 U13395 ( .A1(n15565), .A2(n16345), .ZN(n11651) );
  OAI21_X1 U13396 ( .B1(n16345), .B2(n11652), .A(n11651), .ZN(P1_U3477) );
  NAND2_X1 U13397 ( .A1(n11656), .A2(n11655), .ZN(n11661) );
  INV_X1 U13398 ( .A(n15189), .ZN(n11926) );
  OAI22_X1 U13399 ( .A1(n11668), .A2(n13588), .B1(n11926), .B2(n13587), .ZN(
        n11818) );
  NAND2_X1 U13400 ( .A1(n16132), .A2(n13578), .ZN(n11658) );
  NAND2_X1 U13401 ( .A1(n15189), .A2(n13265), .ZN(n11657) );
  NAND2_X1 U13402 ( .A1(n11658), .A2(n11657), .ZN(n11659) );
  XNOR2_X1 U13403 ( .A(n11659), .B(n11815), .ZN(n11817) );
  XOR2_X1 U13404 ( .A(n11818), .B(n11817), .Z(n11660) );
  NAND2_X1 U13405 ( .A1(n11661), .A2(n11660), .ZN(n11821) );
  OAI211_X1 U13406 ( .C1(n11661), .C2(n11660), .A(n11821), .B(n16356), .ZN(
        n11667) );
  INV_X1 U13407 ( .A(n11662), .ZN(n11663) );
  OAI22_X1 U13408 ( .A1(n15132), .A2(n11663), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8732), .ZN(n11664) );
  AOI21_X1 U13409 ( .B1(n15167), .B2(n11665), .A(n11664), .ZN(n11666) );
  OAI211_X1 U13410 ( .C1(n11668), .C2(n16353), .A(n11667), .B(n11666), .ZN(
        P1_U3213) );
  INV_X1 U13411 ( .A(n14685), .ZN(n14649) );
  AND2_X1 U13412 ( .A1(n13717), .A2(n14649), .ZN(n11669) );
  NAND2_X1 U13413 ( .A1(n11671), .A2(n12412), .ZN(n11674) );
  AOI22_X1 U13414 ( .A1(n13406), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n11672), 
        .B2(n13405), .ZN(n11673) );
  NAND2_X1 U13415 ( .A1(n11674), .A2(n11673), .ZN(n13729) );
  XNOR2_X1 U13416 ( .A(n13729), .B(n11911), .ZN(n13633) );
  XNOR2_X1 U13417 ( .A(n11851), .B(n13633), .ZN(n11675) );
  NAND2_X1 U13418 ( .A1(n11675), .A2(n14924), .ZN(n11684) );
  NAND2_X1 U13419 ( .A1(n13523), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n11682) );
  NAND2_X1 U13420 ( .A1(n7425), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n11681) );
  INV_X1 U13421 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n11676) );
  NAND2_X1 U13422 ( .A1(n11677), .A2(n11676), .ZN(n11678) );
  AND2_X1 U13423 ( .A1(n11864), .A2(n11678), .ZN(n11910) );
  NAND2_X1 U13424 ( .A1(n13522), .A2(n11910), .ZN(n11680) );
  NAND2_X1 U13425 ( .A1(n13517), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n11679) );
  NAND4_X1 U13426 ( .A1(n11682), .A2(n11681), .A3(n11680), .A4(n11679), .ZN(
        n14682) );
  AOI22_X1 U13427 ( .A1(n14885), .A2(n14682), .B1(n14685), .B2(n14883), .ZN(
        n11683) );
  NAND2_X1 U13428 ( .A1(n11684), .A2(n11683), .ZN(n16193) );
  MUX2_X1 U13429 ( .A(n16193), .B(P2_REG2_REG_8__SCAN_IN), .S(n14938), .Z(
        n11696) );
  INV_X1 U13430 ( .A(n13729), .ZN(n16189) );
  NAND2_X1 U13431 ( .A1(n11685), .A2(n16189), .ZN(n11891) );
  OR2_X1 U13432 ( .A1(n11685), .A2(n16189), .ZN(n11686) );
  NAND2_X1 U13433 ( .A1(n11891), .A2(n11686), .ZN(n16190) );
  NAND2_X1 U13434 ( .A1(n11688), .A2(n11687), .ZN(n11690) );
  OR2_X1 U13435 ( .A1(n13717), .A2(n14685), .ZN(n11689) );
  INV_X1 U13436 ( .A(n13633), .ZN(n11691) );
  NAND2_X1 U13437 ( .A1(n11692), .A2(n11691), .ZN(n16187) );
  NAND3_X1 U13438 ( .A1(n16188), .A2(n16187), .A3(n14870), .ZN(n11694) );
  AOI22_X1 U13439 ( .A1(n14849), .A2(n13729), .B1(n11746), .B2(n14929), .ZN(
        n11693) );
  OAI211_X1 U13440 ( .C1(n14846), .C2(n16190), .A(n11694), .B(n11693), .ZN(
        n11695) );
  OR2_X1 U13441 ( .A1(n11696), .A2(n11695), .ZN(P2_U3257) );
  INV_X1 U13442 ( .A(n13621), .ZN(n11698) );
  AOI21_X1 U13443 ( .B1(n14902), .B2(n11698), .A(n11697), .ZN(n11700) );
  INV_X1 U13444 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n11699) );
  OAI22_X1 U13445 ( .A1(n14938), .A2(n11700), .B1(n11699), .B2(n14840), .ZN(
        n11701) );
  AOI21_X1 U13446 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n14938), .A(n11701), .ZN(
        n11704) );
  OAI21_X1 U13447 ( .B1(n14849), .B2(n14936), .A(n11702), .ZN(n11703) );
  OAI211_X1 U13448 ( .C1(n14933), .C2(n13621), .A(n11704), .B(n11703), .ZN(
        P2_U3265) );
  INV_X1 U13449 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n16258) );
  AOI22_X1 U13450 ( .A1(n15775), .A2(n16258), .B1(n11707), .B2(n11706), .ZN(
        n11709) );
  INV_X1 U13451 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n16284) );
  MUX2_X1 U13452 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n16284), .S(n12081), .Z(
        n11708) );
  OAI21_X1 U13453 ( .B1(n11709), .B2(n11708), .A(n15776), .ZN(n11720) );
  AOI21_X1 U13454 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n11711), .A(n11710), 
        .ZN(n15773) );
  INV_X1 U13455 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11712) );
  MUX2_X1 U13456 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n11712), .S(n15779), .Z(
        n15774) );
  NAND2_X1 U13457 ( .A1(n15773), .A2(n15774), .ZN(n15772) );
  OAI21_X1 U13458 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n15779), .A(n15772), 
        .ZN(n11714) );
  INV_X1 U13459 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n12085) );
  MUX2_X1 U13460 ( .A(n12085), .B(P1_REG2_REG_13__SCAN_IN), .S(n12081), .Z(
        n11713) );
  NOR2_X1 U13461 ( .A1(n11714), .A2(n11713), .ZN(n12092) );
  AOI211_X1 U13462 ( .C1(n11714), .C2(n11713), .A(n15767), .B(n12092), .ZN(
        n11718) );
  NOR2_X1 U13463 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8665), .ZN(n11715) );
  AOI21_X1 U13464 ( .B1(n15757), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n11715), 
        .ZN(n11716) );
  OAI21_X1 U13465 ( .B1(n15765), .B2(n12086), .A(n11716), .ZN(n11717) );
  NOR2_X1 U13466 ( .A1(n11718), .A2(n11717), .ZN(n11719) );
  OAI21_X1 U13467 ( .B1(n11720), .B2(n12080), .A(n11719), .ZN(P1_U3256) );
  INV_X1 U13468 ( .A(n11721), .ZN(n11722) );
  AOI21_X1 U13469 ( .B1(n11724), .B2(n11723), .A(n11722), .ZN(n11732) );
  INV_X1 U13470 ( .A(n11725), .ZN(n11730) );
  OAI21_X1 U13471 ( .B1(n14017), .B2(n11727), .A(n11726), .ZN(n11729) );
  OAI22_X1 U13472 ( .A1(n11946), .A2(n14032), .B1(n14015), .B2(n16055), .ZN(
        n11728) );
  AOI211_X1 U13473 ( .C1(n11730), .C2(n14023), .A(n11729), .B(n11728), .ZN(
        n11731) );
  OAI21_X1 U13474 ( .B1(n11732), .B2(n14041), .A(n11731), .ZN(P3_U3170) );
  INV_X1 U13475 ( .A(n12507), .ZN(n11736) );
  NAND2_X1 U13476 ( .A1(n11733), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n11734) );
  XNOR2_X1 U13477 ( .A(n11734), .B(P2_IR_REG_16__SCAN_IN), .ZN(n12508) );
  INV_X1 U13478 ( .A(n12508), .ZN(n12342) );
  OAI222_X1 U13479 ( .A1(n13255), .A2(n11735), .B1(n15061), .B2(n11736), .C1(
        n12342), .C2(P2_U3088), .ZN(P2_U3311) );
  INV_X1 U13480 ( .A(n15206), .ZN(n12636) );
  OAI222_X1 U13481 ( .A1(n15597), .A2(n11737), .B1(n15604), .B2(n11736), .C1(
        n12636), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U13482 ( .A(n11738), .ZN(n11739) );
  NOR2_X1 U13483 ( .A1(n11740), .A2(n11739), .ZN(n11742) );
  XNOR2_X1 U13484 ( .A(n13729), .B(n14553), .ZN(n11905) );
  NAND2_X1 U13485 ( .A1(n14684), .A2(n14552), .ZN(n11904) );
  XNOR2_X1 U13486 ( .A(n11905), .B(n11904), .ZN(n11741) );
  NOR3_X1 U13487 ( .A1(n11743), .A2(n11742), .A3(n11741), .ZN(n11744) );
  OAI21_X1 U13488 ( .B1(n7565), .B2(n11744), .A(n14658), .ZN(n11751) );
  INV_X1 U13489 ( .A(n11745), .ZN(n11749) );
  INV_X1 U13490 ( .A(n11746), .ZN(n11747) );
  OAI22_X1 U13491 ( .A1(n14638), .A2(n11747), .B1(n14649), .B2(n14661), .ZN(
        n11748) );
  AOI211_X1 U13492 ( .C1(n14627), .C2(n14682), .A(n11749), .B(n11748), .ZN(
        n11750) );
  OAI211_X1 U13493 ( .C1(n16189), .C2(n14670), .A(n11751), .B(n11750), .ZN(
        P2_U3193) );
  OAI21_X1 U13494 ( .B1(n11753), .B2(n11754), .A(n11752), .ZN(n16104) );
  INV_X1 U13495 ( .A(n16104), .ZN(n11763) );
  AOI21_X1 U13496 ( .B1(n11755), .B2(n11754), .A(n16053), .ZN(n11758) );
  INV_X1 U13497 ( .A(n14054), .ZN(n12260) );
  OAI22_X1 U13498 ( .A1(n12260), .A2(n16056), .B1(n11946), .B2(n16054), .ZN(
        n11756) );
  AOI21_X1 U13499 ( .B1(n11758), .B2(n11757), .A(n11756), .ZN(n16105) );
  MUX2_X1 U13500 ( .A(n16105), .B(n11759), .S(n14341), .Z(n11762) );
  INV_X1 U13501 ( .A(n11951), .ZN(n11760) );
  AOI22_X1 U13502 ( .A1(n16096), .A2(n16101), .B1(n16094), .B2(n11760), .ZN(
        n11761) );
  OAI211_X1 U13503 ( .C1(n14288), .C2(n11763), .A(n11762), .B(n11761), .ZN(
        P3_U3227) );
  INV_X1 U13504 ( .A(n11764), .ZN(n11765) );
  OAI222_X1 U13505 ( .A1(P3_U3151), .A2(n11767), .B1(n13926), .B2(n11766), 
        .C1(n13924), .C2(n11765), .ZN(P3_U3274) );
  INV_X1 U13506 ( .A(n12534), .ZN(n11774) );
  INV_X1 U13507 ( .A(n15216), .ZN(n15222) );
  OAI222_X1 U13508 ( .A1(n15597), .A2(n11768), .B1(n15604), .B2(n11774), .C1(
        P1_U3086), .C2(n15222), .ZN(P1_U3338) );
  OAI21_X1 U13509 ( .B1(n11771), .B2(n11770), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n11772) );
  MUX2_X1 U13510 ( .A(P2_IR_REG_31__SCAN_IN), .B(n11772), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n11773) );
  AND2_X1 U13511 ( .A1(n12233), .A2(n11773), .ZN(n12670) );
  INV_X1 U13512 ( .A(n12670), .ZN(n12451) );
  OAI222_X1 U13513 ( .A1(n13255), .A2(n11775), .B1(n15061), .B2(n11774), .C1(
        P2_U3088), .C2(n12451), .ZN(P2_U3310) );
  XNOR2_X1 U13514 ( .A(n11776), .B(n11781), .ZN(n16121) );
  AND2_X1 U13515 ( .A1(n11777), .A2(n16122), .ZN(n11779) );
  OR2_X1 U13516 ( .A1(n11779), .A2(n11778), .ZN(n16124) );
  AOI22_X1 U13517 ( .A1(n14849), .A2(n16122), .B1(n14929), .B2(n14647), .ZN(
        n11780) );
  OAI21_X1 U13518 ( .B1(n14846), .B2(n16124), .A(n11780), .ZN(n11789) );
  NAND2_X1 U13519 ( .A1(n11782), .A2(n11781), .ZN(n11783) );
  NAND2_X1 U13520 ( .A1(n11784), .A2(n11783), .ZN(n11785) );
  NAND2_X1 U13521 ( .A1(n11785), .A2(n14924), .ZN(n11787) );
  AOI22_X1 U13522 ( .A1(n14883), .A2(n14687), .B1(n14685), .B2(n14885), .ZN(
        n11786) );
  NAND2_X1 U13523 ( .A1(n11787), .A2(n11786), .ZN(n16127) );
  MUX2_X1 U13524 ( .A(n16127), .B(P2_REG2_REG_6__SCAN_IN), .S(n14938), .Z(
        n11788) );
  AOI211_X1 U13525 ( .C1(n14870), .C2(n16121), .A(n11789), .B(n11788), .ZN(
        n11790) );
  INV_X1 U13526 ( .A(n11790), .ZN(P2_U3259) );
  NAND2_X1 U13527 ( .A1(n14055), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n11791) );
  OAI21_X1 U13528 ( .B1(n11792), .B2(n14055), .A(n11791), .ZN(P3_U3521) );
  MUX2_X1 U13529 ( .A(n11793), .B(P3_REG1_REG_4__SCAN_IN), .S(n9764), .Z(
        n11794) );
  AOI21_X1 U13530 ( .B1(n12441), .B2(n7933), .A(n11794), .ZN(n11795) );
  INV_X1 U13531 ( .A(n11795), .ZN(P3_U3463) );
  INV_X1 U13532 ( .A(n11796), .ZN(n11799) );
  OAI22_X1 U13533 ( .A1(n11797), .A2(P3_U3151), .B1(SI_22_), .B2(n13926), .ZN(
        n11798) );
  AOI21_X1 U13534 ( .B1(n11799), .B2(n14474), .A(n11798), .ZN(P3_U3273) );
  OAI21_X1 U13535 ( .B1(n11802), .B2(n11801), .A(n11800), .ZN(n16089) );
  OAI21_X1 U13536 ( .B1(n11805), .B2(n11804), .A(n11803), .ZN(n11807) );
  AOI222_X1 U13537 ( .A1(n9714), .A2(n11807), .B1(n14056), .B2(n14304), .C1(
        n11806), .C2(n14384), .ZN(n16090) );
  INV_X1 U13538 ( .A(n16090), .ZN(n11808) );
  AOI21_X1 U13539 ( .B1(n16103), .B2(n16089), .A(n11808), .ZN(n11814) );
  INV_X1 U13540 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n11809) );
  OAI22_X1 U13541 ( .A1(n14464), .A2(n11810), .B1(n11809), .B2(n16242), .ZN(
        n11811) );
  INV_X1 U13542 ( .A(n11811), .ZN(n11812) );
  OAI21_X1 U13543 ( .B1(n11814), .B2(n16239), .A(n11812), .ZN(P3_U3405) );
  AOI22_X1 U13544 ( .A1(n12441), .A2(n16097), .B1(n9764), .B2(
        P3_REG1_REG_5__SCAN_IN), .ZN(n11813) );
  OAI21_X1 U13545 ( .B1(n11814), .B2(n9764), .A(n11813), .ZN(P3_U3464) );
  INV_X1 U13546 ( .A(n16162), .ZN(n16175) );
  OAI22_X1 U13547 ( .A1(n16175), .A2(n13594), .B1(n11931), .B2(n13588), .ZN(
        n11816) );
  XNOR2_X1 U13548 ( .A(n11816), .B(n11815), .ZN(n11974) );
  OAI22_X1 U13549 ( .A1(n16175), .A2(n13588), .B1(n11931), .B2(n13587), .ZN(
        n11975) );
  XNOR2_X1 U13550 ( .A(n11974), .B(n11975), .ZN(n11823) );
  INV_X1 U13551 ( .A(n11817), .ZN(n11820) );
  INV_X1 U13552 ( .A(n11818), .ZN(n11819) );
  AOI21_X1 U13553 ( .B1(n11823), .B2(n11822), .A(n11978), .ZN(n11830) );
  NAND2_X1 U13554 ( .A1(n15187), .A2(n15457), .ZN(n16161) );
  NAND2_X1 U13555 ( .A1(n15189), .A2(n15455), .ZN(n16153) );
  NAND2_X1 U13556 ( .A1(n16161), .A2(n16153), .ZN(n11824) );
  NAND2_X1 U13557 ( .A1(n15153), .A2(n11824), .ZN(n11825) );
  OAI211_X1 U13558 ( .C1(n16361), .C2(n11827), .A(n11826), .B(n11825), .ZN(
        n11828) );
  AOI21_X1 U13559 ( .B1(n16162), .B2(n15173), .A(n11828), .ZN(n11829) );
  OAI21_X1 U13560 ( .B1(n11830), .B2(n15175), .A(n11829), .ZN(P1_U3221) );
  XNOR2_X1 U13561 ( .A(n11831), .B(n11832), .ZN(n11833) );
  NAND2_X1 U13562 ( .A1(n11833), .A2(n16041), .ZN(n11838) );
  INV_X1 U13563 ( .A(n14056), .ZN(n12051) );
  OAI22_X1 U13564 ( .A1(n11834), .A2(n14015), .B1(n14032), .B2(n12051), .ZN(
        n11835) );
  AOI211_X1 U13565 ( .C1(n16037), .C2(n16097), .A(n11836), .B(n11835), .ZN(
        n11837) );
  OAI211_X1 U13566 ( .C1(n16093), .C2(n14036), .A(n11838), .B(n11837), .ZN(
        P3_U3167) );
  OAI21_X1 U13567 ( .B1(n11840), .B2(n7939), .A(n11839), .ZN(n11993) );
  INV_X1 U13568 ( .A(n11993), .ZN(n11849) );
  INV_X1 U13569 ( .A(n14053), .ZN(n12404) );
  OAI211_X1 U13570 ( .C1(n11843), .C2(n11842), .A(n11841), .B(n9714), .ZN(
        n11844) );
  OAI21_X1 U13571 ( .B1(n12404), .B2(n16056), .A(n11844), .ZN(n11991) );
  NAND2_X1 U13572 ( .A1(n11991), .A2(n16100), .ZN(n11848) );
  NOR2_X1 U13573 ( .A1(n16100), .A2(n9381), .ZN(n11846) );
  OAI22_X1 U13574 ( .A1(n14337), .A2(n11995), .B1(n12056), .B2(n16059), .ZN(
        n11845) );
  AOI211_X1 U13575 ( .C1(n12291), .C2(n14056), .A(n11846), .B(n11845), .ZN(
        n11847) );
  OAI211_X1 U13576 ( .C1(n11849), .C2(n14288), .A(n11848), .B(n11847), .ZN(
        P3_U3226) );
  NAND2_X1 U13577 ( .A1(n13729), .A2(n11911), .ZN(n11850) );
  NAND2_X1 U13578 ( .A1(n11851), .A2(n11850), .ZN(n11853) );
  OR2_X1 U13579 ( .A1(n13729), .A2(n11911), .ZN(n11852) );
  NAND2_X1 U13580 ( .A1(n11853), .A2(n11852), .ZN(n11896) );
  NAND2_X1 U13581 ( .A1(n11854), .A2(n12412), .ZN(n11857) );
  AOI22_X1 U13582 ( .A1(n11855), .A2(n13405), .B1(n13406), .B2(
        P1_DATAO_REG_9__SCAN_IN), .ZN(n11856) );
  INV_X1 U13583 ( .A(n14682), .ZN(n13736) );
  XNOR2_X1 U13584 ( .A(n13734), .B(n13736), .ZN(n13634) );
  INV_X1 U13585 ( .A(n13634), .ZN(n11888) );
  NAND2_X1 U13586 ( .A1(n11896), .A2(n11888), .ZN(n11859) );
  OR2_X1 U13587 ( .A1(n13734), .A2(n13736), .ZN(n11858) );
  NAND2_X1 U13588 ( .A1(n11860), .A2(n12412), .ZN(n11862) );
  AOI22_X1 U13589 ( .A1(n15742), .A2(n13405), .B1(n13406), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n11861) );
  NAND2_X1 U13590 ( .A1(n13523), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n11869) );
  NAND2_X1 U13591 ( .A1(n7425), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n11868) );
  NAND2_X1 U13592 ( .A1(n11864), .A2(n11863), .ZN(n11865) );
  AND2_X1 U13593 ( .A1(n11875), .A2(n11865), .ZN(n12065) );
  NAND2_X1 U13594 ( .A1(n12110), .A2(n12065), .ZN(n11867) );
  NAND2_X1 U13595 ( .A1(n13517), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n11866) );
  NAND4_X1 U13596 ( .A1(n11869), .A2(n11868), .A3(n11867), .A4(n11866), .ZN(
        n14681) );
  INV_X1 U13597 ( .A(n14681), .ZN(n12303) );
  XNOR2_X1 U13598 ( .A(n13747), .B(n12303), .ZN(n13635) );
  XNOR2_X1 U13599 ( .A(n12025), .B(n13635), .ZN(n11883) );
  NAND2_X1 U13600 ( .A1(n13729), .A2(n14684), .ZN(n11870) );
  NAND2_X1 U13601 ( .A1(n11871), .A2(n13635), .ZN(n12019) );
  OR2_X1 U13602 ( .A1(n11871), .A2(n13635), .ZN(n11872) );
  NAND2_X1 U13603 ( .A1(n12019), .A2(n11872), .ZN(n11969) );
  NAND2_X1 U13604 ( .A1(n13517), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n11880) );
  NAND2_X1 U13605 ( .A1(n13523), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n11879) );
  INV_X1 U13606 ( .A(n11875), .ZN(n11873) );
  NAND2_X1 U13607 ( .A1(n11873), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n12031) );
  INV_X1 U13608 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n11874) );
  NAND2_X1 U13609 ( .A1(n11875), .A2(n11874), .ZN(n11876) );
  AND2_X1 U13610 ( .A1(n12031), .A2(n11876), .ZN(n12302) );
  NAND2_X1 U13611 ( .A1(n13522), .A2(n12302), .ZN(n11878) );
  NAND2_X1 U13612 ( .A1(n7425), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n11877) );
  NAND4_X1 U13613 ( .A1(n11880), .A2(n11879), .A3(n11878), .A4(n11877), .ZN(
        n14680) );
  AOI22_X1 U13614 ( .A1(n14883), .A2(n14682), .B1(n14680), .B2(n14885), .ZN(
        n11881) );
  OAI21_X1 U13615 ( .B1(n11969), .B2(n10661), .A(n11881), .ZN(n11882) );
  AOI21_X1 U13616 ( .B1(n11883), .B2(n14924), .A(n11882), .ZN(n11968) );
  AOI21_X1 U13617 ( .B1(n13747), .B2(n11892), .A(n12040), .ZN(n11966) );
  INV_X1 U13618 ( .A(n13747), .ZN(n12070) );
  AOI22_X1 U13619 ( .A1(n14938), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n12065), 
        .B2(n14929), .ZN(n11884) );
  OAI21_X1 U13620 ( .B1(n12070), .B2(n14932), .A(n11884), .ZN(n11886) );
  NOR2_X1 U13621 ( .A1(n11969), .A2(n14933), .ZN(n11885) );
  AOI211_X1 U13622 ( .C1(n11966), .C2(n14936), .A(n11886), .B(n11885), .ZN(
        n11887) );
  OAI21_X1 U13623 ( .B1(n14938), .B2(n11968), .A(n11887), .ZN(P2_U3255) );
  XNOR2_X1 U13624 ( .A(n11889), .B(n11888), .ZN(n16205) );
  AOI21_X1 U13625 ( .B1(n11891), .B2(n13734), .A(n10363), .ZN(n11893) );
  NAND2_X1 U13626 ( .A1(n11893), .A2(n11892), .ZN(n16206) );
  NOR2_X1 U13627 ( .A1(n11894), .A2(n7415), .ZN(n14832) );
  INV_X1 U13628 ( .A(n14832), .ZN(n14733) );
  AOI22_X1 U13629 ( .A1(n14849), .A2(n13734), .B1(n11910), .B2(n14929), .ZN(
        n11895) );
  OAI21_X1 U13630 ( .B1(n16206), .B2(n14733), .A(n11895), .ZN(n11902) );
  XNOR2_X1 U13631 ( .A(n11896), .B(n13634), .ZN(n11897) );
  NAND2_X1 U13632 ( .A1(n11897), .A2(n14924), .ZN(n11900) );
  NAND2_X1 U13633 ( .A1(n16205), .A2(n14902), .ZN(n11899) );
  AOI22_X1 U13634 ( .A1(n14885), .A2(n14681), .B1(n14684), .B2(n14883), .ZN(
        n11898) );
  NAND3_X1 U13635 ( .A1(n11900), .A2(n11899), .A3(n11898), .ZN(n16210) );
  MUX2_X1 U13636 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n16210), .S(n14843), .Z(
        n11901) );
  AOI211_X1 U13637 ( .C1(n14908), .C2(n16205), .A(n11902), .B(n11901), .ZN(
        n11903) );
  INV_X1 U13638 ( .A(n11903), .ZN(P2_U3256) );
  INV_X1 U13639 ( .A(n13734), .ZN(n16208) );
  XNOR2_X1 U13640 ( .A(n13734), .B(n14553), .ZN(n12059) );
  NAND2_X1 U13641 ( .A1(n14682), .A2(n14552), .ZN(n12057) );
  XNOR2_X1 U13642 ( .A(n12059), .B(n12057), .ZN(n11908) );
  INV_X1 U13643 ( .A(n11904), .ZN(n11906) );
  OAI21_X1 U13644 ( .B1(n11908), .B2(n11907), .A(n12061), .ZN(n11909) );
  NAND2_X1 U13645 ( .A1(n11909), .A2(n14658), .ZN(n11916) );
  INV_X1 U13646 ( .A(n11910), .ZN(n11912) );
  OAI22_X1 U13647 ( .A1(n14638), .A2(n11912), .B1(n11911), .B2(n14661), .ZN(
        n11913) );
  AOI211_X1 U13648 ( .C1(n14627), .C2(n14681), .A(n11914), .B(n11913), .ZN(
        n11915) );
  OAI211_X1 U13649 ( .C1(n16208), .C2(n14670), .A(n11916), .B(n11915), .ZN(
        P2_U3203) );
  OR2_X1 U13650 ( .A1(n16132), .A2(n15189), .ZN(n11918) );
  INV_X1 U13651 ( .A(n16157), .ZN(n16149) );
  NAND2_X1 U13652 ( .A1(n16162), .A2(n15188), .ZN(n11919) );
  NAND2_X1 U13653 ( .A1(n16152), .A2(n11919), .ZN(n11922) );
  INV_X1 U13654 ( .A(n11922), .ZN(n11921) );
  NAND2_X1 U13655 ( .A1(n11922), .A2(n11930), .ZN(n11923) );
  NAND2_X1 U13656 ( .A1(n12012), .A2(n11923), .ZN(n16202) );
  INV_X1 U13657 ( .A(n16202), .ZN(n11941) );
  NAND2_X1 U13658 ( .A1(n16132), .A2(n11926), .ZN(n11927) );
  OR2_X1 U13659 ( .A1(n16162), .A2(n11931), .ZN(n11929) );
  XNOR2_X1 U13660 ( .A(n12005), .B(n11930), .ZN(n11934) );
  OAI22_X1 U13661 ( .A1(n11931), .A2(n15406), .B1(n12271), .B2(n15408), .ZN(
        n11932) );
  AOI21_X1 U13662 ( .B1(n16202), .B2(n16160), .A(n11932), .ZN(n11933) );
  OAI21_X1 U13663 ( .B1(n16280), .B2(n11934), .A(n11933), .ZN(n16200) );
  NAND2_X1 U13664 ( .A1(n16200), .A2(n16179), .ZN(n11940) );
  INV_X1 U13665 ( .A(n11935), .ZN(n11985) );
  OAI22_X1 U13666 ( .A1(n16179), .A2(n11936), .B1(n11985), .B2(n16110), .ZN(
        n11938) );
  AND2_X2 U13667 ( .A1(n16163), .A2(n16175), .ZN(n16165) );
  OAI21_X1 U13668 ( .B1(n16197), .B2(n16165), .A(n12000), .ZN(n16199) );
  NOR2_X1 U13669 ( .A1(n16199), .A2(n15416), .ZN(n11937) );
  AOI211_X1 U13670 ( .C1(n16265), .C2(n12010), .A(n11938), .B(n11937), .ZN(
        n11939) );
  OAI211_X1 U13671 ( .C1(n11941), .C2(n15435), .A(n11940), .B(n11939), .ZN(
        P1_U3284) );
  AOI21_X1 U13672 ( .B1(n11943), .B2(n11942), .A(n14041), .ZN(n11945) );
  NAND2_X1 U13673 ( .A1(n11945), .A2(n11944), .ZN(n11950) );
  NAND2_X1 U13674 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n15987) );
  INV_X1 U13675 ( .A(n15987), .ZN(n11948) );
  OAI22_X1 U13676 ( .A1(n12260), .A2(n14032), .B1(n14015), .B2(n11946), .ZN(
        n11947) );
  AOI211_X1 U13677 ( .C1(n16037), .C2(n16101), .A(n11948), .B(n11947), .ZN(
        n11949) );
  OAI211_X1 U13678 ( .C1(n11951), .C2(n14036), .A(n11950), .B(n11949), .ZN(
        P3_U3179) );
  NAND2_X1 U13679 ( .A1(n11952), .A2(n14474), .ZN(n11954) );
  OAI211_X1 U13680 ( .C1(n11955), .C2(n13926), .A(n11954), .B(n11953), .ZN(
        P3_U3272) );
  OAI21_X1 U13681 ( .B1(n11957), .B2(n7568), .A(n11956), .ZN(n11958) );
  AOI22_X1 U13682 ( .A1(n11958), .A2(n9714), .B1(n14304), .B2(n14052), .ZN(
        n12073) );
  OAI21_X1 U13683 ( .B1(n11961), .B2(n11960), .A(n11959), .ZN(n12071) );
  OAI22_X1 U13684 ( .A1(n14337), .A2(n12075), .B1(n7460), .B2(n16059), .ZN(
        n11962) );
  AOI21_X1 U13685 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n14341), .A(n11962), .ZN(
        n11963) );
  OAI21_X1 U13686 ( .B1(n12260), .B2(n14284), .A(n11963), .ZN(n11964) );
  AOI21_X1 U13687 ( .B1(n12071), .B2(n14339), .A(n11964), .ZN(n11965) );
  OAI21_X1 U13688 ( .B1(n12073), .B2(n14341), .A(n11965), .ZN(P3_U3225) );
  AOI22_X1 U13689 ( .A1(n11966), .A2(n15027), .B1(n15026), .B2(n13747), .ZN(
        n11967) );
  OAI211_X1 U13690 ( .C1(n15031), .C2(n11969), .A(n11968), .B(n11967), .ZN(
        n11971) );
  NAND2_X1 U13691 ( .A1(n11971), .A2(n16293), .ZN(n11970) );
  OAI21_X1 U13692 ( .B1(n16293), .B2(n10987), .A(n11970), .ZN(P2_U3509) );
  INV_X1 U13693 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n11973) );
  NAND2_X1 U13694 ( .A1(n11971), .A2(n7419), .ZN(n11972) );
  OAI21_X1 U13695 ( .B1(n7419), .B2(n11973), .A(n11972), .ZN(P2_U3460) );
  INV_X1 U13696 ( .A(n11974), .ZN(n11977) );
  INV_X1 U13697 ( .A(n11975), .ZN(n11976) );
  NAND2_X1 U13698 ( .A1(n12010), .A2(n13578), .ZN(n11980) );
  NAND2_X1 U13699 ( .A1(n15187), .A2(n13265), .ZN(n11979) );
  NAND2_X1 U13700 ( .A1(n11980), .A2(n11979), .ZN(n11981) );
  XNOR2_X1 U13701 ( .A(n11981), .B(n13268), .ZN(n12267) );
  AND2_X1 U13702 ( .A1(n15187), .A2(n13572), .ZN(n11982) );
  AOI21_X1 U13703 ( .B1(n12010), .B2(n13265), .A(n11982), .ZN(n12270) );
  XNOR2_X1 U13704 ( .A(n12267), .B(n12270), .ZN(n11983) );
  OAI211_X1 U13705 ( .C1(n11984), .C2(n11983), .A(n12268), .B(n16356), .ZN(
        n11990) );
  NOR2_X1 U13706 ( .A1(n16361), .A2(n11985), .ZN(n11988) );
  OAI22_X1 U13707 ( .A1(n15170), .A2(n12271), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11986), .ZN(n11987) );
  AOI211_X1 U13708 ( .C1(n16349), .C2(n15188), .A(n11988), .B(n11987), .ZN(
        n11989) );
  OAI211_X1 U13709 ( .C1(n16197), .C2(n16353), .A(n11990), .B(n11989), .ZN(
        P1_U3231) );
  NOR2_X1 U13710 ( .A1(n12051), .A2(n16054), .ZN(n11992) );
  AOI211_X1 U13711 ( .C1(n16103), .C2(n11993), .A(n11992), .B(n11991), .ZN(
        n11999) );
  INV_X1 U13712 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n11994) );
  OAI22_X1 U13713 ( .A1(n14464), .A2(n11995), .B1(n11994), .B2(n16242), .ZN(
        n11996) );
  INV_X1 U13714 ( .A(n11996), .ZN(n11997) );
  OAI21_X1 U13715 ( .B1(n11999), .B2(n16239), .A(n11997), .ZN(P3_U3411) );
  AOI22_X1 U13716 ( .A1(n12441), .A2(n12053), .B1(n9764), .B2(
        P3_REG1_REG_7__SCAN_IN), .ZN(n11998) );
  OAI21_X1 U13717 ( .B1(n11999), .B2(n9764), .A(n11998), .ZN(P3_U3466) );
  NAND2_X1 U13718 ( .A1(n12000), .A2(n12272), .ZN(n12001) );
  NAND2_X1 U13719 ( .A1(n12001), .A2(n16247), .ZN(n12002) );
  OR2_X1 U13720 ( .A1(n7564), .A2(n12002), .ZN(n12004) );
  NAND2_X1 U13721 ( .A1(n15185), .A2(n15457), .ZN(n12003) );
  AND2_X1 U13722 ( .A1(n12004), .A2(n12003), .ZN(n16214) );
  OR2_X1 U13723 ( .A1(n12010), .A2(n12006), .ZN(n12007) );
  XNOR2_X1 U13724 ( .A(n12163), .B(n12167), .ZN(n12009) );
  AOI22_X1 U13725 ( .A1(n12009), .A2(n16330), .B1(n15455), .B2(n15187), .ZN(
        n16215) );
  OAI21_X1 U13726 ( .B1(n7429), .B2(n16214), .A(n16215), .ZN(n12016) );
  XNOR2_X1 U13727 ( .A(n12168), .B(n12167), .ZN(n16218) );
  NAND2_X1 U13728 ( .A1(n16218), .A2(n15366), .ZN(n12014) );
  AOI22_X1 U13729 ( .A1(n16264), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n12281), 
        .B2(n16262), .ZN(n12013) );
  OAI211_X1 U13730 ( .C1(n16216), .C2(n16114), .A(n12014), .B(n12013), .ZN(
        n12015) );
  AOI21_X1 U13731 ( .B1(n16179), .B2(n12016), .A(n12015), .ZN(n12017) );
  INV_X1 U13732 ( .A(n12017), .ZN(P1_U3283) );
  NAND2_X1 U13733 ( .A1(n13747), .A2(n14681), .ZN(n12018) );
  NAND2_X1 U13734 ( .A1(n12019), .A2(n12018), .ZN(n12098) );
  NAND2_X1 U13735 ( .A1(n12020), .A2(n12412), .ZN(n12023) );
  AOI22_X1 U13736 ( .A1(n12021), .A2(n13405), .B1(n13406), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n12022) );
  INV_X1 U13737 ( .A(n14680), .ZN(n12115) );
  XNOR2_X1 U13738 ( .A(n13753), .B(n12115), .ZN(n13637) );
  XNOR2_X1 U13739 ( .A(n12098), .B(n8035), .ZN(n12310) );
  INV_X1 U13740 ( .A(n13635), .ZN(n12024) );
  OR2_X1 U13741 ( .A1(n13747), .A2(n12303), .ZN(n12026) );
  INV_X1 U13742 ( .A(n12119), .ZN(n12116) );
  AOI21_X1 U13743 ( .B1(n13637), .B2(n12028), .A(n12116), .ZN(n12038) );
  NAND2_X1 U13744 ( .A1(n13517), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n12036) );
  NAND2_X1 U13745 ( .A1(n13523), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n12035) );
  INV_X1 U13746 ( .A(n12031), .ZN(n12029) );
  NAND2_X1 U13747 ( .A1(n12029), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n12108) );
  INV_X1 U13748 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n12030) );
  NAND2_X1 U13749 ( .A1(n12031), .A2(n12030), .ZN(n12032) );
  AND2_X1 U13750 ( .A1(n12108), .A2(n12032), .ZN(n12371) );
  NAND2_X1 U13751 ( .A1(n13522), .A2(n12371), .ZN(n12034) );
  NAND2_X1 U13752 ( .A1(n7425), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n12033) );
  NAND4_X1 U13753 ( .A1(n12036), .A2(n12035), .A3(n12034), .A4(n12033), .ZN(
        n14679) );
  AOI22_X1 U13754 ( .A1(n14883), .A2(n14681), .B1(n14679), .B2(n14885), .ZN(
        n12037) );
  OAI21_X1 U13755 ( .B1(n12038), .B2(n14821), .A(n12037), .ZN(n12039) );
  AOI21_X1 U13756 ( .B1(n14902), .B2(n12310), .A(n12039), .ZN(n12313) );
  INV_X1 U13757 ( .A(n13753), .ZN(n12309) );
  INV_X1 U13758 ( .A(n12040), .ZN(n12042) );
  NAND2_X1 U13759 ( .A1(n12309), .A2(n12040), .ZN(n12123) );
  INV_X1 U13760 ( .A(n12123), .ZN(n12041) );
  AOI21_X1 U13761 ( .B1(n13753), .B2(n12042), .A(n12041), .ZN(n12311) );
  NAND2_X1 U13762 ( .A1(n12311), .A2(n14936), .ZN(n12044) );
  AOI22_X1 U13763 ( .A1(n14938), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n12302), 
        .B2(n14929), .ZN(n12043) );
  OAI211_X1 U13764 ( .C1(n12309), .C2(n14932), .A(n12044), .B(n12043), .ZN(
        n12045) );
  AOI21_X1 U13765 ( .B1(n12310), .B2(n14908), .A(n12045), .ZN(n12046) );
  OAI21_X1 U13766 ( .B1(n12313), .B2(n14938), .A(n12046), .ZN(P2_U3254) );
  OAI211_X1 U13767 ( .C1(n12049), .C2(n12048), .A(n12047), .B(n16041), .ZN(
        n12055) );
  INV_X1 U13768 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n12050) );
  NOR2_X1 U13769 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12050), .ZN(n16003) );
  OAI22_X1 U13770 ( .A1(n12051), .A2(n14015), .B1(n14032), .B2(n12404), .ZN(
        n12052) );
  AOI211_X1 U13771 ( .C1(n16037), .C2(n12053), .A(n16003), .B(n12052), .ZN(
        n12054) );
  OAI211_X1 U13772 ( .C1(n12056), .C2(n14036), .A(n12055), .B(n12054), .ZN(
        P3_U3153) );
  XNOR2_X1 U13773 ( .A(n13747), .B(n14553), .ZN(n12296) );
  NAND2_X1 U13774 ( .A1(n14681), .A2(n14552), .ZN(n12294) );
  XNOR2_X1 U13775 ( .A(n12296), .B(n12294), .ZN(n12063) );
  INV_X1 U13776 ( .A(n12057), .ZN(n12058) );
  OAI21_X1 U13777 ( .B1(n12063), .B2(n12062), .A(n12295), .ZN(n12064) );
  NAND2_X1 U13778 ( .A1(n12064), .A2(n14658), .ZN(n12069) );
  AND2_X1 U13779 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n15740) );
  INV_X1 U13780 ( .A(n12065), .ZN(n12066) );
  OAI22_X1 U13781 ( .A1(n14638), .A2(n12066), .B1(n13736), .B2(n14661), .ZN(
        n12067) );
  AOI211_X1 U13782 ( .C1(n14627), .C2(n14680), .A(n15740), .B(n12067), .ZN(
        n12068) );
  OAI211_X1 U13783 ( .C1(n12070), .C2(n14670), .A(n12069), .B(n12068), .ZN(
        P2_U3189) );
  AOI22_X1 U13784 ( .A1(n12071), .A2(n16103), .B1(n14384), .B2(n14054), .ZN(
        n12072) );
  AND2_X1 U13785 ( .A1(n12073), .A2(n12072), .ZN(n12079) );
  INV_X1 U13786 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n12074) );
  OAI22_X1 U13787 ( .A1(n14464), .A2(n12075), .B1(n12074), .B2(n16242), .ZN(
        n12076) );
  INV_X1 U13788 ( .A(n12076), .ZN(n12077) );
  OAI21_X1 U13789 ( .B1(n12079), .B2(n16239), .A(n12077), .ZN(P3_U3414) );
  AOI22_X1 U13790 ( .A1(n12441), .A2(n12263), .B1(n9764), .B2(
        P3_REG1_REG_8__SCAN_IN), .ZN(n12078) );
  OAI21_X1 U13791 ( .B1(n12079), .B2(n9764), .A(n12078), .ZN(P3_U3467) );
  AOI21_X1 U13792 ( .B1(n12081), .B2(P1_REG1_REG_13__SCAN_IN), .A(n12080), 
        .ZN(n12084) );
  INV_X1 U13793 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n12082) );
  MUX2_X1 U13794 ( .A(n12082), .B(P1_REG1_REG_14__SCAN_IN), .S(n12619), .Z(
        n12083) );
  NOR2_X1 U13795 ( .A1(n12084), .A2(n12083), .ZN(n12618) );
  AOI211_X1 U13796 ( .C1(n12084), .C2(n12083), .A(n15240), .B(n12618), .ZN(
        n12097) );
  INV_X1 U13797 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n12626) );
  MUX2_X1 U13798 ( .A(n12626), .B(P1_REG2_REG_14__SCAN_IN), .S(n12619), .Z(
        n12088) );
  NOR2_X1 U13799 ( .A1(n12086), .A2(n12085), .ZN(n12090) );
  INV_X1 U13800 ( .A(n12090), .ZN(n12087) );
  NAND2_X1 U13801 ( .A1(n12088), .A2(n12087), .ZN(n12091) );
  MUX2_X1 U13802 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n12626), .S(n12619), .Z(
        n12089) );
  OAI21_X1 U13803 ( .B1(n12092), .B2(n12090), .A(n12089), .ZN(n12624) );
  OAI211_X1 U13804 ( .C1(n12092), .C2(n12091), .A(n12624), .B(n15780), .ZN(
        n12095) );
  NOR2_X1 U13805 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n15086), .ZN(n12093) );
  AOI21_X1 U13806 ( .B1(n15757), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n12093), 
        .ZN(n12094) );
  OAI211_X1 U13807 ( .C1(n15765), .C2(n12625), .A(n12095), .B(n12094), .ZN(
        n12096) );
  OR2_X1 U13808 ( .A1(n12097), .A2(n12096), .ZN(P1_U3257) );
  NAND2_X1 U13809 ( .A1(n12098), .A2(n13637), .ZN(n12100) );
  NAND2_X1 U13810 ( .A1(n13753), .A2(n14680), .ZN(n12099) );
  NAND2_X1 U13811 ( .A1(n12100), .A2(n12099), .ZN(n12105) );
  NAND2_X1 U13812 ( .A1(n12101), .A2(n12412), .ZN(n12103) );
  AOI22_X1 U13813 ( .A1(n13406), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n13405), 
        .B2(n12243), .ZN(n12102) );
  INV_X1 U13814 ( .A(n14679), .ZN(n13760) );
  OR2_X1 U13815 ( .A1(n13758), .A2(n13760), .ZN(n12186) );
  NAND2_X1 U13816 ( .A1(n13758), .A2(n13760), .ZN(n12104) );
  NAND2_X1 U13817 ( .A1(n12186), .A2(n12104), .ZN(n13638) );
  NAND2_X1 U13818 ( .A1(n12105), .A2(n13638), .ZN(n12182) );
  OR2_X1 U13819 ( .A1(n12105), .A2(n13638), .ZN(n12106) );
  NAND2_X1 U13820 ( .A1(n13517), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n12114) );
  NAND2_X1 U13821 ( .A1(n13523), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n12113) );
  INV_X1 U13822 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n12107) );
  NAND2_X1 U13823 ( .A1(n12108), .A2(n12107), .ZN(n12109) );
  AND2_X1 U13824 ( .A1(n12190), .A2(n12109), .ZN(n12477) );
  NAND2_X1 U13825 ( .A1(n12110), .A2(n12477), .ZN(n12112) );
  NAND2_X1 U13826 ( .A1(n7425), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n12111) );
  NAND4_X1 U13827 ( .A1(n12114), .A2(n12113), .A3(n12112), .A4(n12111), .ZN(
        n14678) );
  OAI22_X1 U13828 ( .A1(n12115), .A2(n14914), .B1(n12587), .B2(n14916), .ZN(
        n12122) );
  AND2_X1 U13829 ( .A1(n13753), .A2(n12115), .ZN(n12117) );
  OAI21_X1 U13830 ( .B1(n12116), .B2(n12117), .A(n13638), .ZN(n12120) );
  NOR2_X1 U13831 ( .A1(n13638), .A2(n12117), .ZN(n12118) );
  AND3_X1 U13832 ( .A1(n12120), .A2(n14924), .A3(n12187), .ZN(n12121) );
  AOI211_X1 U13833 ( .C1(n12352), .C2(n14902), .A(n12122), .B(n12121), .ZN(
        n12355) );
  INV_X1 U13834 ( .A(n13758), .ZN(n12126) );
  INV_X1 U13835 ( .A(n12200), .ZN(n12201) );
  AOI21_X1 U13836 ( .B1(n13758), .B2(n12123), .A(n12201), .ZN(n12353) );
  NAND2_X1 U13837 ( .A1(n12353), .A2(n14936), .ZN(n12125) );
  AOI22_X1 U13838 ( .A1(n14938), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n12371), 
        .B2(n14929), .ZN(n12124) );
  OAI211_X1 U13839 ( .C1(n12126), .C2(n14932), .A(n12125), .B(n12124), .ZN(
        n12127) );
  AOI21_X1 U13840 ( .B1(n12352), .B2(n14908), .A(n12127), .ZN(n12128) );
  OAI21_X1 U13841 ( .B1(n12355), .B2(n14938), .A(n12128), .ZN(P2_U3253) );
  AOI21_X1 U13842 ( .B1(n12130), .B2(n12129), .A(n7561), .ZN(n12146) );
  INV_X1 U13843 ( .A(n12131), .ZN(n12139) );
  INV_X1 U13844 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n12132) );
  NOR2_X1 U13845 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12132), .ZN(n13197) );
  INV_X1 U13846 ( .A(n13197), .ZN(n12133) );
  OAI21_X1 U13847 ( .B1(n16027), .B2(n15890), .A(n12133), .ZN(n12138) );
  AOI211_X1 U13848 ( .C1(n12136), .C2(n12135), .A(n15960), .B(n12134), .ZN(
        n12137) );
  AOI211_X1 U13849 ( .C1(n16020), .C2(n12139), .A(n12138), .B(n12137), .ZN(
        n12145) );
  AOI21_X1 U13850 ( .B1(n12142), .B2(n12141), .A(n12140), .ZN(n12143) );
  OR2_X1 U13851 ( .A1(n12143), .A2(n16009), .ZN(n12144) );
  OAI211_X1 U13852 ( .C1(n12146), .C2(n16013), .A(n12145), .B(n12144), .ZN(
        P3_U3194) );
  AOI21_X1 U13853 ( .B1(n12148), .B2(n12500), .A(n12147), .ZN(n12161) );
  XNOR2_X1 U13854 ( .A(n12150), .B(n12149), .ZN(n12159) );
  INV_X1 U13855 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n12151) );
  NOR2_X1 U13856 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12151), .ZN(n12644) );
  AOI21_X1 U13857 ( .B1(n15646), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n12644), 
        .ZN(n12152) );
  OAI21_X1 U13858 ( .B1(n15997), .B2(n12153), .A(n12152), .ZN(n12158) );
  AOI21_X1 U13859 ( .B1(n9448), .B2(n12155), .A(n12154), .ZN(n12156) );
  NOR2_X1 U13860 ( .A1(n12156), .A2(n16013), .ZN(n12157) );
  AOI211_X1 U13861 ( .C1(n16017), .C2(n12159), .A(n12158), .B(n12157), .ZN(
        n12160) );
  OAI21_X1 U13862 ( .B1(n12161), .B2(n16009), .A(n12160), .ZN(P3_U3193) );
  INV_X1 U13863 ( .A(n12167), .ZN(n12162) );
  NAND2_X1 U13864 ( .A1(n12163), .A2(n12162), .ZN(n12165) );
  OR2_X1 U13865 ( .A1(n12272), .A2(n12271), .ZN(n12164) );
  XNOR2_X1 U13866 ( .A(n12483), .B(n12169), .ZN(n16228) );
  INV_X1 U13867 ( .A(n16228), .ZN(n12180) );
  OAI21_X1 U13868 ( .B1(n12170), .B2(n12169), .A(n12488), .ZN(n16225) );
  INV_X1 U13869 ( .A(n16225), .ZN(n12178) );
  OAI211_X1 U13870 ( .C1(n16224), .C2(n7564), .A(n16247), .B(n16245), .ZN(
        n16223) );
  NAND2_X1 U13871 ( .A1(n15184), .A2(n15457), .ZN(n12172) );
  NAND2_X1 U13872 ( .A1(n15186), .A2(n15455), .ZN(n12171) );
  AND2_X1 U13873 ( .A1(n12172), .A2(n12171), .ZN(n16222) );
  NAND2_X1 U13874 ( .A1(n16264), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n12174) );
  NAND2_X1 U13875 ( .A1(n16262), .A2(n12395), .ZN(n12173) );
  OAI211_X1 U13876 ( .C1(n16264), .C2(n16222), .A(n12174), .B(n12173), .ZN(
        n12175) );
  AOI21_X1 U13877 ( .B1(n12484), .B2(n16265), .A(n12175), .ZN(n12176) );
  OAI21_X1 U13878 ( .B1(n16223), .B2(n16181), .A(n12176), .ZN(n12177) );
  AOI21_X1 U13879 ( .B1(n12178), .B2(n15366), .A(n12177), .ZN(n12179) );
  OAI21_X1 U13880 ( .B1(n15462), .B2(n12180), .A(n12179), .ZN(P1_U3282) );
  NAND2_X1 U13881 ( .A1(n13758), .A2(n14679), .ZN(n12181) );
  NAND2_X1 U13882 ( .A1(n12182), .A2(n12181), .ZN(n12222) );
  NAND2_X1 U13883 ( .A1(n12183), .A2(n12412), .ZN(n12185) );
  AOI22_X1 U13884 ( .A1(n13406), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n13405), 
        .B2(n15717), .ZN(n12184) );
  XNOR2_X1 U13885 ( .A(n13770), .B(n12587), .ZN(n13639) );
  XNOR2_X1 U13886 ( .A(n12222), .B(n13639), .ZN(n12199) );
  XNOR2_X1 U13887 ( .A(n12208), .B(n13639), .ZN(n12197) );
  INV_X1 U13888 ( .A(n12190), .ZN(n12188) );
  NAND2_X1 U13889 ( .A1(n12188), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n12215) );
  INV_X1 U13890 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n12189) );
  NAND2_X1 U13891 ( .A1(n12190), .A2(n12189), .ZN(n12191) );
  NAND2_X1 U13892 ( .A1(n12215), .A2(n12191), .ZN(n12588) );
  OR2_X1 U13893 ( .A1(n13504), .A2(n12588), .ZN(n12195) );
  NAND2_X1 U13894 ( .A1(n13523), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n12194) );
  NAND2_X1 U13895 ( .A1(n13517), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n12193) );
  NAND2_X1 U13896 ( .A1(n7425), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n12192) );
  NAND4_X1 U13897 ( .A1(n12195), .A2(n12194), .A3(n12193), .A4(n12192), .ZN(
        n14677) );
  OAI22_X1 U13898 ( .A1(n13776), .A2(n14916), .B1(n13760), .B2(n14914), .ZN(
        n12196) );
  AOI21_X1 U13899 ( .B1(n12197), .B2(n14924), .A(n12196), .ZN(n12198) );
  OAI21_X1 U13900 ( .B1(n12199), .B2(n10661), .A(n12198), .ZN(n16289) );
  INV_X1 U13901 ( .A(n16289), .ZN(n12206) );
  INV_X1 U13902 ( .A(n12199), .ZN(n16291) );
  INV_X1 U13903 ( .A(n13770), .ZN(n16288) );
  OAI211_X1 U13904 ( .C1(n16288), .C2(n12201), .A(n15027), .B(n12227), .ZN(
        n16287) );
  AOI22_X1 U13905 ( .A1(n14938), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n12477), 
        .B2(n14929), .ZN(n12203) );
  NAND2_X1 U13906 ( .A1(n13770), .A2(n14849), .ZN(n12202) );
  OAI211_X1 U13907 ( .C1(n16287), .C2(n14733), .A(n12203), .B(n12202), .ZN(
        n12204) );
  AOI21_X1 U13908 ( .B1(n16291), .B2(n14908), .A(n12204), .ZN(n12205) );
  OAI21_X1 U13909 ( .B1(n12206), .B2(n14938), .A(n12205), .ZN(P2_U3252) );
  INV_X1 U13910 ( .A(n13639), .ZN(n12207) );
  NAND2_X1 U13911 ( .A1(n12208), .A2(n12207), .ZN(n12210) );
  OR2_X1 U13912 ( .A1(n13770), .A2(n12587), .ZN(n12209) );
  NAND2_X1 U13913 ( .A1(n12211), .A2(n12412), .ZN(n12213) );
  INV_X1 U13914 ( .A(n15680), .ZN(n15689) );
  AOI22_X1 U13915 ( .A1(n13406), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n13405), 
        .B2(n15689), .ZN(n12212) );
  XNOR2_X1 U13916 ( .A(n13774), .B(n13776), .ZN(n13641) );
  XNOR2_X1 U13917 ( .A(n12418), .B(n13641), .ZN(n12221) );
  INV_X1 U13918 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n12214) );
  NAND2_X1 U13919 ( .A1(n12215), .A2(n12214), .ZN(n12216) );
  NAND2_X1 U13920 ( .A1(n12422), .A2(n12216), .ZN(n12613) );
  AOI22_X1 U13921 ( .A1(n13517), .A2(P2_REG0_REG_15__SCAN_IN), .B1(n13523), 
        .B2(P2_REG2_REG_15__SCAN_IN), .ZN(n12218) );
  NAND2_X1 U13922 ( .A1(n7425), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n12217) );
  OAI211_X1 U13923 ( .C1(n12613), .C2(n13504), .A(n12218), .B(n12217), .ZN(
        n14676) );
  NAND2_X1 U13924 ( .A1(n14676), .A2(n14885), .ZN(n12219) );
  OAI21_X1 U13925 ( .B1(n12587), .B2(n14914), .A(n12219), .ZN(n12220) );
  AOI21_X1 U13926 ( .B1(n12221), .B2(n14924), .A(n12220), .ZN(n16312) );
  NAND2_X1 U13927 ( .A1(n12222), .A2(n13639), .ZN(n12224) );
  NAND2_X1 U13928 ( .A1(n13770), .A2(n14678), .ZN(n12223) );
  NAND2_X1 U13929 ( .A1(n12224), .A2(n12223), .ZN(n12225) );
  NAND2_X1 U13930 ( .A1(n12225), .A2(n13641), .ZN(n12411) );
  OR2_X1 U13931 ( .A1(n12225), .A2(n13641), .ZN(n12226) );
  AND2_X1 U13932 ( .A1(n12411), .A2(n12226), .ZN(n16311) );
  NAND2_X1 U13933 ( .A1(n13774), .A2(n12227), .ZN(n12228) );
  NAND2_X1 U13934 ( .A1(n12430), .A2(n12228), .ZN(n16308) );
  INV_X1 U13935 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n12248) );
  OAI22_X1 U13936 ( .A1(n14843), .A2(n12248), .B1(n12588), .B2(n14840), .ZN(
        n12229) );
  AOI21_X1 U13937 ( .B1(n13774), .B2(n14849), .A(n12229), .ZN(n12230) );
  OAI21_X1 U13938 ( .B1(n16308), .B2(n14846), .A(n12230), .ZN(n12231) );
  AOI21_X1 U13939 ( .B1(n16311), .B2(n14870), .A(n12231), .ZN(n12232) );
  OAI21_X1 U13940 ( .B1(n16312), .B2(n14938), .A(n12232), .ZN(P2_U3251) );
  INV_X1 U13941 ( .A(n13398), .ZN(n12236) );
  NAND2_X1 U13942 ( .A1(n12233), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n12234) );
  XNOR2_X1 U13943 ( .A(n12234), .B(P2_IR_REG_18__SCAN_IN), .ZN(n15695) );
  INV_X1 U13944 ( .A(n15695), .ZN(n15702) );
  OAI222_X1 U13945 ( .A1(n13255), .A2(n12235), .B1(n15061), .B2(n12236), .C1(
        n15702), .C2(P2_U3088), .ZN(P2_U3309) );
  INV_X1 U13946 ( .A(n15233), .ZN(n15227) );
  OAI222_X1 U13947 ( .A1(n15597), .A2(n12237), .B1(P1_U3086), .B2(n15227), 
        .C1(n12236), .C2(n15604), .ZN(P1_U3337) );
  OAI21_X1 U13948 ( .B1(n12243), .B2(P2_REG1_REG_12__SCAN_IN), .A(n12238), 
        .ZN(n15729) );
  INV_X1 U13949 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n16292) );
  MUX2_X1 U13950 ( .A(n16292), .B(P2_REG1_REG_13__SCAN_IN), .S(n15717), .Z(
        n15730) );
  NOR2_X1 U13951 ( .A1(n15729), .A2(n15730), .ZN(n15727) );
  AOI21_X1 U13952 ( .B1(n15717), .B2(P2_REG1_REG_13__SCAN_IN), .A(n15727), 
        .ZN(n15687) );
  INV_X1 U13953 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n12240) );
  NAND2_X1 U13954 ( .A1(n15680), .A2(n12240), .ZN(n12239) );
  OAI21_X1 U13955 ( .B1(n15680), .B2(n12240), .A(n12239), .ZN(n15686) );
  NOR2_X1 U13956 ( .A1(n15687), .A2(n15686), .ZN(n15685) );
  AOI21_X1 U13957 ( .B1(n15689), .B2(P2_REG1_REG_14__SCAN_IN), .A(n15685), 
        .ZN(n12338) );
  INV_X1 U13958 ( .A(n12338), .ZN(n12241) );
  XNOR2_X1 U13959 ( .A(n12241), .B(n12414), .ZN(n12336) );
  XOR2_X1 U13960 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n12336), .Z(n12256) );
  NAND2_X1 U13961 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3088), .ZN(n12612)
         );
  OAI21_X1 U13962 ( .B1(n15724), .B2(n12337), .A(n12612), .ZN(n12254) );
  INV_X1 U13963 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n12252) );
  NOR2_X1 U13964 ( .A1(n12248), .A2(n15680), .ZN(n15679) );
  NAND2_X1 U13965 ( .A1(n15717), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n12247) );
  NOR2_X1 U13966 ( .A1(n12243), .A2(n12242), .ZN(n12245) );
  NOR2_X1 U13967 ( .A1(n12245), .A2(n12244), .ZN(n15721) );
  INV_X1 U13968 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n12246) );
  NAND2_X1 U13969 ( .A1(n15725), .A2(n12246), .ZN(n15715) );
  NAND3_X1 U13970 ( .A1(n15721), .A2(n12247), .A3(n15715), .ZN(n15719) );
  NAND2_X1 U13971 ( .A1(n12247), .A2(n15719), .ZN(n15681) );
  OR2_X1 U13972 ( .A1(n15679), .A2(n15681), .ZN(n12250) );
  NAND2_X1 U13973 ( .A1(n15680), .A2(n12248), .ZN(n12249) );
  NAND2_X1 U13974 ( .A1(n12250), .A2(n12249), .ZN(n12343) );
  XNOR2_X1 U13975 ( .A(n12343), .B(n12337), .ZN(n12251) );
  NOR2_X1 U13976 ( .A1(n12251), .A2(n12252), .ZN(n12344) );
  AOI211_X1 U13977 ( .C1(n12252), .C2(n12251), .A(n15736), .B(n12344), .ZN(
        n12253) );
  AOI211_X1 U13978 ( .C1(n15683), .C2(P2_ADDR_REG_15__SCAN_IN), .A(n12254), 
        .B(n12253), .ZN(n12255) );
  OAI21_X1 U13979 ( .B1(n12256), .B2(n15728), .A(n12255), .ZN(P2_U3229) );
  OAI211_X1 U13980 ( .C1(n12259), .C2(n12258), .A(n12257), .B(n16041), .ZN(
        n12265) );
  OAI22_X1 U13981 ( .A1(n12260), .A2(n14015), .B1(n14032), .B2(n12332), .ZN(
        n12261) );
  AOI211_X1 U13982 ( .C1(n16037), .C2(n12263), .A(n12262), .B(n12261), .ZN(
        n12264) );
  OAI211_X1 U13983 ( .C1(n7460), .C2(n14036), .A(n12265), .B(n12264), .ZN(
        P3_U3161) );
  INV_X1 U13984 ( .A(n13404), .ZN(n13251) );
  AND2_X1 U13985 ( .A1(n7415), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13658) );
  AOI21_X1 U13986 ( .B1(P1_DATAO_REG_19__SCAN_IN), .B2(n15059), .A(n13658), 
        .ZN(n12266) );
  OAI21_X1 U13987 ( .B1(n13251), .B2(n15061), .A(n12266), .ZN(P2_U3308) );
  INV_X1 U13988 ( .A(n12267), .ZN(n12269) );
  OAI21_X1 U13989 ( .B1(n12270), .B2(n12269), .A(n12268), .ZN(n12277) );
  OAI22_X1 U13990 ( .A1(n16216), .A2(n13588), .B1(n12271), .B2(n13587), .ZN(
        n12386) );
  NAND2_X1 U13991 ( .A1(n12272), .A2(n13578), .ZN(n12274) );
  NAND2_X1 U13992 ( .A1(n15186), .A2(n13265), .ZN(n12273) );
  NAND2_X1 U13993 ( .A1(n12274), .A2(n12273), .ZN(n12275) );
  XNOR2_X1 U13994 ( .A(n12275), .B(n13268), .ZN(n12385) );
  XOR2_X1 U13995 ( .A(n12386), .B(n12385), .Z(n12276) );
  NAND2_X1 U13996 ( .A1(n12277), .A2(n12276), .ZN(n12389) );
  OAI211_X1 U13997 ( .C1(n12277), .C2(n12276), .A(n12389), .B(n16356), .ZN(
        n12283) );
  NAND2_X1 U13998 ( .A1(n16349), .A2(n15187), .ZN(n12279) );
  OAI211_X1 U13999 ( .C1(n15170), .C2(n12489), .A(n12279), .B(n12278), .ZN(
        n12280) );
  AOI21_X1 U14000 ( .B1(n12281), .B2(n15167), .A(n12280), .ZN(n12282) );
  OAI211_X1 U14001 ( .C1(n16216), .C2(n16353), .A(n12283), .B(n12282), .ZN(
        P1_U3217) );
  NAND2_X1 U14002 ( .A1(n12284), .A2(n9420), .ZN(n12285) );
  NAND2_X1 U14003 ( .A1(n12286), .A2(n12285), .ZN(n12437) );
  INV_X1 U14004 ( .A(n14051), .ZN(n12642) );
  OAI211_X1 U14005 ( .C1(n8368), .C2(n9420), .A(n9714), .B(n12287), .ZN(n12288) );
  OAI21_X1 U14006 ( .B1(n12642), .B2(n16056), .A(n12288), .ZN(n12438) );
  NAND2_X1 U14007 ( .A1(n12438), .A2(n16100), .ZN(n12293) );
  NOR2_X1 U14008 ( .A1(n16100), .A2(n9408), .ZN(n12290) );
  OAI22_X1 U14009 ( .A1(n14337), .A2(n12444), .B1(n12402), .B2(n16059), .ZN(
        n12289) );
  AOI211_X1 U14010 ( .C1(n12291), .C2(n14053), .A(n12290), .B(n12289), .ZN(
        n12292) );
  OAI211_X1 U14011 ( .C1(n14288), .C2(n12437), .A(n12293), .B(n12292), .ZN(
        P3_U3224) );
  XNOR2_X1 U14012 ( .A(n13753), .B(n14553), .ZN(n12364) );
  NAND2_X1 U14013 ( .A1(n14680), .A2(n14552), .ZN(n12362) );
  XNOR2_X1 U14014 ( .A(n12364), .B(n12362), .ZN(n12299) );
  INV_X1 U14015 ( .A(n12294), .ZN(n12297) );
  OAI21_X1 U14016 ( .B1(n12297), .B2(n12296), .A(n12295), .ZN(n12298) );
  OAI21_X1 U14017 ( .B1(n12299), .B2(n12298), .A(n12366), .ZN(n12300) );
  NAND2_X1 U14018 ( .A1(n12300), .A2(n14658), .ZN(n12308) );
  INV_X1 U14019 ( .A(n12301), .ZN(n12306) );
  INV_X1 U14020 ( .A(n12302), .ZN(n12304) );
  OAI22_X1 U14021 ( .A1(n14638), .A2(n12304), .B1(n12303), .B2(n14661), .ZN(
        n12305) );
  AOI211_X1 U14022 ( .C1(n14627), .C2(n14679), .A(n12306), .B(n12305), .ZN(
        n12307) );
  OAI211_X1 U14023 ( .C1(n12309), .C2(n14670), .A(n12308), .B(n12307), .ZN(
        P2_U3208) );
  INV_X1 U14024 ( .A(n12310), .ZN(n12314) );
  AOI22_X1 U14025 ( .A1(n12311), .A2(n15027), .B1(n15026), .B2(n13753), .ZN(
        n12312) );
  OAI211_X1 U14026 ( .C1(n12314), .C2(n15031), .A(n12313), .B(n12312), .ZN(
        n12317) );
  NAND2_X1 U14027 ( .A1(n12317), .A2(n16293), .ZN(n12315) );
  OAI21_X1 U14028 ( .B1(n16293), .B2(n12316), .A(n12315), .ZN(P2_U3510) );
  INV_X1 U14029 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n12319) );
  NAND2_X1 U14030 ( .A1(n12317), .A2(n7419), .ZN(n12318) );
  OAI21_X1 U14031 ( .B1(n7419), .B2(n12319), .A(n12318), .ZN(P2_U3463) );
  OAI211_X1 U14032 ( .C1(n12321), .C2(n12325), .A(n12320), .B(n9714), .ZN(
        n12324) );
  NAND2_X1 U14033 ( .A1(n12322), .A2(n14304), .ZN(n12323) );
  AND2_X1 U14034 ( .A1(n12324), .A2(n12323), .ZN(n12468) );
  NAND2_X1 U14035 ( .A1(n12326), .A2(n12325), .ZN(n12327) );
  NAND2_X1 U14036 ( .A1(n12328), .A2(n12327), .ZN(n12466) );
  OAI22_X1 U14037 ( .A1(n14337), .A2(n12473), .B1(n12329), .B2(n16059), .ZN(
        n12330) );
  AOI21_X1 U14038 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n14341), .A(n12330), 
        .ZN(n12331) );
  OAI21_X1 U14039 ( .B1(n12332), .B2(n14284), .A(n12331), .ZN(n12333) );
  AOI21_X1 U14040 ( .B1(n12466), .B2(n14339), .A(n12333), .ZN(n12334) );
  OAI21_X1 U14041 ( .B1(n12468), .B2(n14341), .A(n12334), .ZN(P3_U3223) );
  INV_X1 U14042 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n12335) );
  OAI22_X1 U14043 ( .A1(n12338), .A2(n12337), .B1(n12336), .B2(n12335), .ZN(
        n12340) );
  XNOR2_X1 U14044 ( .A(n12342), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n12339) );
  NAND2_X1 U14045 ( .A1(n12339), .A2(n12340), .ZN(n12448) );
  OAI211_X1 U14046 ( .C1(n12340), .C2(n12339), .A(n15743), .B(n12448), .ZN(
        n12351) );
  INV_X1 U14047 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n14586) );
  OR2_X1 U14048 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14586), .ZN(n12341) );
  OAI21_X1 U14049 ( .B1(n15724), .B2(n12342), .A(n12341), .ZN(n12349) );
  INV_X1 U14050 ( .A(n12343), .ZN(n12345) );
  AOI21_X1 U14051 ( .B1(n12345), .B2(n12414), .A(n12344), .ZN(n12347) );
  NAND2_X1 U14052 ( .A1(n12508), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n12456) );
  OAI21_X1 U14053 ( .B1(n12508), .B2(P2_REG2_REG_16__SCAN_IN), .A(n12456), 
        .ZN(n12346) );
  NOR2_X1 U14054 ( .A1(n12347), .A2(n12346), .ZN(n12454) );
  AOI211_X1 U14055 ( .C1(n12347), .C2(n12346), .A(n12454), .B(n15736), .ZN(
        n12348) );
  AOI211_X1 U14056 ( .C1(n15683), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n12349), 
        .B(n12348), .ZN(n12350) );
  NAND2_X1 U14057 ( .A1(n12351), .A2(n12350), .ZN(P2_U3230) );
  INV_X1 U14058 ( .A(n12352), .ZN(n12356) );
  AOI22_X1 U14059 ( .A1(n12353), .A2(n15027), .B1(n15026), .B2(n13758), .ZN(
        n12354) );
  OAI211_X1 U14060 ( .C1(n15031), .C2(n12356), .A(n12355), .B(n12354), .ZN(
        n12359) );
  NAND2_X1 U14061 ( .A1(n12359), .A2(n16293), .ZN(n12357) );
  OAI21_X1 U14062 ( .B1(n16293), .B2(n12358), .A(n12357), .ZN(P2_U3511) );
  INV_X1 U14063 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n12361) );
  NAND2_X1 U14064 ( .A1(n12359), .A2(n7419), .ZN(n12360) );
  OAI21_X1 U14065 ( .B1(n7419), .B2(n12361), .A(n12360), .ZN(P2_U3466) );
  INV_X1 U14066 ( .A(n12362), .ZN(n12363) );
  XNOR2_X1 U14067 ( .A(n13758), .B(n14553), .ZN(n12368) );
  AND2_X1 U14068 ( .A1(n14679), .A2(n14552), .ZN(n12367) );
  NOR2_X1 U14069 ( .A1(n12368), .A2(n12367), .ZN(n12475) );
  INV_X1 U14070 ( .A(n12475), .ZN(n12369) );
  NAND2_X1 U14071 ( .A1(n12368), .A2(n12367), .ZN(n12474) );
  NAND2_X1 U14072 ( .A1(n12369), .A2(n12474), .ZN(n12370) );
  XNOR2_X1 U14073 ( .A(n12476), .B(n12370), .ZN(n12376) );
  AOI22_X1 U14074 ( .A1(n14648), .A2(n14680), .B1(n14667), .B2(n12371), .ZN(
        n12373) );
  OAI211_X1 U14075 ( .C1(n12587), .C2(n14663), .A(n12373), .B(n12372), .ZN(
        n12374) );
  AOI21_X1 U14076 ( .B1(n13758), .B2(n14651), .A(n12374), .ZN(n12375) );
  OAI21_X1 U14077 ( .B1(n12376), .B2(n14642), .A(n12375), .ZN(P2_U3196) );
  INV_X1 U14078 ( .A(n12377), .ZN(n12379) );
  OAI222_X1 U14079 ( .A1(n13924), .A2(n12379), .B1(n13926), .B2(n12724), .C1(
        P3_U3151), .C2(n12378), .ZN(P3_U3270) );
  INV_X1 U14080 ( .A(n12380), .ZN(n12382) );
  OAI222_X1 U14081 ( .A1(P3_U3151), .A2(n12383), .B1(n13924), .B2(n12382), 
        .C1(n12381), .C2(n13926), .ZN(P3_U3271) );
  OAI22_X1 U14082 ( .A1(n16224), .A2(n13594), .B1(n12489), .B2(n13588), .ZN(
        n12384) );
  XNOR2_X1 U14083 ( .A(n12384), .B(n13268), .ZN(n12563) );
  OAI22_X1 U14084 ( .A1(n16224), .A2(n13588), .B1(n12489), .B2(n13587), .ZN(
        n12564) );
  XNOR2_X1 U14085 ( .A(n12563), .B(n12564), .ZN(n12391) );
  INV_X1 U14086 ( .A(n12385), .ZN(n12388) );
  INV_X1 U14087 ( .A(n12386), .ZN(n12387) );
  AOI21_X1 U14088 ( .B1(n12391), .B2(n12390), .A(n12567), .ZN(n12397) );
  OAI22_X1 U14089 ( .A1(n15132), .A2(n16222), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12392), .ZN(n12394) );
  NOR2_X1 U14090 ( .A1(n16224), .A2(n16353), .ZN(n12393) );
  AOI211_X1 U14091 ( .C1(n15167), .C2(n12395), .A(n12394), .B(n12393), .ZN(
        n12396) );
  OAI21_X1 U14092 ( .B1(n12397), .B2(n15175), .A(n12396), .ZN(P1_U3236) );
  INV_X1 U14093 ( .A(n12398), .ZN(n12399) );
  AOI21_X1 U14094 ( .B1(n12401), .B2(n12400), .A(n12399), .ZN(n12409) );
  INV_X1 U14095 ( .A(n12402), .ZN(n12407) );
  OR2_X1 U14096 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12403), .ZN(n16025) );
  OAI21_X1 U14097 ( .B1(n14017), .B2(n12444), .A(n16025), .ZN(n12406) );
  OAI22_X1 U14098 ( .A1(n12404), .A2(n14015), .B1(n14032), .B2(n12642), .ZN(
        n12405) );
  AOI211_X1 U14099 ( .C1(n12407), .C2(n14023), .A(n12406), .B(n12405), .ZN(
        n12408) );
  OAI21_X1 U14100 ( .B1(n12409), .B2(n14041), .A(n12408), .ZN(P3_U3171) );
  NAND2_X1 U14101 ( .A1(n13774), .A2(n14677), .ZN(n12410) );
  NAND2_X1 U14102 ( .A1(n12413), .A2(n13615), .ZN(n12416) );
  AOI22_X1 U14103 ( .A1(n13406), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n13405), 
        .B2(n12414), .ZN(n12415) );
  XNOR2_X1 U14104 ( .A(n15025), .B(n14676), .ZN(n13642) );
  XNOR2_X1 U14105 ( .A(n12520), .B(n13642), .ZN(n15024) );
  NAND2_X1 U14106 ( .A1(n13774), .A2(n13776), .ZN(n12417) );
  NAND2_X1 U14107 ( .A1(n12418), .A2(n12417), .ZN(n12420) );
  OR2_X1 U14108 ( .A1(n13774), .A2(n13776), .ZN(n12419) );
  XNOR2_X1 U14109 ( .A(n12506), .B(n13642), .ZN(n12428) );
  INV_X1 U14110 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n12426) );
  NAND2_X1 U14111 ( .A1(n12422), .A2(n14586), .ZN(n12423) );
  NAND2_X1 U14112 ( .A1(n12512), .A2(n12423), .ZN(n14588) );
  OR2_X1 U14113 ( .A1(n14588), .A2(n13504), .ZN(n12425) );
  AOI22_X1 U14114 ( .A1(n13517), .A2(P2_REG0_REG_16__SCAN_IN), .B1(n13523), 
        .B2(P2_REG2_REG_16__SCAN_IN), .ZN(n12424) );
  OAI211_X1 U14115 ( .C1(n13612), .C2(n12426), .A(n12425), .B(n12424), .ZN(
        n14675) );
  AOI22_X1 U14116 ( .A1(n14675), .A2(n14885), .B1(n14883), .B2(n14677), .ZN(
        n12427) );
  OAI21_X1 U14117 ( .B1(n12428), .B2(n14821), .A(n12427), .ZN(n12429) );
  AOI21_X1 U14118 ( .B1(n14902), .B2(n15024), .A(n12429), .ZN(n15030) );
  INV_X1 U14119 ( .A(n15025), .ZN(n12434) );
  AOI21_X1 U14120 ( .B1(n15025), .B2(n12430), .A(n7974), .ZN(n15028) );
  NAND2_X1 U14121 ( .A1(n15028), .A2(n14936), .ZN(n12433) );
  INV_X1 U14122 ( .A(n12613), .ZN(n12431) );
  AOI22_X1 U14123 ( .A1(n14938), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n12431), 
        .B2(n14929), .ZN(n12432) );
  OAI211_X1 U14124 ( .C1(n12434), .C2(n14932), .A(n12433), .B(n12432), .ZN(
        n12435) );
  AOI21_X1 U14125 ( .B1(n15024), .B2(n14908), .A(n12435), .ZN(n12436) );
  OAI21_X1 U14126 ( .B1(n15030), .B2(n14938), .A(n12436), .ZN(P2_U3250) );
  NOR2_X1 U14127 ( .A1(n12437), .A2(n14391), .ZN(n12439) );
  AOI211_X1 U14128 ( .C1(n14384), .C2(n14053), .A(n12439), .B(n12438), .ZN(
        n12447) );
  AOI22_X1 U14129 ( .A1(n12441), .A2(n12440), .B1(n9764), .B2(
        P3_REG1_REG_9__SCAN_IN), .ZN(n12442) );
  OAI21_X1 U14130 ( .B1(n12447), .B2(n9764), .A(n12442), .ZN(P3_U3468) );
  INV_X1 U14131 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n12443) );
  OAI22_X1 U14132 ( .A1(n14464), .A2(n12444), .B1(n12443), .B2(n16242), .ZN(
        n12445) );
  INV_X1 U14133 ( .A(n12445), .ZN(n12446) );
  OAI21_X1 U14134 ( .B1(n12447), .B2(n16239), .A(n12446), .ZN(P3_U3417) );
  NAND2_X1 U14135 ( .A1(n12508), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n12449) );
  NAND2_X1 U14136 ( .A1(n12449), .A2(n12448), .ZN(n12665) );
  INV_X1 U14137 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n12450) );
  XNOR2_X1 U14138 ( .A(n12670), .B(n12450), .ZN(n12664) );
  XNOR2_X1 U14139 ( .A(n12665), .B(n12664), .ZN(n12461) );
  NAND2_X1 U14140 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3088), .ZN(n14596)
         );
  INV_X1 U14141 ( .A(n14596), .ZN(n12453) );
  NOR2_X1 U14142 ( .A1(n15724), .A2(n12451), .ZN(n12452) );
  AOI211_X1 U14143 ( .C1(P2_ADDR_REG_17__SCAN_IN), .C2(n15683), .A(n12453), 
        .B(n12452), .ZN(n12460) );
  INV_X1 U14144 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n12557) );
  XNOR2_X1 U14145 ( .A(n12670), .B(n12557), .ZN(n12458) );
  INV_X1 U14146 ( .A(n12454), .ZN(n12455) );
  NAND2_X1 U14147 ( .A1(n12456), .A2(n12455), .ZN(n12457) );
  NAND2_X1 U14148 ( .A1(n12457), .A2(n12458), .ZN(n12672) );
  OAI211_X1 U14149 ( .C1(n12458), .C2(n12457), .A(n15718), .B(n12672), .ZN(
        n12459) );
  OAI211_X1 U14150 ( .C1(n12461), .C2(n15728), .A(n12460), .B(n12459), .ZN(
        P2_U3231) );
  INV_X1 U14151 ( .A(n12462), .ZN(n12465) );
  OAI222_X1 U14152 ( .A1(n13924), .A2(n12465), .B1(n13926), .B2(n12464), .C1(
        P3_U3151), .C2(n12463), .ZN(P3_U3269) );
  AOI22_X1 U14153 ( .A1(n12466), .A2(n16103), .B1(n14384), .B2(n14052), .ZN(
        n12467) );
  AND2_X1 U14154 ( .A1(n12468), .A2(n12467), .ZN(n12471) );
  INV_X1 U14155 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n12469) );
  MUX2_X1 U14156 ( .A(n12471), .B(n12469), .S(n9764), .Z(n12470) );
  OAI21_X1 U14157 ( .B1(n14418), .B2(n12473), .A(n12470), .ZN(P3_U3469) );
  MUX2_X1 U14158 ( .A(n12471), .B(n9425), .S(n16239), .Z(n12472) );
  OAI21_X1 U14159 ( .B1(n14464), .B2(n12473), .A(n12472), .ZN(P3_U3420) );
  XNOR2_X1 U14160 ( .A(n13770), .B(n14553), .ZN(n12580) );
  NAND2_X1 U14161 ( .A1(n14678), .A2(n14552), .ZN(n12579) );
  XNOR2_X1 U14162 ( .A(n12580), .B(n12579), .ZN(n12582) );
  XNOR2_X1 U14163 ( .A(n12583), .B(n12582), .ZN(n12481) );
  AOI22_X1 U14164 ( .A1(n14648), .A2(n14679), .B1(n14667), .B2(n12477), .ZN(
        n12478) );
  NAND2_X1 U14165 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n15722)
         );
  OAI211_X1 U14166 ( .C1(n13776), .C2(n14663), .A(n12478), .B(n15722), .ZN(
        n12479) );
  AOI21_X1 U14167 ( .B1(n13770), .B2(n14651), .A(n12479), .ZN(n12480) );
  OAI21_X1 U14168 ( .B1(n12481), .B2(n14642), .A(n12480), .ZN(P2_U3206) );
  NOR2_X1 U14169 ( .A1(n12484), .A2(n12489), .ZN(n12482) );
  OR2_X1 U14170 ( .A1(n16266), .A2(n12687), .ZN(n12487) );
  XNOR2_X1 U14171 ( .A(n12649), .B(n12659), .ZN(n16281) );
  XNOR2_X1 U14172 ( .A(n7567), .B(n12659), .ZN(n16283) );
  NAND2_X1 U14173 ( .A1(n16283), .A2(n15366), .ZN(n12494) );
  XNOR2_X1 U14174 ( .A(n16277), .B(n16246), .ZN(n12490) );
  OAI222_X1 U14175 ( .A1(n16198), .A2(n12490), .B1(n15406), .B2(n12687), .C1(
        n15408), .C2(n12699), .ZN(n16276) );
  AOI22_X1 U14176 ( .A1(n16264), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n12690), 
        .B2(n16262), .ZN(n12491) );
  OAI21_X1 U14177 ( .B1(n12693), .B2(n16114), .A(n12491), .ZN(n12492) );
  AOI21_X1 U14178 ( .B1(n16276), .B2(n16269), .A(n12492), .ZN(n12493) );
  OAI211_X1 U14179 ( .C1(n16281), .C2(n15462), .A(n12494), .B(n12493), .ZN(
        P1_U3280) );
  XNOR2_X1 U14180 ( .A(n12495), .B(n12498), .ZN(n12496) );
  AOI222_X1 U14181 ( .A1(n9714), .A2(n12496), .B1(n14050), .B2(n14304), .C1(
        n14051), .C2(n14384), .ZN(n12715) );
  OAI21_X1 U14182 ( .B1(n12499), .B2(n12498), .A(n12497), .ZN(n12713) );
  NOR2_X1 U14183 ( .A1(n16100), .A2(n12500), .ZN(n12503) );
  OAI22_X1 U14184 ( .A1(n14337), .A2(n12501), .B1(n12647), .B2(n16059), .ZN(
        n12502) );
  AOI211_X1 U14185 ( .C1(n12713), .C2(n14339), .A(n12503), .B(n12502), .ZN(
        n12504) );
  OAI21_X1 U14186 ( .B1(n12715), .B2(n14341), .A(n12504), .ZN(P3_U3222) );
  INV_X1 U14187 ( .A(n14676), .ZN(n14587) );
  NOR2_X1 U14188 ( .A1(n15025), .A2(n14587), .ZN(n12505) );
  NAND2_X1 U14189 ( .A1(n12507), .A2(n13615), .ZN(n12510) );
  AOI22_X1 U14190 ( .A1(n13406), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n12508), 
        .B2(n13405), .ZN(n12509) );
  XNOR2_X1 U14191 ( .A(n15017), .B(n14675), .ZN(n13643) );
  XNOR2_X1 U14192 ( .A(n12533), .B(n13643), .ZN(n12516) );
  INV_X1 U14193 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n12511) );
  NAND2_X1 U14194 ( .A1(n12512), .A2(n12511), .ZN(n12513) );
  NAND2_X1 U14195 ( .A1(n12540), .A2(n12513), .ZN(n14598) );
  AOI22_X1 U14196 ( .A1(n7425), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n13523), 
        .B2(P2_REG2_REG_17__SCAN_IN), .ZN(n12515) );
  NAND2_X1 U14197 ( .A1(n13517), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n12514) );
  OAI211_X1 U14198 ( .C1(n14598), .C2(n13504), .A(n12515), .B(n12514), .ZN(
        n14674) );
  AOI222_X1 U14199 ( .A1(n14924), .A2(n12516), .B1(n14674), .B2(n14885), .C1(
        n14676), .C2(n14883), .ZN(n15023) );
  XOR2_X1 U14200 ( .A(n12554), .B(n15017), .Z(n15018) );
  INV_X1 U14201 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n12517) );
  OAI22_X1 U14202 ( .A1(n14843), .A2(n12517), .B1(n14588), .B2(n14840), .ZN(
        n12519) );
  NOR2_X1 U14203 ( .A1(n7973), .A2(n14932), .ZN(n12518) );
  AOI211_X1 U14204 ( .C1(n15018), .C2(n14936), .A(n12519), .B(n12518), .ZN(
        n12525) );
  OR2_X1 U14205 ( .A1(n15025), .A2(n14676), .ZN(n12521) );
  NAND2_X1 U14206 ( .A1(n12523), .A2(n13643), .ZN(n15019) );
  NAND3_X1 U14207 ( .A1(n7629), .A2(n15019), .A3(n14870), .ZN(n12524) );
  OAI211_X1 U14208 ( .C1(n15023), .C2(n14938), .A(n12525), .B(n12524), .ZN(
        P2_U3249) );
  INV_X1 U14209 ( .A(n13417), .ZN(n12531) );
  OAI222_X1 U14210 ( .A1(P1_U3086), .A2(n12527), .B1(n15604), .B2(n12531), 
        .C1(n12526), .C2(n15597), .ZN(P1_U3335) );
  INV_X1 U14211 ( .A(n12528), .ZN(n12530) );
  INV_X1 U14212 ( .A(SI_27_), .ZN(n12529) );
  OAI222_X1 U14213 ( .A1(n13924), .A2(n12530), .B1(n13926), .B2(n12529), .C1(
        P3_U3151), .C2(n14141), .ZN(P3_U3268) );
  OAI222_X1 U14214 ( .A1(n13255), .A2(n13418), .B1(P2_U3088), .B2(n13912), 
        .C1(n15061), .C2(n12531), .ZN(P2_U3307) );
  INV_X1 U14215 ( .A(n14675), .ZN(n14597) );
  AND2_X1 U14216 ( .A1(n15017), .A2(n14597), .ZN(n12532) );
  NAND2_X1 U14217 ( .A1(n12534), .A2(n13615), .ZN(n12536) );
  AOI22_X1 U14218 ( .A1(n13406), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n13405), 
        .B2(n12670), .ZN(n12535) );
  OR2_X1 U14219 ( .A1(n15011), .A2(n14674), .ZN(n13533) );
  NAND2_X1 U14220 ( .A1(n15011), .A2(n14674), .ZN(n12537) );
  NAND2_X1 U14221 ( .A1(n13533), .A2(n12537), .ZN(n13645) );
  XNOR2_X1 U14222 ( .A(n13403), .B(n8152), .ZN(n12538) );
  NAND2_X1 U14223 ( .A1(n12538), .A2(n14924), .ZN(n12550) );
  INV_X1 U14224 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n14637) );
  NAND2_X1 U14225 ( .A1(n12540), .A2(n14637), .ZN(n12541) );
  NAND2_X1 U14226 ( .A1(n13423), .A2(n12541), .ZN(n14928) );
  OR2_X1 U14227 ( .A1(n14928), .A2(n13504), .ZN(n12548) );
  INV_X1 U14228 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n12544) );
  NAND2_X1 U14229 ( .A1(n13517), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n12543) );
  NAND2_X1 U14230 ( .A1(n7425), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n12542) );
  OAI211_X1 U14231 ( .C1(n12545), .C2(n12544), .A(n12543), .B(n12542), .ZN(
        n12546) );
  INV_X1 U14232 ( .A(n12546), .ZN(n12547) );
  NAND2_X1 U14233 ( .A1(n12548), .A2(n12547), .ZN(n14673) );
  AOI22_X1 U14234 ( .A1(n14673), .A2(n14885), .B1(n14883), .B2(n14675), .ZN(
        n12549) );
  NAND2_X1 U14235 ( .A1(n12550), .A2(n12549), .ZN(n15015) );
  INV_X1 U14236 ( .A(n15015), .ZN(n12562) );
  NAND2_X1 U14237 ( .A1(n15017), .A2(n14675), .ZN(n12551) );
  NAND2_X1 U14238 ( .A1(n12552), .A2(n13645), .ZN(n12553) );
  NAND2_X1 U14239 ( .A1(n13534), .A2(n12553), .ZN(n15010) );
  INV_X1 U14240 ( .A(n13530), .ZN(n14927) );
  NAND2_X1 U14241 ( .A1(n15011), .A2(n12555), .ZN(n12556) );
  NAND2_X1 U14242 ( .A1(n14927), .A2(n12556), .ZN(n15013) );
  OAI22_X1 U14243 ( .A1(n14843), .A2(n12557), .B1(n14598), .B2(n14840), .ZN(
        n12558) );
  AOI21_X1 U14244 ( .B1(n15011), .B2(n14849), .A(n12558), .ZN(n12559) );
  OAI21_X1 U14245 ( .B1(n15013), .B2(n14846), .A(n12559), .ZN(n12560) );
  AOI21_X1 U14246 ( .B1(n15010), .B2(n14870), .A(n12560), .ZN(n12561) );
  OAI21_X1 U14247 ( .B1(n12562), .B2(n14938), .A(n12561), .ZN(P2_U3248) );
  INV_X1 U14248 ( .A(n12563), .ZN(n12566) );
  INV_X1 U14249 ( .A(n12564), .ZN(n12565) );
  OAI22_X1 U14250 ( .A1(n16249), .A2(n13594), .B1(n12687), .B2(n13588), .ZN(
        n12568) );
  XNOR2_X1 U14251 ( .A(n12568), .B(n13268), .ZN(n12677) );
  AND2_X1 U14252 ( .A1(n15184), .A2(n13572), .ZN(n12569) );
  AOI21_X1 U14253 ( .B1(n16266), .B2(n13265), .A(n12569), .ZN(n12680) );
  XNOR2_X1 U14254 ( .A(n12677), .B(n12680), .ZN(n12570) );
  OAI211_X1 U14255 ( .C1(n12571), .C2(n12570), .A(n12678), .B(n16356), .ZN(
        n12576) );
  NAND2_X1 U14256 ( .A1(n15183), .A2(n15457), .ZN(n12573) );
  NAND2_X1 U14257 ( .A1(n15185), .A2(n15455), .ZN(n12572) );
  AND2_X1 U14258 ( .A1(n12573), .A2(n12572), .ZN(n16253) );
  NAND2_X1 U14259 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n15782)
         );
  OAI21_X1 U14260 ( .B1(n15132), .B2(n16253), .A(n15782), .ZN(n12574) );
  AOI21_X1 U14261 ( .B1(n15167), .B2(n16263), .A(n12574), .ZN(n12575) );
  OAI211_X1 U14262 ( .C1(n16249), .C2(n16353), .A(n12576), .B(n12575), .ZN(
        P1_U3224) );
  AND2_X1 U14263 ( .A1(n14677), .A2(n14552), .ZN(n12578) );
  XNOR2_X1 U14264 ( .A(n13774), .B(n14553), .ZN(n12577) );
  NOR2_X1 U14265 ( .A1(n12577), .A2(n12578), .ZN(n12610) );
  AOI21_X1 U14266 ( .B1(n12578), .B2(n12577), .A(n12610), .ZN(n12585) );
  INV_X1 U14267 ( .A(n12579), .ZN(n12581) );
  OAI21_X1 U14268 ( .B1(n12585), .B2(n12584), .A(n12611), .ZN(n12586) );
  NAND2_X1 U14269 ( .A1(n12586), .A2(n14658), .ZN(n12592) );
  NAND2_X1 U14270 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n15692)
         );
  INV_X1 U14271 ( .A(n15692), .ZN(n12590) );
  OAI22_X1 U14272 ( .A1(n14638), .A2(n12588), .B1(n12587), .B2(n14661), .ZN(
        n12589) );
  AOI211_X1 U14273 ( .C1(n14627), .C2(n14676), .A(n12590), .B(n12589), .ZN(
        n12591) );
  OAI211_X1 U14274 ( .C1(n7975), .C2(n14670), .A(n12592), .B(n12591), .ZN(
        P2_U3187) );
  INV_X1 U14275 ( .A(n13432), .ZN(n12595) );
  OAI222_X1 U14276 ( .A1(n15597), .A2(n12594), .B1(n15604), .B2(n12595), .C1(
        P1_U3086), .C2(n12593), .ZN(P1_U3334) );
  OAI222_X1 U14277 ( .A1(n13255), .A2(n13433), .B1(n15061), .B2(n12595), .C1(
        n13899), .C2(P2_U3088), .ZN(P2_U3306) );
  OAI21_X1 U14278 ( .B1(n12596), .B2(n12600), .A(n13178), .ZN(n16235) );
  INV_X1 U14279 ( .A(n16235), .ZN(n12609) );
  INV_X1 U14280 ( .A(n12597), .ZN(n12598) );
  NAND2_X1 U14281 ( .A1(n16100), .A2(n12598), .ZN(n14263) );
  XOR2_X1 U14282 ( .A(n12600), .B(n12599), .Z(n12605) );
  INV_X1 U14283 ( .A(n14256), .ZN(n12603) );
  OAI22_X1 U14284 ( .A1(n13200), .A2(n16054), .B1(n12601), .B2(n16056), .ZN(
        n12602) );
  AOI21_X1 U14285 ( .B1(n16235), .B2(n12603), .A(n12602), .ZN(n12604) );
  OAI21_X1 U14286 ( .B1(n12605), .B2(n16053), .A(n12604), .ZN(n16233) );
  NAND2_X1 U14287 ( .A1(n16233), .A2(n16100), .ZN(n12608) );
  OAI22_X1 U14288 ( .A1(n14337), .A2(n16232), .B1(n13198), .B2(n16059), .ZN(
        n12606) );
  AOI21_X1 U14289 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n14341), .A(n12606), 
        .ZN(n12607) );
  OAI211_X1 U14290 ( .C1(n12609), .C2(n14263), .A(n12608), .B(n12607), .ZN(
        P3_U3221) );
  NAND2_X1 U14291 ( .A1(n14676), .A2(n14552), .ZN(n14479) );
  XNOR2_X1 U14292 ( .A(n15025), .B(n14553), .ZN(n14478) );
  XOR2_X1 U14293 ( .A(n14479), .B(n14478), .Z(n14481) );
  XNOR2_X1 U14294 ( .A(n14482), .B(n14481), .ZN(n12617) );
  OAI21_X1 U14295 ( .B1(n14663), .B2(n14597), .A(n12612), .ZN(n12615) );
  OAI22_X1 U14296 ( .A1(n14638), .A2(n12613), .B1(n13776), .B2(n14661), .ZN(
        n12614) );
  AOI211_X1 U14297 ( .C1(n15025), .C2(n14651), .A(n12615), .B(n12614), .ZN(
        n12616) );
  OAI21_X1 U14298 ( .B1(n12617), .B2(n14642), .A(n12616), .ZN(P2_U3213) );
  INV_X1 U14299 ( .A(n12620), .ZN(n12621) );
  INV_X1 U14300 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n16340) );
  XNOR2_X1 U14301 ( .A(n15206), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n12622) );
  NOR2_X1 U14302 ( .A1(n12622), .A2(n12623), .ZN(n15205) );
  AOI211_X1 U14303 ( .C1(n12623), .C2(n12622), .A(n15205), .B(n15240), .ZN(
        n12638) );
  OAI21_X1 U14304 ( .B1(n12626), .B2(n12625), .A(n12624), .ZN(n12628) );
  INV_X1 U14305 ( .A(n12628), .ZN(n12629) );
  XNOR2_X1 U14306 ( .A(n12628), .B(n12627), .ZN(n15764) );
  NOR2_X1 U14307 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n15764), .ZN(n15763) );
  AOI21_X1 U14308 ( .B1(n12629), .B2(n15766), .A(n15763), .ZN(n12632) );
  NAND2_X1 U14309 ( .A1(n15206), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n15199) );
  INV_X1 U14310 ( .A(n15199), .ZN(n12630) );
  AOI21_X1 U14311 ( .B1(n8618), .B2(n12636), .A(n12630), .ZN(n12631) );
  NAND2_X1 U14312 ( .A1(n12631), .A2(n12632), .ZN(n15198) );
  OAI211_X1 U14313 ( .C1(n12632), .C2(n12631), .A(n15780), .B(n15198), .ZN(
        n12635) );
  NAND2_X1 U14314 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n16358)
         );
  INV_X1 U14315 ( .A(n16358), .ZN(n12633) );
  AOI21_X1 U14316 ( .B1(n15757), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n12633), 
        .ZN(n12634) );
  OAI211_X1 U14317 ( .C1(n15765), .C2(n12636), .A(n12635), .B(n12634), .ZN(
        n12637) );
  OR2_X1 U14318 ( .A1(n12638), .A2(n12637), .ZN(P1_U3259) );
  OAI211_X1 U14319 ( .C1(n12641), .C2(n12640), .A(n12639), .B(n16041), .ZN(
        n12646) );
  OAI22_X1 U14320 ( .A1(n12642), .A2(n14015), .B1(n14032), .B2(n13230), .ZN(
        n12643) );
  AOI211_X1 U14321 ( .C1(n16037), .C2(n12712), .A(n12644), .B(n12643), .ZN(
        n12645) );
  OAI211_X1 U14322 ( .C1(n12647), .C2(n14036), .A(n12646), .B(n12645), .ZN(
        P3_U3176) );
  INV_X1 U14323 ( .A(n15462), .ZN(n15418) );
  XNOR2_X1 U14324 ( .A(n12698), .B(n12697), .ZN(n16304) );
  INV_X1 U14325 ( .A(n15089), .ZN(n16298) );
  OR2_X1 U14326 ( .A1(n16277), .A2(n16246), .ZN(n12651) );
  INV_X1 U14327 ( .A(n12651), .ZN(n12652) );
  OAI211_X1 U14328 ( .C1(n16298), .C2(n12652), .A(n16247), .B(n12695), .ZN(
        n16297) );
  NAND2_X1 U14329 ( .A1(n16348), .A2(n15457), .ZN(n12654) );
  NAND2_X1 U14330 ( .A1(n15183), .A2(n15455), .ZN(n12653) );
  AND2_X1 U14331 ( .A1(n12654), .A2(n12653), .ZN(n16296) );
  INV_X1 U14332 ( .A(n15088), .ZN(n12655) );
  OAI22_X1 U14333 ( .A1(n16264), .A2(n16296), .B1(n12655), .B2(n16110), .ZN(
        n12657) );
  NOR2_X1 U14334 ( .A1(n16298), .A2(n16114), .ZN(n12656) );
  AOI211_X1 U14335 ( .C1(n16264), .C2(P1_REG2_REG_14__SCAN_IN), .A(n12657), 
        .B(n12656), .ZN(n12658) );
  OAI21_X1 U14336 ( .B1(n16181), .B2(n16297), .A(n12658), .ZN(n12662) );
  AND2_X1 U14337 ( .A1(n12660), .A2(n12697), .ZN(n16300) );
  NOR3_X1 U14338 ( .A1(n16301), .A2(n16300), .A3(n15466), .ZN(n12661) );
  AOI211_X1 U14339 ( .C1(n15418), .C2(n16304), .A(n12662), .B(n12661), .ZN(
        n12663) );
  INV_X1 U14340 ( .A(n12663), .ZN(P1_U3279) );
  NAND2_X1 U14341 ( .A1(n12665), .A2(n12664), .ZN(n12667) );
  NAND2_X1 U14342 ( .A1(n12670), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n12666) );
  NAND2_X1 U14343 ( .A1(n12667), .A2(n12666), .ZN(n15701) );
  XNOR2_X1 U14344 ( .A(n15701), .B(n15695), .ZN(n15705) );
  XOR2_X1 U14345 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n15705), .Z(n12676) );
  NOR2_X1 U14346 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14637), .ZN(n12669) );
  NOR2_X1 U14347 ( .A1(n15724), .A2(n15702), .ZN(n12668) );
  AOI211_X1 U14348 ( .C1(P2_ADDR_REG_18__SCAN_IN), .C2(n15683), .A(n12669), 
        .B(n12668), .ZN(n12675) );
  NAND2_X1 U14349 ( .A1(n12670), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n12671) );
  NAND2_X1 U14350 ( .A1(n12672), .A2(n12671), .ZN(n15694) );
  XNOR2_X1 U14351 ( .A(n15694), .B(n15695), .ZN(n15696) );
  XNOR2_X1 U14352 ( .A(n15696), .B(P2_REG2_REG_18__SCAN_IN), .ZN(n12673) );
  NAND2_X1 U14353 ( .A1(n12673), .A2(n15718), .ZN(n12674) );
  OAI211_X1 U14354 ( .C1(n12676), .C2(n15728), .A(n12675), .B(n12674), .ZN(
        P2_U3232) );
  INV_X1 U14355 ( .A(n12677), .ZN(n12679) );
  OAI21_X1 U14356 ( .B1(n12680), .B2(n12679), .A(n12678), .ZN(n12686) );
  OAI22_X1 U14357 ( .A1(n12693), .A2(n13588), .B1(n12681), .B2(n13587), .ZN(
        n13261) );
  NAND2_X1 U14358 ( .A1(n16277), .A2(n13578), .ZN(n12683) );
  NAND2_X1 U14359 ( .A1(n15183), .A2(n13265), .ZN(n12682) );
  NAND2_X1 U14360 ( .A1(n12683), .A2(n12682), .ZN(n12684) );
  XNOR2_X1 U14361 ( .A(n12684), .B(n13268), .ZN(n13260) );
  XOR2_X1 U14362 ( .A(n13261), .B(n13260), .Z(n12685) );
  OAI211_X1 U14363 ( .C1(n12686), .C2(n12685), .A(n13264), .B(n16356), .ZN(
        n12692) );
  OAI22_X1 U14364 ( .A1(n15170), .A2(n12699), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8665), .ZN(n12689) );
  NOR2_X1 U14365 ( .A1(n15159), .A2(n12687), .ZN(n12688) );
  AOI211_X1 U14366 ( .C1(n15167), .C2(n12690), .A(n12689), .B(n12688), .ZN(
        n12691) );
  OAI211_X1 U14367 ( .C1(n12693), .C2(n16353), .A(n12692), .B(n12691), .ZN(
        P1_U3234) );
  NAND2_X1 U14368 ( .A1(n12694), .A2(n12702), .ZN(n13331) );
  OAI21_X1 U14369 ( .B1(n12694), .B2(n12702), .A(n13331), .ZN(n16338) );
  AOI21_X1 U14370 ( .B1(n13354), .B2(n12695), .A(n16198), .ZN(n12696) );
  NAND2_X1 U14371 ( .A1(n12696), .A2(n15453), .ZN(n16332) );
  NAND2_X1 U14372 ( .A1(n12698), .A2(n12697), .ZN(n12701) );
  NAND2_X1 U14373 ( .A1(n15089), .A2(n12699), .ZN(n12700) );
  NAND2_X1 U14374 ( .A1(n12703), .A2(n12702), .ZN(n16329) );
  NAND3_X1 U14375 ( .A1(n13356), .A2(n16329), .A3(n15418), .ZN(n12709) );
  NAND2_X1 U14376 ( .A1(n16322), .A2(n15457), .ZN(n12705) );
  NAND2_X1 U14377 ( .A1(n16321), .A2(n15455), .ZN(n12704) );
  AND2_X1 U14378 ( .A1(n12705), .A2(n12704), .ZN(n16331) );
  OAI22_X1 U14379 ( .A1(n16264), .A2(n16331), .B1(n16328), .B2(n16110), .ZN(
        n12707) );
  INV_X1 U14380 ( .A(n13354), .ZN(n16334) );
  NOR2_X1 U14381 ( .A1(n16334), .A2(n16114), .ZN(n12706) );
  AOI211_X1 U14382 ( .C1(n16275), .C2(P1_REG2_REG_15__SCAN_IN), .A(n12707), 
        .B(n12706), .ZN(n12708) );
  OAI211_X1 U14383 ( .C1(n16332), .C2(n16181), .A(n12709), .B(n12708), .ZN(
        n12710) );
  AOI21_X1 U14384 ( .B1(n16338), .B2(n15366), .A(n12710), .ZN(n12711) );
  INV_X1 U14385 ( .A(n12711), .ZN(P1_U3278) );
  AOI22_X1 U14386 ( .A1(n12713), .A2(n16103), .B1(n12712), .B2(n16102), .ZN(
        n12714) );
  NAND2_X1 U14387 ( .A1(n12715), .A2(n12714), .ZN(n16221) );
  MUX2_X1 U14388 ( .A(P3_REG1_REG_11__SCAN_IN), .B(n16221), .S(n16238), .Z(
        n13171) );
  XNOR2_X1 U14389 ( .A(P3_WR_REG_SCAN_IN), .B(keyinput_0), .ZN(n12719) );
  XNOR2_X1 U14390 ( .A(SI_31_), .B(keyinput_1), .ZN(n12718) );
  XNOR2_X1 U14391 ( .A(SI_30_), .B(keyinput_2), .ZN(n12717) );
  XNOR2_X1 U14392 ( .A(SI_29_), .B(keyinput_3), .ZN(n12716) );
  OAI211_X1 U14393 ( .C1(n12719), .C2(n12718), .A(n12717), .B(n12716), .ZN(
        n12723) );
  XNOR2_X1 U14394 ( .A(SI_26_), .B(keyinput_6), .ZN(n12722) );
  XNOR2_X1 U14395 ( .A(SI_28_), .B(keyinput_4), .ZN(n12721) );
  XNOR2_X1 U14396 ( .A(SI_27_), .B(keyinput_5), .ZN(n12720) );
  NAND4_X1 U14397 ( .A1(n12723), .A2(n12722), .A3(n12721), .A4(n12720), .ZN(
        n12727) );
  XNOR2_X1 U14398 ( .A(n12724), .B(keyinput_7), .ZN(n12726) );
  XNOR2_X1 U14399 ( .A(SI_24_), .B(keyinput_8), .ZN(n12725) );
  NAND3_X1 U14400 ( .A1(n12727), .A2(n12726), .A3(n12725), .ZN(n12731) );
  XNOR2_X1 U14401 ( .A(SI_23_), .B(keyinput_9), .ZN(n12729) );
  XNOR2_X1 U14402 ( .A(SI_22_), .B(keyinput_10), .ZN(n12728) );
  NOR2_X1 U14403 ( .A1(n12729), .A2(n12728), .ZN(n12730) );
  NAND2_X1 U14404 ( .A1(n12731), .A2(n12730), .ZN(n12735) );
  XNOR2_X1 U14405 ( .A(n12956), .B(keyinput_13), .ZN(n12734) );
  XNOR2_X1 U14406 ( .A(SI_20_), .B(keyinput_12), .ZN(n12733) );
  XNOR2_X1 U14407 ( .A(SI_21_), .B(keyinput_11), .ZN(n12732) );
  NAND4_X1 U14408 ( .A1(n12735), .A2(n12734), .A3(n12733), .A4(n12732), .ZN(
        n12743) );
  XNOR2_X1 U14409 ( .A(n12736), .B(keyinput_14), .ZN(n12742) );
  XNOR2_X1 U14410 ( .A(n12737), .B(keyinput_15), .ZN(n12740) );
  XNOR2_X1 U14411 ( .A(SI_15_), .B(keyinput_17), .ZN(n12739) );
  XNOR2_X1 U14412 ( .A(SI_16_), .B(keyinput_16), .ZN(n12738) );
  NAND3_X1 U14413 ( .A1(n12740), .A2(n12739), .A3(n12738), .ZN(n12741) );
  AOI21_X1 U14414 ( .B1(n12743), .B2(n12742), .A(n12741), .ZN(n12754) );
  XNOR2_X1 U14415 ( .A(SI_14_), .B(keyinput_18), .ZN(n12753) );
  OAI22_X1 U14416 ( .A1(n12971), .A2(keyinput_19), .B1(n12745), .B2(
        keyinput_22), .ZN(n12744) );
  AOI221_X1 U14417 ( .B1(n12971), .B2(keyinput_19), .C1(keyinput_22), .C2(
        n12745), .A(n12744), .ZN(n12752) );
  INV_X1 U14418 ( .A(keyinput_23), .ZN(n12746) );
  NAND2_X1 U14419 ( .A1(n12746), .A2(SI_9_), .ZN(n12748) );
  AOI22_X1 U14420 ( .A1(n12974), .A2(keyinput_23), .B1(n12973), .B2(
        keyinput_21), .ZN(n12747) );
  OAI211_X1 U14421 ( .C1(n12973), .C2(keyinput_21), .A(n12748), .B(n12747), 
        .ZN(n12750) );
  XNOR2_X1 U14422 ( .A(SI_12_), .B(keyinput_20), .ZN(n12749) );
  NOR2_X1 U14423 ( .A1(n12750), .A2(n12749), .ZN(n12751) );
  OAI211_X1 U14424 ( .C1(n12754), .C2(n12753), .A(n12752), .B(n12751), .ZN(
        n12760) );
  XNOR2_X1 U14425 ( .A(SI_8_), .B(keyinput_24), .ZN(n12756) );
  XNOR2_X1 U14426 ( .A(SI_6_), .B(keyinput_26), .ZN(n12755) );
  NOR2_X1 U14427 ( .A1(n12756), .A2(n12755), .ZN(n12759) );
  XNOR2_X1 U14428 ( .A(SI_5_), .B(keyinput_27), .ZN(n12758) );
  XNOR2_X1 U14429 ( .A(SI_7_), .B(keyinput_25), .ZN(n12757) );
  NAND4_X1 U14430 ( .A1(n12760), .A2(n12759), .A3(n12758), .A4(n12757), .ZN(
        n12765) );
  XNOR2_X1 U14431 ( .A(n12761), .B(keyinput_30), .ZN(n12764) );
  XNOR2_X1 U14432 ( .A(SI_4_), .B(keyinput_28), .ZN(n12763) );
  XNOR2_X1 U14433 ( .A(SI_3_), .B(keyinput_29), .ZN(n12762) );
  NAND4_X1 U14434 ( .A1(n12765), .A2(n12764), .A3(n12763), .A4(n12762), .ZN(
        n12767) );
  XNOR2_X1 U14435 ( .A(SI_1_), .B(keyinput_31), .ZN(n12766) );
  NAND2_X1 U14436 ( .A1(n12767), .A2(n12766), .ZN(n12769) );
  XNOR2_X1 U14437 ( .A(SI_0_), .B(keyinput_32), .ZN(n12768) );
  NAND2_X1 U14438 ( .A1(n12769), .A2(n12768), .ZN(n12775) );
  XNOR2_X1 U14439 ( .A(P3_RD_REG_SCAN_IN), .B(keyinput_33), .ZN(n12771) );
  XNOR2_X1 U14440 ( .A(P3_REG3_REG_27__SCAN_IN), .B(keyinput_36), .ZN(n12770)
         );
  NOR2_X1 U14441 ( .A1(n12771), .A2(n12770), .ZN(n12774) );
  XNOR2_X1 U14442 ( .A(P3_REG3_REG_7__SCAN_IN), .B(keyinput_35), .ZN(n12773)
         );
  XNOR2_X1 U14443 ( .A(P3_STATE_REG_SCAN_IN), .B(keyinput_34), .ZN(n12772) );
  NAND4_X1 U14444 ( .A1(n12775), .A2(n12774), .A3(n12773), .A4(n12772), .ZN(
        n12786) );
  INV_X1 U14445 ( .A(keyinput_37), .ZN(n12776) );
  XNOR2_X1 U14446 ( .A(n12776), .B(P3_REG3_REG_14__SCAN_IN), .ZN(n12780) );
  XNOR2_X1 U14447 ( .A(P3_REG3_REG_3__SCAN_IN), .B(keyinput_40), .ZN(n12779)
         );
  XNOR2_X1 U14448 ( .A(P3_REG3_REG_10__SCAN_IN), .B(keyinput_39), .ZN(n12778)
         );
  XNOR2_X1 U14449 ( .A(P3_REG3_REG_23__SCAN_IN), .B(keyinput_38), .ZN(n12777)
         );
  NAND4_X1 U14450 ( .A1(n12780), .A2(n12779), .A3(n12778), .A4(n12777), .ZN(
        n12783) );
  XNOR2_X1 U14451 ( .A(P3_REG3_REG_19__SCAN_IN), .B(keyinput_41), .ZN(n12782)
         );
  XNOR2_X1 U14452 ( .A(P3_REG3_REG_28__SCAN_IN), .B(keyinput_42), .ZN(n12781)
         );
  NOR3_X1 U14453 ( .A1(n12783), .A2(n12782), .A3(n12781), .ZN(n12785) );
  XNOR2_X1 U14454 ( .A(P3_REG3_REG_8__SCAN_IN), .B(keyinput_43), .ZN(n12784)
         );
  AOI21_X1 U14455 ( .B1(n12786), .B2(n12785), .A(n12784), .ZN(n12790) );
  XNOR2_X1 U14456 ( .A(P3_REG3_REG_1__SCAN_IN), .B(keyinput_44), .ZN(n12789)
         );
  XNOR2_X1 U14457 ( .A(n12787), .B(keyinput_45), .ZN(n12788) );
  OAI21_X1 U14458 ( .B1(n12790), .B2(n12789), .A(n12788), .ZN(n12792) );
  XNOR2_X1 U14459 ( .A(P3_REG3_REG_12__SCAN_IN), .B(keyinput_46), .ZN(n12791)
         );
  NAND2_X1 U14460 ( .A1(n12792), .A2(n12791), .ZN(n12796) );
  XNOR2_X1 U14461 ( .A(P3_REG3_REG_25__SCAN_IN), .B(keyinput_47), .ZN(n12794)
         );
  XNOR2_X1 U14462 ( .A(P3_REG3_REG_16__SCAN_IN), .B(keyinput_48), .ZN(n12793)
         );
  NOR2_X1 U14463 ( .A1(n12794), .A2(n12793), .ZN(n12795) );
  NAND2_X1 U14464 ( .A1(n12796), .A2(n12795), .ZN(n12801) );
  XNOR2_X1 U14465 ( .A(n13020), .B(keyinput_50), .ZN(n12800) );
  INV_X1 U14466 ( .A(keyinput_49), .ZN(n12797) );
  XNOR2_X1 U14467 ( .A(n12797), .B(P3_REG3_REG_5__SCAN_IN), .ZN(n12799) );
  XNOR2_X1 U14468 ( .A(P3_REG3_REG_24__SCAN_IN), .B(keyinput_51), .ZN(n12798)
         );
  NAND4_X1 U14469 ( .A1(n12801), .A2(n12800), .A3(n12799), .A4(n12798), .ZN(
        n12811) );
  XNOR2_X1 U14470 ( .A(P3_REG3_REG_4__SCAN_IN), .B(keyinput_52), .ZN(n12810)
         );
  XNOR2_X1 U14471 ( .A(n12802), .B(keyinput_55), .ZN(n12808) );
  INV_X1 U14472 ( .A(keyinput_56), .ZN(n12803) );
  XNOR2_X1 U14473 ( .A(n12803), .B(P3_REG3_REG_13__SCAN_IN), .ZN(n12807) );
  INV_X1 U14474 ( .A(keyinput_54), .ZN(n12804) );
  XNOR2_X1 U14475 ( .A(n12804), .B(P3_REG3_REG_0__SCAN_IN), .ZN(n12806) );
  XNOR2_X1 U14476 ( .A(P3_REG3_REG_9__SCAN_IN), .B(keyinput_53), .ZN(n12805)
         );
  NAND4_X1 U14477 ( .A1(n12808), .A2(n12807), .A3(n12806), .A4(n12805), .ZN(
        n12809) );
  AOI21_X1 U14478 ( .B1(n12811), .B2(n12810), .A(n12809), .ZN(n12816) );
  XNOR2_X1 U14479 ( .A(P3_REG3_REG_22__SCAN_IN), .B(keyinput_57), .ZN(n12815)
         );
  INV_X1 U14480 ( .A(keyinput_59), .ZN(n12812) );
  XNOR2_X1 U14481 ( .A(n12812), .B(P3_REG3_REG_2__SCAN_IN), .ZN(n12814) );
  XNOR2_X1 U14482 ( .A(P3_REG3_REG_11__SCAN_IN), .B(keyinput_58), .ZN(n12813)
         );
  OAI211_X1 U14483 ( .C1(n12816), .C2(n12815), .A(n12814), .B(n12813), .ZN(
        n12822) );
  INV_X1 U14484 ( .A(keyinput_62), .ZN(n12817) );
  XNOR2_X1 U14485 ( .A(n12817), .B(P3_REG3_REG_26__SCAN_IN), .ZN(n12821) );
  INV_X1 U14486 ( .A(keyinput_61), .ZN(n12818) );
  XNOR2_X1 U14487 ( .A(n12818), .B(P3_REG3_REG_6__SCAN_IN), .ZN(n12820) );
  XNOR2_X1 U14488 ( .A(P3_REG3_REG_18__SCAN_IN), .B(keyinput_60), .ZN(n12819)
         );
  NAND4_X1 U14489 ( .A1(n12822), .A2(n12821), .A3(n12820), .A4(n12819), .ZN(
        n12826) );
  INV_X1 U14490 ( .A(keyinput_64), .ZN(n12823) );
  XNOR2_X1 U14491 ( .A(n12823), .B(P3_B_REG_SCAN_IN), .ZN(n12825) );
  XNOR2_X1 U14492 ( .A(P3_REG3_REG_15__SCAN_IN), .B(keyinput_63), .ZN(n12824)
         );
  NAND3_X1 U14493 ( .A1(n12826), .A2(n12825), .A3(n12824), .ZN(n12832) );
  XNOR2_X1 U14494 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(keyinput_66), .ZN(n12828)
         );
  XNOR2_X1 U14495 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(keyinput_67), .ZN(n12827)
         );
  NOR2_X1 U14496 ( .A1(n12828), .A2(n12827), .ZN(n12831) );
  XNOR2_X1 U14497 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(keyinput_68), .ZN(n12830)
         );
  XNOR2_X1 U14498 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(keyinput_65), .ZN(n12829)
         );
  NAND4_X1 U14499 ( .A1(n12832), .A2(n12831), .A3(n12830), .A4(n12829), .ZN(
        n12834) );
  XNOR2_X1 U14500 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(keyinput_69), .ZN(n12833)
         );
  NAND2_X1 U14501 ( .A1(n12834), .A2(n12833), .ZN(n12837) );
  XNOR2_X1 U14502 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(keyinput_70), .ZN(n12836)
         );
  XNOR2_X1 U14503 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(keyinput_71), .ZN(n12835)
         );
  NAND3_X1 U14504 ( .A1(n12837), .A2(n12836), .A3(n12835), .ZN(n12840) );
  XNOR2_X1 U14505 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(keyinput_72), .ZN(n12839)
         );
  XNOR2_X1 U14506 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(keyinput_73), .ZN(n12838)
         );
  AOI21_X1 U14507 ( .B1(n12840), .B2(n12839), .A(n12838), .ZN(n12845) );
  INV_X1 U14508 ( .A(keyinput_76), .ZN(n12841) );
  XNOR2_X1 U14509 ( .A(n12841), .B(P3_DATAO_REG_20__SCAN_IN), .ZN(n12844) );
  XNOR2_X1 U14510 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(keyinput_75), .ZN(n12843)
         );
  XNOR2_X1 U14511 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(keyinput_74), .ZN(n12842)
         );
  OR4_X1 U14512 ( .A1(n12845), .A2(n12844), .A3(n12843), .A4(n12842), .ZN(
        n12847) );
  XNOR2_X1 U14513 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(keyinput_77), .ZN(n12846)
         );
  NAND2_X1 U14514 ( .A1(n12847), .A2(n12846), .ZN(n12850) );
  XNOR2_X1 U14515 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(keyinput_78), .ZN(n12849)
         );
  XNOR2_X1 U14516 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(keyinput_79), .ZN(n12848)
         );
  AOI21_X1 U14517 ( .B1(n12850), .B2(n12849), .A(n12848), .ZN(n12854) );
  XNOR2_X1 U14518 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(keyinput_80), .ZN(n12853)
         );
  INV_X1 U14519 ( .A(keyinput_81), .ZN(n12851) );
  XNOR2_X1 U14520 ( .A(n12851), .B(P3_DATAO_REG_15__SCAN_IN), .ZN(n12852) );
  OAI21_X1 U14521 ( .B1(n12854), .B2(n12853), .A(n12852), .ZN(n12870) );
  INV_X1 U14522 ( .A(keyinput_82), .ZN(n12862) );
  INV_X1 U14523 ( .A(P3_DATAO_REG_9__SCAN_IN), .ZN(n12856) );
  NAND2_X1 U14524 ( .A1(n12856), .A2(keyinput_87), .ZN(n12861) );
  INV_X1 U14525 ( .A(P3_DATAO_REG_14__SCAN_IN), .ZN(n12855) );
  OAI22_X1 U14526 ( .A1(n12856), .A2(keyinput_87), .B1(n12855), .B2(
        keyinput_82), .ZN(n12859) );
  OAI22_X1 U14527 ( .A1(P3_DATAO_REG_8__SCAN_IN), .A2(keyinput_88), .B1(
        keyinput_83), .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n12858) );
  INV_X1 U14528 ( .A(P3_DATAO_REG_10__SCAN_IN), .ZN(n13079) );
  OAI22_X1 U14529 ( .A1(n13079), .A2(keyinput_86), .B1(keyinput_85), .B2(
        P3_DATAO_REG_11__SCAN_IN), .ZN(n12857) );
  NOR3_X1 U14530 ( .A1(n12859), .A2(n12858), .A3(n12857), .ZN(n12860) );
  OAI211_X1 U14531 ( .C1(n12862), .C2(P3_DATAO_REG_14__SCAN_IN), .A(n12861), 
        .B(n12860), .ZN(n12863) );
  INV_X1 U14532 ( .A(n12863), .ZN(n12867) );
  AOI22_X1 U14533 ( .A1(P3_DATAO_REG_13__SCAN_IN), .A2(keyinput_83), .B1(
        P3_DATAO_REG_11__SCAN_IN), .B2(keyinput_85), .ZN(n12866) );
  AOI22_X1 U14534 ( .A1(n13079), .A2(keyinput_86), .B1(P3_DATAO_REG_8__SCAN_IN), .B2(keyinput_88), .ZN(n12865) );
  XNOR2_X1 U14535 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(keyinput_84), .ZN(n12864)
         );
  AND4_X1 U14536 ( .A1(n12867), .A2(n12866), .A3(n12865), .A4(n12864), .ZN(
        n12869) );
  XNOR2_X1 U14537 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(keyinput_89), .ZN(n12868)
         );
  AOI21_X1 U14538 ( .B1(n12870), .B2(n12869), .A(n12868), .ZN(n12881) );
  XNOR2_X1 U14539 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(keyinput_90), .ZN(n12872)
         );
  XNOR2_X1 U14540 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(keyinput_91), .ZN(n12871)
         );
  NOR2_X1 U14541 ( .A1(n12872), .A2(n12871), .ZN(n12878) );
  INV_X1 U14542 ( .A(keyinput_94), .ZN(n12873) );
  XNOR2_X1 U14543 ( .A(n12873), .B(P3_DATAO_REG_2__SCAN_IN), .ZN(n12877) );
  INV_X1 U14544 ( .A(keyinput_92), .ZN(n12874) );
  XNOR2_X1 U14545 ( .A(n12874), .B(P3_DATAO_REG_4__SCAN_IN), .ZN(n12876) );
  XNOR2_X1 U14546 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(keyinput_93), .ZN(n12875)
         );
  NAND4_X1 U14547 ( .A1(n12878), .A2(n12877), .A3(n12876), .A4(n12875), .ZN(
        n12880) );
  XNOR2_X1 U14548 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(keyinput_95), .ZN(n12879)
         );
  OAI21_X1 U14549 ( .B1(n12881), .B2(n12880), .A(n12879), .ZN(n12883) );
  XNOR2_X1 U14550 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(keyinput_96), .ZN(n12882)
         );
  NAND2_X1 U14551 ( .A1(n12883), .A2(n12882), .ZN(n12885) );
  XNOR2_X1 U14552 ( .A(P3_ADDR_REG_0__SCAN_IN), .B(keyinput_97), .ZN(n12884)
         );
  NAND2_X1 U14553 ( .A1(n12885), .A2(n12884), .ZN(n12891) );
  XNOR2_X1 U14554 ( .A(P3_ADDR_REG_2__SCAN_IN), .B(keyinput_99), .ZN(n12887)
         );
  XNOR2_X1 U14555 ( .A(P3_ADDR_REG_4__SCAN_IN), .B(keyinput_101), .ZN(n12886)
         );
  NOR2_X1 U14556 ( .A1(n12887), .A2(n12886), .ZN(n12890) );
  XNOR2_X1 U14557 ( .A(P3_ADDR_REG_3__SCAN_IN), .B(keyinput_100), .ZN(n12889)
         );
  XNOR2_X1 U14558 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(keyinput_98), .ZN(n12888)
         );
  NAND4_X1 U14559 ( .A1(n12891), .A2(n12890), .A3(n12889), .A4(n12888), .ZN(
        n12895) );
  INV_X1 U14560 ( .A(keyinput_102), .ZN(n12892) );
  XNOR2_X1 U14561 ( .A(n12892), .B(P3_ADDR_REG_5__SCAN_IN), .ZN(n12894) );
  XNOR2_X1 U14562 ( .A(P3_ADDR_REG_6__SCAN_IN), .B(keyinput_103), .ZN(n12893)
         );
  AOI21_X1 U14563 ( .B1(n12895), .B2(n12894), .A(n12893), .ZN(n12902) );
  INV_X1 U14564 ( .A(keyinput_107), .ZN(n12896) );
  XNOR2_X1 U14565 ( .A(n12896), .B(P1_IR_REG_0__SCAN_IN), .ZN(n12898) );
  XNOR2_X1 U14566 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(keyinput_104), .ZN(n12897)
         );
  NAND2_X1 U14567 ( .A1(n12898), .A2(n12897), .ZN(n12901) );
  XNOR2_X1 U14568 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(keyinput_105), .ZN(n12900)
         );
  XNOR2_X1 U14569 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(keyinput_106), .ZN(n12899)
         );
  OR4_X1 U14570 ( .A1(n12902), .A2(n12901), .A3(n12900), .A4(n12899), .ZN(
        n12905) );
  INV_X1 U14571 ( .A(keyinput_108), .ZN(n12903) );
  XNOR2_X1 U14572 ( .A(n12903), .B(P1_IR_REG_1__SCAN_IN), .ZN(n12904) );
  NAND2_X1 U14573 ( .A1(n12905), .A2(n12904), .ZN(n12907) );
  XNOR2_X1 U14574 ( .A(n13132), .B(keyinput_109), .ZN(n12906) );
  NAND2_X1 U14575 ( .A1(n12907), .A2(n12906), .ZN(n12909) );
  XNOR2_X1 U14576 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_110), .ZN(n12908) );
  NAND2_X1 U14577 ( .A1(n12909), .A2(n12908), .ZN(n12913) );
  INV_X1 U14578 ( .A(keyinput_112), .ZN(n12910) );
  XNOR2_X1 U14579 ( .A(n12910), .B(P1_IR_REG_5__SCAN_IN), .ZN(n12912) );
  XNOR2_X1 U14580 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_111), .ZN(n12911) );
  NAND3_X1 U14581 ( .A1(n12913), .A2(n12912), .A3(n12911), .ZN(n12922) );
  XNOR2_X1 U14582 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_113), .ZN(n12921) );
  XNOR2_X1 U14583 ( .A(n12914), .B(keyinput_116), .ZN(n12919) );
  INV_X1 U14584 ( .A(keyinput_117), .ZN(n12915) );
  XNOR2_X1 U14585 ( .A(n12915), .B(P1_IR_REG_10__SCAN_IN), .ZN(n12918) );
  XNOR2_X1 U14586 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_114), .ZN(n12917) );
  XNOR2_X1 U14587 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_115), .ZN(n12916) );
  NAND4_X1 U14588 ( .A1(n12919), .A2(n12918), .A3(n12917), .A4(n12916), .ZN(
        n12920) );
  AOI21_X1 U14589 ( .B1(n12922), .B2(n12921), .A(n12920), .ZN(n12929) );
  XNOR2_X1 U14590 ( .A(n12923), .B(keyinput_118), .ZN(n12928) );
  XNOR2_X1 U14591 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_120), .ZN(n12925)
         );
  XNOR2_X1 U14592 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_119), .ZN(n12924)
         );
  NAND2_X1 U14593 ( .A1(n12925), .A2(n12924), .ZN(n12927) );
  XNOR2_X1 U14594 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_121), .ZN(n12926)
         );
  XNOR2_X1 U14595 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_122), .ZN(n12932)
         );
  XNOR2_X1 U14596 ( .A(n12930), .B(keyinput_123), .ZN(n12931) );
  AOI21_X1 U14597 ( .B1(n12933), .B2(n12932), .A(n12931), .ZN(n12937) );
  XNOR2_X1 U14598 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_124), .ZN(n12936)
         );
  XNOR2_X1 U14599 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_126), .ZN(n12935)
         );
  XNOR2_X1 U14600 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_125), .ZN(n12934)
         );
  OAI211_X1 U14601 ( .C1(n12937), .C2(n12936), .A(n12935), .B(n12934), .ZN(
        n13169) );
  XNOR2_X1 U14602 ( .A(SI_31_), .B(keyinput_129), .ZN(n12942) );
  XNOR2_X1 U14603 ( .A(P3_WR_REG_SCAN_IN), .B(keyinput_128), .ZN(n12941) );
  INV_X1 U14604 ( .A(keyinput_130), .ZN(n12938) );
  XNOR2_X1 U14605 ( .A(n12938), .B(SI_30_), .ZN(n12940) );
  XNOR2_X1 U14606 ( .A(n13925), .B(keyinput_131), .ZN(n12939) );
  OAI211_X1 U14607 ( .C1(n12942), .C2(n12941), .A(n12940), .B(n12939), .ZN(
        n12947) );
  INV_X1 U14608 ( .A(keyinput_134), .ZN(n12943) );
  XNOR2_X1 U14609 ( .A(n12943), .B(SI_26_), .ZN(n12946) );
  XNOR2_X1 U14610 ( .A(n13249), .B(keyinput_132), .ZN(n12945) );
  XNOR2_X1 U14611 ( .A(SI_27_), .B(keyinput_133), .ZN(n12944) );
  NAND4_X1 U14612 ( .A1(n12947), .A2(n12946), .A3(n12945), .A4(n12944), .ZN(
        n12951) );
  INV_X1 U14613 ( .A(keyinput_136), .ZN(n12948) );
  XNOR2_X1 U14614 ( .A(n12948), .B(SI_24_), .ZN(n12950) );
  XNOR2_X1 U14615 ( .A(SI_25_), .B(keyinput_135), .ZN(n12949) );
  NAND3_X1 U14616 ( .A1(n12951), .A2(n12950), .A3(n12949), .ZN(n12954) );
  XNOR2_X1 U14617 ( .A(SI_23_), .B(keyinput_137), .ZN(n12953) );
  XNOR2_X1 U14618 ( .A(SI_22_), .B(keyinput_138), .ZN(n12952) );
  NAND3_X1 U14619 ( .A1(n12954), .A2(n12953), .A3(n12952), .ZN(n12960) );
  INV_X1 U14620 ( .A(keyinput_139), .ZN(n12955) );
  XNOR2_X1 U14621 ( .A(n12955), .B(SI_21_), .ZN(n12959) );
  XNOR2_X1 U14622 ( .A(n12956), .B(keyinput_141), .ZN(n12958) );
  XNOR2_X1 U14623 ( .A(SI_20_), .B(keyinput_140), .ZN(n12957) );
  NAND4_X1 U14624 ( .A1(n12960), .A2(n12959), .A3(n12958), .A4(n12957), .ZN(
        n12962) );
  XNOR2_X1 U14625 ( .A(SI_18_), .B(keyinput_142), .ZN(n12961) );
  NAND2_X1 U14626 ( .A1(n12962), .A2(n12961), .ZN(n12966) );
  XNOR2_X1 U14627 ( .A(SI_15_), .B(keyinput_145), .ZN(n12965) );
  XNOR2_X1 U14628 ( .A(SI_16_), .B(keyinput_144), .ZN(n12964) );
  XNOR2_X1 U14629 ( .A(SI_17_), .B(keyinput_143), .ZN(n12963) );
  NAND4_X1 U14630 ( .A1(n12966), .A2(n12965), .A3(n12964), .A4(n12963), .ZN(
        n12968) );
  XNOR2_X1 U14631 ( .A(n7846), .B(keyinput_146), .ZN(n12967) );
  NAND2_X1 U14632 ( .A1(n12968), .A2(n12967), .ZN(n12985) );
  AOI22_X1 U14633 ( .A1(n12971), .A2(keyinput_147), .B1(keyinput_148), .B2(
        n12970), .ZN(n12969) );
  OAI221_X1 U14634 ( .B1(n12971), .B2(keyinput_147), .C1(n12970), .C2(
        keyinput_148), .A(n12969), .ZN(n12977) );
  AOI22_X1 U14635 ( .A1(n12974), .A2(keyinput_151), .B1(n12973), .B2(
        keyinput_149), .ZN(n12972) );
  OAI221_X1 U14636 ( .B1(n12974), .B2(keyinput_151), .C1(n12973), .C2(
        keyinput_149), .A(n12972), .ZN(n12976) );
  XNOR2_X1 U14637 ( .A(SI_10_), .B(keyinput_150), .ZN(n12975) );
  NOR3_X1 U14638 ( .A1(n12977), .A2(n12976), .A3(n12975), .ZN(n12984) );
  INV_X1 U14639 ( .A(keyinput_152), .ZN(n12978) );
  XNOR2_X1 U14640 ( .A(n12978), .B(SI_8_), .ZN(n12982) );
  XNOR2_X1 U14641 ( .A(SI_7_), .B(keyinput_153), .ZN(n12981) );
  XNOR2_X1 U14642 ( .A(SI_5_), .B(keyinput_155), .ZN(n12980) );
  XNOR2_X1 U14643 ( .A(SI_6_), .B(keyinput_154), .ZN(n12979) );
  NAND4_X1 U14644 ( .A1(n12982), .A2(n12981), .A3(n12980), .A4(n12979), .ZN(
        n12983) );
  AOI21_X1 U14645 ( .B1(n12985), .B2(n12984), .A(n12983), .ZN(n12992) );
  XNOR2_X1 U14646 ( .A(SI_3_), .B(keyinput_157), .ZN(n12988) );
  XNOR2_X1 U14647 ( .A(SI_4_), .B(keyinput_156), .ZN(n12987) );
  XNOR2_X1 U14648 ( .A(SI_2_), .B(keyinput_158), .ZN(n12986) );
  NAND3_X1 U14649 ( .A1(n12988), .A2(n12987), .A3(n12986), .ZN(n12991) );
  XNOR2_X1 U14650 ( .A(n12989), .B(keyinput_159), .ZN(n12990) );
  OAI21_X1 U14651 ( .B1(n12992), .B2(n12991), .A(n12990), .ZN(n13000) );
  XNOR2_X1 U14652 ( .A(SI_0_), .B(keyinput_160), .ZN(n12999) );
  INV_X1 U14653 ( .A(keyinput_164), .ZN(n12993) );
  XNOR2_X1 U14654 ( .A(n12993), .B(P3_REG3_REG_27__SCAN_IN), .ZN(n12997) );
  XNOR2_X1 U14655 ( .A(P3_STATE_REG_SCAN_IN), .B(keyinput_162), .ZN(n12996) );
  XNOR2_X1 U14656 ( .A(keyinput_161), .B(P3_RD_REG_SCAN_IN), .ZN(n12995) );
  XNOR2_X1 U14657 ( .A(P3_REG3_REG_7__SCAN_IN), .B(keyinput_163), .ZN(n12994)
         );
  NAND4_X1 U14658 ( .A1(n12997), .A2(n12996), .A3(n12995), .A4(n12994), .ZN(
        n12998) );
  AOI21_X1 U14659 ( .B1(n13000), .B2(n12999), .A(n12998), .ZN(n13010) );
  XNOR2_X1 U14660 ( .A(P3_REG3_REG_3__SCAN_IN), .B(keyinput_168), .ZN(n13002)
         );
  XNOR2_X1 U14661 ( .A(P3_REG3_REG_28__SCAN_IN), .B(keyinput_170), .ZN(n13001)
         );
  NOR2_X1 U14662 ( .A1(n13002), .A2(n13001), .ZN(n13008) );
  XNOR2_X1 U14663 ( .A(P3_REG3_REG_10__SCAN_IN), .B(keyinput_167), .ZN(n13004)
         );
  XNOR2_X1 U14664 ( .A(P3_REG3_REG_19__SCAN_IN), .B(keyinput_169), .ZN(n13003)
         );
  NOR2_X1 U14665 ( .A1(n13004), .A2(n13003), .ZN(n13007) );
  XNOR2_X1 U14666 ( .A(P3_REG3_REG_23__SCAN_IN), .B(keyinput_166), .ZN(n13006)
         );
  XNOR2_X1 U14667 ( .A(P3_REG3_REG_14__SCAN_IN), .B(keyinput_165), .ZN(n13005)
         );
  NAND4_X1 U14668 ( .A1(n13008), .A2(n13007), .A3(n13006), .A4(n13005), .ZN(
        n13009) );
  OR2_X1 U14669 ( .A1(n13010), .A2(n13009), .ZN(n13013) );
  XNOR2_X1 U14670 ( .A(P3_REG3_REG_8__SCAN_IN), .B(keyinput_171), .ZN(n13012)
         );
  XNOR2_X1 U14671 ( .A(P3_REG3_REG_1__SCAN_IN), .B(keyinput_172), .ZN(n13011)
         );
  AOI21_X1 U14672 ( .B1(n13013), .B2(n13012), .A(n13011), .ZN(n13016) );
  XNOR2_X1 U14673 ( .A(P3_REG3_REG_21__SCAN_IN), .B(keyinput_173), .ZN(n13015)
         );
  XNOR2_X1 U14674 ( .A(P3_REG3_REG_12__SCAN_IN), .B(keyinput_174), .ZN(n13014)
         );
  OAI21_X1 U14675 ( .B1(n13016), .B2(n13015), .A(n13014), .ZN(n13019) );
  XNOR2_X1 U14676 ( .A(P3_REG3_REG_25__SCAN_IN), .B(keyinput_175), .ZN(n13018)
         );
  XNOR2_X1 U14677 ( .A(P3_REG3_REG_16__SCAN_IN), .B(keyinput_176), .ZN(n13017)
         );
  NAND3_X1 U14678 ( .A1(n13019), .A2(n13018), .A3(n13017), .ZN(n13028) );
  XNOR2_X1 U14679 ( .A(n13020), .B(keyinput_178), .ZN(n13025) );
  INV_X1 U14680 ( .A(keyinput_177), .ZN(n13021) );
  XNOR2_X1 U14681 ( .A(n13021), .B(P3_REG3_REG_5__SCAN_IN), .ZN(n13024) );
  INV_X1 U14682 ( .A(keyinput_179), .ZN(n13022) );
  XNOR2_X1 U14683 ( .A(n13022), .B(P3_REG3_REG_24__SCAN_IN), .ZN(n13023) );
  AND3_X1 U14684 ( .A1(n13025), .A2(n13024), .A3(n13023), .ZN(n13027) );
  XNOR2_X1 U14685 ( .A(P3_REG3_REG_4__SCAN_IN), .B(keyinput_180), .ZN(n13026)
         );
  AOI21_X1 U14686 ( .B1(n13028), .B2(n13027), .A(n13026), .ZN(n13036) );
  INV_X1 U14687 ( .A(keyinput_184), .ZN(n13029) );
  XNOR2_X1 U14688 ( .A(n13029), .B(P3_REG3_REG_13__SCAN_IN), .ZN(n13033) );
  XNOR2_X1 U14689 ( .A(P3_REG3_REG_9__SCAN_IN), .B(keyinput_181), .ZN(n13032)
         );
  XNOR2_X1 U14690 ( .A(P3_REG3_REG_0__SCAN_IN), .B(keyinput_182), .ZN(n13031)
         );
  XNOR2_X1 U14691 ( .A(P3_REG3_REG_20__SCAN_IN), .B(keyinput_183), .ZN(n13030)
         );
  NAND4_X1 U14692 ( .A1(n13033), .A2(n13032), .A3(n13031), .A4(n13030), .ZN(
        n13035) );
  XNOR2_X1 U14693 ( .A(P3_REG3_REG_22__SCAN_IN), .B(keyinput_185), .ZN(n13034)
         );
  OAI21_X1 U14694 ( .B1(n13036), .B2(n13035), .A(n13034), .ZN(n13039) );
  XNOR2_X1 U14695 ( .A(P3_REG3_REG_11__SCAN_IN), .B(keyinput_186), .ZN(n13038)
         );
  XNOR2_X1 U14696 ( .A(P3_REG3_REG_2__SCAN_IN), .B(keyinput_187), .ZN(n13037)
         );
  NAND3_X1 U14697 ( .A1(n13039), .A2(n13038), .A3(n13037), .ZN(n13044) );
  INV_X1 U14698 ( .A(keyinput_189), .ZN(n13040) );
  XNOR2_X1 U14699 ( .A(n13040), .B(P3_REG3_REG_6__SCAN_IN), .ZN(n13043) );
  XNOR2_X1 U14700 ( .A(P3_REG3_REG_18__SCAN_IN), .B(keyinput_188), .ZN(n13042)
         );
  XNOR2_X1 U14701 ( .A(P3_REG3_REG_26__SCAN_IN), .B(keyinput_190), .ZN(n13041)
         );
  NAND4_X1 U14702 ( .A1(n13044), .A2(n13043), .A3(n13042), .A4(n13041), .ZN(
        n13055) );
  INV_X1 U14703 ( .A(keyinput_192), .ZN(n13045) );
  XNOR2_X1 U14704 ( .A(n13045), .B(P3_B_REG_SCAN_IN), .ZN(n13047) );
  XNOR2_X1 U14705 ( .A(P3_REG3_REG_15__SCAN_IN), .B(keyinput_191), .ZN(n13046)
         );
  AND2_X1 U14706 ( .A1(n13047), .A2(n13046), .ZN(n13054) );
  INV_X1 U14707 ( .A(keyinput_196), .ZN(n13048) );
  XNOR2_X1 U14708 ( .A(n13048), .B(P3_DATAO_REG_28__SCAN_IN), .ZN(n13052) );
  XNOR2_X1 U14709 ( .A(keyinput_194), .B(P3_DATAO_REG_30__SCAN_IN), .ZN(n13051) );
  XNOR2_X1 U14710 ( .A(keyinput_193), .B(P3_DATAO_REG_31__SCAN_IN), .ZN(n13050) );
  XNOR2_X1 U14711 ( .A(keyinput_195), .B(P3_DATAO_REG_29__SCAN_IN), .ZN(n13049) );
  NAND4_X1 U14712 ( .A1(n13052), .A2(n13051), .A3(n13050), .A4(n13049), .ZN(
        n13053) );
  AOI21_X1 U14713 ( .B1(n13055), .B2(n13054), .A(n13053), .ZN(n13059) );
  XNOR2_X1 U14714 ( .A(keyinput_197), .B(P3_DATAO_REG_27__SCAN_IN), .ZN(n13058) );
  XNOR2_X1 U14715 ( .A(keyinput_198), .B(P3_DATAO_REG_26__SCAN_IN), .ZN(n13057) );
  XNOR2_X1 U14716 ( .A(keyinput_199), .B(P3_DATAO_REG_25__SCAN_IN), .ZN(n13056) );
  OAI211_X1 U14717 ( .C1(n13059), .C2(n13058), .A(n13057), .B(n13056), .ZN(
        n13063) );
  INV_X1 U14718 ( .A(keyinput_200), .ZN(n13060) );
  XNOR2_X1 U14719 ( .A(n13060), .B(P3_DATAO_REG_24__SCAN_IN), .ZN(n13062) );
  XNOR2_X1 U14720 ( .A(keyinput_201), .B(P3_DATAO_REG_23__SCAN_IN), .ZN(n13061) );
  AOI21_X1 U14721 ( .B1(n13063), .B2(n13062), .A(n13061), .ZN(n13069) );
  XNOR2_X1 U14722 ( .A(keyinput_203), .B(P3_DATAO_REG_21__SCAN_IN), .ZN(n13066) );
  XNOR2_X1 U14723 ( .A(keyinput_202), .B(P3_DATAO_REG_22__SCAN_IN), .ZN(n13065) );
  XNOR2_X1 U14724 ( .A(keyinput_204), .B(P3_DATAO_REG_20__SCAN_IN), .ZN(n13064) );
  NAND3_X1 U14725 ( .A1(n13066), .A2(n13065), .A3(n13064), .ZN(n13068) );
  XNOR2_X1 U14726 ( .A(keyinput_205), .B(P3_DATAO_REG_19__SCAN_IN), .ZN(n13067) );
  OAI21_X1 U14727 ( .B1(n13069), .B2(n13068), .A(n13067), .ZN(n13073) );
  INV_X1 U14728 ( .A(keyinput_206), .ZN(n13070) );
  XNOR2_X1 U14729 ( .A(n13070), .B(P3_DATAO_REG_18__SCAN_IN), .ZN(n13072) );
  XNOR2_X1 U14730 ( .A(keyinput_207), .B(P3_DATAO_REG_17__SCAN_IN), .ZN(n13071) );
  AOI21_X1 U14731 ( .B1(n13073), .B2(n13072), .A(n13071), .ZN(n13077) );
  XNOR2_X1 U14732 ( .A(keyinput_208), .B(P3_DATAO_REG_16__SCAN_IN), .ZN(n13076) );
  INV_X1 U14733 ( .A(keyinput_209), .ZN(n13074) );
  XNOR2_X1 U14734 ( .A(n13074), .B(P3_DATAO_REG_15__SCAN_IN), .ZN(n13075) );
  OAI21_X1 U14735 ( .B1(n13077), .B2(n13076), .A(n13075), .ZN(n13096) );
  INV_X1 U14736 ( .A(P3_DATAO_REG_8__SCAN_IN), .ZN(n13086) );
  INV_X1 U14737 ( .A(keyinput_211), .ZN(n13078) );
  NAND2_X1 U14738 ( .A1(n13078), .A2(P3_DATAO_REG_13__SCAN_IN), .ZN(n13085) );
  AOI22_X1 U14739 ( .A1(n13079), .A2(keyinput_214), .B1(keyinput_216), .B2(
        n13086), .ZN(n13083) );
  INV_X1 U14740 ( .A(P3_DATAO_REG_13__SCAN_IN), .ZN(n13080) );
  AOI22_X1 U14741 ( .A1(keyinput_213), .A2(P3_DATAO_REG_11__SCAN_IN), .B1(
        n13080), .B2(keyinput_211), .ZN(n13082) );
  INV_X1 U14742 ( .A(P3_DATAO_REG_12__SCAN_IN), .ZN(n13090) );
  AOI22_X1 U14743 ( .A1(keyinput_215), .A2(P3_DATAO_REG_9__SCAN_IN), .B1(
        n13090), .B2(keyinput_212), .ZN(n13081) );
  AND3_X1 U14744 ( .A1(n13083), .A2(n13082), .A3(n13081), .ZN(n13084) );
  OAI211_X1 U14745 ( .C1(n13086), .C2(keyinput_216), .A(n13085), .B(n13084), 
        .ZN(n13087) );
  INV_X1 U14746 ( .A(n13087), .ZN(n13095) );
  INV_X1 U14747 ( .A(keyinput_214), .ZN(n13088) );
  NAND2_X1 U14748 ( .A1(n13088), .A2(P3_DATAO_REG_10__SCAN_IN), .ZN(n13089) );
  OAI21_X1 U14749 ( .B1(n13090), .B2(keyinput_212), .A(n13089), .ZN(n13092) );
  OAI22_X1 U14750 ( .A1(keyinput_213), .A2(P3_DATAO_REG_11__SCAN_IN), .B1(
        keyinput_215), .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n13091) );
  NOR2_X1 U14751 ( .A1(n13092), .A2(n13091), .ZN(n13094) );
  XNOR2_X1 U14752 ( .A(keyinput_210), .B(P3_DATAO_REG_14__SCAN_IN), .ZN(n13093) );
  NAND4_X1 U14753 ( .A1(n13096), .A2(n13095), .A3(n13094), .A4(n13093), .ZN(
        n13107) );
  XNOR2_X1 U14754 ( .A(keyinput_217), .B(P3_DATAO_REG_7__SCAN_IN), .ZN(n13106)
         );
  XNOR2_X1 U14755 ( .A(keyinput_221), .B(P3_DATAO_REG_3__SCAN_IN), .ZN(n13098)
         );
  XNOR2_X1 U14756 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(keyinput_219), .ZN(n13097)
         );
  NOR2_X1 U14757 ( .A1(n13098), .A2(n13097), .ZN(n13104) );
  INV_X1 U14758 ( .A(keyinput_220), .ZN(n13099) );
  XNOR2_X1 U14759 ( .A(n13099), .B(P3_DATAO_REG_4__SCAN_IN), .ZN(n13103) );
  INV_X1 U14760 ( .A(keyinput_218), .ZN(n13100) );
  XNOR2_X1 U14761 ( .A(n13100), .B(P3_DATAO_REG_6__SCAN_IN), .ZN(n13102) );
  XNOR2_X1 U14762 ( .A(keyinput_222), .B(P3_DATAO_REG_2__SCAN_IN), .ZN(n13101)
         );
  NAND4_X1 U14763 ( .A1(n13104), .A2(n13103), .A3(n13102), .A4(n13101), .ZN(
        n13105) );
  AOI21_X1 U14764 ( .B1(n13107), .B2(n13106), .A(n13105), .ZN(n13111) );
  INV_X1 U14765 ( .A(keyinput_223), .ZN(n13108) );
  XNOR2_X1 U14766 ( .A(n13108), .B(P3_DATAO_REG_1__SCAN_IN), .ZN(n13110) );
  XNOR2_X1 U14767 ( .A(keyinput_224), .B(P3_DATAO_REG_0__SCAN_IN), .ZN(n13109)
         );
  OAI21_X1 U14768 ( .B1(n13111), .B2(n13110), .A(n13109), .ZN(n13113) );
  XNOR2_X1 U14769 ( .A(P3_ADDR_REG_0__SCAN_IN), .B(keyinput_225), .ZN(n13112)
         );
  NAND2_X1 U14770 ( .A1(n13113), .A2(n13112), .ZN(n13120) );
  INV_X1 U14771 ( .A(keyinput_229), .ZN(n13114) );
  XNOR2_X1 U14772 ( .A(n13114), .B(P3_ADDR_REG_4__SCAN_IN), .ZN(n13118) );
  XNOR2_X1 U14773 ( .A(keyinput_227), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n13117)
         );
  XNOR2_X1 U14774 ( .A(keyinput_226), .B(P3_ADDR_REG_1__SCAN_IN), .ZN(n13116)
         );
  XNOR2_X1 U14775 ( .A(keyinput_228), .B(P3_ADDR_REG_3__SCAN_IN), .ZN(n13115)
         );
  AND4_X1 U14776 ( .A1(n13118), .A2(n13117), .A3(n13116), .A4(n13115), .ZN(
        n13119) );
  NAND2_X1 U14777 ( .A1(n13120), .A2(n13119), .ZN(n13123) );
  XNOR2_X1 U14778 ( .A(keyinput_230), .B(P3_ADDR_REG_5__SCAN_IN), .ZN(n13122)
         );
  XNOR2_X1 U14779 ( .A(P3_ADDR_REG_6__SCAN_IN), .B(keyinput_231), .ZN(n13121)
         );
  AOI21_X1 U14780 ( .B1(n13123), .B2(n13122), .A(n13121), .ZN(n13131) );
  INV_X1 U14781 ( .A(keyinput_235), .ZN(n13124) );
  XNOR2_X1 U14782 ( .A(n13124), .B(P1_IR_REG_0__SCAN_IN), .ZN(n13128) );
  XNOR2_X1 U14783 ( .A(keyinput_234), .B(P3_ADDR_REG_9__SCAN_IN), .ZN(n13127)
         );
  XNOR2_X1 U14784 ( .A(keyinput_233), .B(P3_ADDR_REG_8__SCAN_IN), .ZN(n13126)
         );
  XNOR2_X1 U14785 ( .A(keyinput_232), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n13125)
         );
  NAND4_X1 U14786 ( .A1(n13128), .A2(n13127), .A3(n13126), .A4(n13125), .ZN(
        n13130) );
  XNOR2_X1 U14787 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_236), .ZN(n13129) );
  OAI21_X1 U14788 ( .B1(n13131), .B2(n13130), .A(n13129), .ZN(n13135) );
  XNOR2_X1 U14789 ( .A(n13132), .B(keyinput_237), .ZN(n13134) );
  XNOR2_X1 U14790 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_238), .ZN(n13133) );
  AOI21_X1 U14791 ( .B1(n13135), .B2(n13134), .A(n13133), .ZN(n13138) );
  XNOR2_X1 U14792 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_239), .ZN(n13137) );
  XNOR2_X1 U14793 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_240), .ZN(n13136) );
  OR3_X1 U14794 ( .A1(n13138), .A2(n13137), .A3(n13136), .ZN(n13146) );
  XNOR2_X1 U14795 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_241), .ZN(n13145) );
  XNOR2_X1 U14796 ( .A(n8602), .B(keyinput_242), .ZN(n13143) );
  INV_X1 U14797 ( .A(keyinput_245), .ZN(n13139) );
  XNOR2_X1 U14798 ( .A(n13139), .B(P1_IR_REG_10__SCAN_IN), .ZN(n13142) );
  XNOR2_X1 U14799 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_244), .ZN(n13141) );
  XNOR2_X1 U14800 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_243), .ZN(n13140) );
  NAND4_X1 U14801 ( .A1(n13143), .A2(n13142), .A3(n13141), .A4(n13140), .ZN(
        n13144) );
  AOI21_X1 U14802 ( .B1(n13146), .B2(n13145), .A(n13144), .ZN(n13157) );
  XNOR2_X1 U14803 ( .A(n13147), .B(keyinput_247), .ZN(n13153) );
  XNOR2_X1 U14804 ( .A(n13148), .B(keyinput_248), .ZN(n13152) );
  INV_X1 U14805 ( .A(keyinput_249), .ZN(n13149) );
  XNOR2_X1 U14806 ( .A(n13149), .B(P1_IR_REG_14__SCAN_IN), .ZN(n13151) );
  XNOR2_X1 U14807 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_246), .ZN(n13150)
         );
  NAND4_X1 U14808 ( .A1(n13153), .A2(n13152), .A3(n13151), .A4(n13150), .ZN(
        n13156) );
  XNOR2_X1 U14809 ( .A(n13154), .B(keyinput_250), .ZN(n13155) );
  OAI21_X1 U14810 ( .B1(n13157), .B2(n13156), .A(n13155), .ZN(n13161) );
  XNOR2_X1 U14811 ( .A(n12930), .B(keyinput_251), .ZN(n13160) );
  XNOR2_X1 U14812 ( .A(n13158), .B(keyinput_252), .ZN(n13159) );
  AOI21_X1 U14813 ( .B1(n13161), .B2(n13160), .A(n13159), .ZN(n13166) );
  XNOR2_X1 U14814 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_253), .ZN(n13163)
         );
  XNOR2_X1 U14815 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_254), .ZN(n13162)
         );
  NAND2_X1 U14816 ( .A1(n13163), .A2(n13162), .ZN(n13165) );
  XNOR2_X1 U14817 ( .A(keyinput_127), .B(keyinput_255), .ZN(n13164) );
  OAI21_X1 U14818 ( .B1(n13166), .B2(n13165), .A(n13164), .ZN(n13168) );
  XNOR2_X1 U14819 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_127), .ZN(n13167)
         );
  NAND3_X1 U14820 ( .A1(n13169), .A2(n13168), .A3(n13167), .ZN(n13170) );
  XNOR2_X1 U14821 ( .A(n13171), .B(n13170), .ZN(P3_U3470) );
  CLKBUF_X1 U14822 ( .A(n13172), .Z(n13173) );
  XNOR2_X1 U14823 ( .A(n13173), .B(n13176), .ZN(n13174) );
  OAI222_X1 U14824 ( .A1(n16054), .A2(n13230), .B1(n16056), .B2(n13211), .C1(
        n16053), .C2(n13174), .ZN(n13219) );
  INV_X1 U14825 ( .A(n13219), .ZN(n13185) );
  INV_X1 U14826 ( .A(n13175), .ZN(n13180) );
  AOI21_X1 U14827 ( .B1(n13178), .B2(n13177), .A(n13176), .ZN(n13179) );
  NOR2_X1 U14828 ( .A1(n13180), .A2(n13179), .ZN(n13220) );
  INV_X1 U14829 ( .A(n13181), .ZN(n13232) );
  AOI22_X1 U14830 ( .A1(n14341), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n16094), 
        .B2(n13232), .ZN(n13182) );
  OAI21_X1 U14831 ( .B1(n13235), .B2(n14337), .A(n13182), .ZN(n13183) );
  AOI21_X1 U14832 ( .B1(n13220), .B2(n14339), .A(n13183), .ZN(n13184) );
  OAI21_X1 U14833 ( .B1(n13185), .B2(n14341), .A(n13184), .ZN(P3_U3220) );
  XNOR2_X1 U14834 ( .A(n13186), .B(n9734), .ZN(n13187) );
  AOI222_X1 U14835 ( .A1(n9714), .A2(n13187), .B1(n14049), .B2(n14384), .C1(
        n14047), .C2(n14304), .ZN(n14421) );
  XNOR2_X1 U14836 ( .A(n13189), .B(n13188), .ZN(n14419) );
  INV_X1 U14837 ( .A(n13190), .ZN(n13940) );
  AOI22_X1 U14838 ( .A1(n14341), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n16094), 
        .B2(n13940), .ZN(n13191) );
  OAI21_X1 U14839 ( .B1(n14422), .B2(n14337), .A(n13191), .ZN(n13192) );
  AOI21_X1 U14840 ( .B1(n14419), .B2(n14339), .A(n13192), .ZN(n13193) );
  OAI21_X1 U14841 ( .B1(n14421), .B2(n14341), .A(n13193), .ZN(P3_U3219) );
  OAI21_X1 U14842 ( .B1(n13196), .B2(n13195), .A(n13194), .ZN(n13206) );
  AOI21_X1 U14843 ( .B1(n16039), .B2(n14049), .A(n13197), .ZN(n13204) );
  INV_X1 U14844 ( .A(n13198), .ZN(n13199) );
  NAND2_X1 U14845 ( .A1(n14023), .A2(n13199), .ZN(n13203) );
  OR2_X1 U14846 ( .A1(n14017), .A2(n16232), .ZN(n13202) );
  OR2_X1 U14847 ( .A1(n14015), .A2(n13200), .ZN(n13201) );
  NAND4_X1 U14848 ( .A1(n13204), .A2(n13203), .A3(n13202), .A4(n13201), .ZN(
        n13205) );
  AOI21_X1 U14849 ( .B1(n13206), .B2(n16041), .A(n13205), .ZN(n13207) );
  INV_X1 U14850 ( .A(n13207), .ZN(P3_U3164) );
  XNOR2_X1 U14851 ( .A(n13208), .B(n13209), .ZN(n13210) );
  OAI222_X1 U14852 ( .A1(n16054), .A2(n13211), .B1(n16056), .B2(n14317), .C1(
        n13210), .C2(n16053), .ZN(n14414) );
  INV_X1 U14853 ( .A(n14414), .ZN(n13218) );
  OAI21_X1 U14854 ( .B1(n13214), .B2(n13213), .A(n13212), .ZN(n14415) );
  NOR2_X1 U14855 ( .A1(n14463), .A2(n14337), .ZN(n13216) );
  OAI22_X1 U14856 ( .A1(n16100), .A2(n14078), .B1(n14037), .B2(n16059), .ZN(
        n13215) );
  AOI211_X1 U14857 ( .C1(n14415), .C2(n14339), .A(n13216), .B(n13215), .ZN(
        n13217) );
  OAI21_X1 U14858 ( .B1(n13218), .B2(n14341), .A(n13217), .ZN(P3_U3218) );
  INV_X1 U14859 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n13221) );
  AOI21_X1 U14860 ( .B1(n13220), .B2(n16103), .A(n13219), .ZN(n13223) );
  MUX2_X1 U14861 ( .A(n13221), .B(n13223), .S(n16242), .Z(n13222) );
  OAI21_X1 U14862 ( .B1(n14464), .B2(n13235), .A(n13222), .ZN(P3_U3429) );
  MUX2_X1 U14863 ( .A(n9479), .B(n13223), .S(n16238), .Z(n13224) );
  OAI21_X1 U14864 ( .B1(n14418), .B2(n13235), .A(n13224), .ZN(P3_U3472) );
  AOI21_X1 U14865 ( .B1(n13226), .B2(n13225), .A(n14041), .ZN(n13228) );
  NAND2_X1 U14866 ( .A1(n13228), .A2(n13227), .ZN(n13234) );
  AND2_X1 U14867 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n14070) );
  AOI21_X1 U14868 ( .B1(n16039), .B2(n14048), .A(n14070), .ZN(n13229) );
  OAI21_X1 U14869 ( .B1(n13230), .B2(n14015), .A(n13229), .ZN(n13231) );
  AOI21_X1 U14870 ( .B1(n13232), .B2(n14023), .A(n13231), .ZN(n13233) );
  OAI211_X1 U14871 ( .C1(n14017), .C2(n13235), .A(n13234), .B(n13233), .ZN(
        P3_U3174) );
  INV_X1 U14872 ( .A(n13387), .ZN(n13238) );
  AOI21_X1 U14873 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n15601), .A(n13236), 
        .ZN(n13237) );
  OAI21_X1 U14874 ( .B1(n13238), .B2(n15604), .A(n13237), .ZN(P1_U3332) );
  INV_X1 U14875 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n13239) );
  INV_X1 U14876 ( .A(n13462), .ZN(n13241) );
  OAI222_X1 U14877 ( .A1(n15597), .A2(n13239), .B1(n15604), .B2(n13241), .C1(
        P1_U3086), .C2(n10504), .ZN(P1_U3331) );
  INV_X1 U14878 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n13463) );
  OAI222_X1 U14879 ( .A1(n13255), .A2(n13463), .B1(n15061), .B2(n13241), .C1(
        n13240), .C2(P2_U3088), .ZN(P2_U3303) );
  NAND2_X1 U14880 ( .A1(n13387), .A2(n13242), .ZN(n13244) );
  INV_X1 U14881 ( .A(n13243), .ZN(n13900) );
  AND2_X1 U14882 ( .A1(n13900), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13903) );
  INV_X1 U14883 ( .A(n13903), .ZN(n13896) );
  OAI211_X1 U14884 ( .C1(n13388), .C2(n13255), .A(n13244), .B(n13896), .ZN(
        P2_U3304) );
  INV_X1 U14885 ( .A(n13372), .ZN(n15062) );
  OAI222_X1 U14886 ( .A1(n15597), .A2(n13246), .B1(n15604), .B2(n15062), .C1(
        P1_U3086), .C2(n13245), .ZN(P1_U3327) );
  INV_X1 U14887 ( .A(n13247), .ZN(n13250) );
  OAI222_X1 U14888 ( .A1(n13924), .A2(n13250), .B1(n13926), .B2(n13249), .C1(
        P3_U3151), .C2(n13248), .ZN(P3_U3267) );
  OAI222_X1 U14889 ( .A1(n15597), .A2(n13252), .B1(n15604), .B2(n13251), .C1(
        P1_U3086), .C2(n15244), .ZN(P1_U3336) );
  INV_X1 U14890 ( .A(n13446), .ZN(n13254) );
  OAI222_X1 U14891 ( .A1(n13255), .A2(n13447), .B1(n15061), .B2(n13254), .C1(
        n13902), .C2(P2_U3088), .ZN(P2_U3305) );
  NAND2_X1 U14892 ( .A1(n15542), .A2(n13578), .ZN(n13257) );
  NAND2_X1 U14893 ( .A1(n15182), .A2(n13265), .ZN(n13256) );
  NAND2_X1 U14894 ( .A1(n13257), .A2(n13256), .ZN(n13259) );
  XNOR2_X1 U14895 ( .A(n13259), .B(n13268), .ZN(n13293) );
  INV_X1 U14896 ( .A(n15542), .ZN(n15428) );
  INV_X1 U14897 ( .A(n15182), .ZN(n15407) );
  OAI22_X1 U14898 ( .A1(n15428), .A2(n13588), .B1(n15407), .B2(n13587), .ZN(
        n13292) );
  INV_X1 U14899 ( .A(n13260), .ZN(n13263) );
  INV_X1 U14900 ( .A(n13261), .ZN(n13262) );
  AOI22_X1 U14901 ( .A1(n15089), .A2(n13265), .B1(n13572), .B2(n16321), .ZN(
        n13271) );
  NAND2_X1 U14902 ( .A1(n15089), .A2(n13578), .ZN(n13267) );
  NAND2_X1 U14903 ( .A1(n16321), .A2(n13265), .ZN(n13266) );
  NAND2_X1 U14904 ( .A1(n13267), .A2(n13266), .ZN(n13269) );
  XNOR2_X1 U14905 ( .A(n13269), .B(n13268), .ZN(n13273) );
  XOR2_X1 U14906 ( .A(n13271), .B(n13273), .Z(n15085) );
  INV_X1 U14907 ( .A(n13271), .ZN(n13272) );
  NAND2_X1 U14908 ( .A1(n13354), .A2(n13578), .ZN(n13276) );
  NAND2_X1 U14909 ( .A1(n16348), .A2(n13265), .ZN(n13275) );
  NAND2_X1 U14910 ( .A1(n13276), .A2(n13275), .ZN(n13277) );
  XNOR2_X1 U14911 ( .A(n13277), .B(n13268), .ZN(n13279) );
  AOI22_X1 U14912 ( .A1(n13354), .A2(n13265), .B1(n13572), .B2(n16348), .ZN(
        n16320) );
  OAI22_X1 U14913 ( .A1(n16354), .A2(n13588), .B1(n13357), .B2(n13587), .ZN(
        n13283) );
  NAND2_X1 U14914 ( .A1(n15454), .A2(n13578), .ZN(n13281) );
  NAND2_X1 U14915 ( .A1(n16322), .A2(n13265), .ZN(n13280) );
  NAND2_X1 U14916 ( .A1(n13281), .A2(n13280), .ZN(n13282) );
  XNOR2_X1 U14917 ( .A(n13282), .B(n13268), .ZN(n13284) );
  XOR2_X1 U14918 ( .A(n13283), .B(n13284), .Z(n16346) );
  NAND2_X1 U14919 ( .A1(n16347), .A2(n16346), .ZN(n13286) );
  OR2_X1 U14920 ( .A1(n13284), .A2(n13283), .ZN(n13285) );
  INV_X1 U14921 ( .A(n15550), .ZN(n13332) );
  OAI22_X1 U14922 ( .A1(n13332), .A2(n13588), .B1(n15158), .B2(n13587), .ZN(
        n13290) );
  NAND2_X1 U14923 ( .A1(n15550), .A2(n13578), .ZN(n13288) );
  NAND2_X1 U14924 ( .A1(n16350), .A2(n13265), .ZN(n13287) );
  NAND2_X1 U14925 ( .A1(n13288), .A2(n13287), .ZN(n13289) );
  XNOR2_X1 U14926 ( .A(n13289), .B(n13268), .ZN(n13291) );
  XOR2_X1 U14927 ( .A(n13290), .B(n13291), .Z(n15130) );
  XOR2_X1 U14928 ( .A(n13292), .B(n13293), .Z(n15157) );
  INV_X1 U14929 ( .A(n15534), .ZN(n15412) );
  INV_X1 U14930 ( .A(n15421), .ZN(n13361) );
  OAI22_X1 U14931 ( .A1(n15412), .A2(n13588), .B1(n13361), .B2(n13587), .ZN(
        n13297) );
  NAND2_X1 U14932 ( .A1(n15534), .A2(n13578), .ZN(n13295) );
  NAND2_X1 U14933 ( .A1(n15421), .A2(n13265), .ZN(n13294) );
  NAND2_X1 U14934 ( .A1(n13295), .A2(n13294), .ZN(n13296) );
  XNOR2_X1 U14935 ( .A(n13296), .B(n13268), .ZN(n13298) );
  XOR2_X1 U14936 ( .A(n13297), .B(n13298), .Z(n15106) );
  NAND2_X1 U14937 ( .A1(n13300), .A2(n13299), .ZN(n15146) );
  INV_X1 U14938 ( .A(n15146), .ZN(n13306) );
  AND2_X1 U14939 ( .A1(n15375), .A2(n13572), .ZN(n13301) );
  AOI21_X1 U14940 ( .B1(n15528), .B2(n13265), .A(n13301), .ZN(n13307) );
  NAND2_X1 U14941 ( .A1(n15528), .A2(n13578), .ZN(n13303) );
  NAND2_X1 U14942 ( .A1(n15375), .A2(n13265), .ZN(n13302) );
  NAND2_X1 U14943 ( .A1(n13303), .A2(n13302), .ZN(n13304) );
  XNOR2_X1 U14944 ( .A(n13304), .B(n13268), .ZN(n13309) );
  XOR2_X1 U14945 ( .A(n13307), .B(n13309), .Z(n15145) );
  INV_X1 U14946 ( .A(n15145), .ZN(n13305) );
  INV_X1 U14947 ( .A(n13307), .ZN(n13308) );
  NAND2_X1 U14948 ( .A1(n13309), .A2(n13308), .ZN(n13310) );
  AOI22_X1 U14949 ( .A1(n15525), .A2(n13578), .B1(n13265), .B2(n15181), .ZN(
        n13311) );
  XNOR2_X1 U14950 ( .A(n13311), .B(n13268), .ZN(n13314) );
  AOI22_X1 U14951 ( .A1(n15525), .A2(n13265), .B1(n13572), .B2(n15181), .ZN(
        n13313) );
  XNOR2_X1 U14952 ( .A(n13314), .B(n13313), .ZN(n15115) );
  INV_X1 U14953 ( .A(n15115), .ZN(n13312) );
  NAND2_X1 U14954 ( .A1(n13314), .A2(n13313), .ZN(n13315) );
  OAI22_X1 U14955 ( .A1(n7417), .A2(n13594), .B1(n15097), .B2(n13588), .ZN(
        n13316) );
  XNOR2_X1 U14956 ( .A(n13316), .B(n13268), .ZN(n13553) );
  OAI22_X1 U14957 ( .A1(n7417), .A2(n13588), .B1(n15097), .B2(n13587), .ZN(
        n13552) );
  XNOR2_X1 U14958 ( .A(n13553), .B(n13552), .ZN(n13318) );
  AOI21_X1 U14959 ( .B1(n13317), .B2(n13318), .A(n15175), .ZN(n13320) );
  INV_X1 U14960 ( .A(n13318), .ZN(n13319) );
  NAND2_X1 U14961 ( .A1(n13320), .A2(n13555), .ZN(n13325) );
  INV_X1 U14962 ( .A(n15180), .ZN(n15324) );
  OAI22_X1 U14963 ( .A1(n13364), .A2(n15406), .B1(n15324), .B2(n15408), .ZN(
        n15354) );
  INV_X1 U14964 ( .A(n15361), .ZN(n13322) );
  OAI22_X1 U14965 ( .A1(n16361), .A2(n13322), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13321), .ZN(n13323) );
  AOI21_X1 U14966 ( .B1(n15354), .B2(n15153), .A(n13323), .ZN(n13324) );
  OAI211_X1 U14967 ( .C1(n16353), .C2(n7417), .A(n13325), .B(n13324), .ZN(
        P1_U3235) );
  INV_X1 U14968 ( .A(n13326), .ZN(n13327) );
  OAI222_X1 U14969 ( .A1(n9278), .A2(P3_U3151), .B1(n13926), .B2(n13328), .C1(
        n13924), .C2(n13327), .ZN(P3_U3265) );
  INV_X1 U14970 ( .A(n13616), .ZN(n13605) );
  OAI222_X1 U14971 ( .A1(n15061), .A2(n13605), .B1(P2_U3088), .B2(n13329), 
        .C1(n13617), .C2(n13255), .ZN(P2_U3297) );
  INV_X1 U14972 ( .A(n7417), .ZN(n15362) );
  INV_X1 U14973 ( .A(n15375), .ZN(n15409) );
  INV_X1 U14974 ( .A(n15528), .ZN(n15393) );
  OAI21_X1 U14975 ( .B1(n13354), .B2(n16348), .A(n13331), .ZN(n15450) );
  NAND2_X1 U14976 ( .A1(n15428), .A2(n15407), .ZN(n13334) );
  INV_X1 U14977 ( .A(n15402), .ZN(n13335) );
  INV_X1 U14978 ( .A(n15369), .ZN(n15373) );
  INV_X1 U14979 ( .A(n13337), .ZN(n15358) );
  NAND2_X1 U14980 ( .A1(n15359), .A2(n15358), .ZN(n15357) );
  OAI21_X1 U14981 ( .B1(n15362), .B2(n15374), .A(n15357), .ZN(n15341) );
  INV_X1 U14982 ( .A(n15321), .ZN(n15308) );
  INV_X1 U14983 ( .A(n15293), .ZN(n15302) );
  INV_X1 U14984 ( .A(n15265), .ZN(n13341) );
  OAI21_X1 U14985 ( .B1(n15079), .B2(n15480), .A(n15268), .ZN(n13343) );
  INV_X1 U14986 ( .A(n13368), .ZN(n13342) );
  OR2_X1 U14987 ( .A1(n15534), .A2(n15404), .ZN(n15405) );
  OR2_X1 U14988 ( .A1(n15405), .A2(n15528), .ZN(n15388) );
  NAND2_X1 U14989 ( .A1(n7417), .A2(n15378), .ZN(n15360) );
  OR2_X1 U14990 ( .A1(n15349), .A2(n15360), .ZN(n15343) );
  INV_X1 U14991 ( .A(n15498), .ZN(n15318) );
  INV_X1 U14992 ( .A(n15491), .ZN(n15301) );
  NAND2_X1 U14993 ( .A1(n13344), .A2(n15269), .ZN(n13345) );
  NOR2_X1 U14994 ( .A1(n15594), .A2(n13346), .ZN(n13347) );
  NOR2_X1 U14995 ( .A1(n15408), .A2(n13347), .ZN(n15250) );
  NAND2_X1 U14996 ( .A1(n15178), .A2(n15250), .ZN(n15473) );
  OAI22_X1 U14997 ( .A1(n13349), .A2(n15473), .B1(n13348), .B2(n16110), .ZN(
        n13350) );
  AOI21_X1 U14998 ( .B1(P1_REG2_REG_29__SCAN_IN), .B2(n16275), .A(n13350), 
        .ZN(n13351) );
  OAI21_X1 U14999 ( .B1(n15474), .B2(n16114), .A(n13351), .ZN(n13352) );
  AOI21_X1 U15000 ( .B1(n15476), .B2(n16073), .A(n13352), .ZN(n13371) );
  OR2_X1 U15001 ( .A1(n13354), .A2(n13353), .ZN(n13355) );
  INV_X1 U15002 ( .A(n15443), .ZN(n13359) );
  AND2_X1 U15003 ( .A1(n15550), .A2(n15158), .ZN(n13358) );
  NAND2_X1 U15004 ( .A1(n15424), .A2(n15423), .ZN(n15422) );
  OR2_X1 U15005 ( .A1(n15542), .A2(n15407), .ZN(n13360) );
  NAND2_X1 U15006 ( .A1(n15534), .A2(n13361), .ZN(n13362) );
  OR2_X1 U15007 ( .A1(n15528), .A2(n15409), .ZN(n13363) );
  OR2_X1 U15008 ( .A1(n15525), .A2(n13364), .ZN(n13365) );
  INV_X1 U15009 ( .A(n15342), .ZN(n13366) );
  INV_X1 U15010 ( .A(n15349), .ZN(n15511) );
  INV_X1 U15011 ( .A(n15312), .ZN(n15125) );
  NOR2_X1 U15012 ( .A1(n15480), .A2(n15282), .ZN(n13367) );
  NAND2_X1 U15013 ( .A1(n15477), .A2(n16179), .ZN(n13370) );
  OAI211_X1 U15014 ( .C1(n15478), .C2(n15466), .A(n13371), .B(n13370), .ZN(
        P1_U3356) );
  NAND2_X1 U15015 ( .A1(n13372), .A2(n13615), .ZN(n13375) );
  OR2_X1 U15016 ( .A1(n13618), .A2(n13373), .ZN(n13374) );
  NAND2_X1 U15017 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(P2_REG3_REG_19__SCAN_IN), 
        .ZN(n13376) );
  INV_X1 U15018 ( .A(n13436), .ZN(n13377) );
  NAND2_X1 U15019 ( .A1(n13377), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n13450) );
  INV_X1 U15020 ( .A(n13466), .ZN(n13378) );
  NAND2_X1 U15021 ( .A1(n13378), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n13479) );
  INV_X1 U15022 ( .A(n13479), .ZN(n13379) );
  NAND2_X1 U15023 ( .A1(n13379), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n13490) );
  INV_X1 U15024 ( .A(n13501), .ZN(n13380) );
  NAND2_X1 U15025 ( .A1(n13380), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n13503) );
  INV_X1 U15026 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n13381) );
  NAND2_X1 U15027 ( .A1(n13503), .A2(n13381), .ZN(n13382) );
  INV_X1 U15028 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n13385) );
  NAND2_X1 U15029 ( .A1(n13523), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n13384) );
  NAND2_X1 U15030 ( .A1(n13517), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n13383) );
  OAI211_X1 U15031 ( .C1(n13385), .C2(n13612), .A(n13384), .B(n13383), .ZN(
        n13386) );
  AOI21_X1 U15032 ( .B1(n14743), .B2(n13522), .A(n13386), .ZN(n14752) );
  NAND2_X1 U15033 ( .A1(n13387), .A2(n13615), .ZN(n13390) );
  OR2_X1 U15034 ( .A1(n13618), .A2(n13388), .ZN(n13389) );
  NAND2_X2 U15035 ( .A1(n13390), .A2(n13389), .ZN(n14975) );
  NAND2_X1 U15036 ( .A1(n13452), .A2(n14534), .ZN(n13391) );
  AND2_X1 U15037 ( .A1(n13466), .A2(n13391), .ZN(n14826) );
  NAND2_X1 U15038 ( .A1(n14826), .A2(n13522), .ZN(n13397) );
  INV_X1 U15039 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n13394) );
  NAND2_X1 U15040 ( .A1(n13523), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n13393) );
  NAND2_X1 U15041 ( .A1(n13517), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n13392) );
  OAI211_X1 U15042 ( .C1(n13394), .C2(n13612), .A(n13393), .B(n13392), .ZN(
        n13395) );
  INV_X1 U15043 ( .A(n13395), .ZN(n13396) );
  NAND2_X1 U15044 ( .A1(n13398), .A2(n13615), .ZN(n13400) );
  AOI22_X1 U15045 ( .A1(n13406), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n13405), 
        .B2(n15695), .ZN(n13399) );
  XNOR2_X1 U15046 ( .A(n15005), .B(n14673), .ZN(n14919) );
  INV_X1 U15047 ( .A(n14674), .ZN(n14915) );
  NAND2_X1 U15048 ( .A1(n15011), .A2(n14915), .ZN(n13402) );
  NOR2_X1 U15049 ( .A1(n15011), .A2(n14915), .ZN(n13401) );
  NAND2_X1 U15050 ( .A1(n13404), .A2(n13615), .ZN(n13408) );
  AOI22_X1 U15051 ( .A1(n13406), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n13405), 
        .B2(n7415), .ZN(n13407) );
  XNOR2_X1 U15052 ( .A(n13423), .B(P2_REG3_REG_19__SCAN_IN), .ZN(n14904) );
  NAND2_X1 U15053 ( .A1(n14904), .A2(n13522), .ZN(n13414) );
  INV_X1 U15054 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13411) );
  NAND2_X1 U15055 ( .A1(n13523), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n13410) );
  NAND2_X1 U15056 ( .A1(n13517), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n13409) );
  OAI211_X1 U15057 ( .C1(n13612), .C2(n13411), .A(n13410), .B(n13409), .ZN(
        n13412) );
  INV_X1 U15058 ( .A(n13412), .ZN(n13413) );
  NAND2_X1 U15059 ( .A1(n13414), .A2(n13413), .ZN(n14884) );
  INV_X1 U15060 ( .A(n14884), .ZN(n14917) );
  OR2_X1 U15061 ( .A1(n15001), .A2(n14917), .ZN(n13416) );
  NAND2_X1 U15062 ( .A1(n15001), .A2(n14917), .ZN(n13415) );
  NAND2_X1 U15063 ( .A1(n13416), .A2(n13415), .ZN(n14896) );
  INV_X1 U15064 ( .A(n14673), .ZN(n14894) );
  AND2_X1 U15065 ( .A1(n15005), .A2(n14894), .ZN(n14897) );
  NAND2_X1 U15066 ( .A1(n13417), .A2(n13615), .ZN(n13420) );
  OR2_X1 U15067 ( .A1(n13618), .A2(n13418), .ZN(n13419) );
  INV_X1 U15068 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n13422) );
  INV_X1 U15069 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13421) );
  OAI21_X1 U15070 ( .B1(n13423), .B2(n13422), .A(n13421), .ZN(n13424) );
  AND2_X1 U15071 ( .A1(n13424), .A2(n13436), .ZN(n14877) );
  NAND2_X1 U15072 ( .A1(n14877), .A2(n13522), .ZN(n13430) );
  INV_X1 U15073 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n13427) );
  NAND2_X1 U15074 ( .A1(n13523), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n13426) );
  NAND2_X1 U15075 ( .A1(n13517), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n13425) );
  OAI211_X1 U15076 ( .C1(n13427), .C2(n13612), .A(n13426), .B(n13425), .ZN(
        n13428) );
  INV_X1 U15077 ( .A(n13428), .ZN(n13429) );
  XNOR2_X1 U15078 ( .A(n14993), .B(n14857), .ZN(n14881) );
  NAND2_X1 U15079 ( .A1(n14882), .A2(n14881), .ZN(n14880) );
  INV_X1 U15080 ( .A(n14857), .ZN(n14895) );
  NAND2_X1 U15081 ( .A1(n14993), .A2(n14895), .ZN(n13431) );
  NAND2_X1 U15082 ( .A1(n14880), .A2(n13431), .ZN(n14855) );
  NAND2_X1 U15083 ( .A1(n13432), .A2(n13615), .ZN(n13435) );
  OR2_X1 U15084 ( .A1(n13618), .A2(n13433), .ZN(n13434) );
  INV_X1 U15085 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n14570) );
  NAND2_X1 U15086 ( .A1(n13436), .A2(n14570), .ZN(n13437) );
  NAND2_X1 U15087 ( .A1(n13450), .A2(n13437), .ZN(n14865) );
  OR2_X1 U15088 ( .A1(n14865), .A2(n13504), .ZN(n13443) );
  INV_X1 U15089 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n13440) );
  NAND2_X1 U15090 ( .A1(n13523), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n13439) );
  NAND2_X1 U15091 ( .A1(n13517), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n13438) );
  OAI211_X1 U15092 ( .C1(n13612), .C2(n13440), .A(n13439), .B(n13438), .ZN(
        n13441) );
  INV_X1 U15093 ( .A(n13441), .ZN(n13442) );
  OR2_X1 U15094 ( .A1(n14987), .A2(n8168), .ZN(n13445) );
  AND2_X1 U15095 ( .A1(n14987), .A2(n8168), .ZN(n13444) );
  NAND2_X1 U15096 ( .A1(n13446), .A2(n13615), .ZN(n13449) );
  OR2_X1 U15097 ( .A1(n13618), .A2(n13447), .ZN(n13448) );
  NAND2_X1 U15098 ( .A1(n13450), .A2(n14619), .ZN(n13451) );
  NAND2_X1 U15099 ( .A1(n13452), .A2(n13451), .ZN(n14841) );
  OR2_X1 U15100 ( .A1(n14841), .A2(n13504), .ZN(n13458) );
  INV_X1 U15101 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n13455) );
  NAND2_X1 U15102 ( .A1(n13517), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n13454) );
  NAND2_X1 U15103 ( .A1(n13523), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n13453) );
  OAI211_X1 U15104 ( .C1(n13455), .C2(n13612), .A(n13454), .B(n13453), .ZN(
        n13456) );
  INV_X1 U15105 ( .A(n13456), .ZN(n13457) );
  INV_X1 U15106 ( .A(n14858), .ZN(n14571) );
  NAND2_X1 U15107 ( .A1(n14981), .A2(n14571), .ZN(n13459) );
  NAND2_X1 U15108 ( .A1(n14834), .A2(n13459), .ZN(n13461) );
  OR2_X1 U15109 ( .A1(n14981), .A2(n14571), .ZN(n13460) );
  INV_X1 U15110 ( .A(n14837), .ZN(n14620) );
  NAND2_X1 U15111 ( .A1(n13462), .A2(n12412), .ZN(n13465) );
  OR2_X1 U15112 ( .A1(n13618), .A2(n13463), .ZN(n13464) );
  NAND2_X2 U15113 ( .A1(n13465), .A2(n13464), .ZN(n14969) );
  INV_X1 U15114 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n14605) );
  NAND2_X1 U15115 ( .A1(n13466), .A2(n14605), .ZN(n13467) );
  NAND2_X1 U15116 ( .A1(n13479), .A2(n13467), .ZN(n14803) );
  OR2_X1 U15117 ( .A1(n14803), .A2(n13504), .ZN(n13473) );
  INV_X1 U15118 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n13470) );
  NAND2_X1 U15119 ( .A1(n13517), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n13469) );
  NAND2_X1 U15120 ( .A1(n13523), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n13468) );
  OAI211_X1 U15121 ( .C1(n13470), .C2(n13612), .A(n13469), .B(n13468), .ZN(
        n13471) );
  INV_X1 U15122 ( .A(n13471), .ZN(n13472) );
  INV_X1 U15123 ( .A(n14819), .ZN(n14535) );
  NAND2_X1 U15124 ( .A1(n14969), .A2(n14535), .ZN(n13475) );
  OR2_X1 U15125 ( .A1(n14969), .A2(n14535), .ZN(n13474) );
  NAND2_X1 U15126 ( .A1(n13475), .A2(n13474), .ZN(n14807) );
  NAND2_X1 U15127 ( .A1(n15070), .A2(n13615), .ZN(n13477) );
  OR2_X1 U15128 ( .A1(n13618), .A2(n15073), .ZN(n13476) );
  INV_X1 U15129 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13478) );
  NAND2_X1 U15130 ( .A1(n13479), .A2(n13478), .ZN(n13480) );
  NAND2_X1 U15131 ( .A1(n13490), .A2(n13480), .ZN(n14788) );
  INV_X1 U15132 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n13483) );
  NAND2_X1 U15133 ( .A1(n13517), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n13482) );
  NAND2_X1 U15134 ( .A1(n13523), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n13481) );
  OAI211_X1 U15135 ( .C1(n13483), .C2(n13612), .A(n13482), .B(n13481), .ZN(
        n13484) );
  INV_X1 U15136 ( .A(n13484), .ZN(n13485) );
  NAND2_X1 U15137 ( .A1(n14964), .A2(n14662), .ZN(n14770) );
  OR2_X1 U15138 ( .A1(n14964), .A2(n14662), .ZN(n13487) );
  NAND2_X1 U15139 ( .A1(n15067), .A2(n13615), .ZN(n13489) );
  OR2_X1 U15140 ( .A1(n13618), .A2(n15068), .ZN(n13488) );
  NAND2_X1 U15141 ( .A1(n13490), .A2(n14660), .ZN(n13491) );
  NAND2_X1 U15142 ( .A1(n14777), .A2(n13522), .ZN(n13497) );
  INV_X1 U15143 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n13494) );
  NAND2_X1 U15144 ( .A1(n13523), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n13493) );
  NAND2_X1 U15145 ( .A1(n13517), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n13492) );
  OAI211_X1 U15146 ( .C1(n13494), .C2(n13612), .A(n13493), .B(n13492), .ZN(
        n13495) );
  INV_X1 U15147 ( .A(n13495), .ZN(n13496) );
  NAND2_X1 U15148 ( .A1(n13497), .A2(n13496), .ZN(n14795) );
  INV_X1 U15149 ( .A(n14795), .ZN(n14751) );
  XNOR2_X1 U15150 ( .A(n14959), .B(n14751), .ZN(n14771) );
  INV_X1 U15151 ( .A(n14771), .ZN(n14768) );
  NAND2_X1 U15152 ( .A1(n14959), .A2(n14751), .ZN(n14754) );
  NAND2_X1 U15153 ( .A1(n15063), .A2(n13615), .ZN(n13500) );
  OR2_X1 U15154 ( .A1(n13618), .A2(n15065), .ZN(n13499) );
  NAND2_X2 U15155 ( .A1(n13500), .A2(n13499), .ZN(n14954) );
  INV_X1 U15156 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n14526) );
  NAND2_X1 U15157 ( .A1(n13501), .A2(n14526), .ZN(n13502) );
  NAND2_X1 U15158 ( .A1(n13503), .A2(n13502), .ZN(n14760) );
  INV_X1 U15159 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n13507) );
  NAND2_X1 U15160 ( .A1(n13517), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n13506) );
  NAND2_X1 U15161 ( .A1(n13523), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n13505) );
  OAI211_X1 U15162 ( .C1(n13507), .C2(n13612), .A(n13506), .B(n13505), .ZN(
        n13508) );
  INV_X1 U15163 ( .A(n13508), .ZN(n13509) );
  INV_X1 U15164 ( .A(n14774), .ZN(n14664) );
  NAND2_X1 U15165 ( .A1(n14954), .A2(n14664), .ZN(n13511) );
  NAND2_X1 U15166 ( .A1(n14949), .A2(n14672), .ZN(n13549) );
  NAND2_X1 U15167 ( .A1(n13549), .A2(n13512), .ZN(n13651) );
  NAND2_X1 U15168 ( .A1(n13513), .A2(n13615), .ZN(n13515) );
  OR2_X1 U15169 ( .A1(n13618), .A2(n15057), .ZN(n13514) );
  INV_X1 U15170 ( .A(n13516), .ZN(n13531) );
  INV_X1 U15171 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n13520) );
  NAND2_X1 U15172 ( .A1(n13517), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n13519) );
  NAND2_X1 U15173 ( .A1(n13523), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n13518) );
  OAI211_X1 U15174 ( .C1(n13520), .C2(n13612), .A(n13519), .B(n13518), .ZN(
        n13521) );
  AOI21_X1 U15175 ( .B1(n13531), .B2(n13522), .A(n13521), .ZN(n13869) );
  XNOR2_X1 U15176 ( .A(n14944), .B(n14740), .ZN(n13653) );
  AOI21_X1 U15177 ( .B1(n13906), .B2(P2_B_REG_SCAN_IN), .A(n14916), .ZN(n14723) );
  NAND2_X1 U15178 ( .A1(n7425), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n13526) );
  NAND2_X1 U15179 ( .A1(n13523), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n13525) );
  NAND2_X1 U15180 ( .A1(n10328), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n13524) );
  INV_X1 U15181 ( .A(n13866), .ZN(n14671) );
  AOI22_X1 U15182 ( .A1(n14672), .A2(n14883), .B1(n14723), .B2(n14671), .ZN(
        n13527) );
  INV_X1 U15183 ( .A(n14993), .ZN(n14879) );
  INV_X1 U15184 ( .A(n14964), .ZN(n14791) );
  AOI22_X1 U15185 ( .A1(n13531), .A2(n14929), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n14938), .ZN(n13532) );
  OAI21_X1 U15186 ( .B1(n13871), .B2(n14932), .A(n13532), .ZN(n13551) );
  XNOR2_X1 U15187 ( .A(n14981), .B(n14858), .ZN(n14851) );
  AND2_X1 U15188 ( .A1(n13534), .A2(n13533), .ZN(n14918) );
  OR2_X1 U15189 ( .A1(n15005), .A2(n14673), .ZN(n13535) );
  NAND2_X1 U15190 ( .A1(n14893), .A2(n14896), .ZN(n13537) );
  OR2_X1 U15191 ( .A1(n15001), .A2(n14884), .ZN(n13536) );
  NOR2_X1 U15192 ( .A1(n14993), .A2(n14857), .ZN(n13538) );
  NAND2_X1 U15193 ( .A1(n14881), .A2(n14857), .ZN(n13539) );
  AND2_X1 U15194 ( .A1(n14987), .A2(n14886), .ZN(n13540) );
  NAND2_X1 U15195 ( .A1(n14981), .A2(n14858), .ZN(n13541) );
  OR2_X1 U15196 ( .A1(n14975), .A2(n14837), .ZN(n13542) );
  INV_X1 U15197 ( .A(n14794), .ZN(n13543) );
  NAND2_X1 U15198 ( .A1(n14784), .A2(n13543), .ZN(n13545) );
  OR2_X1 U15199 ( .A1(n14964), .A2(n14811), .ZN(n13544) );
  NAND2_X1 U15200 ( .A1(n14769), .A2(n14771), .ZN(n13547) );
  OR2_X1 U15201 ( .A1(n14959), .A2(n14795), .ZN(n13546) );
  NAND2_X1 U15202 ( .A1(n14954), .A2(n14774), .ZN(n13548) );
  NAND2_X1 U15203 ( .A1(n14736), .A2(n13549), .ZN(n13550) );
  NAND2_X1 U15204 ( .A1(n13553), .A2(n13552), .ZN(n13554) );
  AOI22_X1 U15205 ( .A1(n15349), .A2(n13578), .B1(n13265), .B2(n15180), .ZN(
        n13556) );
  XNOR2_X1 U15206 ( .A(n13556), .B(n13268), .ZN(n13559) );
  AOI22_X1 U15207 ( .A1(n15349), .A2(n13265), .B1(n13572), .B2(n15180), .ZN(
        n13558) );
  XNOR2_X1 U15208 ( .A(n13559), .B(n13558), .ZN(n15096) );
  INV_X1 U15209 ( .A(n15096), .ZN(n13557) );
  NAND2_X1 U15210 ( .A1(n13559), .A2(n13558), .ZN(n13560) );
  NAND2_X1 U15211 ( .A1(n15093), .A2(n13560), .ZN(n15138) );
  OAI22_X1 U15212 ( .A1(n15503), .A2(n13588), .B1(n8259), .B2(n13587), .ZN(
        n13565) );
  NAND2_X1 U15213 ( .A1(n15334), .A2(n13578), .ZN(n13562) );
  NAND2_X1 U15214 ( .A1(n15311), .A2(n13265), .ZN(n13561) );
  NAND2_X1 U15215 ( .A1(n13562), .A2(n13561), .ZN(n13563) );
  XNOR2_X1 U15216 ( .A(n13563), .B(n13268), .ZN(n13564) );
  XOR2_X1 U15217 ( .A(n13565), .B(n13564), .Z(n15139) );
  NAND2_X1 U15218 ( .A1(n15138), .A2(n15139), .ZN(n15137) );
  INV_X1 U15219 ( .A(n13564), .ZN(n13567) );
  INV_X1 U15220 ( .A(n13565), .ZN(n13566) );
  NAND2_X1 U15221 ( .A1(n13567), .A2(n13566), .ZN(n13568) );
  NAND2_X1 U15222 ( .A1(n15137), .A2(n13568), .ZN(n15121) );
  NAND2_X1 U15223 ( .A1(n15498), .A2(n13578), .ZN(n13570) );
  NAND2_X1 U15224 ( .A1(n15329), .A2(n13265), .ZN(n13569) );
  NAND2_X1 U15225 ( .A1(n13570), .A2(n13569), .ZN(n13571) );
  XNOR2_X1 U15226 ( .A(n13571), .B(n13268), .ZN(n13573) );
  AOI22_X1 U15227 ( .A1(n15498), .A2(n13265), .B1(n13572), .B2(n15329), .ZN(
        n13574) );
  XNOR2_X1 U15228 ( .A(n13573), .B(n13574), .ZN(n15122) );
  NAND2_X1 U15229 ( .A1(n15121), .A2(n15122), .ZN(n13577) );
  INV_X1 U15230 ( .A(n13573), .ZN(n13575) );
  NAND2_X1 U15231 ( .A1(n13575), .A2(n13574), .ZN(n13576) );
  NAND2_X1 U15232 ( .A1(n13577), .A2(n13576), .ZN(n15165) );
  OAI22_X1 U15233 ( .A1(n15301), .A2(n13588), .B1(n15125), .B2(n13587), .ZN(
        n13583) );
  NAND2_X1 U15234 ( .A1(n15491), .A2(n13578), .ZN(n13580) );
  NAND2_X1 U15235 ( .A1(n15312), .A2(n13265), .ZN(n13579) );
  NAND2_X1 U15236 ( .A1(n13580), .A2(n13579), .ZN(n13581) );
  XNOR2_X1 U15237 ( .A(n13581), .B(n11815), .ZN(n13582) );
  XOR2_X1 U15238 ( .A(n13583), .B(n13582), .Z(n15166) );
  INV_X1 U15239 ( .A(n13582), .ZN(n13585) );
  INV_X1 U15240 ( .A(n13583), .ZN(n13584) );
  NAND2_X1 U15241 ( .A1(n13585), .A2(n13584), .ZN(n13586) );
  OAI22_X1 U15242 ( .A1(n15485), .A2(n13588), .B1(n15171), .B2(n13587), .ZN(
        n13591) );
  OAI22_X1 U15243 ( .A1(n15485), .A2(n13594), .B1(n15171), .B2(n13588), .ZN(
        n13589) );
  XNOR2_X1 U15244 ( .A(n13589), .B(n11815), .ZN(n13590) );
  INV_X1 U15245 ( .A(n13590), .ZN(n13593) );
  INV_X1 U15246 ( .A(n13591), .ZN(n13592) );
  OAI22_X1 U15247 ( .A1(n15480), .A2(n13594), .B1(n15079), .B2(n13588), .ZN(
        n13597) );
  OAI22_X1 U15248 ( .A1(n15480), .A2(n13588), .B1(n15079), .B2(n13587), .ZN(
        n13595) );
  XNOR2_X1 U15249 ( .A(n13595), .B(n11815), .ZN(n13596) );
  XOR2_X1 U15250 ( .A(n13597), .B(n13596), .Z(n13598) );
  OAI22_X1 U15251 ( .A1(n15171), .A2(n15406), .B1(n13599), .B2(n15408), .ZN(
        n15263) );
  AOI22_X1 U15252 ( .A1(n15153), .A2(n15263), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13600) );
  OAI21_X1 U15253 ( .B1(n15272), .B2(n16361), .A(n13600), .ZN(n13601) );
  AOI21_X1 U15254 ( .B1(n15274), .B2(n15173), .A(n13601), .ZN(n13602) );
  OAI21_X1 U15255 ( .B1(n13603), .B2(n15175), .A(n13602), .ZN(P1_U3220) );
  OAI222_X1 U15256 ( .A1(n15604), .A2(n13605), .B1(P1_U3086), .B2(n8381), .C1(
        n13604), .C2(n15597), .ZN(P1_U3325) );
  NAND2_X1 U15257 ( .A1(n15051), .A2(n13615), .ZN(n13608) );
  OR2_X1 U15258 ( .A1(n13618), .A2(n13606), .ZN(n13607) );
  INV_X1 U15259 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n13611) );
  NAND2_X1 U15260 ( .A1(n13523), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n13610) );
  NAND2_X1 U15261 ( .A1(n13517), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n13609) );
  OAI211_X1 U15262 ( .C1(n13612), .C2(n13611), .A(n13610), .B(n13609), .ZN(
        n14724) );
  INV_X1 U15263 ( .A(n14724), .ZN(n13613) );
  NAND2_X1 U15264 ( .A1(n14725), .A2(n13613), .ZN(n13892) );
  OR2_X1 U15265 ( .A1(n14725), .A2(n13613), .ZN(n13614) );
  NAND2_X1 U15266 ( .A1(n13892), .A2(n13614), .ZN(n13883) );
  INV_X1 U15267 ( .A(n13883), .ZN(n13657) );
  NAND2_X1 U15268 ( .A1(n13616), .A2(n13615), .ZN(n13620) );
  OR2_X1 U15269 ( .A1(n13618), .A2(n13617), .ZN(n13619) );
  INV_X1 U15270 ( .A(n14942), .ZN(n13867) );
  XNOR2_X1 U15271 ( .A(n13867), .B(n13866), .ZN(n13655) );
  XNOR2_X1 U15272 ( .A(n14987), .B(n14886), .ZN(n14862) );
  AND2_X1 U15273 ( .A1(n13621), .A2(n8074), .ZN(n13624) );
  NAND4_X1 U15274 ( .A1(n13625), .A2(n13624), .A3(n13623), .A4(n13622), .ZN(
        n13627) );
  NOR2_X1 U15275 ( .A1(n13627), .A2(n13626), .ZN(n13630) );
  NAND4_X1 U15276 ( .A1(n13629), .A2(n13630), .A3(n13631), .A4(n13628), .ZN(
        n13632) );
  OR4_X1 U15277 ( .A1(n13635), .A2(n13634), .A3(n13633), .A4(n13632), .ZN(
        n13636) );
  OR4_X1 U15278 ( .A1(n13639), .A2(n13638), .A3(n13637), .A4(n13636), .ZN(
        n13640) );
  NOR2_X1 U15279 ( .A1(n13641), .A2(n13640), .ZN(n13644) );
  NAND4_X1 U15280 ( .A1(n13645), .A2(n13644), .A3(n13643), .A4(n13642), .ZN(
        n13646) );
  NOR2_X1 U15281 ( .A1(n14896), .A2(n13646), .ZN(n13647) );
  NAND4_X1 U15282 ( .A1(n14862), .A2(n13647), .A3(n14881), .A4(n14919), .ZN(
        n13648) );
  NOR2_X1 U15283 ( .A1(n14807), .A2(n13648), .ZN(n13649) );
  NAND4_X1 U15284 ( .A1(n14794), .A2(n13649), .A3(n14851), .A4(n14818), .ZN(
        n13650) );
  NOR2_X1 U15285 ( .A1(n14771), .A2(n13650), .ZN(n13652) );
  NAND4_X1 U15286 ( .A1(n13653), .A2(n13652), .A3(n13651), .A4(n14753), .ZN(
        n13654) );
  NOR2_X1 U15287 ( .A1(n13655), .A2(n13654), .ZN(n13656) );
  NAND2_X1 U15288 ( .A1(n13657), .A2(n13656), .ZN(n13918) );
  NAND3_X1 U15289 ( .A1(n13900), .A2(n13658), .A3(n13899), .ZN(n13911) );
  INV_X1 U15290 ( .A(n13911), .ZN(n13661) );
  MUX2_X1 U15291 ( .A(n13899), .B(n13902), .S(n13912), .Z(n13660) );
  NAND2_X1 U15292 ( .A1(n13900), .A2(n13658), .ZN(n13659) );
  NOR2_X1 U15293 ( .A1(n13660), .A2(n13659), .ZN(n13909) );
  AOI21_X1 U15294 ( .B1(n13918), .B2(n13661), .A(n13909), .ZN(n13921) );
  NAND2_X1 U15295 ( .A1(n13664), .A2(n13870), .ZN(n13673) );
  NAND2_X1 U15296 ( .A1(n13669), .A2(n13667), .ZN(n13671) );
  NOR2_X1 U15297 ( .A1(n13666), .A2(n13665), .ZN(n13670) );
  NAND2_X1 U15298 ( .A1(n13673), .A2(n13672), .ZN(n13683) );
  NAND2_X1 U15299 ( .A1(n14691), .A2(n13716), .ZN(n13675) );
  NAND2_X1 U15300 ( .A1(n7432), .A2(n13676), .ZN(n13674) );
  NAND2_X1 U15301 ( .A1(n13675), .A2(n13674), .ZN(n13682) );
  AOI22_X1 U15302 ( .A1(n7423), .A2(n13676), .B1(n13716), .B2(n14626), .ZN(
        n13685) );
  NAND2_X1 U15303 ( .A1(n7423), .A2(n13716), .ZN(n13679) );
  NAND2_X1 U15304 ( .A1(n13679), .A2(n13678), .ZN(n13684) );
  OAI22_X1 U15305 ( .A1(n13683), .A2(n13682), .B1(n13685), .B2(n13684), .ZN(
        n13688) );
  AOI22_X1 U15306 ( .A1(n14691), .A2(n13676), .B1(n13716), .B2(n7432), .ZN(
        n13681) );
  AOI21_X1 U15307 ( .B1(n13683), .B2(n13682), .A(n13681), .ZN(n13687) );
  NAND2_X1 U15308 ( .A1(n13685), .A2(n13684), .ZN(n13686) );
  NAND2_X1 U15309 ( .A1(n14689), .A2(n13716), .ZN(n13690) );
  NAND2_X1 U15310 ( .A1(n13695), .A2(n13676), .ZN(n13689) );
  NAND2_X1 U15311 ( .A1(n13690), .A2(n13689), .ZN(n13697) );
  AOI22_X1 U15312 ( .A1(n14688), .A2(n13676), .B1(n13691), .B2(n13716), .ZN(
        n13701) );
  NAND2_X1 U15313 ( .A1(n14688), .A2(n13857), .ZN(n13693) );
  BUF_X4 U15314 ( .A(n13870), .Z(n13868) );
  NAND2_X1 U15315 ( .A1(n13691), .A2(n13868), .ZN(n13692) );
  NAND2_X1 U15316 ( .A1(n13693), .A2(n13692), .ZN(n13700) );
  OAI22_X1 U15317 ( .A1(n13698), .A2(n13697), .B1(n13701), .B2(n13700), .ZN(
        n13694) );
  AOI22_X1 U15318 ( .A1(n14689), .A2(n13676), .B1(n13857), .B2(n13695), .ZN(
        n13696) );
  AOI21_X1 U15319 ( .B1(n13698), .B2(n13697), .A(n13696), .ZN(n13699) );
  NAND2_X1 U15320 ( .A1(n13701), .A2(n13700), .ZN(n13702) );
  NAND2_X1 U15321 ( .A1(n13703), .A2(n13702), .ZN(n13709) );
  NAND2_X1 U15322 ( .A1(n13706), .A2(n13676), .ZN(n13705) );
  NAND2_X1 U15323 ( .A1(n14687), .A2(n13857), .ZN(n13704) );
  NAND2_X1 U15324 ( .A1(n13705), .A2(n13704), .ZN(n13708) );
  AOI22_X1 U15325 ( .A1(n13706), .A2(n13857), .B1(n14687), .B2(n13868), .ZN(
        n13707) );
  NAND2_X1 U15326 ( .A1(n16122), .A2(n13857), .ZN(n13711) );
  NAND2_X1 U15327 ( .A1(n14686), .A2(n13868), .ZN(n13710) );
  NAND2_X1 U15328 ( .A1(n13711), .A2(n13710), .ZN(n13713) );
  AOI22_X1 U15329 ( .A1(n16122), .A2(n13868), .B1(n13857), .B2(n14686), .ZN(
        n13712) );
  NAND2_X1 U15330 ( .A1(n13717), .A2(n13868), .ZN(n13715) );
  NAND2_X1 U15331 ( .A1(n14685), .A2(n13857), .ZN(n13714) );
  NAND2_X1 U15332 ( .A1(n13715), .A2(n13714), .ZN(n13722) );
  NAND2_X1 U15333 ( .A1(n13721), .A2(n13722), .ZN(n13720) );
  NAND2_X1 U15334 ( .A1(n13717), .A2(n13857), .ZN(n13718) );
  OAI21_X1 U15335 ( .B1(n14649), .B2(n13891), .A(n13718), .ZN(n13719) );
  NAND2_X1 U15336 ( .A1(n13720), .A2(n13719), .ZN(n13726) );
  NAND2_X1 U15337 ( .A1(n13724), .A2(n13723), .ZN(n13725) );
  NAND2_X1 U15338 ( .A1(n13729), .A2(n13891), .ZN(n13728) );
  NAND2_X1 U15339 ( .A1(n14684), .A2(n13868), .ZN(n13727) );
  AOI22_X1 U15340 ( .A1(n13729), .A2(n13868), .B1(n13891), .B2(n14684), .ZN(
        n13730) );
  INV_X1 U15341 ( .A(n13730), .ZN(n13731) );
  NAND2_X1 U15342 ( .A1(n13734), .A2(n13868), .ZN(n13733) );
  NAND2_X1 U15343 ( .A1(n14682), .A2(n13891), .ZN(n13732) );
  NAND2_X1 U15344 ( .A1(n13733), .A2(n13732), .ZN(n13740) );
  NAND2_X1 U15345 ( .A1(n13734), .A2(n13891), .ZN(n13735) );
  OAI21_X1 U15346 ( .B1(n13736), .B2(n13891), .A(n13735), .ZN(n13737) );
  NAND2_X1 U15347 ( .A1(n13738), .A2(n13737), .ZN(n13744) );
  INV_X1 U15348 ( .A(n13739), .ZN(n13742) );
  INV_X1 U15349 ( .A(n13740), .ZN(n13741) );
  NAND2_X1 U15350 ( .A1(n13742), .A2(n13741), .ZN(n13743) );
  NAND2_X1 U15351 ( .A1(n13747), .A2(n13857), .ZN(n13746) );
  NAND2_X1 U15352 ( .A1(n14681), .A2(n13868), .ZN(n13745) );
  NAND2_X1 U15353 ( .A1(n13746), .A2(n13745), .ZN(n13749) );
  AOI22_X1 U15354 ( .A1(n13747), .A2(n13868), .B1(n13891), .B2(n14681), .ZN(
        n13748) );
  NAND2_X1 U15355 ( .A1(n13753), .A2(n13868), .ZN(n13752) );
  NAND2_X1 U15356 ( .A1(n14680), .A2(n13857), .ZN(n13751) );
  NAND2_X1 U15357 ( .A1(n13752), .A2(n13751), .ZN(n13755) );
  AOI22_X1 U15358 ( .A1(n13753), .A2(n13891), .B1(n14680), .B2(n13868), .ZN(
        n13754) );
  NAND2_X1 U15359 ( .A1(n13758), .A2(n13857), .ZN(n13757) );
  NAND2_X1 U15360 ( .A1(n14679), .A2(n13868), .ZN(n13756) );
  NAND2_X1 U15361 ( .A1(n13757), .A2(n13756), .ZN(n13764) );
  NAND2_X1 U15362 ( .A1(n13758), .A2(n13868), .ZN(n13759) );
  OAI21_X1 U15363 ( .B1(n13760), .B2(n13870), .A(n13759), .ZN(n13761) );
  INV_X1 U15364 ( .A(n13763), .ZN(n13766) );
  INV_X1 U15365 ( .A(n13764), .ZN(n13765) );
  NAND2_X1 U15366 ( .A1(n13766), .A2(n13765), .ZN(n13767) );
  NAND2_X1 U15367 ( .A1(n13770), .A2(n13868), .ZN(n13769) );
  NAND2_X1 U15368 ( .A1(n14678), .A2(n13857), .ZN(n13768) );
  AOI22_X1 U15369 ( .A1(n13770), .A2(n13891), .B1(n14678), .B2(n13868), .ZN(
        n13771) );
  NAND2_X1 U15370 ( .A1(n13774), .A2(n13857), .ZN(n13773) );
  NAND2_X1 U15371 ( .A1(n14677), .A2(n13868), .ZN(n13772) );
  NAND2_X1 U15372 ( .A1(n13774), .A2(n13868), .ZN(n13775) );
  OAI21_X1 U15373 ( .B1(n13776), .B2(n13870), .A(n13775), .ZN(n13777) );
  NAND2_X1 U15374 ( .A1(n15025), .A2(n13868), .ZN(n13779) );
  NAND2_X1 U15375 ( .A1(n14676), .A2(n13857), .ZN(n13778) );
  NAND2_X1 U15376 ( .A1(n13779), .A2(n13778), .ZN(n13782) );
  AOI22_X1 U15377 ( .A1(n15025), .A2(n13891), .B1(n14676), .B2(n13868), .ZN(
        n13780) );
  AOI21_X1 U15378 ( .B1(n13783), .B2(n13782), .A(n13780), .ZN(n13781) );
  NOR2_X1 U15379 ( .A1(n13783), .A2(n13782), .ZN(n13784) );
  NAND2_X1 U15380 ( .A1(n15017), .A2(n13891), .ZN(n13786) );
  NAND2_X1 U15381 ( .A1(n14675), .A2(n13868), .ZN(n13785) );
  NAND2_X1 U15382 ( .A1(n15017), .A2(n13868), .ZN(n13787) );
  OAI21_X1 U15383 ( .B1(n14597), .B2(n13870), .A(n13787), .ZN(n13788) );
  NAND2_X1 U15384 ( .A1(n15011), .A2(n13868), .ZN(n13790) );
  NAND2_X1 U15385 ( .A1(n14674), .A2(n13891), .ZN(n13789) );
  NAND2_X1 U15386 ( .A1(n13790), .A2(n13789), .ZN(n13793) );
  AOI22_X1 U15387 ( .A1(n15011), .A2(n13891), .B1(n14674), .B2(n13868), .ZN(
        n13791) );
  AOI21_X1 U15388 ( .B1(n13794), .B2(n13793), .A(n13791), .ZN(n13792) );
  NAND2_X1 U15389 ( .A1(n15005), .A2(n13891), .ZN(n13796) );
  NAND2_X1 U15390 ( .A1(n14673), .A2(n13868), .ZN(n13795) );
  AOI22_X1 U15391 ( .A1(n15005), .A2(n13868), .B1(n13891), .B2(n14673), .ZN(
        n13797) );
  NAND2_X1 U15392 ( .A1(n15001), .A2(n13868), .ZN(n13799) );
  NAND2_X1 U15393 ( .A1(n14884), .A2(n13891), .ZN(n13798) );
  NAND2_X1 U15394 ( .A1(n13799), .A2(n13798), .ZN(n13804) );
  NAND2_X1 U15395 ( .A1(n13803), .A2(n13804), .ZN(n13802) );
  NAND2_X1 U15396 ( .A1(n15001), .A2(n13891), .ZN(n13800) );
  OAI21_X1 U15397 ( .B1(n14917), .B2(n13857), .A(n13800), .ZN(n13801) );
  NAND2_X1 U15398 ( .A1(n13802), .A2(n13801), .ZN(n13808) );
  INV_X1 U15399 ( .A(n13803), .ZN(n13806) );
  INV_X1 U15400 ( .A(n13804), .ZN(n13805) );
  NAND2_X1 U15401 ( .A1(n13806), .A2(n13805), .ZN(n13807) );
  NAND2_X1 U15402 ( .A1(n14993), .A2(n13891), .ZN(n13810) );
  NAND2_X1 U15403 ( .A1(n14857), .A2(n13868), .ZN(n13809) );
  NAND2_X1 U15404 ( .A1(n13810), .A2(n13809), .ZN(n13812) );
  AOI22_X1 U15405 ( .A1(n14993), .A2(n13868), .B1(n13857), .B2(n14857), .ZN(
        n13811) );
  AOI21_X1 U15406 ( .B1(n13813), .B2(n13812), .A(n13811), .ZN(n13814) );
  NAND2_X1 U15407 ( .A1(n14987), .A2(n13868), .ZN(n13816) );
  NAND2_X1 U15408 ( .A1(n14886), .A2(n13891), .ZN(n13815) );
  NAND2_X1 U15409 ( .A1(n13816), .A2(n13815), .ZN(n13820) );
  NAND2_X1 U15410 ( .A1(n14987), .A2(n13891), .ZN(n13818) );
  NAND2_X1 U15411 ( .A1(n14886), .A2(n13868), .ZN(n13817) );
  NAND2_X1 U15412 ( .A1(n13818), .A2(n13817), .ZN(n13819) );
  INV_X1 U15413 ( .A(n13820), .ZN(n13821) );
  NAND2_X1 U15414 ( .A1(n14981), .A2(n13891), .ZN(n13823) );
  NAND2_X1 U15415 ( .A1(n14858), .A2(n13868), .ZN(n13822) );
  NAND2_X1 U15416 ( .A1(n13823), .A2(n13822), .ZN(n13825) );
  AOI22_X1 U15417 ( .A1(n14981), .A2(n13868), .B1(n13891), .B2(n14858), .ZN(
        n13824) );
  AOI21_X1 U15418 ( .B1(n13826), .B2(n13825), .A(n13824), .ZN(n13828) );
  NOR2_X1 U15419 ( .A1(n13826), .A2(n13825), .ZN(n13827) );
  NAND2_X1 U15420 ( .A1(n14975), .A2(n13868), .ZN(n13830) );
  NAND2_X1 U15421 ( .A1(n14837), .A2(n13891), .ZN(n13829) );
  NAND2_X1 U15422 ( .A1(n13830), .A2(n13829), .ZN(n13834) );
  NAND2_X1 U15423 ( .A1(n14975), .A2(n13891), .ZN(n13831) );
  OAI21_X1 U15424 ( .B1(n14620), .B2(n13857), .A(n13831), .ZN(n13832) );
  NAND2_X1 U15425 ( .A1(n14969), .A2(n13891), .ZN(n13836) );
  NAND2_X1 U15426 ( .A1(n14819), .A2(n13868), .ZN(n13835) );
  AOI22_X1 U15427 ( .A1(n14969), .A2(n13868), .B1(n13857), .B2(n14819), .ZN(
        n13837) );
  NAND2_X1 U15428 ( .A1(n14964), .A2(n13868), .ZN(n13840) );
  NAND2_X1 U15429 ( .A1(n14811), .A2(n13891), .ZN(n13839) );
  NAND2_X1 U15430 ( .A1(n13840), .A2(n13839), .ZN(n13842) );
  AOI22_X1 U15431 ( .A1(n14964), .A2(n13891), .B1(n14811), .B2(n13868), .ZN(
        n13841) );
  NAND2_X1 U15432 ( .A1(n14959), .A2(n13891), .ZN(n13845) );
  NAND2_X1 U15433 ( .A1(n14795), .A2(n13868), .ZN(n13844) );
  NAND2_X1 U15434 ( .A1(n13845), .A2(n13844), .ZN(n13850) );
  NAND2_X1 U15435 ( .A1(n14959), .A2(n13868), .ZN(n13847) );
  NAND2_X1 U15436 ( .A1(n14795), .A2(n13891), .ZN(n13846) );
  NAND2_X1 U15437 ( .A1(n13847), .A2(n13846), .ZN(n13848) );
  NAND2_X1 U15438 ( .A1(n13849), .A2(n13848), .ZN(n13854) );
  INV_X1 U15439 ( .A(n13850), .ZN(n13851) );
  NAND2_X1 U15440 ( .A1(n13852), .A2(n13851), .ZN(n13853) );
  NAND2_X1 U15441 ( .A1(n14954), .A2(n13870), .ZN(n13856) );
  NAND2_X1 U15442 ( .A1(n14774), .A2(n13891), .ZN(n13855) );
  NAND2_X1 U15443 ( .A1(n13856), .A2(n13855), .ZN(n13859) );
  AOI22_X1 U15444 ( .A1(n14949), .A2(n13857), .B1(n14672), .B2(n13676), .ZN(
        n13875) );
  OAI22_X1 U15445 ( .A1(n7418), .A2(n13857), .B1(n14752), .B2(n13870), .ZN(
        n13874) );
  AOI22_X1 U15446 ( .A1(n14954), .A2(n13857), .B1(n14774), .B2(n13676), .ZN(
        n13858) );
  NOR2_X1 U15447 ( .A1(n13861), .A2(n8074), .ZN(n13864) );
  INV_X1 U15448 ( .A(n13862), .ZN(n13863) );
  AOI211_X1 U15449 ( .C1(n14724), .C2(n13868), .A(n13864), .B(n13863), .ZN(
        n13865) );
  OAI22_X1 U15450 ( .A1(n14942), .A2(n13870), .B1(n13866), .B2(n13865), .ZN(
        n13885) );
  AOI22_X1 U15451 ( .A1(n13867), .A2(n13868), .B1(n13857), .B2(n14671), .ZN(
        n13884) );
  AOI22_X1 U15452 ( .A1(n14944), .A2(n13868), .B1(n13857), .B2(n14740), .ZN(
        n13878) );
  OAI22_X1 U15453 ( .A1(n13871), .A2(n13870), .B1(n13869), .B2(n13857), .ZN(
        n13879) );
  AOI22_X1 U15454 ( .A1(n13885), .A2(n13884), .B1(n13878), .B2(n13879), .ZN(
        n13872) );
  NOR2_X1 U15455 ( .A1(n13872), .A2(n13883), .ZN(n13880) );
  INV_X1 U15456 ( .A(n13874), .ZN(n13877) );
  INV_X1 U15457 ( .A(n13875), .ZN(n13876) );
  OAI22_X1 U15458 ( .A1(n13879), .A2(n13878), .B1(n13877), .B2(n13876), .ZN(
        n13882) );
  INV_X1 U15459 ( .A(n13880), .ZN(n13881) );
  OAI21_X1 U15460 ( .B1(n13883), .B2(n13882), .A(n13881), .ZN(n13889) );
  INV_X1 U15461 ( .A(n13884), .ZN(n13887) );
  INV_X1 U15462 ( .A(n13885), .ZN(n13886) );
  NOR2_X1 U15463 ( .A1(n13892), .A2(n13891), .ZN(n13910) );
  NAND2_X1 U15464 ( .A1(n14724), .A2(n13857), .ZN(n13893) );
  NOR2_X1 U15465 ( .A1(n14725), .A2(n13893), .ZN(n13898) );
  AOI22_X1 U15466 ( .A1(n13895), .A2(n13902), .B1(n13894), .B2(n15711), .ZN(
        n13897) );
  NOR4_X1 U15467 ( .A1(n13910), .A2(n13898), .A3(n13897), .A4(n13896), .ZN(
        n13920) );
  NAND4_X1 U15468 ( .A1(n13900), .A2(P2_STATE_REG_SCAN_IN), .A3(n13899), .A4(
        n15711), .ZN(n13917) );
  AOI21_X1 U15469 ( .B1(n13903), .B2(n13902), .A(n13901), .ZN(n13908) );
  INV_X1 U15470 ( .A(n13904), .ZN(n13905) );
  NAND4_X1 U15471 ( .A1(n14883), .A2(n13906), .A3(n15647), .A4(n13905), .ZN(
        n13907) );
  AOI22_X1 U15472 ( .A1(n13910), .A2(n13909), .B1(n13908), .B2(n13907), .ZN(
        n13916) );
  INV_X1 U15473 ( .A(n13910), .ZN(n13913) );
  AOI21_X1 U15474 ( .B1(n13913), .B2(n13912), .A(n13911), .ZN(n13914) );
  NAND2_X1 U15475 ( .A1(n13914), .A2(n13918), .ZN(n13915) );
  OAI211_X1 U15476 ( .C1(n13918), .C2(n13917), .A(n13916), .B(n13915), .ZN(
        n13919) );
  INV_X1 U15477 ( .A(n13922), .ZN(n13923) );
  OAI222_X1 U15478 ( .A1(n13927), .A2(P3_U3151), .B1(n13926), .B2(n13925), 
        .C1(n13924), .C2(n13923), .ZN(P3_U3266) );
  AOI22_X1 U15479 ( .A1(n14351), .A2(n14034), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13930) );
  NAND2_X1 U15480 ( .A1(n14184), .A2(n14023), .ZN(n13929) );
  OAI211_X1 U15481 ( .C1(n14044), .C2(n14032), .A(n13930), .B(n13929), .ZN(
        n13931) );
  AOI21_X1 U15482 ( .B1(n14352), .B2(n16037), .A(n13931), .ZN(n13932) );
  OAI21_X1 U15483 ( .B1(n13933), .B2(n14041), .A(n13932), .ZN(P3_U3154) );
  OAI211_X1 U15484 ( .C1(n13936), .C2(n13935), .A(n13934), .B(n16041), .ZN(
        n13942) );
  AOI21_X1 U15485 ( .B1(n14034), .B2(n14049), .A(n13937), .ZN(n13938) );
  OAI21_X1 U15486 ( .B1(n14331), .B2(n14032), .A(n13938), .ZN(n13939) );
  AOI21_X1 U15487 ( .B1(n13940), .B2(n14023), .A(n13939), .ZN(n13941) );
  OAI211_X1 U15488 ( .C1(n14017), .C2(n14422), .A(n13942), .B(n13941), .ZN(
        P3_U3155) );
  XNOR2_X1 U15489 ( .A(n13943), .B(n13988), .ZN(n13990) );
  XNOR2_X1 U15490 ( .A(n13990), .B(n14252), .ZN(n13948) );
  AOI22_X1 U15491 ( .A1(n14360), .A2(n16039), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13945) );
  NAND2_X1 U15492 ( .A1(n14023), .A2(n14242), .ZN(n13944) );
  OAI211_X1 U15493 ( .C1(n14244), .C2(n14015), .A(n13945), .B(n13944), .ZN(
        n13946) );
  AOI21_X1 U15494 ( .B1(n14372), .B2(n16037), .A(n13946), .ZN(n13947) );
  OAI21_X1 U15495 ( .B1(n13948), .B2(n14041), .A(n13947), .ZN(P3_U3156) );
  XNOR2_X1 U15496 ( .A(n13950), .B(n13949), .ZN(n13955) );
  NAND2_X1 U15497 ( .A1(n16039), .A2(n14383), .ZN(n13951) );
  NAND2_X1 U15498 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n14151)
         );
  OAI211_X1 U15499 ( .C1(n14316), .C2(n14015), .A(n13951), .B(n14151), .ZN(
        n13953) );
  NOR2_X1 U15500 ( .A1(n14297), .A2(n14017), .ZN(n13952) );
  AOI211_X1 U15501 ( .C1(n14295), .C2(n14023), .A(n13953), .B(n13952), .ZN(
        n13954) );
  OAI21_X1 U15502 ( .B1(n13955), .B2(n14041), .A(n13954), .ZN(P3_U3159) );
  INV_X1 U15503 ( .A(n13956), .ZN(n13957) );
  NOR2_X1 U15504 ( .A1(n13958), .A2(n13957), .ZN(n13959) );
  XNOR2_X1 U15505 ( .A(n13960), .B(n13959), .ZN(n13965) );
  AOI22_X1 U15506 ( .A1(n14034), .A2(n14383), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13962) );
  NAND2_X1 U15507 ( .A1(n14023), .A2(n14266), .ZN(n13961) );
  OAI211_X1 U15508 ( .C1(n14244), .C2(n14032), .A(n13962), .B(n13961), .ZN(
        n13963) );
  AOI21_X1 U15509 ( .B1(n14385), .B2(n16037), .A(n13963), .ZN(n13964) );
  OAI21_X1 U15510 ( .B1(n13965), .B2(n14041), .A(n13964), .ZN(P3_U3163) );
  XOR2_X1 U15511 ( .A(n13967), .B(n13966), .Z(n13972) );
  AOI22_X1 U15512 ( .A1(n14351), .A2(n16039), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13969) );
  NAND2_X1 U15513 ( .A1(n14206), .A2(n14023), .ZN(n13968) );
  OAI211_X1 U15514 ( .C1(n14208), .C2(n14015), .A(n13969), .B(n13968), .ZN(
        n13970) );
  AOI21_X1 U15515 ( .B1(n14361), .B2(n16037), .A(n13970), .ZN(n13971) );
  OAI21_X1 U15516 ( .B1(n13972), .B2(n14041), .A(n13971), .ZN(P3_U3165) );
  XNOR2_X1 U15517 ( .A(n13974), .B(n13973), .ZN(n13980) );
  NAND2_X1 U15518 ( .A1(n16039), .A2(n14306), .ZN(n13976) );
  OAI211_X1 U15519 ( .C1(n14331), .C2(n14015), .A(n13976), .B(n13975), .ZN(
        n13978) );
  NOR2_X1 U15520 ( .A1(n14459), .A2(n14017), .ZN(n13977) );
  AOI211_X1 U15521 ( .C1(n14335), .C2(n14023), .A(n13978), .B(n13977), .ZN(
        n13979) );
  OAI21_X1 U15522 ( .B1(n13980), .B2(n14041), .A(n13979), .ZN(P3_U3166) );
  XNOR2_X1 U15523 ( .A(n13982), .B(n13981), .ZN(n13987) );
  NAND2_X1 U15524 ( .A1(n16039), .A2(n14290), .ZN(n13983) );
  NAND2_X1 U15525 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n14098)
         );
  OAI211_X1 U15526 ( .C1(n14317), .C2(n14015), .A(n13983), .B(n14098), .ZN(
        n13985) );
  NOR2_X1 U15527 ( .A1(n14455), .A2(n14017), .ZN(n13984) );
  AOI211_X1 U15528 ( .C1(n14321), .C2(n14023), .A(n13985), .B(n13984), .ZN(
        n13986) );
  OAI21_X1 U15529 ( .B1(n13987), .B2(n14041), .A(n13986), .ZN(P3_U3168) );
  OAI22_X1 U15530 ( .A1(n13990), .A2(n14223), .B1(n13989), .B2(n13988), .ZN(
        n13993) );
  XNOR2_X1 U15531 ( .A(n13991), .B(n14208), .ZN(n13992) );
  XNOR2_X1 U15532 ( .A(n13993), .B(n13992), .ZN(n13998) );
  AOI22_X1 U15533 ( .A1(n8346), .A2(n16039), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13995) );
  NAND2_X1 U15534 ( .A1(n14226), .A2(n14023), .ZN(n13994) );
  OAI211_X1 U15535 ( .C1(n14252), .C2(n14015), .A(n13995), .B(n13994), .ZN(
        n13996) );
  AOI21_X1 U15536 ( .B1(n14227), .B2(n16037), .A(n13996), .ZN(n13997) );
  OAI21_X1 U15537 ( .B1(n13998), .B2(n14041), .A(n13997), .ZN(P3_U3169) );
  XNOR2_X1 U15538 ( .A(n14000), .B(n13999), .ZN(n14005) );
  AOI22_X1 U15539 ( .A1(n16039), .A2(n14045), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n14002) );
  NAND2_X1 U15540 ( .A1(n14023), .A2(n14282), .ZN(n14001) );
  OAI211_X1 U15541 ( .C1(n14390), .C2(n14015), .A(n14002), .B(n14001), .ZN(
        n14003) );
  AOI21_X1 U15542 ( .B1(n14389), .B2(n16037), .A(n14003), .ZN(n14004) );
  OAI21_X1 U15543 ( .B1(n14005), .B2(n14041), .A(n14004), .ZN(P3_U3173) );
  XNOR2_X1 U15544 ( .A(n14006), .B(n14371), .ZN(n14011) );
  AOI22_X1 U15545 ( .A1(n14034), .A2(n14045), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n14008) );
  NAND2_X1 U15546 ( .A1(n14023), .A2(n14257), .ZN(n14007) );
  OAI211_X1 U15547 ( .C1(n14252), .C2(n14032), .A(n14008), .B(n14007), .ZN(
        n14009) );
  AOI21_X1 U15548 ( .B1(n14377), .B2(n16037), .A(n14009), .ZN(n14010) );
  OAI21_X1 U15549 ( .B1(n14011), .B2(n14041), .A(n14010), .ZN(P3_U3175) );
  XNOR2_X1 U15550 ( .A(n14013), .B(n14012), .ZN(n14021) );
  NAND2_X1 U15551 ( .A1(n16039), .A2(n14305), .ZN(n14014) );
  NAND2_X1 U15552 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n14126)
         );
  OAI211_X1 U15553 ( .C1(n14330), .C2(n14015), .A(n14014), .B(n14126), .ZN(
        n14019) );
  INV_X1 U15554 ( .A(n14016), .ZN(n14451) );
  NOR2_X1 U15555 ( .A1(n14451), .A2(n14017), .ZN(n14018) );
  AOI211_X1 U15556 ( .C1(n14310), .C2(n14023), .A(n14019), .B(n14018), .ZN(
        n14020) );
  OAI21_X1 U15557 ( .B1(n14021), .B2(n14041), .A(n14020), .ZN(P3_U3178) );
  AOI22_X1 U15558 ( .A1(n8346), .A2(n14034), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n14025) );
  NAND2_X1 U15559 ( .A1(n14195), .A2(n14023), .ZN(n14024) );
  OAI211_X1 U15560 ( .C1(n14174), .C2(n14032), .A(n14025), .B(n14024), .ZN(
        n14026) );
  AOI21_X1 U15561 ( .B1(n14356), .B2(n16037), .A(n14026), .ZN(n14027) );
  XNOR2_X1 U15562 ( .A(n14028), .B(n14047), .ZN(n14029) );
  XNOR2_X1 U15563 ( .A(n14030), .B(n14029), .ZN(n14042) );
  INV_X1 U15564 ( .A(n14463), .ZN(n14039) );
  INV_X1 U15565 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n14031) );
  NOR2_X1 U15566 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14031), .ZN(n14083) );
  NOR2_X1 U15567 ( .A1(n14032), .A2(n14317), .ZN(n14033) );
  AOI211_X1 U15568 ( .C1(n14034), .C2(n14048), .A(n14083), .B(n14033), .ZN(
        n14035) );
  OAI21_X1 U15569 ( .B1(n14037), .B2(n14036), .A(n14035), .ZN(n14038) );
  AOI21_X1 U15570 ( .B1(n14039), .B2(n16037), .A(n14038), .ZN(n14040) );
  OAI21_X1 U15571 ( .B1(n14042), .B2(n14041), .A(n14040), .ZN(P3_U3181) );
  MUX2_X1 U15572 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n14043), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U15573 ( .A(n14178), .B(P3_DATAO_REG_29__SCAN_IN), .S(n14055), .Z(
        P3_U3520) );
  MUX2_X1 U15574 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n9706), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U15575 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n14346), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U15576 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n14351), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U15577 ( .A(n8346), .B(P3_DATAO_REG_25__SCAN_IN), .S(n14055), .Z(
        P3_U3516) );
  MUX2_X1 U15578 ( .A(n14360), .B(P3_DATAO_REG_24__SCAN_IN), .S(n14055), .Z(
        P3_U3515) );
  MUX2_X1 U15579 ( .A(n14223), .B(P3_DATAO_REG_23__SCAN_IN), .S(n14055), .Z(
        P3_U3514) );
  MUX2_X1 U15580 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n14371), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U15581 ( .A(n14045), .B(P3_DATAO_REG_21__SCAN_IN), .S(n14055), .Z(
        P3_U3512) );
  MUX2_X1 U15582 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n14383), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U15583 ( .A(n14305), .B(P3_DATAO_REG_19__SCAN_IN), .S(n14055), .Z(
        P3_U3510) );
  MUX2_X1 U15584 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n14290), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U15585 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n14306), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U15586 ( .A(n14046), .B(P3_DATAO_REG_16__SCAN_IN), .S(n14055), .Z(
        P3_U3507) );
  MUX2_X1 U15587 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n14047), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U15588 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n14048), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U15589 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n14049), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U15590 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n14050), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U15591 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n14051), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U15592 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n14052), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U15593 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n14053), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U15594 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n14054), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U15595 ( .A(n14056), .B(P3_DATAO_REG_6__SCAN_IN), .S(n14055), .Z(
        P3_U3497) );
  MUX2_X1 U15596 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n14057), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U15597 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n14058), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U15598 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n16040), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U15599 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n14059), .S(P3_U3897), .Z(
        P3_U3491) );
  AOI21_X1 U15600 ( .B1(n9479), .B2(n14061), .A(n14060), .ZN(n14076) );
  OAI21_X1 U15601 ( .B1(n14064), .B2(n14063), .A(n14062), .ZN(n14074) );
  AOI21_X1 U15602 ( .B1(n14067), .B2(n14066), .A(n14065), .ZN(n14068) );
  NOR2_X1 U15603 ( .A1(n16009), .A2(n14068), .ZN(n14069) );
  AOI211_X1 U15604 ( .C1(n15646), .C2(P3_ADDR_REG_13__SCAN_IN), .A(n14070), 
        .B(n14069), .ZN(n14071) );
  OAI21_X1 U15605 ( .B1(n14072), .B2(n15997), .A(n14071), .ZN(n14073) );
  AOI21_X1 U15606 ( .B1(n14074), .B2(n16017), .A(n14073), .ZN(n14075) );
  OAI21_X1 U15607 ( .B1(n14076), .B2(n16013), .A(n14075), .ZN(P3_U3195) );
  AOI21_X1 U15608 ( .B1(n14079), .B2(n14078), .A(n14077), .ZN(n14093) );
  OAI21_X1 U15609 ( .B1(n14082), .B2(n14081), .A(n14080), .ZN(n14091) );
  AOI21_X1 U15610 ( .B1(n15646), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n14083), 
        .ZN(n14084) );
  OAI21_X1 U15611 ( .B1(n15997), .B2(n14085), .A(n14084), .ZN(n14090) );
  AOI21_X1 U15612 ( .B1(n14416), .B2(n14087), .A(n14086), .ZN(n14088) );
  NOR2_X1 U15613 ( .A1(n14088), .A2(n16013), .ZN(n14089) );
  AOI211_X1 U15614 ( .C1(n16017), .C2(n14091), .A(n14090), .B(n14089), .ZN(
        n14092) );
  OAI21_X1 U15615 ( .B1(n14093), .B2(n16009), .A(n14092), .ZN(P3_U3197) );
  OR2_X1 U15616 ( .A1(n14094), .A2(n14412), .ZN(n14095) );
  NOR2_X1 U15617 ( .A1(n14408), .A2(n14097), .ZN(n14127) );
  AOI21_X1 U15618 ( .B1(n14408), .B2(n14097), .A(n14127), .ZN(n14114) );
  INV_X1 U15619 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n15939) );
  OAI21_X1 U15620 ( .B1(n16027), .B2(n15939), .A(n14098), .ZN(n14105) );
  MUX2_X1 U15621 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n14141), .Z(n14121) );
  XNOR2_X1 U15622 ( .A(n14121), .B(n14129), .ZN(n14102) );
  NOR2_X1 U15623 ( .A1(n14103), .A2(n14102), .ZN(n14120) );
  AOI211_X1 U15624 ( .C1(n14103), .C2(n14102), .A(n15960), .B(n14120), .ZN(
        n14104) );
  AOI211_X1 U15625 ( .C1(n16020), .C2(n7984), .A(n14105), .B(n14104), .ZN(
        n14113) );
  INV_X1 U15626 ( .A(n14109), .ZN(n14108) );
  NOR2_X1 U15627 ( .A1(n14108), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n14111) );
  OAI21_X1 U15628 ( .B1(n14111), .B2(n14115), .A(n15973), .ZN(n14112) );
  OAI211_X1 U15629 ( .C1(n14114), .C2(n16013), .A(n14113), .B(n14112), .ZN(
        P3_U3199) );
  NOR2_X1 U15630 ( .A1(n7984), .A2(n7489), .ZN(n14116) );
  NAND2_X1 U15631 ( .A1(P3_REG2_REG_18__SCAN_IN), .A2(n14148), .ZN(n14117) );
  OAI21_X1 U15632 ( .B1(n14148), .B2(P3_REG2_REG_18__SCAN_IN), .A(n14117), 
        .ZN(n14118) );
  NOR2_X1 U15633 ( .A1(n14119), .A2(n14118), .ZN(n14147) );
  AOI21_X1 U15634 ( .B1(n14119), .B2(n14118), .A(n14147), .ZN(n14134) );
  MUX2_X1 U15635 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n14141), .Z(n14123) );
  AOI21_X1 U15636 ( .B1(n14121), .B2(n14129), .A(n14120), .ZN(n14140) );
  XNOR2_X1 U15637 ( .A(n14140), .B(n14139), .ZN(n14122) );
  NOR2_X1 U15638 ( .A1(n14122), .A2(n14123), .ZN(n14138) );
  AOI21_X1 U15639 ( .B1(n14123), .B2(n14122), .A(n14138), .ZN(n14124) );
  INV_X1 U15640 ( .A(n14124), .ZN(n14132) );
  NAND2_X1 U15641 ( .A1(n15646), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n14125) );
  OAI211_X1 U15642 ( .C1(n15997), .C2(n14148), .A(n14126), .B(n14125), .ZN(
        n14131) );
  NAND2_X1 U15643 ( .A1(n14148), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n14135) );
  OAI21_X1 U15644 ( .B1(n14148), .B2(P3_REG1_REG_18__SCAN_IN), .A(n14135), 
        .ZN(n14130) );
  OAI21_X1 U15645 ( .B1(n14134), .B2(n16009), .A(n14133), .ZN(P3_U3200) );
  NAND2_X1 U15646 ( .A1(n14136), .A2(n14135), .ZN(n14137) );
  XNOR2_X1 U15647 ( .A(n14145), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n14142) );
  XNOR2_X1 U15648 ( .A(n14137), .B(n14142), .ZN(n14155) );
  XNOR2_X1 U15649 ( .A(n14145), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n14146) );
  MUX2_X1 U15650 ( .A(n14146), .B(n14142), .S(n14141), .Z(n14143) );
  XNOR2_X1 U15651 ( .A(n14144), .B(n14143), .ZN(n14153) );
  NOR2_X1 U15652 ( .A1(n15997), .A2(n14145), .ZN(n14152) );
  INV_X1 U15653 ( .A(n14146), .ZN(n14149) );
  NAND2_X1 U15654 ( .A1(n15646), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n14150) );
  OAI21_X1 U15655 ( .B1(n14155), .B2(n16013), .A(n14154), .ZN(P3_U3201) );
  INV_X1 U15656 ( .A(n14156), .ZN(n14425) );
  AOI21_X1 U15657 ( .B1(n16094), .B2(n14164), .A(n14341), .ZN(n14159) );
  OR2_X1 U15658 ( .A1(n14158), .A2(n14157), .ZN(n14423) );
  NAND2_X1 U15659 ( .A1(n14159), .A2(n14423), .ZN(n14161) );
  OAI21_X1 U15660 ( .B1(P3_REG2_REG_31__SCAN_IN), .B2(n16100), .A(n14161), 
        .ZN(n14160) );
  OAI21_X1 U15661 ( .B1(n14425), .B2(n14337), .A(n14160), .ZN(P3_U3202) );
  OAI21_X1 U15662 ( .B1(P3_REG2_REG_30__SCAN_IN), .B2(n16100), .A(n14161), 
        .ZN(n14162) );
  OAI21_X1 U15663 ( .B1(n14428), .B2(n14337), .A(n14162), .ZN(P3_U3203) );
  INV_X1 U15664 ( .A(n14163), .ZN(n14170) );
  AOI22_X1 U15665 ( .A1(n14164), .A2(n16094), .B1(P3_REG2_REG_29__SCAN_IN), 
        .B2(n14341), .ZN(n14165) );
  OAI21_X1 U15666 ( .B1(n14166), .B2(n14337), .A(n14165), .ZN(n14167) );
  AOI21_X1 U15667 ( .B1(n14168), .B2(n14339), .A(n14167), .ZN(n14169) );
  OAI21_X1 U15668 ( .B1(n14170), .B2(n14341), .A(n14169), .ZN(P3_U3204) );
  XOR2_X1 U15669 ( .A(n14176), .B(n14171), .Z(n14350) );
  AOI22_X1 U15670 ( .A1(n14172), .A2(n16094), .B1(n14341), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n14173) );
  OAI21_X1 U15671 ( .B1(n14174), .B2(n14284), .A(n14173), .ZN(n14180) );
  INV_X1 U15672 ( .A(n14175), .ZN(n14177) );
  OAI21_X1 U15673 ( .B1(n14350), .B2(n14288), .A(n14181), .ZN(P3_U3205) );
  XNOR2_X1 U15674 ( .A(n14182), .B(n14188), .ZN(n14183) );
  AOI22_X1 U15675 ( .A1(n14183), .A2(n9714), .B1(n14304), .B2(n9706), .ZN(
        n14354) );
  AOI22_X1 U15676 ( .A1(n14184), .A2(n16094), .B1(n14341), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n14185) );
  OAI21_X1 U15677 ( .B1(n14186), .B2(n14284), .A(n14185), .ZN(n14191) );
  AOI21_X1 U15678 ( .B1(n14189), .B2(n14188), .A(n14187), .ZN(n14355) );
  NOR2_X1 U15679 ( .A1(n14355), .A2(n14288), .ZN(n14190) );
  AOI211_X1 U15680 ( .C1(n16096), .C2(n14352), .A(n14191), .B(n14190), .ZN(
        n14192) );
  OAI21_X1 U15681 ( .B1(n14341), .B2(n14354), .A(n14192), .ZN(P3_U3206) );
  XNOR2_X1 U15682 ( .A(n14193), .B(n14199), .ZN(n14194) );
  AOI22_X1 U15683 ( .A1(n14194), .A2(n9714), .B1(n14304), .B2(n14346), .ZN(
        n14358) );
  AOI22_X1 U15684 ( .A1(n14195), .A2(n16094), .B1(n14341), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n14196) );
  OAI21_X1 U15685 ( .B1(n14197), .B2(n14284), .A(n14196), .ZN(n14202) );
  OAI21_X1 U15686 ( .B1(n14200), .B2(n14199), .A(n14198), .ZN(n14359) );
  NOR2_X1 U15687 ( .A1(n14359), .A2(n14288), .ZN(n14201) );
  AOI211_X1 U15688 ( .C1(n16096), .C2(n14356), .A(n14202), .B(n14201), .ZN(
        n14203) );
  OAI21_X1 U15689 ( .B1(n14358), .B2(n14341), .A(n14203), .ZN(P3_U3207) );
  XNOR2_X1 U15690 ( .A(n14205), .B(n14204), .ZN(n14364) );
  AOI22_X1 U15691 ( .A1(n14206), .A2(n16094), .B1(n14341), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n14207) );
  OAI21_X1 U15692 ( .B1(n14208), .B2(n14284), .A(n14207), .ZN(n14215) );
  INV_X1 U15693 ( .A(n14209), .ZN(n14211) );
  AOI21_X1 U15694 ( .B1(n14211), .B2(n14210), .A(n16053), .ZN(n14213) );
  AOI22_X1 U15695 ( .A1(n14213), .A2(n14212), .B1(n14304), .B2(n14351), .ZN(
        n14363) );
  NOR2_X1 U15696 ( .A1(n14363), .A2(n14341), .ZN(n14214) );
  AOI211_X1 U15697 ( .C1(n16096), .C2(n14361), .A(n14215), .B(n14214), .ZN(
        n14216) );
  OAI21_X1 U15698 ( .B1(n14288), .B2(n14364), .A(n14216), .ZN(P3_U3208) );
  NOR2_X1 U15699 ( .A1(n14217), .A2(n14221), .ZN(n14218) );
  XOR2_X1 U15700 ( .A(n14221), .B(n14220), .Z(n14222) );
  NAND2_X1 U15701 ( .A1(n14222), .A2(n9714), .ZN(n14225) );
  AOI22_X1 U15702 ( .A1(n8346), .A2(n14304), .B1(n14384), .B2(n14223), .ZN(
        n14224) );
  OAI211_X1 U15703 ( .C1(n14256), .C2(n14366), .A(n14225), .B(n14224), .ZN(
        n14367) );
  AOI22_X1 U15704 ( .A1(n14226), .A2(n16094), .B1(n14341), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n14229) );
  NAND2_X1 U15705 ( .A1(n14227), .A2(n16096), .ZN(n14228) );
  OAI211_X1 U15706 ( .C1(n14366), .C2(n14263), .A(n14229), .B(n14228), .ZN(
        n14230) );
  AOI21_X1 U15707 ( .B1(n14367), .B2(n16100), .A(n14230), .ZN(n14231) );
  INV_X1 U15708 ( .A(n14231), .ZN(P3_U3209) );
  NAND2_X1 U15709 ( .A1(n14233), .A2(n14232), .ZN(n14234) );
  NAND2_X1 U15710 ( .A1(n14235), .A2(n14234), .ZN(n14374) );
  NAND2_X1 U15711 ( .A1(n14237), .A2(n14236), .ZN(n14238) );
  NAND2_X1 U15712 ( .A1(n14238), .A2(n9714), .ZN(n14239) );
  OR2_X1 U15713 ( .A1(n7524), .A2(n14239), .ZN(n14241) );
  NAND2_X1 U15714 ( .A1(n14360), .A2(n14304), .ZN(n14240) );
  NAND2_X1 U15715 ( .A1(n14241), .A2(n14240), .ZN(n14376) );
  NAND2_X1 U15716 ( .A1(n14376), .A2(n16100), .ZN(n14247) );
  AOI22_X1 U15717 ( .A1(n14341), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n16094), 
        .B2(n14242), .ZN(n14243) );
  OAI21_X1 U15718 ( .B1(n14244), .B2(n14284), .A(n14243), .ZN(n14245) );
  AOI21_X1 U15719 ( .B1(n14372), .B2(n16096), .A(n14245), .ZN(n14246) );
  OAI211_X1 U15720 ( .C1(n14374), .C2(n14288), .A(n14247), .B(n14246), .ZN(
        P3_U3210) );
  XNOR2_X1 U15721 ( .A(n14248), .B(n7950), .ZN(n14378) );
  OAI21_X1 U15722 ( .B1(n14251), .B2(n14250), .A(n14249), .ZN(n14254) );
  OAI22_X1 U15723 ( .A1(n14252), .A2(n16056), .B1(n14281), .B2(n16054), .ZN(
        n14253) );
  AOI21_X1 U15724 ( .B1(n14254), .B2(n9714), .A(n14253), .ZN(n14255) );
  OAI21_X1 U15725 ( .B1(n14256), .B2(n14378), .A(n14255), .ZN(n14379) );
  NAND2_X1 U15726 ( .A1(n14379), .A2(n16100), .ZN(n14262) );
  INV_X1 U15727 ( .A(n14257), .ZN(n14258) );
  OAI22_X1 U15728 ( .A1(n16100), .A2(n14259), .B1(n14258), .B2(n16059), .ZN(
        n14260) );
  AOI21_X1 U15729 ( .B1(n14377), .B2(n16096), .A(n14260), .ZN(n14261) );
  OAI211_X1 U15730 ( .C1(n14378), .C2(n14263), .A(n14262), .B(n14261), .ZN(
        P3_U3211) );
  XNOR2_X1 U15731 ( .A(n14264), .B(n14269), .ZN(n14265) );
  AOI22_X1 U15732 ( .A1(n14265), .A2(n9714), .B1(n14304), .B2(n14371), .ZN(
        n14387) );
  AOI22_X1 U15733 ( .A1(n14341), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n16094), 
        .B2(n14266), .ZN(n14267) );
  OAI21_X1 U15734 ( .B1(n14268), .B2(n14284), .A(n14267), .ZN(n14272) );
  XNOR2_X1 U15735 ( .A(n14270), .B(n14269), .ZN(n14388) );
  NOR2_X1 U15736 ( .A1(n14388), .A2(n14288), .ZN(n14271) );
  AOI211_X1 U15737 ( .C1(n16096), .C2(n14385), .A(n14272), .B(n14271), .ZN(
        n14273) );
  OAI21_X1 U15738 ( .B1(n14341), .B2(n14387), .A(n14273), .ZN(P3_U3212) );
  INV_X1 U15739 ( .A(n14292), .ZN(n14275) );
  OAI21_X1 U15740 ( .B1(n14275), .B2(n14274), .A(n7542), .ZN(n14277) );
  NAND2_X1 U15741 ( .A1(n14277), .A2(n14276), .ZN(n14392) );
  OAI211_X1 U15742 ( .C1(n14279), .C2(n7542), .A(n9714), .B(n14278), .ZN(
        n14280) );
  OAI21_X1 U15743 ( .B1(n14281), .B2(n16056), .A(n14280), .ZN(n14394) );
  NAND2_X1 U15744 ( .A1(n14394), .A2(n16100), .ZN(n14287) );
  AOI22_X1 U15745 ( .A1(n14341), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n16094), 
        .B2(n14282), .ZN(n14283) );
  OAI21_X1 U15746 ( .B1(n14390), .B2(n14284), .A(n14283), .ZN(n14285) );
  AOI21_X1 U15747 ( .B1(n14389), .B2(n16096), .A(n14285), .ZN(n14286) );
  OAI211_X1 U15748 ( .C1(n14288), .C2(n14392), .A(n14287), .B(n14286), .ZN(
        P3_U3213) );
  XOR2_X1 U15749 ( .A(n14289), .B(n14293), .Z(n14291) );
  AOI222_X1 U15750 ( .A1(n9714), .A2(n14291), .B1(n14290), .B2(n14384), .C1(
        n14383), .C2(n14304), .ZN(n14400) );
  OAI21_X1 U15751 ( .B1(n14294), .B2(n14293), .A(n14292), .ZN(n14398) );
  AOI22_X1 U15752 ( .A1(n14341), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n16094), 
        .B2(n14295), .ZN(n14296) );
  OAI21_X1 U15753 ( .B1(n14297), .B2(n14337), .A(n14296), .ZN(n14298) );
  AOI21_X1 U15754 ( .B1(n14398), .B2(n14339), .A(n14298), .ZN(n14299) );
  OAI21_X1 U15755 ( .B1(n14400), .B2(n14341), .A(n14299), .ZN(P3_U3214) );
  NOR2_X1 U15756 ( .A1(n8363), .A2(n14300), .ZN(n14303) );
  OAI21_X1 U15757 ( .B1(n14303), .B2(n14302), .A(n14301), .ZN(n14307) );
  AOI222_X1 U15758 ( .A1(n9714), .A2(n14307), .B1(n14306), .B2(n14384), .C1(
        n14305), .C2(n14304), .ZN(n14401) );
  OAI21_X1 U15759 ( .B1(n14309), .B2(n9576), .A(n14308), .ZN(n14403) );
  AOI22_X1 U15760 ( .A1(n14341), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n16094), 
        .B2(n14310), .ZN(n14311) );
  OAI21_X1 U15761 ( .B1(n14451), .B2(n14337), .A(n14311), .ZN(n14312) );
  AOI21_X1 U15762 ( .B1(n14403), .B2(n14339), .A(n14312), .ZN(n14313) );
  OAI21_X1 U15763 ( .B1(n14401), .B2(n14341), .A(n14313), .ZN(P3_U3215) );
  XNOR2_X1 U15764 ( .A(n14314), .B(n14319), .ZN(n14315) );
  OAI222_X1 U15765 ( .A1(n16054), .A2(n14317), .B1(n16056), .B2(n14316), .C1(
        n16053), .C2(n14315), .ZN(n14406) );
  INV_X1 U15766 ( .A(n14406), .ZN(n14325) );
  OAI21_X1 U15767 ( .B1(n14320), .B2(n14319), .A(n14318), .ZN(n14407) );
  AOI22_X1 U15768 ( .A1(n14341), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n16094), 
        .B2(n14321), .ZN(n14322) );
  OAI21_X1 U15769 ( .B1(n14455), .B2(n14337), .A(n14322), .ZN(n14323) );
  AOI21_X1 U15770 ( .B1(n14407), .B2(n14339), .A(n14323), .ZN(n14324) );
  OAI21_X1 U15771 ( .B1(n14325), .B2(n14341), .A(n14324), .ZN(P3_U3216) );
  INV_X1 U15772 ( .A(n14326), .ZN(n14327) );
  AOI21_X1 U15773 ( .B1(n14333), .B2(n14328), .A(n14327), .ZN(n14329) );
  OAI222_X1 U15774 ( .A1(n16054), .A2(n14331), .B1(n16056), .B2(n14330), .C1(
        n16053), .C2(n14329), .ZN(n14410) );
  INV_X1 U15775 ( .A(n14410), .ZN(n14342) );
  OAI21_X1 U15776 ( .B1(n14334), .B2(n14333), .A(n14332), .ZN(n14411) );
  AOI22_X1 U15777 ( .A1(n14341), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n16094), 
        .B2(n14335), .ZN(n14336) );
  OAI21_X1 U15778 ( .B1(n14459), .B2(n14337), .A(n14336), .ZN(n14338) );
  AOI21_X1 U15779 ( .B1(n14411), .B2(n14339), .A(n14338), .ZN(n14340) );
  OAI21_X1 U15780 ( .B1(n14342), .B2(n14341), .A(n14340), .ZN(P3_U3217) );
  NOR2_X1 U15781 ( .A1(n14423), .A2(n9764), .ZN(n14344) );
  AOI21_X1 U15782 ( .B1(P3_REG1_REG_31__SCAN_IN), .B2(n9764), .A(n14344), .ZN(
        n14343) );
  OAI21_X1 U15783 ( .B1(n14425), .B2(n14418), .A(n14343), .ZN(P3_U3490) );
  AOI21_X1 U15784 ( .B1(P3_REG1_REG_30__SCAN_IN), .B2(n9764), .A(n14344), .ZN(
        n14345) );
  OAI21_X1 U15785 ( .B1(n14428), .B2(n14418), .A(n14345), .ZN(P3_U3489) );
  AOI22_X1 U15786 ( .A1(n14347), .A2(n16102), .B1(n14384), .B2(n14346), .ZN(
        n14348) );
  OAI211_X1 U15787 ( .C1(n14391), .C2(n14350), .A(n14349), .B(n14348), .ZN(
        n14429) );
  MUX2_X1 U15788 ( .A(P3_REG1_REG_28__SCAN_IN), .B(n14429), .S(n16238), .Z(
        P3_U3487) );
  AOI22_X1 U15789 ( .A1(n14352), .A2(n16102), .B1(n14384), .B2(n14351), .ZN(
        n14353) );
  OAI211_X1 U15790 ( .C1(n14391), .C2(n14355), .A(n14354), .B(n14353), .ZN(
        n14430) );
  MUX2_X1 U15791 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n14430), .S(n16238), .Z(
        P3_U3486) );
  AOI22_X1 U15792 ( .A1(n14356), .A2(n16102), .B1(n14384), .B2(n8346), .ZN(
        n14357) );
  OAI211_X1 U15793 ( .C1(n14391), .C2(n14359), .A(n14358), .B(n14357), .ZN(
        n14431) );
  MUX2_X1 U15794 ( .A(P3_REG1_REG_26__SCAN_IN), .B(n14431), .S(n16238), .Z(
        P3_U3485) );
  AOI22_X1 U15795 ( .A1(n14361), .A2(n16102), .B1(n14384), .B2(n14360), .ZN(
        n14362) );
  OAI211_X1 U15796 ( .C1(n14391), .C2(n14364), .A(n14363), .B(n14362), .ZN(
        n14432) );
  MUX2_X1 U15797 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n14432), .S(n16238), .Z(
        P3_U3484) );
  INV_X1 U15798 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n14369) );
  INV_X1 U15799 ( .A(n14365), .ZN(n16236) );
  INV_X1 U15800 ( .A(n14366), .ZN(n14368) );
  AOI21_X1 U15801 ( .B1(n16236), .B2(n14368), .A(n14367), .ZN(n14433) );
  MUX2_X1 U15802 ( .A(n14369), .B(n14433), .S(n16238), .Z(n14370) );
  OAI21_X1 U15803 ( .B1(n14436), .B2(n14418), .A(n14370), .ZN(P3_U3483) );
  AOI22_X1 U15804 ( .A1(n14372), .A2(n16102), .B1(n14384), .B2(n14371), .ZN(
        n14373) );
  OAI21_X1 U15805 ( .B1(n14374), .B2(n14391), .A(n14373), .ZN(n14375) );
  MUX2_X1 U15806 ( .A(n14437), .B(P3_REG1_REG_23__SCAN_IN), .S(n9764), .Z(
        P3_U3482) );
  INV_X1 U15807 ( .A(n14377), .ZN(n14441) );
  INV_X1 U15808 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n14381) );
  INV_X1 U15809 ( .A(n14378), .ZN(n14380) );
  AOI21_X1 U15810 ( .B1(n16236), .B2(n14380), .A(n14379), .ZN(n14438) );
  MUX2_X1 U15811 ( .A(n14381), .B(n14438), .S(n16238), .Z(n14382) );
  OAI21_X1 U15812 ( .B1(n14441), .B2(n14418), .A(n14382), .ZN(P3_U3481) );
  AOI22_X1 U15813 ( .A1(n14385), .A2(n16102), .B1(n14384), .B2(n14383), .ZN(
        n14386) );
  OAI211_X1 U15814 ( .C1(n14391), .C2(n14388), .A(n14387), .B(n14386), .ZN(
        n14442) );
  MUX2_X1 U15815 ( .A(P3_REG1_REG_21__SCAN_IN), .B(n14442), .S(n16238), .Z(
        P3_U3480) );
  INV_X1 U15816 ( .A(n14389), .ZN(n14446) );
  OAI22_X1 U15817 ( .A1(n14392), .A2(n14391), .B1(n14390), .B2(n16054), .ZN(
        n14393) );
  NOR2_X1 U15818 ( .A1(n14394), .A2(n14393), .ZN(n14444) );
  INV_X1 U15819 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n14395) );
  MUX2_X1 U15820 ( .A(n14444), .B(n14395), .S(n9764), .Z(n14396) );
  OAI21_X1 U15821 ( .B1(n14446), .B2(n14418), .A(n14396), .ZN(P3_U3479) );
  AOI22_X1 U15822 ( .A1(n14398), .A2(n16103), .B1(n16102), .B2(n14397), .ZN(
        n14399) );
  NAND2_X1 U15823 ( .A1(n14400), .A2(n14399), .ZN(n14447) );
  MUX2_X1 U15824 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n14447), .S(n16238), .Z(
        P3_U3478) );
  INV_X1 U15825 ( .A(n14401), .ZN(n14402) );
  AOI21_X1 U15826 ( .B1(n16103), .B2(n14403), .A(n14402), .ZN(n14448) );
  MUX2_X1 U15827 ( .A(n14404), .B(n14448), .S(n16238), .Z(n14405) );
  OAI21_X1 U15828 ( .B1(n14451), .B2(n14418), .A(n14405), .ZN(P3_U3477) );
  AOI21_X1 U15829 ( .B1(n16103), .B2(n14407), .A(n14406), .ZN(n14452) );
  MUX2_X1 U15830 ( .A(n14408), .B(n14452), .S(n16238), .Z(n14409) );
  OAI21_X1 U15831 ( .B1(n14418), .B2(n14455), .A(n14409), .ZN(P3_U3476) );
  AOI21_X1 U15832 ( .B1(n16103), .B2(n14411), .A(n14410), .ZN(n14456) );
  MUX2_X1 U15833 ( .A(n14412), .B(n14456), .S(n16238), .Z(n14413) );
  OAI21_X1 U15834 ( .B1(n14459), .B2(n14418), .A(n14413), .ZN(P3_U3475) );
  AOI21_X1 U15835 ( .B1(n16103), .B2(n14415), .A(n14414), .ZN(n14460) );
  MUX2_X1 U15836 ( .A(n14416), .B(n14460), .S(n16238), .Z(n14417) );
  OAI21_X1 U15837 ( .B1(n14418), .B2(n14463), .A(n14417), .ZN(P3_U3474) );
  NAND2_X1 U15838 ( .A1(n14419), .A2(n16103), .ZN(n14420) );
  OAI211_X1 U15839 ( .C1(n16231), .C2(n14422), .A(n14421), .B(n14420), .ZN(
        n14465) );
  MUX2_X1 U15840 ( .A(P3_REG1_REG_14__SCAN_IN), .B(n14465), .S(n16238), .Z(
        P3_U3473) );
  NOR2_X1 U15841 ( .A1(n14423), .A2(n16239), .ZN(n14426) );
  AOI21_X1 U15842 ( .B1(P3_REG0_REG_31__SCAN_IN), .B2(n16239), .A(n14426), 
        .ZN(n14424) );
  OAI21_X1 U15843 ( .B1(n14425), .B2(n14464), .A(n14424), .ZN(P3_U3458) );
  AOI21_X1 U15844 ( .B1(n16239), .B2(P3_REG0_REG_30__SCAN_IN), .A(n14426), 
        .ZN(n14427) );
  OAI21_X1 U15845 ( .B1(n14428), .B2(n14464), .A(n14427), .ZN(P3_U3457) );
  MUX2_X1 U15846 ( .A(P3_REG0_REG_28__SCAN_IN), .B(n14429), .S(n16242), .Z(
        P3_U3455) );
  MUX2_X1 U15847 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n14430), .S(n16242), .Z(
        P3_U3454) );
  MUX2_X1 U15848 ( .A(P3_REG0_REG_26__SCAN_IN), .B(n14431), .S(n16242), .Z(
        P3_U3453) );
  MUX2_X1 U15849 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n14432), .S(n16242), .Z(
        P3_U3452) );
  INV_X1 U15850 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n14434) );
  MUX2_X1 U15851 ( .A(n14434), .B(n14433), .S(n16242), .Z(n14435) );
  OAI21_X1 U15852 ( .B1(n14436), .B2(n14464), .A(n14435), .ZN(P3_U3451) );
  MUX2_X1 U15853 ( .A(n14437), .B(P3_REG0_REG_23__SCAN_IN), .S(n16239), .Z(
        P3_U3450) );
  INV_X1 U15854 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n14439) );
  MUX2_X1 U15855 ( .A(n14439), .B(n14438), .S(n16242), .Z(n14440) );
  OAI21_X1 U15856 ( .B1(n14441), .B2(n14464), .A(n14440), .ZN(P3_U3449) );
  MUX2_X1 U15857 ( .A(P3_REG0_REG_21__SCAN_IN), .B(n14442), .S(n16242), .Z(
        P3_U3448) );
  INV_X1 U15858 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n14443) );
  MUX2_X1 U15859 ( .A(n14444), .B(n14443), .S(n16239), .Z(n14445) );
  OAI21_X1 U15860 ( .B1(n14446), .B2(n14464), .A(n14445), .ZN(P3_U3447) );
  MUX2_X1 U15861 ( .A(P3_REG0_REG_19__SCAN_IN), .B(n14447), .S(n16242), .Z(
        P3_U3446) );
  MUX2_X1 U15862 ( .A(n14449), .B(n14448), .S(n16242), .Z(n14450) );
  OAI21_X1 U15863 ( .B1(n14451), .B2(n14464), .A(n14450), .ZN(P3_U3444) );
  MUX2_X1 U15864 ( .A(n14453), .B(n14452), .S(n16242), .Z(n14454) );
  OAI21_X1 U15865 ( .B1(n14464), .B2(n14455), .A(n14454), .ZN(P3_U3441) );
  INV_X1 U15866 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n14457) );
  MUX2_X1 U15867 ( .A(n14457), .B(n14456), .S(n16242), .Z(n14458) );
  OAI21_X1 U15868 ( .B1(n14459), .B2(n14464), .A(n14458), .ZN(P3_U3438) );
  INV_X1 U15869 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n14461) );
  MUX2_X1 U15870 ( .A(n14461), .B(n14460), .S(n16242), .Z(n14462) );
  OAI21_X1 U15871 ( .B1(n14464), .B2(n14463), .A(n14462), .ZN(P3_U3435) );
  MUX2_X1 U15872 ( .A(P3_REG0_REG_14__SCAN_IN), .B(n14465), .S(n16242), .Z(
        P3_U3432) );
  MUX2_X1 U15873 ( .A(P3_D_REG_1__SCAN_IN), .B(n14466), .S(n14467), .Z(
        P3_U3377) );
  MUX2_X1 U15874 ( .A(P3_D_REG_0__SCAN_IN), .B(n14468), .S(n14467), .Z(
        P3_U3376) );
  NAND3_X1 U15875 ( .A1(n14470), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n14472) );
  OAI22_X1 U15876 ( .A1(n14469), .A2(n14472), .B1(n14471), .B2(n13926), .ZN(
        n14473) );
  AOI21_X1 U15877 ( .B1(n14475), .B2(n14474), .A(n14473), .ZN(n14476) );
  INV_X1 U15878 ( .A(n14476), .ZN(P3_U3264) );
  MUX2_X1 U15879 ( .A(n14477), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  INV_X1 U15880 ( .A(n14478), .ZN(n14480) );
  XNOR2_X1 U15881 ( .A(n15017), .B(n14487), .ZN(n14484) );
  NAND2_X1 U15882 ( .A1(n14675), .A2(n14552), .ZN(n14483) );
  NAND2_X1 U15883 ( .A1(n14484), .A2(n14483), .ZN(n14485) );
  OAI21_X1 U15884 ( .B1(n14484), .B2(n14483), .A(n14485), .ZN(n14585) );
  INV_X1 U15885 ( .A(n14485), .ZN(n14486) );
  XNOR2_X1 U15886 ( .A(n15011), .B(n14487), .ZN(n14489) );
  NAND2_X1 U15887 ( .A1(n14674), .A2(n11126), .ZN(n14488) );
  NAND2_X1 U15888 ( .A1(n14489), .A2(n14488), .ZN(n14490) );
  OAI21_X1 U15889 ( .B1(n14489), .B2(n14488), .A(n14490), .ZN(n14594) );
  INV_X1 U15890 ( .A(n14490), .ZN(n14491) );
  NAND2_X1 U15891 ( .A1(n14673), .A2(n11126), .ZN(n14492) );
  XNOR2_X1 U15892 ( .A(n14493), .B(n14492), .ZN(n14635) );
  INV_X1 U15893 ( .A(n14492), .ZN(n14494) );
  NAND2_X1 U15894 ( .A1(n14884), .A2(n11126), .ZN(n14496) );
  INV_X1 U15895 ( .A(n14495), .ZN(n14497) );
  XNOR2_X1 U15896 ( .A(n14993), .B(n14553), .ZN(n14499) );
  NAND2_X1 U15897 ( .A1(n14857), .A2(n11126), .ZN(n14498) );
  XNOR2_X1 U15898 ( .A(n14499), .B(n14498), .ZN(n14610) );
  INV_X1 U15899 ( .A(n14498), .ZN(n14500) );
  NAND2_X1 U15900 ( .A1(n14886), .A2(n11126), .ZN(n14502) );
  XNOR2_X1 U15901 ( .A(n14987), .B(n14553), .ZN(n14501) );
  XOR2_X1 U15902 ( .A(n14502), .B(n14501), .Z(n14568) );
  INV_X1 U15903 ( .A(n14501), .ZN(n14503) );
  XNOR2_X1 U15904 ( .A(n14981), .B(n14525), .ZN(n14505) );
  XNOR2_X1 U15905 ( .A(n14504), .B(n14505), .ZN(n14618) );
  NAND2_X1 U15906 ( .A1(n14858), .A2(n11126), .ZN(n14617) );
  INV_X1 U15907 ( .A(n14504), .ZN(n14507) );
  INV_X1 U15908 ( .A(n14505), .ZN(n14506) );
  OAI22_X1 U15909 ( .A1(n14618), .A2(n14617), .B1(n14507), .B2(n14506), .ZN(
        n14508) );
  XNOR2_X1 U15910 ( .A(n14975), .B(n14525), .ZN(n14509) );
  XNOR2_X1 U15911 ( .A(n14508), .B(n14509), .ZN(n14532) );
  NAND2_X1 U15912 ( .A1(n14837), .A2(n11126), .ZN(n14533) );
  INV_X1 U15913 ( .A(n14508), .ZN(n14511) );
  INV_X1 U15914 ( .A(n14509), .ZN(n14510) );
  XNOR2_X1 U15915 ( .A(n14969), .B(n14553), .ZN(n14512) );
  NAND2_X1 U15916 ( .A1(n14819), .A2(n14552), .ZN(n14513) );
  XNOR2_X1 U15917 ( .A(n14512), .B(n14513), .ZN(n14603) );
  NAND2_X1 U15918 ( .A1(n14604), .A2(n14603), .ZN(n14516) );
  INV_X1 U15919 ( .A(n14513), .ZN(n14514) );
  NAND2_X1 U15920 ( .A1(n14512), .A2(n14514), .ZN(n14515) );
  XNOR2_X1 U15921 ( .A(n14964), .B(n14525), .ZN(n14517) );
  NAND2_X1 U15922 ( .A1(n14811), .A2(n11126), .ZN(n14518) );
  XNOR2_X1 U15923 ( .A(n14517), .B(n14518), .ZN(n14576) );
  INV_X1 U15924 ( .A(n14517), .ZN(n14519) );
  NOR2_X1 U15925 ( .A1(n14519), .A2(n14518), .ZN(n14520) );
  AND2_X1 U15926 ( .A1(n14795), .A2(n14552), .ZN(n14522) );
  XNOR2_X1 U15927 ( .A(n14959), .B(n14525), .ZN(n14521) );
  NOR2_X1 U15928 ( .A1(n14521), .A2(n14522), .ZN(n14523) );
  AOI21_X1 U15929 ( .B1(n14522), .B2(n14521), .A(n14523), .ZN(n14657) );
  NAND2_X1 U15930 ( .A1(n14656), .A2(n14657), .ZN(n14655) );
  INV_X1 U15931 ( .A(n14523), .ZN(n14524) );
  NAND2_X1 U15932 ( .A1(n14655), .A2(n14524), .ZN(n14551) );
  NAND2_X1 U15933 ( .A1(n14774), .A2(n11126), .ZN(n14548) );
  XNOR2_X1 U15934 ( .A(n14954), .B(n14525), .ZN(n14547) );
  XOR2_X1 U15935 ( .A(n14548), .B(n14547), .Z(n14550) );
  XNOR2_X1 U15936 ( .A(n14551), .B(n14550), .ZN(n14531) );
  NOR2_X1 U15937 ( .A1(n14751), .A2(n14661), .ZN(n14528) );
  OAI22_X1 U15938 ( .A1(n14760), .A2(n14638), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14526), .ZN(n14527) );
  AOI211_X1 U15939 ( .C1(n14672), .C2(n14627), .A(n14528), .B(n14527), .ZN(
        n14530) );
  NAND2_X1 U15940 ( .A1(n14954), .A2(n14651), .ZN(n14529) );
  OAI211_X1 U15941 ( .C1(n14531), .C2(n14642), .A(n14530), .B(n14529), .ZN(
        P2_U3186) );
  XNOR2_X1 U15942 ( .A(n14532), .B(n14533), .ZN(n14540) );
  OAI22_X1 U15943 ( .A1(n14535), .A2(n14663), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14534), .ZN(n14538) );
  INV_X1 U15944 ( .A(n14826), .ZN(n14536) );
  OAI22_X1 U15945 ( .A1(n14571), .A2(n14661), .B1(n14536), .B2(n14638), .ZN(
        n14537) );
  AOI211_X1 U15946 ( .C1(n14975), .C2(n14651), .A(n14538), .B(n14537), .ZN(
        n14539) );
  OAI21_X1 U15947 ( .B1(n14540), .B2(n14642), .A(n14539), .ZN(P2_U3188) );
  XNOR2_X1 U15948 ( .A(n14542), .B(n14541), .ZN(n14546) );
  AOI22_X1 U15949 ( .A1(n14648), .A2(n14673), .B1(n14667), .B2(n14904), .ZN(
        n14543) );
  NAND2_X1 U15950 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3088), .ZN(n15713)
         );
  OAI211_X1 U15951 ( .C1(n14895), .C2(n14663), .A(n14543), .B(n15713), .ZN(
        n14544) );
  AOI21_X1 U15952 ( .B1(n15001), .B2(n14651), .A(n14544), .ZN(n14545) );
  OAI21_X1 U15953 ( .B1(n14546), .B2(n14642), .A(n14545), .ZN(P2_U3191) );
  INV_X1 U15954 ( .A(n14547), .ZN(n14549) );
  MUX2_X1 U15955 ( .A(n14949), .B(n14737), .S(n14552), .Z(n14554) );
  XNOR2_X1 U15956 ( .A(n14554), .B(n14553), .ZN(n14555) );
  XNOR2_X1 U15957 ( .A(n14556), .B(n14555), .ZN(n14561) );
  AOI22_X1 U15958 ( .A1(n14743), .A2(n14667), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14557) );
  OAI21_X1 U15959 ( .B1(n14664), .B2(n14661), .A(n14557), .ZN(n14559) );
  NOR2_X1 U15960 ( .A1(n7418), .A2(n14670), .ZN(n14558) );
  AOI211_X1 U15961 ( .C1(n14627), .C2(n14740), .A(n14559), .B(n14558), .ZN(
        n14560) );
  OAI21_X1 U15962 ( .B1(n14561), .B2(n14642), .A(n14560), .ZN(P2_U3192) );
  AOI22_X1 U15963 ( .A1(n14651), .A2(n7432), .B1(n14625), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n14567) );
  AOI22_X1 U15964 ( .A1(n14648), .A2(n13669), .B1(n14627), .B2(n7423), .ZN(
        n14566) );
  NOR2_X1 U15965 ( .A1(n14563), .A2(n14562), .ZN(n14564) );
  OAI21_X1 U15966 ( .B1(n14630), .B2(n14564), .A(n14658), .ZN(n14565) );
  NAND3_X1 U15967 ( .A1(n14567), .A2(n14566), .A3(n14565), .ZN(P2_U3194) );
  XNOR2_X1 U15968 ( .A(n14569), .B(n14568), .ZN(n14575) );
  OAI22_X1 U15969 ( .A1(n14571), .A2(n14663), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14570), .ZN(n14573) );
  OAI22_X1 U15970 ( .A1(n14638), .A2(n14865), .B1(n14895), .B2(n14661), .ZN(
        n14572) );
  AOI211_X1 U15971 ( .C1(n14987), .C2(n14651), .A(n14573), .B(n14572), .ZN(
        n14574) );
  OAI21_X1 U15972 ( .B1(n14575), .B2(n14642), .A(n14574), .ZN(P2_U3195) );
  XNOR2_X1 U15973 ( .A(n14577), .B(n14576), .ZN(n14582) );
  NAND2_X1 U15974 ( .A1(n14795), .A2(n14627), .ZN(n14579) );
  AOI22_X1 U15975 ( .A1(n14819), .A2(n14648), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14578) );
  OAI211_X1 U15976 ( .C1(n14638), .C2(n14788), .A(n14579), .B(n14578), .ZN(
        n14580) );
  AOI21_X1 U15977 ( .B1(n14964), .B2(n14651), .A(n14580), .ZN(n14581) );
  OAI21_X1 U15978 ( .B1(n14582), .B2(n14642), .A(n14581), .ZN(P2_U3197) );
  AOI21_X1 U15979 ( .B1(n14585), .B2(n14584), .A(n14583), .ZN(n14592) );
  OAI22_X1 U15980 ( .A1(n14663), .A2(n14915), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14586), .ZN(n14590) );
  OAI22_X1 U15981 ( .A1(n14638), .A2(n14588), .B1(n14587), .B2(n14661), .ZN(
        n14589) );
  AOI211_X1 U15982 ( .C1(n15017), .C2(n14651), .A(n14590), .B(n14589), .ZN(
        n14591) );
  OAI21_X1 U15983 ( .B1(n14592), .B2(n14642), .A(n14591), .ZN(P2_U3198) );
  AOI21_X1 U15984 ( .B1(n14595), .B2(n14594), .A(n14593), .ZN(n14602) );
  OAI21_X1 U15985 ( .B1(n14663), .B2(n14894), .A(n14596), .ZN(n14600) );
  OAI22_X1 U15986 ( .A1(n14638), .A2(n14598), .B1(n14597), .B2(n14661), .ZN(
        n14599) );
  AOI211_X1 U15987 ( .C1(n15011), .C2(n14651), .A(n14600), .B(n14599), .ZN(
        n14601) );
  OAI21_X1 U15988 ( .B1(n14602), .B2(n14642), .A(n14601), .ZN(P2_U3200) );
  XNOR2_X1 U15989 ( .A(n14604), .B(n14603), .ZN(n14609) );
  OAI22_X1 U15990 ( .A1(n14620), .A2(n14661), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14605), .ZN(n14607) );
  OAI22_X1 U15991 ( .A1(n14662), .A2(n14663), .B1(n14638), .B2(n14803), .ZN(
        n14606) );
  AOI211_X1 U15992 ( .C1(n14969), .C2(n14651), .A(n14607), .B(n14606), .ZN(
        n14608) );
  OAI21_X1 U15993 ( .B1(n14609), .B2(n14642), .A(n14608), .ZN(P2_U3201) );
  XNOR2_X1 U15994 ( .A(n14611), .B(n14610), .ZN(n14616) );
  OAI22_X1 U15995 ( .A1(n14663), .A2(n8168), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13421), .ZN(n14614) );
  INV_X1 U15996 ( .A(n14877), .ZN(n14612) );
  OAI22_X1 U15997 ( .A1(n14638), .A2(n14612), .B1(n14917), .B2(n14661), .ZN(
        n14613) );
  AOI211_X1 U15998 ( .C1(n14993), .C2(n14651), .A(n14614), .B(n14613), .ZN(
        n14615) );
  OAI21_X1 U15999 ( .B1(n14616), .B2(n14642), .A(n14615), .ZN(P2_U3205) );
  XNOR2_X1 U16000 ( .A(n14618), .B(n14617), .ZN(n14624) );
  OAI22_X1 U16001 ( .A1(n14620), .A2(n14663), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14619), .ZN(n14622) );
  OAI22_X1 U16002 ( .A1(n14638), .A2(n14841), .B1(n8168), .B2(n14661), .ZN(
        n14621) );
  AOI211_X1 U16003 ( .C1(n14981), .C2(n14651), .A(n14622), .B(n14621), .ZN(
        n14623) );
  OAI21_X1 U16004 ( .B1(n14624), .B2(n14642), .A(n14623), .ZN(P2_U3207) );
  AOI22_X1 U16005 ( .A1(n14651), .A2(n14626), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n14625), .ZN(n14634) );
  AOI22_X1 U16006 ( .A1(n14648), .A2(n7580), .B1(n14627), .B2(n14689), .ZN(
        n14633) );
  NOR3_X1 U16007 ( .A1(n14630), .A2(n14629), .A3(n14628), .ZN(n14631) );
  OAI21_X1 U16008 ( .B1(n7570), .B2(n14631), .A(n14658), .ZN(n14632) );
  NAND3_X1 U16009 ( .A1(n14634), .A2(n14633), .A3(n14632), .ZN(P2_U3209) );
  XNOR2_X1 U16010 ( .A(n14636), .B(n14635), .ZN(n14643) );
  OAI22_X1 U16011 ( .A1(n14663), .A2(n14917), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14637), .ZN(n14640) );
  OAI22_X1 U16012 ( .A1(n14638), .A2(n14928), .B1(n14915), .B2(n14661), .ZN(
        n14639) );
  AOI211_X1 U16013 ( .C1(n15005), .C2(n14651), .A(n14640), .B(n14639), .ZN(
        n14641) );
  OAI21_X1 U16014 ( .B1(n14643), .B2(n14642), .A(n14641), .ZN(P2_U3210) );
  OAI211_X1 U16015 ( .C1(n14646), .C2(n14645), .A(n14644), .B(n14658), .ZN(
        n14654) );
  AOI22_X1 U16016 ( .A1(n14648), .A2(n14687), .B1(n14667), .B2(n14647), .ZN(
        n14653) );
  NAND2_X1 U16017 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n15665) );
  OAI21_X1 U16018 ( .B1(n14663), .B2(n14649), .A(n15665), .ZN(n14650) );
  AOI21_X1 U16019 ( .B1(n16122), .B2(n14651), .A(n14650), .ZN(n14652) );
  NAND3_X1 U16020 ( .A1(n14654), .A2(n14653), .A3(n14652), .ZN(P2_U3211) );
  INV_X1 U16021 ( .A(n14959), .ZN(n14780) );
  OAI21_X1 U16022 ( .B1(n14657), .B2(n14656), .A(n14655), .ZN(n14659) );
  NAND2_X1 U16023 ( .A1(n14659), .A2(n14658), .ZN(n14669) );
  OAI22_X1 U16024 ( .A1(n14662), .A2(n14661), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14660), .ZN(n14666) );
  NOR2_X1 U16025 ( .A1(n14664), .A2(n14663), .ZN(n14665) );
  AOI211_X1 U16026 ( .C1(n14667), .C2(n14777), .A(n14666), .B(n14665), .ZN(
        n14668) );
  OAI211_X1 U16027 ( .C1(n14780), .C2(n14670), .A(n14669), .B(n14668), .ZN(
        P2_U3212) );
  MUX2_X1 U16028 ( .A(n14724), .B(P2_DATAO_REG_31__SCAN_IN), .S(n14683), .Z(
        P2_U3562) );
  MUX2_X1 U16029 ( .A(n14671), .B(P2_DATAO_REG_30__SCAN_IN), .S(n14683), .Z(
        P2_U3561) );
  MUX2_X1 U16030 ( .A(n14740), .B(P2_DATAO_REG_29__SCAN_IN), .S(n14683), .Z(
        P2_U3560) );
  MUX2_X1 U16031 ( .A(n14672), .B(P2_DATAO_REG_28__SCAN_IN), .S(n14683), .Z(
        P2_U3559) );
  MUX2_X1 U16032 ( .A(n14774), .B(P2_DATAO_REG_27__SCAN_IN), .S(n14683), .Z(
        P2_U3558) );
  MUX2_X1 U16033 ( .A(n14795), .B(P2_DATAO_REG_26__SCAN_IN), .S(n14683), .Z(
        P2_U3557) );
  MUX2_X1 U16034 ( .A(n14811), .B(P2_DATAO_REG_25__SCAN_IN), .S(n14683), .Z(
        P2_U3556) );
  MUX2_X1 U16035 ( .A(n14819), .B(P2_DATAO_REG_24__SCAN_IN), .S(n14683), .Z(
        P2_U3555) );
  MUX2_X1 U16036 ( .A(n14837), .B(P2_DATAO_REG_23__SCAN_IN), .S(n14683), .Z(
        P2_U3554) );
  MUX2_X1 U16037 ( .A(n14858), .B(P2_DATAO_REG_22__SCAN_IN), .S(n14683), .Z(
        P2_U3553) );
  MUX2_X1 U16038 ( .A(n14886), .B(P2_DATAO_REG_21__SCAN_IN), .S(n14683), .Z(
        P2_U3552) );
  MUX2_X1 U16039 ( .A(n14857), .B(P2_DATAO_REG_20__SCAN_IN), .S(n14683), .Z(
        P2_U3551) );
  MUX2_X1 U16040 ( .A(n14884), .B(P2_DATAO_REG_19__SCAN_IN), .S(n14683), .Z(
        P2_U3550) );
  MUX2_X1 U16041 ( .A(n14673), .B(P2_DATAO_REG_18__SCAN_IN), .S(n14683), .Z(
        P2_U3549) );
  MUX2_X1 U16042 ( .A(n14674), .B(P2_DATAO_REG_17__SCAN_IN), .S(n14683), .Z(
        P2_U3548) );
  MUX2_X1 U16043 ( .A(n14675), .B(P2_DATAO_REG_16__SCAN_IN), .S(n14683), .Z(
        P2_U3547) );
  MUX2_X1 U16044 ( .A(n14676), .B(P2_DATAO_REG_15__SCAN_IN), .S(n14683), .Z(
        P2_U3546) );
  MUX2_X1 U16045 ( .A(n14677), .B(P2_DATAO_REG_14__SCAN_IN), .S(n14683), .Z(
        P2_U3545) );
  MUX2_X1 U16046 ( .A(n14678), .B(P2_DATAO_REG_13__SCAN_IN), .S(n14683), .Z(
        P2_U3544) );
  MUX2_X1 U16047 ( .A(n14679), .B(P2_DATAO_REG_12__SCAN_IN), .S(n14683), .Z(
        P2_U3543) );
  MUX2_X1 U16048 ( .A(n14680), .B(P2_DATAO_REG_11__SCAN_IN), .S(n14683), .Z(
        P2_U3542) );
  MUX2_X1 U16049 ( .A(n14681), .B(P2_DATAO_REG_10__SCAN_IN), .S(n14683), .Z(
        P2_U3541) );
  MUX2_X1 U16050 ( .A(n14682), .B(P2_DATAO_REG_9__SCAN_IN), .S(n14683), .Z(
        P2_U3540) );
  MUX2_X1 U16051 ( .A(n14684), .B(P2_DATAO_REG_8__SCAN_IN), .S(n14683), .Z(
        P2_U3539) );
  MUX2_X1 U16052 ( .A(n14685), .B(P2_DATAO_REG_7__SCAN_IN), .S(n14683), .Z(
        P2_U3538) );
  MUX2_X1 U16053 ( .A(n14686), .B(P2_DATAO_REG_6__SCAN_IN), .S(n14683), .Z(
        P2_U3537) );
  MUX2_X1 U16054 ( .A(n14687), .B(P2_DATAO_REG_5__SCAN_IN), .S(n14683), .Z(
        P2_U3536) );
  MUX2_X1 U16055 ( .A(n14688), .B(P2_DATAO_REG_4__SCAN_IN), .S(n14683), .Z(
        P2_U3535) );
  MUX2_X1 U16056 ( .A(n14689), .B(P2_DATAO_REG_3__SCAN_IN), .S(n14683), .Z(
        P2_U3534) );
  MUX2_X1 U16057 ( .A(n7423), .B(P2_DATAO_REG_2__SCAN_IN), .S(n14683), .Z(
        P2_U3533) );
  MUX2_X1 U16058 ( .A(n7580), .B(P2_DATAO_REG_1__SCAN_IN), .S(n14683), .Z(
        P2_U3532) );
  MUX2_X1 U16059 ( .A(n13669), .B(P2_DATAO_REG_0__SCAN_IN), .S(n14683), .Z(
        P2_U3531) );
  INV_X1 U16060 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n14692) );
  OAI22_X1 U16061 ( .A1(n15724), .A2(n14698), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14692), .ZN(n14693) );
  AOI21_X1 U16062 ( .B1(n15683), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n14693), .ZN(
        n14705) );
  MUX2_X1 U16063 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n10547), .S(n14698), .Z(
        n14696) );
  INV_X1 U16064 ( .A(n14694), .ZN(n14695) );
  NAND2_X1 U16065 ( .A1(n14696), .A2(n14695), .ZN(n14697) );
  OAI211_X1 U16066 ( .C1(n15657), .C2(n14697), .A(n15743), .B(n14711), .ZN(
        n14704) );
  MUX2_X1 U16067 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n14699), .S(n14698), .Z(
        n14700) );
  NAND3_X1 U16068 ( .A1(n15654), .A2(n14701), .A3(n14700), .ZN(n14702) );
  NAND3_X1 U16069 ( .A1(n15718), .A2(n14717), .A3(n14702), .ZN(n14703) );
  NAND3_X1 U16070 ( .A1(n14705), .A2(n14704), .A3(n14703), .ZN(P2_U3216) );
  OAI22_X1 U16071 ( .A1(n15724), .A2(n14714), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14706), .ZN(n14707) );
  AOI21_X1 U16072 ( .B1(n15683), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n14707), .ZN(
        n14722) );
  INV_X1 U16073 ( .A(n14708), .ZN(n14713) );
  NAND3_X1 U16074 ( .A1(n14711), .A2(n14710), .A3(n14709), .ZN(n14712) );
  NAND3_X1 U16075 ( .A1(n15743), .A2(n14713), .A3(n14712), .ZN(n14721) );
  MUX2_X1 U16076 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10559), .S(n14714), .Z(
        n14715) );
  NAND3_X1 U16077 ( .A1(n14717), .A2(n14716), .A3(n14715), .ZN(n14718) );
  NAND3_X1 U16078 ( .A1(n15718), .A2(n14719), .A3(n14718), .ZN(n14720) );
  NAND3_X1 U16079 ( .A1(n14722), .A2(n14721), .A3(n14720), .ZN(P2_U3217) );
  NAND2_X1 U16080 ( .A1(n14729), .A2(n14942), .ZN(n14728) );
  NAND2_X1 U16081 ( .A1(n14724), .A2(n14723), .ZN(n14940) );
  NOR2_X1 U16082 ( .A1(n14938), .A2(n14940), .ZN(n14731) );
  NOR2_X1 U16083 ( .A1(n7966), .A2(n14932), .ZN(n14726) );
  AOI211_X1 U16084 ( .C1(P2_REG2_REG_31__SCAN_IN), .C2(n14938), .A(n14731), 
        .B(n14726), .ZN(n14727) );
  OAI21_X1 U16085 ( .B1(n14733), .B2(n14939), .A(n14727), .ZN(P2_U3234) );
  OAI211_X1 U16086 ( .C1(n14729), .C2(n14942), .A(n14728), .B(n15027), .ZN(
        n14941) );
  NOR2_X1 U16087 ( .A1(n14942), .A2(n14932), .ZN(n14730) );
  AOI211_X1 U16088 ( .C1(n14938), .C2(P2_REG2_REG_30__SCAN_IN), .A(n14731), 
        .B(n14730), .ZN(n14732) );
  OAI21_X1 U16089 ( .B1(n14733), .B2(n14941), .A(n14732), .ZN(P2_U3235) );
  AND2_X2 U16090 ( .A1(n14736), .A2(n14735), .ZN(n14951) );
  INV_X1 U16091 ( .A(n14951), .ZN(n14749) );
  AOI22_X1 U16092 ( .A1(n14740), .A2(n14885), .B1(n14883), .B2(n14774), .ZN(
        n14741) );
  INV_X1 U16093 ( .A(n14953), .ZN(n14746) );
  OAI211_X1 U16094 ( .C1(n14759), .C2(n7418), .A(n15027), .B(n7467), .ZN(
        n14948) );
  INV_X1 U16095 ( .A(n14743), .ZN(n14744) );
  OAI22_X1 U16096 ( .A1(n14948), .A2(n7415), .B1(n14840), .B2(n14744), .ZN(
        n14745) );
  OAI21_X1 U16097 ( .B1(n14746), .B2(n14745), .A(n14843), .ZN(n14748) );
  AOI22_X1 U16098 ( .A1(n14949), .A2(n14849), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n14938), .ZN(n14747) );
  XOR2_X1 U16099 ( .A(n14750), .B(n14753), .Z(n14764) );
  OAI22_X1 U16100 ( .A1(n14752), .A2(n14916), .B1(n14751), .B2(n14914), .ZN(
        n14758) );
  NAND3_X1 U16101 ( .A1(n14773), .A2(n7820), .A3(n14754), .ZN(n14755) );
  AOI21_X1 U16102 ( .B1(n14756), .B2(n14755), .A(n14821), .ZN(n14757) );
  AOI21_X1 U16103 ( .B1(n14954), .B2(n7511), .A(n14759), .ZN(n14955) );
  INV_X1 U16104 ( .A(n14954), .ZN(n14763) );
  INV_X1 U16105 ( .A(n14760), .ZN(n14761) );
  AOI22_X1 U16106 ( .A1(n14761), .A2(n14929), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n14938), .ZN(n14762) );
  OAI21_X1 U16107 ( .B1(n14763), .B2(n14932), .A(n14762), .ZN(n14766) );
  INV_X1 U16108 ( .A(n14764), .ZN(n14958) );
  NOR2_X1 U16109 ( .A1(n14958), .A2(n14933), .ZN(n14765) );
  AOI211_X1 U16110 ( .C1(n14955), .C2(n14936), .A(n14766), .B(n14765), .ZN(
        n14767) );
  OAI21_X1 U16111 ( .B1(n14957), .B2(n14938), .A(n14767), .ZN(P2_U3238) );
  XNOR2_X1 U16112 ( .A(n14769), .B(n14768), .ZN(n14963) );
  NAND3_X1 U16113 ( .A1(n14792), .A2(n14771), .A3(n14770), .ZN(n14772) );
  NAND2_X1 U16114 ( .A1(n14773), .A2(n14772), .ZN(n14775) );
  AOI222_X1 U16115 ( .A1(n14924), .A2(n14775), .B1(n14774), .B2(n14885), .C1(
        n14811), .C2(n14883), .ZN(n14962) );
  INV_X1 U16116 ( .A(n14962), .ZN(n14782) );
  NAND2_X1 U16117 ( .A1(n14785), .A2(n14959), .ZN(n14776) );
  AND2_X1 U16118 ( .A1(n7511), .A2(n14776), .ZN(n14960) );
  NAND2_X1 U16119 ( .A1(n14960), .A2(n14936), .ZN(n14779) );
  AOI22_X1 U16120 ( .A1(n14777), .A2(n14929), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n14938), .ZN(n14778) );
  OAI211_X1 U16121 ( .C1(n14780), .C2(n14932), .A(n14779), .B(n14778), .ZN(
        n14781) );
  AOI21_X1 U16122 ( .B1(n14782), .B2(n14843), .A(n14781), .ZN(n14783) );
  OAI21_X1 U16123 ( .B1(n14891), .B2(n14963), .A(n14783), .ZN(P2_U3239) );
  XNOR2_X1 U16124 ( .A(n14784), .B(n14794), .ZN(n14968) );
  INV_X1 U16125 ( .A(n14802), .ZN(n14787) );
  INV_X1 U16126 ( .A(n14785), .ZN(n14786) );
  AOI21_X1 U16127 ( .B1(n14964), .B2(n14787), .A(n14786), .ZN(n14965) );
  INV_X1 U16128 ( .A(n14788), .ZN(n14789) );
  AOI22_X1 U16129 ( .A1(n14789), .A2(n14929), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n14938), .ZN(n14790) );
  OAI21_X1 U16130 ( .B1(n14791), .B2(n14932), .A(n14790), .ZN(n14798) );
  OAI21_X1 U16131 ( .B1(n14794), .B2(n14793), .A(n14792), .ZN(n14796) );
  AOI211_X1 U16132 ( .C1(n14965), .C2(n14936), .A(n14798), .B(n14797), .ZN(
        n14799) );
  OAI21_X1 U16133 ( .B1(n14968), .B2(n14891), .A(n14799), .ZN(P2_U3240) );
  XOR2_X1 U16134 ( .A(n14800), .B(n7827), .Z(n14973) );
  AND2_X1 U16135 ( .A1(n14824), .A2(n14969), .ZN(n14801) );
  NOR2_X1 U16136 ( .A1(n14802), .A2(n14801), .ZN(n14970) );
  INV_X1 U16137 ( .A(n14969), .ZN(n14806) );
  INV_X1 U16138 ( .A(n14803), .ZN(n14804) );
  AOI22_X1 U16139 ( .A1(n14804), .A2(n14929), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n14938), .ZN(n14805) );
  OAI21_X1 U16140 ( .B1(n14806), .B2(n14932), .A(n14805), .ZN(n14814) );
  INV_X1 U16141 ( .A(n14807), .ZN(n14810) );
  INV_X1 U16142 ( .A(n7825), .ZN(n14809) );
  OAI21_X1 U16143 ( .B1(n14810), .B2(n14809), .A(n14808), .ZN(n14812) );
  AOI222_X1 U16144 ( .A1(n14924), .A2(n14812), .B1(n14811), .B2(n14885), .C1(
        n14837), .C2(n14883), .ZN(n14972) );
  NOR2_X1 U16145 ( .A1(n14972), .A2(n14938), .ZN(n14813) );
  AOI211_X1 U16146 ( .C1(n14970), .C2(n14936), .A(n14814), .B(n14813), .ZN(
        n14815) );
  OAI21_X1 U16147 ( .B1(n14973), .B2(n14891), .A(n14815), .ZN(P2_U3241) );
  XNOR2_X1 U16148 ( .A(n14816), .B(n14818), .ZN(n14829) );
  XNOR2_X1 U16149 ( .A(n14817), .B(n14818), .ZN(n14822) );
  AOI22_X1 U16150 ( .A1(n14819), .A2(n14885), .B1(n14883), .B2(n14858), .ZN(
        n14820) );
  OAI21_X1 U16151 ( .B1(n14822), .B2(n14821), .A(n14820), .ZN(n14823) );
  AOI21_X1 U16152 ( .B1(n14902), .B2(n14829), .A(n14823), .ZN(n14976) );
  INV_X1 U16153 ( .A(n14824), .ZN(n14825) );
  AOI211_X1 U16154 ( .C1(n14975), .C2(n14845), .A(n10363), .B(n14825), .ZN(
        n14974) );
  INV_X1 U16155 ( .A(n14975), .ZN(n14828) );
  AOI22_X1 U16156 ( .A1(n14938), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n14826), 
        .B2(n14929), .ZN(n14827) );
  OAI21_X1 U16157 ( .B1(n14828), .B2(n14932), .A(n14827), .ZN(n14831) );
  INV_X1 U16158 ( .A(n14829), .ZN(n14978) );
  NOR2_X1 U16159 ( .A1(n14978), .A2(n14933), .ZN(n14830) );
  AOI211_X1 U16160 ( .C1(n14974), .C2(n14832), .A(n14831), .B(n14830), .ZN(
        n14833) );
  OAI21_X1 U16161 ( .B1(n14938), .B2(n14976), .A(n14833), .ZN(P2_U3242) );
  INV_X1 U16162 ( .A(n14834), .ZN(n14835) );
  XNOR2_X1 U16163 ( .A(n14851), .B(n14835), .ZN(n14836) );
  NAND2_X1 U16164 ( .A1(n14836), .A2(n14924), .ZN(n14839) );
  AOI22_X1 U16165 ( .A1(n14837), .A2(n14885), .B1(n14883), .B2(n14886), .ZN(
        n14838) );
  NAND2_X1 U16166 ( .A1(n14839), .A2(n14838), .ZN(n14985) );
  INV_X1 U16167 ( .A(n14985), .ZN(n14854) );
  INV_X1 U16168 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n14842) );
  OAI22_X1 U16169 ( .A1(n14843), .A2(n14842), .B1(n14841), .B2(n14840), .ZN(
        n14848) );
  NAND2_X1 U16170 ( .A1(n14981), .A2(n14864), .ZN(n14844) );
  NAND2_X1 U16171 ( .A1(n14845), .A2(n14844), .ZN(n14982) );
  NOR2_X1 U16172 ( .A1(n14982), .A2(n14846), .ZN(n14847) );
  AOI211_X1 U16173 ( .C1(n14849), .C2(n14981), .A(n14848), .B(n14847), .ZN(
        n14853) );
  NAND2_X1 U16174 ( .A1(n14851), .A2(n14850), .ZN(n14979) );
  NAND3_X1 U16175 ( .A1(n14980), .A2(n14979), .A3(n14870), .ZN(n14852) );
  OAI211_X1 U16176 ( .C1(n14854), .C2(n14938), .A(n14853), .B(n14852), .ZN(
        P2_U3243) );
  XNOR2_X1 U16177 ( .A(n14855), .B(n14862), .ZN(n14856) );
  NAND2_X1 U16178 ( .A1(n14856), .A2(n14924), .ZN(n14860) );
  AOI22_X1 U16179 ( .A1(n14858), .A2(n14885), .B1(n14883), .B2(n14857), .ZN(
        n14859) );
  NAND2_X1 U16180 ( .A1(n14860), .A2(n14859), .ZN(n14992) );
  INV_X1 U16181 ( .A(n14992), .ZN(n14872) );
  XNOR2_X1 U16182 ( .A(n14862), .B(n14861), .ZN(n14986) );
  NAND2_X1 U16183 ( .A1(n14987), .A2(n14874), .ZN(n14863) );
  AND2_X1 U16184 ( .A1(n14864), .A2(n14863), .ZN(n14988) );
  NAND2_X1 U16185 ( .A1(n14988), .A2(n14936), .ZN(n14868) );
  INV_X1 U16186 ( .A(n14865), .ZN(n14866) );
  AOI22_X1 U16187 ( .A1(n14938), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n14866), 
        .B2(n14929), .ZN(n14867) );
  OAI211_X1 U16188 ( .C1(n8169), .C2(n14932), .A(n14868), .B(n14867), .ZN(
        n14869) );
  AOI21_X1 U16189 ( .B1(n14986), .B2(n14870), .A(n14869), .ZN(n14871) );
  OAI21_X1 U16190 ( .B1(n14872), .B2(n14938), .A(n14871), .ZN(P2_U3244) );
  XNOR2_X1 U16191 ( .A(n14881), .B(n14873), .ZN(n14997) );
  INV_X1 U16192 ( .A(n14892), .ZN(n14876) );
  INV_X1 U16193 ( .A(n14874), .ZN(n14875) );
  AOI21_X1 U16194 ( .B1(n14993), .B2(n14876), .A(n14875), .ZN(n14994) );
  AOI22_X1 U16195 ( .A1(n14938), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n14877), 
        .B2(n14929), .ZN(n14878) );
  OAI21_X1 U16196 ( .B1(n14879), .B2(n14932), .A(n14878), .ZN(n14889) );
  OAI21_X1 U16197 ( .B1(n14882), .B2(n14881), .A(n14880), .ZN(n14887) );
  AOI222_X1 U16198 ( .A1(n14924), .A2(n14887), .B1(n14886), .B2(n14885), .C1(
        n14884), .C2(n14883), .ZN(n14996) );
  NOR2_X1 U16199 ( .A1(n14996), .A2(n14938), .ZN(n14888) );
  AOI211_X1 U16200 ( .C1(n14994), .C2(n14936), .A(n14889), .B(n14888), .ZN(
        n14890) );
  OAI21_X1 U16201 ( .B1(n14891), .B2(n14997), .A(n14890), .ZN(P2_U3245) );
  AOI211_X1 U16202 ( .C1(n15001), .C2(n14925), .A(n10363), .B(n14892), .ZN(
        n15000) );
  XNOR2_X1 U16203 ( .A(n14893), .B(n14896), .ZN(n14999) );
  OAI22_X1 U16204 ( .A1(n14895), .A2(n14916), .B1(n14894), .B2(n14914), .ZN(
        n14901) );
  OAI21_X1 U16205 ( .B1(n14911), .B2(n14897), .A(n14896), .ZN(n14898) );
  AND3_X1 U16206 ( .A1(n14899), .A2(n14924), .A3(n14898), .ZN(n14900) );
  AOI211_X1 U16207 ( .C1(n14902), .C2(n14999), .A(n14901), .B(n14900), .ZN(
        n15003) );
  INV_X1 U16208 ( .A(n15003), .ZN(n14903) );
  AOI21_X1 U16209 ( .B1(n15000), .B2(n15711), .A(n14903), .ZN(n14910) );
  INV_X1 U16210 ( .A(n15001), .ZN(n14906) );
  AOI22_X1 U16211 ( .A1(n14938), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n14904), 
        .B2(n14929), .ZN(n14905) );
  OAI21_X1 U16212 ( .B1(n14906), .B2(n14932), .A(n14905), .ZN(n14907) );
  AOI21_X1 U16213 ( .B1(n14999), .B2(n14908), .A(n14907), .ZN(n14909) );
  OAI21_X1 U16214 ( .B1(n14910), .B2(n14938), .A(n14909), .ZN(P2_U3246) );
  OAI21_X1 U16215 ( .B1(n14913), .B2(n14919), .A(n14912), .ZN(n14923) );
  OAI22_X1 U16216 ( .A1(n14917), .A2(n14916), .B1(n14915), .B2(n14914), .ZN(
        n14922) );
  INV_X1 U16217 ( .A(n14918), .ZN(n14920) );
  XNOR2_X1 U16218 ( .A(n14920), .B(n14919), .ZN(n15009) );
  NOR2_X1 U16219 ( .A1(n15009), .A2(n10661), .ZN(n14921) );
  AOI211_X1 U16220 ( .C1(n14924), .C2(n14923), .A(n14922), .B(n14921), .ZN(
        n15008) );
  INV_X1 U16221 ( .A(n14925), .ZN(n14926) );
  AOI21_X1 U16222 ( .B1(n15005), .B2(n14927), .A(n14926), .ZN(n15006) );
  INV_X1 U16223 ( .A(n14928), .ZN(n14930) );
  AOI22_X1 U16224 ( .A1(n14938), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14930), 
        .B2(n14929), .ZN(n14931) );
  OAI21_X1 U16225 ( .B1(n13529), .B2(n14932), .A(n14931), .ZN(n14935) );
  NOR2_X1 U16226 ( .A1(n15009), .A2(n14933), .ZN(n14934) );
  AOI211_X1 U16227 ( .C1(n15006), .C2(n14936), .A(n14935), .B(n14934), .ZN(
        n14937) );
  OAI21_X1 U16228 ( .B1(n15008), .B2(n14938), .A(n14937), .ZN(P2_U3247) );
  MUX2_X1 U16229 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n15034), .S(n16293), .Z(
        P2_U3530) );
  OAI211_X1 U16230 ( .C1(n14942), .C2(n16307), .A(n14941), .B(n14940), .ZN(
        n15035) );
  MUX2_X1 U16231 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n15035), .S(n16293), .Z(
        P2_U3529) );
  AOI21_X1 U16232 ( .B1(n15026), .B2(n14944), .A(n14943), .ZN(n14945) );
  OAI21_X1 U16233 ( .B1(n7418), .B2(n16307), .A(n14948), .ZN(n14950) );
  AOI21_X1 U16234 ( .B1(n14951), .B2(n13663), .A(n14950), .ZN(n14952) );
  NAND2_X1 U16235 ( .A1(n14953), .A2(n14952), .ZN(n15037) );
  MUX2_X1 U16236 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n15037), .S(n16293), .Z(
        P2_U3527) );
  AOI22_X1 U16237 ( .A1(n14955), .A2(n15027), .B1(n15026), .B2(n14954), .ZN(
        n14956) );
  MUX2_X1 U16238 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n15038), .S(n16293), .Z(
        P2_U3526) );
  AOI22_X1 U16239 ( .A1(n14960), .A2(n15027), .B1(n15026), .B2(n14959), .ZN(
        n14961) );
  OAI211_X1 U16240 ( .C1(n14998), .C2(n14963), .A(n14962), .B(n14961), .ZN(
        n15039) );
  MUX2_X1 U16241 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n15039), .S(n16293), .Z(
        P2_U3525) );
  AOI22_X1 U16242 ( .A1(n14965), .A2(n15027), .B1(n15026), .B2(n14964), .ZN(
        n14966) );
  OAI211_X1 U16243 ( .C1(n14998), .C2(n14968), .A(n14967), .B(n14966), .ZN(
        n15040) );
  MUX2_X1 U16244 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n15040), .S(n16293), .Z(
        P2_U3524) );
  AOI22_X1 U16245 ( .A1(n14970), .A2(n15027), .B1(n15026), .B2(n14969), .ZN(
        n14971) );
  OAI211_X1 U16246 ( .C1(n14973), .C2(n14998), .A(n14972), .B(n14971), .ZN(
        n15041) );
  MUX2_X1 U16247 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n15041), .S(n16293), .Z(
        P2_U3523) );
  AOI21_X1 U16248 ( .B1(n15026), .B2(n14975), .A(n14974), .ZN(n14977) );
  OAI211_X1 U16249 ( .C1(n14978), .C2(n15031), .A(n14977), .B(n14976), .ZN(
        n15042) );
  MUX2_X1 U16250 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n15042), .S(n16293), .Z(
        P2_U3522) );
  AND3_X1 U16251 ( .A1(n14980), .A2(n14979), .A3(n16310), .ZN(n14984) );
  OAI22_X1 U16252 ( .A1(n14982), .A2(n10363), .B1(n7971), .B2(n16307), .ZN(
        n14983) );
  MUX2_X1 U16253 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n15043), .S(n16293), .Z(
        P2_U3521) );
  NAND2_X1 U16254 ( .A1(n14986), .A2(n16310), .ZN(n14990) );
  AOI22_X1 U16255 ( .A1(n14988), .A2(n15027), .B1(n15026), .B2(n14987), .ZN(
        n14989) );
  NAND2_X1 U16256 ( .A1(n14990), .A2(n14989), .ZN(n14991) );
  MUX2_X1 U16257 ( .A(n15044), .B(P2_REG1_REG_21__SCAN_IN), .S(n16314), .Z(
        P2_U3520) );
  AOI22_X1 U16258 ( .A1(n14994), .A2(n15027), .B1(n15026), .B2(n14993), .ZN(
        n14995) );
  OAI211_X1 U16259 ( .C1(n14998), .C2(n14997), .A(n14996), .B(n14995), .ZN(
        n15045) );
  MUX2_X1 U16260 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n15045), .S(n16293), .Z(
        P2_U3519) );
  INV_X1 U16261 ( .A(n14999), .ZN(n15004) );
  AOI21_X1 U16262 ( .B1(n15026), .B2(n15001), .A(n15000), .ZN(n15002) );
  OAI211_X1 U16263 ( .C1(n15004), .C2(n15031), .A(n15003), .B(n15002), .ZN(
        n15046) );
  MUX2_X1 U16264 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n15046), .S(n16293), .Z(
        P2_U3518) );
  AOI22_X1 U16265 ( .A1(n15006), .A2(n15027), .B1(n15026), .B2(n15005), .ZN(
        n15007) );
  OAI211_X1 U16266 ( .C1(n15031), .C2(n15009), .A(n15008), .B(n15007), .ZN(
        n15047) );
  MUX2_X1 U16267 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n15047), .S(n16293), .Z(
        P2_U3517) );
  AND2_X1 U16268 ( .A1(n15010), .A2(n16310), .ZN(n15016) );
  INV_X1 U16269 ( .A(n15011), .ZN(n15012) );
  OAI22_X1 U16270 ( .A1(n15013), .A2(n10363), .B1(n15012), .B2(n16307), .ZN(
        n15014) );
  MUX2_X1 U16271 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n15048), .S(n16293), .Z(
        P2_U3516) );
  AOI22_X1 U16272 ( .A1(n15018), .A2(n15027), .B1(n15026), .B2(n15017), .ZN(
        n15022) );
  NAND3_X1 U16273 ( .A1(n7629), .A2(n15019), .A3(n16310), .ZN(n15021) );
  NAND3_X1 U16274 ( .A1(n15023), .A2(n15022), .A3(n15021), .ZN(n15049) );
  MUX2_X1 U16275 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n15049), .S(n16293), .Z(
        P2_U3515) );
  INV_X1 U16276 ( .A(n15024), .ZN(n15032) );
  AOI22_X1 U16277 ( .A1(n15028), .A2(n15027), .B1(n15026), .B2(n15025), .ZN(
        n15029) );
  OAI211_X1 U16278 ( .C1(n15032), .C2(n15031), .A(n15030), .B(n15029), .ZN(
        n15050) );
  MUX2_X1 U16279 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n15050), .S(n16293), .Z(
        P2_U3514) );
  MUX2_X1 U16280 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n15033), .S(n16293), .Z(
        P2_U3503) );
  MUX2_X1 U16281 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n15035), .S(n7419), .Z(
        P2_U3497) );
  MUX2_X1 U16282 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n15037), .S(n7419), .Z(
        P2_U3495) );
  MUX2_X1 U16283 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n15038), .S(n7419), .Z(
        P2_U3494) );
  MUX2_X1 U16284 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n15039), .S(n7419), .Z(
        P2_U3493) );
  MUX2_X1 U16285 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n15040), .S(n7419), .Z(
        P2_U3492) );
  MUX2_X1 U16286 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n15041), .S(n7419), .Z(
        P2_U3491) );
  MUX2_X1 U16287 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n15042), .S(n7419), .Z(
        P2_U3490) );
  MUX2_X1 U16288 ( .A(n15043), .B(P2_REG0_REG_22__SCAN_IN), .S(n16315), .Z(
        P2_U3489) );
  MUX2_X1 U16289 ( .A(n15044), .B(P2_REG0_REG_21__SCAN_IN), .S(n16315), .Z(
        P2_U3488) );
  MUX2_X1 U16290 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n15045), .S(n7419), .Z(
        P2_U3487) );
  MUX2_X1 U16291 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n15046), .S(n7419), .Z(
        P2_U3486) );
  MUX2_X1 U16292 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n15047), .S(n7419), .Z(
        P2_U3484) );
  MUX2_X1 U16293 ( .A(n15048), .B(P2_REG0_REG_17__SCAN_IN), .S(n16315), .Z(
        P2_U3481) );
  MUX2_X1 U16294 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n15049), .S(n7419), .Z(
        P2_U3478) );
  MUX2_X1 U16295 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n15050), .S(n7419), .Z(
        P2_U3475) );
  INV_X1 U16296 ( .A(n15051), .ZN(n15591) );
  INV_X1 U16297 ( .A(n15052), .ZN(n15053) );
  NOR4_X1 U16298 ( .A1(n15053), .A2(P2_IR_REG_30__SCAN_IN), .A3(n10411), .A4(
        P2_U3088), .ZN(n15054) );
  AOI21_X1 U16299 ( .B1(n15059), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n15054), 
        .ZN(n15055) );
  OAI21_X1 U16300 ( .B1(n15591), .B2(n15061), .A(n15055), .ZN(P2_U3296) );
  INV_X1 U16301 ( .A(n13513), .ZN(n15592) );
  OAI222_X1 U16302 ( .A1(n13255), .A2(n15057), .B1(n15061), .B2(n15592), .C1(
        n15056), .C2(P2_U3088), .ZN(P2_U3298) );
  AOI21_X1 U16303 ( .B1(n15059), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n15058), 
        .ZN(n15060) );
  OAI21_X1 U16304 ( .B1(n15062), .B2(n15061), .A(n15060), .ZN(P2_U3299) );
  INV_X1 U16305 ( .A(n15063), .ZN(n15595) );
  OAI222_X1 U16306 ( .A1(n13255), .A2(n15065), .B1(n15061), .B2(n15595), .C1(
        n15064), .C2(P2_U3088), .ZN(P2_U3300) );
  INV_X1 U16307 ( .A(n15066), .ZN(n15069) );
  INV_X1 U16308 ( .A(n15067), .ZN(n15599) );
  OAI222_X1 U16309 ( .A1(n15069), .A2(P2_U3088), .B1(n15061), .B2(n15599), 
        .C1(n15068), .C2(n13255), .ZN(P2_U3301) );
  INV_X1 U16310 ( .A(n15070), .ZN(n15605) );
  INV_X1 U16311 ( .A(n15071), .ZN(n15072) );
  OAI222_X1 U16312 ( .A1(n13255), .A2(n15073), .B1(n15061), .B2(n15605), .C1(
        n15072), .C2(P2_U3088), .ZN(P2_U3302) );
  INV_X1 U16313 ( .A(n15074), .ZN(n15075) );
  MUX2_X1 U16314 ( .A(n15075), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  AOI22_X1 U16315 ( .A1(n16349), .A2(n15312), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n15078) );
  NAND2_X1 U16316 ( .A1(n15167), .A2(n15287), .ZN(n15077) );
  OAI211_X1 U16317 ( .C1(n15079), .C2(n15170), .A(n15078), .B(n15077), .ZN(
        n15080) );
  AOI21_X1 U16318 ( .B1(n15288), .B2(n15173), .A(n15080), .ZN(n15081) );
  INV_X1 U16319 ( .A(n15082), .ZN(n15083) );
  AOI21_X1 U16320 ( .B1(n15085), .B2(n15084), .A(n15083), .ZN(n15092) );
  OAI22_X1 U16321 ( .A1(n15132), .A2(n16296), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15086), .ZN(n15087) );
  AOI21_X1 U16322 ( .B1(n15167), .B2(n15088), .A(n15087), .ZN(n15091) );
  NAND2_X1 U16323 ( .A1(n15089), .A2(n15173), .ZN(n15090) );
  OAI211_X1 U16324 ( .C1(n15092), .C2(n15175), .A(n15091), .B(n15090), .ZN(
        P1_U3215) );
  INV_X1 U16325 ( .A(n15093), .ZN(n15094) );
  AOI21_X1 U16326 ( .B1(n15096), .B2(n15095), .A(n15094), .ZN(n15104) );
  OR2_X1 U16327 ( .A1(n15097), .A2(n15406), .ZN(n15099) );
  NAND2_X1 U16328 ( .A1(n15311), .A2(n15457), .ZN(n15098) );
  AND2_X1 U16329 ( .A1(n15099), .A2(n15098), .ZN(n15509) );
  OAI22_X1 U16330 ( .A1(n15132), .A2(n15509), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15100), .ZN(n15102) );
  NOR2_X1 U16331 ( .A1(n15511), .A2(n16353), .ZN(n15101) );
  AOI211_X1 U16332 ( .C1(n15167), .C2(n15345), .A(n15102), .B(n15101), .ZN(
        n15103) );
  OAI21_X1 U16333 ( .B1(n15104), .B2(n15175), .A(n15103), .ZN(P1_U3216) );
  XOR2_X1 U16334 ( .A(n15106), .B(n15105), .Z(n15111) );
  NAND2_X1 U16335 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n15247)
         );
  OAI21_X1 U16336 ( .B1(n15159), .B2(n15407), .A(n15247), .ZN(n15107) );
  AOI21_X1 U16337 ( .B1(n16351), .B2(n15375), .A(n15107), .ZN(n15108) );
  OAI21_X1 U16338 ( .B1(n15410), .B2(n16361), .A(n15108), .ZN(n15109) );
  AOI21_X1 U16339 ( .B1(n15534), .B2(n15173), .A(n15109), .ZN(n15110) );
  OAI21_X1 U16340 ( .B1(n15111), .B2(n15175), .A(n15110), .ZN(P1_U3219) );
  INV_X1 U16341 ( .A(n15112), .ZN(n15113) );
  AOI21_X1 U16342 ( .B1(n15115), .B2(n15114), .A(n15113), .ZN(n15120) );
  AOI22_X1 U16343 ( .A1(n16351), .A2(n15374), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n15117) );
  NAND2_X1 U16344 ( .A1(n15167), .A2(n15380), .ZN(n15116) );
  OAI211_X1 U16345 ( .C1(n15409), .C2(n15159), .A(n15117), .B(n15116), .ZN(
        n15118) );
  AOI21_X1 U16346 ( .B1(n15525), .B2(n15173), .A(n15118), .ZN(n15119) );
  OAI21_X1 U16347 ( .B1(n15120), .B2(n15175), .A(n15119), .ZN(P1_U3223) );
  XOR2_X1 U16348 ( .A(n15122), .B(n15121), .Z(n15128) );
  AOI22_X1 U16349 ( .A1(n16349), .A2(n15311), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n15124) );
  NAND2_X1 U16350 ( .A1(n15167), .A2(n15315), .ZN(n15123) );
  OAI211_X1 U16351 ( .C1(n15125), .C2(n15170), .A(n15124), .B(n15123), .ZN(
        n15126) );
  AOI21_X1 U16352 ( .B1(n15498), .B2(n15173), .A(n15126), .ZN(n15127) );
  OAI21_X1 U16353 ( .B1(n15128), .B2(n15175), .A(n15127), .ZN(P1_U3225) );
  XOR2_X1 U16354 ( .A(n15129), .B(n15130), .Z(n15136) );
  NOR2_X1 U16355 ( .A1(n16361), .A2(n15439), .ZN(n15134) );
  AND2_X1 U16356 ( .A1(n16322), .A2(n15455), .ZN(n15131) );
  AOI21_X1 U16357 ( .B1(n15182), .B2(n15457), .A(n15131), .ZN(n15548) );
  NAND2_X1 U16358 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n15203)
         );
  OAI21_X1 U16359 ( .B1(n15548), .B2(n15132), .A(n15203), .ZN(n15133) );
  AOI211_X1 U16360 ( .C1(n15550), .C2(n15173), .A(n15134), .B(n15133), .ZN(
        n15135) );
  OAI21_X1 U16361 ( .B1(n15136), .B2(n15175), .A(n15135), .ZN(P1_U3228) );
  OAI21_X1 U16362 ( .B1(n15139), .B2(n15138), .A(n15137), .ZN(n15140) );
  NAND2_X1 U16363 ( .A1(n15140), .A2(n16356), .ZN(n15144) );
  AOI22_X1 U16364 ( .A1(n16351), .A2(n15329), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n15141) );
  OAI21_X1 U16365 ( .B1(n15324), .B2(n15159), .A(n15141), .ZN(n15142) );
  AOI21_X1 U16366 ( .B1(n15333), .B2(n15167), .A(n15142), .ZN(n15143) );
  OAI211_X1 U16367 ( .C1(n15503), .C2(n16353), .A(n15144), .B(n15143), .ZN(
        P1_U3229) );
  AOI21_X1 U16368 ( .B1(n15146), .B2(n15145), .A(n15175), .ZN(n15148) );
  NAND2_X1 U16369 ( .A1(n15148), .A2(n15147), .ZN(n15155) );
  NAND2_X1 U16370 ( .A1(n15181), .A2(n15457), .ZN(n15150) );
  NAND2_X1 U16371 ( .A1(n15421), .A2(n15455), .ZN(n15149) );
  NAND2_X1 U16372 ( .A1(n15150), .A2(n15149), .ZN(n15386) );
  INV_X1 U16373 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n15151) );
  OAI22_X1 U16374 ( .A1(n16361), .A2(n15390), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15151), .ZN(n15152) );
  AOI21_X1 U16375 ( .B1(n15386), .B2(n15153), .A(n15152), .ZN(n15154) );
  OAI211_X1 U16376 ( .C1(n15393), .C2(n16353), .A(n15155), .B(n15154), .ZN(
        P1_U3233) );
  XOR2_X1 U16377 ( .A(n15157), .B(n15156), .Z(n15164) );
  NAND2_X1 U16378 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n15213)
         );
  OAI21_X1 U16379 ( .B1(n15159), .B2(n15158), .A(n15213), .ZN(n15160) );
  AOI21_X1 U16380 ( .B1(n16351), .B2(n15421), .A(n15160), .ZN(n15161) );
  OAI21_X1 U16381 ( .B1(n15429), .B2(n16361), .A(n15161), .ZN(n15162) );
  AOI21_X1 U16382 ( .B1(n15542), .B2(n15173), .A(n15162), .ZN(n15163) );
  OAI21_X1 U16383 ( .B1(n15164), .B2(n15175), .A(n15163), .ZN(P1_U3238) );
  XOR2_X1 U16384 ( .A(n15166), .B(n15165), .Z(n15176) );
  AOI22_X1 U16385 ( .A1(n16349), .A2(n15329), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n15169) );
  NAND2_X1 U16386 ( .A1(n15167), .A2(n15299), .ZN(n15168) );
  OAI211_X1 U16387 ( .C1(n15171), .C2(n15170), .A(n15169), .B(n15168), .ZN(
        n15172) );
  AOI21_X1 U16388 ( .B1(n15491), .B2(n15173), .A(n15172), .ZN(n15174) );
  OAI21_X1 U16389 ( .B1(n15176), .B2(n15175), .A(n15174), .ZN(P1_U3240) );
  MUX2_X1 U16390 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n15177), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U16391 ( .A(n15178), .B(P1_DATAO_REG_30__SCAN_IN), .S(n15196), .Z(
        P1_U3590) );
  MUX2_X1 U16392 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n15179), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16393 ( .A(n15282), .B(P1_DATAO_REG_28__SCAN_IN), .S(n15196), .Z(
        P1_U3588) );
  MUX2_X1 U16394 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n15295), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16395 ( .A(n15312), .B(P1_DATAO_REG_26__SCAN_IN), .S(n15196), .Z(
        P1_U3586) );
  MUX2_X1 U16396 ( .A(n15329), .B(P1_DATAO_REG_25__SCAN_IN), .S(n15196), .Z(
        P1_U3585) );
  MUX2_X1 U16397 ( .A(n15311), .B(P1_DATAO_REG_24__SCAN_IN), .S(n15196), .Z(
        P1_U3584) );
  MUX2_X1 U16398 ( .A(n15180), .B(P1_DATAO_REG_23__SCAN_IN), .S(n15196), .Z(
        P1_U3583) );
  MUX2_X1 U16399 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n15374), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16400 ( .A(n15181), .B(P1_DATAO_REG_21__SCAN_IN), .S(n15196), .Z(
        P1_U3581) );
  MUX2_X1 U16401 ( .A(n15375), .B(P1_DATAO_REG_20__SCAN_IN), .S(n15196), .Z(
        P1_U3580) );
  MUX2_X1 U16402 ( .A(n15421), .B(P1_DATAO_REG_19__SCAN_IN), .S(n15196), .Z(
        P1_U3579) );
  MUX2_X1 U16403 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n15182), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16404 ( .A(n16350), .B(P1_DATAO_REG_17__SCAN_IN), .S(n15196), .Z(
        P1_U3577) );
  MUX2_X1 U16405 ( .A(n16322), .B(P1_DATAO_REG_16__SCAN_IN), .S(n15196), .Z(
        P1_U3576) );
  MUX2_X1 U16406 ( .A(n16348), .B(P1_DATAO_REG_15__SCAN_IN), .S(n15196), .Z(
        P1_U3575) );
  MUX2_X1 U16407 ( .A(n16321), .B(P1_DATAO_REG_14__SCAN_IN), .S(n15196), .Z(
        P1_U3574) );
  MUX2_X1 U16408 ( .A(n15183), .B(P1_DATAO_REG_13__SCAN_IN), .S(n15196), .Z(
        P1_U3573) );
  MUX2_X1 U16409 ( .A(n15184), .B(P1_DATAO_REG_12__SCAN_IN), .S(n15196), .Z(
        P1_U3572) );
  MUX2_X1 U16410 ( .A(n15185), .B(P1_DATAO_REG_11__SCAN_IN), .S(n15196), .Z(
        P1_U3571) );
  MUX2_X1 U16411 ( .A(n15186), .B(P1_DATAO_REG_10__SCAN_IN), .S(n15196), .Z(
        P1_U3570) );
  MUX2_X1 U16412 ( .A(n15187), .B(P1_DATAO_REG_9__SCAN_IN), .S(n15196), .Z(
        P1_U3569) );
  MUX2_X1 U16413 ( .A(n15188), .B(P1_DATAO_REG_8__SCAN_IN), .S(n15196), .Z(
        P1_U3568) );
  MUX2_X1 U16414 ( .A(n15189), .B(P1_DATAO_REG_7__SCAN_IN), .S(n15196), .Z(
        P1_U3567) );
  MUX2_X1 U16415 ( .A(n15190), .B(P1_DATAO_REG_6__SCAN_IN), .S(n15196), .Z(
        P1_U3566) );
  MUX2_X1 U16416 ( .A(n15191), .B(P1_DATAO_REG_5__SCAN_IN), .S(n15196), .Z(
        P1_U3565) );
  MUX2_X1 U16417 ( .A(n15192), .B(P1_DATAO_REG_4__SCAN_IN), .S(n15196), .Z(
        P1_U3564) );
  MUX2_X1 U16418 ( .A(n15193), .B(P1_DATAO_REG_3__SCAN_IN), .S(n15196), .Z(
        P1_U3563) );
  MUX2_X1 U16419 ( .A(n15194), .B(P1_DATAO_REG_2__SCAN_IN), .S(n15196), .Z(
        P1_U3562) );
  MUX2_X1 U16420 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n15195), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U16421 ( .A(n15197), .B(P1_DATAO_REG_0__SCAN_IN), .S(n15196), .Z(
        P1_U3560) );
  NAND2_X1 U16422 ( .A1(n15199), .A2(n15198), .ZN(n15202) );
  INV_X1 U16423 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n15223) );
  NOR2_X1 U16424 ( .A1(n15222), .A2(n15223), .ZN(n15200) );
  AOI21_X1 U16425 ( .B1(n15223), .B2(n15222), .A(n15200), .ZN(n15201) );
  NAND2_X1 U16426 ( .A1(n15201), .A2(n15202), .ZN(n15221) );
  OAI211_X1 U16427 ( .C1(n15202), .C2(n15201), .A(n15780), .B(n15221), .ZN(
        n15212) );
  INV_X1 U16428 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n15204) );
  OAI21_X1 U16429 ( .B1(n15784), .B2(n15204), .A(n15203), .ZN(n15210) );
  XNOR2_X1 U16430 ( .A(n15216), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n15207) );
  AOI211_X1 U16431 ( .C1(n15208), .C2(n15207), .A(n15215), .B(n15240), .ZN(
        n15209) );
  AOI211_X1 U16432 ( .C1(n15778), .C2(n15216), .A(n15210), .B(n15209), .ZN(
        n15211) );
  NAND2_X1 U16433 ( .A1(n15212), .A2(n15211), .ZN(P1_U3260) );
  INV_X1 U16434 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n15214) );
  OAI21_X1 U16435 ( .B1(n15784), .B2(n15214), .A(n15213), .ZN(n15220) );
  INV_X1 U16436 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n15218) );
  NOR2_X1 U16437 ( .A1(n15218), .A2(n15217), .ZN(n15230) );
  AOI211_X1 U16438 ( .C1(n15218), .C2(n15217), .A(n15230), .B(n15240), .ZN(
        n15219) );
  AOI211_X1 U16439 ( .C1(n15778), .C2(n15233), .A(n15220), .B(n15219), .ZN(
        n15226) );
  OAI21_X1 U16440 ( .B1(n15223), .B2(n15222), .A(n15221), .ZN(n15232) );
  XNOR2_X1 U16441 ( .A(n15227), .B(n15232), .ZN(n15224) );
  NAND2_X1 U16442 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n15224), .ZN(n15234) );
  OAI211_X1 U16443 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n15224), .A(n15780), 
        .B(n15234), .ZN(n15225) );
  NAND2_X1 U16444 ( .A1(n15226), .A2(n15225), .ZN(P1_U3261) );
  NOR2_X1 U16445 ( .A1(n15228), .A2(n15227), .ZN(n15229) );
  NOR2_X1 U16446 ( .A1(n15230), .A2(n15229), .ZN(n15231) );
  XNOR2_X1 U16447 ( .A(n15231), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n15243) );
  NAND2_X1 U16448 ( .A1(n15233), .A2(n15232), .ZN(n15235) );
  NAND2_X1 U16449 ( .A1(n15235), .A2(n15234), .ZN(n15236) );
  XOR2_X1 U16450 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n15236), .Z(n15242) );
  INV_X1 U16451 ( .A(n15242), .ZN(n15238) );
  AOI21_X1 U16452 ( .B1(n15238), .B2(n15237), .A(n15778), .ZN(n15239) );
  OAI21_X1 U16453 ( .B1(n15243), .B2(n15240), .A(n15239), .ZN(n15241) );
  INV_X1 U16454 ( .A(n15241), .ZN(n15246) );
  AOI22_X1 U16455 ( .A1(n15243), .A2(n15776), .B1(n15780), .B2(n15242), .ZN(
        n15245) );
  MUX2_X1 U16456 ( .A(n15246), .B(n15245), .S(n15244), .Z(n15248) );
  OAI211_X1 U16457 ( .C1(n8392), .C2(n15784), .A(n15248), .B(n15247), .ZN(
        P1_U3262) );
  NOR2_X1 U16458 ( .A1(n15257), .A2(n15258), .ZN(n15256) );
  XNOR2_X1 U16459 ( .A(n15256), .B(n15253), .ZN(n15249) );
  NAND2_X1 U16460 ( .A1(n15249), .A2(n16247), .ZN(n15467) );
  INV_X1 U16461 ( .A(n15250), .ZN(n15251) );
  OR2_X1 U16462 ( .A1(n15252), .A2(n15251), .ZN(n15470) );
  NOR2_X1 U16463 ( .A1(n16264), .A2(n15470), .ZN(n15259) );
  INV_X1 U16464 ( .A(n15253), .ZN(n15468) );
  NOR2_X1 U16465 ( .A1(n15468), .A2(n16114), .ZN(n15254) );
  AOI211_X1 U16466 ( .C1(n16264), .C2(P1_REG2_REG_31__SCAN_IN), .A(n15259), 
        .B(n15254), .ZN(n15255) );
  OAI21_X1 U16467 ( .B1(n15467), .B2(n16181), .A(n15255), .ZN(P1_U3263) );
  AOI21_X1 U16468 ( .B1(n15258), .B2(n15257), .A(n15256), .ZN(n15469) );
  NAND2_X1 U16469 ( .A1(n15469), .A2(n16073), .ZN(n15261) );
  AOI21_X1 U16470 ( .B1(n16275), .B2(P1_REG2_REG_30__SCAN_IN), .A(n15259), 
        .ZN(n15260) );
  OAI211_X1 U16471 ( .C1(n15472), .C2(n16114), .A(n15261), .B(n15260), .ZN(
        P1_U3264) );
  XNOR2_X1 U16472 ( .A(n15262), .B(n15265), .ZN(n15264) );
  AOI21_X1 U16473 ( .B1(n15264), .B2(n16330), .A(n15263), .ZN(n15483) );
  NAND2_X1 U16474 ( .A1(n15266), .A2(n15265), .ZN(n15267) );
  AOI21_X1 U16475 ( .B1(n7437), .B2(n15274), .A(n16198), .ZN(n15270) );
  NAND2_X1 U16476 ( .A1(n15270), .A2(n15269), .ZN(n15479) );
  NAND2_X1 U16477 ( .A1(n16264), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n15271) );
  OAI21_X1 U16478 ( .B1(n16110), .B2(n15272), .A(n15271), .ZN(n15273) );
  AOI21_X1 U16479 ( .B1(n15274), .B2(n16265), .A(n15273), .ZN(n15275) );
  OAI21_X1 U16480 ( .B1(n15479), .B2(n16181), .A(n15275), .ZN(n15276) );
  AOI21_X1 U16481 ( .B1(n15482), .B2(n15366), .A(n15276), .ZN(n15277) );
  OAI21_X1 U16482 ( .B1(n15483), .B2(n16264), .A(n15277), .ZN(P1_U3265) );
  XNOR2_X1 U16483 ( .A(n15278), .B(n15280), .ZN(n15286) );
  OAI21_X1 U16484 ( .B1(n15281), .B2(n15280), .A(n15279), .ZN(n15488) );
  INV_X1 U16485 ( .A(n15488), .ZN(n15284) );
  AOI22_X1 U16486 ( .A1(n15455), .A2(n15312), .B1(n15282), .B2(n15457), .ZN(
        n15283) );
  OAI21_X1 U16487 ( .B1(n15284), .B2(n16254), .A(n15283), .ZN(n15285) );
  OAI21_X1 U16488 ( .B1(n15297), .B2(n15485), .A(n7437), .ZN(n15486) );
  AOI22_X1 U16489 ( .A1(n16264), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n15287), 
        .B2(n16262), .ZN(n15290) );
  NAND2_X1 U16490 ( .A1(n15288), .A2(n16265), .ZN(n15289) );
  OAI211_X1 U16491 ( .C1(n15486), .C2(n15416), .A(n15290), .B(n15289), .ZN(
        n15291) );
  AOI21_X1 U16492 ( .B1(n15488), .B2(n16270), .A(n15291), .ZN(n15292) );
  OAI21_X1 U16493 ( .B1(n15490), .B2(n16264), .A(n15292), .ZN(P1_U3266) );
  XNOR2_X1 U16494 ( .A(n15294), .B(n15293), .ZN(n15296) );
  AOI222_X1 U16495 ( .A1(n16330), .A2(n15296), .B1(n15295), .B2(n15457), .C1(
        n15329), .C2(n15455), .ZN(n15494) );
  INV_X1 U16496 ( .A(n15309), .ZN(n15298) );
  AOI21_X1 U16497 ( .B1(n15491), .B2(n15298), .A(n15297), .ZN(n15492) );
  AOI22_X1 U16498 ( .A1(n16264), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n15299), 
        .B2(n16262), .ZN(n15300) );
  OAI21_X1 U16499 ( .B1(n15301), .B2(n16114), .A(n15300), .ZN(n15305) );
  XNOR2_X1 U16500 ( .A(n15303), .B(n15302), .ZN(n15495) );
  NOR2_X1 U16501 ( .A1(n15495), .A2(n15466), .ZN(n15304) );
  AOI211_X1 U16502 ( .C1(n15492), .C2(n16073), .A(n15305), .B(n15304), .ZN(
        n15306) );
  OAI21_X1 U16503 ( .B1(n16264), .B2(n15494), .A(n15306), .ZN(P1_U3267) );
  OAI21_X1 U16504 ( .B1(n7539), .B2(n15308), .A(n15307), .ZN(n15502) );
  INV_X1 U16505 ( .A(n15331), .ZN(n15310) );
  AOI211_X1 U16506 ( .C1(n15498), .C2(n15310), .A(n16198), .B(n15309), .ZN(
        n15496) );
  NAND2_X1 U16507 ( .A1(n15311), .A2(n15455), .ZN(n15314) );
  NAND2_X1 U16508 ( .A1(n15312), .A2(n15457), .ZN(n15313) );
  NAND2_X1 U16509 ( .A1(n15314), .A2(n15313), .ZN(n15497) );
  AOI22_X1 U16510 ( .A1(n16179), .A2(n15497), .B1(n15315), .B2(n16262), .ZN(
        n15317) );
  NAND2_X1 U16511 ( .A1(n16264), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n15316) );
  OAI211_X1 U16512 ( .C1(n15318), .C2(n16114), .A(n15317), .B(n15316), .ZN(
        n15319) );
  AOI21_X1 U16513 ( .B1(n15496), .B2(n16269), .A(n15319), .ZN(n15323) );
  OAI21_X1 U16514 ( .B1(n7528), .B2(n15321), .A(n15320), .ZN(n15499) );
  NAND2_X1 U16515 ( .A1(n15499), .A2(n15418), .ZN(n15322) );
  OAI211_X1 U16516 ( .C1(n15502), .C2(n15466), .A(n15323), .B(n15322), .ZN(
        P1_U3268) );
  NOR2_X1 U16517 ( .A1(n15324), .A2(n15406), .ZN(n15328) );
  AOI211_X1 U16518 ( .C1(n15330), .C2(n15326), .A(n16280), .B(n15325), .ZN(
        n15327) );
  AOI211_X1 U16519 ( .C1(n15457), .C2(n15329), .A(n15328), .B(n15327), .ZN(
        n15507) );
  OAI21_X1 U16520 ( .B1(n15330), .B2(n7497), .A(n8297), .ZN(n15506) );
  AND2_X1 U16521 ( .A1(n15343), .A2(n15334), .ZN(n15332) );
  OR2_X1 U16522 ( .A1(n15332), .A2(n15331), .ZN(n15504) );
  AOI22_X1 U16523 ( .A1(n16264), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n15333), 
        .B2(n16262), .ZN(n15336) );
  NAND2_X1 U16524 ( .A1(n15334), .A2(n16265), .ZN(n15335) );
  OAI211_X1 U16525 ( .C1(n15504), .C2(n15416), .A(n15336), .B(n15335), .ZN(
        n15337) );
  AOI21_X1 U16526 ( .B1(n15506), .B2(n15366), .A(n15337), .ZN(n15338) );
  OAI21_X1 U16527 ( .B1(n16264), .B2(n15507), .A(n15338), .ZN(P1_U3269) );
  XNOR2_X1 U16528 ( .A(n15339), .B(n15342), .ZN(n15515) );
  AOI21_X1 U16529 ( .B1(n15342), .B2(n15341), .A(n15340), .ZN(n15513) );
  AOI21_X1 U16530 ( .B1(n15349), .B2(n15360), .A(n16198), .ZN(n15344) );
  NAND2_X1 U16531 ( .A1(n15344), .A2(n15343), .ZN(n15510) );
  NAND2_X1 U16532 ( .A1(n16264), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n15347) );
  NAND2_X1 U16533 ( .A1(n16262), .A2(n15345), .ZN(n15346) );
  OAI211_X1 U16534 ( .C1(n16264), .C2(n15509), .A(n15347), .B(n15346), .ZN(
        n15348) );
  AOI21_X1 U16535 ( .B1(n15349), .B2(n16265), .A(n15348), .ZN(n15350) );
  OAI21_X1 U16536 ( .B1(n15510), .B2(n16181), .A(n15350), .ZN(n15351) );
  AOI21_X1 U16537 ( .B1(n15513), .B2(n15366), .A(n15351), .ZN(n15352) );
  OAI21_X1 U16538 ( .B1(n15515), .B2(n15462), .A(n15352), .ZN(P1_U3270) );
  AOI21_X1 U16539 ( .B1(n15358), .B2(n15353), .A(n7657), .ZN(n15356) );
  INV_X1 U16540 ( .A(n15354), .ZN(n15355) );
  OAI21_X1 U16541 ( .B1(n15356), .B2(n16280), .A(n15355), .ZN(n15519) );
  INV_X1 U16542 ( .A(n15519), .ZN(n15368) );
  OAI21_X1 U16543 ( .B1(n15359), .B2(n15358), .A(n15357), .ZN(n15520) );
  OAI21_X1 U16544 ( .B1(n7417), .B2(n15378), .A(n15360), .ZN(n15517) );
  AOI22_X1 U16545 ( .A1(n16264), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n15361), 
        .B2(n16262), .ZN(n15364) );
  NAND2_X1 U16546 ( .A1(n15362), .A2(n16265), .ZN(n15363) );
  OAI211_X1 U16547 ( .C1(n15517), .C2(n15416), .A(n15364), .B(n15363), .ZN(
        n15365) );
  AOI21_X1 U16548 ( .B1(n15520), .B2(n15366), .A(n15365), .ZN(n15367) );
  OAI21_X1 U16549 ( .B1(n16264), .B2(n15368), .A(n15367), .ZN(P1_U3271) );
  XNOR2_X1 U16550 ( .A(n15370), .B(n15369), .ZN(n15527) );
  OAI211_X1 U16551 ( .C1(n15373), .C2(n15372), .A(n15371), .B(n16330), .ZN(
        n15377) );
  AOI22_X1 U16552 ( .A1(n15375), .A2(n15455), .B1(n15457), .B2(n15374), .ZN(
        n15376) );
  NAND2_X1 U16553 ( .A1(n15377), .A2(n15376), .ZN(n15523) );
  AND2_X1 U16554 ( .A1(n15525), .A2(n15388), .ZN(n15379) );
  OR2_X1 U16555 ( .A1(n15379), .A2(n15378), .ZN(n15522) );
  AOI22_X1 U16556 ( .A1(n15380), .A2(n16262), .B1(n16264), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n15382) );
  NAND2_X1 U16557 ( .A1(n15525), .A2(n16265), .ZN(n15381) );
  OAI211_X1 U16558 ( .C1(n15522), .C2(n15416), .A(n15382), .B(n15381), .ZN(
        n15383) );
  AOI21_X1 U16559 ( .B1(n15523), .B2(n16179), .A(n15383), .ZN(n15384) );
  OAI21_X1 U16560 ( .B1(n15527), .B2(n15466), .A(n15384), .ZN(P1_U3272) );
  AOI21_X1 U16561 ( .B1(n15385), .B2(n15396), .A(n16280), .ZN(n15387) );
  AOI21_X1 U16562 ( .B1(n15387), .B2(n7438), .A(n15386), .ZN(n15531) );
  INV_X1 U16563 ( .A(n15388), .ZN(n15389) );
  AOI21_X1 U16564 ( .B1(n15528), .B2(n15405), .A(n15389), .ZN(n15529) );
  INV_X1 U16565 ( .A(n15390), .ZN(n15391) );
  AOI22_X1 U16566 ( .A1(n15391), .A2(n16262), .B1(n16264), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n15392) );
  OAI21_X1 U16567 ( .B1(n15393), .B2(n16114), .A(n15392), .ZN(n15398) );
  OAI21_X1 U16568 ( .B1(n15394), .B2(n15396), .A(n15395), .ZN(n15532) );
  NOR2_X1 U16569 ( .A1(n15532), .A2(n15466), .ZN(n15397) );
  AOI211_X1 U16570 ( .C1(n15529), .C2(n16073), .A(n15398), .B(n15397), .ZN(
        n15399) );
  OAI21_X1 U16571 ( .B1(n16264), .B2(n15531), .A(n15399), .ZN(P1_U3273) );
  XNOR2_X1 U16572 ( .A(n15400), .B(n15402), .ZN(n15540) );
  OAI21_X1 U16573 ( .B1(n15403), .B2(n15402), .A(n15401), .ZN(n15538) );
  INV_X1 U16574 ( .A(n15404), .ZN(n15427) );
  OAI21_X1 U16575 ( .B1(n15412), .B2(n15427), .A(n15405), .ZN(n15536) );
  OAI22_X1 U16576 ( .A1(n15409), .A2(n15408), .B1(n15407), .B2(n15406), .ZN(
        n15533) );
  INV_X1 U16577 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n15411) );
  OAI22_X1 U16578 ( .A1(n16179), .A2(n15411), .B1(n15410), .B2(n16110), .ZN(
        n15414) );
  NOR2_X1 U16579 ( .A1(n15412), .A2(n16114), .ZN(n15413) );
  AOI211_X1 U16580 ( .C1(n16179), .C2(n15533), .A(n15414), .B(n15413), .ZN(
        n15415) );
  OAI21_X1 U16581 ( .B1(n15416), .B2(n15536), .A(n15415), .ZN(n15417) );
  AOI21_X1 U16582 ( .B1(n15418), .B2(n15538), .A(n15417), .ZN(n15419) );
  OAI21_X1 U16583 ( .B1(n15540), .B2(n15466), .A(n15419), .ZN(P1_U3274) );
  XOR2_X1 U16584 ( .A(n15423), .B(n15420), .Z(n15546) );
  AOI22_X1 U16585 ( .A1(n15421), .A2(n15457), .B1(n15455), .B2(n16350), .ZN(
        n15426) );
  OAI211_X1 U16586 ( .C1(n15424), .C2(n15423), .A(n15422), .B(n16330), .ZN(
        n15425) );
  OAI211_X1 U16587 ( .C1(n15546), .C2(n16254), .A(n15426), .B(n15425), .ZN(
        n15541) );
  NAND2_X1 U16588 ( .A1(n15541), .A2(n16179), .ZN(n15434) );
  AOI21_X1 U16589 ( .B1(n15542), .B2(n15438), .A(n15427), .ZN(n15543) );
  NOR2_X1 U16590 ( .A1(n15428), .A2(n16114), .ZN(n15432) );
  INV_X1 U16591 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n15430) );
  OAI22_X1 U16592 ( .A1(n16179), .A2(n15430), .B1(n15429), .B2(n16110), .ZN(
        n15431) );
  AOI211_X1 U16593 ( .C1(n15543), .C2(n16073), .A(n15432), .B(n15431), .ZN(
        n15433) );
  OAI211_X1 U16594 ( .C1(n15546), .C2(n15435), .A(n15434), .B(n15433), .ZN(
        P1_U3275) );
  XNOR2_X1 U16595 ( .A(n15436), .B(n15443), .ZN(n15557) );
  NAND2_X1 U16596 ( .A1(n15550), .A2(n15451), .ZN(n15437) );
  NAND2_X1 U16597 ( .A1(n15438), .A2(n15437), .ZN(n15552) );
  INV_X1 U16598 ( .A(n15552), .ZN(n15448) );
  NAND2_X1 U16599 ( .A1(n15550), .A2(n16265), .ZN(n15442) );
  OAI22_X1 U16600 ( .A1(n15548), .A2(n16264), .B1(n15439), .B2(n16110), .ZN(
        n15440) );
  INV_X1 U16601 ( .A(n15440), .ZN(n15441) );
  OAI211_X1 U16602 ( .C1(n16179), .C2(n15223), .A(n15442), .B(n15441), .ZN(
        n15447) );
  NOR2_X1 U16603 ( .A1(n15444), .A2(n15443), .ZN(n15547) );
  INV_X1 U16604 ( .A(n15554), .ZN(n15445) );
  NOR3_X1 U16605 ( .A1(n15547), .A2(n15445), .A3(n15466), .ZN(n15446) );
  AOI211_X1 U16606 ( .C1(n15448), .C2(n16073), .A(n15447), .B(n15446), .ZN(
        n15449) );
  OAI21_X1 U16607 ( .B1(n15557), .B2(n15462), .A(n15449), .ZN(P1_U3276) );
  XOR2_X1 U16608 ( .A(n15461), .B(n15450), .Z(n15564) );
  INV_X1 U16609 ( .A(n15451), .ZN(n15452) );
  AOI21_X1 U16610 ( .B1(n15454), .B2(n15453), .A(n15452), .ZN(n15562) );
  AND2_X1 U16611 ( .A1(n16348), .A2(n15455), .ZN(n15456) );
  AOI21_X1 U16612 ( .B1(n16350), .B2(n15457), .A(n15456), .ZN(n15558) );
  OAI22_X1 U16613 ( .A1(n16264), .A2(n15558), .B1(n16360), .B2(n16110), .ZN(
        n15458) );
  AOI21_X1 U16614 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n16264), .A(n15458), 
        .ZN(n15459) );
  OAI21_X1 U16615 ( .B1(n16354), .B2(n16114), .A(n15459), .ZN(n15464) );
  AOI21_X1 U16616 ( .B1(n15461), .B2(n15460), .A(n7563), .ZN(n15559) );
  NOR2_X1 U16617 ( .A1(n15559), .A2(n15462), .ZN(n15463) );
  AOI211_X1 U16618 ( .C1(n15562), .C2(n16073), .A(n15464), .B(n15463), .ZN(
        n15465) );
  OAI21_X1 U16619 ( .B1(n15564), .B2(n15466), .A(n15465), .ZN(P1_U3277) );
  OAI211_X1 U16620 ( .C1(n15468), .C2(n16333), .A(n15467), .B(n15470), .ZN(
        n15566) );
  MUX2_X1 U16621 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n15566), .S(n16341), .Z(
        P1_U3559) );
  NAND2_X1 U16622 ( .A1(n15469), .A2(n16247), .ZN(n15471) );
  OAI211_X1 U16623 ( .C1(n15472), .C2(n16333), .A(n15471), .B(n15470), .ZN(
        n15567) );
  MUX2_X1 U16624 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n15567), .S(n16341), .Z(
        P1_U3558) );
  OAI21_X1 U16625 ( .B1(n15474), .B2(n16333), .A(n15473), .ZN(n15475) );
  MUX2_X1 U16626 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n15568), .S(n16341), .Z(
        P1_U3557) );
  OAI21_X1 U16627 ( .B1(n15480), .B2(n16333), .A(n15479), .ZN(n15481) );
  NAND2_X1 U16628 ( .A1(n15484), .A2(n15483), .ZN(n15569) );
  MUX2_X1 U16629 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n15569), .S(n16341), .Z(
        P1_U3556) );
  OAI22_X1 U16630 ( .A1(n15486), .A2(n16198), .B1(n15485), .B2(n16333), .ZN(
        n15487) );
  AOI21_X1 U16631 ( .B1(n15488), .B2(n16257), .A(n15487), .ZN(n15489) );
  NAND2_X1 U16632 ( .A1(n15490), .A2(n15489), .ZN(n15570) );
  MUX2_X1 U16633 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15570), .S(n16341), .Z(
        P1_U3555) );
  AOI22_X1 U16634 ( .A1(n15492), .A2(n16247), .B1(n16278), .B2(n15491), .ZN(
        n15493) );
  OAI211_X1 U16635 ( .C1(n15495), .C2(n16299), .A(n15494), .B(n15493), .ZN(
        n15571) );
  MUX2_X1 U16636 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15571), .S(n16341), .Z(
        P1_U3554) );
  AOI211_X1 U16637 ( .C1(n16278), .C2(n15498), .A(n15497), .B(n15496), .ZN(
        n15501) );
  NAND2_X1 U16638 ( .A1(n15499), .A2(n16330), .ZN(n15500) );
  OAI211_X1 U16639 ( .C1(n15502), .C2(n16299), .A(n15501), .B(n15500), .ZN(
        n15572) );
  MUX2_X1 U16640 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n15572), .S(n16341), .Z(
        P1_U3553) );
  OAI22_X1 U16641 ( .A1(n15504), .A2(n16198), .B1(n15503), .B2(n16333), .ZN(
        n15505) );
  AOI21_X1 U16642 ( .B1(n15506), .B2(n16337), .A(n15505), .ZN(n15508) );
  NAND2_X1 U16643 ( .A1(n15508), .A2(n15507), .ZN(n15573) );
  MUX2_X1 U16644 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n15573), .S(n16341), .Z(
        P1_U3552) );
  OAI211_X1 U16645 ( .C1(n15511), .C2(n16333), .A(n15510), .B(n15509), .ZN(
        n15512) );
  AOI21_X1 U16646 ( .B1(n15513), .B2(n16337), .A(n15512), .ZN(n15514) );
  OAI21_X1 U16647 ( .B1(n16280), .B2(n15515), .A(n15514), .ZN(n15574) );
  MUX2_X1 U16648 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15574), .S(n16341), .Z(
        P1_U3551) );
  OAI22_X1 U16649 ( .A1(n15517), .A2(n16198), .B1(n7417), .B2(n16333), .ZN(
        n15518) );
  AOI211_X1 U16650 ( .C1(n15520), .C2(n16337), .A(n15519), .B(n15518), .ZN(
        n15521) );
  INV_X1 U16651 ( .A(n15521), .ZN(n15575) );
  MUX2_X1 U16652 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15575), .S(n16341), .Z(
        P1_U3550) );
  NOR2_X1 U16653 ( .A1(n15522), .A2(n16198), .ZN(n15524) );
  AOI211_X1 U16654 ( .C1(n16278), .C2(n15525), .A(n15524), .B(n15523), .ZN(
        n15526) );
  OAI21_X1 U16655 ( .B1(n15527), .B2(n16299), .A(n15526), .ZN(n15576) );
  MUX2_X1 U16656 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n15576), .S(n16341), .Z(
        P1_U3549) );
  AOI22_X1 U16657 ( .A1(n15529), .A2(n16247), .B1(n16278), .B2(n15528), .ZN(
        n15530) );
  OAI211_X1 U16658 ( .C1(n15532), .C2(n16299), .A(n15531), .B(n15530), .ZN(
        n15577) );
  MUX2_X1 U16659 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n15577), .S(n16341), .Z(
        P1_U3548) );
  AOI21_X1 U16660 ( .B1(n15534), .B2(n16278), .A(n15533), .ZN(n15535) );
  OAI21_X1 U16661 ( .B1(n15536), .B2(n16198), .A(n15535), .ZN(n15537) );
  AOI21_X1 U16662 ( .B1(n15538), .B2(n16330), .A(n15537), .ZN(n15539) );
  OAI21_X1 U16663 ( .B1(n15540), .B2(n16299), .A(n15539), .ZN(n15578) );
  MUX2_X1 U16664 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15578), .S(n16341), .Z(
        P1_U3547) );
  INV_X1 U16665 ( .A(n15541), .ZN(n15545) );
  AOI22_X1 U16666 ( .A1(n15543), .A2(n16247), .B1(n16278), .B2(n15542), .ZN(
        n15544) );
  OAI211_X1 U16667 ( .C1(n15546), .C2(n16135), .A(n15545), .B(n15544), .ZN(
        n15579) );
  MUX2_X1 U16668 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15579), .S(n16341), .Z(
        P1_U3546) );
  NOR2_X1 U16669 ( .A1(n15547), .A2(n16299), .ZN(n15555) );
  INV_X1 U16670 ( .A(n15548), .ZN(n15549) );
  AOI21_X1 U16671 ( .B1(n15550), .B2(n16278), .A(n15549), .ZN(n15551) );
  OAI21_X1 U16672 ( .B1(n15552), .B2(n16198), .A(n15551), .ZN(n15553) );
  AOI21_X1 U16673 ( .B1(n15555), .B2(n15554), .A(n15553), .ZN(n15556) );
  OAI21_X1 U16674 ( .B1(n16280), .B2(n15557), .A(n15556), .ZN(n15580) );
  MUX2_X1 U16675 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15580), .S(n16341), .Z(
        P1_U3545) );
  OAI21_X1 U16676 ( .B1(n16354), .B2(n16333), .A(n15558), .ZN(n15561) );
  NOR2_X1 U16677 ( .A1(n15559), .A2(n16280), .ZN(n15560) );
  AOI211_X1 U16678 ( .C1(n16247), .C2(n15562), .A(n15561), .B(n15560), .ZN(
        n15563) );
  OAI21_X1 U16679 ( .B1(n15564), .B2(n16299), .A(n15563), .ZN(n15581) );
  MUX2_X1 U16680 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15581), .S(n16341), .Z(
        P1_U3544) );
  MUX2_X1 U16681 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n15565), .S(n16341), .Z(
        P1_U3534) );
  MUX2_X1 U16682 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n15566), .S(n16345), .Z(
        P1_U3527) );
  MUX2_X1 U16683 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n15567), .S(n16345), .Z(
        P1_U3526) );
  MUX2_X1 U16684 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n15568), .S(n16345), .Z(
        P1_U3525) );
  MUX2_X1 U16685 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n15569), .S(n16345), .Z(
        P1_U3524) );
  MUX2_X1 U16686 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n15570), .S(n16345), .Z(
        P1_U3523) );
  MUX2_X1 U16687 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15571), .S(n16345), .Z(
        P1_U3522) );
  MUX2_X1 U16688 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n15572), .S(n16345), .Z(
        P1_U3521) );
  MUX2_X1 U16689 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n15573), .S(n16345), .Z(
        P1_U3520) );
  MUX2_X1 U16690 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15574), .S(n16345), .Z(
        P1_U3519) );
  MUX2_X1 U16691 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15575), .S(n16345), .Z(
        P1_U3518) );
  MUX2_X1 U16692 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n15576), .S(n16345), .Z(
        P1_U3517) );
  MUX2_X1 U16693 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n15577), .S(n16345), .Z(
        P1_U3516) );
  MUX2_X1 U16694 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15578), .S(n16345), .Z(
        P1_U3515) );
  MUX2_X1 U16695 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15579), .S(n16345), .Z(
        P1_U3513) );
  MUX2_X1 U16696 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15580), .S(n16345), .Z(
        P1_U3510) );
  MUX2_X1 U16697 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15581), .S(n16345), .Z(
        P1_U3507) );
  INV_X1 U16698 ( .A(n15582), .ZN(n15584) );
  MUX2_X1 U16699 ( .A(P1_D_REG_1__SCAN_IN), .B(n15585), .S(n15640), .Z(
        P1_U3446) );
  MUX2_X1 U16700 ( .A(P1_D_REG_0__SCAN_IN), .B(n15586), .S(n15640), .Z(
        P1_U3445) );
  NOR4_X1 U16701 ( .A1(n15588), .A2(P1_IR_REG_30__SCAN_IN), .A3(n7671), .A4(
        P1_U3086), .ZN(n15589) );
  AOI21_X1 U16702 ( .B1(n15601), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n15589), 
        .ZN(n15590) );
  OAI21_X1 U16703 ( .B1(n15591), .B2(n15604), .A(n15590), .ZN(P1_U3324) );
  OAI222_X1 U16704 ( .A1(n15597), .A2(n15593), .B1(n15604), .B2(n15592), .C1(
        n8380), .C2(P1_U3086), .ZN(P1_U3326) );
  OAI222_X1 U16705 ( .A1(n15597), .A2(n15596), .B1(n15604), .B2(n15595), .C1(
        P1_U3086), .C2(n15594), .ZN(P1_U3328) );
  OAI222_X1 U16706 ( .A1(P1_U3086), .A2(n15600), .B1(n15604), .B2(n15599), 
        .C1(n15598), .C2(n15597), .ZN(P1_U3329) );
  AOI22_X1 U16707 ( .A1(n15602), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n15601), .ZN(n15603) );
  OAI21_X1 U16708 ( .B1(n15605), .B2(n15604), .A(n15603), .ZN(P1_U3330) );
  MUX2_X1 U16709 ( .A(n15607), .B(n15606), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  MUX2_X1 U16710 ( .A(n15608), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16711 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n15609) );
  NOR2_X1 U16712 ( .A1(n15640), .A2(n15609), .ZN(P1_U3323) );
  INV_X1 U16713 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n15610) );
  NOR2_X1 U16714 ( .A1(n15640), .A2(n15610), .ZN(P1_U3322) );
  INV_X1 U16715 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n15611) );
  NOR2_X1 U16716 ( .A1(n15640), .A2(n15611), .ZN(P1_U3321) );
  INV_X1 U16717 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n15612) );
  NOR2_X1 U16718 ( .A1(n15640), .A2(n15612), .ZN(P1_U3320) );
  INV_X1 U16719 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n15613) );
  NOR2_X1 U16720 ( .A1(n15640), .A2(n15613), .ZN(P1_U3319) );
  INV_X1 U16721 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n15614) );
  NOR2_X1 U16722 ( .A1(n15640), .A2(n15614), .ZN(P1_U3318) );
  INV_X1 U16723 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n15615) );
  NOR2_X1 U16724 ( .A1(n15625), .A2(n15615), .ZN(P1_U3317) );
  INV_X1 U16725 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n15616) );
  NOR2_X1 U16726 ( .A1(n15625), .A2(n15616), .ZN(P1_U3316) );
  INV_X1 U16727 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n15617) );
  NOR2_X1 U16728 ( .A1(n15625), .A2(n15617), .ZN(P1_U3315) );
  INV_X1 U16729 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n15618) );
  NOR2_X1 U16730 ( .A1(n15625), .A2(n15618), .ZN(P1_U3314) );
  INV_X1 U16731 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n15619) );
  NOR2_X1 U16732 ( .A1(n15625), .A2(n15619), .ZN(P1_U3313) );
  INV_X1 U16733 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n15620) );
  NOR2_X1 U16734 ( .A1(n15625), .A2(n15620), .ZN(P1_U3312) );
  INV_X1 U16735 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n15621) );
  NOR2_X1 U16736 ( .A1(n15625), .A2(n15621), .ZN(P1_U3311) );
  INV_X1 U16737 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n15622) );
  NOR2_X1 U16738 ( .A1(n15625), .A2(n15622), .ZN(P1_U3310) );
  INV_X1 U16739 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n15623) );
  NOR2_X1 U16740 ( .A1(n15625), .A2(n15623), .ZN(P1_U3309) );
  INV_X1 U16741 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n15624) );
  NOR2_X1 U16742 ( .A1(n15625), .A2(n15624), .ZN(P1_U3308) );
  INV_X1 U16743 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n15626) );
  NOR2_X1 U16744 ( .A1(n15640), .A2(n15626), .ZN(P1_U3307) );
  INV_X1 U16745 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n15627) );
  NOR2_X1 U16746 ( .A1(n15640), .A2(n15627), .ZN(P1_U3306) );
  INV_X1 U16747 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n15628) );
  NOR2_X1 U16748 ( .A1(n15640), .A2(n15628), .ZN(P1_U3305) );
  INV_X1 U16749 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n15629) );
  NOR2_X1 U16750 ( .A1(n15640), .A2(n15629), .ZN(P1_U3304) );
  INV_X1 U16751 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n15630) );
  NOR2_X1 U16752 ( .A1(n15640), .A2(n15630), .ZN(P1_U3303) );
  INV_X1 U16753 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n15631) );
  NOR2_X1 U16754 ( .A1(n15640), .A2(n15631), .ZN(P1_U3302) );
  INV_X1 U16755 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n15632) );
  NOR2_X1 U16756 ( .A1(n15640), .A2(n15632), .ZN(P1_U3301) );
  INV_X1 U16757 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n15633) );
  NOR2_X1 U16758 ( .A1(n15640), .A2(n15633), .ZN(P1_U3300) );
  INV_X1 U16759 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n15634) );
  NOR2_X1 U16760 ( .A1(n15640), .A2(n15634), .ZN(P1_U3299) );
  INV_X1 U16761 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n15635) );
  NOR2_X1 U16762 ( .A1(n15640), .A2(n15635), .ZN(P1_U3298) );
  INV_X1 U16763 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n15636) );
  NOR2_X1 U16764 ( .A1(n15640), .A2(n15636), .ZN(P1_U3297) );
  INV_X1 U16765 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n15637) );
  NOR2_X1 U16766 ( .A1(n15640), .A2(n15637), .ZN(P1_U3296) );
  INV_X1 U16767 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n15638) );
  NOR2_X1 U16768 ( .A1(n15640), .A2(n15638), .ZN(P1_U3295) );
  INV_X1 U16769 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n15639) );
  NOR2_X1 U16770 ( .A1(n15640), .A2(n15639), .ZN(P1_U3294) );
  OAI21_X1 U16771 ( .B1(n15647), .B2(P2_D_REG_1__SCAN_IN), .A(n15641), .ZN(
        n15642) );
  INV_X1 U16772 ( .A(n15642), .ZN(P2_U3417) );
  INV_X1 U16773 ( .A(n15643), .ZN(n15644) );
  AND2_X1 U16774 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15645), .ZN(P2_U3295) );
  AND2_X1 U16775 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15645), .ZN(P2_U3294) );
  AND2_X1 U16776 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15645), .ZN(P2_U3293) );
  AND2_X1 U16777 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15645), .ZN(P2_U3292) );
  AND2_X1 U16778 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15645), .ZN(P2_U3291) );
  AND2_X1 U16779 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15645), .ZN(P2_U3290) );
  AND2_X1 U16780 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15645), .ZN(P2_U3289) );
  AND2_X1 U16781 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15645), .ZN(P2_U3288) );
  AND2_X1 U16782 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15645), .ZN(P2_U3287) );
  AND2_X1 U16783 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15645), .ZN(P2_U3286) );
  AND2_X1 U16784 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15645), .ZN(P2_U3285) );
  AND2_X1 U16785 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15645), .ZN(P2_U3284) );
  AND2_X1 U16786 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15645), .ZN(P2_U3283) );
  AND2_X1 U16787 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15645), .ZN(P2_U3282) );
  AND2_X1 U16788 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15645), .ZN(P2_U3281) );
  AND2_X1 U16789 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15645), .ZN(P2_U3280) );
  AND2_X1 U16790 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15645), .ZN(P2_U3279) );
  AND2_X1 U16791 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15645), .ZN(P2_U3278) );
  AND2_X1 U16792 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15645), .ZN(P2_U3277) );
  AND2_X1 U16793 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15645), .ZN(P2_U3276) );
  AND2_X1 U16794 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15645), .ZN(P2_U3275) );
  AND2_X1 U16795 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15645), .ZN(P2_U3274) );
  AND2_X1 U16796 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15645), .ZN(P2_U3273) );
  AND2_X1 U16797 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15645), .ZN(P2_U3272) );
  AND2_X1 U16798 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15645), .ZN(P2_U3271) );
  AND2_X1 U16799 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15645), .ZN(P2_U3270) );
  AND2_X1 U16800 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15645), .ZN(P2_U3269) );
  AND2_X1 U16801 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15645), .ZN(P2_U3268) );
  AND2_X1 U16802 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15645), .ZN(P2_U3267) );
  AND2_X1 U16803 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15645), .ZN(P2_U3266) );
  NOR2_X1 U16804 ( .A1(n15683), .A2(P2_U3947), .ZN(P2_U3087) );
  NOR2_X1 U16805 ( .A1(P3_U3897), .A2(n15646), .ZN(P3_U3150) );
  OAI22_X1 U16806 ( .A1(n15649), .A2(n15648), .B1(P2_D_REG_0__SCAN_IN), .B2(
        n15647), .ZN(n15650) );
  INV_X1 U16807 ( .A(n15650), .ZN(P2_U3416) );
  OAI22_X1 U16808 ( .A1(n15724), .A2(n15652), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15651), .ZN(n15653) );
  AOI21_X1 U16809 ( .B1(P2_ADDR_REG_1__SCAN_IN), .B2(n15683), .A(n15653), .ZN(
        n15664) );
  OAI211_X1 U16810 ( .C1(n15656), .C2(n15655), .A(n15718), .B(n15654), .ZN(
        n15663) );
  INV_X1 U16811 ( .A(n15657), .ZN(n15661) );
  OAI21_X1 U16812 ( .B1(n10546), .B2(n15659), .A(n15658), .ZN(n15660) );
  NAND3_X1 U16813 ( .A1(n15743), .A2(n15661), .A3(n15660), .ZN(n15662) );
  NAND3_X1 U16814 ( .A1(n15664), .A2(n15663), .A3(n15662), .ZN(P2_U3215) );
  NAND2_X1 U16815 ( .A1(n15683), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n15666) );
  OAI211_X1 U16816 ( .C1(n15724), .C2(n15667), .A(n15666), .B(n15665), .ZN(
        n15668) );
  INV_X1 U16817 ( .A(n15668), .ZN(n15678) );
  OAI211_X1 U16818 ( .C1(n15671), .C2(n15670), .A(n15718), .B(n15669), .ZN(
        n15677) );
  AOI211_X1 U16819 ( .C1(n15674), .C2(n15673), .A(n15728), .B(n15672), .ZN(
        n15675) );
  INV_X1 U16820 ( .A(n15675), .ZN(n15676) );
  NAND3_X1 U16821 ( .A1(n15678), .A2(n15677), .A3(n15676), .ZN(P2_U3220) );
  AOI21_X1 U16822 ( .B1(n12248), .B2(n15680), .A(n15679), .ZN(n15682) );
  XOR2_X1 U16823 ( .A(n15682), .B(n15681), .Z(n15684) );
  AOI22_X1 U16824 ( .A1(n15684), .A2(n15718), .B1(n15683), .B2(
        P2_ADDR_REG_14__SCAN_IN), .ZN(n15693) );
  AOI211_X1 U16825 ( .C1(n15687), .C2(n15686), .A(n15728), .B(n15685), .ZN(
        n15688) );
  INV_X1 U16826 ( .A(n15688), .ZN(n15691) );
  NAND2_X1 U16827 ( .A1(n15741), .A2(n15689), .ZN(n15690) );
  NAND4_X1 U16828 ( .A1(n15693), .A2(n15692), .A3(n15691), .A4(n15690), .ZN(
        P2_U3228) );
  OAI22_X1 U16829 ( .A1(n15696), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n15695), 
        .B2(n15694), .ZN(n15699) );
  INV_X1 U16830 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n15697) );
  XNOR2_X1 U16831 ( .A(n7415), .B(n15697), .ZN(n15698) );
  XNOR2_X1 U16832 ( .A(n15699), .B(n15698), .ZN(n15700) );
  NAND2_X1 U16833 ( .A1(n15700), .A2(n15718), .ZN(n15710) );
  INV_X1 U16834 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n15704) );
  INV_X1 U16835 ( .A(n15701), .ZN(n15703) );
  OAI22_X1 U16836 ( .A1(n15705), .A2(n15704), .B1(n15703), .B2(n15702), .ZN(
        n15707) );
  XNOR2_X1 U16837 ( .A(n7415), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n15706) );
  XNOR2_X1 U16838 ( .A(n15707), .B(n15706), .ZN(n15708) );
  NAND2_X1 U16839 ( .A1(n15708), .A2(n15743), .ZN(n15709) );
  OAI211_X1 U16840 ( .C1(n15724), .C2(n15711), .A(n15710), .B(n15709), .ZN(
        n15712) );
  INV_X1 U16841 ( .A(n15712), .ZN(n15714) );
  OAI211_X1 U16842 ( .C1(n8393), .C2(n15749), .A(n15714), .B(n15713), .ZN(
        P2_U3233) );
  INV_X1 U16843 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n15897) );
  INV_X1 U16844 ( .A(n15715), .ZN(n15716) );
  AOI21_X1 U16845 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n15717), .A(n15716), 
        .ZN(n15720) );
  OAI211_X1 U16846 ( .C1(n15721), .C2(n15720), .A(n15719), .B(n15718), .ZN(
        n15723) );
  OAI211_X1 U16847 ( .C1(n15725), .C2(n15724), .A(n15723), .B(n15722), .ZN(
        n15726) );
  INV_X1 U16848 ( .A(n15726), .ZN(n15733) );
  AOI211_X1 U16849 ( .C1(n15730), .C2(n15729), .A(n15728), .B(n15727), .ZN(
        n15731) );
  INV_X1 U16850 ( .A(n15731), .ZN(n15732) );
  OAI211_X1 U16851 ( .C1(n15749), .C2(n15897), .A(n15733), .B(n15732), .ZN(
        P2_U3227) );
  INV_X1 U16852 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n15872) );
  INV_X1 U16853 ( .A(n15734), .ZN(n15735) );
  AOI211_X1 U16854 ( .C1(n15738), .C2(n15737), .A(n15736), .B(n15735), .ZN(
        n15739) );
  AOI211_X1 U16855 ( .C1(n15742), .C2(n15741), .A(n15740), .B(n15739), .ZN(
        n15748) );
  OAI211_X1 U16856 ( .C1(n15746), .C2(n15745), .A(n15744), .B(n15743), .ZN(
        n15747) );
  OAI211_X1 U16857 ( .C1(n15749), .C2(n15872), .A(n15748), .B(n15747), .ZN(
        P2_U3224) );
  NOR2_X1 U16858 ( .A1(n15750), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n15754) );
  NOR2_X1 U16859 ( .A1(n15752), .A2(n15751), .ZN(n15753) );
  MUX2_X1 U16860 ( .A(n15754), .B(n15753), .S(P1_IR_REG_0__SCAN_IN), .Z(n15755) );
  OR2_X1 U16861 ( .A1(n15756), .A2(n15755), .ZN(n15760) );
  AOI22_X1 U16862 ( .A1(n15757), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n15758) );
  OAI21_X1 U16863 ( .B1(n15760), .B2(n15759), .A(n15758), .ZN(P1_U3243) );
  OAI21_X1 U16864 ( .B1(n15762), .B2(n16340), .A(n15761), .ZN(n15770) );
  AOI21_X1 U16865 ( .B1(n15764), .B2(P1_REG2_REG_15__SCAN_IN), .A(n15763), 
        .ZN(n15768) );
  OAI22_X1 U16866 ( .A1(n15768), .A2(n15767), .B1(n15766), .B2(n15765), .ZN(
        n15769) );
  AOI21_X1 U16867 ( .B1(n15770), .B2(n15776), .A(n15769), .ZN(n15771) );
  NAND2_X1 U16868 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n16326)
         );
  OAI211_X1 U16869 ( .C1(n15922), .C2(n15784), .A(n15771), .B(n16326), .ZN(
        P1_U3258) );
  INV_X1 U16870 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n15785) );
  OAI21_X1 U16871 ( .B1(n15774), .B2(n15773), .A(n15772), .ZN(n15781) );
  XNOR2_X1 U16872 ( .A(n15775), .B(n16258), .ZN(n15777) );
  AOI222_X1 U16873 ( .A1(n15781), .A2(n15780), .B1(n15779), .B2(n15778), .C1(
        n15777), .C2(n15776), .ZN(n15783) );
  OAI211_X1 U16874 ( .C1(n15785), .C2(n15784), .A(n15783), .B(n15782), .ZN(
        P1_U3255) );
  AOI21_X1 U16875 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n15967), .A(n7576), .ZN(
        n15787) );
  INV_X1 U16876 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15786) );
  NOR2_X1 U16877 ( .A1(n15787), .A2(n15786), .ZN(n15958) );
  AOI21_X1 U16878 ( .B1(n15787), .B2(n15786), .A(n15958), .ZN(SUB_1596_U53) );
  NOR2_X1 U16879 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n15788), .ZN(n15789) );
  XNOR2_X1 U16880 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n15797), .ZN(n15800) );
  NAND2_X1 U16881 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n15791), .ZN(n15793) );
  NAND2_X1 U16882 ( .A1(n15959), .A2(n15958), .ZN(n15792) );
  NAND2_X1 U16883 ( .A1(n15793), .A2(n15792), .ZN(n15801) );
  NOR2_X1 U16884 ( .A1(n15801), .A2(n15800), .ZN(n15802) );
  AOI21_X1 U16885 ( .B1(n15800), .B2(n15801), .A(n15802), .ZN(n15794) );
  INV_X1 U16886 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n15804) );
  XNOR2_X1 U16887 ( .A(n15794), .B(n15804), .ZN(SUB_1596_U61) );
  NOR2_X1 U16888 ( .A1(n15796), .A2(n15795), .ZN(n15799) );
  XNOR2_X1 U16889 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n15805), .ZN(n15808) );
  NAND2_X1 U16890 ( .A1(n15801), .A2(n15800), .ZN(n15803) );
  AOI21_X1 U16891 ( .B1(n15804), .B2(n15803), .A(n15802), .ZN(n15809) );
  XNOR2_X1 U16892 ( .A(n15808), .B(n15809), .ZN(n15810) );
  XNOR2_X1 U16893 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15810), .ZN(SUB_1596_U60)
         );
  NOR2_X1 U16894 ( .A1(n15809), .A2(n15808), .ZN(n15812) );
  NOR2_X1 U16895 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(n15810), .ZN(n15811) );
  NOR2_X1 U16896 ( .A1(n15812), .A2(n15811), .ZN(n15817) );
  XOR2_X1 U16897 ( .A(n15818), .B(n15817), .Z(SUB_1596_U59) );
  NOR2_X1 U16898 ( .A1(n15813), .A2(n10860), .ZN(n15815) );
  INV_X1 U16899 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n15816) );
  INV_X1 U16900 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n15821) );
  AOI22_X1 U16901 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .B1(n15816), .B2(n15821), .ZN(n15822) );
  XNOR2_X1 U16902 ( .A(n15823), .B(n15822), .ZN(n15828) );
  NAND2_X1 U16903 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n15819), .ZN(n15820) );
  XOR2_X1 U16904 ( .A(n15830), .B(P2_ADDR_REG_5__SCAN_IN), .Z(SUB_1596_U58) );
  NOR2_X1 U16905 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n15821), .ZN(n15825) );
  NOR2_X1 U16906 ( .A1(n15823), .A2(n15822), .ZN(n15824) );
  NAND2_X1 U16907 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n15989), .ZN(n15826) );
  OAI21_X1 U16908 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(n15989), .A(n15826), .ZN(
        n15827) );
  XOR2_X1 U16909 ( .A(n15835), .B(n15827), .Z(n15831) );
  AND2_X1 U16910 ( .A1(n15832), .A2(n15831), .ZN(n15956) );
  NOR2_X1 U16911 ( .A1(n15955), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n15833) );
  INV_X1 U16912 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n15841) );
  OR2_X1 U16913 ( .A1(n15989), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n15834) );
  XOR2_X1 U16914 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n15840), .Z(n15842) );
  XNOR2_X1 U16915 ( .A(n15841), .B(n15842), .ZN(n15837) );
  XOR2_X1 U16916 ( .A(n15838), .B(n15837), .Z(SUB_1596_U56) );
  NAND2_X1 U16917 ( .A1(n15836), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n15839) );
  NAND2_X1 U16918 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n15840), .ZN(n15844) );
  NAND2_X1 U16919 ( .A1(n15842), .A2(n15841), .ZN(n15843) );
  NAND2_X1 U16920 ( .A1(n15844), .A2(n15843), .ZN(n15851) );
  INV_X1 U16921 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n15854) );
  NAND2_X1 U16922 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n15854), .ZN(n15845) );
  OAI21_X1 U16923 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n15854), .A(n15845), .ZN(
        n15852) );
  XOR2_X1 U16924 ( .A(n15851), .B(n15852), .Z(n15848) );
  XOR2_X1 U16925 ( .A(n15846), .B(P2_ADDR_REG_8__SCAN_IN), .Z(SUB_1596_U55) );
  NAND2_X1 U16926 ( .A1(n15846), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n15850) );
  NAND2_X1 U16927 ( .A1(n15848), .A2(n15847), .ZN(n15849) );
  NOR2_X1 U16928 ( .A1(n15852), .A2(n15851), .ZN(n15853) );
  INV_X1 U16929 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n16028) );
  NAND2_X1 U16930 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n16028), .ZN(n15855) );
  OAI21_X1 U16931 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n16028), .A(n15855), .ZN(
        n15857) );
  XOR2_X1 U16932 ( .A(n15858), .B(n15857), .Z(n15861) );
  NAND2_X1 U16933 ( .A1(n15861), .A2(n15860), .ZN(n15862) );
  OAI21_X1 U16934 ( .B1(n15860), .B2(n15861), .A(n15862), .ZN(n15856) );
  XNOR2_X1 U16935 ( .A(n15856), .B(P2_ADDR_REG_9__SCAN_IN), .ZN(SUB_1596_U54)
         );
  NOR2_X1 U16936 ( .A1(n15858), .A2(n15857), .ZN(n15859) );
  XNOR2_X1 U16937 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n15865) );
  XNOR2_X1 U16938 ( .A(n15866), .B(n15865), .ZN(n15870) );
  OAI21_X1 U16939 ( .B1(n15870), .B2(n15869), .A(n15871), .ZN(n15864) );
  XNOR2_X1 U16940 ( .A(n15864), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(SUB_1596_U70)
         );
  INV_X1 U16941 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n15877) );
  XNOR2_X1 U16942 ( .A(n15877), .B(P1_ADDR_REG_11__SCAN_IN), .ZN(n15875) );
  NAND2_X1 U16943 ( .A1(n15866), .A2(n15865), .ZN(n15867) );
  XOR2_X1 U16944 ( .A(n15875), .B(n15874), .Z(n15879) );
  AOI21_X1 U16945 ( .B1(n15879), .B2(n15878), .A(n15880), .ZN(n15873) );
  XNOR2_X1 U16946 ( .A(n15873), .B(n15881), .ZN(SUB_1596_U69) );
  NOR2_X1 U16947 ( .A1(n15875), .A2(n15874), .ZN(n15876) );
  XNOR2_X1 U16948 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n15887) );
  XNOR2_X1 U16949 ( .A(n15888), .B(n15887), .ZN(n15882) );
  XNOR2_X1 U16950 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n15884), .ZN(SUB_1596_U68)
         );
  NOR2_X1 U16951 ( .A1(n15883), .A2(n15882), .ZN(n15886) );
  XNOR2_X1 U16952 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n15891) );
  NAND2_X1 U16953 ( .A1(n15888), .A2(n15887), .ZN(n15889) );
  XNOR2_X1 U16954 ( .A(n15891), .B(n15900), .ZN(n15894) );
  AOI21_X1 U16955 ( .B1(n15893), .B2(n15894), .A(n15895), .ZN(n15892) );
  XNOR2_X1 U16956 ( .A(n15892), .B(n15897), .ZN(SUB_1596_U67) );
  NAND2_X1 U16957 ( .A1(n15894), .A2(n15893), .ZN(n15896) );
  INV_X1 U16958 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n15901) );
  INV_X1 U16959 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n15898) );
  NAND2_X1 U16960 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n15898), .ZN(n15899) );
  AOI22_X1 U16961 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n15901), .B1(n15900), 
        .B2(n15899), .ZN(n15905) );
  INV_X1 U16962 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n15902) );
  INV_X1 U16963 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n15907) );
  XOR2_X1 U16964 ( .A(n15902), .B(n15907), .Z(n15904) );
  XNOR2_X1 U16965 ( .A(n15905), .B(n15904), .ZN(n15909) );
  AOI21_X1 U16966 ( .B1(n15910), .B2(n15909), .A(n15911), .ZN(n15903) );
  INV_X1 U16967 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n15913) );
  XNOR2_X1 U16968 ( .A(n15903), .B(n15913), .ZN(SUB_1596_U66) );
  NOR2_X1 U16969 ( .A1(n15905), .A2(n15904), .ZN(n15906) );
  AOI21_X1 U16970 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n15907), .A(n15906), 
        .ZN(n15920) );
  INV_X1 U16971 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n15908) );
  XNOR2_X1 U16972 ( .A(n15908), .B(n15922), .ZN(n15919) );
  XOR2_X1 U16973 ( .A(n15920), .B(n15919), .Z(n15915) );
  NAND2_X1 U16974 ( .A1(n15910), .A2(n15909), .ZN(n15912) );
  NOR2_X1 U16975 ( .A1(n15918), .A2(n15917), .ZN(n15916) );
  XOR2_X1 U16976 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n15916), .Z(SUB_1596_U65)
         );
  NAND2_X1 U16977 ( .A1(n15920), .A2(n15919), .ZN(n15921) );
  XOR2_X1 U16978 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n15929), .Z(n15930) );
  XOR2_X1 U16979 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n15930), .Z(n15924) );
  NOR2_X1 U16980 ( .A1(n15928), .A2(n15926), .ZN(n15925) );
  XOR2_X1 U16981 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n15925), .Z(SUB_1596_U64)
         );
  NOR2_X1 U16982 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n15929), .ZN(n15932) );
  XNOR2_X1 U16983 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n15937), .ZN(n15938) );
  XOR2_X1 U16984 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n15938), .Z(n15933) );
  XOR2_X1 U16985 ( .A(n15933), .B(P2_ADDR_REG_17__SCAN_IN), .Z(n15934) );
  XOR2_X1 U16986 ( .A(n15935), .B(n15934), .Z(SUB_1596_U63) );
  NAND2_X1 U16987 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n15933), .ZN(n15936) );
  NOR2_X1 U16988 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n15937), .ZN(n15941) );
  NOR2_X1 U16989 ( .A1(n15939), .A2(n15938), .ZN(n15940) );
  NOR2_X1 U16990 ( .A1(n15941), .A2(n15940), .ZN(n15947) );
  XNOR2_X1 U16991 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n15948) );
  XOR2_X1 U16992 ( .A(n15947), .B(n15948), .Z(n15944) );
  XOR2_X1 U16993 ( .A(n15942), .B(P2_ADDR_REG_18__SCAN_IN), .Z(SUB_1596_U62)
         );
  NAND2_X1 U16994 ( .A1(n15942), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n15946) );
  NAND2_X1 U16995 ( .A1(n15944), .A2(n15943), .ZN(n15945) );
  NAND2_X1 U16996 ( .A1(n15946), .A2(n15945), .ZN(n15954) );
  NAND2_X1 U16997 ( .A1(n15948), .A2(n15947), .ZN(n15949) );
  OAI21_X1 U16998 ( .B1(n15214), .B2(P3_ADDR_REG_18__SCAN_IN), .A(n15949), 
        .ZN(n15952) );
  XNOR2_X1 U16999 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n15950) );
  XNOR2_X1 U17000 ( .A(n15950), .B(n7637), .ZN(n15951) );
  XNOR2_X1 U17001 ( .A(n15952), .B(n15951), .ZN(n15953) );
  XNOR2_X1 U17002 ( .A(n15954), .B(n15953), .ZN(SUB_1596_U4) );
  NOR2_X1 U17003 ( .A1(n15956), .A2(n15955), .ZN(n15957) );
  XOR2_X1 U17004 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n15957), .Z(SUB_1596_U57) );
  XOR2_X1 U17005 ( .A(n15959), .B(n15958), .Z(SUB_1596_U5) );
  NAND3_X1 U17006 ( .A1(n16013), .A2(n16009), .A3(n15960), .ZN(n15964) );
  OAI21_X1 U17007 ( .B1(P3_IR_REG_0__SCAN_IN), .B2(n15962), .A(n15961), .ZN(
        n15963) );
  NAND2_X1 U17008 ( .A1(n15964), .A2(n15963), .ZN(n15966) );
  AOI22_X1 U17009 ( .A1(n16020), .A2(P3_IR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n15965) );
  OAI211_X1 U17010 ( .C1(n15967), .C2(n16027), .A(n15966), .B(n15965), .ZN(
        P3_U3182) );
  XNOR2_X1 U17011 ( .A(n15969), .B(n15968), .ZN(n15986) );
  AND3_X1 U17012 ( .A1(n15972), .A2(n15971), .A3(n15970), .ZN(n15974) );
  OAI21_X1 U17013 ( .B1(n15975), .B2(n15974), .A(n15973), .ZN(n15983) );
  AND3_X1 U17014 ( .A1(n15978), .A2(n15977), .A3(n15976), .ZN(n15980) );
  OAI21_X1 U17015 ( .B1(n15981), .B2(n15980), .A(n15979), .ZN(n15982) );
  OAI211_X1 U17016 ( .C1(n15997), .C2(n15984), .A(n15983), .B(n15982), .ZN(
        n15985) );
  AOI21_X1 U17017 ( .B1(n15986), .B2(n16017), .A(n15985), .ZN(n15988) );
  OAI211_X1 U17018 ( .C1(n15989), .C2(n16027), .A(n15988), .B(n15987), .ZN(
        P3_U3188) );
  INV_X1 U17019 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n16006) );
  XNOR2_X1 U17020 ( .A(n15991), .B(n15990), .ZN(n16002) );
  AOI21_X1 U17021 ( .B1(n9381), .B2(n15993), .A(n15992), .ZN(n15994) );
  NOR2_X1 U17022 ( .A1(n15994), .A2(n16009), .ZN(n16001) );
  AOI21_X1 U17023 ( .B1(n9378), .B2(n15996), .A(n15995), .ZN(n15999) );
  OAI22_X1 U17024 ( .A1(n15999), .A2(n16013), .B1(n15998), .B2(n15997), .ZN(
        n16000) );
  AOI211_X1 U17025 ( .C1(n16017), .C2(n16002), .A(n16001), .B(n16000), .ZN(
        n16005) );
  INV_X1 U17026 ( .A(n16003), .ZN(n16004) );
  OAI211_X1 U17027 ( .C1(n16006), .C2(n16027), .A(n16005), .B(n16004), .ZN(
        P3_U3189) );
  AOI21_X1 U17028 ( .B1(n9408), .B2(n16008), .A(n16007), .ZN(n16010) );
  OR2_X1 U17029 ( .A1(n16010), .A2(n16009), .ZN(n16024) );
  AOI21_X1 U17030 ( .B1(n9405), .B2(n16012), .A(n16011), .ZN(n16014) );
  OR2_X1 U17031 ( .A1(n16014), .A2(n16013), .ZN(n16023) );
  XNOR2_X1 U17032 ( .A(n16016), .B(n16015), .ZN(n16018) );
  NAND2_X1 U17033 ( .A1(n16018), .A2(n16017), .ZN(n16022) );
  NAND2_X1 U17034 ( .A1(n16020), .A2(n16019), .ZN(n16021) );
  AND4_X1 U17035 ( .A1(n16024), .A2(n16023), .A3(n16022), .A4(n16021), .ZN(
        n16026) );
  OAI211_X1 U17036 ( .C1(n16028), .C2(n16027), .A(n16026), .B(n16025), .ZN(
        P3_U3191) );
  INV_X1 U17037 ( .A(P3_RD_REG_SCAN_IN), .ZN(n16029) );
  OAI221_X1 U17038 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .C1(n8391), .C2(n16030), .A(n16029), .ZN(U29) );
  OAI22_X1 U17039 ( .A1(n16033), .A2(n16135), .B1(n16032), .B2(n16031), .ZN(
        n16034) );
  NOR2_X1 U17040 ( .A1(n16035), .A2(n16034), .ZN(n16036) );
  AOI22_X1 U17041 ( .A1(n16341), .A2(n16036), .B1(n15751), .B2(n16339), .ZN(
        P1_U3528) );
  AOI22_X1 U17042 ( .A1(n16345), .A2(n16036), .B1(n8785), .B2(n16342), .ZN(
        P1_U3459) );
  AOI222_X1 U17043 ( .A1(n16042), .A2(n16041), .B1(n16040), .B2(n16039), .C1(
        n16038), .C2(n16037), .ZN(n16043) );
  OAI21_X1 U17044 ( .B1(n16045), .B2(n16044), .A(n16043), .ZN(P3_U3172) );
  INV_X1 U17045 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n16046) );
  AOI22_X1 U17046 ( .A1(n16242), .A2(n16047), .B1(n16046), .B2(n16239), .ZN(
        P3_U3393) );
  XNOR2_X1 U17047 ( .A(n16048), .B(n16050), .ZN(n16065) );
  NOR2_X1 U17048 ( .A1(n16049), .A2(n16231), .ZN(n16058) );
  XNOR2_X1 U17049 ( .A(n16051), .B(n16050), .ZN(n16052) );
  OAI222_X1 U17050 ( .A1(n16056), .A2(n16055), .B1(n16054), .B2(n7579), .C1(
        n16053), .C2(n16052), .ZN(n16063) );
  AOI211_X1 U17051 ( .C1(n16065), .C2(n16103), .A(n16058), .B(n16063), .ZN(
        n16057) );
  AOI22_X1 U17052 ( .A1(n16238), .A2(n16057), .B1(n10169), .B2(n9764), .ZN(
        P3_U3461) );
  AOI22_X1 U17053 ( .A1(n16242), .A2(n16057), .B1(n9303), .B2(n16239), .ZN(
        P3_U3396) );
  INV_X1 U17054 ( .A(n16058), .ZN(n16062) );
  OAI22_X1 U17055 ( .A1(n16062), .A2(n16061), .B1(n16060), .B2(n16059), .ZN(
        n16064) );
  AOI211_X1 U17056 ( .C1(n16065), .C2(n16088), .A(n16064), .B(n16063), .ZN(
        n16066) );
  AOI22_X1 U17057 ( .A1(n14341), .A2(n16067), .B1(n16066), .B2(n16100), .ZN(
        P3_U3231) );
  INV_X1 U17058 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n16068) );
  AOI22_X1 U17059 ( .A1(n16345), .A2(n16069), .B1(n16068), .B2(n16342), .ZN(
        P1_U3465) );
  INV_X1 U17060 ( .A(n16070), .ZN(n16071) );
  AOI21_X1 U17061 ( .B1(n16160), .B2(n16079), .A(n16071), .ZN(n16081) );
  NAND2_X1 U17062 ( .A1(n16073), .A2(n16072), .ZN(n16076) );
  AOI22_X1 U17063 ( .A1(n16264), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n16262), 
        .B2(n10958), .ZN(n16075) );
  OAI211_X1 U17064 ( .C1(n16077), .C2(n16114), .A(n16076), .B(n16075), .ZN(
        n16078) );
  AOI21_X1 U17065 ( .B1(n16270), .B2(n16079), .A(n16078), .ZN(n16080) );
  OAI21_X1 U17066 ( .B1(n16275), .B2(n16081), .A(n16080), .ZN(P1_U3290) );
  OAI22_X1 U17067 ( .A1(n16082), .A2(n16198), .B1(n8053), .B2(n16333), .ZN(
        n16084) );
  AOI211_X1 U17068 ( .C1(n16337), .C2(n16085), .A(n16084), .B(n16083), .ZN(
        n16087) );
  AOI22_X1 U17069 ( .A1(n16341), .A2(n16087), .B1(n10607), .B2(n16339), .ZN(
        P1_U3532) );
  INV_X1 U17070 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n16086) );
  AOI22_X1 U17071 ( .A1(n16345), .A2(n16087), .B1(n16086), .B2(n16342), .ZN(
        P1_U3471) );
  INV_X1 U17072 ( .A(n16088), .ZN(n16092) );
  INV_X1 U17073 ( .A(n16089), .ZN(n16091) );
  OAI21_X1 U17074 ( .B1(n16092), .B2(n16091), .A(n16090), .ZN(n16098) );
  INV_X1 U17075 ( .A(n16093), .ZN(n16095) );
  AOI222_X1 U17076 ( .A1(n16098), .A2(n16100), .B1(n16097), .B2(n16096), .C1(
        n16095), .C2(n16094), .ZN(n16099) );
  OAI21_X1 U17077 ( .B1(n16100), .B2(n9344), .A(n16099), .ZN(P3_U3228) );
  AOI22_X1 U17078 ( .A1(n16104), .A2(n16103), .B1(n16102), .B2(n16101), .ZN(
        n16106) );
  AND2_X1 U17079 ( .A1(n16106), .A2(n16105), .ZN(n16108) );
  INV_X1 U17080 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n16107) );
  AOI22_X1 U17081 ( .A1(n16238), .A2(n16108), .B1(n16107), .B2(n9764), .ZN(
        P3_U3465) );
  AOI22_X1 U17082 ( .A1(n16242), .A2(n16108), .B1(n9359), .B2(n16239), .ZN(
        P3_U3408) );
  NOR2_X1 U17083 ( .A1(n16110), .A2(n16109), .ZN(n16111) );
  AOI21_X1 U17084 ( .B1(n16264), .B2(P1_REG2_REG_6__SCAN_IN), .A(n16111), .ZN(
        n16112) );
  OAI21_X1 U17085 ( .B1(n16114), .B2(n16113), .A(n16112), .ZN(n16115) );
  INV_X1 U17086 ( .A(n16115), .ZN(n16119) );
  AOI22_X1 U17087 ( .A1(n16117), .A2(n16270), .B1(n16269), .B2(n16116), .ZN(
        n16118) );
  OAI211_X1 U17088 ( .C1(n16275), .C2(n16120), .A(n16119), .B(n16118), .ZN(
        P1_U3287) );
  AND2_X1 U17089 ( .A1(n16121), .A2(n16310), .ZN(n16126) );
  INV_X1 U17090 ( .A(n16122), .ZN(n16123) );
  OAI22_X1 U17091 ( .A1(n16124), .A2(n10363), .B1(n16123), .B2(n16307), .ZN(
        n16125) );
  NOR3_X1 U17092 ( .A1(n16127), .A2(n16126), .A3(n16125), .ZN(n16130) );
  AOI22_X1 U17093 ( .A1(n16293), .A2(n16130), .B1(n16128), .B2(n16314), .ZN(
        P2_U3505) );
  INV_X1 U17094 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n16129) );
  AOI22_X1 U17095 ( .A1(n7419), .A2(n16130), .B1(n16129), .B2(n16315), .ZN(
        P2_U3448) );
  INV_X1 U17096 ( .A(n16136), .ZN(n16138) );
  AOI21_X1 U17097 ( .B1(n16278), .B2(n16132), .A(n16131), .ZN(n16133) );
  OAI211_X1 U17098 ( .C1(n16136), .C2(n16135), .A(n16134), .B(n16133), .ZN(
        n16137) );
  AOI21_X1 U17099 ( .B1(n16160), .B2(n16138), .A(n16137), .ZN(n16140) );
  AOI22_X1 U17100 ( .A1(n16341), .A2(n16140), .B1(n10682), .B2(n16339), .ZN(
        P1_U3535) );
  INV_X1 U17101 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n16139) );
  AOI22_X1 U17102 ( .A1(n16345), .A2(n16140), .B1(n16139), .B2(n16342), .ZN(
        P1_U3480) );
  OAI22_X1 U17103 ( .A1(n16142), .A2(n10363), .B1(n16141), .B2(n16307), .ZN(
        n16144) );
  AOI211_X1 U17104 ( .C1(n16145), .C2(n16310), .A(n16144), .B(n16143), .ZN(
        n16148) );
  AOI22_X1 U17105 ( .A1(n16293), .A2(n16148), .B1(n16146), .B2(n16314), .ZN(
        P2_U3506) );
  INV_X1 U17106 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n16147) );
  AOI22_X1 U17107 ( .A1(n7419), .A2(n16148), .B1(n16147), .B2(n16315), .ZN(
        P2_U3451) );
  NAND2_X1 U17108 ( .A1(n16150), .A2(n16149), .ZN(n16151) );
  INV_X1 U17109 ( .A(n16153), .ZN(n16159) );
  INV_X1 U17110 ( .A(n16154), .ZN(n16155) );
  AOI211_X1 U17111 ( .C1(n16157), .C2(n16156), .A(n16280), .B(n16155), .ZN(
        n16158) );
  AOI211_X1 U17112 ( .C1(n16160), .C2(n16178), .A(n16159), .B(n16158), .ZN(
        n16186) );
  INV_X1 U17113 ( .A(n16161), .ZN(n16171) );
  AOI21_X1 U17114 ( .B1(n16162), .B2(n16278), .A(n16171), .ZN(n16167) );
  OAI21_X1 U17115 ( .B1(n16163), .B2(n16175), .A(n16247), .ZN(n16164) );
  OR2_X1 U17116 ( .A1(n16165), .A2(n16164), .ZN(n16182) );
  NAND2_X1 U17117 ( .A1(n16178), .A2(n16257), .ZN(n16166) );
  AOI22_X1 U17118 ( .A1(n16341), .A2(n16169), .B1(n10757), .B2(n16339), .ZN(
        P1_U3536) );
  INV_X1 U17119 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n16168) );
  AOI22_X1 U17120 ( .A1(n16345), .A2(n16169), .B1(n16168), .B2(n16342), .ZN(
        P1_U3483) );
  INV_X1 U17121 ( .A(n16170), .ZN(n16177) );
  AOI21_X1 U17122 ( .B1(n16262), .B2(n16172), .A(n16171), .ZN(n16173) );
  OAI21_X1 U17123 ( .B1(n16175), .B2(n16174), .A(n16173), .ZN(n16176) );
  AOI21_X1 U17124 ( .B1(n16178), .B2(n16177), .A(n16176), .ZN(n16185) );
  OAI22_X1 U17125 ( .A1(n16182), .A2(n16181), .B1(n16180), .B2(n16179), .ZN(
        n16183) );
  INV_X1 U17126 ( .A(n16183), .ZN(n16184) );
  OAI221_X1 U17127 ( .B1(n16275), .B2(n16186), .C1(n16275), .C2(n16185), .A(
        n16184), .ZN(P1_U3285) );
  AND3_X1 U17128 ( .A1(n16188), .A2(n16187), .A3(n16310), .ZN(n16192) );
  OAI22_X1 U17129 ( .A1(n16190), .A2(n10363), .B1(n16189), .B2(n16307), .ZN(
        n16191) );
  NOR3_X1 U17130 ( .A1(n16193), .A2(n16192), .A3(n16191), .ZN(n16196) );
  AOI22_X1 U17131 ( .A1(n16293), .A2(n16196), .B1(n16194), .B2(n16314), .ZN(
        P2_U3507) );
  INV_X1 U17132 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n16195) );
  AOI22_X1 U17133 ( .A1(n7419), .A2(n16196), .B1(n16195), .B2(n16315), .ZN(
        P2_U3454) );
  OAI22_X1 U17134 ( .A1(n16199), .A2(n16198), .B1(n16197), .B2(n16333), .ZN(
        n16201) );
  AOI211_X1 U17135 ( .C1(n16257), .C2(n16202), .A(n16201), .B(n16200), .ZN(
        n16204) );
  AOI22_X1 U17136 ( .A1(n16341), .A2(n16204), .B1(n10754), .B2(n16339), .ZN(
        P1_U3537) );
  INV_X1 U17137 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n16203) );
  AOI22_X1 U17138 ( .A1(n16345), .A2(n16204), .B1(n16203), .B2(n16342), .ZN(
        P1_U3486) );
  NAND2_X1 U17139 ( .A1(n16205), .A2(n13663), .ZN(n16207) );
  OAI211_X1 U17140 ( .C1(n16208), .C2(n16307), .A(n16207), .B(n16206), .ZN(
        n16209) );
  NOR2_X1 U17141 ( .A1(n16210), .A2(n16209), .ZN(n16213) );
  AOI22_X1 U17142 ( .A1(n16293), .A2(n16213), .B1(n16211), .B2(n16314), .ZN(
        P2_U3508) );
  INV_X1 U17143 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n16212) );
  AOI22_X1 U17144 ( .A1(n7419), .A2(n16213), .B1(n16212), .B2(n16315), .ZN(
        P2_U3457) );
  OAI211_X1 U17145 ( .C1(n16216), .C2(n16333), .A(n16215), .B(n16214), .ZN(
        n16217) );
  AOI21_X1 U17146 ( .B1(n16218), .B2(n16337), .A(n16217), .ZN(n16220) );
  AOI22_X1 U17147 ( .A1(n16341), .A2(n16220), .B1(n11173), .B2(n16339), .ZN(
        P1_U3538) );
  INV_X1 U17148 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n16219) );
  AOI22_X1 U17149 ( .A1(n16345), .A2(n16220), .B1(n16219), .B2(n16342), .ZN(
        P1_U3489) );
  MUX2_X1 U17150 ( .A(P3_REG0_REG_11__SCAN_IN), .B(n16221), .S(n16242), .Z(
        P3_U3423) );
  OAI211_X1 U17151 ( .C1(n16224), .C2(n16333), .A(n16223), .B(n16222), .ZN(
        n16227) );
  NOR2_X1 U17152 ( .A1(n16225), .A2(n16299), .ZN(n16226) );
  AOI211_X1 U17153 ( .C1(n16228), .C2(n16330), .A(n16227), .B(n16226), .ZN(
        n16230) );
  AOI22_X1 U17154 ( .A1(n16341), .A2(n16230), .B1(n7716), .B2(n16339), .ZN(
        P1_U3539) );
  INV_X1 U17155 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n16229) );
  AOI22_X1 U17156 ( .A1(n16345), .A2(n16230), .B1(n16229), .B2(n16342), .ZN(
        P1_U3492) );
  NOR2_X1 U17157 ( .A1(n16232), .A2(n16231), .ZN(n16234) );
  AOI211_X1 U17158 ( .C1(n16236), .C2(n16235), .A(n16234), .B(n16233), .ZN(
        n16241) );
  AOI22_X1 U17159 ( .A1(n16238), .A2(n16241), .B1(n16237), .B2(n9764), .ZN(
        P3_U3471) );
  INV_X1 U17160 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n16240) );
  AOI22_X1 U17161 ( .A1(n16242), .A2(n16241), .B1(n16240), .B2(n16239), .ZN(
        P3_U3426) );
  AOI21_X1 U17162 ( .B1(n16251), .B2(n16244), .A(n16243), .ZN(n16255) );
  INV_X1 U17163 ( .A(n16255), .ZN(n16271) );
  INV_X1 U17164 ( .A(n16245), .ZN(n16248) );
  OAI211_X1 U17165 ( .C1(n16248), .C2(n16249), .A(n16247), .B(n16246), .ZN(
        n16267) );
  OAI21_X1 U17166 ( .B1(n16249), .B2(n16333), .A(n16267), .ZN(n16256) );
  OAI211_X1 U17167 ( .C1(n7562), .C2(n16251), .A(n16250), .B(n16330), .ZN(
        n16252) );
  OAI211_X1 U17168 ( .C1(n16255), .C2(n16254), .A(n16253), .B(n16252), .ZN(
        n16261) );
  AOI211_X1 U17169 ( .C1(n16257), .C2(n16271), .A(n16256), .B(n16261), .ZN(
        n16260) );
  AOI22_X1 U17170 ( .A1(n16341), .A2(n16260), .B1(n16258), .B2(n16339), .ZN(
        P1_U3540) );
  INV_X1 U17171 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n16259) );
  AOI22_X1 U17172 ( .A1(n16345), .A2(n16260), .B1(n16259), .B2(n16342), .ZN(
        P1_U3495) );
  INV_X1 U17173 ( .A(n16261), .ZN(n16274) );
  AOI222_X1 U17174 ( .A1(n16266), .A2(n16265), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n16264), .C1(n16263), .C2(n16262), .ZN(n16273) );
  INV_X1 U17175 ( .A(n16267), .ZN(n16268) );
  AOI22_X1 U17176 ( .A1(n16271), .A2(n16270), .B1(n16269), .B2(n16268), .ZN(
        n16272) );
  OAI211_X1 U17177 ( .C1(n16275), .C2(n16274), .A(n16273), .B(n16272), .ZN(
        P1_U3281) );
  AOI21_X1 U17178 ( .B1(n16278), .B2(n16277), .A(n16276), .ZN(n16279) );
  OAI21_X1 U17179 ( .B1(n16281), .B2(n16280), .A(n16279), .ZN(n16282) );
  AOI21_X1 U17180 ( .B1(n16283), .B2(n16337), .A(n16282), .ZN(n16286) );
  AOI22_X1 U17181 ( .A1(n16341), .A2(n16286), .B1(n16284), .B2(n16339), .ZN(
        P1_U3541) );
  INV_X1 U17182 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n16285) );
  AOI22_X1 U17183 ( .A1(n16345), .A2(n16286), .B1(n16285), .B2(n16342), .ZN(
        P1_U3498) );
  OAI21_X1 U17184 ( .B1(n16288), .B2(n16307), .A(n16287), .ZN(n16290) );
  AOI211_X1 U17185 ( .C1(n13663), .C2(n16291), .A(n16290), .B(n16289), .ZN(
        n16295) );
  AOI22_X1 U17186 ( .A1(n16293), .A2(n16295), .B1(n16292), .B2(n16314), .ZN(
        P2_U3512) );
  INV_X1 U17187 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n16294) );
  AOI22_X1 U17188 ( .A1(n7419), .A2(n16295), .B1(n16294), .B2(n16315), .ZN(
        P2_U3469) );
  OAI211_X1 U17189 ( .C1(n16298), .C2(n16333), .A(n16297), .B(n16296), .ZN(
        n16303) );
  NOR3_X1 U17190 ( .A1(n16301), .A2(n16300), .A3(n16299), .ZN(n16302) );
  AOI211_X1 U17191 ( .C1(n16330), .C2(n16304), .A(n16303), .B(n16302), .ZN(
        n16306) );
  AOI22_X1 U17192 ( .A1(n16341), .A2(n16306), .B1(n12082), .B2(n16339), .ZN(
        P1_U3542) );
  INV_X1 U17193 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n16305) );
  AOI22_X1 U17194 ( .A1(n16345), .A2(n16306), .B1(n16305), .B2(n16342), .ZN(
        P1_U3501) );
  OAI22_X1 U17195 ( .A1(n16308), .A2(n10363), .B1(n7975), .B2(n16307), .ZN(
        n16309) );
  AOI21_X1 U17196 ( .B1(n16311), .B2(n16310), .A(n16309), .ZN(n16313) );
  AND2_X1 U17197 ( .A1(n16313), .A2(n16312), .ZN(n16317) );
  AOI22_X1 U17198 ( .A1(n16293), .A2(n16317), .B1(n12240), .B2(n16314), .ZN(
        P2_U3513) );
  INV_X1 U17199 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n16316) );
  AOI22_X1 U17200 ( .A1(n7419), .A2(n16317), .B1(n16316), .B2(n16315), .ZN(
        P2_U3472) );
  OAI21_X1 U17201 ( .B1(n16320), .B2(n16319), .A(n16318), .ZN(n16325) );
  AOI22_X1 U17202 ( .A1(n16351), .A2(n16322), .B1(n16349), .B2(n16321), .ZN(
        n16323) );
  OAI21_X1 U17203 ( .B1(n16334), .B2(n16353), .A(n16323), .ZN(n16324) );
  AOI21_X1 U17204 ( .B1(n16325), .B2(n16356), .A(n16324), .ZN(n16327) );
  OAI211_X1 U17205 ( .C1(n16361), .C2(n16328), .A(n16327), .B(n16326), .ZN(
        P1_U3241) );
  AND3_X1 U17206 ( .A1(n13356), .A2(n16330), .A3(n16329), .ZN(n16336) );
  OAI211_X1 U17207 ( .C1(n16334), .C2(n16333), .A(n16332), .B(n16331), .ZN(
        n16335) );
  AOI211_X1 U17208 ( .C1(n16338), .C2(n16337), .A(n16336), .B(n16335), .ZN(
        n16344) );
  AOI22_X1 U17209 ( .A1(n16341), .A2(n16344), .B1(n16340), .B2(n16339), .ZN(
        P1_U3543) );
  INV_X1 U17210 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n16343) );
  AOI22_X1 U17211 ( .A1(n16345), .A2(n16344), .B1(n16343), .B2(n16342), .ZN(
        P1_U3504) );
  XNOR2_X1 U17212 ( .A(n16347), .B(n16346), .ZN(n16357) );
  AOI22_X1 U17213 ( .A1(n16351), .A2(n16350), .B1(n16349), .B2(n16348), .ZN(
        n16352) );
  OAI21_X1 U17214 ( .B1(n16354), .B2(n16353), .A(n16352), .ZN(n16355) );
  AOI21_X1 U17215 ( .B1(n16357), .B2(n16356), .A(n16355), .ZN(n16359) );
  OAI211_X1 U17216 ( .C1(n16361), .C2(n16360), .A(n16359), .B(n16358), .ZN(
        P1_U3226) );
  AOI21_X1 U17217 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n16362) );
  OAI21_X1 U17218 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(n16362), 
        .ZN(U28) );
  AND3_X1 U7518 ( .A1(n8962), .A2(n8961), .A3(n8960), .ZN(n8964) );
  NAND2_X1 U7549 ( .A1(n11131), .A2(n10432), .ZN(n10312) );
  CLKBUF_X1 U7609 ( .A(n9537), .Z(n9551) );
  CLKBUF_X1 U7754 ( .A(n10131), .Z(n7594) );
  CLKBUF_X1 U7862 ( .A(n10662), .Z(n7415) );
  NAND2_X1 U7873 ( .A1(n10048), .A2(n10047), .ZN(n14176) );
  NAND2_X1 U7881 ( .A1(n14469), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9272) );
  CLKBUF_X3 U7938 ( .A(n13680), .Z(n7432) );
  CLKBUF_X1 U8850 ( .A(n15020), .Z(n7629) );
  CLKBUF_X1 U9631 ( .A(n11260), .Z(n7430) );
endmodule

