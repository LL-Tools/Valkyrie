

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398;

  INV_X4 U4775 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NAND2_X1 U4776 ( .A1(n9384), .A2(n9287), .ZN(n9557) );
  INV_X2 U4778 ( .A(n7313), .ZN(n7748) );
  NAND2_X1 U4779 ( .A1(n8277), .A2(n8078), .ZN(n6648) );
  XNOR2_X1 U4780 ( .A(n5508), .B(n5507), .ZN(n6992) );
  INV_X1 U4781 ( .A(n6998), .ZN(n6946) );
  NAND2_X1 U4782 ( .A1(n5265), .A2(n5264), .ZN(n5858) );
  NAND3_X2 U4783 ( .A1(n4711), .A2(n5890), .A3(n4710), .ZN(n6943) );
  INV_X1 U4784 ( .A(n4271), .ZN(n6950) );
  INV_X1 U4785 ( .A(n6640), .ZN(n6742) );
  INV_X1 U4786 ( .A(n6097), .ZN(n6073) );
  AND2_X1 U4787 ( .A1(n5393), .A2(n5394), .ZN(n5422) );
  CLKBUF_X3 U4788 ( .A(n4271), .Z(n5690) );
  INV_X1 U4789 ( .A(n6354), .ZN(n6599) );
  INV_X1 U4790 ( .A(n6319), .ZN(n6484) );
  INV_X1 U4791 ( .A(n7719), .ZN(n6917) );
  AND2_X1 U4792 ( .A1(n4745), .A2(n4744), .ZN(n6845) );
  OR2_X1 U4793 ( .A1(n5858), .A2(n7458), .ZN(n7296) );
  NAND2_X1 U4794 ( .A1(n4464), .A2(n4939), .ZN(n5508) );
  INV_X1 U4795 ( .A(n10272), .ZN(n7652) );
  INV_X1 U4797 ( .A(n7569), .ZN(n8312) );
  AND2_X1 U4798 ( .A1(n5773), .A2(n5772), .ZN(n9566) );
  AND2_X1 U4799 ( .A1(n4315), .A2(n5290), .ZN(n10219) );
  INV_X1 U4800 ( .A(n7344), .ZN(n7723) );
  OAI21_X1 U4801 ( .B1(n8050), .B2(n5097), .A(n9534), .ZN(n9813) );
  NAND2_X1 U4802 ( .A1(n8542), .A2(n5077), .ZN(n4270) );
  OR2_X1 U4804 ( .A1(n5392), .A2(SI_6_), .ZN(n5393) );
  OR2_X2 U4805 ( .A1(n8680), .A2(n8679), .ZN(n8682) );
  AOI21_X1 U4806 ( .B1(n6671), .B2(n5131), .A(n5130), .ZN(n5129) );
  NAND2_X2 U4807 ( .A1(n7436), .A2(n9307), .ZN(n5180) );
  NAND2_X2 U4808 ( .A1(n10078), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5185) );
  XNOR2_X2 U4809 ( .A(n5940), .B(n5938), .ZN(n7374) );
  OAI21_X2 U4810 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10357), .ZN(n10386) );
  BUF_X8 U4811 ( .A(n6947), .Z(n4271) );
  NAND2_X2 U4812 ( .A1(n4929), .A2(n4928), .ZN(n6947) );
  XNOR2_X1 U4813 ( .A(n4560), .B(n9557), .ZN(n9823) );
  NAND2_X1 U4814 ( .A1(n5857), .A2(n5856), .ZN(n9560) );
  XNOR2_X1 U4815 ( .A(n9580), .B(n4272), .ZN(n9832) );
  INV_X1 U4816 ( .A(n9588), .ZN(n4272) );
  NOR2_X2 U4817 ( .A1(n6736), .A2(n6737), .ZN(n8536) );
  OR2_X1 U4818 ( .A1(n9828), .A2(n9567), .ZN(n9230) );
  OAI21_X1 U4819 ( .B1(n7850), .B2(n4660), .A(n4657), .ZN(n8175) );
  NAND2_X1 U4820 ( .A1(n6556), .A2(n6555), .ZN(n8543) );
  OR3_X1 U4821 ( .A1(n5747), .A2(n5746), .A3(n9034), .ZN(n5766) );
  NAND2_X1 U4822 ( .A1(n6421), .A2(n6420), .ZN(n8946) );
  CLKBUF_X2 U4823 ( .A(n6083), .Z(n6093) );
  INV_X2 U4824 ( .A(n6083), .ZN(n5929) );
  CLKBUF_X2 U4825 ( .A(n5935), .Z(n6083) );
  INV_X2 U4826 ( .A(n7522), .ZN(n6059) );
  INV_X2 U4827 ( .A(n5902), .ZN(n6056) );
  INV_X2 U4828 ( .A(n9267), .ZN(n9242) );
  INV_X1 U4829 ( .A(n7087), .ZN(n7290) );
  AND3_X1 U4830 ( .A1(n6331), .A2(n6330), .A3(n6329), .ZN(n7569) );
  INV_X1 U4831 ( .A(n6354), .ZN(n6341) );
  AND2_X2 U4832 ( .A1(n5184), .A2(n4786), .ZN(n5311) );
  NAND2_X1 U4833 ( .A1(n6998), .A2(n6950), .ZN(n9255) );
  NAND2_X2 U4834 ( .A1(n7014), .A2(n5815), .ZN(n6998) );
  OR2_X1 U4835 ( .A1(n5411), .A2(n7791), .ZN(n5437) );
  NAND3_X1 U4836 ( .A1(n5809), .A2(n5238), .A3(n5028), .ZN(n4694) );
  NOR2_X1 U4837 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5240) );
  OAI21_X1 U4838 ( .B1(n9033), .B2(n5032), .A(n4299), .ZN(n6108) );
  NAND2_X1 U4839 ( .A1(n6085), .A2(n9032), .ZN(n9033) );
  AND2_X1 U4840 ( .A1(n5187), .A2(n5186), .ZN(n9831) );
  OR3_X1 U4841 ( .A1(n8999), .A2(n4691), .A3(n4689), .ZN(n4688) );
  OR2_X1 U4842 ( .A1(n8999), .A2(n4691), .ZN(n4686) );
  AND2_X1 U4843 ( .A1(n5047), .A2(n5046), .ZN(n8999) );
  AND2_X1 U4844 ( .A1(n5091), .A2(n5092), .ZN(n8050) );
  NAND2_X1 U4845 ( .A1(n5091), .A2(n4331), .ZN(n9534) );
  AND2_X1 U4846 ( .A1(n4479), .A2(n4808), .ZN(n9547) );
  NAND2_X1 U4847 ( .A1(n4644), .A2(n5164), .ZN(n8599) );
  NOR2_X1 U4848 ( .A1(n8056), .A2(n9259), .ZN(n9528) );
  NAND2_X1 U4849 ( .A1(n4276), .A2(n4540), .ZN(n9580) );
  NAND2_X1 U4850 ( .A1(n5854), .A2(n4542), .ZN(n4276) );
  NAND2_X1 U4851 ( .A1(n9675), .A2(n9293), .ZN(n9657) );
  OR2_X1 U4852 ( .A1(n8781), .A2(n7467), .ZN(n6749) );
  AOI21_X1 U4853 ( .B1(n9675), .B2(n5175), .A(n5173), .ZN(n9643) );
  NAND2_X1 U4854 ( .A1(n9641), .A2(n5852), .ZN(n5854) );
  AND2_X1 U4855 ( .A1(n6079), .A2(n9031), .ZN(n5050) );
  NAND2_X1 U4856 ( .A1(n9676), .A2(n9677), .ZN(n9675) );
  NAND2_X1 U4857 ( .A1(n4277), .A2(n5081), .ZN(n9666) );
  NAND2_X1 U4858 ( .A1(n4806), .A2(n9215), .ZN(n9676) );
  OAI21_X1 U4859 ( .B1(n5537), .B2(n4801), .A(n4799), .ZN(n4806) );
  NAND2_X1 U4860 ( .A1(n9671), .A2(n5083), .ZN(n4277) );
  NAND2_X1 U4861 ( .A1(n8038), .A2(n8042), .ZN(n6024) );
  XNOR2_X1 U4862 ( .A(n6282), .B(n5798), .ZN(n8965) );
  CLKBUF_X1 U4863 ( .A(n8260), .Z(n4725) );
  INV_X1 U4864 ( .A(n9549), .ZN(n9590) );
  NAND2_X1 U4865 ( .A1(n5797), .A2(n5796), .ZN(n6282) );
  AND2_X2 U4866 ( .A1(n9343), .A2(n9234), .ZN(n9596) );
  AND2_X1 U4867 ( .A1(n8537), .A2(n6732), .ZN(n8555) );
  OAI21_X1 U4868 ( .B1(n9744), .B2(n4553), .A(n4551), .ZN(n9671) );
  NAND2_X1 U4869 ( .A1(n8039), .A2(n8040), .ZN(n8038) );
  OR2_X1 U4870 ( .A1(n8802), .A2(n8368), .ZN(n8537) );
  NAND2_X1 U4871 ( .A1(n9792), .A2(n9793), .ZN(n9791) );
  AND2_X1 U4872 ( .A1(n5754), .A2(n5753), .ZN(n9549) );
  NAND2_X1 U4873 ( .A1(n5843), .A2(n5089), .ZN(n9744) );
  NAND2_X1 U4874 ( .A1(n5745), .A2(n5744), .ZN(n9826) );
  AND2_X2 U4875 ( .A1(n8651), .A2(n8922), .ZN(n8612) );
  NAND2_X2 U4876 ( .A1(n6545), .A2(n6544), .ZN(n8802) );
  XNOR2_X1 U4877 ( .A(n5762), .B(n5761), .ZN(n10090) );
  AND2_X1 U4878 ( .A1(n5748), .A2(n5766), .ZN(n9574) );
  OAI21_X1 U4879 ( .B1(n5739), .B2(n5738), .A(n5737), .ZN(n5757) );
  NAND2_X1 U4880 ( .A1(n4951), .A2(n4949), .ZN(n5762) );
  NAND2_X1 U4881 ( .A1(n5167), .A2(n9297), .ZN(n7913) );
  NAND2_X1 U4882 ( .A1(n5663), .A2(n5662), .ZN(n9991) );
  NAND2_X1 U4883 ( .A1(n6487), .A2(n6486), .ZN(n8834) );
  NAND2_X1 U4884 ( .A1(n5098), .A2(n4292), .ZN(n5840) );
  NAND2_X1 U4885 ( .A1(n7688), .A2(n4273), .ZN(n5098) );
  NAND2_X1 U4886 ( .A1(n7688), .A2(n5835), .ZN(n7859) );
  XNOR2_X1 U4887 ( .A(n5643), .B(n5642), .ZN(n7451) );
  NAND2_X1 U4888 ( .A1(n6465), .A2(n6464), .ZN(n8926) );
  NAND2_X1 U4889 ( .A1(n6930), .A2(n6923), .ZN(n8377) );
  NAND2_X1 U4890 ( .A1(n5601), .A2(n5600), .ZN(n10004) );
  NAND2_X1 U4891 ( .A1(n5586), .A2(n5585), .ZN(n10010) );
  NOR2_X1 U4892 ( .A1(n4275), .A2(n4274), .ZN(n4273) );
  XNOR2_X1 U4893 ( .A(n8938), .B(n6884), .ZN(n8258) );
  NAND2_X1 U4894 ( .A1(n7526), .A2(n7525), .ZN(n7524) );
  XNOR2_X1 U4895 ( .A(n4311), .B(n5592), .ZN(n7307) );
  AOI21_X1 U4896 ( .B1(n5129), .B2(n5132), .A(n5128), .ZN(n5127) );
  INV_X1 U4897 ( .A(n5101), .ZN(n4275) );
  NAND2_X1 U4898 ( .A1(n4649), .A2(n8092), .ZN(n8098) );
  NAND2_X1 U4899 ( .A1(n6456), .A2(n6455), .ZN(n8933) );
  AOI22_X1 U4900 ( .A1(n5967), .A2(n5966), .B1(n9119), .B2(n5965), .ZN(n5968)
         );
  OR2_X1 U4901 ( .A1(n5634), .A2(n9934), .ZN(n5651) );
  NAND2_X1 U4902 ( .A1(n7503), .A2(n4728), .ZN(n7472) );
  NAND2_X1 U4903 ( .A1(n5515), .A2(n5514), .ZN(n10032) );
  NAND2_X1 U4904 ( .A1(n4610), .A2(n5541), .ZN(n5565) );
  NAND2_X1 U4905 ( .A1(n7195), .A2(n7194), .ZN(n8094) );
  NAND2_X1 U4906 ( .A1(n4281), .A2(n5829), .ZN(n7503) );
  AND2_X1 U4907 ( .A1(n5497), .A2(n5496), .ZN(n10040) );
  INV_X1 U4908 ( .A(n5828), .ZN(n4281) );
  NAND2_X1 U4909 ( .A1(n5553), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5577) );
  NAND2_X1 U4910 ( .A1(n5525), .A2(n4615), .ZN(n4610) );
  AND2_X2 U4911 ( .A1(n7745), .A2(n10327), .ZN(n7747) );
  AND2_X1 U4912 ( .A1(n7511), .A2(n10229), .ZN(n7477) );
  INV_X1 U4913 ( .A(n5835), .ZN(n4274) );
  NAND2_X1 U4914 ( .A1(n6412), .A2(n6411), .ZN(n8243) );
  AND2_X1 U4915 ( .A1(n5453), .A2(n5452), .ZN(n7767) );
  NAND2_X1 U4916 ( .A1(n5410), .A2(n5409), .ZN(n10236) );
  NAND2_X1 U4917 ( .A1(n6384), .A2(n6383), .ZN(n10337) );
  NAND2_X1 U4918 ( .A1(n9307), .A2(n9357), .ZN(n7437) );
  NAND2_X1 U4919 ( .A1(n7418), .A2(n4291), .ZN(n7508) );
  NAND2_X1 U4920 ( .A1(n5434), .A2(n5433), .ZN(n10048) );
  XNOR2_X1 U4921 ( .A(n5450), .B(n5449), .ZN(n6979) );
  NAND2_X1 U4922 ( .A1(n5916), .A2(n7290), .ZN(n9398) );
  NAND2_X1 U4923 ( .A1(n5831), .A2(n9071), .ZN(n9357) );
  NAND2_X1 U4924 ( .A1(n5346), .A2(n5347), .ZN(n10198) );
  AND2_X1 U4925 ( .A1(n6352), .A2(n6351), .ZN(n7802) );
  AND4_X1 U4926 ( .A1(n5340), .A2(n5339), .A3(n5338), .A4(n5337), .ZN(n7471)
         );
  NAND2_X1 U4927 ( .A1(n5331), .A2(n4278), .ZN(n9071) );
  NAND2_X1 U4928 ( .A1(n5314), .A2(n4316), .ZN(n9458) );
  AND4_X1 U4929 ( .A1(n6308), .A2(n6307), .A3(n6306), .A4(n6305), .ZN(n7314)
         );
  AND2_X1 U4930 ( .A1(n5329), .A2(n5330), .ZN(n4278) );
  AND4_X1 U4931 ( .A1(n5298), .A2(n5297), .A3(n5296), .A4(n5295), .ZN(n7441)
         );
  AOI21_X1 U4932 ( .B1(n4403), .B2(n4959), .A(n4950), .ZN(n4949) );
  NAND2_X1 U4933 ( .A1(n4437), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5471) );
  CLKBUF_X3 U4934 ( .A(n9255), .Z(n4282) );
  AND2_X2 U4935 ( .A1(n10082), .A2(n10085), .ZN(n5336) );
  INV_X4 U4936 ( .A(n4785), .ZN(n5786) );
  INV_X1 U4937 ( .A(n5455), .ZN(n4437) );
  INV_X2 U4938 ( .A(n5317), .ZN(n9253) );
  INV_X1 U4939 ( .A(n5184), .ZN(n10082) );
  INV_X1 U4940 ( .A(n9283), .ZN(n7735) );
  AND2_X2 U4941 ( .A1(n5184), .A2(n10085), .ZN(n5730) );
  NAND2_X2 U4942 ( .A1(n6264), .A2(n8971), .ZN(n6319) );
  NAND2_X1 U4943 ( .A1(n6998), .A2(n5690), .ZN(n5317) );
  NAND2_X1 U4944 ( .A1(n5435), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5455) );
  NAND2_X1 U4945 ( .A1(n5245), .A2(n10078), .ZN(n10085) );
  INV_X1 U4946 ( .A(n5437), .ZN(n5435) );
  OAI21_X1 U4947 ( .B1(n6290), .B2(P2_IR_REG_27__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6245) );
  AND2_X1 U4948 ( .A1(n6171), .A2(n6170), .ZN(n6268) );
  NAND2_X1 U4949 ( .A1(n4693), .A2(n4692), .ZN(n10078) );
  NAND2_X1 U4950 ( .A1(n4721), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5253) );
  XNOR2_X1 U4951 ( .A(n5813), .B(n4736), .ZN(n9435) );
  NAND2_X1 U4952 ( .A1(n5324), .A2(n5323), .ZN(n5357) );
  OAI21_X2 U4953 ( .B1(n5868), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5865) );
  XNOR2_X1 U4954 ( .A(n6202), .B(n6133), .ZN(n7211) );
  NOR2_X1 U4955 ( .A1(n4798), .A2(n4360), .ZN(n4692) );
  INV_X1 U4956 ( .A(n4694), .ZN(n4693) );
  INV_X1 U4957 ( .A(n6176), .ZN(n6145) );
  AND2_X1 U4958 ( .A1(n5810), .A2(n5465), .ZN(n5491) );
  NAND2_X1 U4959 ( .A1(n5027), .A2(n5252), .ZN(n4798) );
  NOR2_X1 U4960 ( .A1(n6162), .A2(n6161), .ZN(n6163) );
  AND4_X2 U4961 ( .A1(n5232), .A2(n5231), .A3(n5624), .A4(n5230), .ZN(n5809)
         );
  INV_X1 U4962 ( .A(n5241), .ZN(n5027) );
  NAND3_X1 U4963 ( .A1(n6276), .A2(n4923), .A3(n4922), .ZN(n4929) );
  NAND4_X1 U4964 ( .A1(n5240), .A2(n5375), .A3(n5362), .A4(n5405), .ZN(n5241)
         );
  AND2_X1 U4965 ( .A1(n4280), .A2(n4279), .ZN(n5232) );
  NAND3_X1 U4966 ( .A1(n5254), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4928) );
  NAND2_X1 U4967 ( .A1(n5332), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5349) );
  INV_X1 U4968 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5405) );
  NOR2_X1 U4969 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5234) );
  INV_X1 U4970 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6212) );
  INV_X1 U4971 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5623) );
  AND2_X1 U4972 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5332) );
  NOR2_X1 U4973 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n4279) );
  NOR2_X1 U4974 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4280) );
  INV_X1 U4975 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5229) );
  INV_X1 U4976 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5490) );
  INV_X1 U4977 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5362) );
  NOR2_X2 U4978 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4790) );
  INV_X1 U4979 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4922) );
  INV_X1 U4980 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4923) );
  INV_X1 U4981 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n6276) );
  INV_X1 U4982 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5254) );
  NOR2_X1 U4983 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n5235) );
  NOR2_X1 U4984 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n5236) );
  INV_X2 U4985 ( .A(n9071), .ZN(n10224) );
  NAND2_X1 U4986 ( .A1(n7472), .A2(n5832), .ZN(n7475) );
  XNOR2_X2 U4987 ( .A(n5251), .B(n5250), .ZN(n5815) );
  XNOR2_X2 U4988 ( .A(n5253), .B(n5252), .ZN(n7014) );
  NAND2_X1 U4989 ( .A1(n5180), .A2(n9357), .ZN(n7468) );
  BUF_X8 U4990 ( .A(n5730), .Z(n4283) );
  OR2_X2 U4991 ( .A1(n10285), .A2(n10313), .ZN(n10277) );
  NAND3_X2 U4992 ( .A1(n4350), .A2(n6288), .A3(n6289), .ZN(n10285) );
  AND2_X4 U4993 ( .A1(n6943), .A2(n6114), .ZN(n5985) );
  AND2_X4 U4994 ( .A1(n8967), .A2(n8155), .ZN(n6345) );
  NOR2_X4 U4995 ( .A1(n8000), .A2(n8946), .ZN(n8736) );
  OR2_X2 U4996 ( .A1(n8748), .A2(n8243), .ZN(n8000) );
  OR2_X1 U4997 ( .A1(n8059), .A2(n9550), .ZN(n9349) );
  INV_X1 U4998 ( .A(n4935), .ZN(n4934) );
  OAI21_X1 U4999 ( .B1(n4937), .B2(n4936), .A(n5659), .ZN(n4935) );
  NAND2_X1 U5000 ( .A1(n9333), .A2(n9293), .ZN(n5849) );
  NAND2_X1 U5001 ( .A1(n5619), .A2(n5618), .ZN(n5641) );
  NAND2_X1 U5002 ( .A1(n5523), .A2(n5222), .ZN(n5525) );
  INV_X1 U5003 ( .A(n5311), .ZN(n5801) );
  NAND2_X1 U5004 ( .A1(n4369), .A2(n4911), .ZN(n4906) );
  NOR2_X1 U5005 ( .A1(n4913), .A2(n6681), .ZN(n4909) );
  AOI21_X1 U5006 ( .B1(n6702), .B2(n6742), .A(n4623), .ZN(n4622) );
  NAND2_X1 U5007 ( .A1(n4891), .A2(n6703), .ZN(n4890) );
  NAND2_X1 U5008 ( .A1(n4624), .A2(n6697), .ZN(n4623) );
  INV_X1 U5009 ( .A(n8587), .ZN(n4606) );
  NOR2_X1 U5010 ( .A1(n8125), .A2(n6730), .ZN(n4608) );
  INV_X1 U5011 ( .A(n4900), .ZN(n4899) );
  NAND2_X1 U5012 ( .A1(n4735), .A2(n4327), .ZN(n6752) );
  OAI211_X1 U5013 ( .C1(n9245), .C2(n9244), .A(n9240), .B(n4887), .ZN(n4886)
         );
  MUX2_X1 U5014 ( .A(n9239), .B(n9238), .S(n9267), .Z(n9240) );
  AOI21_X1 U5015 ( .B1(n4945), .B2(n4947), .A(n4943), .ZN(n4942) );
  INV_X1 U5016 ( .A(n5592), .ZN(n4943) );
  INV_X1 U5017 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5566) );
  NOR2_X1 U5018 ( .A1(n5152), .A2(n5149), .ZN(n5148) );
  INV_X1 U5019 ( .A(n6588), .ZN(n5149) );
  INV_X1 U5020 ( .A(n6749), .ZN(n5152) );
  NAND2_X1 U5021 ( .A1(n6587), .A2(n8397), .ZN(n6588) );
  XNOR2_X1 U5022 ( .A(n8149), .B(n8397), .ZN(n8130) );
  OR2_X1 U5023 ( .A1(n6580), .A2(n6579), .ZN(n6591) );
  NAND2_X1 U5024 ( .A1(n8536), .A2(n8537), .ZN(n4683) );
  AND2_X1 U5025 ( .A1(n8543), .A2(n8129), .ZN(n6737) );
  NAND2_X1 U5026 ( .A1(n8917), .A2(n8224), .ZN(n4835) );
  AND2_X1 U5027 ( .A1(n4831), .A2(n8596), .ZN(n4830) );
  NAND2_X1 U5028 ( .A1(n4833), .A2(n4832), .ZN(n4831) );
  INV_X1 U5029 ( .A(n4834), .ZN(n4832) );
  NOR2_X1 U5030 ( .A1(n8604), .A2(n8823), .ZN(n5072) );
  AOI21_X1 U5031 ( .B1(n4640), .B2(n4334), .A(n4639), .ZN(n4638) );
  INV_X1 U5032 ( .A(n6695), .ZN(n4643) );
  NAND2_X1 U5033 ( .A1(n4637), .A2(n4640), .ZN(n4636) );
  NAND2_X1 U5034 ( .A1(n4819), .A2(n4524), .ZN(n4523) );
  NAND2_X1 U5035 ( .A1(n5206), .A2(n5204), .ZN(n5203) );
  OR2_X1 U5036 ( .A1(n6423), .A2(n6422), .ZN(n6435) );
  NAND2_X1 U5037 ( .A1(n8312), .A2(n6340), .ZN(n6628) );
  NAND2_X1 U5038 ( .A1(n7539), .A2(n7594), .ZN(n7541) );
  NAND2_X1 U5039 ( .A1(n6646), .A2(n6644), .ZN(n7540) );
  INV_X1 U5040 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n6159) );
  INV_X1 U5041 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6140) );
  NOR2_X1 U5042 ( .A1(n9381), .A2(n4812), .ZN(n4811) );
  INV_X1 U5043 ( .A(n9343), .ZN(n4812) );
  NAND2_X1 U5044 ( .A1(n5710), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5747) );
  INV_X1 U5045 ( .A(n5711), .ZN(n5710) );
  NOR2_X1 U5046 ( .A1(n5855), .A2(n4547), .ZN(n4546) );
  INV_X1 U5047 ( .A(n9422), .ZN(n4547) );
  NOR2_X1 U5048 ( .A1(n5577), .A2(n5576), .ZN(n4440) );
  NAND2_X1 U5049 ( .A1(n7524), .A2(n5087), .ZN(n7688) );
  NOR2_X1 U5050 ( .A1(n9409), .A2(n5088), .ZN(n5087) );
  INV_X1 U5051 ( .A(n5834), .ZN(n5088) );
  INV_X1 U5052 ( .A(n9458), .ZN(n5831) );
  NAND2_X1 U5053 ( .A1(n9458), .A2(n10224), .ZN(n9307) );
  NOR2_X2 U5054 ( .A1(n9954), .A2(n5237), .ZN(n5238) );
  NAND2_X1 U5055 ( .A1(n5707), .A2(n5706), .ZN(n5724) );
  NAND2_X1 U5056 ( .A1(n5687), .A2(n5680), .ZN(n5688) );
  NAND2_X1 U5057 ( .A1(n5674), .A2(SI_21_), .ZN(n5675) );
  AOI21_X1 U5058 ( .B1(n4934), .B2(n4936), .A(n4932), .ZN(n4931) );
  INV_X1 U5059 ( .A(n5661), .ZN(n4932) );
  NAND2_X1 U5060 ( .A1(n5617), .A2(n4934), .ZN(n4580) );
  AND2_X1 U5061 ( .A1(n5661), .A2(n5647), .ZN(n5659) );
  NAND2_X1 U5062 ( .A1(n5641), .A2(n5621), .ZN(n5642) );
  NAND2_X1 U5063 ( .A1(n5613), .A2(n5612), .ZN(n5617) );
  NAND2_X1 U5064 ( .A1(n4463), .A2(n5506), .ZN(n5523) );
  NAND2_X1 U5065 ( .A1(n5445), .A2(n5444), .ZN(n5482) );
  XNOR2_X1 U5066 ( .A(n5396), .B(SI_7_), .ZN(n5391) );
  NAND2_X1 U5067 ( .A1(n8098), .A2(n4647), .ZN(n8308) );
  NOR2_X1 U5068 ( .A1(n7396), .A2(n4648), .ZN(n4647) );
  INV_X1 U5069 ( .A(n6782), .ZN(n4648) );
  AND2_X1 U5070 ( .A1(n7719), .A2(n7723), .ZN(n6932) );
  AND2_X1 U5071 ( .A1(n6917), .A2(n6639), .ZN(n7334) );
  NOR2_X1 U5072 ( .A1(n8504), .A2(n5147), .ZN(n5146) );
  AOI21_X1 U5073 ( .B1(n8616), .B2(n6573), .A(n6514), .ZN(n8346) );
  AND2_X1 U5074 ( .A1(n6507), .A2(n6506), .ZN(n8223) );
  NAND2_X1 U5075 ( .A1(n8397), .A2(n8324), .ZN(n8110) );
  NAND2_X1 U5076 ( .A1(n8140), .A2(n8130), .ZN(n8144) );
  NAND2_X1 U5077 ( .A1(n8128), .A2(n5223), .ZN(n8533) );
  NAND2_X1 U5078 ( .A1(n6527), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6548) );
  INV_X1 U5079 ( .A(n6528), .ZN(n6527) );
  NAND2_X1 U5080 ( .A1(n4529), .A2(n4528), .ZN(n8626) );
  NAND2_X1 U5081 ( .A1(n4371), .A2(n4532), .ZN(n4528) );
  NAND2_X1 U5082 ( .A1(n8660), .A2(n4345), .ZN(n4529) );
  NAND2_X1 U5083 ( .A1(n7955), .A2(n7954), .ZN(n8746) );
  NAND2_X1 U5084 ( .A1(n6628), .A2(n7575), .ZN(n7561) );
  OAI21_X1 U5085 ( .B1(n4709), .B2(n7625), .A(n7629), .ZN(n5967) );
  OR2_X2 U5086 ( .A1(n5184), .A2(n10085), .ZN(n4785) );
  AND2_X1 U5087 ( .A1(n9283), .A2(n9302), .ZN(n6944) );
  NOR2_X1 U5088 ( .A1(n6120), .A2(n6110), .ZN(n7292) );
  NOR2_X1 U5089 ( .A1(n9805), .A2(n9252), .ZN(n9431) );
  INV_X1 U5090 ( .A(n10085), .ZN(n4786) );
  NOR2_X1 U5091 ( .A1(n7268), .A2(n7267), .ZN(n7356) );
  XNOR2_X1 U5092 ( .A(n9497), .B(n9496), .ZN(n9473) );
  XNOR2_X1 U5093 ( .A(n4581), .B(n9681), .ZN(n9520) );
  NAND2_X1 U5094 ( .A1(n4583), .A2(n4582), .ZN(n4581) );
  NAND2_X1 U5095 ( .A1(n9511), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4582) );
  INV_X1 U5096 ( .A(n9510), .ZN(n4583) );
  OR2_X1 U5097 ( .A1(n9259), .A2(n9263), .ZN(n9350) );
  NAND2_X1 U5098 ( .A1(n4478), .A2(n4477), .ZN(n4483) );
  NAND2_X1 U5099 ( .A1(n9595), .A2(n4811), .ZN(n4808) );
  INV_X1 U5100 ( .A(n4810), .ZN(n4809) );
  OAI21_X1 U5101 ( .B1(n9381), .B2(n4813), .A(n9284), .ZN(n4810) );
  OR2_X1 U5102 ( .A1(n9395), .A2(n9394), .ZN(n9563) );
  AND2_X2 U5103 ( .A1(n9581), .A2(n9586), .ZN(n9582) );
  AOI21_X1 U5104 ( .B1(n5170), .B2(n4486), .A(n4789), .ZN(n4788) );
  NAND2_X1 U5105 ( .A1(n4355), .A2(n9676), .ZN(n4743) );
  NAND2_X1 U5106 ( .A1(n5650), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5664) );
  INV_X1 U5107 ( .A(n4439), .ZN(n5697) );
  OR2_X1 U5108 ( .A1(n9994), .A2(n9647), .ZN(n9334) );
  AOI21_X1 U5109 ( .B1(n5083), .B2(n5085), .A(n4864), .ZN(n5081) );
  NOR2_X1 U5110 ( .A1(n5562), .A2(n5090), .ZN(n5089) );
  INV_X1 U5111 ( .A(n5842), .ZN(n5090) );
  INV_X1 U5112 ( .A(n9278), .ZN(n6110) );
  NAND2_X1 U5113 ( .A1(n5865), .A2(n5864), .ZN(n5045) );
  OR2_X1 U5114 ( .A1(n5404), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5407) );
  OR2_X1 U5115 ( .A1(n5407), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5431) );
  AOI21_X1 U5116 ( .B1(n10080), .B2(n6328), .A(n6608), .ZN(n8900) );
  OR2_X1 U5117 ( .A1(n9553), .A2(n5801), .ZN(n5773) );
  INV_X1 U5118 ( .A(n6637), .ZN(n4915) );
  OAI21_X1 U5119 ( .B1(n6629), .B2(n6742), .A(n4916), .ZN(n6649) );
  NAND2_X1 U5120 ( .A1(n4917), .A2(n6742), .ZN(n4916) );
  NAND2_X1 U5121 ( .A1(n6628), .A2(n6648), .ZN(n4917) );
  NAND2_X1 U5122 ( .A1(n6683), .A2(n6742), .ZN(n4912) );
  NAND2_X1 U5123 ( .A1(n4374), .A2(n4911), .ZN(n4905) );
  NOR2_X1 U5124 ( .A1(n6710), .A2(n6709), .ZN(n4603) );
  OAI21_X1 U5125 ( .B1(n6711), .B2(n4604), .A(n4601), .ZN(n4599) );
  NAND2_X1 U5126 ( .A1(n4608), .A2(n4600), .ZN(n4597) );
  INV_X1 U5127 ( .A(n6731), .ZN(n4600) );
  NOR2_X1 U5128 ( .A1(n6735), .A2(n6736), .ZN(n4607) );
  INV_X1 U5129 ( .A(n6738), .ZN(n4920) );
  AND2_X1 U5130 ( .A1(n4863), .A2(n9218), .ZN(n4862) );
  INV_X1 U5131 ( .A(n9217), .ZN(n4863) );
  INV_X1 U5132 ( .A(n9670), .ZN(n4425) );
  OR2_X1 U5133 ( .A1(n6698), .A2(n4642), .ZN(n4641) );
  NAND2_X1 U5134 ( .A1(n6616), .A2(n6695), .ZN(n4642) );
  NAND2_X1 U5135 ( .A1(n9260), .A2(n9258), .ZN(n4729) );
  INV_X1 U5136 ( .A(n9292), .ZN(n5172) );
  NAND2_X1 U5137 ( .A1(n7409), .A2(n9457), .ZN(n9162) );
  NOR2_X1 U5138 ( .A1(n5642), .A2(n4938), .ZN(n4937) );
  INV_X1 U5139 ( .A(n5616), .ZN(n4938) );
  NAND2_X1 U5140 ( .A1(n5645), .A2(n5644), .ZN(n5661) );
  AOI21_X1 U5141 ( .B1(n4942), .B2(n4944), .A(n4364), .ZN(n4940) );
  INV_X1 U5142 ( .A(n4945), .ZN(n4944) );
  NAND2_X1 U5143 ( .A1(n5487), .A2(n5486), .ZN(n5506) );
  NOR2_X1 U5144 ( .A1(n4713), .A2(n4469), .ZN(n4468) );
  OAI21_X1 U5145 ( .B1(n4271), .B2(n4779), .A(n4778), .ZN(n5396) );
  NAND2_X1 U5146 ( .A1(n4271), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n4778) );
  OAI21_X1 U5147 ( .B1(n5690), .B2(n5361), .A(n5360), .ZN(n5392) );
  NAND2_X1 U5148 ( .A1(n5690), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n5360) );
  AND2_X1 U5149 ( .A1(n5126), .A2(n4383), .ZN(n4661) );
  NAND2_X1 U5150 ( .A1(n4661), .A2(n4659), .ZN(n4658) );
  INV_X1 U5151 ( .A(n6823), .ZN(n4659) );
  NAND2_X1 U5152 ( .A1(n4726), .A2(n8262), .ZN(n6844) );
  NAND2_X1 U5153 ( .A1(n8258), .A2(n8259), .ZN(n4726) );
  NAND2_X1 U5154 ( .A1(n8322), .A2(n5114), .ZN(n5113) );
  INV_X1 U5155 ( .A(n8191), .ZN(n5114) );
  OR2_X1 U5156 ( .A1(n4667), .A2(n6855), .ZN(n4666) );
  AOI21_X1 U5157 ( .B1(n5110), .B2(n5108), .A(n5107), .ZN(n5106) );
  INV_X1 U5158 ( .A(n6851), .ZN(n5107) );
  INV_X1 U5159 ( .A(n6845), .ZN(n5108) );
  AND2_X1 U5160 ( .A1(n6468), .A2(n6467), .ZN(n6488) );
  INV_X1 U5161 ( .A(n7334), .ZN(n6773) );
  NAND2_X1 U5162 ( .A1(n8175), .A2(n6841), .ZN(n8260) );
  AOI22_X1 U5163 ( .A1(n6627), .A2(n7609), .B1(n7333), .B2(n7719), .ZN(n6759)
         );
  AOI21_X1 U5164 ( .B1(n4899), .B2(n4901), .A(n4366), .ZN(n4897) );
  NOR2_X1 U5165 ( .A1(n6917), .A2(n4900), .ZN(n4895) );
  NAND2_X1 U5166 ( .A1(n6756), .A2(n6751), .ZN(n6755) );
  INV_X1 U5167 ( .A(n7200), .ZN(n4977) );
  NOR2_X1 U5168 ( .A1(n8781), .A2(n5076), .ZN(n5075) );
  INV_X1 U5169 ( .A(n5077), .ZN(n5076) );
  NAND2_X1 U5170 ( .A1(n4963), .A2(n4961), .ZN(n6740) );
  NOR2_X1 U5171 ( .A1(n8367), .A2(n4962), .ZN(n4961) );
  INV_X1 U5172 ( .A(n6567), .ZN(n4962) );
  OR2_X1 U5173 ( .A1(n8802), .A2(n8400), .ZN(n8126) );
  OR2_X1 U5174 ( .A1(n8555), .A2(n8551), .ZN(n8127) );
  NAND2_X1 U5175 ( .A1(n8582), .A2(n5138), .ZN(n5137) );
  INV_X1 U5176 ( .A(n4683), .ZN(n5225) );
  NAND2_X1 U5177 ( .A1(n8555), .A2(n6728), .ZN(n5141) );
  INV_X1 U5178 ( .A(n8933), .ZN(n5079) );
  NOR2_X1 U5179 ( .A1(n8938), .A2(n8739), .ZN(n5080) );
  NAND2_X1 U5180 ( .A1(n4300), .A2(n8757), .ZN(n4820) );
  INV_X1 U5181 ( .A(n6435), .ZN(n6434) );
  NOR2_X1 U5182 ( .A1(n6446), .A2(n9891), .ZN(n4678) );
  NOR2_X1 U5183 ( .A1(n7989), .A2(n5209), .ZN(n5208) );
  INV_X1 U5184 ( .A(n7956), .ZN(n5209) );
  AND2_X1 U5185 ( .A1(n7993), .A2(n5210), .ZN(n5206) );
  NAND2_X1 U5186 ( .A1(n6413), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6423) );
  INV_X1 U5187 ( .A(n6414), .ZN(n6413) );
  NAND2_X1 U5188 ( .A1(n7552), .A2(n6658), .ZN(n6375) );
  INV_X1 U5189 ( .A(n6343), .ZN(n4684) );
  AND2_X1 U5190 ( .A1(n8671), .A2(n8650), .ZN(n8651) );
  NOR2_X1 U5191 ( .A1(n8688), .A2(n8926), .ZN(n8671) );
  NAND2_X1 U5192 ( .A1(n6238), .A2(n9861), .ZN(n6148) );
  NOR2_X1 U5193 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n6155) );
  INV_X1 U5194 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6267) );
  NAND2_X1 U5195 ( .A1(n6040), .A2(n4284), .ZN(n4700) );
  INV_X1 U5196 ( .A(n4729), .ZN(n9392) );
  OAI21_X1 U5197 ( .B1(n4884), .B2(n4885), .A(n9249), .ZN(n9262) );
  AND2_X1 U5198 ( .A1(n4729), .A2(n9805), .ZN(n9266) );
  INV_X1 U5199 ( .A(n10134), .ZN(n4841) );
  INV_X1 U5200 ( .A(n10133), .ZN(n4840) );
  INV_X1 U5201 ( .A(n7359), .ZN(n5005) );
  NAND2_X1 U5202 ( .A1(n4484), .A2(n9384), .ZN(n4478) );
  NAND2_X1 U5203 ( .A1(n9595), .A2(n4480), .ZN(n4477) );
  NOR2_X1 U5204 ( .A1(n5774), .A2(n4481), .ZN(n4480) );
  INV_X1 U5205 ( .A(n4811), .ZN(n4481) );
  NAND2_X1 U5206 ( .A1(n4887), .A2(n4809), .ZN(n4484) );
  NAND2_X1 U5207 ( .A1(n5026), .A2(n9154), .ZN(n5025) );
  OR2_X1 U5208 ( .A1(n9980), .A2(n9093), .ZN(n9342) );
  OR2_X1 U5209 ( .A1(n9640), .A2(n5174), .ZN(n5173) );
  NOR2_X1 U5210 ( .A1(n9999), .A2(n10004), .ZN(n5018) );
  INV_X1 U5211 ( .A(n4802), .ZN(n4801) );
  NOR2_X1 U5212 ( .A1(n5182), .A2(n9209), .ZN(n4802) );
  NOR2_X1 U5213 ( .A1(n4358), .A2(n4805), .ZN(n4804) );
  INV_X1 U5214 ( .A(n9198), .ZN(n4805) );
  NAND2_X1 U5215 ( .A1(n5537), .A2(n9198), .ZN(n9746) );
  OR2_X1 U5216 ( .A1(n10029), .A2(n8045), .ZN(n9198) );
  NOR2_X1 U5217 ( .A1(n9313), .A2(n5169), .ZN(n5168) );
  INV_X1 U5218 ( .A(n9175), .ZN(n5169) );
  INV_X1 U5219 ( .A(n8024), .ZN(n4710) );
  INV_X1 U5220 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5869) );
  INV_X1 U5221 ( .A(n4937), .ZN(n4474) );
  NOR2_X1 U5222 ( .A1(n5526), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n5572) );
  AND2_X1 U5223 ( .A1(n5581), .A2(n5570), .ZN(n5583) );
  XNOR2_X1 U5224 ( .A(n5539), .B(SI_14_), .ZN(n5538) );
  NAND2_X1 U5225 ( .A1(n5510), .A2(n5509), .ZN(n5524) );
  AND2_X1 U5226 ( .A1(n5477), .A2(n5478), .ZN(n5481) );
  NOR2_X1 U5227 ( .A1(n5217), .A2(n4353), .ZN(n4939) );
  AND2_X1 U5228 ( .A1(n5462), .A2(n5461), .ZN(n5477) );
  XNOR2_X1 U5229 ( .A(n5483), .B(SI_11_), .ZN(n5478) );
  AND2_X1 U5230 ( .A1(n5462), .A2(n5430), .ZN(n5444) );
  NAND2_X1 U5231 ( .A1(n4467), .A2(n4466), .ZN(n5423) );
  NAND2_X1 U5232 ( .A1(n5423), .A2(n5388), .ZN(n5371) );
  NAND2_X1 U5233 ( .A1(n4767), .A2(n5321), .ZN(n5355) );
  AOI21_X1 U5234 ( .B1(n8342), .B2(n8341), .A(n6873), .ZN(n6877) );
  NAND2_X1 U5235 ( .A1(n4372), .A2(n4288), .ZN(n5118) );
  NAND2_X1 U5236 ( .A1(n5122), .A2(n6893), .ZN(n5121) );
  INV_X1 U5237 ( .A(n5123), .ZN(n5122) );
  NAND2_X1 U5238 ( .A1(n4288), .A2(n6893), .ZN(n5119) );
  AND2_X1 U5239 ( .A1(n6807), .A2(n6802), .ZN(n5125) );
  AOI21_X1 U5240 ( .B1(n5125), .B2(n4674), .A(n4673), .ZN(n4672) );
  INV_X1 U5241 ( .A(n6808), .ZN(n4673) );
  AND2_X1 U5242 ( .A1(n5111), .A2(n8287), .ZN(n5110) );
  NAND2_X1 U5243 ( .A1(n6845), .A2(n6846), .ZN(n5111) );
  NAND2_X1 U5244 ( .A1(n7660), .A2(n6818), .ZN(n7850) );
  NAND2_X1 U5245 ( .A1(n4682), .A2(n4681), .ZN(n6414) );
  NOR2_X1 U5246 ( .A1(n6404), .A2(n7976), .ZN(n4681) );
  INV_X1 U5247 ( .A(n4682), .ZN(n6405) );
  NAND2_X1 U5248 ( .A1(n8308), .A2(n6789), .ZN(n8307) );
  NOR2_X1 U5249 ( .A1(n8900), .A2(n8104), .ZN(n6757) );
  INV_X1 U5250 ( .A(n6755), .ZN(n6754) );
  INV_X1 U5251 ( .A(n5148), .ZN(n5143) );
  AND2_X1 U5252 ( .A1(n6566), .A2(n6565), .ZN(n8129) );
  OR2_X1 U5253 ( .A1(n8371), .A2(n6561), .ZN(n6566) );
  AOI21_X1 U5254 ( .B1(n8561), .B2(n6332), .A(n6553), .ZN(n8368) );
  AOI21_X1 U5255 ( .B1(n8576), .B2(n6573), .A(n6543), .ZN(n8299) );
  AND2_X1 U5256 ( .A1(n6524), .A2(n6523), .ZN(n8224) );
  OR2_X1 U5257 ( .A1(n8345), .A2(n6561), .ZN(n6524) );
  AND3_X1 U5258 ( .A1(n6472), .A2(n6471), .A3(n6470), .ZN(n8288) );
  AND4_X1 U5259 ( .A1(n6440), .A2(n6439), .A3(n6438), .A4(n6437), .ZN(n8384)
         );
  AND4_X1 U5260 ( .A1(n6428), .A2(n6427), .A3(n6426), .A4(n6425), .ZN(n8171)
         );
  NAND2_X1 U5261 ( .A1(n6311), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6300) );
  XOR2_X1 U5262 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n7211), .Z(n7200) );
  OR2_X1 U5263 ( .A1(n7164), .A2(n4979), .ZN(n4978) );
  AND2_X1 U5264 ( .A1(n6251), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4979) );
  NAND2_X1 U5265 ( .A1(n6252), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4975) );
  OAI21_X1 U5266 ( .B1(n4978), .B2(n4456), .A(n4454), .ZN(n4458) );
  NOR2_X1 U5267 ( .A1(n7213), .A2(n4455), .ZN(n4454) );
  NOR2_X1 U5268 ( .A1(n4977), .A2(n4456), .ZN(n4455) );
  INV_X1 U5269 ( .A(n4975), .ZN(n4456) );
  NAND2_X1 U5270 ( .A1(n4978), .A2(n4977), .ZN(n4976) );
  AND2_X1 U5271 ( .A1(n4458), .A2(n4457), .ZN(n7252) );
  NAND2_X1 U5272 ( .A1(n6253), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4457) );
  AND2_X1 U5273 ( .A1(n7279), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4973) );
  INV_X1 U5274 ( .A(n7496), .ZN(n4971) );
  OR2_X1 U5275 ( .A1(n6990), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4991) );
  NAND2_X1 U5276 ( .A1(n7811), .A2(n7810), .ZN(n7809) );
  AND2_X1 U5277 ( .A1(n4991), .A2(n4449), .ZN(n4448) );
  INV_X1 U5278 ( .A(n8033), .ZN(n4449) );
  AOI21_X1 U5279 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n6395), .A(n7675), .ZN(
        n7811) );
  XNOR2_X1 U5280 ( .A(n6257), .B(n8456), .ZN(n8454) );
  OR2_X1 U5281 ( .A1(n8466), .A2(n8476), .ZN(n4983) );
  AND2_X1 U5282 ( .A1(n6454), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4989) );
  NOR2_X1 U5283 ( .A1(n8475), .A2(n4452), .ZN(n6259) );
  AND2_X1 U5284 ( .A1(n6473), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4452) );
  AND2_X1 U5285 ( .A1(n6581), .A2(n6591), .ZN(n8510) );
  NAND2_X1 U5286 ( .A1(n8907), .A2(n8129), .ZN(n5199) );
  OR2_X1 U5287 ( .A1(n6548), .A2(n6547), .ZN(n6559) );
  NOR2_X1 U5288 ( .A1(n8555), .A2(n6728), .ZN(n4760) );
  NAND2_X1 U5289 ( .A1(n5136), .A2(n5141), .ZN(n5135) );
  NAND2_X1 U5290 ( .A1(n6554), .A2(n6536), .ZN(n5136) );
  AND2_X1 U5291 ( .A1(n8571), .A2(n8555), .ZN(n6554) );
  NAND2_X1 U5292 ( .A1(n8582), .A2(n10290), .ZN(n4645) );
  AND2_X1 U5293 ( .A1(n8553), .A2(n6726), .ZN(n8571) );
  NOR2_X1 U5294 ( .A1(n8124), .A2(n4838), .ZN(n4834) );
  AOI21_X1 U5295 ( .B1(n4834), .B2(n8123), .A(n4836), .ZN(n4833) );
  NOR2_X1 U5296 ( .A1(n8823), .A2(n8404), .ZN(n4836) );
  AND2_X1 U5297 ( .A1(n8583), .A2(n6721), .ZN(n8598) );
  NAND2_X1 U5298 ( .A1(n5166), .A2(n8123), .ZN(n8627) );
  AND2_X1 U5299 ( .A1(n6704), .A2(n6714), .ZN(n8641) );
  NAND2_X1 U5300 ( .A1(n8684), .A2(n8121), .ZN(n8660) );
  INV_X1 U5301 ( .A(n4523), .ZN(n4520) );
  NAND2_X1 U5302 ( .A1(n4522), .A2(n5201), .ZN(n4521) );
  INV_X1 U5303 ( .A(n4820), .ZN(n4821) );
  AND2_X1 U5304 ( .A1(n6694), .A2(n6701), .ZN(n8721) );
  OR2_X1 U5305 ( .A1(n8243), .A2(n8412), .ZN(n5210) );
  NAND2_X1 U5306 ( .A1(n7957), .A2(n5208), .ZN(n5207) );
  NAND2_X1 U5307 ( .A1(n5207), .A2(n5206), .ZN(n8719) );
  NAND2_X1 U5308 ( .A1(n8746), .A2(n8757), .ZN(n7957) );
  INV_X1 U5309 ( .A(n5129), .ZN(n4635) );
  NOR2_X1 U5310 ( .A1(n4632), .A2(n4631), .ZN(n4633) );
  NAND2_X1 U5311 ( .A1(n7926), .A2(n6672), .ZN(n8756) );
  NOR2_X1 U5312 ( .A1(n7930), .A2(n4527), .ZN(n4526) );
  INV_X1 U5313 ( .A(n7928), .ZN(n4527) );
  NAND2_X1 U5314 ( .A1(n7830), .A2(n4816), .ZN(n7895) );
  NOR2_X1 U5315 ( .A1(n6385), .A2(n4817), .ZN(n4816) );
  INV_X1 U5316 ( .A(n7829), .ZN(n4817) );
  AND2_X1 U5317 ( .A1(n6673), .A2(n6668), .ZN(n7899) );
  NAND2_X1 U5318 ( .A1(n7892), .A2(n7899), .ZN(n7891) );
  OR2_X1 U5319 ( .A1(n6369), .A2(n9937), .ZN(n6377) );
  NAND2_X1 U5320 ( .A1(n7548), .A2(n7551), .ZN(n7830) );
  NAND2_X1 U5321 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6343) );
  NAND2_X1 U5322 ( .A1(n4684), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6356) );
  NAND2_X1 U5323 ( .A1(n7561), .A2(n4518), .ZN(n4517) );
  INV_X1 U5324 ( .A(n7543), .ZN(n4518) );
  AND2_X1 U5325 ( .A1(n7561), .A2(n7540), .ZN(n4515) );
  NOR2_X1 U5326 ( .A1(n10277), .A2(n8090), .ZN(n7604) );
  OR2_X1 U5327 ( .A1(n6607), .A2(n6949), .ZN(n6288) );
  OR2_X1 U5328 ( .A1(n10328), .A2(n7723), .ZN(n7328) );
  NAND2_X1 U5329 ( .A1(n9254), .A2(n6328), .ZN(n4724) );
  NAND2_X1 U5330 ( .A1(n8508), .A2(n10331), .ZN(n4656) );
  NAND2_X1 U5331 ( .A1(n6517), .A2(n6516), .ZN(n8604) );
  NAND2_X1 U5332 ( .A1(n6500), .A2(n6499), .ZN(n8634) );
  INV_X1 U5333 ( .A(n8090), .ZN(n5133) );
  AND2_X1 U5334 ( .A1(n6291), .A2(n8961), .ZN(n4628) );
  OAI21_X1 U5335 ( .B1(n8961), .B2(n6291), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n4626) );
  NAND2_X1 U5336 ( .A1(n6291), .A2(n6293), .ZN(n6294) );
  INV_X1 U5337 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6244) );
  NAND2_X1 U5338 ( .A1(n6613), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6240) );
  CLKBUF_X1 U5339 ( .A(n6195), .Z(n6201) );
  XNOR2_X1 U5340 ( .A(n4707), .B(n4424), .ZN(n7625) );
  OAI21_X1 U5341 ( .B1(n7636), .B2(n5902), .A(n4708), .ZN(n4707) );
  NAND2_X1 U5342 ( .A1(n9123), .A2(n6097), .ZN(n4708) );
  INV_X1 U5343 ( .A(n4349), .ZN(n5035) );
  NAND2_X1 U5344 ( .A1(n6024), .A2(n6023), .ZN(n8990) );
  NAND2_X1 U5345 ( .A1(n4439), .A2(n5696), .ZN(n5711) );
  OR2_X1 U5346 ( .A1(n6051), .A2(n6050), .ZN(n9009) );
  NAND2_X1 U5347 ( .A1(n8980), .A2(n8981), .ZN(n5036) );
  AND2_X1 U5348 ( .A1(n4338), .A2(n4704), .ZN(n4702) );
  NAND2_X1 U5349 ( .A1(n4705), .A2(n6040), .ZN(n4704) );
  INV_X1 U5350 ( .A(n4706), .ZN(n4705) );
  INV_X1 U5351 ( .A(n6023), .ZN(n4718) );
  INV_X1 U5352 ( .A(n6024), .ZN(n4719) );
  NOR2_X1 U5353 ( .A1(n4321), .A2(n4700), .ZN(n4699) );
  AND2_X1 U5354 ( .A1(n7292), .A2(n9281), .ZN(n6117) );
  INV_X1 U5355 ( .A(n9142), .ZN(n5055) );
  NOR2_X1 U5356 ( .A1(n5057), .A2(n6029), .ZN(n9143) );
  NAND2_X1 U5357 ( .A1(n4585), .A2(n7018), .ZN(n7128) );
  NAND2_X1 U5358 ( .A1(n7125), .A2(n7124), .ZN(n4585) );
  AOI21_X1 U5359 ( .B1(n7019), .B2(n7128), .A(n7020), .ZN(n7037) );
  NAND2_X1 U5360 ( .A1(n7038), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5003) );
  NAND2_X1 U5361 ( .A1(n7104), .A2(n7105), .ZN(n4844) );
  NAND2_X1 U5362 ( .A1(n7095), .A2(n4842), .ZN(n10134) );
  NAND2_X1 U5363 ( .A1(n7091), .A2(n7703), .ZN(n4842) );
  AND2_X1 U5364 ( .A1(n10131), .A2(n10130), .ZN(n10128) );
  OR2_X1 U5365 ( .A1(n7356), .A2(n4395), .ZN(n4494) );
  NOR2_X1 U5366 ( .A1(n7614), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n4849) );
  NOR2_X1 U5367 ( .A1(n7364), .A2(n7363), .ZN(n7611) );
  INV_X1 U5368 ( .A(n7615), .ZN(n5007) );
  INV_X1 U5369 ( .A(n7616), .ZN(n5006) );
  OAI21_X1 U5370 ( .B1(n7364), .B2(n4594), .A(n4593), .ZN(n10152) );
  INV_X1 U5371 ( .A(n4595), .ZN(n4594) );
  AOI21_X1 U5372 ( .B1(n4595), .B2(n4849), .A(n4307), .ZN(n4593) );
  AOI21_X1 U5373 ( .B1(n7363), .B2(n4596), .A(n9463), .ZN(n4595) );
  NAND2_X1 U5374 ( .A1(n10152), .A2(n10151), .ZN(n4846) );
  OAI21_X1 U5375 ( .B1(n9473), .B2(n4499), .A(n4501), .ZN(n4498) );
  NAND2_X1 U5376 ( .A1(n10163), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4499) );
  NAND2_X1 U5377 ( .A1(n4500), .A2(n4294), .ZN(n4496) );
  AND2_X1 U5378 ( .A1(n4497), .A2(n4496), .ZN(n10158) );
  NOR2_X1 U5379 ( .A1(n4498), .A2(n10159), .ZN(n4497) );
  NOR2_X1 U5380 ( .A1(n9482), .A2(n4839), .ZN(n9484) );
  NOR2_X1 U5381 ( .A1(n9472), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n4839) );
  INV_X1 U5382 ( .A(n10170), .ZN(n4508) );
  NAND2_X1 U5383 ( .A1(n5800), .A2(n5799), .ZN(n9259) );
  AOI21_X1 U5384 ( .B1(n5093), .B2(n9395), .A(n4362), .ZN(n5092) );
  NAND2_X1 U5385 ( .A1(n9560), .A2(n5093), .ZN(n5091) );
  AOI21_X1 U5386 ( .B1(n4365), .B2(n4543), .A(n4541), .ZN(n4540) );
  NOR2_X1 U5387 ( .A1(n9589), .A2(n9977), .ZN(n4541) );
  INV_X1 U5388 ( .A(n4546), .ZN(n4545) );
  AOI21_X1 U5389 ( .B1(n4544), .B2(n4546), .A(n4328), .ZN(n4543) );
  INV_X1 U5390 ( .A(n4549), .ZN(n4544) );
  NOR2_X1 U5391 ( .A1(n5086), .A2(n4550), .ZN(n4549) );
  INV_X1 U5392 ( .A(n5853), .ZN(n4550) );
  INV_X1 U5393 ( .A(n5228), .ZN(n5086) );
  AOI21_X1 U5394 ( .B1(n5850), .B2(n5084), .A(n4348), .ZN(n5083) );
  INV_X1 U5395 ( .A(n5846), .ZN(n5084) );
  INV_X1 U5396 ( .A(n5850), .ZN(n5085) );
  INV_X1 U5397 ( .A(n4552), .ZN(n4551) );
  OAI21_X1 U5398 ( .B1(n5215), .B2(n4553), .A(n5845), .ZN(n4552) );
  INV_X1 U5399 ( .A(n5844), .ZN(n4553) );
  INV_X1 U5400 ( .A(n5849), .ZN(n9677) );
  AOI21_X1 U5401 ( .B1(n9205), .B2(n9295), .A(n9206), .ZN(n5182) );
  NAND2_X1 U5402 ( .A1(n5537), .A2(n4804), .ZN(n4803) );
  NAND2_X1 U5403 ( .A1(n9744), .A2(n5215), .ZN(n9731) );
  INV_X1 U5404 ( .A(n5555), .ZN(n5553) );
  AOI21_X1 U5405 ( .B1(n4536), .B2(n4539), .A(n4333), .ZN(n4533) );
  AND2_X1 U5406 ( .A1(n9196), .A2(n9764), .ZN(n9793) );
  NOR2_X1 U5407 ( .A1(n9358), .A2(n5179), .ZN(n5178) );
  INV_X1 U5408 ( .A(n9363), .ZN(n5367) );
  INV_X1 U5409 ( .A(n9357), .ZN(n5179) );
  NAND2_X1 U5410 ( .A1(n9534), .A2(n4775), .ZN(n5861) );
  AND2_X1 U5411 ( .A1(n9535), .A2(n4776), .ZN(n4775) );
  AND2_X1 U5412 ( .A1(n9533), .A2(n10234), .ZN(n4776) );
  NAND2_X1 U5413 ( .A1(n9429), .A2(n10234), .ZN(n4748) );
  NAND2_X1 U5414 ( .A1(n4791), .A2(n9799), .ZN(n4793) );
  XNOR2_X1 U5415 ( .A(n5808), .B(n9429), .ZN(n4791) );
  NAND2_X1 U5416 ( .A1(n5729), .A2(n5728), .ZN(n9828) );
  NAND2_X1 U5417 ( .A1(n5379), .A2(n5378), .ZN(n7698) );
  INV_X1 U5418 ( .A(n9123), .ZN(n10229) );
  NAND2_X1 U5419 ( .A1(n5859), .A2(n6109), .ZN(n10047) );
  AND2_X1 U5420 ( .A1(n7735), .A2(n9432), .ZN(n7088) );
  AND2_X1 U5421 ( .A1(n5809), .A2(n4324), .ZN(n4794) );
  AND2_X1 U5422 ( .A1(n5250), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n4796) );
  INV_X1 U5423 ( .A(n4798), .ZN(n4797) );
  NOR2_X1 U5424 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n5242), .ZN(n4795) );
  NAND2_X1 U5425 ( .A1(n5738), .A2(n5737), .ZN(n4960) );
  INV_X1 U5426 ( .A(n4577), .ZN(n4576) );
  OAI21_X1 U5427 ( .B1(n4290), .B2(n4578), .A(n5687), .ZN(n4577) );
  NAND2_X1 U5428 ( .A1(n5675), .A2(n4579), .ZN(n4578) );
  AND2_X1 U5429 ( .A1(n5706), .A2(n5693), .ZN(n5704) );
  NAND2_X1 U5430 ( .A1(n5617), .A2(n5616), .ZN(n5643) );
  XNOR2_X1 U5431 ( .A(n5565), .B(n5564), .ZN(n7119) );
  XNOR2_X1 U5432 ( .A(n5371), .B(n5369), .ZN(n6965) );
  OR2_X1 U5433 ( .A1(n4491), .A2(n5466), .ZN(n5288) );
  NOR2_X1 U5434 ( .A1(n10107), .A2(n10106), .ZN(n10108) );
  NAND2_X1 U5435 ( .A1(n4426), .A2(n10111), .ZN(n10112) );
  XNOR2_X1 U5436 ( .A(n6877), .B(n4669), .ZN(n8182) );
  INV_X1 U5437 ( .A(n6876), .ZN(n4669) );
  NAND2_X1 U5438 ( .A1(n8098), .A2(n6782), .ZN(n7395) );
  OR2_X1 U5439 ( .A1(n8377), .A2(n7313), .ZN(n8353) );
  NAND2_X1 U5440 ( .A1(n6930), .A2(n6932), .ZN(n8374) );
  INV_X1 U5441 ( .A(n6765), .ZN(n5155) );
  INV_X1 U5442 ( .A(n8129), .ZN(n8399) );
  NOR2_X1 U5443 ( .A1(n7276), .A2(n7275), .ZN(n7274) );
  NOR2_X1 U5444 ( .A1(n7237), .A2(n4974), .ZN(n7276) );
  AND2_X1 U5445 ( .A1(n6365), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4974) );
  INV_X1 U5446 ( .A(n4967), .ZN(n4966) );
  OAI21_X1 U5447 ( .B1(n6270), .B2(n10261), .A(n10260), .ZN(n4967) );
  NAND2_X1 U5448 ( .A1(n8110), .A2(n8109), .ZN(n8111) );
  XNOR2_X1 U5449 ( .A(n4741), .B(n4740), .ZN(n8112) );
  INV_X1 U5450 ( .A(n10279), .ZN(n10267) );
  NOR2_X1 U5451 ( .A1(n10276), .A2(n7726), .ZN(n10286) );
  AND2_X1 U5452 ( .A1(n10352), .A2(n10338), .ZN(n8873) );
  AND2_X1 U5453 ( .A1(n8770), .A2(n8773), .ZN(n8897) );
  NAND2_X1 U5454 ( .A1(n6576), .A2(n6575), .ZN(n8149) );
  NAND2_X1 U5455 ( .A1(n4826), .A2(n4825), .ZN(n4824) );
  INV_X1 U5456 ( .A(n8796), .ZN(n4825) );
  INV_X1 U5457 ( .A(n8795), .ZN(n4826) );
  AND2_X1 U5458 ( .A1(n10345), .A2(n10338), .ZN(n8947) );
  INV_X1 U5459 ( .A(n8947), .ZN(n8956) );
  AOI21_X1 U5460 ( .B1(n9633), .B2(n5311), .A(n5686), .ZN(n9648) );
  AOI21_X1 U5461 ( .B1(n5063), .B2(n5061), .A(n5060), .ZN(n5059) );
  AND2_X1 U5462 ( .A1(n5658), .A2(n5657), .ZN(n9647) );
  INV_X1 U5463 ( .A(n10040), .ZN(n7951) );
  NAND2_X1 U5464 ( .A1(n4766), .A2(n9031), .ZN(n4765) );
  INV_X1 U5465 ( .A(n9032), .ZN(n4766) );
  INV_X1 U5466 ( .A(n10016), .ZN(n9734) );
  AND2_X1 U5467 ( .A1(n5611), .A2(n5610), .ZN(n9054) );
  NAND2_X1 U5468 ( .A1(n5649), .A2(n5648), .ZN(n9994) );
  NAND2_X1 U5469 ( .A1(n5682), .A2(n5681), .ZN(n9984) );
  NAND2_X1 U5470 ( .A1(n6112), .A2(n9755), .ZN(n9138) );
  NOR2_X1 U5471 ( .A1(n9431), .A2(n4413), .ZN(n4867) );
  OR2_X1 U5472 ( .A1(n9441), .A2(n9442), .ZN(n4747) );
  AND2_X1 U5473 ( .A1(n5807), .A2(n5806), .ZN(n9263) );
  INV_X1 U5474 ( .A(n9550), .ZN(n9446) );
  INV_X1 U5475 ( .A(n9648), .ZN(n9448) );
  INV_X1 U5476 ( .A(n9220), .ZN(n9658) );
  INV_X1 U5477 ( .A(n9054), .ZN(n9714) );
  OR2_X1 U5478 ( .A1(n10128), .A2(n4323), .ZN(n5001) );
  NAND2_X1 U5479 ( .A1(n7360), .A2(n7359), .ZN(n7615) );
  INV_X1 U5480 ( .A(n4494), .ZN(n7360) );
  NOR2_X1 U5481 ( .A1(n4320), .A2(n9465), .ZN(n9482) );
  XNOR2_X1 U5482 ( .A(n9484), .B(n9500), .ZN(n10165) );
  NAND2_X1 U5483 ( .A1(n10165), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n10164) );
  OAI21_X1 U5484 ( .B1(n9520), .B2(n9519), .A(n9518), .ZN(n5010) );
  AOI21_X1 U5485 ( .B1(n9517), .B2(n10190), .A(n10188), .ZN(n9518) );
  NAND2_X1 U5486 ( .A1(n4490), .A2(n4488), .ZN(n4487) );
  NAND2_X1 U5487 ( .A1(n9520), .A2(n10143), .ZN(n4490) );
  NAND2_X1 U5488 ( .A1(n4489), .A2(n10190), .ZN(n4488) );
  INV_X1 U5489 ( .A(n9517), .ZN(n4489) );
  NAND2_X1 U5490 ( .A1(n4808), .A2(n4809), .ZN(n9548) );
  AOI21_X1 U5491 ( .B1(n9447), .B2(n9796), .A(n9568), .ZN(n9569) );
  AOI22_X1 U5492 ( .A1(n9590), .A2(n9796), .B1(n9794), .B2(n9589), .ZN(n5186)
         );
  NAND2_X1 U5493 ( .A1(n5188), .A2(n9799), .ZN(n5187) );
  NAND2_X1 U5494 ( .A1(n5094), .A2(n9393), .ZN(n4560) );
  NAND2_X1 U5495 ( .A1(n4568), .A2(n4567), .ZN(n4566) );
  OAI21_X1 U5496 ( .B1(n4568), .B2(n6606), .A(n4563), .ZN(n4562) );
  XNOR2_X1 U5497 ( .A(n5432), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7266) );
  NOR2_X1 U5498 ( .A1(n10378), .A2(n4421), .ZN(n10377) );
  NOR2_X1 U5499 ( .A1(n10377), .A2(n10376), .ZN(n10375) );
  NOR2_X1 U5500 ( .A1(n6649), .A2(n4914), .ZN(n6653) );
  NAND2_X1 U5501 ( .A1(n4915), .A2(n7599), .ZN(n4914) );
  INV_X1 U5502 ( .A(n4912), .ZN(n4910) );
  NAND2_X1 U5503 ( .A1(n4368), .A2(n4908), .ZN(n4907) );
  OR2_X1 U5504 ( .A1(n6683), .A2(n4913), .ZN(n4908) );
  NOR2_X1 U5505 ( .A1(n8732), .A2(n6687), .ZN(n4911) );
  NAND2_X1 U5506 ( .A1(n4620), .A2(n4619), .ZN(n4618) );
  OR2_X1 U5507 ( .A1(n8933), .A2(n4308), .ZN(n4619) );
  NAND2_X1 U5508 ( .A1(n8933), .A2(n4402), .ZN(n4620) );
  NOR2_X1 U5509 ( .A1(n4880), .A2(n4879), .ZN(n4878) );
  INV_X1 U5510 ( .A(n9167), .ZN(n4879) );
  INV_X1 U5511 ( .A(n9166), .ZN(n4880) );
  NAND2_X1 U5512 ( .A1(n8643), .A2(n6640), .ZN(n4624) );
  OR2_X1 U5513 ( .A1(n6694), .A2(n6742), .ZN(n4892) );
  NAND2_X1 U5514 ( .A1(n4883), .A2(n4881), .ZN(n9173) );
  AOI21_X1 U5515 ( .B1(n9160), .B2(n4882), .A(n9165), .ZN(n4881) );
  INV_X1 U5516 ( .A(n9242), .ZN(n4882) );
  AOI21_X1 U5517 ( .B1(n4750), .B2(n4749), .A(n4639), .ZN(n6706) );
  NOR2_X1 U5518 ( .A1(n6713), .A2(n6705), .ZN(n4749) );
  AND2_X1 U5519 ( .A1(n4609), .A2(n4602), .ZN(n4601) );
  NAND2_X1 U5520 ( .A1(n4606), .A2(n4603), .ZN(n4602) );
  NAND2_X1 U5521 ( .A1(n4606), .A2(n4605), .ZN(n4604) );
  INV_X1 U5522 ( .A(n6709), .ZN(n4605) );
  AND2_X1 U5523 ( .A1(n9201), .A2(n4875), .ZN(n4874) );
  NAND2_X1 U5524 ( .A1(n4329), .A2(n9319), .ZN(n4875) );
  NAND2_X1 U5525 ( .A1(n4864), .A2(n4860), .ZN(n4859) );
  INV_X1 U5526 ( .A(n9218), .ZN(n4860) );
  NAND2_X1 U5527 ( .A1(n4920), .A2(n8520), .ZN(n4919) );
  AND2_X1 U5528 ( .A1(n8130), .A2(n6741), .ZN(n4918) );
  AND3_X1 U5529 ( .A1(n4607), .A2(n4598), .A3(n4597), .ZN(n4921) );
  NAND2_X1 U5530 ( .A1(n4856), .A2(n4347), .ZN(n4854) );
  OR2_X1 U5531 ( .A1(n4862), .A2(n9663), .ZN(n4861) );
  MUX2_X1 U5532 ( .A(n9236), .B(n9561), .S(n9267), .Z(n9246) );
  NAND2_X1 U5533 ( .A1(n4756), .A2(n4903), .ZN(n4900) );
  NOR2_X1 U5534 ( .A1(n4901), .A2(n6742), .ZN(n4757) );
  NAND2_X1 U5535 ( .A1(n8900), .A2(n8104), .ZN(n6756) );
  NOR2_X1 U5536 ( .A1(n8720), .A2(n5208), .ZN(n5204) );
  INV_X1 U5537 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6139) );
  INV_X1 U5538 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6179) );
  OR2_X1 U5539 ( .A1(n6192), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n6218) );
  INV_X1 U5540 ( .A(SI_23_), .ZN(n9838) );
  INV_X1 U5541 ( .A(n5641), .ZN(n4936) );
  INV_X1 U5542 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5485) );
  NAND2_X1 U5543 ( .A1(n4723), .A2(n4722), .ZN(n5483) );
  OR2_X1 U5544 ( .A1(n4271), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n4723) );
  NAND2_X1 U5545 ( .A1(n4271), .A2(n6989), .ZN(n4722) );
  NAND2_X1 U5546 ( .A1(n4271), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5323) );
  OR2_X1 U5547 ( .A1(n4271), .A2(n5322), .ZN(n5324) );
  NOR2_X1 U5548 ( .A1(n6510), .A2(n8225), .ZN(n4680) );
  NOR2_X1 U5549 ( .A1(n6389), .A2(n6388), .ZN(n4682) );
  NAND2_X1 U5550 ( .A1(n8439), .A2(n4772), .ZN(n6257) );
  OR2_X1 U5551 ( .A1(n7062), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4772) );
  NOR2_X1 U5552 ( .A1(n8149), .A2(n8793), .ZN(n5077) );
  NOR2_X1 U5553 ( .A1(n8520), .A2(n8536), .ZN(n5195) );
  OAI21_X1 U5554 ( .B1(n8520), .B2(n5199), .A(n5198), .ZN(n5197) );
  OR2_X1 U5555 ( .A1(n8793), .A2(n8398), .ZN(n5198) );
  NAND2_X1 U5556 ( .A1(n5195), .A2(n5193), .ZN(n5192) );
  INV_X1 U5557 ( .A(n5223), .ZN(n5193) );
  NAND2_X1 U5558 ( .A1(n4680), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6528) );
  NAND2_X1 U5559 ( .A1(n8834), .A2(n8406), .ZN(n4532) );
  INV_X1 U5560 ( .A(n8122), .ZN(n4530) );
  NOR2_X1 U5561 ( .A1(n8834), .A2(n8406), .ZN(n4815) );
  NAND2_X1 U5562 ( .A1(n6488), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6501) );
  NOR2_X1 U5563 ( .A1(n8700), .A2(n4525), .ZN(n4524) );
  INV_X1 U5564 ( .A(n8118), .ZN(n4525) );
  INV_X1 U5565 ( .A(n6696), .ZN(n6616) );
  OR2_X1 U5566 ( .A1(n8933), .A2(n8386), .ZN(n6696) );
  NAND2_X1 U5567 ( .A1(n8933), .A2(n8386), .ZN(n6695) );
  INV_X1 U5568 ( .A(n6668), .ZN(n4634) );
  INV_X1 U5569 ( .A(n5127), .ZN(n4632) );
  NOR2_X1 U5570 ( .A1(n7828), .A2(n10337), .ZN(n5066) );
  AND2_X1 U5571 ( .A1(n6659), .A2(n6658), .ZN(n7547) );
  AND2_X1 U5572 ( .A1(n6630), .A2(n7575), .ZN(n6629) );
  AND2_X1 U5573 ( .A1(n8542), .A2(n8530), .ZN(n8525) );
  NOR2_X1 U5574 ( .A1(n8575), .A2(n5070), .ZN(n5068) );
  AND2_X1 U5575 ( .A1(n8736), .A2(n8943), .ZN(n8737) );
  AND2_X1 U5576 ( .A1(n6145), .A2(n6144), .ZN(n6171) );
  INV_X1 U5577 ( .A(n6171), .ZN(n6151) );
  OR2_X1 U5578 ( .A1(n9050), .A2(n6036), .ZN(n6039) );
  AOI21_X1 U5579 ( .B1(n5929), .B2(n9460), .A(n5928), .ZN(n5930) );
  OR2_X1 U5580 ( .A1(n10219), .A2(n6073), .ZN(n5925) );
  INV_X1 U5581 ( .A(n4702), .ZN(n4701) );
  INV_X1 U5582 ( .A(n4700), .ZN(n4698) );
  OAI21_X1 U5583 ( .B1(n5901), .B2(n9283), .A(n6097), .ZN(n5935) );
  NOR2_X1 U5584 ( .A1(n5054), .A2(n5053), .ZN(n5052) );
  INV_X1 U5585 ( .A(n9030), .ZN(n5054) );
  INV_X1 U5586 ( .A(n9088), .ZN(n5048) );
  NAND2_X1 U5587 ( .A1(n7266), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5002) );
  INV_X1 U5588 ( .A(n4849), .ZN(n4596) );
  INV_X1 U5589 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n4847) );
  NOR2_X1 U5590 ( .A1(n10141), .A2(n4492), .ZN(n9497) );
  AND2_X1 U5591 ( .A1(n9471), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4492) );
  NAND2_X1 U5592 ( .A1(n10187), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4995) );
  AND2_X1 U5593 ( .A1(n4543), .A2(n4318), .ZN(n4542) );
  NAND2_X1 U5594 ( .A1(n5173), .A2(n5172), .ZN(n4485) );
  OR2_X1 U5595 ( .A1(n10004), .A2(n9054), .ZN(n9214) );
  NAND2_X1 U5596 ( .A1(n5021), .A2(n10021), .ZN(n5020) );
  NOR2_X1 U5597 ( .A1(n5517), .A2(n5516), .ZN(n4438) );
  INV_X1 U5598 ( .A(n9746), .ZN(n5183) );
  NOR2_X1 U5599 ( .A1(n10029), .A2(n10032), .ZN(n5021) );
  AND2_X1 U5600 ( .A1(n9785), .A2(n4537), .ZN(n4536) );
  NAND2_X1 U5601 ( .A1(n4538), .A2(n5841), .ZN(n4537) );
  INV_X1 U5602 ( .A(n5841), .ZN(n4539) );
  INV_X1 U5603 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5516) );
  INV_X1 U5604 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5498) );
  OR2_X1 U5605 ( .A1(n5499), .A2(n5498), .ZN(n5517) );
  NAND2_X1 U5606 ( .A1(n4436), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5499) );
  INV_X1 U5607 ( .A(n5471), .ZN(n4436) );
  AOI21_X1 U5608 ( .B1(n5101), .B2(n5100), .A(n4352), .ZN(n5099) );
  INV_X1 U5609 ( .A(n5836), .ZN(n5100) );
  NOR2_X1 U5610 ( .A1(n7527), .A2(n10236), .ZN(n5014) );
  INV_X1 U5611 ( .A(n9162), .ZN(n5830) );
  AND2_X1 U5612 ( .A1(n9406), .A2(n7502), .ZN(n4728) );
  XNOR2_X1 U5613 ( .A(n10219), .B(n4554), .ZN(n9402) );
  INV_X1 U5614 ( .A(n7323), .ZN(n7082) );
  AND2_X1 U5615 ( .A1(n9745), .A2(n9295), .ZN(n9721) );
  NOR2_X1 U5616 ( .A1(n5690), .A2(n6956), .ZN(n4889) );
  NOR2_X1 U5617 ( .A1(n6603), .A2(n4571), .ZN(n4570) );
  INV_X1 U5618 ( .A(n6281), .ZN(n4571) );
  NAND2_X1 U5619 ( .A1(n5234), .A2(n5233), .ZN(n9954) );
  INV_X1 U5620 ( .A(n5688), .ZN(n4579) );
  NAND2_X1 U5621 ( .A1(n4940), .A2(n4476), .ZN(n5613) );
  OR2_X1 U5622 ( .A1(n4303), .A2(n5582), .ZN(n4945) );
  NAND2_X1 U5623 ( .A1(n5564), .A2(n5563), .ZN(n4948) );
  NOR2_X1 U5624 ( .A1(n5542), .A2(n4616), .ZN(n4615) );
  INV_X1 U5625 ( .A(n5524), .ZN(n4616) );
  INV_X1 U5626 ( .A(n5538), .ZN(n5542) );
  NAND2_X1 U5627 ( .A1(n4614), .A2(n5541), .ZN(n4613) );
  INV_X1 U5628 ( .A(n5564), .ZN(n4614) );
  NAND2_X1 U5629 ( .A1(n5448), .A2(SI_10_), .ZN(n5479) );
  XNOR2_X1 U5630 ( .A(n5359), .B(SI_5_), .ZN(n5358) );
  XNOR2_X1 U5631 ( .A(n5357), .B(SI_4_), .ZN(n5342) );
  OAI211_X1 U5632 ( .C1(n4929), .C2(n4927), .A(n4926), .B(n4924), .ZN(n5320)
         );
  NAND2_X1 U5633 ( .A1(n4925), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n4924) );
  INV_X1 U5634 ( .A(n4928), .ZN(n4925) );
  NOR2_X1 U5635 ( .A1(n8366), .A2(n5124), .ZN(n5123) );
  NAND2_X1 U5636 ( .A1(n10090), .A2(n6328), .ZN(n4963) );
  INV_X1 U5637 ( .A(n4661), .ZN(n4660) );
  AND2_X1 U5638 ( .A1(n4658), .A2(n6837), .ZN(n4657) );
  NAND2_X1 U5639 ( .A1(n8082), .A2(n5125), .ZN(n8204) );
  OR2_X1 U5640 ( .A1(n6501), .A2(n8327), .ZN(n6510) );
  INV_X1 U5641 ( .A(n4680), .ZN(n6518) );
  INV_X1 U5642 ( .A(n6879), .ZN(n8297) );
  OR2_X1 U5643 ( .A1(n7314), .A2(n7886), .ZN(n10283) );
  NAND2_X1 U5644 ( .A1(n8193), .A2(n6856), .ZN(n8190) );
  NAND2_X1 U5645 ( .A1(n4373), .A2(n4285), .ZN(n5112) );
  AOI21_X1 U5646 ( .B1(n7849), .B2(n6823), .A(n4410), .ZN(n5126) );
  INV_X1 U5647 ( .A(n5110), .ZN(n5109) );
  OR2_X1 U5648 ( .A1(n7341), .A2(n6929), .ZN(n8385) );
  NOR2_X1 U5649 ( .A1(n6931), .A2(n10303), .ZN(n6930) );
  OR2_X1 U5650 ( .A1(n7341), .A2(n8969), .ZN(n8383) );
  NOR2_X1 U5651 ( .A1(n4419), .A2(n6917), .ZN(n4896) );
  AND2_X1 U5652 ( .A1(n4677), .A2(n4676), .ZN(n8367) );
  INV_X1 U5653 ( .A(n6572), .ZN(n4676) );
  NAND2_X1 U5654 ( .A1(n8527), .A2(n6573), .ZN(n4677) );
  AND2_X1 U5655 ( .A1(n6535), .A2(n6534), .ZN(n6874) );
  OR2_X1 U5656 ( .A1(n8590), .A2(n6561), .ZN(n6535) );
  AND2_X1 U5657 ( .A1(n6482), .A2(n6481), .ZN(n8358) );
  AND4_X1 U5658 ( .A1(n6452), .A2(n6451), .A3(n6450), .A4(n6449), .ZN(n8117)
         );
  AND4_X1 U5659 ( .A1(n6419), .A2(n6418), .A3(n6417), .A4(n6416), .ZN(n7997)
         );
  AND4_X1 U5660 ( .A1(n6401), .A2(n6400), .A3(n6399), .A4(n6398), .ZN(n7973)
         );
  AND4_X1 U5661 ( .A1(n6394), .A2(n6393), .A3(n6392), .A4(n6391), .ZN(n7927)
         );
  AND4_X1 U5662 ( .A1(n6374), .A2(n6373), .A3(n6372), .A4(n6371), .ZN(n8206)
         );
  AND4_X1 U5663 ( .A1(n6361), .A2(n6360), .A3(n6359), .A4(n6358), .ZN(n7580)
         );
  OAI21_X1 U5664 ( .B1(n7250), .B2(n4451), .A(n4450), .ZN(n7239) );
  NAND2_X1 U5665 ( .A1(n4289), .A2(n4770), .ZN(n4451) );
  NAND2_X1 U5666 ( .A1(n7226), .A2(n4289), .ZN(n4450) );
  NOR2_X1 U5667 ( .A1(n7239), .A2(n7238), .ZN(n7237) );
  OAI22_X1 U5668 ( .A1(n7274), .A2(n4459), .B1(n4971), .B2(n4773), .ZN(n7677)
         );
  OR2_X1 U5669 ( .A1(n4773), .A2(n4973), .ZN(n4459) );
  AND2_X1 U5670 ( .A1(n6976), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4773) );
  NOR2_X1 U5671 ( .A1(n7677), .A2(n7676), .ZN(n7675) );
  AND2_X1 U5672 ( .A1(n4987), .A2(n4305), .ZN(n8465) );
  INV_X1 U5673 ( .A(n8466), .ZN(n4981) );
  OAI21_X1 U5674 ( .B1(n8128), .B2(n5194), .A(n5191), .ZN(n8139) );
  INV_X1 U5675 ( .A(n5195), .ZN(n5194) );
  AND2_X1 U5676 ( .A1(n5196), .A2(n5192), .ZN(n5191) );
  INV_X1 U5677 ( .A(n5197), .ZN(n5196) );
  INV_X1 U5678 ( .A(n8130), .ZN(n8141) );
  NAND2_X1 U5679 ( .A1(n6557), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6580) );
  OAI211_X1 U5680 ( .C1(n5137), .C2(n4683), .A(n4755), .B(n6574), .ZN(n8519)
         );
  AND2_X1 U5681 ( .A1(n8520), .A2(n8521), .ZN(n6574) );
  NAND2_X1 U5682 ( .A1(n5137), .A2(n5135), .ZN(n8554) );
  NAND2_X1 U5683 ( .A1(n8554), .A2(n5225), .ZN(n8535) );
  NAND2_X1 U5684 ( .A1(n4833), .A2(n4835), .ZN(n4828) );
  INV_X1 U5685 ( .A(n4835), .ZN(n4827) );
  NAND2_X1 U5686 ( .A1(n8612), .A2(n5072), .ZN(n8602) );
  OR2_X1 U5687 ( .A1(n8604), .A2(n8224), .ZN(n8583) );
  NAND2_X1 U5688 ( .A1(n6712), .A2(n6536), .ZN(n8587) );
  NAND2_X1 U5689 ( .A1(n4376), .A2(n6722), .ZN(n5164) );
  NAND2_X1 U5690 ( .A1(n4636), .A2(n4293), .ZN(n4644) );
  NAND2_X1 U5691 ( .A1(n8612), .A2(n8618), .ZN(n8613) );
  NAND2_X1 U5692 ( .A1(n4636), .A2(n4638), .ZN(n8629) );
  OAI21_X1 U5693 ( .B1(n8696), .B2(n6616), .A(n6695), .ZN(n8680) );
  NAND2_X1 U5694 ( .A1(n8736), .A2(n4297), .ZN(n8688) );
  NAND2_X1 U5695 ( .A1(n6434), .A2(n4306), .ZN(n6476) );
  NAND2_X1 U5696 ( .A1(n4820), .A2(n5201), .ZN(n4819) );
  NAND2_X1 U5697 ( .A1(n8736), .A2(n4287), .ZN(n8703) );
  NAND2_X1 U5698 ( .A1(n8736), .A2(n5080), .ZN(n8724) );
  NOR2_X1 U5699 ( .A1(n8732), .A2(n5163), .ZN(n5162) );
  INV_X1 U5700 ( .A(n6431), .ZN(n5163) );
  NAND2_X1 U5701 ( .A1(n6434), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6447) );
  NAND2_X1 U5702 ( .A1(n6434), .A2(n4678), .ZN(n6457) );
  NAND2_X1 U5703 ( .A1(n7747), .A2(n7823), .ZN(n7843) );
  NAND2_X1 U5704 ( .A1(n7747), .A2(n5066), .ZN(n7903) );
  OR2_X1 U5705 ( .A1(n6377), .A2(n6376), .ZN(n6389) );
  NAND2_X1 U5706 ( .A1(n6375), .A2(n6659), .ZN(n7835) );
  NAND2_X1 U5707 ( .A1(n7830), .A2(n7829), .ZN(n7831) );
  AND2_X1 U5708 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_REG3_REG_5__SCAN_IN), 
        .ZN(n4685) );
  AND2_X1 U5709 ( .A1(n6657), .A2(n6651), .ZN(n7738) );
  INV_X1 U5710 ( .A(n7561), .ZN(n7564) );
  CLKBUF_X1 U5711 ( .A(n7538), .Z(n7339) );
  AND2_X1 U5712 ( .A1(n7933), .A2(n10342), .ZN(n8868) );
  INV_X1 U5713 ( .A(n10326), .ZN(n10338) );
  INV_X1 U5714 ( .A(n7750), .ZN(n10327) );
  OR2_X1 U5715 ( .A1(n6932), .A2(n6915), .ZN(n10326) );
  AND2_X1 U5716 ( .A1(n7331), .A2(n7330), .ZN(n7402) );
  MUX2_X1 U5717 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8979), .S(n6319), .Z(n10313)
         );
  INV_X1 U5718 ( .A(n8868), .ZN(n10331) );
  NAND2_X1 U5719 ( .A1(n6934), .A2(n10312), .ZN(n10303) );
  XNOR2_X1 U5720 ( .A(n6238), .B(P2_IR_REG_22__SCAN_IN), .ZN(n6615) );
  INV_X1 U5721 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6146) );
  INV_X1 U5722 ( .A(n4438), .ZN(n5530) );
  INV_X1 U5723 ( .A(n5968), .ZN(n5061) );
  NAND2_X1 U5724 ( .A1(n4717), .A2(n4716), .ZN(n5060) );
  NAND2_X1 U5725 ( .A1(n5981), .A2(n7789), .ZN(n4716) );
  NAND2_X1 U5726 ( .A1(n5982), .A2(n5983), .ZN(n4717) );
  NAND2_X1 U5727 ( .A1(n4363), .A2(n4284), .ZN(n4706) );
  AND2_X1 U5728 ( .A1(n8998), .A2(n9029), .ZN(n4691) );
  INV_X1 U5729 ( .A(n5933), .ZN(n5043) );
  NAND2_X1 U5730 ( .A1(n7323), .A2(n5985), .ZN(n5913) );
  NAND2_X1 U5731 ( .A1(n5348), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5382) );
  INV_X1 U5732 ( .A(n5349), .ZN(n5348) );
  INV_X1 U5733 ( .A(n7625), .ZN(n9119) );
  CLKBUF_X1 U5734 ( .A(n9121), .Z(n4753) );
  OR3_X1 U5735 ( .A1(n6766), .A2(n7415), .A3(n6104), .ZN(n6120) );
  AOI21_X1 U5736 ( .B1(n9391), .B2(n9390), .A(n4340), .ZN(n9434) );
  NAND2_X1 U5737 ( .A1(n4730), .A2(n9392), .ZN(n9433) );
  NOR2_X1 U5738 ( .A1(n9430), .A2(n9431), .ZN(n4730) );
  AOI21_X1 U5739 ( .B1(n9392), .B2(n9353), .A(n9431), .ZN(n9354) );
  INV_X1 U5740 ( .A(n9435), .ZN(n9442) );
  NOR2_X1 U5741 ( .A1(n9266), .A2(n9265), .ZN(n9268) );
  NAND2_X1 U5742 ( .A1(n9391), .A2(n4731), .ZN(n9270) );
  NOR2_X1 U5743 ( .A1(n4732), .A2(n9264), .ZN(n4731) );
  NOR2_X1 U5744 ( .A1(n9263), .A2(n9267), .ZN(n4732) );
  AND2_X1 U5745 ( .A1(n5703), .A2(n5702), .ZN(n9093) );
  OR2_X1 U5746 ( .A1(n9612), .A2(n5801), .ZN(n5703) );
  AND2_X1 U5747 ( .A1(n5591), .A2(n5590), .ZN(n9722) );
  AND4_X1 U5748 ( .A1(n5416), .A2(n5415), .A3(n5414), .A4(n5413), .ZN(n7780)
         );
  NOR2_X1 U5749 ( .A1(n7037), .A2(n4354), .ZN(n7180) );
  AND2_X1 U5750 ( .A1(n5003), .A2(n4512), .ZN(n4511) );
  INV_X1 U5751 ( .A(n7177), .ZN(n4512) );
  NOR2_X1 U5752 ( .A1(n7050), .A2(n4319), .ZN(n7104) );
  NAND2_X1 U5753 ( .A1(n4592), .A2(n7042), .ZN(n7095) );
  NAND2_X1 U5754 ( .A1(n4844), .A2(n4843), .ZN(n4592) );
  INV_X1 U5755 ( .A(n7041), .ZN(n4843) );
  AND2_X1 U5756 ( .A1(n7097), .A2(n7098), .ZN(n4591) );
  NAND2_X1 U5757 ( .A1(n4841), .A2(n4840), .ZN(n10135) );
  NAND2_X1 U5758 ( .A1(n4841), .A2(n4344), .ZN(n4587) );
  NAND2_X1 U5759 ( .A1(n4590), .A2(n4589), .ZN(n4588) );
  INV_X1 U5760 ( .A(n4591), .ZN(n4590) );
  OAI21_X1 U5761 ( .B1(n10128), .B2(n4513), .A(n4998), .ZN(n7268) );
  OR2_X1 U5762 ( .A1(n4999), .A2(n4323), .ZN(n4513) );
  NAND2_X1 U5763 ( .A1(n7093), .A2(n5002), .ZN(n4998) );
  INV_X1 U5764 ( .A(n5002), .ZN(n4999) );
  NAND2_X1 U5765 ( .A1(n4493), .A2(n5004), .ZN(n10144) );
  AOI21_X1 U5766 ( .B1(n5005), .B2(n5008), .A(n4394), .ZN(n5004) );
  NAND2_X1 U5767 ( .A1(n4494), .A2(n5008), .ZN(n4493) );
  AND2_X1 U5768 ( .A1(n10144), .A2(n10145), .ZN(n10141) );
  NOR2_X1 U5769 ( .A1(n9501), .A2(n10158), .ZN(n10172) );
  OR2_X1 U5770 ( .A1(n9490), .A2(n9491), .ZN(n4851) );
  NAND2_X1 U5771 ( .A1(n10183), .A2(n4995), .ZN(n4506) );
  OR2_X1 U5772 ( .A1(n10170), .A2(n4507), .ZN(n4505) );
  NAND2_X1 U5773 ( .A1(n4995), .A2(n4406), .ZN(n4507) );
  AND2_X1 U5774 ( .A1(n4505), .A2(n4503), .ZN(n9510) );
  NOR2_X1 U5775 ( .A1(n9505), .A2(n4504), .ZN(n4503) );
  INV_X1 U5776 ( .A(n4506), .ZN(n4504) );
  XNOR2_X1 U5777 ( .A(n4584), .B(n9515), .ZN(n9517) );
  NAND2_X1 U5778 ( .A1(n4851), .A2(n4850), .ZN(n4584) );
  NAND2_X1 U5779 ( .A1(n9513), .A2(n9514), .ZN(n4850) );
  NOR2_X1 U5780 ( .A1(n8059), .A2(n5025), .ZN(n5024) );
  NAND2_X1 U5781 ( .A1(n5765), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n5784) );
  INV_X1 U5782 ( .A(n5766), .ZN(n5765) );
  INV_X1 U5783 ( .A(n4484), .ZN(n4479) );
  NAND2_X1 U5784 ( .A1(n9582), .A2(n9154), .ZN(n9571) );
  INV_X1 U5785 ( .A(n5025), .ZN(n5023) );
  NOR2_X1 U5786 ( .A1(n9562), .A2(n9561), .ZN(n9564) );
  AND2_X1 U5787 ( .A1(n4814), .A2(n4813), .ZN(n9562) );
  AND2_X1 U5788 ( .A1(n5718), .A2(n5717), .ZN(n9617) );
  OR2_X1 U5789 ( .A1(n9602), .A2(n5801), .ZN(n5718) );
  AND2_X1 U5790 ( .A1(n9336), .A2(n4485), .ZN(n5170) );
  NAND2_X1 U5791 ( .A1(n9675), .A2(n5171), .ZN(n4787) );
  NAND2_X1 U5792 ( .A1(n9697), .A2(n5018), .ZN(n9685) );
  OAI21_X1 U5793 ( .B1(n4801), .B2(n4804), .A(n4807), .ZN(n4800) );
  NAND2_X1 U5794 ( .A1(n4440), .A2(n5602), .ZN(n5634) );
  INV_X1 U5795 ( .A(n4440), .ZN(n5605) );
  AND2_X1 U5796 ( .A1(n9697), .A2(n9700), .ZN(n9699) );
  AND2_X1 U5797 ( .A1(n9322), .A2(n9205), .ZN(n9728) );
  NAND2_X1 U5798 ( .A1(n4438), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5555) );
  NAND2_X1 U5799 ( .A1(n5843), .A2(n5842), .ZN(n9742) );
  NOR2_X1 U5800 ( .A1(n5216), .A2(n5019), .ZN(n9773) );
  INV_X1 U5801 ( .A(n5021), .ZN(n5019) );
  OAI21_X1 U5802 ( .B1(n8008), .B2(n9190), .A(n9189), .ZN(n9792) );
  NOR2_X1 U5803 ( .A1(n5216), .A2(n10032), .ZN(n9786) );
  AND4_X1 U5804 ( .A1(n5522), .A2(n5521), .A3(n5520), .A4(n5519), .ZN(n9771)
         );
  NAND2_X1 U5805 ( .A1(n5098), .A2(n5099), .ZN(n7912) );
  NOR2_X1 U5806 ( .A1(n7864), .A2(n10043), .ZN(n7910) );
  AND4_X1 U5807 ( .A1(n5442), .A2(n5441), .A3(n5440), .A4(n5439), .ZN(n7858)
         );
  NAND2_X1 U5808 ( .A1(n5014), .A2(n5013), .ZN(n7864) );
  NAND2_X1 U5809 ( .A1(n5380), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5411) );
  INV_X1 U5810 ( .A(n5382), .ZN(n5380) );
  NAND2_X1 U5811 ( .A1(n7524), .A2(n5834), .ZN(n7686) );
  INV_X1 U5812 ( .A(n5014), .ZN(n7866) );
  AND2_X1 U5813 ( .A1(n9362), .A2(n9166), .ZN(n9410) );
  AND4_X1 U5814 ( .A1(n5387), .A2(n5386), .A3(n5385), .A4(n5384), .ZN(n7794)
         );
  NOR2_X1 U5815 ( .A1(n5627), .A2(n5625), .ZN(n4739) );
  NOR2_X1 U5816 ( .A1(n5630), .A2(n5629), .ZN(n4738) );
  NAND2_X1 U5817 ( .A1(n5310), .A2(n9356), .ZN(n7436) );
  NAND2_X1 U5818 ( .A1(n7418), .A2(n7485), .ZN(n5015) );
  INV_X1 U5819 ( .A(n6109), .ZN(n10199) );
  NAND2_X1 U5820 ( .A1(n7421), .A2(n9304), .ZN(n9365) );
  INV_X1 U5821 ( .A(n4727), .ZN(n9404) );
  NAND2_X1 U5822 ( .A1(n9401), .A2(n9398), .ZN(n7423) );
  AND2_X1 U5823 ( .A1(n9267), .A2(n9435), .ZN(n5896) );
  NAND2_X1 U5824 ( .A1(n7323), .A2(n7458), .ZN(n7298) );
  NAND2_X1 U5825 ( .A1(n9257), .A2(n9256), .ZN(n9808) );
  INV_X1 U5826 ( .A(n9560), .ZN(n5096) );
  NAND2_X1 U5827 ( .A1(n9697), .A2(n4286), .ZN(n5224) );
  AND2_X1 U5828 ( .A1(n5575), .A2(n5574), .ZN(n10016) );
  INV_X1 U5829 ( .A(n10033), .ZN(n10239) );
  NOR2_X1 U5830 ( .A1(n6768), .A2(n6767), .ZN(n7417) );
  NAND2_X1 U5831 ( .A1(n4568), .A2(n4564), .ZN(n4563) );
  NAND2_X1 U5832 ( .A1(n4565), .A2(n4567), .ZN(n4564) );
  INV_X1 U5833 ( .A(n4570), .ZN(n4565) );
  AOI21_X1 U5834 ( .B1(n4570), .B2(n4407), .A(n4569), .ZN(n4568) );
  INV_X1 U5835 ( .A(n6602), .ZN(n4569) );
  INV_X1 U5836 ( .A(n6606), .ZN(n4567) );
  NAND2_X1 U5837 ( .A1(n4574), .A2(n4398), .ZN(n5797) );
  XNOR2_X1 U5838 ( .A(n6604), .B(n6603), .ZN(n9254) );
  OAI21_X1 U5839 ( .B1(n6282), .B2(n4407), .A(n6281), .ZN(n6604) );
  NAND2_X1 U5840 ( .A1(n4574), .A2(n5777), .ZN(n4573) );
  INV_X1 U5841 ( .A(n4955), .ZN(n4950) );
  AOI21_X1 U5842 ( .B1(n4959), .B2(n4957), .A(n4956), .ZN(n4955) );
  INV_X1 U5843 ( .A(n5737), .ZN(n4957) );
  INV_X1 U5844 ( .A(n5776), .ZN(n4956) );
  NOR2_X1 U5845 ( .A1(n4958), .A2(n4953), .ZN(n4952) );
  XNOR2_X1 U5846 ( .A(n5877), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5890) );
  OAI21_X1 U5847 ( .B1(n5876), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5877) );
  XNOR2_X1 U5848 ( .A(n5757), .B(n5756), .ZN(n8049) );
  XNOR2_X1 U5849 ( .A(n5739), .B(n5738), .ZN(n8022) );
  XNOR2_X1 U5850 ( .A(n5866), .B(n5869), .ZN(n5891) );
  NAND2_X1 U5851 ( .A1(n5044), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5866) );
  XNOR2_X1 U5852 ( .A(n5724), .B(n5719), .ZN(n7923) );
  NAND2_X1 U5853 ( .A1(n4575), .A2(n5675), .ZN(n5689) );
  NAND2_X1 U5854 ( .A1(n5810), .A2(n5809), .ZN(n5868) );
  XNOR2_X1 U5855 ( .A(n5660), .B(n5659), .ZN(n7518) );
  AOI21_X1 U5856 ( .B1(n4473), .B2(n5612), .A(n4474), .ZN(n4472) );
  XNOR2_X1 U5857 ( .A(n4617), .B(n5583), .ZN(n7148) );
  OAI21_X1 U5858 ( .B1(n5525), .B2(n4613), .A(n4611), .ZN(n4617) );
  INV_X1 U5859 ( .A(n4612), .ZN(n4611) );
  OAI21_X1 U5860 ( .B1(n4615), .B2(n4613), .A(n5563), .ZN(n4612) );
  NAND2_X1 U5861 ( .A1(n5525), .A2(n5524), .ZN(n5543) );
  NAND2_X1 U5862 ( .A1(n5494), .A2(n5229), .ZN(n5526) );
  INV_X1 U5863 ( .A(n5493), .ZN(n5494) );
  NAND2_X1 U5864 ( .A1(n5482), .A2(n5481), .ZN(n4464) );
  XNOR2_X1 U5865 ( .A(n5403), .B(n5418), .ZN(n6960) );
  XNOR2_X1 U5866 ( .A(n5373), .B(n5391), .ZN(n6973) );
  OAI21_X1 U5867 ( .B1(n5283), .B2(n4271), .A(n5284), .ZN(n5304) );
  NAND2_X1 U5868 ( .A1(n5272), .A2(n5259), .ZN(n5261) );
  NAND2_X1 U5869 ( .A1(n6950), .A2(n5258), .ZN(n5259) );
  NOR2_X1 U5870 ( .A1(n10383), .A2(n10109), .ZN(n10110) );
  NAND2_X1 U5871 ( .A1(n4427), .A2(n10113), .ZN(n10114) );
  NAND2_X1 U5872 ( .A1(n8082), .A2(n6802), .ZN(n7644) );
  INV_X1 U5873 ( .A(n8181), .ZN(n4668) );
  OR2_X1 U5874 ( .A1(n7850), .A2(n7849), .ZN(n7969) );
  NAND2_X1 U5875 ( .A1(n6787), .A2(n6788), .ZN(n7396) );
  NAND2_X1 U5876 ( .A1(n8355), .A2(n6855), .ZN(n8193) );
  NAND2_X1 U5877 ( .A1(n5117), .A2(n5115), .ZN(n6926) );
  AOI21_X1 U5878 ( .B1(n5118), .B2(n5119), .A(n5116), .ZN(n5115) );
  INV_X1 U5879 ( .A(n6922), .ZN(n5116) );
  OAI21_X1 U5880 ( .B1(n6888), .B2(n5119), .A(n5118), .ZN(n6928) );
  AOI21_X1 U5881 ( .B1(n4672), .B2(n4675), .A(n4411), .ZN(n4671) );
  INV_X1 U5882 ( .A(n5125), .ZN(n4675) );
  INV_X1 U5883 ( .A(n10285), .ZN(n10320) );
  AND4_X1 U5884 ( .A1(n6410), .A2(n6409), .A3(n6408), .A4(n6407), .ZN(n8232)
         );
  INV_X1 U5885 ( .A(n8258), .ZN(n8261) );
  NAND2_X1 U5886 ( .A1(n5105), .A2(n5110), .ZN(n8352) );
  NAND2_X1 U5887 ( .A1(n4725), .A2(n6845), .ZN(n5105) );
  AND4_X1 U5888 ( .A1(n6382), .A2(n6381), .A3(n6380), .A4(n6379), .ZN(n7893)
         );
  NAND2_X1 U5889 ( .A1(n8190), .A2(n8191), .ZN(n8321) );
  NAND2_X1 U5890 ( .A1(n8321), .A2(n8322), .ZN(n8320) );
  NAND2_X1 U5891 ( .A1(n4662), .A2(n5126), .ZN(n8230) );
  NAND2_X1 U5892 ( .A1(n7850), .A2(n6823), .ZN(n4662) );
  NAND2_X1 U5893 ( .A1(n8094), .A2(n6777), .ZN(n4649) );
  NAND2_X1 U5894 ( .A1(n6798), .A2(n8076), .ZN(n8082) );
  INV_X1 U5895 ( .A(n8374), .ZN(n8387) );
  INV_X1 U5896 ( .A(n8377), .ZN(n8380) );
  INV_X1 U5897 ( .A(n8364), .ZN(n8392) );
  OAI21_X1 U5898 ( .B1(n8144), .B2(n5144), .A(n5142), .ZN(n6609) );
  NOR2_X1 U5899 ( .A1(n5145), .A2(n5146), .ZN(n5144) );
  AOI21_X1 U5900 ( .B1(n5145), .B2(n4296), .A(n4356), .ZN(n5142) );
  NAND2_X1 U5901 ( .A1(n6586), .A2(n6585), .ZN(n8397) );
  INV_X1 U5902 ( .A(n6874), .ZN(n8402) );
  INV_X1 U5903 ( .A(n8224), .ZN(n8403) );
  NAND4_X1 U5904 ( .A1(n6349), .A2(n6348), .A3(n6347), .A4(n6346), .ZN(n8419)
         );
  NAND2_X1 U5905 ( .A1(n6339), .A2(n5221), .ZN(n8420) );
  NAND2_X1 U5906 ( .A1(n6327), .A2(n6326), .ZN(n8421) );
  AND3_X1 U5907 ( .A1(n6325), .A2(n6324), .A3(n6323), .ZN(n6327) );
  NAND4_X1 U5908 ( .A1(n6303), .A2(n6302), .A3(n6301), .A4(n6300), .ZN(n6310)
         );
  OR2_X1 U5909 ( .A1(n6354), .A2(n6297), .ZN(n6303) );
  INV_X2 U5910 ( .A(P2_U3966), .ZN(n8422) );
  INV_X1 U5911 ( .A(n4978), .ZN(n7201) );
  INV_X1 U5912 ( .A(n4976), .ZN(n7199) );
  AND2_X1 U5913 ( .A1(n4976), .A2(n4975), .ZN(n7214) );
  NOR2_X1 U5914 ( .A1(n7250), .A2(n4769), .ZN(n7227) );
  INV_X1 U5915 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9937) );
  INV_X1 U5916 ( .A(n4972), .ZN(n7497) );
  OR2_X1 U5917 ( .A1(n7274), .A2(n4973), .ZN(n4972) );
  NAND2_X1 U5918 ( .A1(n7809), .A2(n4991), .ZN(n8032) );
  NAND2_X1 U5919 ( .A1(n8425), .A2(n8426), .ZN(n8424) );
  NAND2_X1 U5920 ( .A1(n4447), .A2(n4445), .ZN(n8425) );
  NAND2_X1 U5921 ( .A1(n4446), .A2(n4392), .ZN(n4445) );
  NAND2_X1 U5922 ( .A1(n7811), .A2(n4399), .ZN(n4447) );
  INV_X1 U5923 ( .A(n4448), .ZN(n4446) );
  NAND2_X1 U5924 ( .A1(n8440), .A2(n8441), .ZN(n8439) );
  NAND2_X1 U5925 ( .A1(n8424), .A2(n4771), .ZN(n8440) );
  OR2_X1 U5926 ( .A1(n7011), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4771) );
  INV_X1 U5927 ( .A(n8465), .ZN(n4986) );
  INV_X1 U5928 ( .A(n4989), .ZN(n4985) );
  NAND2_X1 U5929 ( .A1(n4453), .A2(n4984), .ZN(n8475) );
  NAND2_X1 U5930 ( .A1(n4989), .A2(n4988), .ZN(n4984) );
  NAND2_X1 U5931 ( .A1(n4980), .A2(n4987), .ZN(n4453) );
  XNOR2_X1 U5932 ( .A(n6259), .B(n7351), .ZN(n8496) );
  INV_X1 U5933 ( .A(n10261), .ZN(n10255) );
  AOI211_X1 U5934 ( .C1(n8504), .C2(n8503), .A(n10328), .B(n8502), .ZN(n8775)
         );
  XNOR2_X1 U5935 ( .A(n8139), .B(n8141), .ZN(n8508) );
  INV_X1 U5936 ( .A(n8149), .ZN(n6587) );
  XNOR2_X1 U5937 ( .A(n6580), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8527) );
  AND2_X1 U5938 ( .A1(n5200), .A2(n5199), .ZN(n8518) );
  NAND2_X1 U5939 ( .A1(n8533), .A2(n8534), .ZN(n5200) );
  AND2_X1 U5940 ( .A1(n6549), .A2(n6559), .ZN(n8561) );
  NAND2_X1 U5941 ( .A1(n8570), .A2(n4760), .ZN(n4759) );
  NAND2_X1 U5942 ( .A1(n8588), .A2(n8587), .ZN(n8811) );
  NAND2_X1 U5943 ( .A1(n4829), .A2(n4833), .ZN(n8597) );
  NAND2_X1 U5944 ( .A1(n8626), .A2(n4834), .ZN(n4829) );
  NAND2_X1 U5945 ( .A1(n8627), .A2(n6718), .ZN(n8620) );
  OAI21_X1 U5946 ( .B1(n8626), .B2(n8123), .A(n4837), .ZN(n8611) );
  NAND2_X1 U5947 ( .A1(n4531), .A2(n8122), .ZN(n8642) );
  NAND2_X1 U5948 ( .A1(n8660), .A2(n4314), .ZN(n4531) );
  NAND2_X1 U5949 ( .A1(n8702), .A2(n8120), .ZN(n8686) );
  NAND2_X1 U5950 ( .A1(n4818), .A2(n5201), .ZN(n8722) );
  NAND2_X1 U5951 ( .A1(n8746), .A2(n4821), .ZN(n4818) );
  NAND2_X1 U5952 ( .A1(n5207), .A2(n5210), .ZN(n7991) );
  NAND2_X1 U5953 ( .A1(n7957), .A2(n7956), .ZN(n7990) );
  OAI21_X1 U5954 ( .B1(n7926), .B2(n5132), .A(n5129), .ZN(n7959) );
  NAND2_X1 U5955 ( .A1(n8756), .A2(n6671), .ZN(n8760) );
  NAND2_X1 U5956 ( .A1(n7929), .A2(n7928), .ZN(n7931) );
  NAND2_X1 U5957 ( .A1(n7895), .A2(n7894), .ZN(n7898) );
  NAND2_X1 U5958 ( .A1(n7749), .A2(n10279), .ZN(n8763) );
  AND2_X1 U5959 ( .A1(n4516), .A2(n4517), .ZN(n7560) );
  OR2_X1 U5960 ( .A1(n6962), .A2(n6322), .ZN(n4742) );
  OR2_X1 U5961 ( .A1(n6607), .A2(n6948), .ZN(n6316) );
  INV_X1 U5962 ( .A(n10284), .ZN(n8769) );
  INV_X1 U5963 ( .A(n7802), .ZN(n8277) );
  OAI211_X1 U5964 ( .C1(n8794), .C2(n8868), .A(n4435), .B(n4433), .ZN(n8904)
         );
  NOR2_X1 U5965 ( .A1(n8791), .A2(n4434), .ZN(n4433) );
  INV_X1 U5966 ( .A(n8792), .ZN(n4435) );
  AND2_X1 U5967 ( .A1(n8793), .A2(n10338), .ZN(n4434) );
  INV_X1 U5968 ( .A(n8604), .ZN(n8917) );
  INV_X1 U5969 ( .A(n8634), .ZN(n8922) );
  AND2_X1 U5970 ( .A1(n6933), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10312) );
  NAND3_X1 U5971 ( .A1(n4629), .A2(n4627), .A3(n4625), .ZN(n8155) );
  OAI21_X1 U5972 ( .B1(n8961), .B2(P2_IR_REG_31__SCAN_IN), .A(n4626), .ZN(
        n4625) );
  CLKBUF_X1 U5973 ( .A(n6264), .Z(n8969) );
  INV_X1 U5974 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6246) );
  INV_X1 U5975 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n9863) );
  XNOR2_X1 U5976 ( .A(n6150), .B(n6149), .ZN(n7925) );
  NAND2_X1 U5977 ( .A1(n6168), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6150) );
  INV_X1 U5978 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7761) );
  INV_X1 U5979 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8101) );
  INV_X1 U5980 ( .A(n6615), .ZN(n8099) );
  INV_X1 U5981 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7610) );
  INV_X1 U5982 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n9938) );
  INV_X1 U5983 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n9943) );
  INV_X1 U5984 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7190) );
  INV_X1 U5985 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7122) );
  INV_X1 U5986 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7064) );
  INV_X1 U5987 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7013) );
  INV_X1 U5988 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9844) );
  OAI211_X1 U5989 ( .C1(n6194), .C2(n4994), .A(n6201), .B(n4992), .ZN(n7172)
         );
  NAND2_X1 U5990 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4994) );
  NAND2_X1 U5991 ( .A1(n6293), .A2(n4993), .ZN(n4992) );
  OAI211_X1 U5992 ( .C1(P2_IR_REG_31__SCAN_IN), .C2(P2_IR_REG_1__SCAN_IN), .A(
        n4444), .B(n4443), .ZN(n7161) );
  NAND3_X1 U5993 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .A3(
        P2_IR_REG_1__SCAN_IN), .ZN(n4443) );
  NAND2_X1 U5994 ( .A1(n4442), .A2(n4441), .ZN(n4444) );
  AND4_X1 U5995 ( .A1(n5352), .A2(n5351), .A3(n5353), .A4(n5354), .ZN(n7636)
         );
  AND2_X1 U5996 ( .A1(n5792), .A2(n5791), .ZN(n9550) );
  OR2_X1 U5997 ( .A1(n8055), .A2(n5801), .ZN(n5792) );
  NAND2_X1 U5998 ( .A1(n4349), .A2(n5032), .ZN(n5031) );
  NOR2_X1 U5999 ( .A1(n5035), .A2(n5030), .ZN(n5034) );
  NAND2_X1 U6000 ( .A1(n10090), .A2(n9253), .ZN(n5764) );
  NAND2_X1 U6001 ( .A1(n5695), .A2(n5694), .ZN(n9980) );
  AND4_X1 U6002 ( .A1(n5476), .A2(n5475), .A3(n5474), .A4(n5473), .ZN(n8009)
         );
  NAND2_X1 U6003 ( .A1(n9098), .A2(n5933), .ZN(n7373) );
  NAND2_X1 U6004 ( .A1(n7373), .A2(n7374), .ZN(n7372) );
  NAND2_X1 U6005 ( .A1(n9131), .A2(n5030), .ZN(n5029) );
  AND3_X1 U6006 ( .A1(n5561), .A2(n5560), .A3(n5559), .ZN(n9769) );
  AND2_X1 U6007 ( .A1(n5736), .A2(n5735), .ZN(n9567) );
  NAND2_X1 U6008 ( .A1(n4688), .A2(n4687), .ZN(n4715) );
  NAND2_X1 U6009 ( .A1(n9059), .A2(n5053), .ZN(n4687) );
  INV_X1 U6010 ( .A(n9059), .ZN(n4689) );
  NAND2_X1 U6011 ( .A1(n4697), .A2(n4695), .ZN(n9081) );
  INV_X1 U6012 ( .A(n4696), .ZN(n4695) );
  AND4_X1 U6013 ( .A1(n5535), .A2(n5534), .A3(n5533), .A4(n5532), .ZN(n8045)
         );
  AND2_X1 U6014 ( .A1(n5671), .A2(n5670), .ZN(n9220) );
  INV_X1 U6015 ( .A(n9150), .ZN(n9113) );
  NAND2_X1 U6016 ( .A1(n5992), .A2(n5991), .ZN(n7874) );
  NAND2_X1 U6017 ( .A1(n5365), .A2(n5364), .ZN(n9123) );
  OR2_X1 U6018 ( .A1(n6116), .A2(n9279), .ZN(n9148) );
  AND2_X1 U6019 ( .A1(n6117), .A2(n9279), .ZN(n9150) );
  INV_X1 U6020 ( .A(n9143), .ZN(n5056) );
  INV_X1 U6021 ( .A(n9093), .ZN(n9629) );
  INV_X1 U6022 ( .A(n9647), .ZN(n9678) );
  INV_X1 U6023 ( .A(n9112), .ZN(n9695) );
  INV_X1 U6024 ( .A(n8045), .ZN(n9797) );
  CLKBUF_X2 U6025 ( .A(P1_U4006), .Z(n9461) );
  INV_X1 U6026 ( .A(n4510), .ZN(n7175) );
  NAND2_X1 U6027 ( .A1(n7030), .A2(n5003), .ZN(n7176) );
  NAND2_X1 U6028 ( .A1(n4510), .A2(n4509), .ZN(n7055) );
  AND2_X1 U6029 ( .A1(n7056), .A2(n4301), .ZN(n4509) );
  INV_X1 U6030 ( .A(n4844), .ZN(n7106) );
  OAI21_X1 U6031 ( .B1(n7111), .B2(n7034), .A(n7113), .ZN(n7035) );
  NOR2_X1 U6032 ( .A1(n7035), .A2(n7036), .ZN(n7090) );
  NOR2_X1 U6033 ( .A1(n7090), .A2(n4514), .ZN(n10131) );
  NOR2_X1 U6034 ( .A1(n7096), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4514) );
  AND3_X1 U6035 ( .A1(n4588), .A2(n4587), .A3(n4586), .ZN(n7361) );
  INV_X1 U6036 ( .A(n7264), .ZN(n4586) );
  NAND2_X1 U6037 ( .A1(n4588), .A2(n4587), .ZN(n7265) );
  NOR2_X1 U6038 ( .A1(n7611), .A2(n4849), .ZN(n9462) );
  NAND2_X1 U6039 ( .A1(n7615), .A2(n5008), .ZN(n9468) );
  NOR2_X1 U6040 ( .A1(n5007), .A2(n5006), .ZN(n7617) );
  INV_X1 U6041 ( .A(n4846), .ZN(n10154) );
  NAND2_X1 U6042 ( .A1(n10148), .A2(n9464), .ZN(n4845) );
  NAND2_X1 U6043 ( .A1(n4496), .A2(n4495), .ZN(n10160) );
  INV_X1 U6044 ( .A(n4498), .ZN(n4495) );
  NAND2_X1 U6045 ( .A1(n9485), .A2(n10164), .ZN(n10178) );
  INV_X1 U6046 ( .A(n4997), .ZN(n10184) );
  NAND2_X1 U6047 ( .A1(n4508), .A2(n4406), .ZN(n4997) );
  INV_X1 U6048 ( .A(n4851), .ZN(n9512) );
  INV_X1 U6049 ( .A(n9808), .ZN(n9529) );
  AOI21_X1 U6050 ( .B1(n9794), .B2(n9447), .A(n8052), .ZN(n8053) );
  INV_X1 U6051 ( .A(n9977), .ZN(n9606) );
  OAI21_X1 U6052 ( .B1(n5854), .B2(n4545), .A(n4543), .ZN(n9594) );
  NAND2_X1 U6053 ( .A1(n4548), .A2(n9422), .ZN(n9609) );
  NAND2_X1 U6054 ( .A1(n5854), .A2(n4549), .ZN(n4548) );
  NAND2_X1 U6055 ( .A1(n5854), .A2(n5853), .ZN(n9624) );
  NAND2_X1 U6056 ( .A1(n9657), .A2(n9334), .ZN(n9644) );
  OAI21_X1 U6057 ( .B1(n9671), .B2(n5085), .A(n5083), .ZN(n9664) );
  NAND2_X1 U6058 ( .A1(n7451), .A2(n9253), .ZN(n5633) );
  NAND2_X1 U6059 ( .A1(n5082), .A2(n5850), .ZN(n9673) );
  NAND2_X1 U6060 ( .A1(n9671), .A2(n5846), .ZN(n5082) );
  NAND2_X1 U6061 ( .A1(n4803), .A2(n5181), .ZN(n9713) );
  INV_X1 U6062 ( .A(n5182), .ZN(n5181) );
  NAND2_X1 U6063 ( .A1(n9731), .A2(n5844), .ZN(n9708) );
  NAND2_X1 U6064 ( .A1(n5552), .A2(n5551), .ZN(n9759) );
  NAND2_X1 U6065 ( .A1(n8010), .A2(n9397), .ZN(n4535) );
  NAND2_X1 U6066 ( .A1(n5469), .A2(n5468), .ZN(n7920) );
  AND2_X1 U6067 ( .A1(n10209), .A2(n7464), .ZN(n9651) );
  NAND2_X1 U6068 ( .A1(n10209), .A2(n10199), .ZN(n9789) );
  INV_X1 U6069 ( .A(n10219), .ZN(n9102) );
  INV_X2 U6070 ( .A(n10209), .ZN(n10211) );
  AND2_X1 U6071 ( .A1(n9651), .A2(n10033), .ZN(n9802) );
  INV_X1 U6072 ( .A(n9789), .ZN(n9758) );
  INV_X1 U6073 ( .A(n9755), .ZN(n10201) );
  NAND2_X2 U6074 ( .A1(n7530), .A2(n9755), .ZN(n10209) );
  OAI21_X1 U6075 ( .B1(n9534), .B2(n4748), .A(n5821), .ZN(n4777) );
  NOR2_X1 U6076 ( .A1(n9825), .A2(n4781), .ZN(n4780) );
  INV_X1 U6077 ( .A(n9824), .ZN(n4782) );
  AND2_X1 U6078 ( .A1(n9826), .A2(n10047), .ZN(n4781) );
  INV_X1 U6079 ( .A(n5190), .ZN(n5189) );
  AND2_X1 U6080 ( .A1(n6943), .A2(n5892), .ZN(n9278) );
  NAND2_X1 U6081 ( .A1(n9278), .A2(n6983), .ZN(n10218) );
  NAND2_X1 U6082 ( .A1(n5244), .A2(n5243), .ZN(n5245) );
  NAND2_X1 U6083 ( .A1(n5242), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5243) );
  INV_X1 U6084 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n9930) );
  INV_X1 U6085 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8083) );
  CLKBUF_X1 U6086 ( .A(n5891), .Z(n8085) );
  INV_X1 U6087 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7757) );
  INV_X1 U6088 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7736) );
  INV_X1 U6089 ( .A(n9302), .ZN(n9432) );
  INV_X1 U6090 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7519) );
  INV_X1 U6091 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7465) );
  INV_X1 U6092 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7382) );
  INV_X1 U6093 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7310) );
  INV_X1 U6094 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7061) );
  INV_X1 U6095 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n7010) );
  INV_X1 U6096 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6989) );
  AND2_X1 U6097 ( .A1(n5408), .A2(n5431), .ZN(n10125) );
  NAND2_X1 U6098 ( .A1(n5299), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4852) );
  OAI21_X1 U6099 ( .B1(n5288), .B2(n5287), .A(n5299), .ZN(n7123) );
  XNOR2_X1 U6100 ( .A(n5256), .B(n5255), .ZN(n7067) );
  OAI21_X1 U6101 ( .B1(n10353), .B2(n10101), .A(n10355), .ZN(n10393) );
  AND2_X1 U6102 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10108), .ZN(n10382) );
  NOR2_X1 U6103 ( .A1(n10118), .A2(n10388), .ZN(n10380) );
  NOR2_X1 U6104 ( .A1(n10375), .A2(n4420), .ZN(n10374) );
  NAND2_X1 U6105 ( .A1(n10374), .A2(n10373), .ZN(n10372) );
  OAI21_X1 U6106 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10372), .ZN(n10370) );
  NAND2_X1 U6107 ( .A1(n10370), .A2(n10371), .ZN(n10369) );
  NAND2_X1 U6108 ( .A1(n10369), .A2(n4428), .ZN(n10367) );
  NAND2_X1 U6109 ( .A1(n10157), .A2(n4429), .ZN(n4428) );
  INV_X1 U6110 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n4429) );
  OAI21_X1 U6111 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10366), .ZN(n10364) );
  OAI21_X1 U6112 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10363), .ZN(n10361) );
  NAND2_X1 U6113 ( .A1(n10361), .A2(n10362), .ZN(n10360) );
  NAND2_X1 U6114 ( .A1(n10360), .A2(n4430), .ZN(n10358) );
  NAND2_X1 U6115 ( .A1(n4432), .A2(n4431), .ZN(n4430) );
  INV_X1 U6116 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n4432) );
  AND2_X1 U6117 ( .A1(n8306), .A2(n4397), .ZN(n4751) );
  NAND2_X1 U6118 ( .A1(n4970), .A2(n7723), .ZN(n4969) );
  AOI21_X1 U6119 ( .B1(n8137), .B2(n10284), .A(n8136), .ZN(n8138) );
  MUX2_X1 U6120 ( .A(n8771), .B(n8897), .S(n10352), .Z(n8772) );
  NAND2_X1 U6121 ( .A1(n4653), .A2(n9952), .ZN(n4652) );
  MUX2_X1 U6122 ( .A(n8798), .B(n8905), .S(n10352), .Z(n8799) );
  MUX2_X1 U6123 ( .A(n8898), .B(n8897), .S(n10345), .Z(n8899) );
  NAND2_X1 U6124 ( .A1(n4655), .A2(n8148), .ZN(n4654) );
  OAI21_X1 U6125 ( .B1(n8905), .B2(n4655), .A(n4822), .ZN(P2_U3514) );
  INV_X1 U6126 ( .A(n4823), .ZN(n4822) );
  OAI22_X1 U6127 ( .A1(n8907), .A2(n8956), .B1(n10345), .B2(n8906), .ZN(n4823)
         );
  AND2_X1 U6128 ( .A1(n9037), .A2(n4405), .ZN(n4783) );
  AND2_X1 U6129 ( .A1(n4746), .A2(n9443), .ZN(n4865) );
  INV_X1 U6130 ( .A(n5001), .ZN(n7094) );
  AOI21_X1 U6131 ( .B1(n10126), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n9521), .ZN(
        n5011) );
  NAND2_X1 U6132 ( .A1(n4487), .A2(n7464), .ZN(n5012) );
  NAND2_X1 U6133 ( .A1(n5010), .A2(n5893), .ZN(n5009) );
  INV_X1 U6134 ( .A(n4557), .ZN(n4559) );
  OAI211_X1 U6135 ( .C1(n9823), .C2(n4558), .A(n4408), .B(n4556), .ZN(P1_U3518) );
  NAND2_X1 U6136 ( .A1(n10245), .A2(n10234), .ZN(n4558) );
  NAND2_X1 U6137 ( .A1(n4557), .A2(n10245), .ZN(n4556) );
  OAI21_X1 U6138 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n10122), .A(n10385), .ZN(
        n10124) );
  AOI21_X1 U6139 ( .B1(n5151), .B2(n5147), .A(n5150), .ZN(n5145) );
  INV_X1 U6140 ( .A(n9131), .ZN(n5032) );
  NAND2_X1 U6141 ( .A1(n6029), .A2(n5055), .ZN(n4284) );
  OR2_X1 U6142 ( .A1(n6615), .A2(n6639), .ZN(n6915) );
  OR2_X1 U6143 ( .A1(n6868), .A2(n8218), .ZN(n4285) );
  XNOR2_X1 U6144 ( .A(n4852), .B(n5300), .ZN(n7031) );
  NOR2_X1 U6145 ( .A1(n4887), .A2(n9394), .ZN(n5093) );
  AND2_X1 U6146 ( .A1(n5018), .A2(n5017), .ZN(n4286) );
  AND2_X1 U6147 ( .A1(n5080), .A2(n5079), .ZN(n4287) );
  NAND2_X1 U6148 ( .A1(n6896), .A2(n6895), .ZN(n4288) );
  NAND2_X1 U6149 ( .A1(n6966), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4289) );
  NAND2_X1 U6150 ( .A1(n8155), .A2(n6298), .ZN(n6354) );
  AND4_X1 U6151 ( .A1(n6315), .A2(n6314), .A3(n6313), .A4(n6312), .ZN(n6778)
         );
  AND2_X1 U6152 ( .A1(n4931), .A2(n5672), .ZN(n4290) );
  INV_X1 U6153 ( .A(n4367), .ZN(n5147) );
  AND2_X1 U6154 ( .A1(n10224), .A2(n7485), .ZN(n4291) );
  INV_X1 U6155 ( .A(n6671), .ZN(n5132) );
  OAI211_X1 U6156 ( .C1(n4523), .C2(n4522), .A(n4357), .B(n4519), .ZN(n8684)
         );
  INV_X1 U6157 ( .A(n9395), .ZN(n5095) );
  AND2_X1 U6158 ( .A1(n5099), .A2(n4336), .ZN(n4292) );
  AND2_X1 U6159 ( .A1(n4638), .A2(n4346), .ZN(n4293) );
  NAND2_X1 U6160 ( .A1(n4404), .A2(n4521), .ZN(n8699) );
  AND2_X1 U6161 ( .A1(n4502), .A2(n9500), .ZN(n4294) );
  INV_X1 U6162 ( .A(n4486), .ZN(n5171) );
  OAI21_X1 U6163 ( .B1(n5173), .B2(n5175), .A(n5172), .ZN(n4486) );
  INV_X1 U6164 ( .A(n4959), .ZN(n4958) );
  AND2_X1 U6165 ( .A1(n4960), .A2(n5756), .ZN(n4959) );
  INV_X1 U6166 ( .A(n8575), .ZN(n8912) );
  NAND2_X1 U6167 ( .A1(n6539), .A2(n6538), .ZN(n8575) );
  AND2_X1 U6168 ( .A1(n5057), .A2(n6029), .ZN(n4295) );
  NAND2_X1 U6169 ( .A1(n5151), .A2(n5148), .ZN(n4296) );
  AND2_X1 U6170 ( .A1(n4287), .A2(n5078), .ZN(n4297) );
  AND3_X1 U6171 ( .A1(n5266), .A2(n5267), .A3(n5269), .ZN(n4298) );
  AND2_X1 U6172 ( .A1(n4370), .A2(n5029), .ZN(n4299) );
  AND2_X1 U6173 ( .A1(n5206), .A2(n5205), .ZN(n4300) );
  NAND2_X1 U6174 ( .A1(n7181), .A2(n7447), .ZN(n4301) );
  INV_X1 U6175 ( .A(n6714), .ZN(n4639) );
  AND2_X1 U6176 ( .A1(n5075), .A2(n5074), .ZN(n4302) );
  AND2_X1 U6177 ( .A1(n4948), .A2(n5583), .ZN(n4303) );
  AND2_X1 U6178 ( .A1(n4286), .A2(n5016), .ZN(n4304) );
  INV_X1 U6179 ( .A(n6679), .ZN(n5130) );
  AND2_X1 U6180 ( .A1(n4982), .A2(n4981), .ZN(n4305) );
  AND2_X1 U6181 ( .A1(n4678), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n4306) );
  AND3_X1 U6182 ( .A1(n6463), .A2(n6462), .A3(n6461), .ZN(n8386) );
  INV_X1 U6183 ( .A(n8386), .ZN(n4621) );
  AND2_X1 U6184 ( .A1(n4848), .A2(n4847), .ZN(n4307) );
  AND2_X1 U6185 ( .A1(n4621), .A2(n6742), .ZN(n4308) );
  AND2_X1 U6186 ( .A1(n5066), .A2(n5065), .ZN(n4309) );
  NAND2_X1 U6187 ( .A1(n7891), .A2(n6668), .ZN(n7926) );
  INV_X1 U6188 ( .A(n4283), .ZN(n5751) );
  INV_X1 U6189 ( .A(n4709), .ZN(n9118) );
  OAI21_X1 U6190 ( .B1(n6083), .B2(n7636), .A(n5958), .ZN(n4709) );
  INV_X1 U6191 ( .A(n8421), .ZN(n6783) );
  AND2_X1 U6192 ( .A1(n4630), .A2(n6291), .ZN(n4310) );
  INV_X1 U6193 ( .A(n7767), .ZN(n10043) );
  AND2_X1 U6194 ( .A1(n8967), .A2(n6299), .ZN(n6311) );
  AND2_X1 U6195 ( .A1(n4941), .A2(n4945), .ZN(n4311) );
  INV_X2 U6196 ( .A(n5985), .ZN(n5902) );
  NOR2_X1 U6197 ( .A1(n9699), .A2(n9698), .ZN(n4312) );
  NAND2_X1 U6198 ( .A1(n4853), .A2(n4555), .ZN(n9460) );
  AND2_X1 U6199 ( .A1(n4853), .A2(n4555), .ZN(n4554) );
  INV_X1 U6200 ( .A(n7263), .ZN(n4589) );
  NAND2_X1 U6201 ( .A1(n6590), .A2(n6589), .ZN(n8781) );
  NAND2_X1 U6202 ( .A1(n5058), .A2(n8992), .ZN(n5057) );
  AND2_X1 U6203 ( .A1(n5140), .A2(n6536), .ZN(n4313) );
  INV_X1 U6204 ( .A(n6311), .ZN(n6368) );
  INV_X1 U6205 ( .A(n5202), .ZN(n5201) );
  INV_X1 U6206 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8961) );
  OR2_X1 U6207 ( .A1(n8675), .A2(n8288), .ZN(n4314) );
  AND2_X1 U6208 ( .A1(n5289), .A2(n4888), .ZN(n4315) );
  NAND2_X1 U6209 ( .A1(n6147), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6238) );
  XNOR2_X1 U6210 ( .A(n8930), .B(n8408), .ZN(n8685) );
  AND3_X1 U6211 ( .A1(n5315), .A2(n5313), .A3(n5316), .ZN(n4316) );
  INV_X1 U6212 ( .A(n4500), .ZN(n9498) );
  OR2_X1 U6213 ( .A1(n9473), .A2(n9474), .ZN(n4500) );
  AND2_X1 U6214 ( .A1(n5940), .A2(n5939), .ZN(n4317) );
  XNOR2_X1 U6215 ( .A(n6240), .B(n6239), .ZN(n7609) );
  INV_X1 U6216 ( .A(n7609), .ZN(n6639) );
  NAND2_X1 U6217 ( .A1(n9977), .A2(n9589), .ZN(n4318) );
  AND2_X1 U6218 ( .A1(n7054), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n4319) );
  AND2_X1 U6219 ( .A1(n4846), .A2(n4845), .ZN(n4320) );
  INV_X1 U6220 ( .A(n9397), .ZN(n4538) );
  NAND2_X1 U6221 ( .A1(n9009), .A2(n6049), .ZN(n4321) );
  NAND2_X1 U6222 ( .A1(n7996), .A2(n6431), .ZN(n8731) );
  NOR2_X1 U6223 ( .A1(n9826), .A2(n9590), .ZN(n9395) );
  INV_X1 U6224 ( .A(n9293), .ZN(n5177) );
  INV_X1 U6225 ( .A(n6644), .ZN(n5160) );
  NAND2_X1 U6226 ( .A1(n4703), .A2(n4706), .ZN(n9038) );
  INV_X1 U6227 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6291) );
  AND2_X1 U6228 ( .A1(n6749), .A2(n4367), .ZN(n8785) );
  INV_X1 U6229 ( .A(n8785), .ZN(n4740) );
  NAND2_X1 U6230 ( .A1(n6433), .A2(n6432), .ZN(n8739) );
  AND2_X1 U6231 ( .A1(n8182), .A2(n4668), .ZN(n4322) );
  AND2_X1 U6232 ( .A1(n10125), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4323) );
  AND3_X1 U6233 ( .A1(n5028), .A2(n5238), .A3(n4796), .ZN(n4324) );
  INV_X1 U6234 ( .A(n9331), .ZN(n4807) );
  NAND2_X1 U6235 ( .A1(n5183), .A2(n5562), .ZN(n9745) );
  INV_X1 U6236 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6208) );
  OR2_X1 U6237 ( .A1(n8887), .A2(n7973), .ZN(n6672) );
  INV_X1 U6238 ( .A(n6672), .ZN(n5131) );
  AND2_X1 U6239 ( .A1(n4803), .A2(n4802), .ZN(n4325) );
  AND3_X1 U6240 ( .A1(n5058), .A2(n8992), .A3(n4698), .ZN(n4326) );
  AND3_X1 U6241 ( .A1(n6750), .A2(n6751), .A3(n5151), .ZN(n4327) );
  AND2_X1 U6242 ( .A1(n9980), .A2(n9629), .ZN(n4328) );
  AND2_X1 U6243 ( .A1(n9294), .A2(n9267), .ZN(n4329) );
  INV_X1 U6244 ( .A(n9805), .ZN(n9524) );
  NAND2_X1 U6245 ( .A1(n4733), .A2(n9251), .ZN(n9805) );
  AND2_X1 U6246 ( .A1(n4500), .A2(n4502), .ZN(n4330) );
  AND2_X1 U6247 ( .A1(n5092), .A2(n5097), .ZN(n4331) );
  OR2_X1 U6248 ( .A1(n9984), .A2(n9648), .ZN(n9336) );
  AND3_X1 U6249 ( .A1(n5028), .A2(n5027), .A3(n5238), .ZN(n4332) );
  OR2_X1 U6250 ( .A1(n8998), .A2(n9029), .ZN(n4690) );
  NOR2_X1 U6251 ( .A1(n8998), .A2(n9029), .ZN(n5053) );
  NAND2_X1 U6252 ( .A1(n5528), .A2(n5527), .ZN(n10029) );
  NAND2_X1 U6253 ( .A1(n5781), .A2(n5780), .ZN(n8059) );
  INV_X1 U6254 ( .A(n8247), .ZN(n5124) );
  AND2_X1 U6255 ( .A1(n10032), .A2(n9450), .ZN(n4333) );
  OR2_X1 U6256 ( .A1(n6698), .A2(n4643), .ZN(n4334) );
  OR2_X1 U6257 ( .A1(n4326), .A2(n4701), .ZN(n4335) );
  OR2_X1 U6258 ( .A1(n7920), .A2(n9451), .ZN(n4336) );
  OR2_X1 U6259 ( .A1(n6088), .A2(n6087), .ZN(n6089) );
  INV_X1 U6260 ( .A(n6089), .ZN(n5030) );
  AND2_X1 U6261 ( .A1(n6739), .A2(n6740), .ZN(n8520) );
  AND2_X1 U6262 ( .A1(n8051), .A2(n4482), .ZN(n4337) );
  AND2_X1 U6263 ( .A1(n10016), .A2(n9750), .ZN(n9206) );
  OR2_X1 U6264 ( .A1(n9819), .A2(n9566), .ZN(n9384) );
  NOR2_X1 U6265 ( .A1(n8504), .A2(n8107), .ZN(n6748) );
  INV_X1 U6266 ( .A(n6748), .ZN(n5151) );
  AND2_X1 U6267 ( .A1(n6039), .A2(n6038), .ZN(n4338) );
  NAND2_X1 U6268 ( .A1(n8612), .A2(n5069), .ZN(n5073) );
  AND2_X1 U6269 ( .A1(n9828), .A2(n9567), .ZN(n9236) );
  XNOR2_X1 U6270 ( .A(n5673), .B(SI_21_), .ZN(n5672) );
  INV_X1 U6271 ( .A(n9557), .ZN(n4887) );
  AND2_X1 U6272 ( .A1(n9582), .A2(n5023), .ZN(n4339) );
  OR2_X1 U6273 ( .A1(n9431), .A2(n9432), .ZN(n4340) );
  NOR2_X1 U6274 ( .A1(n5357), .A2(SI_4_), .ZN(n4341) );
  AND2_X1 U6275 ( .A1(n7896), .A2(n7894), .ZN(n4342) );
  INV_X1 U6276 ( .A(n4947), .ZN(n4946) );
  NAND2_X1 U6277 ( .A1(n5581), .A2(n5563), .ZN(n4947) );
  OR2_X1 U6278 ( .A1(n8634), .A2(n8223), .ZN(n6718) );
  INV_X1 U6279 ( .A(n6718), .ZN(n5165) );
  INV_X1 U6280 ( .A(n4838), .ZN(n4837) );
  AND2_X1 U6281 ( .A1(n4787), .A2(n5170), .ZN(n4343) );
  AND2_X1 U6282 ( .A1(n4840), .A2(n4589), .ZN(n4344) );
  AND2_X1 U6283 ( .A1(n4314), .A2(n4532), .ZN(n4345) );
  AND2_X1 U6284 ( .A1(n6722), .A2(n8123), .ZN(n4346) );
  AND2_X1 U6285 ( .A1(n8217), .A2(n6863), .ZN(n8322) );
  AND2_X1 U6286 ( .A1(n4857), .A2(n4861), .ZN(n4347) );
  INV_X1 U6287 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5252) );
  INV_X1 U6288 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5233) );
  AND2_X1 U6289 ( .A1(n9999), .A2(n9695), .ZN(n4348) );
  INV_X1 U6290 ( .A(n9289), .ZN(n5176) );
  NAND2_X1 U6291 ( .A1(n6096), .A2(n6095), .ZN(n4349) );
  OR2_X1 U6292 ( .A1(n6319), .A2(n7161), .ZN(n4350) );
  AND2_X1 U6293 ( .A1(n6679), .A2(n4910), .ZN(n4351) );
  NAND2_X1 U6294 ( .A1(n4890), .A2(n4622), .ZN(n4750) );
  NAND2_X1 U6295 ( .A1(n4963), .A2(n6567), .ZN(n8793) );
  AND2_X1 U6296 ( .A1(n9174), .A2(n9168), .ZN(n9409) );
  AND2_X1 U6297 ( .A1(n6672), .A2(n8755), .ZN(n7930) );
  NOR2_X1 U6298 ( .A1(n10043), .A2(n9452), .ZN(n4352) );
  NAND2_X1 U6299 ( .A1(n7895), .A2(n4342), .ZN(n7929) );
  AND2_X1 U6300 ( .A1(n5484), .A2(SI_11_), .ZN(n4353) );
  AND2_X1 U6301 ( .A1(n7038), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n4354) );
  AND3_X1 U6302 ( .A1(n4485), .A2(n9677), .A3(n9336), .ZN(n4355) );
  AND2_X1 U6303 ( .A1(n5227), .A2(n4641), .ZN(n4640) );
  INV_X1 U6304 ( .A(n7093), .ZN(n5000) );
  INV_X1 U6305 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5454) );
  AND2_X1 U6306 ( .A1(n5146), .A2(n5143), .ZN(n4356) );
  NAND2_X1 U6307 ( .A1(n9350), .A2(n9386), .ZN(n9535) );
  NOR2_X1 U6308 ( .A1(n5177), .A2(n5176), .ZN(n5175) );
  AND2_X1 U6309 ( .A1(n8679), .A2(n8120), .ZN(n4357) );
  NAND2_X1 U6310 ( .A1(n5562), .A2(n9322), .ZN(n4358) );
  NAND2_X1 U6311 ( .A1(n8999), .A2(n8998), .ZN(n4359) );
  NAND2_X1 U6312 ( .A1(n5250), .A2(n5242), .ZN(n4360) );
  AND2_X1 U6313 ( .A1(n6683), .A2(n6684), .ZN(n7989) );
  INV_X1 U6314 ( .A(n7989), .ZN(n5128) );
  INV_X1 U6315 ( .A(n5070), .ZN(n5069) );
  NAND2_X1 U6316 ( .A1(n5072), .A2(n5071), .ZN(n5070) );
  NAND2_X1 U6317 ( .A1(n5056), .A2(n5055), .ZN(n4361) );
  NOR2_X1 U6318 ( .A1(n9819), .A2(n9447), .ZN(n4362) );
  AND2_X1 U6319 ( .A1(n9342), .A2(n9378), .ZN(n9616) );
  INV_X1 U6320 ( .A(n9616), .ZN(n4789) );
  NOR2_X1 U6321 ( .A1(n6029), .A2(n5055), .ZN(n4363) );
  AND2_X1 U6322 ( .A1(n5594), .A2(SI_17_), .ZN(n4364) );
  AND2_X1 U6323 ( .A1(n4545), .A2(n4318), .ZN(n4365) );
  NOR2_X1 U6324 ( .A1(n6758), .A2(n6640), .ZN(n4366) );
  NAND2_X1 U6325 ( .A1(n8781), .A2(n7467), .ZN(n4367) );
  OR2_X1 U6326 ( .A1(n4912), .A2(n6684), .ZN(n4368) );
  OR2_X1 U6327 ( .A1(n4351), .A2(n4909), .ZN(n4369) );
  AND2_X1 U6328 ( .A1(n5036), .A2(n4349), .ZN(n4370) );
  OR2_X1 U6329 ( .A1(n4815), .A2(n4530), .ZN(n4371) );
  NAND2_X1 U6330 ( .A1(n5121), .A2(n8157), .ZN(n4372) );
  NAND2_X1 U6331 ( .A1(n6869), .A2(n5113), .ZN(n4373) );
  OR2_X1 U6332 ( .A1(n7993), .A2(n4907), .ZN(n4374) );
  AND2_X1 U6333 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_30__SCAN_IN), .ZN(
        n4375) );
  OR2_X1 U6334 ( .A1(n8619), .A2(n5165), .ZN(n4376) );
  AND2_X1 U6335 ( .A1(n8516), .A2(n8509), .ZN(n4377) );
  AND2_X1 U6336 ( .A1(n5864), .A2(n5233), .ZN(n4378) );
  OR2_X1 U6337 ( .A1(n8575), .A2(n8299), .ZN(n8553) );
  AND3_X1 U6338 ( .A1(n6155), .A2(n6267), .A3(n6146), .ZN(n4379) );
  INV_X1 U6339 ( .A(n9663), .ZN(n4864) );
  AND2_X1 U6340 ( .A1(n5024), .A2(n9586), .ZN(n4380) );
  AND2_X1 U6341 ( .A1(n9642), .A2(n9219), .ZN(n4381) );
  AND2_X1 U6342 ( .A1(n6385), .A2(n6659), .ZN(n4382) );
  AND2_X1 U6343 ( .A1(n9349), .A2(n9288), .ZN(n9427) );
  INV_X1 U6344 ( .A(n9427), .ZN(n5097) );
  AND2_X1 U6345 ( .A1(n8170), .A2(n8168), .ZN(n4383) );
  AND2_X1 U6346 ( .A1(n4285), .A2(n8322), .ZN(n4384) );
  OR2_X1 U6347 ( .A1(n8243), .A2(n7997), .ZN(n6683) );
  INV_X1 U6348 ( .A(n6856), .ZN(n4667) );
  AND2_X1 U6349 ( .A1(n5420), .A2(n5419), .ZN(n4385) );
  AND2_X1 U6350 ( .A1(n5997), .A2(n5991), .ZN(n4386) );
  INV_X1 U6351 ( .A(n5139), .ZN(n5138) );
  AND2_X1 U6352 ( .A1(n4517), .A2(n7544), .ZN(n4387) );
  AND2_X1 U6353 ( .A1(n4997), .A2(n4996), .ZN(n4388) );
  NAND2_X1 U6354 ( .A1(n6397), .A2(n6396), .ZN(n8887) );
  AND2_X1 U6355 ( .A1(n4465), .A2(n5444), .ZN(n4389) );
  NAND2_X1 U6356 ( .A1(n8116), .A2(n5203), .ZN(n5202) );
  INV_X1 U6357 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5250) );
  NOR2_X1 U6358 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n4390) );
  AND2_X1 U6359 ( .A1(n9179), .A2(n5102), .ZN(n5101) );
  INV_X1 U6360 ( .A(n5507), .ZN(n4465) );
  NAND2_X1 U6361 ( .A1(n5506), .A2(n5489), .ZN(n5507) );
  INV_X1 U6362 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9834) );
  INV_X1 U6363 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4993) );
  OR2_X1 U6364 ( .A1(n4830), .A2(n4827), .ZN(n4391) );
  AND2_X2 U6365 ( .A1(n7402), .A2(n7715), .ZN(n10352) );
  INV_X1 U6366 ( .A(n10352), .ZN(n4653) );
  OR2_X1 U6367 ( .A1(n8454), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4987) );
  INV_X1 U6368 ( .A(n8720), .ZN(n5205) );
  NAND2_X1 U6369 ( .A1(n6994), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4392) );
  INV_X1 U6370 ( .A(n5890), .ZN(n5894) );
  INV_X1 U6371 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n4927) );
  INV_X1 U6372 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n4930) );
  NAND2_X1 U6373 ( .A1(n4724), .A2(n6287), .ZN(n8504) );
  INV_X1 U6374 ( .A(n8504), .ZN(n5074) );
  NAND2_X1 U6375 ( .A1(n5161), .A2(n6644), .ZN(n7563) );
  NAND2_X1 U6376 ( .A1(n4535), .A2(n5841), .ZN(n9784) );
  NAND2_X1 U6377 ( .A1(n5443), .A2(n9175), .ZN(n7763) );
  XNOR2_X1 U6378 ( .A(n5614), .B(SI_18_), .ZN(n5612) );
  INV_X1 U6379 ( .A(n5612), .ZN(n4475) );
  AND2_X1 U6380 ( .A1(n6696), .A2(n6695), .ZN(n8700) );
  INV_X1 U6381 ( .A(n8700), .ZN(n8119) );
  XOR2_X1 U6382 ( .A(n6852), .B(n6853), .Z(n4393) );
  INV_X1 U6383 ( .A(n9991), .ZN(n5016) );
  INV_X1 U6384 ( .A(n9994), .ZN(n5017) );
  NAND2_X1 U6385 ( .A1(n6526), .A2(n6525), .ZN(n8813) );
  INV_X1 U6386 ( .A(n8813), .ZN(n5071) );
  AND2_X1 U6387 ( .A1(n9467), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4394) );
  AND2_X1 U6388 ( .A1(n7357), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4395) );
  NAND2_X1 U6389 ( .A1(n5764), .A2(n5763), .ZN(n9819) );
  INV_X1 U6390 ( .A(n9819), .ZN(n5026) );
  NAND2_X1 U6391 ( .A1(n7929), .A2(n4526), .ZN(n7955) );
  OR2_X1 U6392 ( .A1(n5216), .A2(n5020), .ZN(n4396) );
  OR2_X1 U6393 ( .A1(n8912), .A2(n8364), .ZN(n4397) );
  AND2_X1 U6394 ( .A1(n5777), .A2(n5793), .ZN(n4398) );
  AND2_X1 U6395 ( .A1(n7810), .A2(n4392), .ZN(n4399) );
  AND2_X1 U6396 ( .A1(n7809), .A2(n4448), .ZN(n4400) );
  AND2_X1 U6397 ( .A1(n4986), .A2(n4985), .ZN(n4401) );
  AND2_X1 U6398 ( .A1(n6496), .A2(n6495), .ZN(n8199) );
  INV_X1 U6399 ( .A(n8199), .ZN(n8406) );
  AND2_X1 U6400 ( .A1(n7618), .A2(n7616), .ZN(n5008) );
  INV_X1 U6401 ( .A(n4770), .ZN(n4769) );
  NAND2_X1 U6402 ( .A1(n6350), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4770) );
  NAND2_X1 U6403 ( .A1(n8386), .A2(n6640), .ZN(n4402) );
  AND2_X1 U6404 ( .A1(n5723), .A2(n5722), .ZN(n4403) );
  AND2_X1 U6405 ( .A1(n4819), .A2(n8118), .ZN(n4404) );
  AND2_X1 U6406 ( .A1(n6257), .A2(n8456), .ZN(n4990) );
  INV_X1 U6407 ( .A(n4990), .ZN(n4982) );
  OR2_X1 U6408 ( .A1(n9586), .A2(n9153), .ZN(n4405) );
  INV_X1 U6409 ( .A(n9140), .ZN(n9145) );
  NAND2_X1 U6410 ( .A1(n7030), .A2(n4511), .ZN(n4510) );
  NAND2_X1 U6411 ( .A1(n4423), .A2(n4424), .ZN(n9753) );
  AND2_X2 U6412 ( .A1(n7402), .A2(n7332), .ZN(n10345) );
  INV_X1 U6413 ( .A(n10345), .ZN(n4655) );
  INV_X1 U6414 ( .A(n8076), .ZN(n4674) );
  INV_X1 U6415 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n4679) );
  NAND2_X1 U6416 ( .A1(n10175), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4406) );
  NOR2_X1 U6417 ( .A1(n6280), .A2(SI_29_), .ZN(n4407) );
  AND2_X1 U6418 ( .A1(n5893), .A2(n7735), .ZN(n9267) );
  OR2_X1 U6419 ( .A1(n10245), .A2(n5770), .ZN(n4408) );
  INV_X1 U6420 ( .A(n8930), .ZN(n5078) );
  NAND2_X1 U6421 ( .A1(n6387), .A2(n6386), .ZN(n8891) );
  INV_X1 U6422 ( .A(n8891), .ZN(n5065) );
  INV_X1 U6423 ( .A(n10048), .ZN(n5013) );
  INV_X1 U6424 ( .A(n6114), .ZN(n5903) );
  NAND2_X1 U6425 ( .A1(n7597), .A2(n7543), .ZN(n7559) );
  AND2_X1 U6426 ( .A1(n7386), .A2(n5015), .ZN(n4409) );
  NAND2_X1 U6427 ( .A1(n8167), .A2(n6825), .ZN(n4410) );
  NAND2_X1 U6428 ( .A1(n6813), .A2(n6812), .ZN(n4411) );
  AND2_X1 U6429 ( .A1(n5001), .A2(n5000), .ZN(n4412) );
  OR2_X1 U6430 ( .A1(n9273), .A2(n9437), .ZN(n4413) );
  INV_X1 U6431 ( .A(n10183), .ZN(n4996) );
  AND2_X1 U6432 ( .A1(n4570), .A2(n6606), .ZN(n4414) );
  INV_X1 U6433 ( .A(n8476), .ZN(n4988) );
  NOR2_X1 U6434 ( .A1(n7227), .A2(n7226), .ZN(n4415) );
  AND2_X1 U6435 ( .A1(n6278), .A2(n6277), .ZN(n4416) );
  AND2_X1 U6436 ( .A1(n10135), .A2(n4591), .ZN(n4417) );
  AND2_X1 U6437 ( .A1(n4972), .A2(n4971), .ZN(n4418) );
  INV_X1 U6438 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6160) );
  INV_X1 U6439 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6239) );
  INV_X1 U6440 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6165) );
  AND2_X1 U6441 ( .A1(n6915), .A2(n6626), .ZN(n4419) );
  NAND2_X1 U6442 ( .A1(n6614), .A2(n6613), .ZN(n7719) );
  INV_X1 U6443 ( .A(n9467), .ZN(n4848) );
  XNOR2_X1 U6444 ( .A(n6269), .B(P2_IR_REG_19__SCAN_IN), .ZN(n7344) );
  AND2_X1 U6445 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n4420) );
  AND2_X1 U6446 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n4421) );
  AND2_X1 U6447 ( .A1(n4510), .A2(n4301), .ZN(n4422) );
  AND2_X1 U6448 ( .A1(n6241), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6764) );
  INV_X1 U6449 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4736) );
  INV_X1 U6450 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n4431) );
  INV_X1 U6451 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n4779) );
  NAND2_X1 U6452 ( .A1(n6114), .A2(n9283), .ZN(n4423) );
  NAND2_X1 U6453 ( .A1(n6113), .A2(n5903), .ZN(n4424) );
  OR2_X1 U6454 ( .A1(n5893), .A2(n7735), .ZN(n6113) );
  XNOR2_X1 U6455 ( .A(n5812), .B(P1_IR_REG_22__SCAN_IN), .ZN(n9283) );
  AND2_X1 U6456 ( .A1(n9302), .A2(n9435), .ZN(n6114) );
  OAI211_X1 U6457 ( .C1(n9813), .C2(n9753), .A(n9817), .B(n9818), .ZN(n4460)
         );
  NAND2_X1 U6458 ( .A1(n9162), .A2(n9161), .ZN(n9406) );
  NAND2_X1 U6459 ( .A1(n4534), .A2(n4533), .ZN(n9763) );
  NAND2_X1 U6460 ( .A1(n7958), .A2(n6683), .ZN(n7994) );
  NAND2_X1 U6461 ( .A1(n7598), .A2(n7599), .ZN(n5161) );
  AND2_X1 U6462 ( .A1(n9262), .A2(n9263), .ZN(n9250) );
  NAND2_X1 U6463 ( .A1(n9173), .A2(n4878), .ZN(n4877) );
  NAND2_X1 U6464 ( .A1(n4877), .A2(n4876), .ZN(n9169) );
  NAND2_X1 U6465 ( .A1(n9159), .A2(n9242), .ZN(n4883) );
  OAI21_X1 U6466 ( .B1(n9197), .B2(n9319), .A(n4874), .ZN(n4873) );
  NAND2_X1 U6467 ( .A1(n9306), .A2(n9356), .ZN(n4727) );
  NAND4_X1 U6468 ( .A1(n9210), .A2(n9217), .A3(n4425), .A4(n4864), .ZN(n4856)
         );
  NAND2_X1 U6469 ( .A1(n7910), .A2(n7980), .ZN(n8015) );
  OAI21_X1 U6470 ( .B1(n9823), .B2(n9753), .A(n4559), .ZN(n10054) );
  NOR2_X4 U6471 ( .A1(n9732), .A2(n10010), .ZN(n9697) );
  NAND2_X1 U6472 ( .A1(n9822), .A2(n9821), .ZN(n4557) );
  OAI21_X2 U6473 ( .B1(n4694), .B2(n4798), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5251) );
  NAND3_X1 U6474 ( .A1(n6145), .A2(n6163), .A3(n6144), .ZN(n6290) );
  NOR2_X2 U6475 ( .A1(n6143), .A2(n6142), .ZN(n6144) );
  NAND2_X1 U6476 ( .A1(n10381), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n4426) );
  NAND2_X1 U6477 ( .A1(n10392), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n4427) );
  NOR2_X1 U6478 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10382), .ZN(n10109) );
  NOR2_X1 U6479 ( .A1(n9268), .A2(n9242), .ZN(n4870) );
  NOR2_X2 U6480 ( .A1(n5664), .A2(n9022), .ZN(n4439) );
  INV_X1 U6481 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4442) );
  INV_X1 U6482 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4441) );
  INV_X1 U6483 ( .A(n4458), .ZN(n7212) );
  MUX2_X1 U6484 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n4460), .S(n10254), .Z(
        P1_U3551) );
  MUX2_X1 U6485 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n4460), .S(n10245), .Z(
        P1_U3519) );
  NAND2_X1 U6486 ( .A1(n5445), .A2(n4389), .ZN(n4462) );
  NAND2_X1 U6487 ( .A1(n4461), .A2(n4939), .ZN(n4463) );
  OAI21_X1 U6488 ( .B1(n5481), .B2(n5507), .A(n4462), .ZN(n4461) );
  NAND2_X1 U6489 ( .A1(n5422), .A2(n5421), .ZN(n4470) );
  NAND3_X1 U6490 ( .A1(n5422), .A2(n4467), .A3(n4466), .ZN(n4471) );
  NAND2_X1 U6491 ( .A1(n4468), .A2(n4767), .ZN(n4466) );
  NOR2_X1 U6492 ( .A1(n5358), .A2(n4341), .ZN(n4467) );
  INV_X1 U6493 ( .A(n5321), .ZN(n4469) );
  NAND3_X1 U6494 ( .A1(n4471), .A2(n4385), .A3(n4470), .ZN(n5425) );
  NAND2_X1 U6495 ( .A1(n5565), .A2(n4942), .ZN(n4476) );
  INV_X1 U6496 ( .A(n4940), .ZN(n4473) );
  OAI21_X1 U6497 ( .B1(n4476), .B2(n4475), .A(n4472), .ZN(n4933) );
  NAND3_X1 U6498 ( .A1(n4478), .A2(n4477), .A3(n5097), .ZN(n4482) );
  NAND2_X1 U6499 ( .A1(n4483), .A2(n9427), .ZN(n8051) );
  NAND3_X2 U6500 ( .A1(n4790), .A2(n4491), .A3(n5239), .ZN(n5327) );
  NAND2_X1 U6501 ( .A1(n4491), .A2(n4790), .ZN(n5325) );
  NOR2_X4 U6502 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n4491) );
  INV_X1 U6503 ( .A(n9499), .ZN(n4502) );
  NAND2_X1 U6504 ( .A1(n9499), .A2(n10163), .ZN(n4501) );
  NAND2_X1 U6505 ( .A1(n4505), .A2(n4506), .ZN(n9504) );
  NAND2_X1 U6506 ( .A1(n6636), .A2(n10287), .ZN(n7338) );
  NAND2_X1 U6507 ( .A1(n10320), .A2(n6310), .ZN(n10287) );
  NAND2_X1 U6508 ( .A1(n4516), .A2(n4387), .ZN(n7573) );
  NAND3_X1 U6509 ( .A1(n7542), .A2(n7541), .A3(n4515), .ZN(n4516) );
  NAND3_X1 U6510 ( .A1(n7542), .A2(n7540), .A3(n7541), .ZN(n7597) );
  INV_X1 U6511 ( .A(n8746), .ZN(n4522) );
  NAND3_X1 U6512 ( .A1(n4819), .A2(n5202), .A3(n4524), .ZN(n4519) );
  NAND2_X1 U6513 ( .A1(n4521), .A2(n4520), .ZN(n8702) );
  AOI21_X1 U6514 ( .B1(n8797), .B2(n10331), .A(n4824), .ZN(n8905) );
  XNOR2_X1 U6515 ( .A(n8533), .B(n8534), .ZN(n8797) );
  NAND2_X1 U6516 ( .A1(n8010), .A2(n4536), .ZN(n4534) );
  NAND2_X1 U6517 ( .A1(n5786), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n4555) );
  NAND2_X1 U6518 ( .A1(n6282), .A2(n4414), .ZN(n4561) );
  OAI211_X1 U6519 ( .C1(n6282), .C2(n4566), .A(n4562), .B(n4561), .ZN(n10080)
         );
  XNOR2_X1 U6520 ( .A(n4573), .B(n4572), .ZN(n8152) );
  INV_X1 U6521 ( .A(n5793), .ZN(n4572) );
  NAND2_X1 U6522 ( .A1(n5779), .A2(n5778), .ZN(n4574) );
  NAND2_X1 U6523 ( .A1(n4580), .A2(n4290), .ZN(n4575) );
  NAND2_X1 U6524 ( .A1(n4580), .A2(n4931), .ZN(n5676) );
  OAI21_X2 U6525 ( .B1(n4580), .B2(n4578), .A(n4576), .ZN(n5705) );
  NAND3_X1 U6526 ( .A1(n4599), .A2(n4608), .A3(n6724), .ZN(n4598) );
  INV_X1 U6527 ( .A(n6725), .ZN(n4609) );
  NAND2_X1 U6528 ( .A1(n8685), .A2(n4618), .ZN(n6700) );
  INV_X1 U6529 ( .A(n7540), .ZN(n7599) );
  OAI21_X1 U6530 ( .B1(n7335), .B2(n7538), .A(n6641), .ZN(n7598) );
  NAND2_X1 U6531 ( .A1(n7576), .A2(n6629), .ZN(n6353) );
  NAND2_X1 U6532 ( .A1(n5161), .A2(n5159), .ZN(n7576) );
  INV_X1 U6533 ( .A(n6292), .ZN(n4630) );
  NAND2_X1 U6534 ( .A1(n6292), .A2(n4375), .ZN(n4629) );
  NAND2_X1 U6535 ( .A1(n4630), .A2(n4628), .ZN(n4627) );
  AND2_X1 U6536 ( .A1(n5129), .A2(n4634), .ZN(n4631) );
  OAI21_X2 U6537 ( .B1(n7891), .B2(n4635), .A(n4633), .ZN(n7958) );
  INV_X1 U6538 ( .A(n8695), .ZN(n4637) );
  OAI22_X1 U6539 ( .A1(n5139), .A2(n4645), .B1(n5135), .B2(n8734), .ZN(n4646)
         );
  NAND2_X1 U6540 ( .A1(n4759), .A2(n4646), .ZN(n8557) );
  NAND2_X1 U6541 ( .A1(n4650), .A2(n4652), .ZN(n8147) );
  NAND3_X1 U6542 ( .A1(n4377), .A2(n10352), .A3(n4656), .ZN(n4650) );
  NAND2_X1 U6543 ( .A1(n4651), .A2(n4654), .ZN(n8151) );
  NAND3_X1 U6544 ( .A1(n4377), .A2(n10345), .A3(n4656), .ZN(n4651) );
  NAND2_X1 U6545 ( .A1(n5104), .A2(n5103), .ZN(n8355) );
  NAND2_X2 U6546 ( .A1(n4663), .A2(n5112), .ZN(n6872) );
  NAND2_X1 U6547 ( .A1(n4664), .A2(n4384), .ZN(n4663) );
  NAND2_X1 U6548 ( .A1(n4665), .A2(n4666), .ZN(n4664) );
  NAND3_X1 U6549 ( .A1(n5104), .A2(n5103), .A3(n6856), .ZN(n4665) );
  NAND2_X1 U6550 ( .A1(n6798), .A2(n4672), .ZN(n4670) );
  NAND2_X1 U6551 ( .A1(n4670), .A2(n4671), .ZN(n7656) );
  NAND3_X1 U6552 ( .A1(n6145), .A2(n6144), .A3(n4379), .ZN(n6613) );
  NAND2_X1 U6553 ( .A1(n8519), .A2(n6740), .ZN(n8140) );
  NAND2_X2 U6554 ( .A1(n8599), .A2(n8598), .ZN(n8582) );
  NAND2_X1 U6555 ( .A1(n4684), .A2(n4685), .ZN(n6369) );
  AOI21_X2 U6556 ( .B1(n7947), .B2(n6008), .A(n6007), .ZN(n8039) );
  NAND2_X1 U6557 ( .A1(n4686), .A2(n4690), .ZN(n9060) );
  OR2_X1 U6558 ( .A1(n8999), .A2(n8998), .ZN(n9028) );
  OAI21_X1 U6559 ( .B1(n4702), .B2(n4321), .A(n6055), .ZN(n4696) );
  NAND3_X1 U6560 ( .A1(n5058), .A2(n4699), .A3(n8992), .ZN(n4697) );
  NAND3_X1 U6561 ( .A1(n5058), .A2(n8992), .A3(n4284), .ZN(n4703) );
  INV_X1 U6562 ( .A(n5891), .ZN(n4711) );
  OAI21_X1 U6563 ( .B1(n9021), .B2(n9019), .A(n9017), .ZN(n9090) );
  OAI21_X1 U6564 ( .B1(n5062), .B2(n9121), .A(n5059), .ZN(n7707) );
  NAND2_X1 U6565 ( .A1(n7707), .A2(n7706), .ZN(n5992) );
  NAND2_X1 U6566 ( .A1(n9099), .A2(n9100), .ZN(n9098) );
  OAI21_X1 U6567 ( .B1(n7408), .B2(n5957), .A(n5956), .ZN(n9121) );
  NAND2_X1 U6568 ( .A1(n7139), .A2(n7138), .ZN(n7137) );
  AOI21_X1 U6569 ( .B1(n5964), .B2(n5968), .A(n5064), .ZN(n5063) );
  OAI21_X1 U6570 ( .B1(n9081), .B2(n9077), .A(n9078), .ZN(n9021) );
  NAND2_X1 U6571 ( .A1(n5033), .A2(n5031), .ZN(n8983) );
  OAI21_X2 U6572 ( .B1(n5724), .B2(n5723), .A(n5722), .ZN(n5739) );
  XNOR2_X1 U6573 ( .A(n4712), .B(n7344), .ZN(n6627) );
  NAND4_X1 U6574 ( .A1(n6753), .A2(n5226), .A3(n6754), .A4(n8130), .ZN(n4712)
         );
  NAND2_X1 U6575 ( .A1(n4774), .A2(n5307), .ZN(n5318) );
  NOR2_X1 U6576 ( .A1(n6757), .A2(n6748), .ZN(n6753) );
  INV_X1 U6577 ( .A(n5356), .ZN(n4713) );
  OAI21_X1 U6578 ( .B1(n6760), .B2(n7759), .A(n5155), .ZN(n5154) );
  NAND2_X1 U6579 ( .A1(n4714), .A2(n9064), .ZN(P1_U3227) );
  OAI21_X1 U6580 ( .B1(n9058), .B2(n4715), .A(n9145), .ZN(n4714) );
  NOR2_X2 U6581 ( .A1(n9060), .A2(n9059), .ZN(n9058) );
  NAND2_X1 U6582 ( .A1(n9666), .A2(n5851), .ZN(n9641) );
  AND2_X1 U6583 ( .A1(n5924), .A2(n5923), .ZN(n9099) );
  NAND2_X2 U6584 ( .A1(n4719), .A2(n4718), .ZN(n8992) );
  NAND2_X2 U6585 ( .A1(n8990), .A2(n8989), .ZN(n5058) );
  NOR2_X1 U6586 ( .A1(n4739), .A2(n4738), .ZN(n4737) );
  NAND2_X1 U6587 ( .A1(n5992), .A2(n4386), .ZN(n7875) );
  NAND2_X1 U6588 ( .A1(n7875), .A2(n6000), .ZN(n7947) );
  NAND2_X1 U6589 ( .A1(n5809), .A2(n4332), .ZN(n4721) );
  NAND2_X4 U6590 ( .A1(n6113), .A2(n5903), .ZN(n7522) );
  INV_X1 U6591 ( .A(n9402), .ZN(n7425) );
  NAND2_X1 U6592 ( .A1(n5950), .A2(n9065), .ZN(n7408) );
  INV_X1 U6593 ( .A(n6756), .ZN(n4901) );
  NAND2_X1 U6594 ( .A1(n4788), .A2(n4743), .ZN(n9619) );
  INV_X1 U6595 ( .A(n4800), .ZN(n4799) );
  NAND2_X1 U6596 ( .A1(n5425), .A2(n5424), .ZN(n5445) );
  INV_X1 U6597 ( .A(n7441), .ZN(n9459) );
  NAND2_X1 U6598 ( .A1(n9763), .A2(n9765), .ZN(n5843) );
  NAND2_X1 U6599 ( .A1(n5141), .A2(n6537), .ZN(n5139) );
  NAND2_X1 U6600 ( .A1(n9805), .A2(n9252), .ZN(n9260) );
  NAND3_X1 U6601 ( .A1(n9440), .A2(n9439), .A3(n4747), .ZN(n4746) );
  NAND2_X1 U6602 ( .A1(n10080), .A2(n9253), .ZN(n4733) );
  NAND2_X1 U6603 ( .A1(n9433), .A2(n9432), .ZN(n9436) );
  NOR2_X1 U6604 ( .A1(n9438), .A2(n9437), .ZN(n9439) );
  NAND2_X1 U6605 ( .A1(n6755), .A2(n6742), .ZN(n4903) );
  NOR2_X1 U6606 ( .A1(n9269), .A2(n9267), .ZN(n4872) );
  NAND2_X1 U6607 ( .A1(n4734), .A2(n4896), .ZN(n4902) );
  NAND2_X1 U6608 ( .A1(n4897), .A2(n4898), .ZN(n4734) );
  NAND2_X1 U6609 ( .A1(n4758), .A2(n4757), .ZN(n4756) );
  NAND2_X1 U6610 ( .A1(n5134), .A2(n5225), .ZN(n4755) );
  NAND3_X1 U6611 ( .A1(n6747), .A2(n6746), .A3(n8785), .ZN(n4735) );
  NAND2_X2 U6612 ( .A1(n5628), .A2(n4737), .ZN(n5893) );
  NAND2_X1 U6613 ( .A1(n6430), .A2(n6429), .ZN(n7996) );
  INV_X1 U6614 ( .A(n6310), .ZN(n6304) );
  NAND2_X1 U6615 ( .A1(n8144), .A2(n6588), .ZN(n4741) );
  AOI21_X1 U6616 ( .B1(n7737), .B2(n7738), .A(n6364), .ZN(n7552) );
  NAND2_X1 U6617 ( .A1(n7837), .A2(n6663), .ZN(n7892) );
  NAND3_X1 U6618 ( .A1(n6321), .A2(n6320), .A3(n4742), .ZN(n10272) );
  NAND2_X1 U6619 ( .A1(n9570), .A2(n9569), .ZN(n9824) );
  NAND2_X2 U6620 ( .A1(n9597), .A2(n9596), .ZN(n9595) );
  OAI211_X1 U6621 ( .C1(n9753), .C2(n9827), .A(n4782), .B(n4780), .ZN(n10055)
         );
  NAND2_X1 U6622 ( .A1(n5120), .A2(n6893), .ZN(n8158) );
  AOI21_X1 U6623 ( .B1(n5106), .B2(n5109), .A(n4393), .ZN(n5103) );
  NAND2_X1 U6624 ( .A1(n8258), .A2(n6843), .ZN(n4744) );
  NAND2_X1 U6625 ( .A1(n6844), .A2(n8263), .ZN(n4745) );
  NAND2_X1 U6626 ( .A1(n4869), .A2(n4867), .ZN(n4866) );
  NOR2_X1 U6627 ( .A1(n9229), .A2(n4886), .ZN(n4885) );
  NAND2_X1 U6628 ( .A1(n4893), .A2(n4902), .ZN(n6760) );
  NAND2_X1 U6629 ( .A1(n5730), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5266) );
  NAND2_X1 U6630 ( .A1(n6752), .A2(n4899), .ZN(n4898) );
  OAI21_X1 U6631 ( .B1(n4921), .B2(n4919), .A(n4918), .ZN(n6747) );
  NAND2_X1 U6632 ( .A1(n5096), .A2(n5095), .ZN(n5094) );
  NAND2_X1 U6633 ( .A1(n4752), .A2(n4751), .ZN(P2_U3231) );
  NAND2_X1 U6634 ( .A1(n4763), .A2(n4761), .ZN(n4752) );
  NAND2_X1 U6635 ( .A1(n6794), .A2(n8279), .ZN(n8272) );
  OR2_X1 U6636 ( .A1(n5931), .A2(n5930), .ZN(n5932) );
  NOR2_X1 U6637 ( .A1(n9271), .A2(n9270), .ZN(n4871) );
  OAI211_X1 U6638 ( .C1(n4869), .C2(n4868), .A(n4866), .B(n4865), .ZN(P1_U3240) );
  NAND2_X1 U6639 ( .A1(n5739), .A2(n5737), .ZN(n4954) );
  INV_X1 U6640 ( .A(n6753), .ZN(n4758) );
  OAI211_X1 U6641 ( .C1(n4897), .C2(n6917), .A(n6759), .B(n4894), .ZN(n4893)
         );
  NAND2_X1 U6642 ( .A1(n6760), .A2(n6761), .ZN(n5157) );
  NAND2_X1 U6643 ( .A1(n4954), .A2(n4959), .ZN(n5779) );
  NAND2_X1 U6644 ( .A1(n5705), .A2(n5704), .ZN(n5707) );
  NAND3_X1 U6645 ( .A1(n8789), .A2(n5218), .A3(n8790), .ZN(n8903) );
  AOI21_X2 U6646 ( .B1(n8112), .B2(n10290), .A(n8111), .ZN(n8789) );
  INV_X1 U6647 ( .A(n8555), .ZN(n8125) );
  INV_X1 U6648 ( .A(n5135), .ZN(n5134) );
  NAND2_X1 U6649 ( .A1(n7475), .A2(n5833), .ZN(n7526) );
  NAND2_X1 U6650 ( .A1(n8582), .A2(n6537), .ZN(n5140) );
  NAND2_X1 U6651 ( .A1(n6375), .A2(n4382), .ZN(n7837) );
  NAND2_X1 U6652 ( .A1(n4762), .A2(n6878), .ZN(n4761) );
  INV_X1 U6653 ( .A(n8301), .ZN(n4762) );
  OAI22_X1 U6654 ( .A1(n8301), .A2(n8377), .B1(n8299), .B2(n8353), .ZN(n4763)
         );
  INV_X4 U6655 ( .A(n6884), .ZN(n6793) );
  NAND2_X1 U6656 ( .A1(n5157), .A2(n6764), .ZN(n5156) );
  NAND2_X1 U6657 ( .A1(n4764), .A2(n9145), .ZN(n4784) );
  OAI21_X1 U6658 ( .B1(n9058), .B2(n4765), .A(n9033), .ZN(n4764) );
  NAND2_X1 U6659 ( .A1(n5318), .A2(n5319), .ZN(n4767) );
  XNOR2_X1 U6660 ( .A(n4768), .B(n7522), .ZN(n5940) );
  INV_X1 U6661 ( .A(n5934), .ZN(n4768) );
  MUX2_X1 U6662 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n9858), .S(n7161), .Z(n7154)
         );
  NAND2_X1 U6663 ( .A1(n6072), .A2(n6071), .ZN(n5046) );
  NAND2_X1 U6664 ( .A1(n5305), .A2(n5304), .ZN(n4774) );
  NOR2_X1 U6665 ( .A1(n5863), .A2(n4777), .ZN(n4792) );
  NAND2_X2 U6666 ( .A1(n4298), .A2(n5268), .ZN(n7323) );
  INV_X1 U6667 ( .A(n5063), .ZN(n5062) );
  INV_X1 U6668 ( .A(n5980), .ZN(n5064) );
  NAND2_X1 U6669 ( .A1(n4792), .A2(n4793), .ZN(n6770) );
  NAND2_X1 U6670 ( .A1(n9619), .A2(n9342), .ZN(n9597) );
  NOR2_X1 U6671 ( .A1(n9334), .A2(n5176), .ZN(n5174) );
  AND3_X1 U6672 ( .A1(n5291), .A2(n5292), .A3(n5293), .ZN(n4853) );
  NAND2_X1 U6673 ( .A1(n4933), .A2(n5641), .ZN(n5660) );
  XNOR2_X2 U6674 ( .A(n5185), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5184) );
  NAND2_X1 U6675 ( .A1(n5049), .A2(n5048), .ZN(n5047) );
  NAND2_X1 U6676 ( .A1(n4784), .A2(n4783), .ZN(P1_U3223) );
  INV_X1 U6677 ( .A(n5154), .ZN(n5153) );
  NAND2_X1 U6678 ( .A1(n7426), .A2(n7425), .ZN(n7424) );
  NAND2_X1 U6679 ( .A1(n4793), .A2(n5821), .ZN(n9537) );
  AOI21_X1 U6680 ( .B1(n4794), .B2(n4797), .A(n4795), .ZN(n5244) );
  NAND2_X1 U6681 ( .A1(n9595), .A2(n9343), .ZN(n4814) );
  INV_X1 U6682 ( .A(n4814), .ZN(n9587) );
  INV_X1 U6683 ( .A(n9236), .ZN(n4813) );
  NAND3_X1 U6684 ( .A1(n9401), .A2(n9402), .A3(n9398), .ZN(n7421) );
  OAI21_X1 U6685 ( .B1(n8626), .B2(n4828), .A(n4391), .ZN(n8588) );
  NOR2_X1 U6686 ( .A1(n8922), .A2(n8223), .ZN(n4838) );
  MUX2_X1 U6687 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9962), .S(n7031), .Z(n7020)
         );
  NAND3_X1 U6688 ( .A1(n4855), .A2(n9222), .A3(n4854), .ZN(n9228) );
  NAND3_X1 U6689 ( .A1(n9213), .A2(n4857), .A3(n4856), .ZN(n4855) );
  AND2_X1 U6690 ( .A1(n4858), .A2(n4381), .ZN(n4857) );
  OR2_X1 U6691 ( .A1(n4862), .A2(n4859), .ZN(n4858) );
  NAND3_X1 U6692 ( .A1(n9275), .A2(n9276), .A3(n9277), .ZN(n4868) );
  NOR3_X2 U6693 ( .A1(n4872), .A2(n4871), .A3(n4870), .ZN(n4869) );
  AOI21_X1 U6694 ( .B1(n9210), .B2(n9711), .A(n9331), .ZN(n9212) );
  AOI21_X2 U6695 ( .B1(n4873), .B2(n9208), .A(n9207), .ZN(n9210) );
  AND2_X1 U6696 ( .A1(n9362), .A2(n9174), .ZN(n4876) );
  NAND3_X1 U6697 ( .A1(n9247), .A2(n9248), .A3(n9427), .ZN(n4884) );
  NAND2_X1 U6698 ( .A1(n6998), .A2(n4889), .ZN(n4888) );
  NAND3_X1 U6699 ( .A1(n6693), .A2(n8700), .A3(n4892), .ZN(n4891) );
  NAND2_X1 U6700 ( .A1(n6752), .A2(n4895), .ZN(n4894) );
  OR2_X1 U6701 ( .A1(n6682), .A2(n4906), .ZN(n4904) );
  NAND2_X1 U6702 ( .A1(n4904), .A2(n4905), .ZN(n6692) );
  NAND2_X1 U6703 ( .A1(n6684), .A2(n6640), .ZN(n4913) );
  NAND3_X1 U6704 ( .A1(n4929), .A2(n4928), .A3(P1_DATAO_REG_3__SCAN_IN), .ZN(
        n4926) );
  NAND2_X1 U6705 ( .A1(n5565), .A2(n4946), .ZN(n4941) );
  NAND2_X1 U6706 ( .A1(n5724), .A2(n4952), .ZN(n4951) );
  INV_X1 U6707 ( .A(n5722), .ZN(n4953) );
  NAND3_X1 U6708 ( .A1(n4969), .A2(n4964), .A3(n4416), .ZN(P2_U3264) );
  NAND2_X1 U6709 ( .A1(n4965), .A2(n7344), .ZN(n4964) );
  NAND2_X1 U6710 ( .A1(n4968), .A2(n4966), .ZN(n4965) );
  NAND2_X1 U6711 ( .A1(n6272), .A2(n10256), .ZN(n4968) );
  OAI22_X1 U6712 ( .A1(n6272), .A2(n10259), .B1(n10261), .B2(n6271), .ZN(n4970) );
  NOR2_X1 U6713 ( .A1(n4990), .A2(n4983), .ZN(n4980) );
  NAND2_X1 U6714 ( .A1(n4982), .A2(n4987), .ZN(n8467) );
  NAND3_X1 U6715 ( .A1(n5012), .A2(n5011), .A3(n5009), .ZN(P1_U3260) );
  NAND2_X1 U6716 ( .A1(n5015), .A2(n9071), .ZN(n7435) );
  NAND2_X1 U6717 ( .A1(n9697), .A2(n4304), .ZN(n9650) );
  NOR3_X2 U6718 ( .A1(n5216), .A2(n5020), .A3(n9734), .ZN(n5022) );
  INV_X1 U6719 ( .A(n5022), .ZN(n9732) );
  NAND2_X1 U6720 ( .A1(n9581), .A2(n4380), .ZN(n8056) );
  NOR2_X2 U6721 ( .A1(n5327), .A2(n5241), .ZN(n5810) );
  INV_X2 U6722 ( .A(n5327), .ZN(n5028) );
  NAND2_X1 U6723 ( .A1(n9033), .A2(n6089), .ZN(n9133) );
  NAND2_X1 U6724 ( .A1(n9033), .A2(n5034), .ZN(n5033) );
  INV_X1 U6725 ( .A(n6108), .ZN(n6107) );
  OAI21_X1 U6726 ( .B1(n9098), .B2(n5038), .A(n5037), .ZN(n9067) );
  AOI21_X1 U6727 ( .B1(n5043), .B2(n7374), .A(n4317), .ZN(n5037) );
  INV_X1 U6728 ( .A(n7374), .ZN(n5038) );
  NAND2_X1 U6729 ( .A1(n5041), .A2(n5039), .ZN(n5950) );
  INV_X1 U6730 ( .A(n5040), .ZN(n5039) );
  OAI21_X1 U6731 ( .B1(n7374), .B2(n4317), .A(n9066), .ZN(n5040) );
  NAND2_X1 U6732 ( .A1(n9098), .A2(n5042), .ZN(n5041) );
  NOR2_X1 U6733 ( .A1(n5043), .A2(n4317), .ZN(n5042) );
  NAND2_X1 U6734 ( .A1(n5865), .A2(n4378), .ZN(n5044) );
  XNOR2_X1 U6735 ( .A(n5045), .B(P1_IR_REG_23__SCAN_IN), .ZN(n7755) );
  NAND2_X1 U6736 ( .A1(n9090), .A2(n9087), .ZN(n5049) );
  NAND3_X1 U6737 ( .A1(n5047), .A2(n5046), .A3(n5052), .ZN(n5051) );
  NAND2_X1 U6738 ( .A1(n5051), .A2(n5050), .ZN(n6085) );
  INV_X1 U6739 ( .A(n5058), .ZN(n8993) );
  OAI21_X1 U6740 ( .B1(n4753), .B2(n5964), .A(n5968), .ZN(n7773) );
  AND3_X2 U6741 ( .A1(n4309), .A2(n7940), .A3(n7747), .ZN(n8747) );
  NAND2_X1 U6742 ( .A1(n4309), .A2(n7747), .ZN(n5067) );
  INV_X1 U6743 ( .A(n5067), .ZN(n7937) );
  AND2_X2 U6744 ( .A1(n8612), .A2(n5068), .ZN(n8574) );
  INV_X1 U6745 ( .A(n5073), .ZN(n8589) );
  NAND2_X1 U6746 ( .A1(n8542), .A2(n5075), .ZN(n8503) );
  NAND2_X1 U6747 ( .A1(n8542), .A2(n4302), .ZN(n8501) );
  OAI21_X1 U6748 ( .B1(n7859), .B2(n5837), .A(n5836), .ZN(n7762) );
  NAND2_X1 U6749 ( .A1(n5837), .A2(n5836), .ZN(n5102) );
  NAND2_X1 U6750 ( .A1(n8260), .A2(n5106), .ZN(n5104) );
  OAI21_X1 U6751 ( .B1(n4725), .B2(n6846), .A(n6845), .ZN(n8286) );
  XNOR2_X2 U6752 ( .A(n6872), .B(n6870), .ZN(n8342) );
  NAND2_X1 U6753 ( .A1(n6888), .A2(n5118), .ZN(n5117) );
  NAND2_X1 U6754 ( .A1(n6888), .A2(n5123), .ZN(n5120) );
  NAND2_X1 U6755 ( .A1(n6888), .A2(n8247), .ZN(n8365) );
  NAND2_X1 U6756 ( .A1(n6318), .A2(n5133), .ZN(n6633) );
  NAND2_X1 U6757 ( .A1(n6778), .A2(n5133), .ZN(n7594) );
  OAI22_X1 U6758 ( .A1(n10328), .A2(n8063), .B1(n10326), .B2(n5133), .ZN(n7345) );
  NOR2_X1 U6759 ( .A1(n8104), .A2(n7609), .ZN(n5150) );
  XNOR2_X1 U6760 ( .A(n6610), .B(n7344), .ZN(n5158) );
  OAI21_X1 U6761 ( .B1(n5158), .B2(n5156), .A(n5153), .ZN(P2_U3244) );
  NOR2_X1 U6762 ( .A1(n6645), .A2(n5160), .ZN(n5159) );
  NAND2_X1 U6763 ( .A1(n7996), .A2(n5162), .ZN(n6442) );
  INV_X1 U6764 ( .A(n8629), .ZN(n5166) );
  NAND2_X1 U6765 ( .A1(n5443), .A2(n5168), .ZN(n5167) );
  AOI21_X1 U6766 ( .B1(n5180), .B2(n5178), .A(n5367), .ZN(n7520) );
  NAND2_X1 U6767 ( .A1(n5189), .A2(n9831), .ZN(n10056) );
  XNOR2_X1 U6768 ( .A(n9587), .B(n4272), .ZN(n5188) );
  OAI21_X1 U6769 ( .B1(n9832), .B2(n9753), .A(n9830), .ZN(n5190) );
  NAND4_X1 U6770 ( .A1(n6144), .A2(n6163), .A3(n6145), .A4(n4390), .ZN(n6292)
         );
  INV_X1 U6771 ( .A(n9826), .ZN(n9154) );
  INV_X1 U6772 ( .A(n5257), .ZN(n5265) );
  OR2_X1 U6773 ( .A1(n6943), .A2(n6942), .ZN(n6996) );
  AND2_X1 U6774 ( .A1(n5910), .A2(n5909), .ZN(n7139) );
  NAND2_X1 U6775 ( .A1(n6633), .A2(n6641), .ZN(n7538) );
  NAND2_X1 U6776 ( .A1(n8564), .A2(n8574), .ZN(n8558) );
  NAND2_X1 U6777 ( .A1(n6290), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6247) );
  NAND2_X1 U6778 ( .A1(n9565), .A2(n9799), .ZN(n9570) );
  CLKBUF_X1 U6779 ( .A(n8695), .Z(n8696) );
  XNOR2_X1 U6780 ( .A(n5865), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9302) );
  OR2_X2 U6781 ( .A1(n7718), .A2(n6615), .ZN(n6640) );
  NAND2_X1 U6782 ( .A1(n6615), .A2(n7344), .ZN(n6626) );
  XNOR2_X1 U6783 ( .A(n6245), .B(n6244), .ZN(n6264) );
  XNOR2_X1 U6784 ( .A(n6884), .B(n10285), .ZN(n6775) );
  NAND2_X1 U6785 ( .A1(n6636), .A2(n10288), .ZN(n10293) );
  AND2_X1 U6786 ( .A1(n8811), .A2(n8550), .ZN(n8569) );
  INV_X1 U6787 ( .A(n9747), .ZN(n5562) );
  OR2_X1 U6788 ( .A1(n10245), .A2(n5804), .ZN(n5211) );
  OR2_X1 U6789 ( .A1(n10254), .A2(n5899), .ZN(n5212) );
  AND2_X1 U6790 ( .A1(n5814), .A2(n9274), .ZN(n9767) );
  INV_X1 U6791 ( .A(n9767), .ZN(n9799) );
  INV_X1 U6792 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n6133) );
  INV_X1 U6793 ( .A(n9566), .ZN(n9447) );
  AND2_X1 U6794 ( .A1(n8125), .A2(n5214), .ZN(n5213) );
  AND2_X1 U6795 ( .A1(n8568), .A2(n8550), .ZN(n5214) );
  NOR2_X1 U6796 ( .A1(n9728), .A2(n5823), .ZN(n5215) );
  OR2_X2 U6797 ( .A1(n8015), .A2(n7951), .ZN(n5216) );
  NOR2_X1 U6798 ( .A1(n5480), .A2(n5479), .ZN(n5217) );
  OR2_X1 U6799 ( .A1(n8788), .A2(n8778), .ZN(n5218) );
  NOR2_X1 U6800 ( .A1(n9611), .A2(n9610), .ZN(n5219) );
  AND2_X1 U6801 ( .A1(n6106), .A2(n9145), .ZN(n5220) );
  AND3_X1 U6802 ( .A1(n6338), .A2(n6337), .A3(n6336), .ZN(n5221) );
  INV_X1 U6803 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5322) );
  AND2_X1 U6804 ( .A1(n5524), .A2(n5512), .ZN(n5222) );
  INV_X1 U6805 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n5361) );
  INV_X1 U6806 ( .A(n9770), .ZN(n9796) );
  INV_X1 U6807 ( .A(n8420), .ZN(n6340) );
  INV_X1 U6808 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5466) );
  AND2_X1 U6809 ( .A1(n8127), .A2(n8126), .ZN(n5223) );
  AND4_X1 U6810 ( .A1(n8785), .A2(n8536), .A3(n8520), .A4(n6625), .ZN(n5226)
         );
  INV_X1 U6811 ( .A(n7993), .ZN(n6429) );
  AND2_X1 U6812 ( .A1(n8641), .A2(n6498), .ZN(n5227) );
  INV_X1 U6813 ( .A(n8619), .ZN(n6515) );
  NAND2_X1 U6814 ( .A1(n9984), .A2(n9448), .ZN(n5228) );
  INV_X1 U6815 ( .A(n9358), .ZN(n5368) );
  INV_X1 U6816 ( .A(n7834), .ZN(n6385) );
  NAND2_X1 U6817 ( .A1(n5236), .A2(n5235), .ZN(n5237) );
  OR2_X1 U6818 ( .A1(n10236), .A2(n7780), .ZN(n9174) );
  INV_X1 U6819 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6376) );
  INV_X1 U6820 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6293) );
  OR2_X1 U6821 ( .A1(n9006), .A2(n9110), .ZN(n6049) );
  XNOR2_X1 U6822 ( .A(n5927), .B(n6059), .ZN(n5931) );
  NAND2_X1 U6823 ( .A1(n7082), .A2(n7458), .ZN(n7083) );
  INV_X1 U6824 ( .A(SI_12_), .ZN(n5486) );
  INV_X1 U6825 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5375) );
  INV_X1 U6826 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5239) );
  INV_X1 U6827 ( .A(n7643), .ZN(n6807) );
  INV_X1 U6828 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n6404) );
  INV_X1 U6829 ( .A(n6345), .ZN(n6542) );
  INV_X1 U6830 ( .A(n6332), .ZN(n6561) );
  AND2_X1 U6831 ( .A1(n8027), .A2(n8028), .ZN(n8429) );
  INV_X1 U6832 ( .A(n8383), .ZN(n8324) );
  INV_X1 U6833 ( .A(n8542), .ZN(n8526) );
  INV_X1 U6834 ( .A(n6607), .ZN(n6485) );
  NAND2_X1 U6835 ( .A1(n6148), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6166) );
  OAI21_X1 U6836 ( .B1(n6053), .B2(n6052), .A(n9008), .ZN(n6054) );
  NOR2_X1 U6837 ( .A1(n9263), .A2(n9770), .ZN(n8052) );
  NOR2_X1 U6838 ( .A1(n9567), .A2(n9772), .ZN(n9568) );
  INV_X1 U6839 ( .A(SI_15_), .ZN(n9921) );
  INV_X1 U6840 ( .A(n8059), .ZN(n9814) );
  INV_X1 U6841 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5242) );
  NAND2_X1 U6842 ( .A1(n5678), .A2(n5677), .ZN(n5687) );
  NAND2_X1 U6843 ( .A1(n5627), .A2(n5626), .ZN(n5628) );
  NAND2_X1 U6844 ( .A1(n5544), .A2(n9921), .ZN(n5563) );
  INV_X1 U6845 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7976) );
  OR2_X1 U6846 ( .A1(n8491), .A2(n6276), .ZN(n6278) );
  INV_X1 U6847 ( .A(n8571), .ZN(n8568) );
  INV_X1 U6848 ( .A(n8598), .ZN(n8596) );
  OR2_X1 U6849 ( .A1(n8926), .A2(n8407), .ZN(n8122) );
  OR2_X1 U6850 ( .A1(n10276), .A2(n7933), .ZN(n7722) );
  AND2_X1 U6851 ( .A1(n10302), .A2(n10307), .ZN(n6914) );
  INV_X1 U6852 ( .A(n7547), .ZN(n7551) );
  NAND2_X1 U6853 ( .A1(n6166), .A2(n6165), .ZN(n6168) );
  INV_X1 U6854 ( .A(n6054), .ZN(n6055) );
  INV_X1 U6855 ( .A(n7873), .ZN(n5997) );
  AND2_X1 U6856 ( .A1(n6122), .A2(n6121), .ZN(n9146) );
  INV_X1 U6857 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7791) );
  OR2_X1 U6858 ( .A1(n7084), .A2(n9435), .ZN(n6109) );
  AND2_X1 U6859 ( .A1(n7088), .A2(n9435), .ZN(n10033) );
  INV_X1 U6860 ( .A(n9794), .ZN(n9772) );
  OR2_X1 U6861 ( .A1(n5816), .A2(n9279), .ZN(n9770) );
  AND2_X1 U6862 ( .A1(n5776), .A2(n5743), .ZN(n5756) );
  NAND2_X1 U6863 ( .A1(n5563), .A2(n5546), .ZN(n5564) );
  AND2_X1 U6864 ( .A1(n7312), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8372) );
  OR2_X1 U6865 ( .A1(n10303), .A2(n7328), .ZN(n10279) );
  AOI21_X1 U6866 ( .B1(n6250), .B2(P2_REG2_REG_1__SCAN_IN), .A(n7153), .ZN(
        n7166) );
  INV_X1 U6867 ( .A(n10256), .ZN(n10259) );
  AND2_X1 U6868 ( .A1(n6266), .A2(n6265), .ZN(n10256) );
  INV_X1 U6869 ( .A(n10328), .ZN(n8892) );
  INV_X1 U6870 ( .A(n8520), .ZN(n8517) );
  INV_X1 U6871 ( .A(n10281), .ZN(n8766) );
  NAND2_X1 U6872 ( .A1(n10270), .A2(n7722), .ZN(n10284) );
  NOR2_X1 U6873 ( .A1(n10308), .A2(n6914), .ZN(n7715) );
  AND2_X1 U6874 ( .A1(n6908), .A2(n6907), .ZN(n10302) );
  INV_X1 U6875 ( .A(n9146), .ZN(n9134) );
  INV_X1 U6876 ( .A(n5336), .ZN(n5820) );
  AND2_X1 U6877 ( .A1(n5640), .A2(n5639), .ZN(n9112) );
  INV_X1 U6878 ( .A(n10182), .ZN(n10143) );
  INV_X1 U6879 ( .A(n10132), .ZN(n10190) );
  AND2_X1 U6880 ( .A1(n9516), .A2(n5815), .ZN(n10188) );
  NAND2_X1 U6881 ( .A1(n9230), .A2(n4813), .ZN(n9588) );
  AND2_X1 U6882 ( .A1(n6944), .A2(n9279), .ZN(n9794) );
  OR2_X1 U6883 ( .A1(n6111), .A2(n6110), .ZN(n9755) );
  INV_X1 U6884 ( .A(n10047), .ZN(n10237) );
  AND2_X1 U6885 ( .A1(n6111), .A2(n7415), .ZN(n6769) );
  AND2_X1 U6886 ( .A1(n5495), .A2(n5526), .ZN(n9467) );
  NAND2_X1 U6887 ( .A1(n4271), .A2(n5274), .ZN(n5272) );
  OR3_X1 U6888 ( .A1(n7925), .A2(n8023), .A3(n8978), .ZN(n6934) );
  INV_X1 U6889 ( .A(n8491), .ZN(n10258) );
  INV_X1 U6890 ( .A(n6939), .ZN(n6940) );
  INV_X1 U6891 ( .A(n8823), .ZN(n8618) );
  AND2_X1 U6892 ( .A1(n6918), .A2(n10279), .ZN(n8364) );
  NAND2_X1 U6893 ( .A1(n6266), .A2(n8969), .ZN(n10260) );
  INV_X1 U6894 ( .A(n10286), .ZN(n8754) );
  OR2_X1 U6895 ( .A1(n10276), .A2(n7721), .ZN(n10270) );
  INV_X1 U6896 ( .A(n8873), .ZN(n8885) );
  INV_X1 U6897 ( .A(n8543), .ZN(n8907) );
  INV_X1 U6898 ( .A(n8739), .ZN(n8943) );
  NOR2_X1 U6899 ( .A1(n10303), .A2(n10302), .ZN(n10306) );
  INV_X1 U6900 ( .A(n10306), .ZN(n10309) );
  INV_X1 U6901 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7924) );
  INV_X1 U6902 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n9928) );
  INV_X1 U6903 ( .A(n8960), .ZN(n8977) );
  INV_X1 U6904 ( .A(n9828), .ZN(n9586) );
  INV_X1 U6905 ( .A(n7920), .ZN(n7980) );
  NAND2_X1 U6906 ( .A1(n7292), .A2(n6105), .ZN(n9140) );
  INV_X1 U6907 ( .A(n9617), .ZN(n9589) );
  INV_X1 U6908 ( .A(n9722), .ZN(n9694) );
  OR2_X1 U6909 ( .A1(P1_U3083), .A2(n6997), .ZN(n10195) );
  NAND2_X1 U6910 ( .A1(n10209), .A2(n10208), .ZN(n9783) );
  INV_X1 U6911 ( .A(n9802), .ZN(n9762) );
  AND2_X2 U6912 ( .A1(n5898), .A2(n6769), .ZN(n10254) );
  AND2_X2 U6913 ( .A1(n7417), .A2(n6769), .ZN(n10245) );
  INV_X1 U6914 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9908) );
  INV_X1 U6915 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7587) );
  INV_X1 U6916 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7120) );
  NOR2_X1 U6917 ( .A1(n10390), .A2(n10389), .ZN(n10388) );
  NOR2_X1 U6918 ( .A1(n10380), .A2(n10379), .ZN(n10378) );
  NOR2_X1 U6919 ( .A1(n6996), .A2(P1_U3084), .ZN(P1_U4006) );
  NOR2_X1 U6920 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5231) );
  NOR2_X2 U6921 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5624) );
  NOR2_X1 U6922 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5230) );
  NAND2_X1 U6923 ( .A1(n5786), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5249) );
  NAND2_X1 U6924 ( .A1(n5730), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5248) );
  NAND2_X1 U6925 ( .A1(n5311), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5247) );
  NAND2_X1 U6926 ( .A1(n5336), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5246) );
  AND4_X2 U6927 ( .A1(n5249), .A2(n5248), .A3(n5247), .A4(n5246), .ZN(n7087)
         );
  INV_X1 U6928 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6954) );
  INV_X1 U6929 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5256) );
  NAND2_X1 U6930 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5255) );
  OAI22_X1 U6931 ( .A1(n9255), .A2(n6954), .B1(n6998), .B2(n7067), .ZN(n5257)
         );
  AND2_X1 U6932 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5274) );
  NAND2_X1 U6933 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5280) );
  INV_X1 U6934 ( .A(n5280), .ZN(n5258) );
  INV_X1 U6935 ( .A(SI_1_), .ZN(n5260) );
  XNOR2_X1 U6936 ( .A(n5261), .B(n5260), .ZN(n5263) );
  MUX2_X1 U6937 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n4271), .Z(n5262) );
  XNOR2_X1 U6938 ( .A(n5263), .B(n5262), .ZN(n6955) );
  OR2_X1 U6939 ( .A1(n5317), .A2(n6955), .ZN(n5264) );
  NAND2_X1 U6940 ( .A1(n7087), .A2(n5858), .ZN(n7297) );
  NAND2_X1 U6941 ( .A1(n5311), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5269) );
  NAND2_X1 U6942 ( .A1(n5786), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5268) );
  NAND2_X1 U6943 ( .A1(n5336), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5267) );
  INV_X1 U6944 ( .A(SI_0_), .ZN(n5271) );
  INV_X1 U6945 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5270) );
  OAI21_X1 U6946 ( .B1(n6950), .B2(n5271), .A(n5270), .ZN(n5273) );
  AND2_X1 U6947 ( .A1(n5273), .A2(n5272), .ZN(n10095) );
  MUX2_X1 U6948 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10095), .S(n6998), .Z(n7458)
         );
  NAND2_X1 U6949 ( .A1(n7297), .A2(n7083), .ZN(n9401) );
  INV_X1 U6950 ( .A(n5858), .ZN(n5916) );
  NOR2_X1 U6951 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(SI_1_), .ZN(n5277) );
  INV_X1 U6952 ( .A(n5274), .ZN(n5276) );
  NAND2_X1 U6953 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(SI_1_), .ZN(n5275) );
  OAI21_X1 U6954 ( .B1(n5277), .B2(n5276), .A(n5275), .ZN(n5278) );
  NAND2_X1 U6955 ( .A1(n4271), .A2(n5278), .ZN(n5284) );
  NOR2_X1 U6956 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5281) );
  NAND2_X1 U6957 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5279) );
  OAI21_X1 U6958 ( .B1(n5281), .B2(n5280), .A(n5279), .ZN(n5282) );
  INV_X1 U6959 ( .A(n5282), .ZN(n5283) );
  INV_X1 U6960 ( .A(SI_2_), .ZN(n5302) );
  XNOR2_X1 U6961 ( .A(n5304), .B(n5302), .ZN(n5286) );
  MUX2_X1 U6962 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n4271), .Z(n5285) );
  XNOR2_X1 U6963 ( .A(n5286), .B(n5285), .ZN(n6957) );
  OR2_X1 U6964 ( .A1(n5317), .A2(n6957), .ZN(n5290) );
  INV_X1 U6965 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6956) );
  INV_X1 U6966 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5287) );
  NAND2_X1 U6967 ( .A1(n5288), .A2(n5287), .ZN(n5299) );
  OR2_X1 U6968 ( .A1(n6998), .A2(n7123), .ZN(n5289) );
  NAND2_X1 U6969 ( .A1(n5311), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5293) );
  NAND2_X1 U6970 ( .A1(n5336), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5292) );
  NAND2_X1 U6971 ( .A1(n4283), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5291) );
  NAND2_X1 U6972 ( .A1(n4554), .A2(n9102), .ZN(n9304) );
  NAND2_X1 U6973 ( .A1(n5786), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5298) );
  NAND2_X1 U6974 ( .A1(n4283), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5297) );
  NAND2_X1 U6975 ( .A1(n5336), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5296) );
  INV_X1 U6976 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5294) );
  NAND2_X1 U6977 ( .A1(n5311), .A2(n5294), .ZN(n5295) );
  INV_X1 U6978 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5300) );
  INV_X1 U6979 ( .A(SI_3_), .ZN(n5301) );
  XNOR2_X1 U6980 ( .A(n5320), .B(n5301), .ZN(n5319) );
  INV_X1 U6981 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6948) );
  NAND2_X1 U6982 ( .A1(n4271), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5303) );
  OAI211_X1 U6983 ( .C1(n4271), .C2(n6948), .A(n5303), .B(n5302), .ZN(n5305)
         );
  NAND2_X1 U6984 ( .A1(n4271), .A2(n6956), .ZN(n5306) );
  OAI211_X1 U6985 ( .C1(n4271), .C2(P1_DATAO_REG_2__SCAN_IN), .A(n5306), .B(
        SI_2_), .ZN(n5307) );
  XNOR2_X1 U6986 ( .A(n5318), .B(n5319), .ZN(n6962) );
  OR2_X1 U6987 ( .A1(n6962), .A2(n5317), .ZN(n5309) );
  OR2_X1 U6988 ( .A1(n4282), .A2(n4927), .ZN(n5308) );
  OAI211_X2 U6989 ( .C1(n6998), .C2(n7031), .A(n5309), .B(n5308), .ZN(n7387)
         );
  INV_X2 U6990 ( .A(n7387), .ZN(n7485) );
  NAND2_X1 U6991 ( .A1(n9459), .A2(n7485), .ZN(n9306) );
  NAND2_X1 U6992 ( .A1(n7441), .A2(n7387), .ZN(n9356) );
  NAND2_X1 U6993 ( .A1(n9365), .A2(n9404), .ZN(n5310) );
  INV_X1 U6994 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5312) );
  XNOR2_X1 U6995 ( .A(n5312), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n9072) );
  NAND2_X1 U6996 ( .A1(n5311), .A2(n9072), .ZN(n5316) );
  NAND2_X1 U6997 ( .A1(n4283), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5315) );
  NAND2_X1 U6998 ( .A1(n5786), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5314) );
  NAND2_X1 U6999 ( .A1(n5336), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5313) );
  NAND2_X1 U7000 ( .A1(n5320), .A2(SI_3_), .ZN(n5321) );
  XNOR2_X1 U7001 ( .A(n5355), .B(n5342), .ZN(n6951) );
  NAND2_X1 U7002 ( .A1(n9253), .A2(n6951), .ZN(n5331) );
  NAND2_X1 U7003 ( .A1(n5325), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5326) );
  MUX2_X1 U7004 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5326), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5328) );
  NAND2_X1 U7005 ( .A1(n5328), .A2(n5327), .ZN(n7181) );
  OR2_X1 U7006 ( .A1(n6998), .A2(n7181), .ZN(n5330) );
  INV_X1 U7007 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6953) );
  OR2_X1 U7008 ( .A1(n4282), .A2(n6953), .ZN(n5329) );
  NAND2_X1 U7009 ( .A1(n4283), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5340) );
  NAND2_X1 U7010 ( .A1(n5786), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5339) );
  INV_X1 U7011 ( .A(n5332), .ZN(n5334) );
  INV_X1 U7012 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5333) );
  NAND2_X1 U7013 ( .A1(n5334), .A2(n5333), .ZN(n5335) );
  AND2_X1 U7014 ( .A1(n5349), .A2(n5335), .ZN(n10200) );
  NAND2_X1 U7015 ( .A1(n5311), .A2(n10200), .ZN(n5338) );
  NAND2_X1 U7016 ( .A1(n5336), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5337) );
  INV_X2 U7017 ( .A(n4282), .ZN(n5631) );
  NAND2_X1 U7018 ( .A1(n5327), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5341) );
  XNOR2_X1 U7019 ( .A(n5341), .B(P1_IR_REG_5__SCAN_IN), .ZN(n7054) );
  AOI22_X1 U7020 ( .A1(n5631), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6946), .B2(
        n7054), .ZN(n5347) );
  INV_X1 U7021 ( .A(n5342), .ZN(n5343) );
  NAND2_X1 U7022 ( .A1(n5355), .A2(n5343), .ZN(n5344) );
  NAND2_X1 U7023 ( .A1(n5357), .A2(SI_4_), .ZN(n5356) );
  NAND2_X1 U7024 ( .A1(n5344), .A2(n5356), .ZN(n5345) );
  MUX2_X1 U7025 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n4271), .Z(n5359) );
  XNOR2_X1 U7026 ( .A(n5345), .B(n5358), .ZN(n6958) );
  NAND2_X1 U7027 ( .A1(n6958), .A2(n9253), .ZN(n5346) );
  NAND2_X1 U7028 ( .A1(n7471), .A2(n10198), .ZN(n9161) );
  INV_X1 U7029 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7109) );
  NAND2_X1 U7030 ( .A1(n5349), .A2(n7109), .ZN(n5350) );
  AND2_X1 U7031 ( .A1(n5382), .A2(n5350), .ZN(n9126) );
  NAND2_X1 U7032 ( .A1(n5311), .A2(n9126), .ZN(n5354) );
  NAND2_X1 U7033 ( .A1(n5786), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5353) );
  NAND2_X1 U7034 ( .A1(n5336), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5352) );
  NAND2_X1 U7035 ( .A1(n4283), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5351) );
  NAND2_X1 U7036 ( .A1(n5359), .A2(SI_5_), .ZN(n5388) );
  XNOR2_X1 U7037 ( .A(n5392), .B(SI_6_), .ZN(n5369) );
  NAND2_X1 U7038 ( .A1(n6965), .A2(n9253), .ZN(n5365) );
  NAND2_X1 U7039 ( .A1(n5028), .A2(n5362), .ZN(n5374) );
  NAND2_X1 U7040 ( .A1(n5374), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5363) );
  XNOR2_X1 U7041 ( .A(n5363), .B(P1_IR_REG_6__SCAN_IN), .ZN(n7040) );
  AOI22_X1 U7042 ( .A1(n5631), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6946), .B2(
        n7040), .ZN(n5364) );
  NAND2_X1 U7043 ( .A1(n7636), .A2(n9123), .ZN(n9167) );
  NAND2_X1 U7044 ( .A1(n9161), .A2(n9167), .ZN(n9358) );
  INV_X1 U7045 ( .A(n7471), .ZN(n9457) );
  INV_X1 U7046 ( .A(n10198), .ZN(n7409) );
  NAND2_X1 U7047 ( .A1(n9167), .A2(n5830), .ZN(n5366) );
  INV_X1 U7048 ( .A(n7636), .ZN(n9456) );
  NAND2_X1 U7049 ( .A1(n10229), .A2(n9456), .ZN(n9171) );
  AND2_X1 U7050 ( .A1(n5366), .A2(n9171), .ZN(n9363) );
  INV_X1 U7051 ( .A(n5369), .ZN(n5370) );
  NAND2_X1 U7052 ( .A1(n5371), .A2(n5370), .ZN(n5372) );
  NAND2_X1 U7053 ( .A1(n5392), .A2(SI_6_), .ZN(n5389) );
  NAND2_X1 U7054 ( .A1(n5372), .A2(n5389), .ZN(n5373) );
  NAND2_X1 U7055 ( .A1(n6973), .A2(n9253), .ZN(n5379) );
  INV_X1 U7056 ( .A(n5374), .ZN(n5376) );
  NAND2_X1 U7057 ( .A1(n5376), .A2(n5375), .ZN(n5404) );
  NAND2_X1 U7058 ( .A1(n5404), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5377) );
  XNOR2_X1 U7059 ( .A(n5377), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7096) );
  AOI22_X1 U7060 ( .A1(n5631), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6946), .B2(
        n7096), .ZN(n5378) );
  NAND2_X1 U7061 ( .A1(n5786), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5387) );
  NAND2_X1 U7062 ( .A1(n4283), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5386) );
  INV_X1 U7063 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5381) );
  NAND2_X1 U7064 ( .A1(n5382), .A2(n5381), .ZN(n5383) );
  AND2_X1 U7065 ( .A1(n5411), .A2(n5383), .ZN(n7634) );
  NAND2_X1 U7066 ( .A1(n5311), .A2(n7634), .ZN(n5385) );
  NAND2_X1 U7067 ( .A1(n5336), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5384) );
  OR2_X1 U7068 ( .A1(n7698), .A2(n7794), .ZN(n9362) );
  NAND2_X1 U7069 ( .A1(n7698), .A2(n7794), .ZN(n9166) );
  NAND2_X1 U7070 ( .A1(n7520), .A2(n9410), .ZN(n7683) );
  NAND2_X1 U7071 ( .A1(n5389), .A2(n5388), .ZN(n5421) );
  INV_X1 U7072 ( .A(n5421), .ZN(n5390) );
  NAND2_X1 U7073 ( .A1(n5423), .A2(n5390), .ZN(n5395) );
  INV_X1 U7074 ( .A(n5391), .ZN(n5394) );
  NAND2_X1 U7075 ( .A1(n5395), .A2(n5422), .ZN(n5397) );
  NAND2_X1 U7076 ( .A1(n5396), .A2(SI_7_), .ZN(n5419) );
  NAND2_X1 U7077 ( .A1(n5397), .A2(n5419), .ZN(n5403) );
  INV_X1 U7078 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6972) );
  INV_X1 U7079 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5398) );
  MUX2_X1 U7080 ( .A(n6972), .B(n5398), .S(n4271), .Z(n5400) );
  INV_X1 U7081 ( .A(SI_8_), .ZN(n5399) );
  NAND2_X1 U7082 ( .A1(n5400), .A2(n5399), .ZN(n5424) );
  INV_X1 U7083 ( .A(n5400), .ZN(n5401) );
  NAND2_X1 U7084 ( .A1(n5401), .A2(SI_8_), .ZN(n5402) );
  NAND2_X1 U7085 ( .A1(n5424), .A2(n5402), .ZN(n5418) );
  NAND2_X1 U7086 ( .A1(n6960), .A2(n9253), .ZN(n5410) );
  NAND2_X1 U7087 ( .A1(n5407), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5406) );
  MUX2_X1 U7088 ( .A(n5406), .B(P1_IR_REG_31__SCAN_IN), .S(n5405), .Z(n5408)
         );
  AOI22_X1 U7089 ( .A1(n5631), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6946), .B2(
        n10125), .ZN(n5409) );
  NAND2_X1 U7090 ( .A1(n4283), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5416) );
  NAND2_X1 U7091 ( .A1(n5786), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5415) );
  NAND2_X1 U7092 ( .A1(n5411), .A2(n7791), .ZN(n5412) );
  AND2_X1 U7093 ( .A1(n5437), .A2(n5412), .ZN(n7792) );
  NAND2_X1 U7094 ( .A1(n5311), .A2(n7792), .ZN(n5414) );
  NAND2_X1 U7095 ( .A1(n5336), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5413) );
  NAND2_X1 U7096 ( .A1(n10236), .A2(n7780), .ZN(n9168) );
  AND2_X1 U7097 ( .A1(n9166), .A2(n9168), .ZN(n9172) );
  NAND2_X1 U7098 ( .A1(n7683), .A2(n9172), .ZN(n5417) );
  NAND2_X1 U7099 ( .A1(n5417), .A2(n9174), .ZN(n7860) );
  INV_X1 U7100 ( .A(n5418), .ZN(n5420) );
  INV_X1 U7101 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6978) );
  INV_X1 U7102 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5426) );
  MUX2_X1 U7103 ( .A(n6978), .B(n5426), .S(n4271), .Z(n5428) );
  INV_X1 U7104 ( .A(SI_9_), .ZN(n5427) );
  NAND2_X1 U7105 ( .A1(n5428), .A2(n5427), .ZN(n5462) );
  INV_X1 U7106 ( .A(n5428), .ZN(n5429) );
  NAND2_X1 U7107 ( .A1(n5429), .A2(SI_9_), .ZN(n5430) );
  XNOR2_X1 U7108 ( .A(n5445), .B(n5444), .ZN(n6969) );
  NAND2_X1 U7109 ( .A1(n6969), .A2(n9253), .ZN(n5434) );
  NAND2_X1 U7110 ( .A1(n5431), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5432) );
  AOI22_X1 U7111 ( .A1(n5631), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6946), .B2(
        n7266), .ZN(n5433) );
  NAND2_X1 U7112 ( .A1(n4283), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5442) );
  NAND2_X1 U7113 ( .A1(n5786), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5441) );
  INV_X1 U7114 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U7115 ( .A1(n5437), .A2(n5436), .ZN(n5438) );
  AND2_X1 U7116 ( .A1(n5455), .A2(n5438), .ZN(n7779) );
  NAND2_X1 U7117 ( .A1(n5311), .A2(n7779), .ZN(n5440) );
  NAND2_X1 U7118 ( .A1(n5336), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5439) );
  NAND2_X1 U7119 ( .A1(n10048), .A2(n7858), .ZN(n9296) );
  NAND2_X1 U7120 ( .A1(n7860), .A2(n9296), .ZN(n5443) );
  OR2_X1 U7121 ( .A1(n10048), .A2(n7858), .ZN(n9175) );
  NAND2_X1 U7122 ( .A1(n5482), .A2(n5462), .ZN(n5450) );
  INV_X1 U7123 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6982) );
  INV_X1 U7124 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6980) );
  MUX2_X1 U7125 ( .A(n6982), .B(n6980), .S(n4271), .Z(n5447) );
  INV_X1 U7126 ( .A(SI_10_), .ZN(n5446) );
  NAND2_X1 U7127 ( .A1(n5447), .A2(n5446), .ZN(n5461) );
  INV_X1 U7128 ( .A(n5447), .ZN(n5448) );
  AND2_X1 U7129 ( .A1(n5461), .A2(n5479), .ZN(n5449) );
  NAND2_X1 U7130 ( .A1(n6979), .A2(n9253), .ZN(n5453) );
  OR2_X1 U7131 ( .A1(n5810), .A2(n5466), .ZN(n5451) );
  XNOR2_X1 U7132 ( .A(n5451), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7357) );
  AOI22_X1 U7133 ( .A1(n5631), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6946), .B2(
        n7357), .ZN(n5452) );
  NAND2_X1 U7134 ( .A1(n5786), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5460) );
  NAND2_X1 U7135 ( .A1(n5336), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U7136 ( .A1(n5455), .A2(n5454), .ZN(n5456) );
  AND2_X1 U7137 ( .A1(n5471), .A2(n5456), .ZN(n7765) );
  NAND2_X1 U7138 ( .A1(n5311), .A2(n7765), .ZN(n5458) );
  NAND2_X1 U7139 ( .A1(n4283), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5457) );
  NAND4_X1 U7140 ( .A1(n5460), .A2(n5459), .A3(n5458), .A4(n5457), .ZN(n9452)
         );
  AND2_X1 U7141 ( .A1(n7767), .A2(n9452), .ZN(n9313) );
  INV_X1 U7142 ( .A(n9452), .ZN(n7878) );
  NAND2_X1 U7143 ( .A1(n10043), .A2(n7878), .ZN(n9297) );
  NAND2_X1 U7144 ( .A1(n5482), .A2(n5477), .ZN(n5463) );
  AND2_X1 U7145 ( .A1(n5463), .A2(n5479), .ZN(n5464) );
  XNOR2_X1 U7146 ( .A(n5464), .B(n5478), .ZN(n6988) );
  NAND2_X1 U7147 ( .A1(n6988), .A2(n9253), .ZN(n5469) );
  INV_X1 U7148 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5465) );
  OR2_X1 U7149 ( .A1(n5491), .A2(n5466), .ZN(n5467) );
  XNOR2_X1 U7150 ( .A(n5467), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7614) );
  AOI22_X1 U7151 ( .A1(n5631), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6946), .B2(
        n7614), .ZN(n5468) );
  NAND2_X1 U7152 ( .A1(n4283), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5476) );
  NAND2_X1 U7153 ( .A1(n5786), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5475) );
  INV_X1 U7154 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U7155 ( .A1(n5471), .A2(n5470), .ZN(n5472) );
  AND2_X1 U7156 ( .A1(n5499), .A2(n5472), .ZN(n7877) );
  NAND2_X1 U7157 ( .A1(n5311), .A2(n7877), .ZN(n5474) );
  NAND2_X1 U7158 ( .A1(n5336), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5473) );
  AND2_X1 U7159 ( .A1(n7920), .A2(n8009), .ZN(n9187) );
  OR2_X1 U7160 ( .A1(n7920), .A2(n8009), .ZN(n9184) );
  OAI21_X1 U7161 ( .B1(n7913), .B2(n9187), .A(n9184), .ZN(n8008) );
  INV_X1 U7162 ( .A(n5478), .ZN(n5480) );
  INV_X1 U7163 ( .A(n5483), .ZN(n5484) );
  MUX2_X1 U7164 ( .A(n9844), .B(n5485), .S(n4271), .Z(n5487) );
  INV_X1 U7165 ( .A(n5487), .ZN(n5488) );
  NAND2_X1 U7166 ( .A1(n5488), .A2(SI_12_), .ZN(n5489) );
  NAND2_X1 U7167 ( .A1(n6992), .A2(n9253), .ZN(n5497) );
  NAND2_X1 U7168 ( .A1(n5491), .A2(n5490), .ZN(n5493) );
  NAND2_X1 U7169 ( .A1(n5493), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5492) );
  MUX2_X1 U7170 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5492), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n5495) );
  AOI22_X1 U7171 ( .A1(n5631), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6946), .B2(
        n9467), .ZN(n5496) );
  NAND2_X1 U7172 ( .A1(n5786), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5504) );
  NAND2_X1 U7173 ( .A1(n5336), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5503) );
  NAND2_X1 U7174 ( .A1(n5499), .A2(n5498), .ZN(n5500) );
  AND2_X1 U7175 ( .A1(n5517), .A2(n5500), .ZN(n8017) );
  NAND2_X1 U7176 ( .A1(n5311), .A2(n8017), .ZN(n5502) );
  NAND2_X1 U7177 ( .A1(n4283), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5501) );
  NAND4_X1 U7178 ( .A1(n5504), .A2(n5503), .A3(n5502), .A4(n5501), .ZN(n9795)
         );
  AND2_X1 U7179 ( .A1(n10040), .A2(n9795), .ZN(n9190) );
  INV_X1 U7180 ( .A(n9190), .ZN(n5505) );
  INV_X1 U7181 ( .A(n9795), .ZN(n6001) );
  NAND2_X1 U7182 ( .A1(n7951), .A2(n6001), .ZN(n9189) );
  MUX2_X1 U7183 ( .A(n7013), .B(n7010), .S(n4271), .Z(n5510) );
  INV_X1 U7184 ( .A(SI_13_), .ZN(n5509) );
  INV_X1 U7185 ( .A(n5510), .ZN(n5511) );
  NAND2_X1 U7186 ( .A1(n5511), .A2(SI_13_), .ZN(n5512) );
  XNOR2_X1 U7187 ( .A(n5523), .B(n5222), .ZN(n7009) );
  NAND2_X1 U7188 ( .A1(n7009), .A2(n9253), .ZN(n5515) );
  NAND2_X1 U7189 ( .A1(n5526), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5513) );
  XNOR2_X1 U7190 ( .A(n5513), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9471) );
  AOI22_X1 U7191 ( .A1(n5631), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6946), .B2(
        n9471), .ZN(n5514) );
  NAND2_X1 U7192 ( .A1(n5786), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5522) );
  NAND2_X1 U7193 ( .A1(n5336), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5521) );
  NAND2_X1 U7194 ( .A1(n5517), .A2(n5516), .ZN(n5518) );
  AND2_X1 U7195 ( .A1(n5530), .A2(n5518), .ZN(n9787) );
  NAND2_X1 U7196 ( .A1(n5311), .A2(n9787), .ZN(n5520) );
  NAND2_X1 U7197 ( .A1(n4283), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5519) );
  OR2_X1 U7198 ( .A1(n10032), .A2(n9771), .ZN(n9196) );
  NAND2_X1 U7199 ( .A1(n10032), .A2(n9771), .ZN(n9764) );
  MUX2_X1 U7200 ( .A(n7064), .B(n7061), .S(n4271), .Z(n5539) );
  XNOR2_X1 U7201 ( .A(n5543), .B(n5538), .ZN(n7060) );
  NAND2_X1 U7202 ( .A1(n7060), .A2(n9253), .ZN(n5528) );
  OR2_X1 U7203 ( .A1(n5572), .A2(n5466), .ZN(n5548) );
  XNOR2_X1 U7204 ( .A(n5548), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9472) );
  AOI22_X1 U7205 ( .A1(n9472), .A2(n6946), .B1(n5631), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n5527) );
  INV_X1 U7206 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5529) );
  NAND2_X1 U7207 ( .A1(n5530), .A2(n5529), .ZN(n5531) );
  NAND2_X1 U7208 ( .A1(n5555), .A2(n5531), .ZN(n9775) );
  OR2_X1 U7209 ( .A1(n9775), .A2(n5801), .ZN(n5535) );
  NAND2_X1 U7210 ( .A1(n5786), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5534) );
  NAND2_X1 U7211 ( .A1(n5336), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5533) );
  NAND2_X1 U7212 ( .A1(n4283), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5532) );
  NAND2_X1 U7213 ( .A1(n10029), .A2(n8045), .ZN(n9294) );
  NAND2_X1 U7214 ( .A1(n9198), .A2(n9294), .ZN(n9765) );
  INV_X1 U7215 ( .A(n9764), .ZN(n9314) );
  NOR2_X1 U7216 ( .A1(n9765), .A2(n9314), .ZN(n5536) );
  NAND2_X1 U7217 ( .A1(n9791), .A2(n5536), .ZN(n5537) );
  INV_X1 U7218 ( .A(n5539), .ZN(n5540) );
  NAND2_X1 U7219 ( .A1(n5540), .A2(SI_14_), .ZN(n5541) );
  MUX2_X1 U7220 ( .A(n7122), .B(n7120), .S(n4271), .Z(n5544) );
  INV_X1 U7221 ( .A(n5544), .ZN(n5545) );
  NAND2_X1 U7222 ( .A1(n5545), .A2(SI_15_), .ZN(n5546) );
  NAND2_X1 U7223 ( .A1(n7119), .A2(n9253), .ZN(n5552) );
  INV_X1 U7224 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5547) );
  NAND2_X1 U7225 ( .A1(n5548), .A2(n5547), .ZN(n5549) );
  NAND2_X1 U7226 ( .A1(n5549), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5550) );
  XNOR2_X1 U7227 ( .A(n5550), .B(P1_IR_REG_15__SCAN_IN), .ZN(n10163) );
  AOI22_X1 U7228 ( .A1(n10163), .A2(n6946), .B1(n5631), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n5551) );
  INV_X1 U7229 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5554) );
  NAND2_X1 U7230 ( .A1(n5555), .A2(n5554), .ZN(n5556) );
  NAND2_X1 U7231 ( .A1(n5577), .A2(n5556), .ZN(n9756) );
  OR2_X1 U7232 ( .A1(n9756), .A2(n5801), .ZN(n5561) );
  NAND2_X1 U7233 ( .A1(n5786), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5558) );
  NAND2_X1 U7234 ( .A1(n4283), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5557) );
  AND2_X1 U7235 ( .A1(n5558), .A2(n5557), .ZN(n5560) );
  NAND2_X1 U7236 ( .A1(n5336), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5559) );
  OR2_X1 U7237 ( .A1(n9759), .A2(n9769), .ZN(n9321) );
  NAND2_X1 U7238 ( .A1(n9759), .A2(n9769), .ZN(n9295) );
  NAND2_X1 U7239 ( .A1(n9321), .A2(n9295), .ZN(n9747) );
  MUX2_X1 U7240 ( .A(n7190), .B(n5566), .S(n4271), .Z(n5568) );
  INV_X1 U7241 ( .A(SI_16_), .ZN(n5567) );
  NAND2_X1 U7242 ( .A1(n5568), .A2(n5567), .ZN(n5581) );
  INV_X1 U7243 ( .A(n5568), .ZN(n5569) );
  NAND2_X1 U7244 ( .A1(n5569), .A2(SI_16_), .ZN(n5570) );
  NAND2_X1 U7245 ( .A1(n7148), .A2(n9253), .ZN(n5575) );
  NOR2_X1 U7246 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5571) );
  NAND2_X1 U7247 ( .A1(n5572), .A2(n5571), .ZN(n5627) );
  NAND2_X1 U7248 ( .A1(n5627), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5573) );
  XNOR2_X1 U7249 ( .A(n5573), .B(P1_IR_REG_16__SCAN_IN), .ZN(n10175) );
  AOI22_X1 U7250 ( .A1(n10175), .A2(n6946), .B1(n5631), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n5574) );
  INV_X1 U7251 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5576) );
  NAND2_X1 U7252 ( .A1(n5577), .A2(n5576), .ZN(n5578) );
  NAND2_X1 U7253 ( .A1(n5605), .A2(n5578), .ZN(n9719) );
  AOI22_X1 U7254 ( .A1(n5336), .A2(P1_REG0_REG_16__SCAN_IN), .B1(n5786), .B2(
        P1_REG1_REG_16__SCAN_IN), .ZN(n5580) );
  NAND2_X1 U7255 ( .A1(n4283), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5579) );
  OAI211_X1 U7256 ( .C1(n9719), .C2(n5801), .A(n5580), .B(n5579), .ZN(n9750)
         );
  INV_X1 U7257 ( .A(n9750), .ZN(n9147) );
  NAND2_X1 U7258 ( .A1(n9734), .A2(n9147), .ZN(n9205) );
  INV_X1 U7259 ( .A(n5581), .ZN(n5582) );
  MUX2_X1 U7260 ( .A(n9928), .B(n7310), .S(n4271), .Z(n5593) );
  XNOR2_X1 U7261 ( .A(n5593), .B(SI_17_), .ZN(n5592) );
  NAND2_X1 U7262 ( .A1(n7307), .A2(n9253), .ZN(n5586) );
  OR2_X1 U7263 ( .A1(n5627), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n5584) );
  NAND2_X1 U7264 ( .A1(n5584), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5597) );
  XNOR2_X1 U7265 ( .A(n5597), .B(P1_IR_REG_17__SCAN_IN), .ZN(n10187) );
  AOI22_X1 U7266 ( .A1(n10187), .A2(n6946), .B1(n5631), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n5585) );
  XNOR2_X1 U7267 ( .A(n5605), .B(P1_REG3_REG_17__SCAN_IN), .ZN(n9709) );
  NAND2_X1 U7268 ( .A1(n9709), .A2(n5311), .ZN(n5591) );
  INV_X1 U7269 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9489) );
  NAND2_X1 U7270 ( .A1(n4283), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U7271 ( .A1(n5336), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5587) );
  OAI211_X1 U7272 ( .C1(n4785), .C2(n9489), .A(n5588), .B(n5587), .ZN(n5589)
         );
  INV_X1 U7273 ( .A(n5589), .ZN(n5590) );
  AND2_X1 U7274 ( .A1(n10010), .A2(n9722), .ZN(n9209) );
  INV_X1 U7275 ( .A(n5593), .ZN(n5594) );
  INV_X1 U7276 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n5595) );
  MUX2_X1 U7277 ( .A(n5595), .B(n7382), .S(n5690), .Z(n5614) );
  XNOR2_X1 U7278 ( .A(n5613), .B(n4475), .ZN(n7349) );
  NAND2_X1 U7279 ( .A1(n7349), .A2(n9253), .ZN(n5601) );
  INV_X1 U7280 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5596) );
  NAND2_X1 U7281 ( .A1(n5597), .A2(n5596), .ZN(n5598) );
  NAND2_X1 U7282 ( .A1(n5598), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5599) );
  XNOR2_X1 U7283 ( .A(n5599), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9511) );
  AOI22_X1 U7284 ( .A1(n9511), .A2(n6946), .B1(n5631), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n5600) );
  AND2_X1 U7285 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_REG3_REG_18__SCAN_IN), 
        .ZN(n5602) );
  INV_X1 U7286 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5604) );
  INV_X1 U7287 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5603) );
  OAI21_X1 U7288 ( .B1(n5605), .B2(n5604), .A(n5603), .ZN(n5606) );
  NAND2_X1 U7289 ( .A1(n5634), .A2(n5606), .ZN(n9701) );
  OR2_X1 U7290 ( .A1(n9701), .A2(n5801), .ZN(n5611) );
  INV_X1 U7291 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9514) );
  NAND2_X1 U7292 ( .A1(n4283), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5608) );
  NAND2_X1 U7293 ( .A1(n5336), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5607) );
  OAI211_X1 U7294 ( .C1(n4785), .C2(n9514), .A(n5608), .B(n5607), .ZN(n5609)
         );
  INV_X1 U7295 ( .A(n5609), .ZN(n5610) );
  OR2_X1 U7296 ( .A1(n10010), .A2(n9722), .ZN(n9690) );
  NAND2_X1 U7297 ( .A1(n9214), .A2(n9690), .ZN(n9331) );
  NAND2_X1 U7298 ( .A1(n10004), .A2(n9054), .ZN(n9215) );
  INV_X1 U7299 ( .A(n5614), .ZN(n5615) );
  NAND2_X1 U7300 ( .A1(n5615), .A2(SI_18_), .ZN(n5616) );
  MUX2_X1 U7301 ( .A(n9943), .B(n7465), .S(n4271), .Z(n5619) );
  INV_X1 U7302 ( .A(SI_19_), .ZN(n5618) );
  INV_X1 U7303 ( .A(n5619), .ZN(n5620) );
  NAND2_X1 U7304 ( .A1(n5620), .A2(SI_19_), .ZN(n5621) );
  NOR2_X1 U7305 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5622) );
  AND2_X1 U7306 ( .A1(n5624), .A2(n5622), .ZN(n5630) );
  XNOR2_X1 U7307 ( .A(P1_IR_REG_31__SCAN_IN), .B(P1_IR_REG_19__SCAN_IN), .ZN(
        n5629) );
  NAND3_X1 U7308 ( .A1(n5624), .A2(P1_IR_REG_19__SCAN_IN), .A3(n5623), .ZN(
        n5625) );
  NOR2_X1 U7309 ( .A1(n5466), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n5626) );
  AOI22_X1 U7310 ( .A1(n5893), .A2(n6946), .B1(n5631), .B2(
        P2_DATAO_REG_19__SCAN_IN), .ZN(n5632) );
  NAND2_X2 U7311 ( .A1(n5633), .A2(n5632), .ZN(n9999) );
  INV_X1 U7312 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9934) );
  NAND2_X1 U7313 ( .A1(n5634), .A2(n9934), .ZN(n5635) );
  AND2_X1 U7314 ( .A1(n5651), .A2(n5635), .ZN(n9012) );
  NAND2_X1 U7315 ( .A1(n9012), .A2(n5311), .ZN(n5640) );
  INV_X1 U7316 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9515) );
  NAND2_X1 U7317 ( .A1(n4283), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5637) );
  NAND2_X1 U7318 ( .A1(n5336), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5636) );
  OAI211_X1 U7319 ( .C1(n4785), .C2(n9515), .A(n5637), .B(n5636), .ZN(n5638)
         );
  INV_X1 U7320 ( .A(n5638), .ZN(n5639) );
  OR2_X1 U7321 ( .A1(n9999), .A2(n9112), .ZN(n9333) );
  NAND2_X1 U7322 ( .A1(n9999), .A2(n9112), .ZN(n9293) );
  MUX2_X1 U7323 ( .A(n9938), .B(n7519), .S(n5690), .Z(n5645) );
  INV_X1 U7324 ( .A(SI_20_), .ZN(n5644) );
  INV_X1 U7325 ( .A(n5645), .ZN(n5646) );
  NAND2_X1 U7326 ( .A1(n5646), .A2(SI_20_), .ZN(n5647) );
  NAND2_X1 U7327 ( .A1(n7518), .A2(n9253), .ZN(n5649) );
  OR2_X1 U7328 ( .A1(n4282), .A2(n7519), .ZN(n5648) );
  INV_X1 U7329 ( .A(n5651), .ZN(n5650) );
  INV_X1 U7330 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9082) );
  NAND2_X1 U7331 ( .A1(n5651), .A2(n9082), .ZN(n5652) );
  NAND2_X1 U7332 ( .A1(n5664), .A2(n5652), .ZN(n9660) );
  OR2_X1 U7333 ( .A1(n9660), .A2(n5801), .ZN(n5658) );
  INV_X1 U7334 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n5655) );
  NAND2_X1 U7335 ( .A1(n5786), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5654) );
  NAND2_X1 U7336 ( .A1(n4283), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5653) );
  OAI211_X1 U7337 ( .C1(n5655), .C2(n5820), .A(n5654), .B(n5653), .ZN(n5656)
         );
  INV_X1 U7338 ( .A(n5656), .ZN(n5657) );
  NAND2_X1 U7339 ( .A1(n9994), .A2(n9647), .ZN(n9289) );
  MUX2_X1 U7340 ( .A(n7610), .B(n7587), .S(n4271), .Z(n5673) );
  XNOR2_X1 U7341 ( .A(n5676), .B(n5672), .ZN(n7586) );
  NAND2_X1 U7342 ( .A1(n7586), .A2(n9253), .ZN(n5663) );
  OR2_X1 U7343 ( .A1(n4282), .A2(n7587), .ZN(n5662) );
  INV_X1 U7344 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9022) );
  NAND2_X1 U7345 ( .A1(n5664), .A2(n9022), .ZN(n5665) );
  AND2_X1 U7346 ( .A1(n5697), .A2(n5665), .ZN(n9652) );
  NAND2_X1 U7347 ( .A1(n9652), .A2(n5311), .ZN(n5671) );
  INV_X1 U7348 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n5668) );
  NAND2_X1 U7349 ( .A1(n5786), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5667) );
  NAND2_X1 U7350 ( .A1(n4283), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5666) );
  OAI211_X1 U7351 ( .C1(n5668), .C2(n5820), .A(n5667), .B(n5666), .ZN(n5669)
         );
  INV_X1 U7352 ( .A(n5669), .ZN(n5670) );
  XNOR2_X1 U7353 ( .A(n9991), .B(n9220), .ZN(n9640) );
  INV_X1 U7354 ( .A(n5673), .ZN(n5674) );
  MUX2_X1 U7355 ( .A(n8101), .B(n7736), .S(n5690), .Z(n5678) );
  INV_X1 U7356 ( .A(SI_22_), .ZN(n5677) );
  INV_X1 U7357 ( .A(n5678), .ZN(n5679) );
  NAND2_X1 U7358 ( .A1(n5679), .A2(SI_22_), .ZN(n5680) );
  XNOR2_X1 U7359 ( .A(n5689), .B(n5688), .ZN(n7734) );
  NAND2_X1 U7360 ( .A1(n7734), .A2(n9253), .ZN(n5682) );
  OR2_X1 U7361 ( .A1(n4282), .A2(n7736), .ZN(n5681) );
  XNOR2_X1 U7362 ( .A(n5697), .B(P1_REG3_REG_22__SCAN_IN), .ZN(n9633) );
  INV_X1 U7363 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U7364 ( .A1(n5786), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5684) );
  NAND2_X1 U7365 ( .A1(n4283), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5683) );
  OAI211_X1 U7366 ( .C1(n5820), .C2(n5685), .A(n5684), .B(n5683), .ZN(n5686)
         );
  NAND2_X1 U7367 ( .A1(n9984), .A2(n9648), .ZN(n9223) );
  NAND2_X1 U7368 ( .A1(n9991), .A2(n9220), .ZN(n9625) );
  NAND2_X1 U7369 ( .A1(n9223), .A2(n9625), .ZN(n9292) );
  MUX2_X1 U7370 ( .A(n7761), .B(n7757), .S(n4271), .Z(n5691) );
  NAND2_X1 U7371 ( .A1(n5691), .A2(n9838), .ZN(n5706) );
  INV_X1 U7372 ( .A(n5691), .ZN(n5692) );
  NAND2_X1 U7373 ( .A1(n5692), .A2(SI_23_), .ZN(n5693) );
  XNOR2_X1 U7374 ( .A(n5705), .B(n5704), .ZN(n7758) );
  NAND2_X1 U7375 ( .A1(n7758), .A2(n9253), .ZN(n5695) );
  OR2_X1 U7376 ( .A1(n4282), .A2(n7757), .ZN(n5694) );
  AND2_X1 U7377 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(P1_REG3_REG_23__SCAN_IN), 
        .ZN(n5696) );
  INV_X1 U7378 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9091) );
  INV_X1 U7379 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9001) );
  OAI21_X1 U7380 ( .B1(n5697), .B2(n9091), .A(n9001), .ZN(n5698) );
  NAND2_X1 U7381 ( .A1(n5711), .A2(n5698), .ZN(n9612) );
  INV_X1 U7382 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9947) );
  NAND2_X1 U7383 ( .A1(n4283), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5700) );
  NAND2_X1 U7384 ( .A1(n5336), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5699) );
  OAI211_X1 U7385 ( .C1(n4785), .C2(n9947), .A(n5700), .B(n5699), .ZN(n5701)
         );
  INV_X1 U7386 ( .A(n5701), .ZN(n5702) );
  NAND2_X1 U7387 ( .A1(n9980), .A2(n9093), .ZN(n9378) );
  MUX2_X1 U7388 ( .A(n7924), .B(n8083), .S(n5690), .Z(n5720) );
  XNOR2_X1 U7389 ( .A(n5720), .B(SI_24_), .ZN(n5719) );
  NAND2_X1 U7390 ( .A1(n7923), .A2(n9253), .ZN(n5709) );
  OR2_X1 U7391 ( .A1(n4282), .A2(n8083), .ZN(n5708) );
  NAND2_X2 U7392 ( .A1(n5709), .A2(n5708), .ZN(n9977) );
  INV_X1 U7393 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9948) );
  NAND2_X1 U7394 ( .A1(n5711), .A2(n9948), .ZN(n5712) );
  NAND2_X1 U7395 ( .A1(n5747), .A2(n5712), .ZN(n9602) );
  INV_X1 U7396 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n5715) );
  NAND2_X1 U7397 ( .A1(n5786), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5714) );
  NAND2_X1 U7398 ( .A1(n4283), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5713) );
  OAI211_X1 U7399 ( .C1(n5715), .C2(n5820), .A(n5714), .B(n5713), .ZN(n5716)
         );
  INV_X1 U7400 ( .A(n5716), .ZN(n5717) );
  OR2_X2 U7401 ( .A1(n9977), .A2(n9617), .ZN(n9343) );
  NAND2_X1 U7402 ( .A1(n9977), .A2(n9617), .ZN(n9234) );
  INV_X1 U7403 ( .A(n5719), .ZN(n5723) );
  INV_X1 U7404 ( .A(n5720), .ZN(n5721) );
  NAND2_X1 U7405 ( .A1(n5721), .A2(SI_24_), .ZN(n5722) );
  MUX2_X1 U7406 ( .A(n9863), .B(n9930), .S(n4271), .Z(n5725) );
  INV_X1 U7407 ( .A(SI_25_), .ZN(n9895) );
  NAND2_X1 U7408 ( .A1(n5725), .A2(n9895), .ZN(n5737) );
  INV_X1 U7409 ( .A(n5725), .ZN(n5726) );
  NAND2_X1 U7410 ( .A1(n5726), .A2(SI_25_), .ZN(n5727) );
  NAND2_X1 U7411 ( .A1(n5737), .A2(n5727), .ZN(n5738) );
  NAND2_X1 U7412 ( .A1(n8022), .A2(n9253), .ZN(n5729) );
  OR2_X1 U7413 ( .A1(n4282), .A2(n9930), .ZN(n5728) );
  XNOR2_X1 U7414 ( .A(n5747), .B(P1_REG3_REG_25__SCAN_IN), .ZN(n9584) );
  NAND2_X1 U7415 ( .A1(n9584), .A2(n5311), .ZN(n5736) );
  INV_X1 U7416 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n5733) );
  NAND2_X1 U7417 ( .A1(n4283), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5732) );
  NAND2_X1 U7418 ( .A1(n5786), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5731) );
  OAI211_X1 U7419 ( .C1(n5733), .C2(n5820), .A(n5732), .B(n5731), .ZN(n5734)
         );
  INV_X1 U7420 ( .A(n5734), .ZN(n5735) );
  INV_X1 U7421 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8975) );
  MUX2_X1 U7422 ( .A(n8975), .B(n9908), .S(n5690), .Z(n5741) );
  INV_X1 U7423 ( .A(SI_26_), .ZN(n5740) );
  NAND2_X1 U7424 ( .A1(n5741), .A2(n5740), .ZN(n5776) );
  INV_X1 U7425 ( .A(n5741), .ZN(n5742) );
  NAND2_X1 U7426 ( .A1(n5742), .A2(SI_26_), .ZN(n5743) );
  NAND2_X1 U7427 ( .A1(n8049), .A2(n9253), .ZN(n5745) );
  OR2_X1 U7428 ( .A1(n4282), .A2(n9908), .ZN(n5744) );
  INV_X1 U7429 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9034) );
  INV_X1 U7430 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5746) );
  OAI21_X1 U7431 ( .B1(n5747), .B2(n9034), .A(n5746), .ZN(n5748) );
  NAND2_X1 U7432 ( .A1(n9574), .A2(n5311), .ZN(n5754) );
  INV_X1 U7433 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9889) );
  NAND2_X1 U7434 ( .A1(n5786), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5750) );
  NAND2_X1 U7435 ( .A1(n5336), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5749) );
  OAI211_X1 U7436 ( .C1(n5751), .C2(n9889), .A(n5750), .B(n5749), .ZN(n5752)
         );
  INV_X1 U7437 ( .A(n5752), .ZN(n5753) );
  OR2_X1 U7438 ( .A1(n9826), .A2(n9549), .ZN(n5755) );
  NAND2_X1 U7439 ( .A1(n5755), .A2(n9230), .ZN(n9381) );
  NAND2_X1 U7440 ( .A1(n9826), .A2(n9549), .ZN(n9284) );
  INV_X1 U7441 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8973) );
  INV_X1 U7442 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10093) );
  MUX2_X1 U7443 ( .A(n8973), .B(n10093), .S(n5690), .Z(n5759) );
  INV_X1 U7444 ( .A(SI_27_), .ZN(n5758) );
  NAND2_X1 U7445 ( .A1(n5759), .A2(n5758), .ZN(n5775) );
  INV_X1 U7446 ( .A(n5759), .ZN(n5760) );
  NAND2_X1 U7447 ( .A1(n5760), .A2(SI_27_), .ZN(n5777) );
  AND2_X1 U7448 ( .A1(n5775), .A2(n5777), .ZN(n5761) );
  OR2_X1 U7449 ( .A1(n4282), .A2(n10093), .ZN(n5763) );
  INV_X1 U7450 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9896) );
  NAND2_X1 U7451 ( .A1(n5766), .A2(n9896), .ZN(n5767) );
  NAND2_X1 U7452 ( .A1(n5784), .A2(n5767), .ZN(n9553) );
  INV_X1 U7453 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n5770) );
  NAND2_X1 U7454 ( .A1(n5786), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5769) );
  NAND2_X1 U7455 ( .A1(n4283), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5768) );
  OAI211_X1 U7456 ( .C1(n5770), .C2(n5820), .A(n5769), .B(n5768), .ZN(n5771)
         );
  INV_X1 U7457 ( .A(n5771), .ZN(n5772) );
  NAND2_X1 U7458 ( .A1(n9819), .A2(n9566), .ZN(n9287) );
  INV_X1 U7459 ( .A(n9384), .ZN(n5774) );
  AND2_X1 U7460 ( .A1(n5776), .A2(n5775), .ZN(n5778) );
  INV_X1 U7461 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8970) );
  INV_X1 U7462 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8153) );
  MUX2_X1 U7463 ( .A(n8970), .B(n8153), .S(n5690), .Z(n5795) );
  XNOR2_X1 U7464 ( .A(n5795), .B(SI_28_), .ZN(n5793) );
  NAND2_X1 U7465 ( .A1(n8152), .A2(n9253), .ZN(n5781) );
  OR2_X1 U7466 ( .A1(n4282), .A2(n8153), .ZN(n5780) );
  INV_X1 U7467 ( .A(n5784), .ZN(n5782) );
  NAND2_X1 U7468 ( .A1(n5782), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9538) );
  INV_X1 U7469 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5783) );
  NAND2_X1 U7470 ( .A1(n5784), .A2(n5783), .ZN(n5785) );
  NAND2_X1 U7471 ( .A1(n9538), .A2(n5785), .ZN(n8055) );
  INV_X1 U7472 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n5789) );
  NAND2_X1 U7473 ( .A1(n4283), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5788) );
  NAND2_X1 U7474 ( .A1(n5786), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5787) );
  OAI211_X1 U7475 ( .C1(n5789), .C2(n5820), .A(n5788), .B(n5787), .ZN(n5790)
         );
  INV_X1 U7476 ( .A(n5790), .ZN(n5791) );
  NAND2_X1 U7477 ( .A1(n8059), .A2(n9550), .ZN(n9288) );
  NAND2_X1 U7478 ( .A1(n8051), .A2(n9288), .ZN(n5808) );
  INV_X1 U7479 ( .A(SI_28_), .ZN(n5794) );
  NAND2_X1 U7480 ( .A1(n5795), .A2(n5794), .ZN(n5796) );
  INV_X1 U7481 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8966) );
  INV_X1 U7482 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10088) );
  MUX2_X1 U7483 ( .A(n8966), .B(n10088), .S(n4271), .Z(n6279) );
  XNOR2_X1 U7484 ( .A(n6279), .B(SI_29_), .ZN(n5798) );
  NAND2_X1 U7485 ( .A1(n8965), .A2(n9253), .ZN(n5800) );
  OR2_X1 U7486 ( .A1(n4282), .A2(n10088), .ZN(n5799) );
  OR2_X1 U7487 ( .A1(n9538), .A2(n5801), .ZN(n5807) );
  INV_X1 U7488 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5804) );
  NAND2_X1 U7489 ( .A1(n4283), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5803) );
  NAND2_X1 U7490 ( .A1(n5786), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5802) );
  OAI211_X1 U7491 ( .C1(n5804), .C2(n5820), .A(n5803), .B(n5802), .ZN(n5805)
         );
  INV_X1 U7492 ( .A(n5805), .ZN(n5806) );
  NAND2_X1 U7493 ( .A1(n9259), .A2(n9263), .ZN(n9386) );
  INV_X1 U7494 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5870) );
  NAND2_X1 U7495 ( .A1(n5865), .A2(n5870), .ZN(n5811) );
  NAND2_X1 U7496 ( .A1(n5811), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5812) );
  NAND2_X1 U7497 ( .A1(n5893), .A2(n9283), .ZN(n5814) );
  NAND2_X1 U7498 ( .A1(n5868), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5813) );
  NAND2_X1 U7499 ( .A1(n9302), .A2(n9442), .ZN(n9274) );
  INV_X1 U7500 ( .A(n5815), .ZN(n9279) );
  INV_X1 U7501 ( .A(n6944), .ZN(n5816) );
  INV_X1 U7502 ( .A(n7014), .ZN(n9280) );
  AND2_X1 U7503 ( .A1(n9280), .A2(P1_B_REG_SCAN_IN), .ZN(n5817) );
  NOR2_X1 U7504 ( .A1(n9770), .A2(n5817), .ZN(n9522) );
  INV_X1 U7505 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9951) );
  NAND2_X1 U7506 ( .A1(n5786), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5819) );
  NAND2_X1 U7507 ( .A1(n4283), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5818) );
  OAI211_X1 U7508 ( .C1(n5820), .C2(n9951), .A(n5819), .B(n5818), .ZN(n9444)
         );
  AOI22_X1 U7509 ( .A1(n9446), .A2(n9794), .B1(n9522), .B2(n9444), .ZN(n5821)
         );
  NAND2_X1 U7510 ( .A1(n8059), .A2(n9446), .ZN(n9533) );
  INV_X1 U7511 ( .A(n9533), .ZN(n5822) );
  INV_X1 U7512 ( .A(n9753), .ZN(n10234) );
  NAND2_X1 U7513 ( .A1(n5822), .A2(n10234), .ZN(n5862) );
  INV_X1 U7514 ( .A(n9206), .ZN(n9322) );
  INV_X1 U7515 ( .A(n9769), .ZN(n9449) );
  OR2_X1 U7516 ( .A1(n9759), .A2(n9449), .ZN(n9727) );
  INV_X1 U7517 ( .A(n9727), .ZN(n5823) );
  OAI21_X1 U7518 ( .B1(n7298), .B2(n7087), .A(n5916), .ZN(n5825) );
  NAND2_X1 U7519 ( .A1(n7298), .A2(n7087), .ZN(n5824) );
  NAND2_X1 U7520 ( .A1(n5825), .A2(n5824), .ZN(n7426) );
  NAND2_X1 U7521 ( .A1(n7441), .A2(n7485), .ZN(n7438) );
  NAND2_X1 U7522 ( .A1(n4554), .A2(n10219), .ZN(n7383) );
  AND2_X1 U7523 ( .A1(n7438), .A2(n7383), .ZN(n5826) );
  NAND2_X1 U7524 ( .A1(n7424), .A2(n5826), .ZN(n5829) );
  INV_X1 U7525 ( .A(n7438), .ZN(n5827) );
  OAI21_X1 U7526 ( .B1(n4727), .B2(n5827), .A(n7437), .ZN(n5828) );
  NAND2_X1 U7527 ( .A1(n5831), .A2(n10224), .ZN(n7502) );
  NAND2_X1 U7528 ( .A1(n9167), .A2(n9171), .ZN(n9407) );
  NAND2_X1 U7529 ( .A1(n9457), .A2(n10198), .ZN(n7473) );
  AND2_X1 U7530 ( .A1(n9407), .A2(n7473), .ZN(n5832) );
  NAND2_X1 U7531 ( .A1(n7636), .A2(n10229), .ZN(n5833) );
  INV_X1 U7532 ( .A(n9410), .ZN(n7525) );
  INV_X1 U7533 ( .A(n7794), .ZN(n9455) );
  OR2_X1 U7534 ( .A1(n7698), .A2(n9455), .ZN(n5834) );
  INV_X1 U7535 ( .A(n7780), .ZN(n9454) );
  NAND2_X1 U7536 ( .A1(n10236), .A2(n9454), .ZN(n5835) );
  INV_X1 U7537 ( .A(n7858), .ZN(n9453) );
  AND2_X1 U7538 ( .A1(n10048), .A2(n9453), .ZN(n5837) );
  OR2_X1 U7539 ( .A1(n10048), .A2(n9453), .ZN(n5836) );
  INV_X1 U7540 ( .A(n9313), .ZN(n5838) );
  NAND2_X1 U7541 ( .A1(n5838), .A2(n9297), .ZN(n9179) );
  INV_X1 U7542 ( .A(n8009), .ZN(n9451) );
  NAND2_X1 U7543 ( .A1(n7920), .A2(n9451), .ZN(n5839) );
  NAND2_X1 U7544 ( .A1(n5840), .A2(n5839), .ZN(n8010) );
  NAND2_X1 U7545 ( .A1(n5505), .A2(n9189), .ZN(n9397) );
  NAND2_X1 U7546 ( .A1(n7951), .A2(n9795), .ZN(n5841) );
  INV_X1 U7547 ( .A(n9793), .ZN(n9785) );
  INV_X1 U7548 ( .A(n9771), .ZN(n9450) );
  NAND2_X1 U7549 ( .A1(n10029), .A2(n9797), .ZN(n5842) );
  NAND2_X1 U7550 ( .A1(n9734), .A2(n9750), .ZN(n5844) );
  OR2_X1 U7551 ( .A1(n10010), .A2(n9694), .ZN(n5845) );
  NAND2_X1 U7552 ( .A1(n10004), .A2(n9714), .ZN(n9672) );
  NAND2_X1 U7553 ( .A1(n10010), .A2(n9694), .ZN(n9670) );
  AND2_X1 U7554 ( .A1(n9672), .A2(n9670), .ZN(n5846) );
  NAND2_X1 U7555 ( .A1(n9214), .A2(n9215), .ZN(n9704) );
  INV_X1 U7556 ( .A(n9672), .ZN(n5847) );
  OR2_X1 U7557 ( .A1(n9704), .A2(n5847), .ZN(n5848) );
  AND2_X1 U7558 ( .A1(n5849), .A2(n5848), .ZN(n5850) );
  NAND2_X1 U7559 ( .A1(n9334), .A2(n9289), .ZN(n9663) );
  NAND2_X1 U7560 ( .A1(n9994), .A2(n9678), .ZN(n5851) );
  OR2_X1 U7561 ( .A1(n9991), .A2(n9658), .ZN(n5852) );
  NAND2_X1 U7562 ( .A1(n9991), .A2(n9658), .ZN(n5853) );
  OR2_X1 U7563 ( .A1(n9984), .A2(n9448), .ZN(n9422) );
  NOR2_X1 U7564 ( .A1(n9980), .A2(n9629), .ZN(n5855) );
  NAND2_X1 U7565 ( .A1(n9580), .A2(n9588), .ZN(n5857) );
  INV_X1 U7566 ( .A(n9567), .ZN(n9598) );
  OR2_X1 U7567 ( .A1(n9828), .A2(n9598), .ZN(n5856) );
  NAND2_X1 U7568 ( .A1(n9826), .A2(n9590), .ZN(n9393) );
  NOR2_X2 U7569 ( .A1(n7296), .A2(n9102), .ZN(n7418) );
  NOR2_X2 U7570 ( .A1(n7508), .A2(n10198), .ZN(n7511) );
  INV_X1 U7571 ( .A(n7698), .ZN(n7641) );
  NAND2_X1 U7572 ( .A1(n7477), .A2(n7641), .ZN(n7527) );
  INV_X1 U7573 ( .A(n10029), .ZN(n9778) );
  INV_X1 U7574 ( .A(n9759), .ZN(n10021) );
  INV_X1 U7575 ( .A(n10004), .ZN(n9700) );
  INV_X1 U7576 ( .A(n9999), .ZN(n9683) );
  NOR2_X2 U7577 ( .A1(n9650), .A2(n9984), .ZN(n9632) );
  INV_X1 U7578 ( .A(n9980), .ZN(n9615) );
  AND2_X2 U7579 ( .A1(n9632), .A2(n9615), .ZN(n9611) );
  AND2_X2 U7580 ( .A1(n9611), .A2(n9606), .ZN(n9581) );
  AOI21_X1 U7581 ( .B1(n9259), .B2(n8056), .A(n9528), .ZN(n9543) );
  NAND2_X1 U7582 ( .A1(n5893), .A2(n7088), .ZN(n5859) );
  INV_X1 U7583 ( .A(n7088), .ZN(n7084) );
  AOI22_X1 U7584 ( .A1(n9543), .A2(n10033), .B1(n9259), .B2(n10047), .ZN(n5860) );
  OAI211_X1 U7585 ( .C1(n9535), .C2(n5862), .A(n5861), .B(n5860), .ZN(n5863)
         );
  OAI21_X1 U7586 ( .B1(P1_IR_REG_22__SCAN_IN), .B2(P1_IR_REG_21__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5864) );
  INV_X1 U7587 ( .A(P1_B_REG_SCAN_IN), .ZN(n5867) );
  NAND2_X1 U7588 ( .A1(n4711), .A2(n5867), .ZN(n5879) );
  INV_X1 U7589 ( .A(n5868), .ZN(n5873) );
  NAND2_X1 U7590 ( .A1(n5870), .A2(n5869), .ZN(n5871) );
  NOR2_X1 U7591 ( .A1(n9954), .A2(n5871), .ZN(n5872) );
  NAND2_X1 U7592 ( .A1(n5873), .A2(n5872), .ZN(n5876) );
  NAND2_X1 U7593 ( .A1(n5876), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5875) );
  INV_X1 U7594 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5874) );
  XNOR2_X1 U7595 ( .A(n5875), .B(n5874), .ZN(n8024) );
  NAND3_X1 U7596 ( .A1(n8085), .A2(P1_B_REG_SCAN_IN), .A3(n8024), .ZN(n5878)
         );
  NAND3_X1 U7597 ( .A1(n5879), .A2(n5878), .A3(n5890), .ZN(n6983) );
  NOR2_X1 U7598 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .ZN(
        n9957) );
  NOR4_X1 U7599 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n5882) );
  NOR4_X1 U7600 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5881) );
  NOR4_X1 U7601 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5880) );
  AND4_X1 U7602 ( .A1(n9957), .A2(n5882), .A3(n5881), .A4(n5880), .ZN(n5888)
         );
  NOR4_X1 U7603 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n5886) );
  NOR4_X1 U7604 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n5885) );
  NOR4_X1 U7605 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_29__SCAN_IN), .ZN(n5884) );
  NOR4_X1 U7606 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n5883) );
  AND4_X1 U7607 ( .A1(n5886), .A2(n5885), .A3(n5884), .A4(n5883), .ZN(n5887)
         );
  AND2_X1 U7608 ( .A1(n5888), .A2(n5887), .ZN(n5889) );
  OR2_X1 U7609 ( .A1(n6983), .A2(n5889), .ZN(n6103) );
  AND2_X1 U7610 ( .A1(n7755), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5892) );
  OR2_X1 U7611 ( .A1(n5893), .A2(n9442), .ZN(n5901) );
  NAND2_X1 U7612 ( .A1(n5901), .A2(n6944), .ZN(n7291) );
  NAND3_X1 U7613 ( .A1(n6103), .A2(n9278), .A3(n7291), .ZN(n6767) );
  OR2_X1 U7614 ( .A1(n6983), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5895) );
  NAND2_X1 U7615 ( .A1(n8085), .A2(n5894), .ZN(n10074) );
  NAND2_X1 U7616 ( .A1(n5895), .A2(n10074), .ZN(n6766) );
  NOR2_X1 U7617 ( .A1(n6767), .A2(n6766), .ZN(n5898) );
  NAND2_X1 U7618 ( .A1(n5896), .A2(n9432), .ZN(n6111) );
  OR2_X1 U7619 ( .A1(n6983), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5897) );
  NAND2_X1 U7620 ( .A1(n5894), .A2(n8024), .ZN(n6984) );
  NAND2_X1 U7621 ( .A1(n5897), .A2(n6984), .ZN(n7415) );
  NAND2_X1 U7622 ( .A1(n6770), .A2(n10254), .ZN(n5900) );
  INV_X1 U7623 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5899) );
  NAND2_X1 U7624 ( .A1(n5900), .A2(n5212), .ZN(P1_U3552) );
  INV_X2 U7625 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  AND2_X4 U7626 ( .A1(n6943), .A2(n5903), .ZN(n6097) );
  AOI22_X1 U7627 ( .A1(n9819), .A2(n5985), .B1(n5929), .B2(n9447), .ZN(n8981)
         );
  AOI22_X1 U7628 ( .A1(n9819), .A2(n6097), .B1(n5985), .B2(n9447), .ZN(n5904)
         );
  XNOR2_X1 U7629 ( .A(n5904), .B(n7522), .ZN(n8980) );
  NAND2_X1 U7630 ( .A1(n9980), .A2(n6097), .ZN(n5906) );
  NAND2_X1 U7631 ( .A1(n9629), .A2(n5985), .ZN(n5905) );
  NAND2_X1 U7632 ( .A1(n5906), .A2(n5905), .ZN(n5907) );
  XNOR2_X1 U7633 ( .A(n5907), .B(n4720), .ZN(n8998) );
  NOR2_X1 U7634 ( .A1(n9093), .A2(n6093), .ZN(n5908) );
  AOI21_X1 U7635 ( .B1(n9980), .B2(n5985), .A(n5908), .ZN(n9029) );
  OR2_X1 U7636 ( .A1(n7082), .A2(n5935), .ZN(n5910) );
  INV_X1 U7637 ( .A(n6943), .ZN(n5911) );
  AOI22_X1 U7638 ( .A1(n5985), .A2(n7458), .B1(n5911), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n5909) );
  AOI22_X1 U7639 ( .A1(n6097), .A2(n7458), .B1(n5911), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n5912) );
  NAND2_X1 U7640 ( .A1(n5913), .A2(n5912), .ZN(n7138) );
  INV_X1 U7641 ( .A(n7138), .ZN(n5914) );
  NAND2_X1 U7642 ( .A1(n5914), .A2(n7522), .ZN(n5915) );
  NAND2_X1 U7643 ( .A1(n7137), .A2(n5915), .ZN(n7320) );
  OAI22_X1 U7644 ( .A1(n7087), .A2(n5969), .B1(n5916), .B2(n6073), .ZN(n5917)
         );
  XNOR2_X1 U7645 ( .A(n5917), .B(n6059), .ZN(n5921) );
  NAND2_X1 U7646 ( .A1(n7320), .A2(n5921), .ZN(n5920) );
  OR2_X1 U7647 ( .A1(n7087), .A2(n6083), .ZN(n5919) );
  NAND2_X1 U7648 ( .A1(n6056), .A2(n5858), .ZN(n5918) );
  NAND2_X1 U7649 ( .A1(n5919), .A2(n5918), .ZN(n7319) );
  NAND2_X1 U7650 ( .A1(n5920), .A2(n7319), .ZN(n5924) );
  INV_X1 U7651 ( .A(n7320), .ZN(n5922) );
  INV_X1 U7652 ( .A(n5921), .ZN(n7321) );
  NAND2_X1 U7653 ( .A1(n5922), .A2(n7321), .ZN(n5923) );
  NAND2_X1 U7654 ( .A1(n9460), .A2(n5985), .ZN(n5926) );
  NAND2_X1 U7655 ( .A1(n5926), .A2(n5925), .ZN(n5927) );
  NOR2_X1 U7656 ( .A1(n10219), .A2(n5902), .ZN(n5928) );
  NAND2_X1 U7657 ( .A1(n5931), .A2(n5930), .ZN(n5933) );
  AND2_X1 U7658 ( .A1(n5933), .A2(n5932), .ZN(n9100) );
  OAI22_X1 U7659 ( .A1(n7441), .A2(n5969), .B1(n7485), .B2(n6073), .ZN(n5934)
         );
  OR2_X1 U7660 ( .A1(n7441), .A2(n6083), .ZN(n5937) );
  NAND2_X1 U7661 ( .A1(n5985), .A2(n7387), .ZN(n5936) );
  NAND2_X1 U7662 ( .A1(n5937), .A2(n5936), .ZN(n5938) );
  INV_X1 U7663 ( .A(n5938), .ZN(n5939) );
  NAND2_X1 U7664 ( .A1(n9458), .A2(n6056), .ZN(n5942) );
  OR2_X1 U7665 ( .A1(n10224), .A2(n6073), .ZN(n5941) );
  NAND2_X1 U7666 ( .A1(n5942), .A2(n5941), .ZN(n5943) );
  XNOR2_X1 U7667 ( .A(n5943), .B(n7522), .ZN(n5946) );
  NAND2_X1 U7668 ( .A1(n5929), .A2(n9458), .ZN(n5945) );
  INV_X1 U7669 ( .A(n5985), .ZN(n5969) );
  OR2_X1 U7670 ( .A1(n10224), .A2(n5902), .ZN(n5944) );
  NAND2_X1 U7671 ( .A1(n5945), .A2(n5944), .ZN(n5947) );
  NAND2_X1 U7672 ( .A1(n5946), .A2(n5947), .ZN(n9066) );
  INV_X1 U7673 ( .A(n5946), .ZN(n5949) );
  INV_X1 U7674 ( .A(n5947), .ZN(n5948) );
  NAND2_X1 U7675 ( .A1(n5949), .A2(n5948), .ZN(n9065) );
  OAI22_X1 U7676 ( .A1(n7471), .A2(n5902), .B1(n7409), .B2(n6073), .ZN(n5951)
         );
  XNOR2_X1 U7677 ( .A(n5951), .B(n4720), .ZN(n7406) );
  OR2_X1 U7678 ( .A1(n7471), .A2(n6093), .ZN(n5953) );
  NAND2_X1 U7679 ( .A1(n10198), .A2(n6056), .ZN(n5952) );
  AND2_X1 U7680 ( .A1(n5953), .A2(n5952), .ZN(n7405) );
  AND2_X1 U7681 ( .A1(n7406), .A2(n7405), .ZN(n5957) );
  INV_X1 U7682 ( .A(n7406), .ZN(n5955) );
  INV_X1 U7683 ( .A(n7405), .ZN(n5954) );
  NAND2_X1 U7684 ( .A1(n5955), .A2(n5954), .ZN(n5956) );
  NAND2_X1 U7685 ( .A1(n9123), .A2(n6056), .ZN(n5958) );
  NAND2_X1 U7686 ( .A1(n7698), .A2(n6097), .ZN(n5960) );
  OR2_X1 U7687 ( .A1(n7794), .A2(n5902), .ZN(n5959) );
  NAND2_X1 U7688 ( .A1(n5960), .A2(n5959), .ZN(n5961) );
  XNOR2_X1 U7689 ( .A(n5961), .B(n7522), .ZN(n7630) );
  NAND2_X1 U7690 ( .A1(n7698), .A2(n6056), .ZN(n5963) );
  OR2_X1 U7691 ( .A1(n7794), .A2(n6083), .ZN(n5962) );
  NAND2_X1 U7692 ( .A1(n5963), .A2(n5962), .ZN(n7629) );
  NAND2_X1 U7693 ( .A1(n7630), .A2(n7629), .ZN(n7628) );
  OAI21_X1 U7694 ( .B1(n9118), .B2(n9119), .A(n7628), .ZN(n5964) );
  INV_X1 U7695 ( .A(n7630), .ZN(n5966) );
  NOR2_X1 U7696 ( .A1(n7629), .A2(n4709), .ZN(n5965) );
  NAND2_X1 U7697 ( .A1(n10048), .A2(n6097), .ZN(n5971) );
  OR2_X1 U7698 ( .A1(n7858), .A2(n5902), .ZN(n5970) );
  NAND2_X1 U7699 ( .A1(n5971), .A2(n5970), .ZN(n5972) );
  XNOR2_X1 U7700 ( .A(n5972), .B(n7522), .ZN(n7776) );
  NAND2_X1 U7701 ( .A1(n10048), .A2(n6056), .ZN(n5974) );
  OR2_X1 U7702 ( .A1(n7858), .A2(n6093), .ZN(n5973) );
  NAND2_X1 U7703 ( .A1(n5974), .A2(n5973), .ZN(n7775) );
  NAND2_X1 U7704 ( .A1(n10236), .A2(n6097), .ZN(n5976) );
  OR2_X1 U7705 ( .A1(n7780), .A2(n5902), .ZN(n5975) );
  NAND2_X1 U7706 ( .A1(n5976), .A2(n5975), .ZN(n5977) );
  XNOR2_X1 U7707 ( .A(n5977), .B(n7522), .ZN(n7774) );
  NAND2_X1 U7708 ( .A1(n10236), .A2(n6056), .ZN(n5979) );
  OR2_X1 U7709 ( .A1(n7780), .A2(n6083), .ZN(n5978) );
  NAND2_X1 U7710 ( .A1(n5979), .A2(n5978), .ZN(n7771) );
  AOI22_X1 U7711 ( .A1(n7776), .A2(n7775), .B1(n7774), .B2(n7771), .ZN(n5980)
         );
  OAI21_X1 U7712 ( .B1(n7774), .B2(n7771), .A(n7775), .ZN(n5983) );
  INV_X1 U7713 ( .A(n7776), .ZN(n5982) );
  INV_X1 U7714 ( .A(n7774), .ZN(n7789) );
  NOR2_X1 U7715 ( .A1(n7775), .A2(n7771), .ZN(n5981) );
  OAI22_X1 U7716 ( .A1(n7767), .A2(n6073), .B1(n7878), .B2(n5902), .ZN(n5984)
         );
  XNOR2_X1 U7717 ( .A(n5984), .B(n4720), .ZN(n5990) );
  OR2_X1 U7718 ( .A1(n7767), .A2(n5902), .ZN(n5987) );
  NAND2_X1 U7719 ( .A1(n5929), .A2(n9452), .ZN(n5986) );
  NAND2_X1 U7720 ( .A1(n5987), .A2(n5986), .ZN(n5988) );
  XNOR2_X1 U7721 ( .A(n5990), .B(n5988), .ZN(n7706) );
  INV_X1 U7722 ( .A(n5988), .ZN(n5989) );
  NAND2_X1 U7723 ( .A1(n5990), .A2(n5989), .ZN(n5991) );
  NAND2_X1 U7724 ( .A1(n7920), .A2(n6097), .ZN(n5994) );
  OR2_X1 U7725 ( .A1(n8009), .A2(n5902), .ZN(n5993) );
  NAND2_X1 U7726 ( .A1(n5994), .A2(n5993), .ZN(n5995) );
  XNOR2_X1 U7727 ( .A(n5995), .B(n4720), .ZN(n5999) );
  NOR2_X1 U7728 ( .A1(n8009), .A2(n6093), .ZN(n5996) );
  AOI21_X1 U7729 ( .B1(n7920), .B2(n6056), .A(n5996), .ZN(n5998) );
  XNOR2_X1 U7730 ( .A(n5999), .B(n5998), .ZN(n7873) );
  OR2_X1 U7731 ( .A1(n5999), .A2(n5998), .ZN(n6000) );
  OAI22_X1 U7732 ( .A1(n10040), .A2(n6073), .B1(n6001), .B2(n5902), .ZN(n6002)
         );
  XNOR2_X1 U7733 ( .A(n6002), .B(n7522), .ZN(n7945) );
  INV_X1 U7734 ( .A(n7945), .ZN(n6005) );
  OR2_X1 U7735 ( .A1(n10040), .A2(n5902), .ZN(n6004) );
  NAND2_X1 U7736 ( .A1(n5929), .A2(n9795), .ZN(n6003) );
  NAND2_X1 U7737 ( .A1(n6004), .A2(n6003), .ZN(n6006) );
  INV_X1 U7738 ( .A(n6006), .ZN(n7944) );
  NAND2_X1 U7739 ( .A1(n6005), .A2(n7944), .ZN(n6008) );
  AND2_X1 U7740 ( .A1(n7945), .A2(n6006), .ZN(n6007) );
  NAND2_X1 U7741 ( .A1(n10032), .A2(n6097), .ZN(n6010) );
  OR2_X1 U7742 ( .A1(n9771), .A2(n5902), .ZN(n6009) );
  NAND2_X1 U7743 ( .A1(n6010), .A2(n6009), .ZN(n6011) );
  XNOR2_X1 U7744 ( .A(n6011), .B(n7522), .ZN(n6014) );
  NAND2_X1 U7745 ( .A1(n10032), .A2(n5985), .ZN(n6013) );
  OR2_X1 U7746 ( .A1(n9771), .A2(n6083), .ZN(n6012) );
  NAND2_X1 U7747 ( .A1(n6013), .A2(n6012), .ZN(n6015) );
  NAND2_X1 U7748 ( .A1(n6014), .A2(n6015), .ZN(n8040) );
  INV_X1 U7749 ( .A(n6014), .ZN(n6017) );
  INV_X1 U7750 ( .A(n6015), .ZN(n6016) );
  NAND2_X1 U7751 ( .A1(n6017), .A2(n6016), .ZN(n8042) );
  NAND2_X1 U7752 ( .A1(n10029), .A2(n6097), .ZN(n6019) );
  NAND2_X1 U7753 ( .A1(n9797), .A2(n5985), .ZN(n6018) );
  NAND2_X1 U7754 ( .A1(n6019), .A2(n6018), .ZN(n6020) );
  XNOR2_X1 U7755 ( .A(n6020), .B(n4720), .ZN(n6023) );
  NAND2_X1 U7756 ( .A1(n10029), .A2(n5985), .ZN(n6022) );
  NAND2_X1 U7757 ( .A1(n9797), .A2(n5929), .ZN(n6021) );
  NAND2_X1 U7758 ( .A1(n6022), .A2(n6021), .ZN(n8989) );
  NAND2_X1 U7759 ( .A1(n9759), .A2(n6097), .ZN(n6026) );
  NAND2_X1 U7760 ( .A1(n9449), .A2(n6056), .ZN(n6025) );
  NAND2_X1 U7761 ( .A1(n6026), .A2(n6025), .ZN(n6027) );
  XNOR2_X1 U7762 ( .A(n6027), .B(n7522), .ZN(n6029) );
  NOR2_X1 U7763 ( .A1(n9769), .A2(n6093), .ZN(n6028) );
  AOI21_X1 U7764 ( .B1(n9759), .B2(n5985), .A(n6028), .ZN(n9142) );
  AOI22_X1 U7765 ( .A1(n10010), .A2(n6097), .B1(n6056), .B2(n9694), .ZN(n6030)
         );
  XNOR2_X1 U7766 ( .A(n6030), .B(n7522), .ZN(n6035) );
  NOR2_X1 U7767 ( .A1(n9722), .A2(n6083), .ZN(n6031) );
  AOI21_X1 U7768 ( .B1(n10010), .B2(n6056), .A(n6031), .ZN(n9049) );
  OAI22_X1 U7769 ( .A1(n10016), .A2(n6073), .B1(n9147), .B2(n5902), .ZN(n6032)
         );
  XNOR2_X1 U7770 ( .A(n6032), .B(n7522), .ZN(n9045) );
  OAI22_X1 U7771 ( .A1(n10016), .A2(n5902), .B1(n9147), .B2(n6093), .ZN(n9044)
         );
  NAND2_X1 U7772 ( .A1(n9045), .A2(n9044), .ZN(n6033) );
  OAI21_X1 U7773 ( .B1(n6035), .B2(n9049), .A(n6033), .ZN(n6034) );
  INV_X1 U7774 ( .A(n6034), .ZN(n6040) );
  INV_X1 U7775 ( .A(n6035), .ZN(n9050) );
  INV_X1 U7776 ( .A(n9045), .ZN(n9048) );
  INV_X1 U7777 ( .A(n9044), .ZN(n6037) );
  AOI21_X1 U7778 ( .B1(n9048), .B2(n6037), .A(n9049), .ZN(n6036) );
  NAND3_X1 U7779 ( .A1(n9048), .A2(n6037), .A3(n9049), .ZN(n6038) );
  NAND2_X1 U7780 ( .A1(n9999), .A2(n6097), .ZN(n6042) );
  NAND2_X1 U7781 ( .A1(n9695), .A2(n5985), .ZN(n6041) );
  NAND2_X1 U7782 ( .A1(n6042), .A2(n6041), .ZN(n6043) );
  XNOR2_X1 U7783 ( .A(n6043), .B(n4720), .ZN(n6051) );
  NOR2_X1 U7784 ( .A1(n9112), .A2(n6083), .ZN(n6044) );
  AOI21_X1 U7785 ( .B1(n9999), .B2(n5985), .A(n6044), .ZN(n6050) );
  NAND2_X1 U7786 ( .A1(n10004), .A2(n6097), .ZN(n6046) );
  NAND2_X1 U7787 ( .A1(n9714), .A2(n5985), .ZN(n6045) );
  NAND2_X1 U7788 ( .A1(n6046), .A2(n6045), .ZN(n6047) );
  XNOR2_X1 U7789 ( .A(n6047), .B(n4720), .ZN(n9006) );
  NOR2_X1 U7790 ( .A1(n9054), .A2(n6083), .ZN(n6048) );
  AOI21_X1 U7791 ( .B1(n10004), .B2(n5985), .A(n6048), .ZN(n9110) );
  INV_X1 U7792 ( .A(n9009), .ZN(n6053) );
  NAND2_X1 U7793 ( .A1(n9006), .A2(n9110), .ZN(n6052) );
  NAND2_X1 U7794 ( .A1(n6051), .A2(n6050), .ZN(n9008) );
  NAND2_X1 U7795 ( .A1(n9994), .A2(n6097), .ZN(n6058) );
  NAND2_X1 U7796 ( .A1(n9678), .A2(n5985), .ZN(n6057) );
  NAND2_X1 U7797 ( .A1(n6058), .A2(n6057), .ZN(n6060) );
  XNOR2_X1 U7798 ( .A(n6060), .B(n4720), .ZN(n6063) );
  NOR2_X1 U7799 ( .A1(n9647), .A2(n6093), .ZN(n6061) );
  AOI21_X1 U7800 ( .B1(n9994), .B2(n5985), .A(n6061), .ZN(n6062) );
  AND2_X1 U7801 ( .A1(n6063), .A2(n6062), .ZN(n9077) );
  OR2_X1 U7802 ( .A1(n6063), .A2(n6062), .ZN(n9078) );
  NAND2_X1 U7803 ( .A1(n9991), .A2(n6097), .ZN(n6065) );
  OR2_X1 U7804 ( .A1(n9220), .A2(n5902), .ZN(n6064) );
  NAND2_X1 U7805 ( .A1(n6065), .A2(n6064), .ZN(n6066) );
  XNOR2_X1 U7806 ( .A(n6066), .B(n4720), .ZN(n6069) );
  NOR2_X1 U7807 ( .A1(n9220), .A2(n6083), .ZN(n6067) );
  AOI21_X1 U7808 ( .B1(n9991), .B2(n5985), .A(n6067), .ZN(n6068) );
  NOR2_X1 U7809 ( .A1(n6069), .A2(n6068), .ZN(n9019) );
  NAND2_X1 U7810 ( .A1(n6069), .A2(n6068), .ZN(n9017) );
  INV_X1 U7811 ( .A(n9090), .ZN(n6072) );
  AOI22_X1 U7812 ( .A1(n9984), .A2(n5985), .B1(n5929), .B2(n9448), .ZN(n9087)
         );
  INV_X1 U7813 ( .A(n9087), .ZN(n6071) );
  AOI22_X1 U7814 ( .A1(n9984), .A2(n6097), .B1(n5985), .B2(n9448), .ZN(n6070)
         );
  XNOR2_X1 U7815 ( .A(n6070), .B(n7522), .ZN(n9088) );
  OAI22_X1 U7816 ( .A1(n9606), .A2(n6073), .B1(n9617), .B2(n5902), .ZN(n6074)
         );
  XNOR2_X1 U7817 ( .A(n6074), .B(n7522), .ZN(n6075) );
  OAI22_X1 U7818 ( .A1(n9606), .A2(n5902), .B1(n9617), .B2(n6093), .ZN(n6076)
         );
  NAND2_X1 U7819 ( .A1(n6075), .A2(n6076), .ZN(n9030) );
  NAND3_X1 U7820 ( .A1(n9030), .A2(n8998), .A3(n9029), .ZN(n6079) );
  INV_X1 U7821 ( .A(n6075), .ZN(n6078) );
  INV_X1 U7822 ( .A(n6076), .ZN(n6077) );
  NAND2_X1 U7823 ( .A1(n6078), .A2(n6077), .ZN(n9031) );
  NAND2_X1 U7824 ( .A1(n9828), .A2(n6097), .ZN(n6081) );
  OR2_X1 U7825 ( .A1(n9567), .A2(n5902), .ZN(n6080) );
  NAND2_X1 U7826 ( .A1(n6081), .A2(n6080), .ZN(n6082) );
  XNOR2_X1 U7827 ( .A(n6082), .B(n7522), .ZN(n6088) );
  NOR2_X1 U7828 ( .A1(n9567), .A2(n6093), .ZN(n6084) );
  AOI21_X1 U7829 ( .B1(n9828), .B2(n5985), .A(n6084), .ZN(n6086) );
  XNOR2_X1 U7830 ( .A(n6088), .B(n6086), .ZN(n9032) );
  INV_X1 U7831 ( .A(n6086), .ZN(n6087) );
  NAND2_X1 U7832 ( .A1(n9826), .A2(n6097), .ZN(n6091) );
  NAND2_X1 U7833 ( .A1(n9590), .A2(n5985), .ZN(n6090) );
  NAND2_X1 U7834 ( .A1(n6091), .A2(n6090), .ZN(n6092) );
  XNOR2_X1 U7835 ( .A(n6092), .B(n4720), .ZN(n6096) );
  NOR2_X1 U7836 ( .A1(n9549), .A2(n6093), .ZN(n6094) );
  AOI21_X1 U7837 ( .B1(n9826), .B2(n5985), .A(n6094), .ZN(n6095) );
  OR2_X1 U7838 ( .A1(n6096), .A2(n6095), .ZN(n9131) );
  NAND2_X1 U7839 ( .A1(n8059), .A2(n6097), .ZN(n6099) );
  NAND2_X1 U7840 ( .A1(n9446), .A2(n5985), .ZN(n6098) );
  NAND2_X1 U7841 ( .A1(n6099), .A2(n6098), .ZN(n6100) );
  XNOR2_X1 U7842 ( .A(n6100), .B(n7522), .ZN(n6102) );
  AOI22_X1 U7843 ( .A1(n8059), .A2(n5985), .B1(n5929), .B2(n9446), .ZN(n6101)
         );
  XNOR2_X1 U7844 ( .A(n6102), .B(n6101), .ZN(n6127) );
  INV_X1 U7845 ( .A(n6127), .ZN(n6106) );
  INV_X1 U7846 ( .A(n6103), .ZN(n6104) );
  NOR2_X1 U7847 ( .A1(n10047), .A2(n6944), .ZN(n6105) );
  NAND2_X1 U7848 ( .A1(n6107), .A2(n5220), .ZN(n6132) );
  OR2_X1 U7849 ( .A1(n8980), .A2(n8981), .ZN(n6126) );
  NAND4_X1 U7850 ( .A1(n6108), .A2(n6127), .A3(n6126), .A4(n9145), .ZN(n6131)
         );
  NAND2_X1 U7851 ( .A1(n7292), .A2(n10199), .ZN(n6112) );
  INV_X1 U7852 ( .A(n6113), .ZN(n6115) );
  NAND2_X1 U7853 ( .A1(n6115), .A2(n6114), .ZN(n7523) );
  INV_X1 U7854 ( .A(n7523), .ZN(n9281) );
  INV_X1 U7855 ( .A(n6117), .ZN(n6116) );
  NAND2_X1 U7856 ( .A1(n9447), .A2(n9150), .ZN(n6125) );
  INV_X1 U7857 ( .A(n8055), .ZN(n6123) );
  NAND2_X1 U7858 ( .A1(n6120), .A2(n10237), .ZN(n6118) );
  NAND4_X1 U7859 ( .A1(n6118), .A2(n7755), .A3(n7291), .A4(n6943), .ZN(n6119)
         );
  NAND2_X1 U7860 ( .A1(n6119), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6122) );
  NAND3_X1 U7861 ( .A1(n6120), .A2(n10199), .A3(n9278), .ZN(n6121) );
  AOI22_X1 U7862 ( .A1(n6123), .A2(n9134), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n6124) );
  OAI211_X1 U7863 ( .C1(n9263), .C2(n9148), .A(n6125), .B(n6124), .ZN(n6129)
         );
  NOR3_X1 U7864 ( .A1(n6127), .A2(n9140), .A3(n6126), .ZN(n6128) );
  AOI211_X1 U7865 ( .C1(n8059), .C2(n9138), .A(n6129), .B(n6128), .ZN(n6130)
         );
  NAND3_X1 U7866 ( .A1(n6132), .A2(n6131), .A3(n6130), .ZN(P1_U3218) );
  NOR2_X2 U7867 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6194) );
  NAND2_X1 U7868 ( .A1(n6194), .A2(n4993), .ZN(n6195) );
  INV_X1 U7869 ( .A(n6195), .ZN(n6134) );
  NAND2_X1 U7870 ( .A1(n6134), .A2(n6133), .ZN(n6176) );
  NAND2_X1 U7871 ( .A1(n6212), .A2(n6208), .ZN(n6177) );
  INV_X1 U7872 ( .A(n6177), .ZN(n6138) );
  NOR2_X1 U7873 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n6137) );
  NOR2_X1 U7874 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n6136) );
  NOR2_X1 U7875 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n6135) );
  NAND4_X1 U7876 ( .A1(n6138), .A2(n6137), .A3(n6136), .A4(n6135), .ZN(n6143)
         );
  NOR2_X1 U7877 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n6141) );
  NAND4_X1 U7878 ( .A1(n6141), .A2(n6140), .A3(n6179), .A4(n6139), .ZN(n6142)
         );
  NAND2_X1 U7879 ( .A1(n6240), .A2(n6239), .ZN(n6147) );
  INV_X1 U7880 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6149) );
  NOR2_X1 U7881 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n6154) );
  NOR2_X1 U7882 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n6153) );
  NOR2_X1 U7883 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n6152) );
  NAND4_X1 U7884 ( .A1(n6155), .A2(n6154), .A3(n6153), .A4(n6152), .ZN(n6162)
         );
  OR2_X1 U7885 ( .A1(n6151), .A2(n6162), .ZN(n6157) );
  NAND2_X1 U7886 ( .A1(n6157), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6156) );
  XNOR2_X1 U7887 ( .A(n6156), .B(n6160), .ZN(n8023) );
  OAI21_X1 U7888 ( .B1(n6157), .B2(P2_IR_REG_25__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6158) );
  MUX2_X1 U7889 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6158), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6164) );
  NAND2_X1 U7890 ( .A1(n6160), .A2(n6159), .ZN(n6161) );
  NAND2_X1 U7891 ( .A1(n6164), .A2(n6290), .ZN(n8978) );
  OR2_X1 U7892 ( .A1(n6166), .A2(n6165), .ZN(n6167) );
  NAND2_X1 U7893 ( .A1(n6168), .A2(n6167), .ZN(n6933) );
  INV_X1 U7894 ( .A(n10312), .ZN(n6169) );
  NOR2_X2 U7895 ( .A1(n6934), .A2(n6169), .ZN(P2_U3966) );
  INV_X1 U7896 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n6170) );
  INV_X1 U7897 ( .A(n6268), .ZN(n6172) );
  NAND2_X1 U7898 ( .A1(n6172), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6173) );
  XNOR2_X1 U7899 ( .A(n6173), .B(P2_IR_REG_18__SCAN_IN), .ZN(n7351) );
  OR2_X1 U7900 ( .A1(n7351), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U7901 ( .A1(n7351), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6174) );
  AND2_X1 U7902 ( .A1(n6236), .A2(n6174), .ZN(n8488) );
  INV_X1 U7903 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n6479) );
  NAND2_X1 U7904 ( .A1(n6151), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6175) );
  XNOR2_X1 U7905 ( .A(n6175), .B(P2_IR_REG_17__SCAN_IN), .ZN(n6473) );
  INV_X1 U7906 ( .A(n6473), .ZN(n8483) );
  XNOR2_X1 U7907 ( .A(n8483), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8479) );
  NOR2_X1 U7908 ( .A1(n6176), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n6206) );
  NOR2_X1 U7909 ( .A1(n6177), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n6178) );
  NAND2_X1 U7910 ( .A1(n6206), .A2(n6178), .ZN(n6192) );
  INV_X1 U7911 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6223) );
  INV_X1 U7912 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6219) );
  NAND3_X1 U7913 ( .A1(n6223), .A2(n6219), .A3(n6179), .ZN(n6180) );
  NOR2_X1 U7914 ( .A1(n6218), .A2(n6180), .ZN(n6227) );
  INV_X1 U7915 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6181) );
  NAND2_X1 U7916 ( .A1(n6227), .A2(n6181), .ZN(n6185) );
  INV_X1 U7917 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6182) );
  INV_X1 U7918 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6188) );
  INV_X1 U7919 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6186) );
  NAND3_X1 U7920 ( .A1(n6182), .A2(n6188), .A3(n6186), .ZN(n6183) );
  OAI21_X1 U7921 ( .B1(n6185), .B2(n6183), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6184) );
  XNOR2_X1 U7922 ( .A(n6184), .B(P2_IR_REG_16__SCAN_IN), .ZN(n6454) );
  INV_X1 U7923 ( .A(n6454), .ZN(n8469) );
  INV_X1 U7924 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n6234) );
  XNOR2_X1 U7925 ( .A(n6454), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8463) );
  NAND2_X1 U7926 ( .A1(n6185), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6229) );
  NAND2_X1 U7927 ( .A1(n6229), .A2(n6186), .ZN(n6187) );
  NAND2_X1 U7928 ( .A1(n6187), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6191) );
  NAND2_X1 U7929 ( .A1(n6191), .A2(n6188), .ZN(n6189) );
  NAND2_X1 U7930 ( .A1(n6189), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6190) );
  XNOR2_X1 U7931 ( .A(n6190), .B(P2_IR_REG_15__SCAN_IN), .ZN(n6443) );
  XNOR2_X1 U7932 ( .A(n6191), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7062) );
  INV_X1 U7933 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10350) );
  NAND2_X1 U7934 ( .A1(n6192), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6193) );
  XNOR2_X1 U7935 ( .A(n6193), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7279) );
  INV_X1 U7936 ( .A(n7279), .ZN(n7287) );
  INV_X1 U7937 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6196) );
  MUX2_X1 U7938 ( .A(n6196), .B(P2_REG1_REG_2__SCAN_IN), .S(n7172), .Z(n6200)
         );
  INV_X1 U7939 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6297) );
  MUX2_X1 U7940 ( .A(n6297), .B(P2_REG1_REG_1__SCAN_IN), .S(n7161), .Z(n6198)
         );
  AND2_X1 U7941 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(
        n6197) );
  NAND2_X1 U7942 ( .A1(n6198), .A2(n6197), .ZN(n7158) );
  INV_X1 U7943 ( .A(n7161), .ZN(n6250) );
  NAND2_X1 U7944 ( .A1(n6250), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6199) );
  NAND2_X1 U7945 ( .A1(n7158), .A2(n6199), .ZN(n7168) );
  NAND2_X1 U7946 ( .A1(n6200), .A2(n7168), .ZN(n7205) );
  INV_X1 U7947 ( .A(n7172), .ZN(n6251) );
  NAND2_X1 U7948 ( .A1(n6251), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7204) );
  INV_X1 U7949 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7651) );
  NAND2_X1 U7950 ( .A1(n6201), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6202) );
  MUX2_X1 U7951 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n7651), .S(n7211), .Z(n7203)
         );
  AOI21_X1 U7952 ( .B1(n7205), .B2(n7204), .A(n7203), .ZN(n7218) );
  NOR2_X1 U7953 ( .A1(n7211), .A2(n7651), .ZN(n7217) );
  INV_X1 U7954 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6205) );
  NAND2_X1 U7955 ( .A1(n6176), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6204) );
  INV_X1 U7956 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6203) );
  XNOR2_X1 U7957 ( .A(n6204), .B(n6203), .ZN(n7225) );
  MUX2_X1 U7958 ( .A(n6205), .B(P2_REG1_REG_4__SCAN_IN), .S(n7225), .Z(n7216)
         );
  OAI21_X1 U7959 ( .B1(n7218), .B2(n7217), .A(n7216), .ZN(n7256) );
  INV_X1 U7960 ( .A(n7225), .ZN(n6253) );
  NAND2_X1 U7961 ( .A1(n6253), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7255) );
  INV_X1 U7962 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6207) );
  OR2_X1 U7963 ( .A1(n6206), .A2(n6293), .ZN(n6209) );
  XNOR2_X1 U7964 ( .A(n6209), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6350) );
  MUX2_X1 U7965 ( .A(n6207), .B(P2_REG1_REG_5__SCAN_IN), .S(n6350), .Z(n7254)
         );
  AOI21_X1 U7966 ( .B1(n7256), .B2(n7255), .A(n7254), .ZN(n7258) );
  INV_X1 U7967 ( .A(n6350), .ZN(n7262) );
  NOR2_X1 U7968 ( .A1(n7262), .A2(n6207), .ZN(n7230) );
  INV_X1 U7969 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6211) );
  NAND2_X1 U7970 ( .A1(n6209), .A2(n6208), .ZN(n6210) );
  NAND2_X1 U7971 ( .A1(n6210), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6213) );
  XNOR2_X1 U7972 ( .A(n6213), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6966) );
  MUX2_X1 U7973 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6211), .S(n6966), .Z(n7229)
         );
  OAI21_X1 U7974 ( .B1(n7258), .B2(n7230), .A(n7229), .ZN(n7243) );
  NAND2_X1 U7975 ( .A1(n6966), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7242) );
  INV_X1 U7976 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6216) );
  NAND2_X1 U7977 ( .A1(n6213), .A2(n6212), .ZN(n6214) );
  NAND2_X1 U7978 ( .A1(n6214), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6215) );
  XNOR2_X1 U7979 ( .A(n6215), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6365) );
  MUX2_X1 U7980 ( .A(n6216), .B(P2_REG1_REG_7__SCAN_IN), .S(n6365), .Z(n7241)
         );
  AOI21_X1 U7981 ( .B1(n7243), .B2(n7242), .A(n7241), .ZN(n7284) );
  INV_X1 U7982 ( .A(n6365), .ZN(n7249) );
  NOR2_X1 U7983 ( .A1(n7249), .A2(n6216), .ZN(n7278) );
  MUX2_X1 U7984 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n10350), .S(n7279), .Z(n6217)
         );
  OAI21_X1 U7985 ( .B1(n7284), .B2(n7278), .A(n6217), .ZN(n7282) );
  OAI21_X1 U7986 ( .B1(n10350), .B2(n7287), .A(n7282), .ZN(n7491) );
  NAND2_X1 U7987 ( .A1(n6218), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6220) );
  XNOR2_X1 U7988 ( .A(n6220), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6976) );
  XOR2_X1 U7989 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n6976), .Z(n7492) );
  AOI22_X1 U7990 ( .A1(n7491), .A2(n7492), .B1(P2_REG1_REG_9__SCAN_IN), .B2(
        n6976), .ZN(n7670) );
  NAND2_X1 U7991 ( .A1(n6220), .A2(n6219), .ZN(n6221) );
  NAND2_X1 U7992 ( .A1(n6221), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6224) );
  XNOR2_X1 U7993 ( .A(n6224), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6395) );
  XNOR2_X1 U7994 ( .A(n6395), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n7671) );
  INV_X1 U7995 ( .A(n6395), .ZN(n7674) );
  INV_X1 U7996 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6222) );
  OAI22_X1 U7997 ( .A1(n7670), .A2(n7671), .B1(n7674), .B2(n6222), .ZN(n7808)
         );
  NAND2_X1 U7998 ( .A1(n6224), .A2(n6223), .ZN(n6225) );
  NAND2_X1 U7999 ( .A1(n6225), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6226) );
  XNOR2_X1 U8000 ( .A(n6226), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6990) );
  INV_X1 U8001 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n8883) );
  XNOR2_X1 U8002 ( .A(n6990), .B(n8883), .ZN(n7807) );
  AOI22_X1 U8003 ( .A1(n7808), .A2(n7807), .B1(P2_REG1_REG_11__SCAN_IN), .B2(
        n6990), .ZN(n8027) );
  OR2_X1 U8004 ( .A1(n6227), .A2(n6293), .ZN(n6228) );
  XNOR2_X1 U8005 ( .A(n6228), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6994) );
  NOR2_X1 U8006 ( .A1(n6994), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8428) );
  AOI21_X1 U8007 ( .B1(n6994), .B2(P2_REG1_REG_12__SCAN_IN), .A(n8428), .ZN(
        n8028) );
  XNOR2_X1 U8008 ( .A(n6229), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7011) );
  OR2_X1 U8009 ( .A1(n7011), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6231) );
  NAND2_X1 U8010 ( .A1(n7011), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6230) );
  AND2_X1 U8011 ( .A1(n6231), .A2(n6230), .ZN(n8427) );
  OAI21_X1 U8012 ( .B1(n8429), .B2(n8428), .A(n8427), .ZN(n8431) );
  NAND2_X1 U8013 ( .A1(n8431), .A2(n6231), .ZN(n8444) );
  INV_X1 U8014 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8864) );
  XNOR2_X1 U8015 ( .A(n7062), .B(n8864), .ZN(n8445) );
  NAND2_X1 U8016 ( .A1(n8444), .A2(n8445), .ZN(n8443) );
  OAI21_X1 U8017 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n7062), .A(n8443), .ZN(
        n6232) );
  XOR2_X1 U8018 ( .A(n6443), .B(n6232), .Z(n8453) );
  INV_X1 U8019 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n6233) );
  INV_X1 U8020 ( .A(n6443), .ZN(n8456) );
  OAI22_X1 U8021 ( .A1(n8453), .A2(n6233), .B1(n8456), .B2(n6232), .ZN(n8464)
         );
  NOR2_X1 U8022 ( .A1(n8463), .A2(n8464), .ZN(n8462) );
  AOI21_X1 U8023 ( .B1(n8469), .B2(n6234), .A(n8462), .ZN(n8480) );
  NAND2_X1 U8024 ( .A1(n8479), .A2(n8480), .ZN(n8478) );
  OAI21_X1 U8025 ( .B1(n6479), .B2(n8483), .A(n8478), .ZN(n6235) );
  INV_X1 U8026 ( .A(n6235), .ZN(n8487) );
  NAND2_X1 U8027 ( .A1(n8488), .A2(n8487), .ZN(n8486) );
  NAND2_X1 U8028 ( .A1(n8486), .A2(n6236), .ZN(n6237) );
  XNOR2_X1 U8029 ( .A(n6237), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n6270) );
  NAND2_X1 U8030 ( .A1(n6615), .A2(n6639), .ZN(n7341) );
  INV_X1 U8031 ( .A(n7341), .ZN(n6275) );
  INV_X1 U8032 ( .A(n6933), .ZN(n6241) );
  INV_X1 U8033 ( .A(n6764), .ZN(n7759) );
  INV_X1 U8034 ( .A(n6934), .ZN(n6242) );
  NAND2_X1 U8035 ( .A1(n6242), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6243) );
  OAI211_X1 U8036 ( .C1(n10303), .C2(n6275), .A(n7759), .B(n6243), .ZN(n6262)
         );
  XNOR2_X2 U8037 ( .A(n6247), .B(n6246), .ZN(n8971) );
  AND2_X1 U8038 ( .A1(n6319), .A2(n8971), .ZN(n6248) );
  NAND2_X1 U8039 ( .A1(n6262), .A2(n6248), .ZN(n10261) );
  NAND2_X1 U8040 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n6454), .ZN(n6249) );
  OAI21_X1 U8041 ( .B1(n6454), .B2(P2_REG2_REG_16__SCAN_IN), .A(n6249), .ZN(
        n8466) );
  INV_X1 U8042 ( .A(n7211), .ZN(n6252) );
  INV_X1 U8043 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9858) );
  NAND2_X1 U8044 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n7155) );
  NOR2_X1 U8045 ( .A1(n7154), .A2(n7155), .ZN(n7153) );
  INV_X1 U8046 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n8066) );
  MUX2_X1 U8047 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n8066), .S(n7172), .Z(n7165)
         );
  NOR2_X1 U8048 ( .A1(n7166), .A2(n7165), .ZN(n7164) );
  XOR2_X1 U8049 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7225), .Z(n7213) );
  XNOR2_X1 U8050 ( .A(n6350), .B(P2_REG2_REG_5__SCAN_IN), .ZN(n7251) );
  NOR2_X1 U8051 ( .A1(n7252), .A2(n7251), .ZN(n7250) );
  XNOR2_X1 U8052 ( .A(n6966), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n7226) );
  XNOR2_X1 U8053 ( .A(n6365), .B(P2_REG2_REG_7__SCAN_IN), .ZN(n7238) );
  MUX2_X1 U8054 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n7841), .S(n7279), .Z(n6254)
         );
  INV_X1 U8055 ( .A(n6254), .ZN(n7275) );
  XNOR2_X1 U8056 ( .A(n6976), .B(P2_REG2_REG_9__SCAN_IN), .ZN(n7496) );
  XNOR2_X1 U8057 ( .A(n6395), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n7676) );
  INV_X1 U8058 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6255) );
  MUX2_X1 U8059 ( .A(n6255), .B(P2_REG2_REG_11__SCAN_IN), .S(n6990), .Z(n6256)
         );
  INV_X1 U8060 ( .A(n6256), .ZN(n7810) );
  XNOR2_X1 U8061 ( .A(n6994), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n8033) );
  XOR2_X1 U8062 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n7011), .Z(n8426) );
  XOR2_X1 U8063 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n7062), .Z(n8441) );
  NAND2_X1 U8064 ( .A1(n6473), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6258) );
  OAI21_X1 U8065 ( .B1(n6473), .B2(P2_REG2_REG_17__SCAN_IN), .A(n6258), .ZN(
        n8476) );
  INV_X1 U8066 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8495) );
  NAND2_X1 U8067 ( .A1(n8496), .A2(n8495), .ZN(n8494) );
  INV_X1 U8068 ( .A(n7351), .ZN(n8500) );
  NAND2_X1 U8069 ( .A1(n6259), .A2(n8500), .ZN(n6260) );
  NAND2_X1 U8070 ( .A1(n8494), .A2(n6260), .ZN(n6261) );
  INV_X1 U8071 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n9881) );
  XNOR2_X1 U8072 ( .A(n6261), .B(n9881), .ZN(n6272) );
  NAND2_X1 U8073 ( .A1(n6262), .A2(n6319), .ZN(n6263) );
  NAND2_X1 U8074 ( .A1(n6263), .A2(n8422), .ZN(n6266) );
  NOR2_X1 U8075 ( .A1(n8969), .A2(n8971), .ZN(n6265) );
  NAND2_X1 U8076 ( .A1(n6268), .A2(n6267), .ZN(n6611) );
  NAND2_X1 U8077 ( .A1(n6611), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6269) );
  INV_X1 U8078 ( .A(n6270), .ZN(n6271) );
  INV_X1 U8079 ( .A(n10303), .ZN(n6274) );
  AOI21_X1 U8080 ( .B1(n10303), .B2(n7759), .A(n6319), .ZN(n6273) );
  AOI21_X1 U8081 ( .B1(n6275), .B2(n6274), .A(n6273), .ZN(n8491) );
  NAND2_X1 U8082 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n6277) );
  INV_X1 U8083 ( .A(n6279), .ZN(n6280) );
  NAND2_X1 U8084 ( .A1(n6280), .A2(SI_29_), .ZN(n6281) );
  INV_X1 U8085 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8156) );
  INV_X1 U8086 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10084) );
  MUX2_X1 U8087 ( .A(n8156), .B(n10084), .S(n4271), .Z(n6284) );
  INV_X1 U8088 ( .A(SI_30_), .ZN(n6283) );
  NAND2_X1 U8089 ( .A1(n6284), .A2(n6283), .ZN(n6602) );
  INV_X1 U8090 ( .A(n6284), .ZN(n6285) );
  NAND2_X1 U8091 ( .A1(n6285), .A2(SI_30_), .ZN(n6286) );
  NAND2_X1 U8092 ( .A1(n6602), .A2(n6286), .ZN(n6603) );
  NAND2_X1 U8093 ( .A1(n6319), .A2(n6950), .ZN(n6322) );
  INV_X2 U8094 ( .A(n6322), .ZN(n6328) );
  NAND2_X4 U8095 ( .A1(n6319), .A2(n4271), .ZN(n6607) );
  OR2_X1 U8096 ( .A1(n6607), .A2(n8156), .ZN(n6287) );
  OR2_X1 U8097 ( .A1(n6322), .A2(n6955), .ZN(n6289) );
  INV_X1 U8098 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6949) );
  NAND2_X1 U8099 ( .A1(n6292), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6295) );
  OAI21_X1 U8100 ( .B1(n6295), .B2(n6291), .A(n6294), .ZN(n6296) );
  NOR2_X2 U8101 ( .A1(n4310), .A2(n6296), .ZN(n6298) );
  INV_X1 U8102 ( .A(n8155), .ZN(n6299) );
  AND2_X2 U8103 ( .A1(n6298), .A2(n6299), .ZN(n6332) );
  NAND2_X1 U8104 ( .A1(n6332), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6302) );
  INV_X1 U8105 ( .A(n6298), .ZN(n8967) );
  NAND2_X1 U8106 ( .A1(n6345), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6301) );
  NAND2_X1 U8107 ( .A1(n10285), .A2(n6304), .ZN(n6636) );
  NAND2_X1 U8108 ( .A1(n6311), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6308) );
  NAND2_X1 U8109 ( .A1(n6341), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6307) );
  NAND2_X1 U8110 ( .A1(n6332), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6306) );
  NAND2_X1 U8111 ( .A1(n6345), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6305) );
  NAND2_X1 U8112 ( .A1(n6950), .A2(SI_0_), .ZN(n6309) );
  XNOR2_X1 U8113 ( .A(n6309), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8979) );
  NAND2_X1 U8114 ( .A1(n7314), .A2(n10313), .ZN(n10288) );
  NAND2_X1 U8115 ( .A1(n10293), .A2(n10287), .ZN(n7335) );
  NAND2_X1 U8116 ( .A1(n6311), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6315) );
  NAND2_X1 U8117 ( .A1(n6341), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6314) );
  NAND2_X1 U8118 ( .A1(n6332), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6313) );
  NAND2_X1 U8119 ( .A1(n6345), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6312) );
  INV_X1 U8120 ( .A(n6778), .ZN(n6318) );
  OR2_X1 U8121 ( .A1(n6322), .A2(n6957), .ZN(n6317) );
  OAI211_X2 U8122 ( .C1(n6319), .C2(n7172), .A(n6317), .B(n6316), .ZN(n8090)
         );
  NAND2_X1 U8123 ( .A1(n6778), .A2(n8090), .ZN(n6641) );
  OR2_X1 U8124 ( .A1(n6319), .A2(n7211), .ZN(n6321) );
  OR2_X1 U8125 ( .A1(n6607), .A2(n4930), .ZN(n6320) );
  INV_X1 U8126 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6334) );
  NAND2_X1 U8127 ( .A1(n6332), .A2(n6334), .ZN(n6325) );
  NAND2_X1 U8128 ( .A1(n6341), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6324) );
  NAND2_X1 U8129 ( .A1(n6345), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6323) );
  NAND2_X1 U8130 ( .A1(n6311), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6326) );
  NAND2_X1 U8131 ( .A1(n7652), .A2(n8421), .ZN(n6646) );
  NAND2_X1 U8132 ( .A1(n6783), .A2(n10272), .ZN(n6644) );
  NAND2_X1 U8133 ( .A1(n6328), .A2(n6951), .ZN(n6331) );
  OR2_X1 U8134 ( .A1(n6319), .A2(n7225), .ZN(n6330) );
  OR2_X1 U8135 ( .A1(n6607), .A2(n5322), .ZN(n6329) );
  INV_X1 U8136 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6333) );
  NAND2_X1 U8137 ( .A1(n6334), .A2(n6333), .ZN(n6335) );
  AND2_X1 U8138 ( .A1(n6335), .A2(n6343), .ZN(n8311) );
  NAND2_X1 U8139 ( .A1(n6332), .A2(n8311), .ZN(n6339) );
  NAND2_X1 U8140 ( .A1(n6341), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6338) );
  NAND2_X1 U8141 ( .A1(n6345), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6337) );
  NAND2_X1 U8142 ( .A1(n6311), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6336) );
  INV_X1 U8143 ( .A(n6628), .ZN(n6645) );
  NAND2_X1 U8144 ( .A1(n8420), .A2(n7569), .ZN(n7575) );
  NAND2_X1 U8145 ( .A1(n6568), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6349) );
  NAND2_X1 U8146 ( .A1(n6341), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6348) );
  INV_X1 U8147 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6342) );
  NAND2_X1 U8148 ( .A1(n6343), .A2(n6342), .ZN(n6344) );
  AND2_X1 U8149 ( .A1(n6356), .A2(n6344), .ZN(n8276) );
  NAND2_X1 U8150 ( .A1(n6332), .A2(n8276), .ZN(n6347) );
  NAND2_X1 U8151 ( .A1(n6345), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6346) );
  NAND2_X1 U8152 ( .A1(n6958), .A2(n6328), .ZN(n6352) );
  AOI22_X1 U8153 ( .A1(n6485), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6484), .B2(
        n6350), .ZN(n6351) );
  NAND2_X1 U8154 ( .A1(n8419), .A2(n7802), .ZN(n6630) );
  INV_X1 U8155 ( .A(n8419), .ZN(n8078) );
  NAND2_X1 U8156 ( .A1(n6353), .A2(n6648), .ZN(n7737) );
  NAND2_X1 U8157 ( .A1(n6568), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6361) );
  NAND2_X1 U8158 ( .A1(n6599), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6360) );
  INV_X1 U8159 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6355) );
  NAND2_X1 U8160 ( .A1(n6356), .A2(n6355), .ZN(n6357) );
  AND2_X1 U8161 ( .A1(n6369), .A2(n6357), .ZN(n8071) );
  NAND2_X1 U8162 ( .A1(n6573), .A2(n8071), .ZN(n6359) );
  NAND2_X1 U8163 ( .A1(n6345), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6358) );
  NAND2_X1 U8164 ( .A1(n6965), .A2(n6328), .ZN(n6363) );
  AOI22_X1 U8165 ( .A1(n6485), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6484), .B2(
        n6966), .ZN(n6362) );
  NAND2_X1 U8166 ( .A1(n6363), .A2(n6362), .ZN(n7750) );
  NAND2_X1 U8167 ( .A1(n7580), .A2(n7750), .ZN(n6657) );
  INV_X1 U8168 ( .A(n7580), .ZN(n8418) );
  NAND2_X1 U8169 ( .A1(n10327), .A2(n8418), .ZN(n6651) );
  INV_X1 U8170 ( .A(n6657), .ZN(n6364) );
  NAND2_X1 U8171 ( .A1(n6973), .A2(n6328), .ZN(n6367) );
  AOI22_X1 U8172 ( .A1(n6485), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6484), .B2(
        n6365), .ZN(n6366) );
  NAND2_X1 U8173 ( .A1(n6367), .A2(n6366), .ZN(n7828) );
  INV_X4 U8174 ( .A(n6368), .ZN(n6568) );
  NAND2_X1 U8175 ( .A1(n6568), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6374) );
  NAND2_X1 U8176 ( .A1(n6599), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6373) );
  NAND2_X1 U8177 ( .A1(n6369), .A2(n9937), .ZN(n6370) );
  AND2_X1 U8178 ( .A1(n6377), .A2(n6370), .ZN(n7820) );
  NAND2_X1 U8179 ( .A1(n6573), .A2(n7820), .ZN(n6372) );
  NAND2_X1 U8180 ( .A1(n6345), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6371) );
  NAND2_X1 U8181 ( .A1(n7828), .A2(n8206), .ZN(n6658) );
  OR2_X1 U8182 ( .A1(n8206), .A2(n7828), .ZN(n6659) );
  NAND2_X1 U8183 ( .A1(n6568), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6382) );
  NAND2_X1 U8184 ( .A1(n6599), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6381) );
  NAND2_X1 U8185 ( .A1(n6377), .A2(n6376), .ZN(n6378) );
  NAND2_X1 U8186 ( .A1(n6389), .A2(n6378), .ZN(n7844) );
  INV_X1 U8187 ( .A(n7844), .ZN(n8209) );
  NAND2_X1 U8188 ( .A1(n6573), .A2(n8209), .ZN(n6380) );
  NAND2_X1 U8189 ( .A1(n6345), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6379) );
  NAND2_X1 U8190 ( .A1(n6960), .A2(n6328), .ZN(n6384) );
  AOI22_X1 U8191 ( .A1(n6485), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6484), .B2(
        n7279), .ZN(n6383) );
  OR2_X1 U8192 ( .A1(n7893), .A2(n10337), .ZN(n6662) );
  NAND2_X1 U8193 ( .A1(n10337), .A2(n7893), .ZN(n6663) );
  NAND2_X1 U8194 ( .A1(n6662), .A2(n6663), .ZN(n7834) );
  NAND2_X1 U8195 ( .A1(n6969), .A2(n6328), .ZN(n6387) );
  AOI22_X1 U8196 ( .A1(n6485), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6484), .B2(
        n6976), .ZN(n6386) );
  NAND2_X1 U8197 ( .A1(n6568), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6394) );
  NAND2_X1 U8198 ( .A1(n6599), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6393) );
  INV_X1 U8199 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6388) );
  NAND2_X1 U8200 ( .A1(n6389), .A2(n6388), .ZN(n6390) );
  AND2_X1 U8201 ( .A1(n6405), .A2(n6390), .ZN(n7904) );
  NAND2_X1 U8202 ( .A1(n6573), .A2(n7904), .ZN(n6392) );
  NAND2_X1 U8203 ( .A1(n6345), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6391) );
  OR2_X1 U8204 ( .A1(n8891), .A2(n7927), .ZN(n6673) );
  NAND2_X1 U8205 ( .A1(n8891), .A2(n7927), .ZN(n6668) );
  NAND2_X1 U8206 ( .A1(n6979), .A2(n6328), .ZN(n6397) );
  AOI22_X1 U8207 ( .A1(n6485), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6395), .B2(
        n6484), .ZN(n6396) );
  NAND2_X1 U8208 ( .A1(n6568), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6401) );
  NAND2_X1 U8209 ( .A1(n6599), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6400) );
  XNOR2_X1 U8210 ( .A(n6405), .B(P2_REG3_REG_10__SCAN_IN), .ZN(n7938) );
  NAND2_X1 U8211 ( .A1(n6573), .A2(n7938), .ZN(n6399) );
  NAND2_X1 U8212 ( .A1(n6345), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6398) );
  NAND2_X1 U8213 ( .A1(n6988), .A2(n6328), .ZN(n6403) );
  AOI22_X1 U8214 ( .A1(n6990), .A2(n6484), .B1(n6485), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n6402) );
  NAND2_X1 U8215 ( .A1(n6403), .A2(n6402), .ZN(n8751) );
  NAND2_X1 U8216 ( .A1(n6568), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6410) );
  NAND2_X1 U8217 ( .A1(n6599), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6409) );
  OAI21_X1 U8218 ( .B1(n6405), .B2(n6404), .A(n7976), .ZN(n6406) );
  AND2_X1 U8219 ( .A1(n6406), .A2(n6414), .ZN(n8752) );
  NAND2_X1 U8220 ( .A1(n6573), .A2(n8752), .ZN(n6408) );
  NAND2_X1 U8221 ( .A1(n6345), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6407) );
  NAND2_X1 U8222 ( .A1(n8751), .A2(n8232), .ZN(n6680) );
  NAND2_X1 U8223 ( .A1(n8887), .A2(n7973), .ZN(n8755) );
  AND2_X1 U8224 ( .A1(n6680), .A2(n8755), .ZN(n6671) );
  OR2_X1 U8225 ( .A1(n8751), .A2(n8232), .ZN(n6679) );
  NAND2_X1 U8226 ( .A1(n6992), .A2(n6328), .ZN(n6412) );
  AOI22_X1 U8227 ( .A1(n6485), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6994), .B2(
        n6484), .ZN(n6411) );
  NAND2_X1 U8228 ( .A1(n6568), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6419) );
  NAND2_X1 U8229 ( .A1(n6599), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6418) );
  INV_X1 U8230 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8029) );
  NAND2_X1 U8231 ( .A1(n6414), .A2(n8029), .ZN(n6415) );
  AND2_X1 U8232 ( .A1(n6423), .A2(n6415), .ZN(n8235) );
  NAND2_X1 U8233 ( .A1(n6573), .A2(n8235), .ZN(n6417) );
  NAND2_X1 U8234 ( .A1(n6345), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6416) );
  NAND2_X1 U8235 ( .A1(n8243), .A2(n7997), .ZN(n6684) );
  INV_X1 U8236 ( .A(n7994), .ZN(n6430) );
  NAND2_X1 U8237 ( .A1(n7009), .A2(n6328), .ZN(n6421) );
  AOI22_X1 U8238 ( .A1(n7011), .A2(n6484), .B1(n6485), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n6420) );
  NAND2_X1 U8239 ( .A1(n6568), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6428) );
  NAND2_X1 U8240 ( .A1(n6599), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6427) );
  INV_X1 U8241 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6422) );
  NAND2_X1 U8242 ( .A1(n6423), .A2(n6422), .ZN(n6424) );
  AND2_X1 U8243 ( .A1(n6435), .A2(n6424), .ZN(n8332) );
  NAND2_X1 U8244 ( .A1(n6573), .A2(n8332), .ZN(n6426) );
  NAND2_X1 U8245 ( .A1(n6345), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6425) );
  XNOR2_X1 U8246 ( .A(n8946), .B(n8171), .ZN(n7993) );
  NAND2_X1 U8247 ( .A1(n8946), .A2(n8171), .ZN(n6431) );
  NAND2_X1 U8248 ( .A1(n7060), .A2(n6328), .ZN(n6433) );
  AOI22_X1 U8249 ( .A1(n7062), .A2(n6484), .B1(n6485), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n6432) );
  NAND2_X1 U8250 ( .A1(n6568), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6440) );
  NAND2_X1 U8251 ( .A1(n6599), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6439) );
  INV_X1 U8252 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9891) );
  NAND2_X1 U8253 ( .A1(n6435), .A2(n9891), .ZN(n6436) );
  AND2_X1 U8254 ( .A1(n6447), .A2(n6436), .ZN(n8740) );
  NAND2_X1 U8255 ( .A1(n6573), .A2(n8740), .ZN(n6438) );
  NAND2_X1 U8256 ( .A1(n6345), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6437) );
  XNOR2_X1 U8257 ( .A(n8739), .B(n8384), .ZN(n8732) );
  INV_X1 U8258 ( .A(n8732), .ZN(n6441) );
  OR2_X1 U8259 ( .A1(n8739), .A2(n8384), .ZN(n6688) );
  NAND2_X1 U8260 ( .A1(n6442), .A2(n6688), .ZN(n8712) );
  NAND2_X1 U8261 ( .A1(n7119), .A2(n6328), .ZN(n6445) );
  AOI22_X1 U8262 ( .A1(n6443), .A2(n6484), .B1(n6485), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n6444) );
  NAND2_X2 U8263 ( .A1(n6445), .A2(n6444), .ZN(n8938) );
  INV_X1 U8264 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6446) );
  NAND2_X1 U8265 ( .A1(n6447), .A2(n6446), .ZN(n6448) );
  AND2_X1 U8266 ( .A1(n6457), .A2(n6448), .ZN(n8717) );
  NAND2_X1 U8267 ( .A1(n8717), .A2(n6332), .ZN(n6452) );
  NAND2_X1 U8268 ( .A1(n6568), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6451) );
  NAND2_X1 U8269 ( .A1(n6599), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6450) );
  NAND2_X1 U8270 ( .A1(n6345), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6449) );
  NAND2_X1 U8271 ( .A1(n8938), .A2(n8117), .ZN(n6701) );
  NAND2_X1 U8272 ( .A1(n8712), .A2(n6701), .ZN(n6453) );
  OR2_X1 U8273 ( .A1(n8938), .A2(n8117), .ZN(n6694) );
  NAND2_X1 U8274 ( .A1(n6453), .A2(n6694), .ZN(n8695) );
  NAND2_X1 U8275 ( .A1(n7148), .A2(n6328), .ZN(n6456) );
  AOI22_X1 U8276 ( .A1(n6454), .A2(n6484), .B1(n6485), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n6455) );
  NAND2_X1 U8277 ( .A1(n6457), .A2(n4679), .ZN(n6458) );
  NAND2_X1 U8278 ( .A1(n6476), .A2(n6458), .ZN(n8706) );
  OR2_X1 U8279 ( .A1(n8706), .A2(n6561), .ZN(n6463) );
  NAND2_X1 U8280 ( .A1(n6599), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6460) );
  NAND2_X1 U8281 ( .A1(n6568), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6459) );
  AND2_X1 U8282 ( .A1(n6460), .A2(n6459), .ZN(n6462) );
  NAND2_X1 U8283 ( .A1(n6345), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6461) );
  NAND2_X1 U8284 ( .A1(n7349), .A2(n6328), .ZN(n6465) );
  AOI22_X1 U8285 ( .A1(n6485), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6484), .B2(
        n7351), .ZN(n6464) );
  INV_X1 U8286 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8291) );
  INV_X1 U8287 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n6466) );
  OAI21_X1 U8288 ( .B1(n6476), .B2(n8291), .A(n6466), .ZN(n6469) );
  INV_X1 U8289 ( .A(n6476), .ZN(n6468) );
  AND2_X1 U8290 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .ZN(n6467) );
  INV_X1 U8291 ( .A(n6488), .ZN(n6490) );
  AND2_X1 U8292 ( .A1(n6469), .A2(n6490), .ZN(n8672) );
  NAND2_X1 U8293 ( .A1(n8672), .A2(n6573), .ZN(n6472) );
  AOI22_X1 U8294 ( .A1(n6599), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n6568), .B2(
        P2_REG2_REG_18__SCAN_IN), .ZN(n6471) );
  NAND2_X1 U8295 ( .A1(n6345), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6470) );
  NAND2_X1 U8296 ( .A1(n8926), .A2(n8288), .ZN(n8645) );
  NAND2_X1 U8297 ( .A1(n7307), .A2(n6328), .ZN(n6475) );
  AOI22_X1 U8298 ( .A1(n6485), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6484), .B2(
        n6473), .ZN(n6474) );
  NAND2_X2 U8299 ( .A1(n6475), .A2(n6474), .ZN(n8930) );
  XNOR2_X1 U8300 ( .A(n6476), .B(P2_REG3_REG_17__SCAN_IN), .ZN(n8690) );
  NAND2_X1 U8301 ( .A1(n8690), .A2(n6573), .ZN(n6482) );
  NAND2_X1 U8302 ( .A1(n6568), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6478) );
  NAND2_X1 U8303 ( .A1(n6345), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6477) );
  OAI211_X1 U8304 ( .C1(n6354), .C2(n6479), .A(n6478), .B(n6477), .ZN(n6480)
         );
  INV_X1 U8305 ( .A(n6480), .ZN(n6481) );
  NAND2_X1 U8306 ( .A1(n8930), .A2(n8358), .ZN(n6483) );
  NAND2_X1 U8307 ( .A1(n8645), .A2(n6483), .ZN(n6698) );
  NAND2_X1 U8308 ( .A1(n7451), .A2(n6328), .ZN(n6487) );
  AOI22_X1 U8309 ( .A1(n6485), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6484), .B2(
        n7344), .ZN(n6486) );
  INV_X1 U8310 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6489) );
  NAND2_X1 U8311 ( .A1(n6490), .A2(n6489), .ZN(n6491) );
  NAND2_X1 U8312 ( .A1(n6501), .A2(n6491), .ZN(n8654) );
  OR2_X1 U8313 ( .A1(n8654), .A2(n6561), .ZN(n6496) );
  NAND2_X1 U8314 ( .A1(n6599), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6493) );
  NAND2_X1 U8315 ( .A1(n6345), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6492) );
  OAI211_X1 U8316 ( .C1(n6368), .C2(n9881), .A(n6493), .B(n6492), .ZN(n6494)
         );
  INV_X1 U8317 ( .A(n6494), .ZN(n6495) );
  OR2_X1 U8318 ( .A1(n8834), .A2(n8199), .ZN(n6704) );
  NAND2_X1 U8319 ( .A1(n8834), .A2(n8199), .ZN(n6714) );
  OR2_X1 U8320 ( .A1(n8926), .A2(n8288), .ZN(n6697) );
  OR2_X1 U8321 ( .A1(n8930), .A2(n8358), .ZN(n8661) );
  NAND2_X1 U8322 ( .A1(n6697), .A2(n8661), .ZN(n6497) );
  NAND2_X1 U8323 ( .A1(n6497), .A2(n8645), .ZN(n6498) );
  NAND2_X1 U8324 ( .A1(n7518), .A2(n6328), .ZN(n6500) );
  OR2_X1 U8325 ( .A1(n6607), .A2(n9938), .ZN(n6499) );
  INV_X1 U8326 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8327) );
  NAND2_X1 U8327 ( .A1(n6501), .A2(n8327), .ZN(n6502) );
  NAND2_X1 U8328 ( .A1(n6510), .A2(n6502), .ZN(n8323) );
  OR2_X1 U8329 ( .A1(n8323), .A2(n6561), .ZN(n6507) );
  INV_X1 U8330 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8920) );
  NAND2_X1 U8331 ( .A1(n6599), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6504) );
  NAND2_X1 U8332 ( .A1(n6568), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6503) );
  OAI211_X1 U8333 ( .C1(n8920), .C2(n6542), .A(n6504), .B(n6503), .ZN(n6505)
         );
  INV_X1 U8334 ( .A(n6505), .ZN(n6506) );
  NAND2_X1 U8335 ( .A1(n8634), .A2(n8223), .ZN(n6715) );
  NAND2_X1 U8336 ( .A1(n6718), .A2(n6715), .ZN(n8628) );
  NAND2_X1 U8337 ( .A1(n7586), .A2(n6328), .ZN(n6509) );
  OR2_X1 U8338 ( .A1(n6607), .A2(n7610), .ZN(n6508) );
  NAND2_X2 U8339 ( .A1(n6509), .A2(n6508), .ZN(n8823) );
  INV_X1 U8340 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8225) );
  NAND2_X1 U8341 ( .A1(n6510), .A2(n8225), .ZN(n6511) );
  AND2_X1 U8342 ( .A1(n6518), .A2(n6511), .ZN(n8616) );
  INV_X1 U8343 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9967) );
  NAND2_X1 U8344 ( .A1(n6568), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6513) );
  NAND2_X1 U8345 ( .A1(n6345), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6512) );
  OAI211_X1 U8346 ( .C1(n6354), .C2(n9967), .A(n6513), .B(n6512), .ZN(n6514)
         );
  XNOR2_X1 U8347 ( .A(n8823), .B(n8346), .ZN(n8619) );
  NAND2_X1 U8348 ( .A1(n8823), .A2(n8346), .ZN(n6722) );
  NAND2_X1 U8349 ( .A1(n7734), .A2(n6328), .ZN(n6517) );
  OR2_X1 U8350 ( .A1(n6607), .A2(n8101), .ZN(n6516) );
  INV_X1 U8351 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8348) );
  NAND2_X1 U8352 ( .A1(n6518), .A2(n8348), .ZN(n6519) );
  NAND2_X1 U8353 ( .A1(n6528), .A2(n6519), .ZN(n8345) );
  INV_X1 U8354 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8915) );
  NAND2_X1 U8355 ( .A1(n6599), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6521) );
  NAND2_X1 U8356 ( .A1(n6568), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6520) );
  OAI211_X1 U8357 ( .C1(n8915), .C2(n6542), .A(n6521), .B(n6520), .ZN(n6522)
         );
  INV_X1 U8358 ( .A(n6522), .ZN(n6523) );
  NAND2_X1 U8359 ( .A1(n8604), .A2(n8224), .ZN(n6721) );
  NAND2_X1 U8360 ( .A1(n7758), .A2(n6328), .ZN(n6526) );
  OR2_X1 U8361 ( .A1(n6607), .A2(n7761), .ZN(n6525) );
  INV_X1 U8362 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8185) );
  NAND2_X1 U8363 ( .A1(n6528), .A2(n8185), .ZN(n6529) );
  NAND2_X1 U8364 ( .A1(n6548), .A2(n6529), .ZN(n8590) );
  INV_X1 U8365 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n6532) );
  NAND2_X1 U8366 ( .A1(n6599), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6531) );
  NAND2_X1 U8367 ( .A1(n6568), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6530) );
  OAI211_X1 U8368 ( .C1(n6532), .C2(n6542), .A(n6531), .B(n6530), .ZN(n6533)
         );
  INV_X1 U8369 ( .A(n6533), .ZN(n6534) );
  OR2_X1 U8370 ( .A1(n8813), .A2(n6874), .ZN(n6712) );
  NAND2_X1 U8371 ( .A1(n8813), .A2(n6874), .ZN(n6536) );
  INV_X1 U8372 ( .A(n8583), .ZN(n6707) );
  NOR2_X1 U8373 ( .A1(n8587), .A2(n6707), .ZN(n6537) );
  INV_X1 U8374 ( .A(n6536), .ZN(n6727) );
  NAND2_X1 U8375 ( .A1(n7923), .A2(n6328), .ZN(n6539) );
  OR2_X1 U8376 ( .A1(n6607), .A2(n7924), .ZN(n6538) );
  XNOR2_X1 U8377 ( .A(n6548), .B(P2_REG3_REG_24__SCAN_IN), .ZN(n8576) );
  INV_X1 U8378 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8910) );
  NAND2_X1 U8379 ( .A1(n6599), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6541) );
  NAND2_X1 U8380 ( .A1(n6568), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6540) );
  OAI211_X1 U8381 ( .C1(n8910), .C2(n6542), .A(n6541), .B(n6540), .ZN(n6543)
         );
  NAND2_X1 U8382 ( .A1(n8575), .A2(n8299), .ZN(n6726) );
  NAND2_X1 U8383 ( .A1(n8022), .A2(n6328), .ZN(n6545) );
  OR2_X1 U8384 ( .A1(n6607), .A2(n9863), .ZN(n6544) );
  INV_X1 U8385 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8304) );
  INV_X1 U8386 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6546) );
  OAI21_X1 U8387 ( .B1(n6548), .B2(n8304), .A(n6546), .ZN(n6549) );
  NAND2_X1 U8388 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_REG3_REG_24__SCAN_IN), 
        .ZN(n6547) );
  INV_X1 U8389 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n6552) );
  NAND2_X1 U8390 ( .A1(n6599), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6551) );
  NAND2_X1 U8391 ( .A1(n6568), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6550) );
  OAI211_X1 U8392 ( .C1(n6542), .C2(n6552), .A(n6551), .B(n6550), .ZN(n6553)
         );
  NAND2_X1 U8393 ( .A1(n8802), .A2(n8368), .ZN(n6732) );
  NAND2_X1 U8394 ( .A1(n8049), .A2(n6328), .ZN(n6556) );
  OR2_X1 U8395 ( .A1(n6607), .A2(n8975), .ZN(n6555) );
  INV_X1 U8396 ( .A(n6559), .ZN(n6557) );
  INV_X1 U8397 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n6558) );
  NAND2_X1 U8398 ( .A1(n6559), .A2(n6558), .ZN(n6560) );
  NAND2_X1 U8399 ( .A1(n6580), .A2(n6560), .ZN(n8371) );
  INV_X1 U8400 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8906) );
  NAND2_X1 U8401 ( .A1(n6599), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6563) );
  NAND2_X1 U8402 ( .A1(n6568), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6562) );
  OAI211_X1 U8403 ( .C1(n8906), .C2(n6542), .A(n6563), .B(n6562), .ZN(n6564)
         );
  INV_X1 U8404 ( .A(n6564), .ZN(n6565) );
  NOR2_X1 U8405 ( .A1(n8543), .A2(n8129), .ZN(n6736) );
  OR2_X1 U8406 ( .A1(n6607), .A2(n8973), .ZN(n6567) );
  INV_X1 U8407 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n6571) );
  NAND2_X1 U8408 ( .A1(n6599), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6570) );
  NAND2_X1 U8409 ( .A1(n6568), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6569) );
  OAI211_X1 U8410 ( .C1(n6571), .C2(n6542), .A(n6570), .B(n6569), .ZN(n6572)
         );
  NAND2_X1 U8411 ( .A1(n8793), .A2(n8367), .ZN(n6739) );
  INV_X1 U8412 ( .A(n6737), .ZN(n8521) );
  NAND2_X1 U8413 ( .A1(n8152), .A2(n6328), .ZN(n6576) );
  OR2_X1 U8414 ( .A1(n6607), .A2(n8970), .ZN(n6575) );
  INV_X1 U8415 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6578) );
  INV_X1 U8416 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6577) );
  OAI21_X1 U8417 ( .B1(n6580), .B2(n6578), .A(n6577), .ZN(n6581) );
  NAND2_X1 U8418 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n6579) );
  NAND2_X1 U8419 ( .A1(n8510), .A2(n6573), .ZN(n6586) );
  INV_X1 U8420 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9952) );
  NAND2_X1 U8421 ( .A1(n6568), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6583) );
  NAND2_X1 U8422 ( .A1(n6345), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6582) );
  OAI211_X1 U8423 ( .C1(n6354), .C2(n9952), .A(n6583), .B(n6582), .ZN(n6584)
         );
  INV_X1 U8424 ( .A(n6584), .ZN(n6585) );
  INV_X1 U8425 ( .A(n8397), .ZN(n6743) );
  NAND2_X1 U8426 ( .A1(n8965), .A2(n6328), .ZN(n6590) );
  OR2_X1 U8427 ( .A1(n6607), .A2(n8966), .ZN(n6589) );
  INV_X1 U8428 ( .A(n6591), .ZN(n8133) );
  INV_X1 U8429 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6594) );
  NAND2_X1 U8430 ( .A1(n6599), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6593) );
  NAND2_X1 U8431 ( .A1(n6568), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6592) );
  OAI211_X1 U8432 ( .C1(n6594), .C2(n6542), .A(n6593), .B(n6592), .ZN(n6595)
         );
  AOI21_X1 U8433 ( .B1(n8133), .B2(n6573), .A(n6595), .ZN(n7467) );
  NAND2_X1 U8434 ( .A1(n6568), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6598) );
  NAND2_X1 U8435 ( .A1(n6599), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6597) );
  NAND2_X1 U8436 ( .A1(n6345), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6596) );
  AND3_X1 U8437 ( .A1(n6598), .A2(n6597), .A3(n6596), .ZN(n8107) );
  INV_X1 U8438 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8898) );
  NAND2_X1 U8439 ( .A1(n6599), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6601) );
  NAND2_X1 U8440 ( .A1(n6568), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6600) );
  OAI211_X1 U8441 ( .C1(n6542), .C2(n8898), .A(n6601), .B(n6600), .ZN(n8104)
         );
  INV_X1 U8442 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8964) );
  INV_X1 U8443 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10076) );
  MUX2_X1 U8444 ( .A(n8964), .B(n10076), .S(n4271), .Z(n6605) );
  XNOR2_X1 U8445 ( .A(n6605), .B(SI_31_), .ZN(n6606) );
  NOR2_X1 U8446 ( .A1(n6607), .A2(n8964), .ZN(n6608) );
  NAND2_X1 U8447 ( .A1(n8504), .A2(n8107), .ZN(n6751) );
  AOI21_X1 U8448 ( .B1(n6609), .B2(n6754), .A(n6757), .ZN(n6610) );
  OAI21_X1 U8449 ( .B1(n6611), .B2(P2_IR_REG_19__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6612) );
  MUX2_X1 U8450 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6612), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n6614) );
  INV_X1 U8451 ( .A(n6915), .ZN(n10314) );
  NOR2_X1 U8452 ( .A1(n7313), .A2(n7334), .ZN(n6761) );
  INV_X1 U8453 ( .A(n8628), .ZN(n8123) );
  INV_X1 U8454 ( .A(n8641), .ZN(n8646) );
  NAND2_X1 U8455 ( .A1(n6697), .A2(n8645), .ZN(n8662) );
  INV_X1 U8456 ( .A(n8358), .ZN(n8408) );
  INV_X1 U8457 ( .A(n8685), .ZN(n8679) );
  INV_X1 U8458 ( .A(n7314), .ZN(n8423) );
  INV_X1 U8459 ( .A(n10313), .ZN(n7886) );
  NAND2_X1 U8460 ( .A1(n8423), .A2(n7886), .ZN(n6638) );
  NAND2_X1 U8461 ( .A1(n10288), .A2(n6638), .ZN(n10315) );
  NOR4_X1 U8462 ( .A1(n7339), .A2(n10315), .A3(n7338), .A4(n7719), .ZN(n6617)
         );
  NAND3_X1 U8463 ( .A1(n6617), .A2(n7599), .A3(n7564), .ZN(n6618) );
  INV_X1 U8464 ( .A(n7738), .ZN(n7741) );
  NAND2_X1 U8465 ( .A1(n6648), .A2(n6630), .ZN(n7577) );
  NOR4_X1 U8466 ( .A1(n6618), .A2(n7741), .A3(n7834), .A4(n7577), .ZN(n6619)
         );
  NAND4_X1 U8467 ( .A1(n6619), .A2(n7899), .A3(n7930), .A4(n7547), .ZN(n6620)
         );
  NAND2_X1 U8468 ( .A1(n6679), .A2(n6680), .ZN(n8757) );
  NOR4_X1 U8469 ( .A1(n6620), .A2(n7993), .A3(n5128), .A4(n8757), .ZN(n6621)
         );
  NAND4_X1 U8470 ( .A1(n8700), .A2(n8721), .A3(n6621), .A4(n6441), .ZN(n6622)
         );
  NOR4_X1 U8471 ( .A1(n8646), .A2(n8662), .A3(n8679), .A4(n6622), .ZN(n6623)
         );
  NAND4_X1 U8472 ( .A1(n8598), .A2(n8123), .A3(n6623), .A4(n6515), .ZN(n6624)
         );
  NOR4_X1 U8473 ( .A1(n8125), .A2(n8568), .A3(n8587), .A4(n6624), .ZN(n6625)
         );
  INV_X1 U8474 ( .A(n6626), .ZN(n7333) );
  NAND2_X1 U8475 ( .A1(n7344), .A2(n6639), .ZN(n7718) );
  AOI22_X1 U8476 ( .A1(n6649), .A2(n6630), .B1(n6629), .B2(n6646), .ZN(n6632)
         );
  INV_X1 U8477 ( .A(n6651), .ZN(n6631) );
  NOR2_X1 U8478 ( .A1(n6632), .A2(n6631), .ZN(n6655) );
  NAND2_X1 U8479 ( .A1(n10287), .A2(n6633), .ZN(n6642) );
  INV_X1 U8480 ( .A(n6642), .ZN(n6634) );
  NAND2_X1 U8481 ( .A1(n6634), .A2(n6638), .ZN(n6635) );
  OAI211_X1 U8482 ( .C1(n6636), .C2(n6642), .A(n6635), .B(n6641), .ZN(n6637)
         );
  AOI21_X1 U8483 ( .B1(n6639), .B2(n6638), .A(n10293), .ZN(n6643) );
  OAI211_X1 U8484 ( .C1(n6643), .C2(n6642), .A(n6641), .B(n6640), .ZN(n6647)
         );
  AOI211_X1 U8485 ( .C1(n6647), .C2(n6646), .A(n6645), .B(n5160), .ZN(n6650)
         );
  OAI211_X1 U8486 ( .C1(n6650), .C2(n6649), .A(n6657), .B(n6648), .ZN(n6652)
         );
  OAI211_X1 U8487 ( .C1(n6653), .C2(n6640), .A(n6652), .B(n6651), .ZN(n6654)
         );
  OAI21_X1 U8488 ( .B1(n6655), .B2(n6640), .A(n6654), .ZN(n6656) );
  OAI211_X1 U8489 ( .C1(n6657), .C2(n6640), .A(n6656), .B(n7547), .ZN(n6661)
         );
  MUX2_X1 U8490 ( .A(n6659), .B(n6658), .S(n6640), .Z(n6660) );
  AOI21_X1 U8491 ( .B1(n6661), .B2(n6660), .A(n7834), .ZN(n6667) );
  INV_X1 U8492 ( .A(n6662), .ZN(n6665) );
  INV_X1 U8493 ( .A(n6663), .ZN(n6664) );
  MUX2_X1 U8494 ( .A(n6665), .B(n6664), .S(n6640), .Z(n6666) );
  OAI21_X1 U8495 ( .B1(n6667), .B2(n6666), .A(n6668), .ZN(n6678) );
  NAND2_X1 U8496 ( .A1(n8755), .A2(n6668), .ZN(n6670) );
  INV_X1 U8497 ( .A(n6673), .ZN(n6669) );
  AOI211_X1 U8498 ( .C1(n6640), .C2(n6670), .A(n6669), .B(n5131), .ZN(n6677)
         );
  INV_X1 U8499 ( .A(n8755), .ZN(n6674) );
  OAI211_X1 U8500 ( .C1(n6674), .C2(n6673), .A(n6679), .B(n6672), .ZN(n6675)
         );
  MUX2_X1 U8501 ( .A(n5132), .B(n6675), .S(n6640), .Z(n6676) );
  AOI21_X1 U8502 ( .B1(n6678), .B2(n6677), .A(n6676), .ZN(n6682) );
  INV_X1 U8503 ( .A(n6680), .ZN(n6681) );
  NOR2_X1 U8504 ( .A1(n8171), .A2(n6640), .ZN(n6686) );
  INV_X1 U8505 ( .A(n8171), .ZN(n8411) );
  NOR2_X1 U8506 ( .A1(n8411), .A2(n6742), .ZN(n6685) );
  MUX2_X1 U8507 ( .A(n6686), .B(n6685), .S(n8946), .Z(n6687) );
  INV_X1 U8508 ( .A(n8384), .ZN(n8410) );
  NOR2_X1 U8509 ( .A1(n8943), .A2(n8410), .ZN(n6690) );
  INV_X1 U8510 ( .A(n6688), .ZN(n6689) );
  MUX2_X1 U8511 ( .A(n6690), .B(n6689), .S(n6640), .Z(n6691) );
  OAI21_X1 U8512 ( .B1(n6692), .B2(n6691), .A(n8721), .ZN(n6693) );
  INV_X1 U8513 ( .A(n6700), .ZN(n6703) );
  INV_X1 U8514 ( .A(n6697), .ZN(n6705) );
  INV_X1 U8515 ( .A(n6698), .ZN(n6699) );
  OAI21_X1 U8516 ( .B1(n6701), .B2(n6700), .A(n6699), .ZN(n6702) );
  INV_X1 U8517 ( .A(n8661), .ZN(n8643) );
  INV_X1 U8518 ( .A(n6704), .ZN(n6713) );
  OAI211_X1 U8519 ( .C1(n6706), .C2(n5165), .A(n6722), .B(n6715), .ZN(n6711)
         );
  NOR2_X1 U8520 ( .A1(n8823), .A2(n8346), .ZN(n6716) );
  NOR3_X1 U8521 ( .A1(n6707), .A2(n6716), .A3(n6640), .ZN(n6710) );
  INV_X1 U8522 ( .A(n6721), .ZN(n6708) );
  MUX2_X1 U8523 ( .A(n6708), .B(n6707), .S(n6640), .Z(n6709) );
  AOI21_X1 U8524 ( .B1(n8553), .B2(n6712), .A(n6640), .ZN(n6725) );
  AOI21_X1 U8525 ( .B1(n4750), .B2(n8645), .A(n6713), .ZN(n6720) );
  NAND2_X1 U8526 ( .A1(n6715), .A2(n6714), .ZN(n6719) );
  INV_X1 U8527 ( .A(n6716), .ZN(n6717) );
  OAI211_X1 U8528 ( .C1(n6720), .C2(n6719), .A(n6718), .B(n6717), .ZN(n6723)
         );
  NAND4_X1 U8529 ( .A1(n6723), .A2(n6722), .A3(n6721), .A4(n6640), .ZN(n6724)
         );
  INV_X1 U8530 ( .A(n6726), .ZN(n6729) );
  OAI21_X1 U8531 ( .B1(n6729), .B2(n6727), .A(n6640), .ZN(n6731) );
  INV_X1 U8532 ( .A(n8553), .ZN(n6728) );
  MUX2_X1 U8533 ( .A(n6729), .B(n6728), .S(n6640), .Z(n6730) );
  INV_X1 U8534 ( .A(n8537), .ZN(n6734) );
  NAND2_X1 U8535 ( .A1(n8521), .A2(n6732), .ZN(n6733) );
  MUX2_X1 U8536 ( .A(n6734), .B(n6733), .S(n6640), .Z(n6735) );
  MUX2_X1 U8537 ( .A(n6737), .B(n6736), .S(n6640), .Z(n6738) );
  MUX2_X1 U8538 ( .A(n6740), .B(n6739), .S(n6640), .Z(n6741) );
  NAND2_X1 U8539 ( .A1(n8397), .A2(n6640), .ZN(n6745) );
  NAND2_X1 U8540 ( .A1(n6743), .A2(n6742), .ZN(n6744) );
  MUX2_X1 U8541 ( .A(n6745), .B(n6744), .S(n8149), .Z(n6746) );
  MUX2_X1 U8542 ( .A(n6749), .B(n4367), .S(n6640), .Z(n6750) );
  INV_X1 U8543 ( .A(n6757), .ZN(n6758) );
  INV_X1 U8544 ( .A(P2_B_REG_SCAN_IN), .ZN(n9917) );
  INV_X1 U8545 ( .A(n6932), .ZN(n6762) );
  NOR4_X1 U8546 ( .A1(n10303), .A2(n8971), .A3(n6762), .A4(n8383), .ZN(n6763)
         );
  AOI211_X1 U8547 ( .C1(n6764), .C2(n8099), .A(n9917), .B(n6763), .ZN(n6765)
         );
  INV_X1 U8548 ( .A(n6766), .ZN(n6768) );
  NAND2_X1 U8549 ( .A1(n6770), .A2(n10245), .ZN(n6771) );
  NAND2_X1 U8550 ( .A1(n6771), .A2(n5211), .ZN(P1_U3520) );
  INV_X1 U8551 ( .A(n10283), .ZN(n6772) );
  NAND2_X1 U8552 ( .A1(n6772), .A2(n7748), .ZN(n7315) );
  AND2_X4 U8553 ( .A1(n4419), .A2(n6773), .ZN(n6884) );
  NAND2_X1 U8554 ( .A1(n7886), .A2(n6793), .ZN(n6774) );
  AND2_X1 U8555 ( .A1(n7315), .A2(n6774), .ZN(n7194) );
  OR2_X1 U8556 ( .A1(n6304), .A2(n7313), .ZN(n6776) );
  XNOR2_X1 U8557 ( .A(n6775), .B(n6776), .ZN(n7195) );
  INV_X1 U8558 ( .A(n6775), .ZN(n8091) );
  NAND2_X1 U8559 ( .A1(n6776), .A2(n8091), .ZN(n6777) );
  OR2_X1 U8560 ( .A1(n6778), .A2(n7313), .ZN(n6781) );
  XNOR2_X1 U8561 ( .A(n6884), .B(n8090), .ZN(n6779) );
  XNOR2_X1 U8562 ( .A(n6781), .B(n6779), .ZN(n8092) );
  INV_X1 U8563 ( .A(n6779), .ZN(n6780) );
  NAND2_X1 U8564 ( .A1(n6781), .A2(n6780), .ZN(n6782) );
  NOR2_X1 U8565 ( .A1(n6783), .A2(n7313), .ZN(n6784) );
  XNOR2_X1 U8566 ( .A(n6884), .B(n10272), .ZN(n8315) );
  NAND2_X1 U8567 ( .A1(n6784), .A2(n8315), .ZN(n6788) );
  INV_X1 U8568 ( .A(n6784), .ZN(n6786) );
  INV_X1 U8569 ( .A(n8315), .ZN(n6785) );
  NAND2_X1 U8570 ( .A1(n6786), .A2(n6785), .ZN(n6787) );
  NAND2_X1 U8571 ( .A1(n8420), .A2(n7748), .ZN(n6791) );
  XNOR2_X1 U8572 ( .A(n7569), .B(n6793), .ZN(n6790) );
  XNOR2_X1 U8573 ( .A(n6791), .B(n6790), .ZN(n8313) );
  AND2_X1 U8574 ( .A1(n6788), .A2(n8313), .ZN(n6789) );
  INV_X1 U8575 ( .A(n6790), .ZN(n8278) );
  NAND2_X1 U8576 ( .A1(n6791), .A2(n8278), .ZN(n6792) );
  NAND2_X1 U8577 ( .A1(n8307), .A2(n6792), .ZN(n6794) );
  XNOR2_X1 U8578 ( .A(n7802), .B(n6793), .ZN(n6795) );
  NAND2_X1 U8579 ( .A1(n8419), .A2(n7748), .ZN(n6796) );
  XNOR2_X1 U8580 ( .A(n6795), .B(n6796), .ZN(n8279) );
  INV_X1 U8581 ( .A(n6795), .ZN(n8077) );
  NAND2_X1 U8582 ( .A1(n8077), .A2(n6796), .ZN(n6797) );
  NAND2_X1 U8583 ( .A1(n8272), .A2(n6797), .ZN(n6798) );
  XNOR2_X1 U8584 ( .A(n7750), .B(n6884), .ZN(n6799) );
  OR2_X1 U8585 ( .A1(n7580), .A2(n7313), .ZN(n6800) );
  XNOR2_X1 U8586 ( .A(n6799), .B(n6800), .ZN(n8076) );
  INV_X1 U8587 ( .A(n6799), .ZN(n6801) );
  NAND2_X1 U8588 ( .A1(n6801), .A2(n6800), .ZN(n6802) );
  XNOR2_X1 U8589 ( .A(n7828), .B(n6884), .ZN(n6803) );
  NOR2_X1 U8590 ( .A1(n8206), .A2(n7313), .ZN(n6804) );
  NAND2_X1 U8591 ( .A1(n6803), .A2(n6804), .ZN(n6808) );
  INV_X1 U8592 ( .A(n6803), .ZN(n8205) );
  INV_X1 U8593 ( .A(n6804), .ZN(n6805) );
  NAND2_X1 U8594 ( .A1(n8205), .A2(n6805), .ZN(n6806) );
  NAND2_X1 U8595 ( .A1(n6808), .A2(n6806), .ZN(n7643) );
  XNOR2_X1 U8596 ( .A(n10337), .B(n6884), .ZN(n6809) );
  NOR2_X1 U8597 ( .A1(n7893), .A2(n7313), .ZN(n6810) );
  NAND2_X1 U8598 ( .A1(n6809), .A2(n6810), .ZN(n6813) );
  INV_X1 U8599 ( .A(n6809), .ZN(n7657) );
  INV_X1 U8600 ( .A(n6810), .ZN(n6811) );
  NAND2_X1 U8601 ( .A1(n7657), .A2(n6811), .ZN(n6812) );
  XNOR2_X1 U8602 ( .A(n8891), .B(n6793), .ZN(n6817) );
  NOR2_X1 U8603 ( .A1(n7927), .A2(n7313), .ZN(n6815) );
  XNOR2_X1 U8604 ( .A(n6817), .B(n6815), .ZN(n7668) );
  AND2_X1 U8605 ( .A1(n7668), .A2(n6813), .ZN(n6814) );
  NAND2_X1 U8606 ( .A1(n7656), .A2(n6814), .ZN(n7660) );
  INV_X1 U8607 ( .A(n6815), .ZN(n6816) );
  NAND2_X1 U8608 ( .A1(n6817), .A2(n6816), .ZN(n6818) );
  XNOR2_X1 U8609 ( .A(n8887), .B(n6884), .ZN(n6819) );
  NOR2_X1 U8610 ( .A1(n7973), .A2(n7313), .ZN(n6820) );
  NAND2_X1 U8611 ( .A1(n6819), .A2(n6820), .ZN(n6823) );
  INV_X1 U8612 ( .A(n6819), .ZN(n7970) );
  INV_X1 U8613 ( .A(n6820), .ZN(n6821) );
  NAND2_X1 U8614 ( .A1(n7970), .A2(n6821), .ZN(n6822) );
  NAND2_X1 U8615 ( .A1(n6823), .A2(n6822), .ZN(n7849) );
  XNOR2_X1 U8616 ( .A(n8751), .B(n6884), .ZN(n6829) );
  NOR2_X1 U8617 ( .A1(n8232), .A2(n7313), .ZN(n6824) );
  NAND2_X1 U8618 ( .A1(n6829), .A2(n6824), .ZN(n8167) );
  INV_X1 U8619 ( .A(n6829), .ZN(n8231) );
  INV_X1 U8620 ( .A(n6824), .ZN(n6827) );
  NAND2_X1 U8621 ( .A1(n8231), .A2(n6827), .ZN(n6825) );
  XNOR2_X1 U8622 ( .A(n8946), .B(n6793), .ZN(n8172) );
  OR2_X1 U8623 ( .A1(n8171), .A2(n7313), .ZN(n6831) );
  AND2_X1 U8624 ( .A1(n8172), .A2(n6831), .ZN(n6835) );
  INV_X1 U8625 ( .A(n6835), .ZN(n8170) );
  XNOR2_X1 U8626 ( .A(n8243), .B(n6884), .ZN(n8166) );
  INV_X1 U8627 ( .A(n8166), .ZN(n6826) );
  OR2_X1 U8628 ( .A1(n7997), .A2(n7313), .ZN(n8165) );
  NAND2_X1 U8629 ( .A1(n6826), .A2(n8165), .ZN(n8168) );
  NAND2_X1 U8630 ( .A1(n8167), .A2(n8165), .ZN(n6830) );
  NOR2_X1 U8631 ( .A1(n8165), .A2(n6827), .ZN(n6828) );
  AOI22_X1 U8632 ( .A1(n8166), .A2(n6830), .B1(n6829), .B2(n6828), .ZN(n6834)
         );
  XNOR2_X1 U8633 ( .A(n8739), .B(n6793), .ZN(n6840) );
  NOR2_X1 U8634 ( .A1(n8384), .A2(n7313), .ZN(n6838) );
  XNOR2_X1 U8635 ( .A(n6840), .B(n6838), .ZN(n8180) );
  INV_X1 U8636 ( .A(n8172), .ZN(n6833) );
  INV_X1 U8637 ( .A(n6831), .ZN(n6832) );
  NAND2_X1 U8638 ( .A1(n6833), .A2(n6832), .ZN(n8169) );
  OAI211_X1 U8639 ( .C1(n6835), .C2(n6834), .A(n8180), .B(n8169), .ZN(n6836)
         );
  INV_X1 U8640 ( .A(n6836), .ZN(n6837) );
  INV_X1 U8641 ( .A(n6838), .ZN(n6839) );
  NAND2_X1 U8642 ( .A1(n6840), .A2(n6839), .ZN(n6841) );
  XNOR2_X1 U8643 ( .A(n8933), .B(n6884), .ZN(n8263) );
  NOR2_X1 U8644 ( .A1(n8386), .A2(n7313), .ZN(n6842) );
  NOR2_X1 U8645 ( .A1(n8117), .A2(n7313), .ZN(n8259) );
  OAI22_X1 U8646 ( .A1(n8263), .A2(n6842), .B1(n8259), .B2(n8258), .ZN(n6846)
         );
  INV_X1 U8647 ( .A(n6842), .ZN(n8262) );
  AND2_X1 U8648 ( .A1(n6842), .A2(n8259), .ZN(n6843) );
  XNOR2_X1 U8649 ( .A(n8930), .B(n6884), .ZN(n6847) );
  NOR2_X1 U8650 ( .A1(n8358), .A2(n7313), .ZN(n6848) );
  NAND2_X1 U8651 ( .A1(n6847), .A2(n6848), .ZN(n6851) );
  INV_X1 U8652 ( .A(n6847), .ZN(n8354) );
  INV_X1 U8653 ( .A(n6848), .ZN(n6849) );
  NAND2_X1 U8654 ( .A1(n8354), .A2(n6849), .ZN(n6850) );
  AND2_X1 U8655 ( .A1(n6851), .A2(n6850), .ZN(n8287) );
  XNOR2_X1 U8656 ( .A(n8926), .B(n6793), .ZN(n6852) );
  NOR2_X1 U8657 ( .A1(n8288), .A2(n7313), .ZN(n6853) );
  INV_X1 U8658 ( .A(n6852), .ZN(n6854) );
  NAND2_X1 U8659 ( .A1(n6854), .A2(n6853), .ZN(n6855) );
  XNOR2_X1 U8660 ( .A(n8834), .B(n6793), .ZN(n6857) );
  NAND2_X1 U8661 ( .A1(n8406), .A2(n7748), .ZN(n6858) );
  NAND2_X1 U8662 ( .A1(n6857), .A2(n6858), .ZN(n6856) );
  INV_X1 U8663 ( .A(n6857), .ZN(n8195) );
  INV_X1 U8664 ( .A(n6858), .ZN(n6859) );
  NAND2_X1 U8665 ( .A1(n8195), .A2(n6859), .ZN(n8191) );
  XNOR2_X1 U8666 ( .A(n8634), .B(n6884), .ZN(n6860) );
  NOR2_X1 U8667 ( .A1(n8223), .A2(n7313), .ZN(n6861) );
  NAND2_X1 U8668 ( .A1(n6860), .A2(n6861), .ZN(n8217) );
  INV_X1 U8669 ( .A(n6860), .ZN(n8216) );
  INV_X1 U8670 ( .A(n6861), .ZN(n6862) );
  NAND2_X1 U8671 ( .A1(n8216), .A2(n6862), .ZN(n6863) );
  XNOR2_X1 U8672 ( .A(n8823), .B(n6793), .ZN(n6867) );
  INV_X1 U8673 ( .A(n6867), .ZN(n6864) );
  NOR2_X1 U8674 ( .A1(n8346), .A2(n7313), .ZN(n6866) );
  NAND2_X1 U8675 ( .A1(n6864), .A2(n6866), .ZN(n6865) );
  AND2_X1 U8676 ( .A1(n8217), .A2(n6865), .ZN(n6869) );
  INV_X1 U8677 ( .A(n6865), .ZN(n6868) );
  XNOR2_X1 U8678 ( .A(n6867), .B(n6866), .ZN(n8218) );
  XNOR2_X1 U8679 ( .A(n8604), .B(n6793), .ZN(n6870) );
  NAND2_X1 U8680 ( .A1(n8403), .A2(n7748), .ZN(n8341) );
  INV_X1 U8681 ( .A(n6870), .ZN(n6871) );
  NOR2_X1 U8682 ( .A1(n6872), .A2(n6871), .ZN(n6873) );
  XNOR2_X1 U8683 ( .A(n8813), .B(n6884), .ZN(n6876) );
  XNOR2_X1 U8684 ( .A(n8575), .B(n6884), .ZN(n6879) );
  NAND2_X1 U8685 ( .A1(n8402), .A2(n7748), .ZN(n8181) );
  AOI21_X1 U8686 ( .B1(n8297), .B2(n8299), .A(n8181), .ZN(n6875) );
  NAND2_X1 U8687 ( .A1(n8182), .A2(n6875), .ZN(n6883) );
  AND2_X1 U8688 ( .A1(n6877), .A2(n6876), .ZN(n8296) );
  OR2_X1 U8689 ( .A1(n8299), .A2(n7313), .ZN(n8300) );
  NAND2_X1 U8690 ( .A1(n8297), .A2(n8300), .ZN(n6881) );
  INV_X1 U8691 ( .A(n8300), .ZN(n6878) );
  AND2_X1 U8692 ( .A1(n6879), .A2(n6878), .ZN(n6880) );
  AOI21_X1 U8693 ( .B1(n8296), .B2(n6881), .A(n6880), .ZN(n6882) );
  NAND2_X1 U8694 ( .A1(n6883), .A2(n6882), .ZN(n8251) );
  XNOR2_X1 U8695 ( .A(n8802), .B(n6884), .ZN(n6885) );
  NOR2_X1 U8696 ( .A1(n8368), .A2(n7313), .ZN(n6886) );
  AND2_X1 U8697 ( .A1(n6885), .A2(n6886), .ZN(n8248) );
  OR2_X2 U8698 ( .A1(n8251), .A2(n8248), .ZN(n6888) );
  INV_X1 U8699 ( .A(n6885), .ZN(n8249) );
  INV_X1 U8700 ( .A(n6886), .ZN(n6887) );
  NAND2_X1 U8701 ( .A1(n8249), .A2(n6887), .ZN(n8247) );
  XNOR2_X1 U8702 ( .A(n8543), .B(n6793), .ZN(n6889) );
  NAND2_X1 U8703 ( .A1(n8399), .A2(n7748), .ZN(n6890) );
  XNOR2_X1 U8704 ( .A(n6889), .B(n6890), .ZN(n8366) );
  INV_X1 U8705 ( .A(n6889), .ZN(n6892) );
  INV_X1 U8706 ( .A(n6890), .ZN(n6891) );
  NAND2_X1 U8707 ( .A1(n6892), .A2(n6891), .ZN(n6893) );
  XNOR2_X1 U8708 ( .A(n8793), .B(n6793), .ZN(n6894) );
  NOR2_X1 U8709 ( .A1(n8367), .A2(n7313), .ZN(n6895) );
  XNOR2_X1 U8710 ( .A(n6894), .B(n6895), .ZN(n8157) );
  INV_X1 U8711 ( .A(n6894), .ZN(n6896) );
  NAND2_X1 U8712 ( .A1(n8397), .A2(n7748), .ZN(n6897) );
  XNOR2_X1 U8713 ( .A(n6897), .B(n6793), .ZN(n6921) );
  NOR4_X1 U8714 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6901) );
  NOR4_X1 U8715 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6900) );
  NOR4_X1 U8716 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6899) );
  NOR4_X1 U8717 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n6898) );
  NAND4_X1 U8718 ( .A1(n6901), .A2(n6900), .A3(n6899), .A4(n6898), .ZN(n6910)
         );
  NOR2_X1 U8719 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .ZN(
        n6905) );
  NOR4_X1 U8720 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n6904) );
  NOR4_X1 U8721 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n6903) );
  NOR4_X1 U8722 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n6902) );
  NAND4_X1 U8723 ( .A1(n6905), .A2(n6904), .A3(n6903), .A4(n6902), .ZN(n6909)
         );
  INV_X1 U8724 ( .A(n8978), .ZN(n6908) );
  XNOR2_X1 U8725 ( .A(n7925), .B(P2_B_REG_SCAN_IN), .ZN(n6906) );
  NAND2_X1 U8726 ( .A1(n8023), .A2(n6906), .ZN(n6907) );
  OAI21_X1 U8727 ( .B1(n6910), .B2(n6909), .A(n10302), .ZN(n7331) );
  INV_X1 U8728 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10310) );
  NAND2_X1 U8729 ( .A1(n10302), .A2(n10310), .ZN(n6912) );
  AND2_X1 U8730 ( .A1(n8978), .A2(n8023), .ZN(n10311) );
  INV_X1 U8731 ( .A(n10311), .ZN(n6911) );
  NAND2_X1 U8732 ( .A1(n6912), .A2(n6911), .ZN(n7327) );
  INV_X1 U8733 ( .A(n7327), .ZN(n6913) );
  AND2_X1 U8734 ( .A1(n7331), .A2(n6913), .ZN(n7717) );
  AND2_X1 U8735 ( .A1(n7925), .A2(n8978), .ZN(n10308) );
  INV_X1 U8736 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10307) );
  NAND2_X1 U8737 ( .A1(n7717), .A2(n7715), .ZN(n6931) );
  OR2_X1 U8738 ( .A1(n6915), .A2(n7719), .ZN(n7726) );
  INV_X1 U8739 ( .A(n7726), .ZN(n6916) );
  NAND2_X1 U8740 ( .A1(n6930), .A2(n6916), .ZN(n6918) );
  OR2_X2 U8741 ( .A1(n6917), .A2(n6915), .ZN(n10328) );
  NOR3_X1 U8742 ( .A1(n6587), .A2(n6921), .A3(n8392), .ZN(n6919) );
  AOI21_X1 U8743 ( .B1(n6587), .B2(n6921), .A(n6919), .ZN(n6927) );
  NAND3_X1 U8744 ( .A1(n8149), .A2(n8364), .A3(n6921), .ZN(n6920) );
  OAI21_X1 U8745 ( .B1(n8149), .B2(n6921), .A(n6920), .ZN(n6922) );
  NAND2_X1 U8746 ( .A1(n8149), .A2(n8392), .ZN(n6924) );
  AND2_X1 U8747 ( .A1(n10326), .A2(n7341), .ZN(n6923) );
  NAND2_X1 U8748 ( .A1(n6924), .A2(n8377), .ZN(n6925) );
  OAI211_X1 U8749 ( .C1(n6928), .C2(n6927), .A(n6926), .B(n6925), .ZN(n6941)
         );
  INV_X1 U8750 ( .A(n8969), .ZN(n6929) );
  OAI22_X1 U8751 ( .A1(n8367), .A2(n8383), .B1(n7467), .B2(n8385), .ZN(n8143)
         );
  INV_X1 U8752 ( .A(n8143), .ZN(n6938) );
  NAND2_X1 U8753 ( .A1(n6931), .A2(n7328), .ZN(n6936) );
  OR2_X1 U8754 ( .A1(n6932), .A2(n7341), .ZN(n7713) );
  AND3_X1 U8755 ( .A1(n6934), .A2(n6933), .A3(n7713), .ZN(n6935) );
  NAND2_X1 U8756 ( .A1(n6936), .A2(n6935), .ZN(n7312) );
  AOI22_X1 U8757 ( .A1(n8510), .A2(n8372), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n6937) );
  OAI21_X1 U8758 ( .B1(n6938), .B2(n8374), .A(n6937), .ZN(n6939) );
  NAND2_X1 U8759 ( .A1(n6941), .A2(n6940), .ZN(P2_U3222) );
  INV_X1 U8760 ( .A(n7755), .ZN(n6942) );
  NAND2_X1 U8761 ( .A1(n6944), .A2(n7755), .ZN(n6945) );
  NAND2_X1 U8762 ( .A1(n6996), .A2(n6945), .ZN(n7015) );
  OAI21_X1 U8763 ( .B1(n7015), .B2(n6946), .A(P1_STATE_REG_SCAN_IN), .ZN(
        P1_U3083) );
  NAND2_X1 U8764 ( .A1(n6950), .A2(P2_U3152), .ZN(n7308) );
  AND2_X1 U8765 ( .A1(n4271), .A2(P2_U3152), .ZN(n7350) );
  INV_X2 U8766 ( .A(n7350), .ZN(n8974) );
  OAI222_X1 U8767 ( .A1(n7172), .A2(P2_U3152), .B1(n7308), .B2(n6957), .C1(
        n6948), .C2(n8974), .ZN(P2_U3356) );
  OAI222_X1 U8768 ( .A1(n7161), .A2(P2_U3152), .B1(n7308), .B2(n6955), .C1(
        n6949), .C2(n8974), .ZN(P2_U3357) );
  AND2_X1 U8769 ( .A1(n6950), .A2(P1_U3084), .ZN(n7149) );
  NOR2_X1 U8770 ( .A1(n6950), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10089) );
  INV_X2 U8771 ( .A(n10089), .ZN(n10087) );
  OAI222_X1 U8772 ( .A1(n10094), .A2(n4927), .B1(n10087), .B2(n6962), .C1(
        P1_U3084), .C2(n7031), .ZN(P1_U3350) );
  INV_X1 U8773 ( .A(n6951), .ZN(n6952) );
  OAI222_X1 U8774 ( .A1(n8974), .A2(n5322), .B1(n7308), .B2(n6952), .C1(
        P2_U3152), .C2(n7225), .ZN(P2_U3354) );
  OAI222_X1 U8775 ( .A1(n10094), .A2(n6953), .B1(n10087), .B2(n6952), .C1(
        P1_U3084), .C2(n7181), .ZN(P1_U3349) );
  INV_X2 U8776 ( .A(n7149), .ZN(n10094) );
  OAI222_X1 U8777 ( .A1(n7067), .A2(P1_U3084), .B1(n10087), .B2(n6955), .C1(
        n6954), .C2(n10094), .ZN(P1_U3352) );
  OAI222_X1 U8778 ( .A1(n7123), .A2(P1_U3084), .B1(n10087), .B2(n6957), .C1(
        n6956), .C2(n10094), .ZN(P1_U3351) );
  INV_X1 U8779 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6959) );
  INV_X1 U8780 ( .A(n6958), .ZN(n6963) );
  INV_X1 U8781 ( .A(n7054), .ZN(n7033) );
  OAI222_X1 U8782 ( .A1(n10094), .A2(n6959), .B1(n10087), .B2(n6963), .C1(
        P1_U3084), .C2(n7033), .ZN(P1_U3348) );
  INV_X1 U8783 ( .A(n6960), .ZN(n6971) );
  AOI22_X1 U8784 ( .A1(n10125), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n7149), .ZN(n6961) );
  OAI21_X1 U8785 ( .B1(n6971), .B2(n10087), .A(n6961), .ZN(P1_U3345) );
  INV_X1 U8786 ( .A(n7308), .ZN(n8960) );
  OAI222_X1 U8787 ( .A1(n8974), .A2(n4930), .B1(n8977), .B2(n6962), .C1(
        P2_U3152), .C2(n7211), .ZN(P2_U3355) );
  INV_X1 U8788 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6964) );
  OAI222_X1 U8789 ( .A1(n8974), .A2(n6964), .B1(n8977), .B2(n6963), .C1(
        P2_U3152), .C2(n7262), .ZN(P2_U3353) );
  INV_X1 U8790 ( .A(n6965), .ZN(n6967) );
  INV_X1 U8791 ( .A(n6966), .ZN(n7236) );
  OAI222_X1 U8792 ( .A1(n8974), .A2(n5361), .B1(n7308), .B2(n6967), .C1(
        P2_U3152), .C2(n7236), .ZN(P2_U3352) );
  INV_X1 U8793 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6968) );
  INV_X1 U8794 ( .A(n7040), .ZN(n7111) );
  OAI222_X1 U8795 ( .A1(n10094), .A2(n6968), .B1(n10087), .B2(n6967), .C1(
        P1_U3084), .C2(n7111), .ZN(P1_U3347) );
  INV_X1 U8796 ( .A(n6969), .ZN(n6977) );
  AOI22_X1 U8797 ( .A1(n7266), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n7149), .ZN(n6970) );
  OAI21_X1 U8798 ( .B1(n6977), .B2(n10087), .A(n6970), .ZN(P1_U3344) );
  OAI222_X1 U8799 ( .A1(n8974), .A2(n6972), .B1(n8977), .B2(n6971), .C1(
        P2_U3152), .C2(n7287), .ZN(P2_U3350) );
  INV_X1 U8800 ( .A(n6973), .ZN(n6974) );
  OAI222_X1 U8801 ( .A1(n8974), .A2(n4779), .B1(n7308), .B2(n6974), .C1(
        P2_U3152), .C2(n7249), .ZN(P2_U3351) );
  INV_X1 U8802 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6975) );
  INV_X1 U8803 ( .A(n7096), .ZN(n7091) );
  OAI222_X1 U8804 ( .A1(n10094), .A2(n6975), .B1(n10087), .B2(n6974), .C1(
        P1_U3084), .C2(n7091), .ZN(P1_U3346) );
  INV_X1 U8805 ( .A(n6976), .ZN(n7495) );
  OAI222_X1 U8806 ( .A1(n8974), .A2(n6978), .B1(n8977), .B2(n6977), .C1(n7495), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U8807 ( .A(n6979), .ZN(n6981) );
  INV_X1 U8808 ( .A(n7357), .ZN(n7362) );
  OAI222_X1 U8809 ( .A1(n10094), .A2(n6980), .B1(n10087), .B2(n6981), .C1(
        n7362), .C2(P1_U3084), .ZN(P1_U3343) );
  OAI222_X1 U8810 ( .A1(n8974), .A2(n6982), .B1(n7308), .B2(n6981), .C1(n7674), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U8811 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6986) );
  INV_X1 U8812 ( .A(n6984), .ZN(n6985) );
  AOI22_X1 U8813 ( .A1(n10218), .A2(n6986), .B1(n9278), .B2(n6985), .ZN(
        P1_U3441) );
  NAND2_X1 U8814 ( .A1(n8104), .A2(P2_U3966), .ZN(n6987) );
  OAI21_X1 U8815 ( .B1(P2_U3966), .B2(n10076), .A(n6987), .ZN(P2_U3583) );
  INV_X1 U8816 ( .A(n6988), .ZN(n6991) );
  INV_X1 U8817 ( .A(n7614), .ZN(n7612) );
  OAI222_X1 U8818 ( .A1(n10094), .A2(n6989), .B1(n10087), .B2(n6991), .C1(
        n7612), .C2(P1_U3084), .ZN(P1_U3342) );
  INV_X1 U8819 ( .A(n6990), .ZN(n7813) );
  OAI222_X1 U8820 ( .A1(n8974), .A2(n9834), .B1(n7308), .B2(n6991), .C1(n7813), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  INV_X1 U8821 ( .A(n6992), .ZN(n6995) );
  AOI22_X1 U8822 ( .A1(n9467), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n7149), .ZN(n6993) );
  OAI21_X1 U8823 ( .B1(n6995), .B2(n10087), .A(n6993), .ZN(P1_U3341) );
  INV_X1 U8824 ( .A(n6994), .ZN(n8031) );
  OAI222_X1 U8825 ( .A1(n8974), .A2(n9844), .B1(n7308), .B2(n6995), .C1(
        P2_U3152), .C2(n8031), .ZN(P2_U3346) );
  NOR2_X1 U8826 ( .A1(n10258), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8827 ( .A(n6996), .ZN(n6997) );
  INV_X1 U8828 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7008) );
  OR2_X1 U8829 ( .A1(n5815), .A2(n9280), .ZN(n7145) );
  INV_X1 U8830 ( .A(n7145), .ZN(n7001) );
  INV_X1 U8831 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n7005) );
  NAND2_X1 U8832 ( .A1(n6998), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7000) );
  OAI21_X1 U8833 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n7014), .A(n9279), .ZN(
        n7142) );
  INV_X1 U8834 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7143) );
  XNOR2_X1 U8835 ( .A(n7142), .B(n7143), .ZN(n6999) );
  AOI211_X1 U8836 ( .C1(n7001), .C2(n7005), .A(n7000), .B(n6999), .ZN(n7002)
         );
  INV_X1 U8837 ( .A(n7015), .ZN(n7004) );
  AOI22_X1 U8838 ( .A1(n7002), .A2(n7004), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3084), .ZN(n7007) );
  NOR2_X1 U8839 ( .A1(n7145), .A2(P1_U3084), .ZN(n7003) );
  NAND2_X1 U8840 ( .A1(n7004), .A2(n7003), .ZN(n10132) );
  NAND3_X1 U8841 ( .A1(n10190), .A2(P1_IR_REG_0__SCAN_IN), .A3(n7005), .ZN(
        n7006) );
  OAI211_X1 U8842 ( .C1(n10195), .C2(n7008), .A(n7007), .B(n7006), .ZN(
        P1_U3241) );
  INV_X1 U8843 ( .A(n7009), .ZN(n7012) );
  INV_X1 U8844 ( .A(n9471), .ZN(n10148) );
  OAI222_X1 U8845 ( .A1(n10094), .A2(n7010), .B1(n10087), .B2(n7012), .C1(
        n10148), .C2(P1_U3084), .ZN(P1_U3340) );
  INV_X1 U8846 ( .A(n7011), .ZN(n8434) );
  OAI222_X1 U8847 ( .A1(n8974), .A2(n7013), .B1(n7308), .B2(n7012), .C1(n8434), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8848 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n7029) );
  OR2_X1 U8849 ( .A1(n7014), .A2(P1_U3084), .ZN(n10091) );
  NOR2_X1 U8850 ( .A1(n7015), .A2(n10091), .ZN(n9516) );
  INV_X1 U8851 ( .A(n7031), .ZN(n7038) );
  NOR2_X1 U8852 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5294), .ZN(n7375) );
  INV_X1 U8853 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n7016) );
  MUX2_X1 U8854 ( .A(n7016), .B(P1_REG1_REG_1__SCAN_IN), .S(n7067), .Z(n7068)
         );
  AND2_X1 U8855 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n7069) );
  NAND2_X1 U8856 ( .A1(n7068), .A2(n7069), .ZN(n7125) );
  OR2_X1 U8857 ( .A1(n7067), .A2(n7016), .ZN(n7124) );
  INV_X1 U8858 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n7017) );
  MUX2_X1 U8859 ( .A(n7017), .B(P1_REG1_REG_2__SCAN_IN), .S(n7123), .Z(n7018)
         );
  INV_X1 U8860 ( .A(n7123), .ZN(n7136) );
  NAND2_X1 U8861 ( .A1(n7136), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7019) );
  INV_X1 U8862 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9962) );
  AND3_X1 U8863 ( .A1(n7020), .A2(n7128), .A3(n7019), .ZN(n7021) );
  NOR3_X1 U8864 ( .A1(n10132), .A2(n7037), .A3(n7021), .ZN(n7022) );
  AOI211_X1 U8865 ( .C1(n10188), .C2(n7038), .A(n7375), .B(n7022), .ZN(n7028)
         );
  XNOR2_X1 U8866 ( .A(n7031), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n7026) );
  INV_X1 U8867 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7024) );
  MUX2_X1 U8868 ( .A(n7024), .B(P1_REG2_REG_2__SCAN_IN), .S(n7123), .Z(n7132)
         );
  INV_X1 U8869 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7023) );
  XNOR2_X1 U8870 ( .A(n7067), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n7066) );
  AND2_X1 U8871 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n7140) );
  NAND2_X1 U8872 ( .A1(n7066), .A2(n7140), .ZN(n7065) );
  OAI21_X1 U8873 ( .B1(n7023), .B2(n7067), .A(n7065), .ZN(n7131) );
  NAND2_X1 U8874 ( .A1(n7132), .A2(n7131), .ZN(n7130) );
  OAI21_X1 U8875 ( .B1(n7123), .B2(n7024), .A(n7130), .ZN(n7025) );
  NAND2_X1 U8876 ( .A1(n9516), .A2(n9279), .ZN(n10182) );
  NAND2_X1 U8877 ( .A1(n7025), .A2(n7026), .ZN(n7030) );
  OAI211_X1 U8878 ( .C1(n7026), .C2(n7025), .A(n10143), .B(n7030), .ZN(n7027)
         );
  OAI211_X1 U8879 ( .C1(n7029), .C2(n10195), .A(n7028), .B(n7027), .ZN(
        P1_U3244) );
  XNOR2_X1 U8880 ( .A(n7096), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n7036) );
  INV_X1 U8881 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7034) );
  INV_X1 U8882 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7032) );
  INV_X1 U8883 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7447) );
  XNOR2_X1 U8884 ( .A(n7181), .B(n7447), .ZN(n7177) );
  XOR2_X1 U8885 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n7054), .Z(n7056) );
  OAI21_X1 U8886 ( .B1(n7033), .B2(n7032), .A(n7055), .ZN(n7114) );
  XOR2_X1 U8887 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n7040), .Z(n7115) );
  NAND2_X1 U8888 ( .A1(n7114), .A2(n7115), .ZN(n7113) );
  AOI21_X1 U8889 ( .B1(n7036), .B2(n7035), .A(n7090), .ZN(n7049) );
  INV_X1 U8890 ( .A(n7181), .ZN(n7039) );
  INV_X1 U8891 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10247) );
  MUX2_X1 U8892 ( .A(n10247), .B(P1_REG1_REG_4__SCAN_IN), .S(n7181), .Z(n7179)
         );
  NAND2_X1 U8893 ( .A1(n7180), .A2(n7179), .ZN(n7178) );
  OAI21_X1 U8894 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n7039), .A(n7178), .ZN(
        n7052) );
  INV_X1 U8895 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7515) );
  MUX2_X1 U8896 ( .A(n7515), .B(P1_REG1_REG_5__SCAN_IN), .S(n7054), .Z(n7051)
         );
  NOR2_X1 U8897 ( .A1(n7052), .A2(n7051), .ZN(n7050) );
  INV_X1 U8898 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10249) );
  MUX2_X1 U8899 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10249), .S(n7040), .Z(n7105)
         );
  NOR2_X1 U8900 ( .A1(n7040), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7041) );
  INV_X1 U8901 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7703) );
  MUX2_X1 U8902 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n7703), .S(n7096), .Z(n7042)
         );
  INV_X1 U8903 ( .A(n7095), .ZN(n7044) );
  NOR3_X1 U8904 ( .A1(n7106), .A2(n7042), .A3(n7041), .ZN(n7043) );
  OAI21_X1 U8905 ( .B1(n7044), .B2(n7043), .A(n10190), .ZN(n7048) );
  AND2_X1 U8906 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7638) );
  INV_X1 U8907 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n7045) );
  NOR2_X1 U8908 ( .A1(n10195), .A2(n7045), .ZN(n7046) );
  AOI211_X1 U8909 ( .C1(n10188), .C2(n7096), .A(n7638), .B(n7046), .ZN(n7047)
         );
  OAI211_X1 U8910 ( .C1(n7049), .C2(n10182), .A(n7048), .B(n7047), .ZN(
        P1_U3248) );
  INV_X1 U8911 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n7059) );
  NOR2_X1 U8912 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5333), .ZN(n7411) );
  AOI211_X1 U8913 ( .C1(n7052), .C2(n7051), .A(n10132), .B(n7050), .ZN(n7053)
         );
  AOI211_X1 U8914 ( .C1(n10188), .C2(n7054), .A(n7411), .B(n7053), .ZN(n7058)
         );
  OAI211_X1 U8915 ( .C1(n7056), .C2(n4422), .A(n10143), .B(n7055), .ZN(n7057)
         );
  OAI211_X1 U8916 ( .C1(n7059), .C2(n10195), .A(n7058), .B(n7057), .ZN(
        P1_U3246) );
  INV_X1 U8917 ( .A(n7060), .ZN(n7063) );
  INV_X1 U8918 ( .A(n9472), .ZN(n9496) );
  OAI222_X1 U8919 ( .A1(n10094), .A2(n7061), .B1(n10087), .B2(n7063), .C1(
        n9496), .C2(P1_U3084), .ZN(P1_U3339) );
  INV_X1 U8920 ( .A(n7062), .ZN(n8448) );
  OAI222_X1 U8921 ( .A1(n8974), .A2(n7064), .B1(n7308), .B2(n7063), .C1(n8448), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8922 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7075) );
  OAI211_X1 U8923 ( .C1(n7066), .C2(n7140), .A(n10143), .B(n7065), .ZN(n7074)
         );
  INV_X1 U8924 ( .A(n7067), .ZN(n7072) );
  INV_X1 U8925 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7452) );
  OAI211_X1 U8926 ( .C1(n7069), .C2(n7068), .A(n10190), .B(n7125), .ZN(n7070)
         );
  OAI21_X1 U8927 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n7452), .A(n7070), .ZN(n7071) );
  AOI21_X1 U8928 ( .B1(n10188), .B2(n7072), .A(n7071), .ZN(n7073) );
  OAI211_X1 U8929 ( .C1(n7075), .C2(n10195), .A(n7074), .B(n7073), .ZN(
        P1_U3242) );
  NAND2_X1 U8930 ( .A1(n5786), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n7078) );
  NAND2_X1 U8931 ( .A1(n4283), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n7077) );
  NAND2_X1 U8932 ( .A1(n5336), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n7076) );
  AND3_X1 U8933 ( .A1(n7078), .A2(n7077), .A3(n7076), .ZN(n9252) );
  INV_X1 U8934 ( .A(n9252), .ZN(n9523) );
  NAND2_X1 U8935 ( .A1(n9523), .A2(n9461), .ZN(n7079) );
  OAI21_X1 U8936 ( .B1(n9461), .B2(n8964), .A(n7079), .ZN(P1_U3586) );
  INV_X1 U8937 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n7081) );
  NAND2_X1 U8938 ( .A1(n7323), .A2(n9461), .ZN(n7080) );
  OAI21_X1 U8939 ( .B1(n9461), .B2(n7081), .A(n7080), .ZN(P1_U3555) );
  OR2_X1 U8940 ( .A1(n7082), .A2(n7458), .ZN(n9399) );
  INV_X1 U8941 ( .A(n9399), .ZN(n7085) );
  INV_X1 U8942 ( .A(n7083), .ZN(n7299) );
  OAI211_X1 U8943 ( .C1(n7085), .C2(n7299), .A(n7084), .B(n7523), .ZN(n7086)
         );
  OAI21_X1 U8944 ( .B1(n7087), .B2(n9770), .A(n7086), .ZN(n7459) );
  AOI21_X1 U8945 ( .B1(n7458), .B2(n7088), .A(n7459), .ZN(n7152) );
  INV_X1 U8946 ( .A(n10254), .ZN(n10251) );
  NAND2_X1 U8947 ( .A1(n10251), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7089) );
  OAI21_X1 U8948 ( .B1(n7152), .B2(n10251), .A(n7089), .ZN(P1_U3523) );
  INV_X1 U8949 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7092) );
  MUX2_X1 U8950 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n7092), .S(n10125), .Z(n10130) );
  XNOR2_X1 U8951 ( .A(n7266), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n7093) );
  AOI211_X1 U8952 ( .C1(n7094), .C2(n7093), .A(n10182), .B(n4412), .ZN(n7103)
         );
  INV_X1 U8953 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10390) );
  INV_X1 U8954 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10252) );
  MUX2_X1 U8955 ( .A(n10252), .B(P1_REG1_REG_8__SCAN_IN), .S(n10125), .Z(
        n10133) );
  NOR2_X1 U8956 ( .A1(n7266), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7263) );
  AOI21_X1 U8957 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n7266), .A(n7263), .ZN(
        n7097) );
  NAND2_X1 U8958 ( .A1(n10125), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7098) );
  AOI21_X1 U8959 ( .B1(n10135), .B2(n7098), .A(n7097), .ZN(n7099) );
  OAI21_X1 U8960 ( .B1(n4417), .B2(n7099), .A(n10190), .ZN(n7101) );
  AND2_X1 U8961 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7782) );
  AOI21_X1 U8962 ( .B1(n10188), .B2(n7266), .A(n7782), .ZN(n7100) );
  OAI211_X1 U8963 ( .C1(n10390), .C2(n10195), .A(n7101), .B(n7100), .ZN(n7102)
         );
  OR2_X1 U8964 ( .A1(n7103), .A2(n7102), .ZN(P1_U3250) );
  INV_X1 U8965 ( .A(n7104), .ZN(n7108) );
  INV_X1 U8966 ( .A(n7105), .ZN(n7107) );
  AOI21_X1 U8967 ( .B1(n7108), .B2(n7107), .A(n7106), .ZN(n7118) );
  INV_X1 U8968 ( .A(n10195), .ZN(n10126) );
  INV_X1 U8969 ( .A(n10188), .ZN(n10149) );
  NOR2_X1 U8970 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7109), .ZN(n9124) );
  INV_X1 U8971 ( .A(n9124), .ZN(n7110) );
  OAI21_X1 U8972 ( .B1(n10149), .B2(n7111), .A(n7110), .ZN(n7112) );
  AOI21_X1 U8973 ( .B1(n10126), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n7112), .ZN(
        n7117) );
  OAI211_X1 U8974 ( .C1(n7115), .C2(n7114), .A(n10143), .B(n7113), .ZN(n7116)
         );
  OAI211_X1 U8975 ( .C1(n7118), .C2(n10132), .A(n7117), .B(n7116), .ZN(
        P1_U3247) );
  INV_X1 U8976 ( .A(n7119), .ZN(n7121) );
  INV_X1 U8977 ( .A(n10163), .ZN(n9500) );
  OAI222_X1 U8978 ( .A1(n10094), .A2(n7120), .B1(n10087), .B2(n7121), .C1(
        P1_U3084), .C2(n9500), .ZN(P1_U3338) );
  OAI222_X1 U8979 ( .A1(n8974), .A2(n7122), .B1(n7308), .B2(n7121), .C1(
        P2_U3152), .C2(n8456), .ZN(P2_U3343) );
  INV_X1 U8980 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7147) );
  MUX2_X1 U8981 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n7017), .S(n7123), .Z(n7126)
         );
  NAND3_X1 U8982 ( .A1(n7126), .A2(n7125), .A3(n7124), .ZN(n7127) );
  NAND2_X1 U8983 ( .A1(n7128), .A2(n7127), .ZN(n7129) );
  INV_X1 U8984 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7431) );
  OAI22_X1 U8985 ( .A1(n10132), .A2(n7129), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7431), .ZN(n7135) );
  OAI211_X1 U8986 ( .C1(n7132), .C2(n7131), .A(n10143), .B(n7130), .ZN(n7133)
         );
  INV_X1 U8987 ( .A(n7133), .ZN(n7134) );
  AOI211_X1 U8988 ( .C1(n10188), .C2(n7136), .A(n7135), .B(n7134), .ZN(n7146)
         );
  OAI21_X1 U8989 ( .B1(n7139), .B2(n7138), .A(n7137), .ZN(n7293) );
  AND3_X1 U8990 ( .A1(n9279), .A2(n9280), .A3(n7140), .ZN(n7141) );
  AOI21_X1 U8991 ( .B1(n7143), .B2(n7142), .A(n7141), .ZN(n7144) );
  OAI211_X1 U8992 ( .C1(n7293), .C2(n7145), .A(n9461), .B(n7144), .ZN(n7187)
         );
  OAI211_X1 U8993 ( .C1(n7147), .C2(n10195), .A(n7146), .B(n7187), .ZN(
        P1_U3243) );
  INV_X1 U8994 ( .A(n7148), .ZN(n7189) );
  AOI22_X1 U8995 ( .A1(n10175), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n7149), .ZN(n7150) );
  OAI21_X1 U8996 ( .B1(n7189), .B2(n10087), .A(n7150), .ZN(P1_U3337) );
  INV_X1 U8997 ( .A(n10245), .ZN(n10243) );
  NAND2_X1 U8998 ( .A1(n10243), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n7151) );
  OAI21_X1 U8999 ( .B1(n7152), .B2(n10243), .A(n7151), .ZN(P1_U3454) );
  AOI211_X1 U9000 ( .C1(n7155), .C2(n7154), .A(n7153), .B(n10259), .ZN(n7163)
         );
  AOI22_X1 U9001 ( .A1(n10258), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n7160) );
  INV_X1 U9002 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10346) );
  MUX2_X1 U9003 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6297), .S(n7161), .Z(n7156)
         );
  OAI21_X1 U9004 ( .B1(n10346), .B2(n4442), .A(n7156), .ZN(n7157) );
  NAND3_X1 U9005 ( .A1(n10255), .A2(n7158), .A3(n7157), .ZN(n7159) );
  OAI211_X1 U9006 ( .C1(n10260), .C2(n7161), .A(n7160), .B(n7159), .ZN(n7162)
         );
  OR2_X1 U9007 ( .A1(n7163), .A2(n7162), .ZN(P2_U3246) );
  AOI211_X1 U9008 ( .C1(n7166), .C2(n7165), .A(n7164), .B(n10259), .ZN(n7174)
         );
  AOI22_X1 U9009 ( .A1(n10258), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n7171) );
  MUX2_X1 U9010 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6196), .S(n7172), .Z(n7167)
         );
  INV_X1 U9011 ( .A(n7167), .ZN(n7169) );
  OAI211_X1 U9012 ( .C1(n7169), .C2(n7168), .A(n10255), .B(n7205), .ZN(n7170)
         );
  OAI211_X1 U9013 ( .C1(n10260), .C2(n7172), .A(n7171), .B(n7170), .ZN(n7173)
         );
  OR2_X1 U9014 ( .A1(n7174), .A2(n7173), .ZN(P2_U3247) );
  AOI21_X1 U9015 ( .B1(n7177), .B2(n7176), .A(n7175), .ZN(n7185) );
  OAI21_X1 U9016 ( .B1(n7180), .B2(n7179), .A(n7178), .ZN(n7183) );
  AND2_X1 U9017 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9070) );
  NOR2_X1 U9018 ( .A1(n10149), .A2(n7181), .ZN(n7182) );
  AOI211_X1 U9019 ( .C1(n10190), .C2(n7183), .A(n9070), .B(n7182), .ZN(n7184)
         );
  OAI21_X1 U9020 ( .B1(n7185), .B2(n10182), .A(n7184), .ZN(n7186) );
  AOI21_X1 U9021 ( .B1(n10126), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n7186), .ZN(
        n7188) );
  NAND2_X1 U9022 ( .A1(n7188), .A2(n7187), .ZN(P1_U3245) );
  OAI222_X1 U9023 ( .A1(n8974), .A2(n7190), .B1(n7308), .B2(n7189), .C1(n8469), 
        .C2(P2_U3152), .ZN(P2_U3342) );
  NOR2_X1 U9024 ( .A1(n7312), .A2(P2_U3152), .ZN(n8088) );
  INV_X1 U9025 ( .A(n8088), .ZN(n7193) );
  OR2_X1 U9026 ( .A1(n6778), .A2(n8385), .ZN(n7192) );
  OR2_X1 U9027 ( .A1(n7314), .A2(n8383), .ZN(n7191) );
  NAND2_X1 U9028 ( .A1(n7192), .A2(n7191), .ZN(n10294) );
  AOI22_X1 U9029 ( .A1(n7193), .A2(P2_REG3_REG_1__SCAN_IN), .B1(n8387), .B2(
        n10294), .ZN(n7198) );
  OAI21_X1 U9030 ( .B1(n7195), .B2(n7194), .A(n8094), .ZN(n7196) );
  NAND2_X1 U9031 ( .A1(n8380), .A2(n7196), .ZN(n7197) );
  OAI211_X1 U9032 ( .C1(n10320), .C2(n8364), .A(n7198), .B(n7197), .ZN(
        P2_U3224) );
  AOI211_X1 U9033 ( .C1(n7201), .C2(n7200), .A(n7199), .B(n10259), .ZN(n7202)
         );
  INV_X1 U9034 ( .A(n7202), .ZN(n7210) );
  NOR2_X1 U9035 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6334), .ZN(n7208) );
  AND3_X1 U9036 ( .A1(n7205), .A2(n7204), .A3(n7203), .ZN(n7206) );
  NOR3_X1 U9037 ( .A1(n10261), .A2(n7218), .A3(n7206), .ZN(n7207) );
  AOI211_X1 U9038 ( .C1(P2_ADDR_REG_3__SCAN_IN), .C2(n10258), .A(n7208), .B(
        n7207), .ZN(n7209) );
  OAI211_X1 U9039 ( .C1(n10260), .C2(n7211), .A(n7210), .B(n7209), .ZN(
        P2_U3248) );
  AOI211_X1 U9040 ( .C1(n7214), .C2(n7213), .A(n7212), .B(n10259), .ZN(n7215)
         );
  INV_X1 U9041 ( .A(n7215), .ZN(n7224) );
  AND2_X1 U9042 ( .A1(P2_U3152), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7222) );
  INV_X1 U9043 ( .A(n7256), .ZN(n7220) );
  NOR3_X1 U9044 ( .A1(n7218), .A2(n7217), .A3(n7216), .ZN(n7219) );
  NOR3_X1 U9045 ( .A1(n10261), .A2(n7220), .A3(n7219), .ZN(n7221) );
  AOI211_X1 U9046 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n10258), .A(n7222), .B(
        n7221), .ZN(n7223) );
  OAI211_X1 U9047 ( .C1(n10260), .C2(n7225), .A(n7224), .B(n7223), .ZN(
        P2_U3249) );
  AOI211_X1 U9048 ( .C1(n7227), .C2(n7226), .A(n10259), .B(n4415), .ZN(n7228)
         );
  INV_X1 U9049 ( .A(n7228), .ZN(n7235) );
  AND2_X1 U9050 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n8074) );
  INV_X1 U9051 ( .A(n7243), .ZN(n7232) );
  NOR3_X1 U9052 ( .A1(n7258), .A2(n7230), .A3(n7229), .ZN(n7231) );
  NOR3_X1 U9053 ( .A1(n10261), .A2(n7232), .A3(n7231), .ZN(n7233) );
  AOI211_X1 U9054 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n10258), .A(n8074), .B(
        n7233), .ZN(n7234) );
  OAI211_X1 U9055 ( .C1(n10260), .C2(n7236), .A(n7235), .B(n7234), .ZN(
        P2_U3251) );
  AOI211_X1 U9056 ( .C1(n7239), .C2(n7238), .A(n10259), .B(n7237), .ZN(n7240)
         );
  INV_X1 U9057 ( .A(n7240), .ZN(n7248) );
  NOR2_X1 U9058 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9937), .ZN(n7246) );
  AND3_X1 U9059 ( .A1(n7243), .A2(n7242), .A3(n7241), .ZN(n7244) );
  NOR3_X1 U9060 ( .A1(n7284), .A2(n10261), .A3(n7244), .ZN(n7245) );
  AOI211_X1 U9061 ( .C1(P2_ADDR_REG_7__SCAN_IN), .C2(n10258), .A(n7246), .B(
        n7245), .ZN(n7247) );
  OAI211_X1 U9062 ( .C1(n10260), .C2(n7249), .A(n7248), .B(n7247), .ZN(
        P2_U3252) );
  AOI211_X1 U9063 ( .C1(n7252), .C2(n7251), .A(n10259), .B(n7250), .ZN(n7253)
         );
  INV_X1 U9064 ( .A(n7253), .ZN(n7261) );
  AND2_X1 U9065 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8274) );
  AND3_X1 U9066 ( .A1(n7256), .A2(n7255), .A3(n7254), .ZN(n7257) );
  NOR3_X1 U9067 ( .A1(n10261), .A2(n7258), .A3(n7257), .ZN(n7259) );
  AOI211_X1 U9068 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n10258), .A(n8274), .B(
        n7259), .ZN(n7260) );
  OAI211_X1 U9069 ( .C1(n10260), .C2(n7262), .A(n7261), .B(n7260), .ZN(
        P2_U3250) );
  XNOR2_X1 U9070 ( .A(n7357), .B(P1_REG1_REG_10__SCAN_IN), .ZN(n7264) );
  AOI21_X1 U9071 ( .B1(n7265), .B2(n7264), .A(n7361), .ZN(n7273) );
  XNOR2_X1 U9072 ( .A(n7357), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n7267) );
  AOI211_X1 U9073 ( .C1(n7268), .C2(n7267), .A(n10182), .B(n7356), .ZN(n7269)
         );
  INV_X1 U9074 ( .A(n7269), .ZN(n7272) );
  NAND2_X1 U9075 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7708) );
  OAI21_X1 U9076 ( .B1(n10149), .B2(n7362), .A(n7708), .ZN(n7270) );
  AOI21_X1 U9077 ( .B1(n10126), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n7270), .ZN(
        n7271) );
  OAI211_X1 U9078 ( .C1(n7273), .C2(n10132), .A(n7272), .B(n7271), .ZN(
        P1_U3251) );
  AOI211_X1 U9079 ( .C1(n7276), .C2(n7275), .A(n10259), .B(n7274), .ZN(n7289)
         );
  NAND2_X1 U9080 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n8213) );
  INV_X1 U9081 ( .A(n8213), .ZN(n7277) );
  AOI21_X1 U9082 ( .B1(n10258), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n7277), .ZN(
        n7286) );
  INV_X1 U9083 ( .A(n7278), .ZN(n7281) );
  MUX2_X1 U9084 ( .A(n10350), .B(P2_REG1_REG_8__SCAN_IN), .S(n7279), .Z(n7280)
         );
  NAND2_X1 U9085 ( .A1(n7281), .A2(n7280), .ZN(n7283) );
  OAI211_X1 U9086 ( .C1(n7284), .C2(n7283), .A(n7282), .B(n10255), .ZN(n7285)
         );
  OAI211_X1 U9087 ( .C1(n10260), .C2(n7287), .A(n7286), .B(n7285), .ZN(n7288)
         );
  OR2_X1 U9088 ( .A1(n7289), .A2(n7288), .ZN(P2_U3253) );
  INV_X1 U9089 ( .A(n9148), .ZN(n9125) );
  AOI22_X1 U9090 ( .A1(n9125), .A2(n7290), .B1(n7458), .B2(n9138), .ZN(n7295)
         );
  OAI21_X1 U9091 ( .B1(n7292), .B2(n10201), .A(n7291), .ZN(n9103) );
  AOI22_X1 U9092 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n9103), .B1(n7293), .B2(
        n9145), .ZN(n7294) );
  NAND2_X1 U9093 ( .A1(n7295), .A2(n7294), .ZN(P1_U3230) );
  INV_X1 U9094 ( .A(n7296), .ZN(n7420) );
  AOI211_X1 U9095 ( .C1(n7458), .C2(n5858), .A(n10239), .B(n7420), .ZN(n7455)
         );
  NAND2_X1 U9096 ( .A1(n7297), .A2(n9398), .ZN(n7300) );
  XOR2_X1 U9097 ( .A(n7298), .B(n7300), .Z(n7305) );
  AOI22_X1 U9098 ( .A1(n7323), .A2(n9794), .B1(n9796), .B2(n9460), .ZN(n7304)
         );
  INV_X1 U9099 ( .A(n9398), .ZN(n7302) );
  AOI21_X1 U9100 ( .B1(n7300), .B2(n7299), .A(n9767), .ZN(n7301) );
  OAI21_X1 U9101 ( .B1(n7302), .B2(n9401), .A(n7301), .ZN(n7303) );
  OAI211_X1 U9102 ( .C1(n7305), .C2(n9753), .A(n7304), .B(n7303), .ZN(n7453)
         );
  AOI211_X1 U9103 ( .C1(n5858), .C2(n10047), .A(n7455), .B(n7453), .ZN(n7353)
         );
  NAND2_X1 U9104 ( .A1(n10251), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7306) );
  OAI21_X1 U9105 ( .B1(n7353), .B2(n10251), .A(n7306), .ZN(P1_U3524) );
  INV_X1 U9106 ( .A(n7307), .ZN(n7309) );
  OAI222_X1 U9107 ( .A1(n8974), .A2(n9928), .B1(n7308), .B2(n7309), .C1(n8483), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  INV_X1 U9108 ( .A(n10187), .ZN(n9488) );
  OAI222_X1 U9109 ( .A1(n10094), .A2(n7310), .B1(n10087), .B2(n7309), .C1(
        n9488), .C2(P1_U3084), .ZN(P1_U3336) );
  INV_X1 U9110 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7885) );
  NOR2_X1 U9111 ( .A1(n7885), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10257) );
  OR2_X1 U9112 ( .A1(n6304), .A2(n8385), .ZN(n7883) );
  NOR2_X1 U9113 ( .A1(n8374), .A2(n7883), .ZN(n7311) );
  AOI211_X1 U9114 ( .C1(P2_REG3_REG_0__SCAN_IN), .C2(n7312), .A(n10257), .B(
        n7311), .ZN(n7318) );
  OAI22_X1 U9115 ( .A1(n8353), .A2(n7314), .B1(n7886), .B2(n8377), .ZN(n7316)
         );
  NAND2_X1 U9116 ( .A1(n7316), .A2(n7315), .ZN(n7317) );
  OAI211_X1 U9117 ( .C1(n8364), .C2(n7886), .A(n7318), .B(n7317), .ZN(P2_U3234) );
  XNOR2_X1 U9118 ( .A(n7320), .B(n7319), .ZN(n7322) );
  XNOR2_X1 U9119 ( .A(n7321), .B(n7322), .ZN(n7326) );
  AOI22_X1 U9120 ( .A1(n9103), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n9138), .B2(
        n5858), .ZN(n7325) );
  AOI22_X1 U9121 ( .A1(n9125), .A2(n9460), .B1(n9150), .B2(n7323), .ZN(n7324)
         );
  OAI211_X1 U9122 ( .C1(n7326), .C2(n9140), .A(n7325), .B(n7324), .ZN(P1_U3220) );
  NAND3_X1 U9123 ( .A1(n7328), .A2(n7327), .A3(n7713), .ZN(n7329) );
  NOR2_X1 U9124 ( .A1(n10303), .A2(n7329), .ZN(n7330) );
  INV_X1 U9125 ( .A(n7715), .ZN(n7332) );
  INV_X1 U9126 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n7348) );
  OR2_X2 U9127 ( .A1(n7334), .A2(n7333), .ZN(n10290) );
  XNOR2_X1 U9128 ( .A(n7335), .B(n7339), .ZN(n7337) );
  INV_X1 U9129 ( .A(n8385), .ZN(n8360) );
  AOI22_X1 U9130 ( .A1(n8324), .A2(n6310), .B1(n8421), .B2(n8360), .ZN(n8086)
         );
  INV_X1 U9131 ( .A(n8086), .ZN(n7336) );
  AOI21_X1 U9132 ( .B1(n10290), .B2(n7337), .A(n7336), .ZN(n8067) );
  NAND2_X1 U9133 ( .A1(n7338), .A2(n10283), .ZN(n7537) );
  NAND2_X1 U9134 ( .A1(n6304), .A2(n10320), .ZN(n7536) );
  NAND2_X1 U9135 ( .A1(n7537), .A2(n7536), .ZN(n7340) );
  NAND2_X1 U9136 ( .A1(n7340), .A2(n7339), .ZN(n7595) );
  OAI21_X1 U9137 ( .B1(n7340), .B2(n7339), .A(n7595), .ZN(n8062) );
  MUX2_X1 U9138 ( .A(n6615), .B(n7341), .S(n7719), .Z(n7343) );
  AND2_X1 U9139 ( .A1(n6915), .A2(n7723), .ZN(n7342) );
  NAND2_X1 U9140 ( .A1(n7343), .A2(n7342), .ZN(n7933) );
  NAND3_X1 U9141 ( .A1(n8099), .A2(n7344), .A3(n7719), .ZN(n10342) );
  XNOR2_X1 U9142 ( .A(n10277), .B(n8090), .ZN(n8063) );
  AOI21_X1 U9143 ( .B1(n8062), .B2(n10331), .A(n7345), .ZN(n7346) );
  NAND2_X1 U9144 ( .A1(n8067), .A2(n7346), .ZN(n7403) );
  NAND2_X1 U9145 ( .A1(n7403), .A2(n10345), .ZN(n7347) );
  OAI21_X1 U9146 ( .B1(n10345), .B2(n7348), .A(n7347), .ZN(P2_U3457) );
  INV_X1 U9147 ( .A(n7349), .ZN(n7381) );
  AOI22_X1 U9148 ( .A1(n7351), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n7350), .ZN(n7352) );
  OAI21_X1 U9149 ( .B1(n7381), .B2(n8977), .A(n7352), .ZN(P2_U3340) );
  INV_X1 U9150 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7355) );
  OR2_X1 U9151 ( .A1(n7353), .A2(n10243), .ZN(n7354) );
  OAI21_X1 U9152 ( .B1(n10245), .B2(n7355), .A(n7354), .ZN(P1_U3457) );
  INV_X1 U9153 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7358) );
  AOI22_X1 U9154 ( .A1(n7614), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7358), .B2(
        n7612), .ZN(n7359) );
  OAI21_X1 U9155 ( .B1(n7360), .B2(n7359), .A(n7615), .ZN(n7370) );
  INV_X1 U9156 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7368) );
  INV_X1 U9157 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9935) );
  AOI21_X1 U9158 ( .B1(n9935), .B2(n7362), .A(n7361), .ZN(n7364) );
  INV_X1 U9159 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7987) );
  AOI22_X1 U9160 ( .A1(n7614), .A2(n7987), .B1(P1_REG1_REG_11__SCAN_IN), .B2(
        n7612), .ZN(n7363) );
  AOI21_X1 U9161 ( .B1(n7364), .B2(n7363), .A(n7611), .ZN(n7365) );
  OR2_X1 U9162 ( .A1(n7365), .A2(n10132), .ZN(n7367) );
  AND2_X1 U9163 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7880) );
  AOI21_X1 U9164 ( .B1(n10188), .B2(n7614), .A(n7880), .ZN(n7366) );
  OAI211_X1 U9165 ( .C1(n7368), .C2(n10195), .A(n7367), .B(n7366), .ZN(n7369)
         );
  AOI21_X1 U9166 ( .B1(n7370), .B2(n10143), .A(n7369), .ZN(n7371) );
  INV_X1 U9167 ( .A(n7371), .ZN(P1_U3252) );
  OAI21_X1 U9168 ( .B1(n7374), .B2(n7373), .A(n7372), .ZN(n7379) );
  AOI22_X1 U9169 ( .A1(n9125), .A2(n9458), .B1(n9150), .B2(n9460), .ZN(n7377)
         );
  AOI21_X1 U9170 ( .B1(n9138), .B2(n7387), .A(n7375), .ZN(n7376) );
  OAI211_X1 U9171 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9146), .A(n7377), .B(
        n7376), .ZN(n7378) );
  AOI21_X1 U9172 ( .B1(n7379), .B2(n9145), .A(n7378), .ZN(n7380) );
  INV_X1 U9173 ( .A(n7380), .ZN(P1_U3216) );
  INV_X1 U9174 ( .A(n9511), .ZN(n9513) );
  OAI222_X1 U9175 ( .A1(n10094), .A2(n7382), .B1(n10087), .B2(n7381), .C1(
        P1_U3084), .C2(n9513), .ZN(P1_U3335) );
  NAND2_X1 U9176 ( .A1(n7424), .A2(n7383), .ZN(n7384) );
  NAND2_X1 U9177 ( .A1(n7384), .A2(n4727), .ZN(n7439) );
  OAI21_X1 U9178 ( .B1(n7384), .B2(n4727), .A(n7439), .ZN(n7487) );
  INV_X1 U9179 ( .A(n7487), .ZN(n7389) );
  XNOR2_X1 U9180 ( .A(n9365), .B(n9404), .ZN(n7385) );
  AOI222_X1 U9181 ( .A1(n9799), .A2(n7385), .B1(n9458), .B2(n9796), .C1(n9460), 
        .C2(n9794), .ZN(n7490) );
  OR2_X1 U9182 ( .A1(n7418), .A2(n7485), .ZN(n7386) );
  AOI22_X1 U9183 ( .A1(n4409), .A2(n10033), .B1(n7387), .B2(n10047), .ZN(n7388) );
  OAI211_X1 U9184 ( .C1(n9753), .C2(n7389), .A(n7490), .B(n7388), .ZN(n7391)
         );
  NAND2_X1 U9185 ( .A1(n7391), .A2(n10254), .ZN(n7390) );
  OAI21_X1 U9186 ( .B1(n10254), .B2(n9962), .A(n7390), .ZN(P1_U3526) );
  INV_X1 U9187 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7393) );
  NAND2_X1 U9188 ( .A1(n7391), .A2(n10245), .ZN(n7392) );
  OAI21_X1 U9189 ( .B1(n10245), .B2(n7393), .A(n7392), .ZN(P1_U3463) );
  INV_X1 U9190 ( .A(n8308), .ZN(n7394) );
  AOI211_X1 U9191 ( .C1(n7396), .C2(n7395), .A(n8377), .B(n7394), .ZN(n7401)
         );
  MUX2_X1 U9192 ( .A(n8372), .B(P2_U3152), .S(P2_REG3_REG_3__SCAN_IN), .Z(
        n7400) );
  NAND2_X1 U9193 ( .A1(n8420), .A2(n8360), .ZN(n7397) );
  OAI21_X1 U9194 ( .B1(n6778), .B2(n8383), .A(n7397), .ZN(n7601) );
  INV_X1 U9195 ( .A(n7601), .ZN(n7398) );
  OAI22_X1 U9196 ( .A1(n8364), .A2(n7652), .B1(n7398), .B2(n8374), .ZN(n7399)
         );
  OR3_X1 U9197 ( .A1(n7401), .A2(n7400), .A3(n7399), .ZN(P2_U3220) );
  NAND2_X1 U9198 ( .A1(n7403), .A2(n10352), .ZN(n7404) );
  OAI21_X1 U9199 ( .B1(n10352), .B2(n6196), .A(n7404), .ZN(P2_U3522) );
  XNOR2_X1 U9200 ( .A(n7406), .B(n7405), .ZN(n7407) );
  XNOR2_X1 U9201 ( .A(n7408), .B(n7407), .ZN(n7414) );
  AOI22_X1 U9202 ( .A1(n9125), .A2(n9456), .B1(n9150), .B2(n9458), .ZN(n7413)
         );
  INV_X1 U9203 ( .A(n9138), .ZN(n9153) );
  NOR2_X1 U9204 ( .A1(n9153), .A2(n7409), .ZN(n7410) );
  AOI211_X1 U9205 ( .C1(n10200), .C2(n9134), .A(n7411), .B(n7410), .ZN(n7412)
         );
  OAI211_X1 U9206 ( .C1(n7414), .C2(n9140), .A(n7413), .B(n7412), .ZN(P1_U3225) );
  INV_X1 U9207 ( .A(n7415), .ZN(n7416) );
  NAND2_X1 U9208 ( .A1(n7417), .A2(n7416), .ZN(n7530) );
  INV_X1 U9209 ( .A(n5893), .ZN(n7464) );
  INV_X1 U9210 ( .A(n7418), .ZN(n7419) );
  OAI21_X1 U9211 ( .B1(n10219), .B2(n7420), .A(n7419), .ZN(n10220) );
  INV_X1 U9212 ( .A(n7421), .ZN(n7422) );
  AOI21_X1 U9213 ( .B1(n7425), .B2(n7423), .A(n7422), .ZN(n7430) );
  AOI22_X1 U9214 ( .A1(n9794), .A2(n7290), .B1(n9459), .B2(n9796), .ZN(n7429)
         );
  OAI21_X1 U9215 ( .B1(n7426), .B2(n7425), .A(n7424), .ZN(n7427) );
  NAND2_X1 U9216 ( .A1(n7427), .A2(n10234), .ZN(n7428) );
  OAI211_X1 U9217 ( .C1(n7430), .C2(n9767), .A(n7429), .B(n7428), .ZN(n10221)
         );
  NAND2_X1 U9218 ( .A1(n10221), .A2(n10209), .ZN(n7434) );
  OAI22_X1 U9219 ( .A1(n9755), .A2(n7431), .B1(n7024), .B2(n10209), .ZN(n7432)
         );
  AOI21_X1 U9220 ( .B1(n9758), .B2(n9102), .A(n7432), .ZN(n7433) );
  OAI211_X1 U9221 ( .C1(n9762), .C2(n10220), .A(n7434), .B(n7433), .ZN(
        P1_U3289) );
  NAND2_X1 U9222 ( .A1(n7508), .A2(n7435), .ZN(n10225) );
  XNOR2_X1 U9223 ( .A(n7437), .B(n7436), .ZN(n7445) );
  INV_X1 U9224 ( .A(n7437), .ZN(n9403) );
  NAND3_X1 U9225 ( .A1(n7439), .A2(n9403), .A3(n7438), .ZN(n7440) );
  NAND2_X1 U9226 ( .A1(n7440), .A2(n7503), .ZN(n7443) );
  OAI22_X1 U9227 ( .A1(n7441), .A2(n9772), .B1(n7471), .B2(n9770), .ZN(n7442)
         );
  AOI21_X1 U9228 ( .B1(n7443), .B2(n10234), .A(n7442), .ZN(n7444) );
  OAI21_X1 U9229 ( .B1(n7445), .B2(n9767), .A(n7444), .ZN(n10226) );
  NAND2_X1 U9230 ( .A1(n10226), .A2(n10209), .ZN(n7450) );
  INV_X1 U9231 ( .A(n9072), .ZN(n7446) );
  OAI22_X1 U9232 ( .A1(n10209), .A2(n7447), .B1(n7446), .B2(n9755), .ZN(n7448)
         );
  AOI21_X1 U9233 ( .B1(n9758), .B2(n9071), .A(n7448), .ZN(n7449) );
  OAI211_X1 U9234 ( .C1(n9762), .C2(n10225), .A(n7450), .B(n7449), .ZN(
        P1_U3287) );
  INV_X1 U9235 ( .A(n7451), .ZN(n7463) );
  OAI222_X1 U9236 ( .A1(n8974), .A2(n9943), .B1(n8977), .B2(n7463), .C1(n7723), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  NOR2_X1 U9237 ( .A1(n9755), .A2(n7452), .ZN(n7454) );
  AOI211_X1 U9238 ( .C1(n7464), .C2(n7455), .A(n7454), .B(n7453), .ZN(n7457)
         );
  AOI22_X1 U9239 ( .A1(n9758), .A2(n5858), .B1(n10211), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n7456) );
  OAI21_X1 U9240 ( .B1(n7457), .B2(n10211), .A(n7456), .ZN(P1_U3290) );
  INV_X1 U9241 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7462) );
  OAI21_X1 U9242 ( .B1(n9802), .B2(n9758), .A(n7458), .ZN(n7461) );
  AOI22_X1 U9243 ( .A1(n7459), .A2(n10209), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n10201), .ZN(n7460) );
  OAI211_X1 U9244 ( .C1(n10209), .C2(n7462), .A(n7461), .B(n7460), .ZN(
        P1_U3291) );
  OAI222_X1 U9245 ( .A1(n7465), .A2(n10094), .B1(P1_U3084), .B2(n7464), .C1(
        n10087), .C2(n7463), .ZN(P1_U3334) );
  NAND2_X1 U9246 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n8422), .ZN(n7466) );
  OAI21_X1 U9247 ( .B1(n7467), .B2(n8422), .A(n7466), .ZN(P2_U3581) );
  INV_X1 U9248 ( .A(n9406), .ZN(n7506) );
  INV_X1 U9249 ( .A(n9161), .ZN(n9158) );
  AOI21_X1 U9250 ( .B1(n7468), .B2(n7506), .A(n9158), .ZN(n7469) );
  INV_X1 U9251 ( .A(n9407), .ZN(n9163) );
  XNOR2_X1 U9252 ( .A(n7469), .B(n9163), .ZN(n7470) );
  OAI222_X1 U9253 ( .A1(n9772), .A2(n7471), .B1(n9770), .B2(n7794), .C1(n7470), 
        .C2(n9767), .ZN(n10231) );
  INV_X1 U9254 ( .A(n10231), .ZN(n7482) );
  INV_X1 U9255 ( .A(n7472), .ZN(n7504) );
  INV_X1 U9256 ( .A(n7473), .ZN(n7474) );
  OAI21_X1 U9257 ( .B1(n7504), .B2(n7474), .A(n9163), .ZN(n7476) );
  NAND2_X1 U9258 ( .A1(n7476), .A2(n7475), .ZN(n10233) );
  NAND2_X1 U9259 ( .A1(n10209), .A2(n10234), .ZN(n9804) );
  INV_X1 U9260 ( .A(n9804), .ZN(n7488) );
  INV_X1 U9261 ( .A(n7477), .ZN(n7529) );
  OAI21_X1 U9262 ( .B1(n10229), .B2(n7511), .A(n7529), .ZN(n10230) );
  AOI22_X1 U9263 ( .A1(n10211), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n9126), .B2(
        n10201), .ZN(n7479) );
  NAND2_X1 U9264 ( .A1(n9758), .A2(n9123), .ZN(n7478) );
  OAI211_X1 U9265 ( .C1(n9762), .C2(n10230), .A(n7479), .B(n7478), .ZN(n7480)
         );
  AOI21_X1 U9266 ( .B1(n10233), .B2(n7488), .A(n7480), .ZN(n7481) );
  OAI21_X1 U9267 ( .B1(n7482), .B2(n10211), .A(n7481), .ZN(P1_U3285) );
  NAND2_X1 U9268 ( .A1(n9802), .A2(n4409), .ZN(n7484) );
  AOI22_X1 U9269 ( .A1(n10211), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10201), .B2(
        n5294), .ZN(n7483) );
  OAI211_X1 U9270 ( .C1(n7485), .C2(n9789), .A(n7484), .B(n7483), .ZN(n7486)
         );
  AOI21_X1 U9271 ( .B1(n7488), .B2(n7487), .A(n7486), .ZN(n7489) );
  OAI21_X1 U9272 ( .B1(n7490), .B2(n10211), .A(n7489), .ZN(P1_U3288) );
  XOR2_X1 U9273 ( .A(n7492), .B(n7491), .Z(n7500) );
  NAND2_X1 U9274 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7662) );
  INV_X1 U9275 ( .A(n7662), .ZN(n7493) );
  AOI21_X1 U9276 ( .B1(n10258), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7493), .ZN(
        n7494) );
  OAI21_X1 U9277 ( .B1(n7495), .B2(n10260), .A(n7494), .ZN(n7499) );
  AOI211_X1 U9278 ( .C1(n7497), .C2(n7496), .A(n10259), .B(n4418), .ZN(n7498)
         );
  AOI211_X1 U9279 ( .C1(n10255), .C2(n7500), .A(n7499), .B(n7498), .ZN(n7501)
         );
  INV_X1 U9280 ( .A(n7501), .ZN(P2_U3254) );
  NAND2_X1 U9281 ( .A1(n7503), .A2(n7502), .ZN(n7505) );
  AOI21_X1 U9282 ( .B1(n7506), .B2(n7505), .A(n7504), .ZN(n10207) );
  INV_X1 U9283 ( .A(n10207), .ZN(n7513) );
  XNOR2_X1 U9284 ( .A(n7468), .B(n7506), .ZN(n7507) );
  AOI222_X1 U9285 ( .A1(n9799), .A2(n7507), .B1(n9458), .B2(n9794), .C1(n9456), 
        .C2(n9796), .ZN(n10204) );
  NAND2_X1 U9286 ( .A1(n7508), .A2(n10198), .ZN(n7509) );
  NAND2_X1 U9287 ( .A1(n7509), .A2(n10033), .ZN(n7510) );
  NOR2_X1 U9288 ( .A1(n7511), .A2(n7510), .ZN(n10197) );
  AOI21_X1 U9289 ( .B1(n10198), .B2(n10047), .A(n10197), .ZN(n7512) );
  OAI211_X1 U9290 ( .C1(n9753), .C2(n7513), .A(n10204), .B(n7512), .ZN(n7516)
         );
  NAND2_X1 U9291 ( .A1(n7516), .A2(n10254), .ZN(n7514) );
  OAI21_X1 U9292 ( .B1(n10254), .B2(n7515), .A(n7514), .ZN(P1_U3528) );
  INV_X1 U9293 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9885) );
  NAND2_X1 U9294 ( .A1(n7516), .A2(n10245), .ZN(n7517) );
  OAI21_X1 U9295 ( .B1(n10245), .B2(n9885), .A(n7517), .ZN(P1_U3469) );
  INV_X1 U9296 ( .A(n7518), .ZN(n7535) );
  OAI222_X1 U9297 ( .A1(n9435), .A2(P1_U3084), .B1(n10087), .B2(n7535), .C1(
        n7519), .C2(n10094), .ZN(P1_U3333) );
  OAI21_X1 U9298 ( .B1(n9410), .B2(n7520), .A(n7683), .ZN(n7521) );
  AOI222_X1 U9299 ( .A1(n9799), .A2(n7521), .B1(n9456), .B2(n9794), .C1(n9454), 
        .C2(n9796), .ZN(n7700) );
  AND2_X1 U9300 ( .A1(n7523), .A2(n7522), .ZN(n10208) );
  INV_X1 U9301 ( .A(n9783), .ZN(n9738) );
  OAI21_X1 U9302 ( .B1(n7526), .B2(n7525), .A(n7524), .ZN(n7696) );
  INV_X1 U9303 ( .A(n7527), .ZN(n7528) );
  AOI211_X1 U9304 ( .C1(n7698), .C2(n7529), .A(n10239), .B(n7528), .ZN(n7697)
         );
  OR2_X1 U9305 ( .A1(n7530), .A2(n5893), .ZN(n9736) );
  INV_X1 U9306 ( .A(n9736), .ZN(n9780) );
  NAND2_X1 U9307 ( .A1(n7697), .A2(n9780), .ZN(n7532) );
  AOI22_X1 U9308 ( .A1(n10211), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7634), .B2(
        n10201), .ZN(n7531) );
  OAI211_X1 U9309 ( .C1(n7641), .C2(n9789), .A(n7532), .B(n7531), .ZN(n7533)
         );
  AOI21_X1 U9310 ( .B1(n9738), .B2(n7696), .A(n7533), .ZN(n7534) );
  OAI21_X1 U9311 ( .B1(n7700), .B2(n10211), .A(n7534), .ZN(P1_U3284) );
  OAI222_X1 U9312 ( .A1(n8974), .A2(n9938), .B1(P2_U3152), .B2(n7719), .C1(
        n8977), .C2(n7535), .ZN(P2_U3338) );
  NAND3_X1 U9313 ( .A1(n7537), .A2(n7536), .A3(n7594), .ZN(n7542) );
  INV_X1 U9314 ( .A(n7538), .ZN(n7539) );
  NAND2_X1 U9315 ( .A1(n6783), .A2(n7652), .ZN(n7543) );
  NAND2_X1 U9316 ( .A1(n6340), .A2(n7569), .ZN(n7544) );
  NAND2_X1 U9317 ( .A1(n7573), .A2(n7577), .ZN(n7572) );
  NAND2_X1 U9318 ( .A1(n8078), .A2(n7802), .ZN(n7545) );
  NAND2_X1 U9319 ( .A1(n7572), .A2(n7545), .ZN(n7742) );
  NAND2_X1 U9320 ( .A1(n7742), .A2(n7741), .ZN(n7744) );
  NAND2_X1 U9321 ( .A1(n10327), .A2(n7580), .ZN(n7546) );
  NAND2_X1 U9322 ( .A1(n7744), .A2(n7546), .ZN(n7548) );
  OAI21_X1 U9323 ( .B1(n7548), .B2(n7551), .A(n7830), .ZN(n7825) );
  NAND2_X1 U9324 ( .A1(n7604), .A2(n7652), .ZN(n7603) );
  OR2_X2 U9325 ( .A1(n7603), .A2(n8312), .ZN(n7574) );
  NOR2_X4 U9326 ( .A1(n7574), .A2(n8277), .ZN(n7745) );
  INV_X1 U9327 ( .A(n7747), .ZN(n7550) );
  INV_X1 U9328 ( .A(n7828), .ZN(n7823) );
  INV_X1 U9329 ( .A(n7843), .ZN(n7549) );
  AOI211_X1 U9330 ( .C1(n7828), .C2(n7550), .A(n10328), .B(n7549), .ZN(n7819)
         );
  XNOR2_X1 U9331 ( .A(n7552), .B(n7551), .ZN(n7554) );
  OR2_X1 U9332 ( .A1(n7893), .A2(n8385), .ZN(n7553) );
  OAI21_X1 U9333 ( .B1(n7580), .B2(n8383), .A(n7553), .ZN(n7645) );
  AOI21_X1 U9334 ( .B1(n7554), .B2(n10290), .A(n7645), .ZN(n7827) );
  INV_X1 U9335 ( .A(n7827), .ZN(n7555) );
  AOI211_X1 U9336 ( .C1(n10331), .C2(n7825), .A(n7819), .B(n7555), .ZN(n7589)
         );
  INV_X1 U9337 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7556) );
  OAI22_X1 U9338 ( .A1(n8956), .A2(n7823), .B1(n10345), .B2(n7556), .ZN(n7557)
         );
  INV_X1 U9339 ( .A(n7557), .ZN(n7558) );
  OAI21_X1 U9340 ( .B1(n7589), .B2(n4655), .A(n7558), .ZN(P2_U3472) );
  OAI21_X1 U9341 ( .B1(n7559), .B2(n7561), .A(n7560), .ZN(n7731) );
  AOI21_X1 U9342 ( .B1(n7603), .B2(n8312), .A(n10328), .ZN(n7562) );
  AND2_X1 U9343 ( .A1(n7562), .A2(n7574), .ZN(n7725) );
  XNOR2_X1 U9344 ( .A(n7564), .B(n7563), .ZN(n7566) );
  NAND2_X1 U9345 ( .A1(n8419), .A2(n8360), .ZN(n7565) );
  OAI21_X1 U9346 ( .B1(n6783), .B2(n8383), .A(n7565), .ZN(n8310) );
  AOI21_X1 U9347 ( .B1(n7566), .B2(n10290), .A(n8310), .ZN(n7733) );
  INV_X1 U9348 ( .A(n7733), .ZN(n7567) );
  AOI211_X1 U9349 ( .C1(n10331), .C2(n7731), .A(n7725), .B(n7567), .ZN(n7591)
         );
  INV_X1 U9350 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n7568) );
  OAI22_X1 U9351 ( .A1(n8956), .A2(n7569), .B1(n10345), .B2(n7568), .ZN(n7570)
         );
  INV_X1 U9352 ( .A(n7570), .ZN(n7571) );
  OAI21_X1 U9353 ( .B1(n7591), .B2(n4655), .A(n7571), .ZN(P2_U3463) );
  OAI21_X1 U9354 ( .B1(n7573), .B2(n7577), .A(n7572), .ZN(n7804) );
  AOI211_X1 U9355 ( .C1(n8277), .C2(n7574), .A(n10328), .B(n7745), .ZN(n7799)
         );
  NAND2_X1 U9356 ( .A1(n7576), .A2(n7575), .ZN(n7578) );
  XNOR2_X1 U9357 ( .A(n7578), .B(n7577), .ZN(n7581) );
  NAND2_X1 U9358 ( .A1(n8420), .A2(n8324), .ZN(n7579) );
  OAI21_X1 U9359 ( .B1(n7580), .B2(n8385), .A(n7579), .ZN(n8275) );
  AOI21_X1 U9360 ( .B1(n7581), .B2(n10290), .A(n8275), .ZN(n7806) );
  INV_X1 U9361 ( .A(n7806), .ZN(n7582) );
  AOI211_X1 U9362 ( .C1(n10331), .C2(n7804), .A(n7799), .B(n7582), .ZN(n7593)
         );
  INV_X1 U9363 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7583) );
  OAI22_X1 U9364 ( .A1(n8956), .A2(n7802), .B1(n10345), .B2(n7583), .ZN(n7584)
         );
  INV_X1 U9365 ( .A(n7584), .ZN(n7585) );
  OAI21_X1 U9366 ( .B1(n7593), .B2(n4655), .A(n7585), .ZN(P2_U3466) );
  INV_X1 U9367 ( .A(n7586), .ZN(n7608) );
  OAI222_X1 U9368 ( .A1(n9432), .A2(P1_U3084), .B1(n10087), .B2(n7608), .C1(
        n7587), .C2(n10094), .ZN(P1_U3332) );
  AOI22_X1 U9369 ( .A1(n8873), .A2(n7828), .B1(n4653), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n7588) );
  OAI21_X1 U9370 ( .B1(n7589), .B2(n4653), .A(n7588), .ZN(P2_U3527) );
  AOI22_X1 U9371 ( .A1(n8873), .A2(n8312), .B1(n4653), .B2(
        P2_REG1_REG_4__SCAN_IN), .ZN(n7590) );
  OAI21_X1 U9372 ( .B1(n7591), .B2(n4653), .A(n7590), .ZN(P2_U3524) );
  AOI22_X1 U9373 ( .A1(n8873), .A2(n8277), .B1(n4653), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n7592) );
  OAI21_X1 U9374 ( .B1(n7593), .B2(n4653), .A(n7592), .ZN(P2_U3525) );
  NAND3_X1 U9375 ( .A1(n7595), .A2(n7599), .A3(n7594), .ZN(n7596) );
  AND2_X1 U9376 ( .A1(n7597), .A2(n7596), .ZN(n10269) );
  XNOR2_X1 U9377 ( .A(n7599), .B(n7598), .ZN(n7602) );
  NOR2_X1 U9378 ( .A1(n10269), .A2(n7933), .ZN(n7600) );
  AOI211_X1 U9379 ( .C1(n7602), .C2(n10290), .A(n7601), .B(n7600), .ZN(n10275)
         );
  OAI211_X1 U9380 ( .C1(n7604), .C2(n7652), .A(n7603), .B(n8892), .ZN(n10268)
         );
  OAI211_X1 U9381 ( .C1(n10269), .C2(n10342), .A(n10275), .B(n10268), .ZN(
        n7654) );
  INV_X1 U9382 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7605) );
  OAI22_X1 U9383 ( .A1(n8956), .A2(n7652), .B1(n10345), .B2(n7605), .ZN(n7606)
         );
  AOI21_X1 U9384 ( .B1(n7654), .B2(n10345), .A(n7606), .ZN(n7607) );
  INV_X1 U9385 ( .A(n7607), .ZN(P2_U3460) );
  OAI222_X1 U9386 ( .A1(n8974), .A2(n7610), .B1(P2_U3152), .B2(n7609), .C1(
        n8977), .C2(n7608), .ZN(P2_U3337) );
  INV_X1 U9387 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7624) );
  XNOR2_X1 U9388 ( .A(n9467), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n9463) );
  XNOR2_X1 U9389 ( .A(n9463), .B(n9462), .ZN(n7622) );
  NAND2_X1 U9390 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7948) );
  INV_X1 U9391 ( .A(n7948), .ZN(n7621) );
  INV_X1 U9392 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7613) );
  XNOR2_X1 U9393 ( .A(n9467), .B(n7613), .ZN(n7618) );
  OR2_X1 U9394 ( .A1(n7614), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7616) );
  OAI211_X1 U9395 ( .C1(n7618), .C2(n7617), .A(n10143), .B(n9468), .ZN(n7619)
         );
  OAI21_X1 U9396 ( .B1(n10149), .B2(n4848), .A(n7619), .ZN(n7620) );
  AOI211_X1 U9397 ( .C1(n10190), .C2(n7622), .A(n7621), .B(n7620), .ZN(n7623)
         );
  OAI21_X1 U9398 ( .B1(n10195), .B2(n7624), .A(n7623), .ZN(P1_U3253) );
  INV_X1 U9399 ( .A(n4753), .ZN(n7627) );
  OAI21_X1 U9400 ( .B1(n4753), .B2(n4709), .A(n7625), .ZN(n7626) );
  OAI21_X1 U9401 ( .B1(n7627), .B2(n9118), .A(n7626), .ZN(n7632) );
  OAI21_X1 U9402 ( .B1(n7630), .B2(n7629), .A(n7628), .ZN(n7631) );
  XNOR2_X1 U9403 ( .A(n7632), .B(n7631), .ZN(n7633) );
  NAND2_X1 U9404 ( .A1(n7633), .A2(n9145), .ZN(n7640) );
  INV_X1 U9405 ( .A(n7634), .ZN(n7635) );
  OAI22_X1 U9406 ( .A1(n9113), .A2(n7636), .B1(n9146), .B2(n7635), .ZN(n7637)
         );
  AOI211_X1 U9407 ( .C1(n9125), .C2(n9454), .A(n7638), .B(n7637), .ZN(n7639)
         );
  OAI211_X1 U9408 ( .C1(n7641), .C2(n9153), .A(n7640), .B(n7639), .ZN(P1_U3211) );
  INV_X1 U9409 ( .A(n8204), .ZN(n7642) );
  AOI211_X1 U9410 ( .C1(n7644), .C2(n7643), .A(n8377), .B(n7642), .ZN(n7650)
         );
  INV_X1 U9411 ( .A(n7645), .ZN(n7646) );
  OAI22_X1 U9412 ( .A1(n8374), .A2(n7646), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9937), .ZN(n7649) );
  INV_X1 U9413 ( .A(n8372), .ZN(n8389) );
  INV_X1 U9414 ( .A(n7820), .ZN(n7647) );
  OAI22_X1 U9415 ( .A1(n7823), .A2(n8364), .B1(n8389), .B2(n7647), .ZN(n7648)
         );
  OR3_X1 U9416 ( .A1(n7650), .A2(n7649), .A3(n7648), .ZN(P2_U3215) );
  OAI22_X1 U9417 ( .A1(n8885), .A2(n7652), .B1(n10352), .B2(n7651), .ZN(n7653)
         );
  AOI21_X1 U9418 ( .B1(n7654), .B2(n10352), .A(n7653), .ZN(n7655) );
  INV_X1 U9419 ( .A(n7655), .ZN(P2_U3523) );
  INV_X1 U9420 ( .A(n7656), .ZN(n7659) );
  NOR3_X1 U9421 ( .A1(n8353), .A2(n7893), .A3(n7657), .ZN(n7658) );
  AOI21_X1 U9422 ( .B1(n7659), .B2(n8380), .A(n7658), .ZN(n7669) );
  INV_X1 U9423 ( .A(n7660), .ZN(n7666) );
  OR2_X1 U9424 ( .A1(n7893), .A2(n8383), .ZN(n7661) );
  OAI21_X1 U9425 ( .B1(n7973), .B2(n8385), .A(n7661), .ZN(n7901) );
  INV_X1 U9426 ( .A(n7901), .ZN(n7664) );
  AOI22_X1 U9427 ( .A1(n8392), .A2(n8891), .B1(n7904), .B2(n8372), .ZN(n7663)
         );
  OAI211_X1 U9428 ( .C1(n7664), .C2(n8374), .A(n7663), .B(n7662), .ZN(n7665)
         );
  AOI21_X1 U9429 ( .B1(n7666), .B2(n8380), .A(n7665), .ZN(n7667) );
  OAI21_X1 U9430 ( .B1(n7669), .B2(n7668), .A(n7667), .ZN(P2_U3233) );
  XOR2_X1 U9431 ( .A(n7671), .B(n7670), .Z(n7680) );
  NAND2_X1 U9432 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n7853) );
  INV_X1 U9433 ( .A(n7853), .ZN(n7672) );
  AOI21_X1 U9434 ( .B1(n10258), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7672), .ZN(
        n7673) );
  OAI21_X1 U9435 ( .B1(n7674), .B2(n10260), .A(n7673), .ZN(n7679) );
  AOI211_X1 U9436 ( .C1(n7677), .C2(n7676), .A(n10259), .B(n7675), .ZN(n7678)
         );
  AOI211_X1 U9437 ( .C1(n10255), .C2(n7680), .A(n7679), .B(n7678), .ZN(n7681)
         );
  INV_X1 U9438 ( .A(n7681), .ZN(P2_U3255) );
  NAND2_X1 U9439 ( .A1(n7527), .A2(n10236), .ZN(n7682) );
  NAND2_X1 U9440 ( .A1(n7866), .A2(n7682), .ZN(n10240) );
  NAND2_X1 U9441 ( .A1(n7683), .A2(n9166), .ZN(n7684) );
  XNOR2_X1 U9442 ( .A(n7684), .B(n9409), .ZN(n7685) );
  NAND2_X1 U9443 ( .A1(n7685), .A2(n9799), .ZN(n7692) );
  NAND2_X1 U9444 ( .A1(n7686), .A2(n9409), .ZN(n7687) );
  AND2_X1 U9445 ( .A1(n7688), .A2(n7687), .ZN(n7690) );
  OAI22_X1 U9446 ( .A1(n7794), .A2(n9772), .B1(n7858), .B2(n9770), .ZN(n7689)
         );
  AOI21_X1 U9447 ( .B1(n7690), .B2(n10234), .A(n7689), .ZN(n7691) );
  NAND2_X1 U9448 ( .A1(n7692), .A2(n7691), .ZN(n10241) );
  MUX2_X1 U9449 ( .A(n10241), .B(P1_REG2_REG_8__SCAN_IN), .S(n10211), .Z(n7693) );
  INV_X1 U9450 ( .A(n7693), .ZN(n7695) );
  AOI22_X1 U9451 ( .A1(n9758), .A2(n10236), .B1(n7792), .B2(n10201), .ZN(n7694) );
  OAI211_X1 U9452 ( .C1(n9762), .C2(n10240), .A(n7695), .B(n7694), .ZN(
        P1_U3283) );
  INV_X1 U9453 ( .A(n7696), .ZN(n7701) );
  AOI21_X1 U9454 ( .B1(n7698), .B2(n10047), .A(n7697), .ZN(n7699) );
  OAI211_X1 U9455 ( .C1(n9753), .C2(n7701), .A(n7700), .B(n7699), .ZN(n7704)
         );
  NAND2_X1 U9456 ( .A1(n7704), .A2(n10254), .ZN(n7702) );
  OAI21_X1 U9457 ( .B1(n10254), .B2(n7703), .A(n7702), .ZN(P1_U3530) );
  INV_X1 U9458 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9911) );
  NAND2_X1 U9459 ( .A1(n7704), .A2(n10245), .ZN(n7705) );
  OAI21_X1 U9460 ( .B1(n10245), .B2(n9911), .A(n7705), .ZN(P1_U3475) );
  XOR2_X1 U9461 ( .A(n7707), .B(n7706), .Z(n7712) );
  AOI22_X1 U9462 ( .A1(n9150), .A2(n9453), .B1(n9134), .B2(n7765), .ZN(n7709)
         );
  OAI211_X1 U9463 ( .C1(n8009), .C2(n9148), .A(n7709), .B(n7708), .ZN(n7710)
         );
  AOI21_X1 U9464 ( .B1(n10043), .B2(n9138), .A(n7710), .ZN(n7711) );
  OAI21_X1 U9465 ( .B1(n7712), .B2(n9140), .A(n7711), .ZN(P1_U3215) );
  INV_X1 U9466 ( .A(n7713), .ZN(n7714) );
  NOR3_X1 U9467 ( .A1(n10303), .A2(n7715), .A3(n7714), .ZN(n7716) );
  NAND2_X1 U9468 ( .A1(n7717), .A2(n7716), .ZN(n7749) );
  INV_X4 U9469 ( .A(n8763), .ZN(n10276) );
  INV_X1 U9470 ( .A(n7718), .ZN(n7720) );
  NAND2_X1 U9471 ( .A1(n7720), .A2(n7719), .ZN(n7721) );
  INV_X1 U9472 ( .A(n7749), .ZN(n7724) );
  NAND2_X1 U9473 ( .A1(n7724), .A2(n7723), .ZN(n10281) );
  AOI22_X1 U9474 ( .A1(n8766), .A2(n7725), .B1(n8311), .B2(n10267), .ZN(n7729)
         );
  NAND2_X1 U9475 ( .A1(n10286), .A2(n8312), .ZN(n7728) );
  NAND2_X1 U9476 ( .A1(n10276), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7727) );
  NAND3_X1 U9477 ( .A1(n7729), .A2(n7728), .A3(n7727), .ZN(n7730) );
  AOI21_X1 U9478 ( .B1(n10284), .B2(n7731), .A(n7730), .ZN(n7732) );
  OAI21_X1 U9479 ( .B1(n10276), .B2(n7733), .A(n7732), .ZN(P2_U3292) );
  INV_X1 U9480 ( .A(n7734), .ZN(n8100) );
  OAI222_X1 U9481 ( .A1(n10094), .A2(n7736), .B1(n10087), .B2(n8100), .C1(
        P1_U3084), .C2(n7735), .ZN(P1_U3331) );
  XNOR2_X1 U9482 ( .A(n7737), .B(n7738), .ZN(n7740) );
  NAND2_X1 U9483 ( .A1(n8419), .A2(n8324), .ZN(n7739) );
  OAI21_X1 U9484 ( .B1(n8206), .B2(n8385), .A(n7739), .ZN(n8075) );
  AOI21_X1 U9485 ( .B1(n7740), .B2(n10290), .A(n8075), .ZN(n10333) );
  OR2_X1 U9486 ( .A1(n7742), .A2(n7741), .ZN(n7743) );
  NAND2_X1 U9487 ( .A1(n7744), .A2(n7743), .ZN(n10332) );
  NOR2_X1 U9488 ( .A1(n7745), .A2(n10327), .ZN(n7746) );
  OR2_X1 U9489 ( .A1(n7747), .A2(n7746), .ZN(n10329) );
  NOR2_X1 U9490 ( .A1(n7749), .A2(n7748), .ZN(n7908) );
  INV_X1 U9491 ( .A(n7908), .ZN(n8064) );
  NAND2_X1 U9492 ( .A1(n10286), .A2(n7750), .ZN(n7752) );
  AOI22_X1 U9493 ( .A1(n10276), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n8071), .B2(
        n10267), .ZN(n7751) );
  OAI211_X1 U9494 ( .C1(n10329), .C2(n8064), .A(n7752), .B(n7751), .ZN(n7753)
         );
  AOI21_X1 U9495 ( .B1(n10332), .B2(n10284), .A(n7753), .ZN(n7754) );
  OAI21_X1 U9496 ( .B1(n10333), .B2(n10276), .A(n7754), .ZN(P2_U3290) );
  NAND2_X1 U9497 ( .A1(n7758), .A2(n10089), .ZN(n7756) );
  OR2_X1 U9498 ( .A1(n7755), .A2(P1_U3084), .ZN(n9437) );
  OAI211_X1 U9499 ( .C1(n7757), .C2(n10094), .A(n7756), .B(n9437), .ZN(
        P1_U3330) );
  NAND2_X1 U9500 ( .A1(n7758), .A2(n8960), .ZN(n7760) );
  OAI211_X1 U9501 ( .C1(n7761), .C2(n8974), .A(n7760), .B(n7759), .ZN(P2_U3335) );
  INV_X1 U9502 ( .A(n9179), .ZN(n9411) );
  XNOR2_X1 U9503 ( .A(n7762), .B(n9411), .ZN(n10045) );
  XNOR2_X1 U9504 ( .A(n7763), .B(n9411), .ZN(n7764) );
  OAI222_X1 U9505 ( .A1(n9772), .A2(n7858), .B1(n9770), .B2(n8009), .C1(n9767), 
        .C2(n7764), .ZN(n10041) );
  NAND2_X1 U9506 ( .A1(n10041), .A2(n10209), .ZN(n7770) );
  AOI211_X1 U9507 ( .C1(n10043), .C2(n7864), .A(n10239), .B(n7910), .ZN(n10042) );
  AOI22_X1 U9508 ( .A1(n10211), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7765), .B2(
        n10201), .ZN(n7766) );
  OAI21_X1 U9509 ( .B1(n7767), .B2(n9789), .A(n7766), .ZN(n7768) );
  AOI21_X1 U9510 ( .B1(n10042), .B2(n9780), .A(n7768), .ZN(n7769) );
  OAI211_X1 U9511 ( .C1(n10045), .C2(n9804), .A(n7770), .B(n7769), .ZN(
        P1_U3281) );
  INV_X1 U9512 ( .A(n7771), .ZN(n7772) );
  NAND2_X1 U9513 ( .A1(n7773), .A2(n7772), .ZN(n7787) );
  NOR2_X1 U9514 ( .A1(n7773), .A2(n7772), .ZN(n7786) );
  AOI21_X1 U9515 ( .B1(n7774), .B2(n7787), .A(n7786), .ZN(n7778) );
  XNOR2_X1 U9516 ( .A(n7776), .B(n7775), .ZN(n7777) );
  XNOR2_X1 U9517 ( .A(n7778), .B(n7777), .ZN(n7785) );
  INV_X1 U9518 ( .A(n7779), .ZN(n7867) );
  OAI22_X1 U9519 ( .A1(n9113), .A2(n7780), .B1(n9146), .B2(n7867), .ZN(n7781)
         );
  AOI211_X1 U9520 ( .C1(n9125), .C2(n9452), .A(n7782), .B(n7781), .ZN(n7784)
         );
  NAND2_X1 U9521 ( .A1(n9138), .A2(n10048), .ZN(n7783) );
  OAI211_X1 U9522 ( .C1(n7785), .C2(n9140), .A(n7784), .B(n7783), .ZN(P1_U3229) );
  INV_X1 U9523 ( .A(n7786), .ZN(n7788) );
  NAND2_X1 U9524 ( .A1(n7788), .A2(n7787), .ZN(n7790) );
  XNOR2_X1 U9525 ( .A(n7790), .B(n7789), .ZN(n7798) );
  NOR2_X1 U9526 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7791), .ZN(n10127) );
  INV_X1 U9527 ( .A(n7792), .ZN(n7793) );
  OAI22_X1 U9528 ( .A1(n9113), .A2(n7794), .B1(n9146), .B2(n7793), .ZN(n7795)
         );
  AOI211_X1 U9529 ( .C1(n9125), .C2(n9453), .A(n10127), .B(n7795), .ZN(n7797)
         );
  NAND2_X1 U9530 ( .A1(n9138), .A2(n10236), .ZN(n7796) );
  OAI211_X1 U9531 ( .C1(n7798), .C2(n9140), .A(n7797), .B(n7796), .ZN(P1_U3219) );
  AOI22_X1 U9532 ( .A1(n10276), .A2(P2_REG2_REG_5__SCAN_IN), .B1(n8276), .B2(
        n10267), .ZN(n7801) );
  NAND2_X1 U9533 ( .A1(n7799), .A2(n8766), .ZN(n7800) );
  OAI211_X1 U9534 ( .C1(n8754), .C2(n7802), .A(n7801), .B(n7800), .ZN(n7803)
         );
  AOI21_X1 U9535 ( .B1(n10284), .B2(n7804), .A(n7803), .ZN(n7805) );
  OAI21_X1 U9536 ( .B1(n10276), .B2(n7806), .A(n7805), .ZN(P2_U3291) );
  XNOR2_X1 U9537 ( .A(n7808), .B(n7807), .ZN(n7818) );
  OAI21_X1 U9538 ( .B1(n7811), .B2(n7810), .A(n7809), .ZN(n7812) );
  NAND2_X1 U9539 ( .A1(n7812), .A2(n10256), .ZN(n7817) );
  AND2_X1 U9540 ( .A1(P2_U3152), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7815) );
  NOR2_X1 U9541 ( .A1(n10260), .A2(n7813), .ZN(n7814) );
  AOI211_X1 U9542 ( .C1(P2_ADDR_REG_11__SCAN_IN), .C2(n10258), .A(n7815), .B(
        n7814), .ZN(n7816) );
  OAI211_X1 U9543 ( .C1(n7818), .C2(n10261), .A(n7817), .B(n7816), .ZN(
        P2_U3256) );
  NAND2_X1 U9544 ( .A1(n7819), .A2(n8766), .ZN(n7822) );
  AOI22_X1 U9545 ( .A1(n10276), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n7820), .B2(
        n10267), .ZN(n7821) );
  OAI211_X1 U9546 ( .C1(n7823), .C2(n8754), .A(n7822), .B(n7821), .ZN(n7824)
         );
  AOI21_X1 U9547 ( .B1(n10284), .B2(n7825), .A(n7824), .ZN(n7826) );
  OAI21_X1 U9548 ( .B1(n7827), .B2(n10276), .A(n7826), .ZN(P2_U3289) );
  INV_X1 U9549 ( .A(n8206), .ZN(n8417) );
  OR2_X1 U9550 ( .A1(n8417), .A2(n7828), .ZN(n7829) );
  NAND2_X1 U9551 ( .A1(n7831), .A2(n6385), .ZN(n7832) );
  AND2_X1 U9552 ( .A1(n7895), .A2(n7832), .ZN(n7839) );
  INV_X1 U9553 ( .A(n7839), .ZN(n10341) );
  INV_X1 U9554 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7841) );
  INV_X1 U9555 ( .A(n7933), .ZN(n7840) );
  OR2_X1 U9556 ( .A1(n8206), .A2(n8383), .ZN(n7833) );
  OAI21_X1 U9557 ( .B1(n7927), .B2(n8385), .A(n7833), .ZN(n8210) );
  NAND2_X1 U9558 ( .A1(n7835), .A2(n7834), .ZN(n7836) );
  INV_X1 U9559 ( .A(n10290), .ZN(n8734) );
  AOI21_X1 U9560 ( .B1(n7837), .B2(n7836), .A(n8734), .ZN(n7838) );
  AOI211_X1 U9561 ( .C1(n7840), .C2(n7839), .A(n8210), .B(n7838), .ZN(n10340)
         );
  MUX2_X1 U9562 ( .A(n7841), .B(n10340), .S(n8763), .Z(n7848) );
  INV_X1 U9563 ( .A(n7903), .ZN(n7842) );
  AOI211_X1 U9564 ( .C1(n10337), .C2(n7843), .A(n10328), .B(n7842), .ZN(n10336) );
  INV_X1 U9565 ( .A(n10337), .ZN(n7845) );
  OAI22_X1 U9566 ( .A1(n8754), .A2(n7845), .B1(n10279), .B2(n7844), .ZN(n7846)
         );
  AOI21_X1 U9567 ( .B1(n10336), .B2(n8766), .A(n7846), .ZN(n7847) );
  OAI211_X1 U9568 ( .C1(n10341), .C2(n10270), .A(n7848), .B(n7847), .ZN(
        P2_U3288) );
  INV_X1 U9569 ( .A(n8887), .ZN(n7940) );
  AOI21_X1 U9570 ( .B1(n7850), .B2(n7849), .A(n8377), .ZN(n7851) );
  NAND2_X1 U9571 ( .A1(n7851), .A2(n7969), .ZN(n7857) );
  OR2_X1 U9572 ( .A1(n8232), .A2(n8385), .ZN(n7852) );
  OAI21_X1 U9573 ( .B1(n7927), .B2(n8383), .A(n7852), .ZN(n7935) );
  INV_X1 U9574 ( .A(n7935), .ZN(n7854) );
  OAI21_X1 U9575 ( .B1(n8374), .B2(n7854), .A(n7853), .ZN(n7855) );
  AOI21_X1 U9576 ( .B1(n7938), .B2(n8372), .A(n7855), .ZN(n7856) );
  OAI211_X1 U9577 ( .C1(n7940), .C2(n8364), .A(n7857), .B(n7856), .ZN(P2_U3219) );
  XNOR2_X1 U9578 ( .A(n10048), .B(n7858), .ZN(n9413) );
  XNOR2_X1 U9579 ( .A(n7859), .B(n9413), .ZN(n10051) );
  INV_X1 U9580 ( .A(n9413), .ZN(n7862) );
  NAND2_X1 U9581 ( .A1(n9175), .A2(n9296), .ZN(n7861) );
  MUX2_X1 U9582 ( .A(n7862), .B(n7861), .S(n7860), .Z(n7863) );
  AOI222_X1 U9583 ( .A1(n9799), .A2(n7863), .B1(n9452), .B2(n9796), .C1(n9454), 
        .C2(n9794), .ZN(n10050) );
  OR2_X1 U9584 ( .A1(n10050), .A2(n10211), .ZN(n7872) );
  INV_X1 U9585 ( .A(n7864), .ZN(n7865) );
  AOI211_X1 U9586 ( .C1(n10048), .C2(n7866), .A(n10239), .B(n7865), .ZN(n10046) );
  NOR2_X1 U9587 ( .A1(n9789), .A2(n5013), .ZN(n7870) );
  INV_X1 U9588 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7868) );
  OAI22_X1 U9589 ( .A1(n10209), .A2(n7868), .B1(n7867), .B2(n9755), .ZN(n7869)
         );
  AOI211_X1 U9590 ( .C1(n10046), .C2(n9651), .A(n7870), .B(n7869), .ZN(n7871)
         );
  OAI211_X1 U9591 ( .C1(n10051), .C2(n9804), .A(n7872), .B(n7871), .ZN(
        P1_U3282) );
  AOI21_X1 U9592 ( .B1(n7874), .B2(n7873), .A(n9140), .ZN(n7876) );
  NAND2_X1 U9593 ( .A1(n7876), .A2(n7875), .ZN(n7882) );
  INV_X1 U9594 ( .A(n7877), .ZN(n7918) );
  OAI22_X1 U9595 ( .A1(n9113), .A2(n7878), .B1(n9146), .B2(n7918), .ZN(n7879)
         );
  AOI211_X1 U9596 ( .C1(n9125), .C2(n9795), .A(n7880), .B(n7879), .ZN(n7881)
         );
  OAI211_X1 U9597 ( .C1(n7980), .C2(n9153), .A(n7882), .B(n7881), .ZN(P1_U3234) );
  INV_X1 U9598 ( .A(n10315), .ZN(n7890) );
  NAND2_X1 U9599 ( .A1(n10315), .A2(n10290), .ZN(n7884) );
  AND2_X1 U9600 ( .A1(n7884), .A2(n7883), .ZN(n10317) );
  OAI22_X1 U9601 ( .A1(n10276), .A2(n10317), .B1(n7885), .B2(n10279), .ZN(
        n7888) );
  AOI21_X1 U9602 ( .B1(n8754), .B2(n8064), .A(n7886), .ZN(n7887) );
  AOI211_X1 U9603 ( .C1(n10276), .C2(P2_REG2_REG_0__SCAN_IN), .A(n7888), .B(
        n7887), .ZN(n7889) );
  OAI21_X1 U9604 ( .B1(n7890), .B2(n8769), .A(n7889), .ZN(P2_U3296) );
  OAI21_X1 U9605 ( .B1(n7899), .B2(n7892), .A(n7891), .ZN(n7902) );
  INV_X1 U9606 ( .A(n7893), .ZN(n8416) );
  NAND2_X1 U9607 ( .A1(n8416), .A2(n10337), .ZN(n7894) );
  INV_X1 U9608 ( .A(n7899), .ZN(n7896) );
  INV_X1 U9609 ( .A(n7929), .ZN(n7897) );
  AOI21_X1 U9610 ( .B1(n7899), .B2(n7898), .A(n7897), .ZN(n8896) );
  NOR2_X1 U9611 ( .A1(n8896), .A2(n7933), .ZN(n7900) );
  AOI211_X1 U9612 ( .C1(n10290), .C2(n7902), .A(n7901), .B(n7900), .ZN(n8895)
         );
  AOI21_X1 U9613 ( .B1(n8891), .B2(n7903), .A(n7937), .ZN(n8893) );
  AOI22_X1 U9614 ( .A1(n10276), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7904), .B2(
        n10267), .ZN(n7905) );
  OAI21_X1 U9615 ( .B1(n8754), .B2(n5065), .A(n7905), .ZN(n7907) );
  NOR2_X1 U9616 ( .A1(n8896), .A2(n10270), .ZN(n7906) );
  AOI211_X1 U9617 ( .C1(n8893), .C2(n7908), .A(n7907), .B(n7906), .ZN(n7909)
         );
  OAI21_X1 U9618 ( .B1(n8895), .B2(n10276), .A(n7909), .ZN(P2_U3287) );
  OR2_X1 U9619 ( .A1(n7910), .A2(n7980), .ZN(n7911) );
  NAND2_X1 U9620 ( .A1(n8015), .A2(n7911), .ZN(n7981) );
  XNOR2_X1 U9621 ( .A(n7920), .B(n8009), .ZN(n9182) );
  INV_X1 U9622 ( .A(n9182), .ZN(n9415) );
  XNOR2_X1 U9623 ( .A(n7912), .B(n9415), .ZN(n7917) );
  XNOR2_X1 U9624 ( .A(n7913), .B(n9415), .ZN(n7914) );
  NAND2_X1 U9625 ( .A1(n7914), .A2(n9799), .ZN(n7916) );
  AOI22_X1 U9626 ( .A1(n9796), .A2(n9795), .B1(n9452), .B2(n9794), .ZN(n7915)
         );
  OAI211_X1 U9627 ( .C1(n9753), .C2(n7917), .A(n7916), .B(n7915), .ZN(n7983)
         );
  NAND2_X1 U9628 ( .A1(n7983), .A2(n10209), .ZN(n7922) );
  OAI22_X1 U9629 ( .A1(n10209), .A2(n7358), .B1(n7918), .B2(n9755), .ZN(n7919)
         );
  AOI21_X1 U9630 ( .B1(n9758), .B2(n7920), .A(n7919), .ZN(n7921) );
  OAI211_X1 U9631 ( .C1(n7981), .C2(n9762), .A(n7922), .B(n7921), .ZN(P1_U3280) );
  INV_X1 U9632 ( .A(n7923), .ZN(n8084) );
  OAI222_X1 U9633 ( .A1(n7925), .A2(P2_U3152), .B1(n8977), .B2(n8084), .C1(
        n7924), .C2(n8974), .ZN(P2_U3334) );
  XNOR2_X1 U9634 ( .A(n7926), .B(n7930), .ZN(n7936) );
  INV_X1 U9635 ( .A(n7927), .ZN(n8415) );
  OR2_X1 U9636 ( .A1(n8415), .A2(n8891), .ZN(n7928) );
  NAND2_X1 U9637 ( .A1(n7931), .A2(n7930), .ZN(n7932) );
  NAND2_X1 U9638 ( .A1(n7955), .A2(n7932), .ZN(n8890) );
  NOR2_X1 U9639 ( .A1(n8890), .A2(n7933), .ZN(n7934) );
  AOI211_X1 U9640 ( .C1(n7936), .C2(n10290), .A(n7935), .B(n7934), .ZN(n8889)
         );
  AOI211_X1 U9641 ( .C1(n8887), .C2(n5067), .A(n10328), .B(n8747), .ZN(n8886)
         );
  AOI22_X1 U9642 ( .A1(n10276), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n7938), .B2(
        n10267), .ZN(n7939) );
  OAI21_X1 U9643 ( .B1(n8754), .B2(n7940), .A(n7939), .ZN(n7942) );
  NOR2_X1 U9644 ( .A1(n8890), .A2(n10270), .ZN(n7941) );
  AOI211_X1 U9645 ( .C1(n8886), .C2(n8766), .A(n7942), .B(n7941), .ZN(n7943)
         );
  OAI21_X1 U9646 ( .B1(n8889), .B2(n10276), .A(n7943), .ZN(P2_U3286) );
  XNOR2_X1 U9647 ( .A(n7945), .B(n7944), .ZN(n7946) );
  XNOR2_X1 U9648 ( .A(n7947), .B(n7946), .ZN(n7953) );
  AOI22_X1 U9649 ( .A1(n9150), .A2(n9451), .B1(n9134), .B2(n8017), .ZN(n7949)
         );
  OAI211_X1 U9650 ( .C1(n9771), .C2(n9148), .A(n7949), .B(n7948), .ZN(n7950)
         );
  AOI21_X1 U9651 ( .B1(n7951), .B2(n9138), .A(n7950), .ZN(n7952) );
  OAI21_X1 U9652 ( .B1(n7953), .B2(n9140), .A(n7952), .ZN(P1_U3222) );
  INV_X1 U9653 ( .A(n7973), .ZN(n8414) );
  NAND2_X1 U9654 ( .A1(n8887), .A2(n8414), .ZN(n7954) );
  INV_X1 U9655 ( .A(n8232), .ZN(n8413) );
  NAND2_X1 U9656 ( .A1(n8751), .A2(n8413), .ZN(n7956) );
  XNOR2_X1 U9657 ( .A(n7990), .B(n7989), .ZN(n8877) );
  INV_X1 U9658 ( .A(n8877), .ZN(n7968) );
  OAI211_X1 U9659 ( .C1(n7959), .C2(n7989), .A(n7958), .B(n10290), .ZN(n7962)
         );
  OR2_X1 U9660 ( .A1(n8232), .A2(n8383), .ZN(n7961) );
  OR2_X1 U9661 ( .A1(n8171), .A2(n8385), .ZN(n7960) );
  AND2_X1 U9662 ( .A1(n7961), .A2(n7960), .ZN(n8239) );
  NAND2_X1 U9663 ( .A1(n7962), .A2(n8239), .ZN(n8875) );
  INV_X1 U9664 ( .A(n8243), .ZN(n8952) );
  INV_X1 U9665 ( .A(n8751), .ZN(n8957) );
  NAND2_X1 U9666 ( .A1(n8747), .A2(n8957), .ZN(n8748) );
  INV_X1 U9667 ( .A(n8000), .ZN(n7963) );
  AOI211_X1 U9668 ( .C1(n8243), .C2(n8748), .A(n10328), .B(n7963), .ZN(n8876)
         );
  NAND2_X1 U9669 ( .A1(n8876), .A2(n8766), .ZN(n7965) );
  AOI22_X1 U9670 ( .A1(n10276), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n8235), .B2(
        n10267), .ZN(n7964) );
  OAI211_X1 U9671 ( .C1(n8952), .C2(n8754), .A(n7965), .B(n7964), .ZN(n7966)
         );
  AOI21_X1 U9672 ( .B1(n8875), .B2(n8763), .A(n7966), .ZN(n7967) );
  OAI21_X1 U9673 ( .B1(n7968), .B2(n8769), .A(n7967), .ZN(P2_U3284) );
  AOI21_X1 U9674 ( .B1(n7969), .B2(n4410), .A(n8377), .ZN(n7972) );
  NOR3_X1 U9675 ( .A1(n8353), .A2(n7973), .A3(n7970), .ZN(n7971) );
  OAI21_X1 U9676 ( .B1(n7972), .B2(n7971), .A(n8230), .ZN(n7979) );
  OR2_X1 U9677 ( .A1(n7973), .A2(n8383), .ZN(n7975) );
  OR2_X1 U9678 ( .A1(n7997), .A2(n8385), .ZN(n7974) );
  AND2_X1 U9679 ( .A1(n7975), .A2(n7974), .ZN(n8761) );
  OAI22_X1 U9680 ( .A1(n8374), .A2(n8761), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7976), .ZN(n7977) );
  AOI21_X1 U9681 ( .B1(n8752), .B2(n8372), .A(n7977), .ZN(n7978) );
  OAI211_X1 U9682 ( .C1(n8957), .C2(n8364), .A(n7979), .B(n7978), .ZN(P2_U3238) );
  INV_X1 U9683 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7984) );
  OAI22_X1 U9684 ( .A1(n7981), .A2(n10239), .B1(n7980), .B2(n10237), .ZN(n7982) );
  NOR2_X1 U9685 ( .A1(n7983), .A2(n7982), .ZN(n7986) );
  MUX2_X1 U9686 ( .A(n7984), .B(n7986), .S(n10245), .Z(n7985) );
  INV_X1 U9687 ( .A(n7985), .ZN(P1_U3487) );
  MUX2_X1 U9688 ( .A(n7987), .B(n7986), .S(n10254), .Z(n7988) );
  INV_X1 U9689 ( .A(n7988), .ZN(P1_U3534) );
  INV_X1 U9690 ( .A(n7997), .ZN(n8412) );
  NAND2_X1 U9691 ( .A1(n7991), .A2(n6429), .ZN(n7992) );
  NAND2_X1 U9692 ( .A1(n8719), .A2(n7992), .ZN(n8869) );
  NAND2_X1 U9693 ( .A1(n7994), .A2(n7993), .ZN(n7995) );
  AOI21_X1 U9694 ( .B1(n7996), .B2(n7995), .A(n8734), .ZN(n7999) );
  OR2_X1 U9695 ( .A1(n7997), .A2(n8383), .ZN(n7998) );
  OAI21_X1 U9696 ( .B1(n8384), .B2(n8385), .A(n7998), .ZN(n8331) );
  OR2_X1 U9697 ( .A1(n7999), .A2(n8331), .ZN(n8867) );
  INV_X1 U9698 ( .A(n8946), .ZN(n8005) );
  NAND2_X1 U9699 ( .A1(n8000), .A2(n8946), .ZN(n8001) );
  NAND2_X1 U9700 ( .A1(n8001), .A2(n8892), .ZN(n8002) );
  NOR2_X1 U9701 ( .A1(n8736), .A2(n8002), .ZN(n8866) );
  NAND2_X1 U9702 ( .A1(n8866), .A2(n8766), .ZN(n8004) );
  AOI22_X1 U9703 ( .A1(n10276), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n8332), .B2(
        n10267), .ZN(n8003) );
  OAI211_X1 U9704 ( .C1(n8005), .C2(n8754), .A(n8004), .B(n8003), .ZN(n8006)
         );
  AOI21_X1 U9705 ( .B1(n8867), .B2(n8763), .A(n8006), .ZN(n8007) );
  OAI21_X1 U9706 ( .B1(n8769), .B2(n8869), .A(n8007), .ZN(P2_U3283) );
  XNOR2_X1 U9707 ( .A(n8008), .B(n9397), .ZN(n8014) );
  OAI22_X1 U9708 ( .A1(n9771), .A2(n9770), .B1(n8009), .B2(n9772), .ZN(n8013)
         );
  XNOR2_X1 U9709 ( .A(n8010), .B(n9397), .ZN(n8011) );
  NOR2_X1 U9710 ( .A1(n8011), .A2(n9753), .ZN(n8012) );
  AOI211_X1 U9711 ( .C1(n9799), .C2(n8014), .A(n8013), .B(n8012), .ZN(n10039)
         );
  INV_X1 U9712 ( .A(n8015), .ZN(n8016) );
  OAI211_X1 U9713 ( .C1(n10040), .C2(n8016), .A(n5216), .B(n10033), .ZN(n10038) );
  INV_X1 U9714 ( .A(n10038), .ZN(n8020) );
  AOI22_X1 U9715 ( .A1(n10211), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n8017), .B2(
        n10201), .ZN(n8018) );
  OAI21_X1 U9716 ( .B1(n10040), .B2(n9789), .A(n8018), .ZN(n8019) );
  AOI21_X1 U9717 ( .B1(n8020), .B2(n9780), .A(n8019), .ZN(n8021) );
  OAI21_X1 U9718 ( .B1(n10039), .B2(n10211), .A(n8021), .ZN(P1_U3279) );
  INV_X1 U9719 ( .A(n8022), .ZN(n8025) );
  OAI222_X1 U9720 ( .A1(n8974), .A2(n9863), .B1(n8977), .B2(n8025), .C1(n8023), 
        .C2(P2_U3152), .ZN(P2_U3333) );
  OAI222_X1 U9721 ( .A1(n10094), .A2(n9930), .B1(n10087), .B2(n8025), .C1(
        n8024), .C2(P1_U3084), .ZN(P1_U3328) );
  INV_X1 U9722 ( .A(n8429), .ZN(n8026) );
  OAI21_X1 U9723 ( .B1(n8028), .B2(n8027), .A(n8026), .ZN(n8036) );
  NOR2_X1 U9724 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8029), .ZN(n8236) );
  AOI21_X1 U9725 ( .B1(n10258), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n8236), .ZN(
        n8030) );
  OAI21_X1 U9726 ( .B1(n8031), .B2(n10260), .A(n8030), .ZN(n8035) );
  AOI211_X1 U9727 ( .C1(n8033), .C2(n8032), .A(n10259), .B(n4400), .ZN(n8034)
         );
  AOI211_X1 U9728 ( .C1(n10255), .C2(n8036), .A(n8035), .B(n8034), .ZN(n8037)
         );
  INV_X1 U9729 ( .A(n8037), .ZN(P2_U3257) );
  INV_X1 U9730 ( .A(n8038), .ZN(n8043) );
  AOI21_X1 U9731 ( .B1(n8042), .B2(n8040), .A(n8039), .ZN(n8041) );
  AOI21_X1 U9732 ( .B1(n8043), .B2(n8042), .A(n8041), .ZN(n8048) );
  AOI22_X1 U9733 ( .A1(n9150), .A2(n9795), .B1(n9134), .B2(n9787), .ZN(n8044)
         );
  NAND2_X1 U9734 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n10147) );
  OAI211_X1 U9735 ( .C1(n8045), .C2(n9148), .A(n8044), .B(n10147), .ZN(n8046)
         );
  AOI21_X1 U9736 ( .B1(n10032), .B2(n9138), .A(n8046), .ZN(n8047) );
  OAI21_X1 U9737 ( .B1(n8048), .B2(n9140), .A(n8047), .ZN(P1_U3232) );
  INV_X1 U9738 ( .A(n8049), .ZN(n8976) );
  OAI222_X1 U9739 ( .A1(n5894), .A2(P1_U3084), .B1(n10087), .B2(n8976), .C1(
        n9908), .C2(n10094), .ZN(P1_U3327) );
  OAI21_X1 U9740 ( .B1(n4337), .B2(n9767), .A(n8053), .ZN(n9812) );
  NAND2_X1 U9741 ( .A1(n9812), .A2(n10209), .ZN(n8061) );
  INV_X1 U9742 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n8054) );
  OAI22_X1 U9743 ( .A1(n8055), .A2(n9755), .B1(n8054), .B2(n10209), .ZN(n8058)
         );
  OAI21_X1 U9744 ( .B1(n9814), .B2(n4339), .A(n8056), .ZN(n9815) );
  NOR2_X1 U9745 ( .A1(n9815), .A2(n9762), .ZN(n8057) );
  AOI211_X1 U9746 ( .C1(n9758), .C2(n8059), .A(n8058), .B(n8057), .ZN(n8060)
         );
  OAI211_X1 U9747 ( .C1(n9783), .C2(n9813), .A(n8061), .B(n8060), .ZN(P1_U3263) );
  INV_X1 U9748 ( .A(n8062), .ZN(n8070) );
  INV_X1 U9749 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n8087) );
  OAI22_X1 U9750 ( .A1(n8064), .A2(n8063), .B1(n8087), .B2(n10279), .ZN(n8065)
         );
  AOI21_X1 U9751 ( .B1(n10286), .B2(n8090), .A(n8065), .ZN(n8069) );
  MUX2_X1 U9752 ( .A(n8067), .B(n8066), .S(n10276), .Z(n8068) );
  OAI211_X1 U9753 ( .C1(n8769), .C2(n8070), .A(n8069), .B(n8068), .ZN(P2_U3294) );
  INV_X1 U9754 ( .A(n8071), .ZN(n8072) );
  OAI22_X1 U9755 ( .A1(n10327), .A2(n8364), .B1(n8389), .B2(n8072), .ZN(n8073)
         );
  AOI211_X1 U9756 ( .C1(n8387), .C2(n8075), .A(n8074), .B(n8073), .ZN(n8081)
         );
  OAI22_X1 U9757 ( .A1(n8353), .A2(n8078), .B1(n8377), .B2(n8077), .ZN(n8079)
         );
  NAND3_X1 U9758 ( .A1(n8272), .A2(n4674), .A3(n8079), .ZN(n8080) );
  OAI211_X1 U9759 ( .C1(n8377), .C2(n8082), .A(n8081), .B(n8080), .ZN(P2_U3241) );
  OAI222_X1 U9760 ( .A1(n8085), .A2(P1_U3084), .B1(n10087), .B2(n8084), .C1(
        n8083), .C2(n10094), .ZN(P1_U3329) );
  OAI22_X1 U9761 ( .A1(n8088), .A2(n8087), .B1(n8374), .B2(n8086), .ZN(n8089)
         );
  AOI21_X1 U9762 ( .B1(n8090), .B2(n8392), .A(n8089), .ZN(n8097) );
  OAI22_X1 U9763 ( .A1(n8353), .A2(n6304), .B1(n8377), .B2(n8091), .ZN(n8095)
         );
  INV_X1 U9764 ( .A(n8092), .ZN(n8093) );
  NAND3_X1 U9765 ( .A1(n8095), .A2(n8094), .A3(n8093), .ZN(n8096) );
  OAI211_X1 U9766 ( .C1(n8377), .C2(n8098), .A(n8097), .B(n8096), .ZN(P2_U3239) );
  OAI222_X1 U9767 ( .A1(n8974), .A2(n8101), .B1(n8977), .B2(n8100), .C1(n8099), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  INV_X1 U9768 ( .A(n8802), .ZN(n8564) );
  INV_X1 U9769 ( .A(n8938), .ZN(n8725) );
  INV_X1 U9770 ( .A(n8834), .ZN(n8650) );
  NOR2_X2 U9771 ( .A1(n8558), .A2(n8543), .ZN(n8542) );
  INV_X1 U9772 ( .A(n8793), .ZN(n8530) );
  XNOR2_X1 U9773 ( .A(n8900), .B(n8501), .ZN(n8102) );
  NAND2_X1 U9774 ( .A1(n8102), .A2(n8892), .ZN(n8770) );
  NOR2_X1 U9775 ( .A1(n8971), .A2(n9917), .ZN(n8103) );
  NOR2_X1 U9776 ( .A1(n8385), .A2(n8103), .ZN(n8108) );
  NAND2_X1 U9777 ( .A1(n8104), .A2(n8108), .ZN(n8773) );
  NOR2_X1 U9778 ( .A1(n10276), .A2(n8773), .ZN(n8505) );
  NOR2_X1 U9779 ( .A1(n8900), .A2(n8754), .ZN(n8105) );
  AOI211_X1 U9780 ( .C1(n10276), .C2(P2_REG2_REG_31__SCAN_IN), .A(n8505), .B(
        n8105), .ZN(n8106) );
  OAI21_X1 U9781 ( .B1(n8770), .B2(n10281), .A(n8106), .ZN(P2_U3265) );
  INV_X1 U9782 ( .A(n8107), .ZN(n8396) );
  NAND2_X1 U9783 ( .A1(n8396), .A2(n8108), .ZN(n8109) );
  NOR2_X1 U9784 ( .A1(n8739), .A2(n8410), .ZN(n8720) );
  NAND2_X1 U9785 ( .A1(n8946), .A2(n8411), .ZN(n8718) );
  NAND2_X1 U9786 ( .A1(n8718), .A2(n8384), .ZN(n8113) );
  NAND2_X1 U9787 ( .A1(n8113), .A2(n8739), .ZN(n8114) );
  OAI21_X1 U9788 ( .B1(n8384), .B2(n8718), .A(n8114), .ZN(n8115) );
  NOR2_X1 U9789 ( .A1(n8721), .A2(n8115), .ZN(n8116) );
  INV_X1 U9790 ( .A(n8117), .ZN(n8409) );
  OR2_X1 U9791 ( .A1(n8938), .A2(n8409), .ZN(n8118) );
  NAND2_X1 U9792 ( .A1(n8933), .A2(n4621), .ZN(n8120) );
  OR2_X1 U9793 ( .A1(n8930), .A2(n8408), .ZN(n8121) );
  INV_X1 U9794 ( .A(n8926), .ZN(n8675) );
  INV_X1 U9795 ( .A(n8288), .ZN(n8407) );
  NOR2_X1 U9796 ( .A1(n8618), .A2(n8346), .ZN(n8124) );
  INV_X1 U9797 ( .A(n8346), .ZN(n8404) );
  NAND2_X1 U9798 ( .A1(n8813), .A2(n8402), .ZN(n8550) );
  NAND2_X1 U9799 ( .A1(n8811), .A2(n5213), .ZN(n8128) );
  INV_X1 U9800 ( .A(n8299), .ZN(n8401) );
  OR2_X1 U9801 ( .A1(n8575), .A2(n8401), .ZN(n8551) );
  INV_X1 U9802 ( .A(n8368), .ZN(n8400) );
  INV_X1 U9803 ( .A(n8536), .ZN(n8534) );
  INV_X1 U9804 ( .A(n8367), .ZN(n8398) );
  NAND2_X1 U9805 ( .A1(n8139), .A2(n8141), .ZN(n8788) );
  NOR2_X1 U9806 ( .A1(n8149), .A2(n8397), .ZN(n8779) );
  INV_X1 U9807 ( .A(n8779), .ZN(n8780) );
  NAND2_X1 U9808 ( .A1(n8788), .A2(n8780), .ZN(n8131) );
  XNOR2_X1 U9809 ( .A(n8131), .B(n4740), .ZN(n8137) );
  AOI21_X1 U9810 ( .B1(n8781), .B2(n4270), .A(n10328), .ZN(n8132) );
  NAND2_X1 U9811 ( .A1(n8503), .A2(n8132), .ZN(n8782) );
  AOI22_X1 U9812 ( .A1(n8133), .A2(n10267), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n10276), .ZN(n8135) );
  NAND2_X1 U9813 ( .A1(n8781), .A2(n10286), .ZN(n8134) );
  OAI211_X1 U9814 ( .C1(n8782), .C2(n10281), .A(n8135), .B(n8134), .ZN(n8136)
         );
  OAI21_X1 U9815 ( .B1(n8789), .B2(n10276), .A(n8138), .ZN(P2_U3267) );
  INV_X1 U9816 ( .A(n8140), .ZN(n8142) );
  AOI21_X1 U9817 ( .B1(n8142), .B2(n8141), .A(n8734), .ZN(n8145) );
  AOI21_X1 U9818 ( .B1(n8145), .B2(n8144), .A(n8143), .ZN(n8516) );
  OAI211_X1 U9819 ( .C1(n6587), .C2(n8525), .A(n4270), .B(n8892), .ZN(n8509)
         );
  NAND2_X1 U9820 ( .A1(n8149), .A2(n8873), .ZN(n8146) );
  NAND2_X1 U9821 ( .A1(n8147), .A2(n8146), .ZN(P2_U3548) );
  INV_X1 U9822 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8148) );
  NAND2_X1 U9823 ( .A1(n8149), .A2(n8947), .ZN(n8150) );
  NAND2_X1 U9824 ( .A1(n8151), .A2(n8150), .ZN(P2_U3516) );
  INV_X1 U9825 ( .A(n8152), .ZN(n8968) );
  OAI222_X1 U9826 ( .A1(n10094), .A2(n8153), .B1(n10087), .B2(n8968), .C1(
        n5815), .C2(P1_U3084), .ZN(P1_U3325) );
  INV_X1 U9827 ( .A(n9254), .ZN(n10083) );
  OAI222_X1 U9828 ( .A1(n8974), .A2(n8156), .B1(n8977), .B2(n10083), .C1(n8155), .C2(P2_U3152), .ZN(P2_U3328) );
  XNOR2_X1 U9829 ( .A(n8158), .B(n8157), .ZN(n8164) );
  NAND2_X1 U9830 ( .A1(n8397), .A2(n8360), .ZN(n8160) );
  NAND2_X1 U9831 ( .A1(n8399), .A2(n8324), .ZN(n8159) );
  AND2_X1 U9832 ( .A1(n8160), .A2(n8159), .ZN(n8522) );
  AOI22_X1 U9833 ( .A1(n8527), .A2(n8372), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n8161) );
  OAI21_X1 U9834 ( .B1(n8522), .B2(n8374), .A(n8161), .ZN(n8162) );
  AOI21_X1 U9835 ( .B1(n8793), .B2(n8392), .A(n8162), .ZN(n8163) );
  OAI21_X1 U9836 ( .B1(n8164), .B2(n8377), .A(n8163), .ZN(P2_U3216) );
  XNOR2_X1 U9837 ( .A(n8166), .B(n8165), .ZN(n8246) );
  NAND3_X1 U9838 ( .A1(n8230), .A2(n8246), .A3(n8167), .ZN(n8240) );
  NAND2_X1 U9839 ( .A1(n8240), .A2(n8168), .ZN(n8336) );
  NAND2_X1 U9840 ( .A1(n8170), .A2(n8169), .ZN(n8337) );
  NOR2_X1 U9841 ( .A1(n8336), .A2(n8337), .ZN(n8335) );
  NOR3_X1 U9842 ( .A1(n8172), .A2(n8171), .A3(n8353), .ZN(n8173) );
  AOI21_X1 U9843 ( .B1(n8335), .B2(n8380), .A(n8173), .ZN(n8179) );
  AOI22_X1 U9844 ( .A1(n8360), .A2(n8409), .B1(n8411), .B2(n8324), .ZN(n8733)
         );
  NAND2_X1 U9845 ( .A1(n8372), .A2(n8740), .ZN(n8174) );
  NAND2_X1 U9846 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8446) );
  OAI211_X1 U9847 ( .C1(n8374), .C2(n8733), .A(n8174), .B(n8446), .ZN(n8177)
         );
  NOR2_X1 U9848 ( .A1(n8175), .A2(n8377), .ZN(n8176) );
  AOI211_X1 U9849 ( .C1(n8739), .C2(n8392), .A(n8177), .B(n8176), .ZN(n8178)
         );
  OAI21_X1 U9850 ( .B1(n8180), .B2(n8179), .A(n8178), .ZN(P2_U3217) );
  INV_X1 U9851 ( .A(n8353), .ZN(n8379) );
  AOI22_X1 U9852 ( .A1(n8182), .A2(n8380), .B1(n8379), .B2(n8402), .ZN(n8189)
         );
  OR2_X1 U9853 ( .A1(n8299), .A2(n8385), .ZN(n8184) );
  NAND2_X1 U9854 ( .A1(n8403), .A2(n8324), .ZN(n8183) );
  NAND2_X1 U9855 ( .A1(n8184), .A2(n8183), .ZN(n8585) );
  OAI22_X1 U9856 ( .A1(n8389), .A2(n8590), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8185), .ZN(n8186) );
  AOI21_X1 U9857 ( .B1(n8585), .B2(n8387), .A(n8186), .ZN(n8188) );
  NAND2_X1 U9858 ( .A1(n8813), .A2(n8392), .ZN(n8187) );
  OAI211_X1 U9859 ( .C1(n4322), .C2(n8189), .A(n8188), .B(n8187), .ZN(P2_U3218) );
  INV_X1 U9860 ( .A(n8321), .ZN(n8196) );
  INV_X1 U9861 ( .A(n8190), .ZN(n8192) );
  NAND2_X1 U9862 ( .A1(n8192), .A2(n8191), .ZN(n8194) );
  AOI22_X1 U9863 ( .A1(n8196), .A2(n8195), .B1(n8194), .B2(n8193), .ZN(n8203)
         );
  INV_X1 U9864 ( .A(n8223), .ZN(n8405) );
  AOI22_X1 U9865 ( .A1(n8405), .A2(n8360), .B1(n8324), .B2(n8407), .ZN(n8648)
         );
  INV_X1 U9866 ( .A(n8648), .ZN(n8197) );
  AOI22_X1 U9867 ( .A1(n8387), .A2(n8197), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3152), .ZN(n8198) );
  OAI21_X1 U9868 ( .B1(n8654), .B2(n8389), .A(n8198), .ZN(n8201) );
  NOR3_X1 U9869 ( .A1(n8321), .A2(n8199), .A3(n8353), .ZN(n8200) );
  AOI211_X1 U9870 ( .C1(n8834), .C2(n8392), .A(n8201), .B(n8200), .ZN(n8202)
         );
  OAI21_X1 U9871 ( .B1(n8203), .B2(n8377), .A(n8202), .ZN(P2_U3221) );
  AOI21_X1 U9872 ( .B1(n8204), .B2(n4411), .A(n8377), .ZN(n8208) );
  NOR3_X1 U9873 ( .A1(n8353), .A2(n8206), .A3(n8205), .ZN(n8207) );
  OAI21_X1 U9874 ( .B1(n8208), .B2(n8207), .A(n7656), .ZN(n8214) );
  AOI22_X1 U9875 ( .A1(n8392), .A2(n10337), .B1(n8372), .B2(n8209), .ZN(n8212)
         );
  NAND2_X1 U9876 ( .A1(n8387), .A2(n8210), .ZN(n8211) );
  NAND4_X1 U9877 ( .A1(n8214), .A2(n8213), .A3(n8212), .A4(n8211), .ZN(
        P2_U3223) );
  INV_X1 U9878 ( .A(n8218), .ZN(n8215) );
  AOI21_X1 U9879 ( .B1(n8320), .B2(n8215), .A(n8377), .ZN(n8222) );
  NOR3_X1 U9880 ( .A1(n8216), .A2(n8223), .A3(n8353), .ZN(n8221) );
  NAND2_X1 U9881 ( .A1(n8320), .A2(n8217), .ZN(n8219) );
  NAND2_X1 U9882 ( .A1(n8219), .A2(n8218), .ZN(n8220) );
  OAI21_X1 U9883 ( .B1(n8222), .B2(n8221), .A(n8220), .ZN(n8229) );
  OAI22_X1 U9884 ( .A1(n8224), .A2(n8385), .B1(n8223), .B2(n8383), .ZN(n8621)
         );
  INV_X1 U9885 ( .A(n8621), .ZN(n8226) );
  OAI22_X1 U9886 ( .A1(n8226), .A2(n8374), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8225), .ZN(n8227) );
  AOI21_X1 U9887 ( .B1(n8616), .B2(n8372), .A(n8227), .ZN(n8228) );
  OAI211_X1 U9888 ( .C1(n8618), .C2(n8364), .A(n8229), .B(n8228), .ZN(P2_U3225) );
  INV_X1 U9889 ( .A(n8230), .ZN(n8234) );
  NOR3_X1 U9890 ( .A1(n8353), .A2(n8232), .A3(n8231), .ZN(n8233) );
  AOI21_X1 U9891 ( .B1(n8234), .B2(n8380), .A(n8233), .ZN(n8245) );
  NAND2_X1 U9892 ( .A1(n8372), .A2(n8235), .ZN(n8238) );
  INV_X1 U9893 ( .A(n8236), .ZN(n8237) );
  OAI211_X1 U9894 ( .C1(n8374), .C2(n8239), .A(n8238), .B(n8237), .ZN(n8242)
         );
  NOR2_X1 U9895 ( .A1(n8240), .A2(n8377), .ZN(n8241) );
  AOI211_X1 U9896 ( .C1(n8243), .C2(n8392), .A(n8242), .B(n8241), .ZN(n8244)
         );
  OAI21_X1 U9897 ( .B1(n8246), .B2(n8245), .A(n8244), .ZN(P2_U3226) );
  OR3_X1 U9898 ( .A1(n5124), .A2(n8248), .A3(n8377), .ZN(n8253) );
  NOR3_X1 U9899 ( .A1(n8249), .A2(n8368), .A3(n8353), .ZN(n8250) );
  AOI21_X1 U9900 ( .B1(n8380), .B2(n5124), .A(n8250), .ZN(n8252) );
  MUX2_X1 U9901 ( .A(n8253), .B(n8252), .S(n8251), .Z(n8257) );
  AOI22_X1 U9902 ( .A1(n8399), .A2(n8360), .B1(n8324), .B2(n8401), .ZN(n8556)
         );
  AOI22_X1 U9903 ( .A1(n8561), .A2(n8372), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8254) );
  OAI21_X1 U9904 ( .B1(n8556), .B2(n8374), .A(n8254), .ZN(n8255) );
  AOI21_X1 U9905 ( .B1(n8802), .B2(n8392), .A(n8255), .ZN(n8256) );
  NAND2_X1 U9906 ( .A1(n8257), .A2(n8256), .ZN(P2_U3227) );
  XNOR2_X1 U9907 ( .A(n4725), .B(n8258), .ZN(n8381) );
  NAND2_X1 U9908 ( .A1(n8381), .A2(n8259), .ZN(n8382) );
  OAI21_X1 U9909 ( .B1(n8261), .B2(n4725), .A(n8382), .ZN(n8265) );
  XNOR2_X1 U9910 ( .A(n8263), .B(n8262), .ZN(n8264) );
  XNOR2_X1 U9911 ( .A(n8265), .B(n8264), .ZN(n8271) );
  OR2_X1 U9912 ( .A1(n8358), .A2(n8385), .ZN(n8267) );
  NAND2_X1 U9913 ( .A1(n8409), .A2(n8324), .ZN(n8266) );
  NAND2_X1 U9914 ( .A1(n8267), .A2(n8266), .ZN(n8697) );
  AOI22_X1 U9915 ( .A1(n8387), .A2(n8697), .B1(P2_REG3_REG_16__SCAN_IN), .B2(
        P2_U3152), .ZN(n8268) );
  OAI21_X1 U9916 ( .B1(n8706), .B2(n8389), .A(n8268), .ZN(n8269) );
  AOI21_X1 U9917 ( .B1(n8933), .B2(n8392), .A(n8269), .ZN(n8270) );
  OAI21_X1 U9918 ( .B1(n8271), .B2(n8377), .A(n8270), .ZN(P2_U3228) );
  INV_X1 U9919 ( .A(n8272), .ZN(n8273) );
  NAND2_X1 U9920 ( .A1(n8273), .A2(n8380), .ZN(n8285) );
  AOI21_X1 U9921 ( .B1(n8387), .B2(n8275), .A(n8274), .ZN(n8284) );
  AOI22_X1 U9922 ( .A1(n8392), .A2(n8277), .B1(n8276), .B2(n8372), .ZN(n8283)
         );
  OAI22_X1 U9923 ( .A1(n8353), .A2(n6340), .B1(n8377), .B2(n8278), .ZN(n8281)
         );
  INV_X1 U9924 ( .A(n8279), .ZN(n8280) );
  NAND3_X1 U9925 ( .A1(n8281), .A2(n8307), .A3(n8280), .ZN(n8282) );
  NAND4_X1 U9926 ( .A1(n8285), .A2(n8284), .A3(n8283), .A4(n8282), .ZN(
        P2_U3229) );
  OAI211_X1 U9927 ( .C1(n8287), .C2(n8286), .A(n8352), .B(n8380), .ZN(n8295)
         );
  OR2_X1 U9928 ( .A1(n8288), .A2(n8385), .ZN(n8290) );
  NAND2_X1 U9929 ( .A1(n4621), .A2(n8324), .ZN(n8289) );
  NAND2_X1 U9930 ( .A1(n8290), .A2(n8289), .ZN(n8681) );
  INV_X1 U9931 ( .A(n8681), .ZN(n8292) );
  OAI22_X1 U9932 ( .A1(n8374), .A2(n8292), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8291), .ZN(n8293) );
  AOI21_X1 U9933 ( .B1(n8690), .B2(n8372), .A(n8293), .ZN(n8294) );
  OAI211_X1 U9934 ( .C1(n5078), .C2(n8364), .A(n8295), .B(n8294), .ZN(P2_U3230) );
  NOR2_X1 U9935 ( .A1(n4322), .A2(n8296), .ZN(n8298) );
  XNOR2_X1 U9936 ( .A(n8298), .B(n8297), .ZN(n8301) );
  OR2_X1 U9937 ( .A1(n8368), .A2(n8385), .ZN(n8303) );
  NAND2_X1 U9938 ( .A1(n8402), .A2(n8324), .ZN(n8302) );
  AND2_X1 U9939 ( .A1(n8303), .A2(n8302), .ZN(n8572) );
  OAI22_X1 U9940 ( .A1(n8572), .A2(n8374), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8304), .ZN(n8305) );
  AOI21_X1 U9941 ( .B1(n8576), .B2(n8372), .A(n8305), .ZN(n8306) );
  OAI21_X1 U9942 ( .B1(n8313), .B2(n8308), .A(n8307), .ZN(n8309) );
  NAND2_X1 U9943 ( .A1(n8309), .A2(n8380), .ZN(n8319) );
  AOI22_X1 U9944 ( .A1(n8387), .A2(n8310), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3152), .ZN(n8318) );
  AOI22_X1 U9945 ( .A1(n8392), .A2(n8312), .B1(n8311), .B2(n8372), .ZN(n8317)
         );
  INV_X1 U9946 ( .A(n8313), .ZN(n8314) );
  NAND4_X1 U9947 ( .A1(n8379), .A2(n8315), .A3(n8314), .A4(n8421), .ZN(n8316)
         );
  NAND4_X1 U9948 ( .A1(n8319), .A2(n8318), .A3(n8317), .A4(n8316), .ZN(
        P2_U3232) );
  OAI211_X1 U9949 ( .C1(n8322), .C2(n8321), .A(n8320), .B(n8380), .ZN(n8330)
         );
  INV_X1 U9950 ( .A(n8323), .ZN(n8635) );
  OR2_X1 U9951 ( .A1(n8346), .A2(n8385), .ZN(n8326) );
  NAND2_X1 U9952 ( .A1(n8406), .A2(n8324), .ZN(n8325) );
  AND2_X1 U9953 ( .A1(n8326), .A2(n8325), .ZN(n8631) );
  OAI22_X1 U9954 ( .A1(n8631), .A2(n8374), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8327), .ZN(n8328) );
  AOI21_X1 U9955 ( .B1(n8635), .B2(n8372), .A(n8328), .ZN(n8329) );
  OAI211_X1 U9956 ( .C1(n8922), .C2(n8364), .A(n8330), .B(n8329), .ZN(P2_U3235) );
  INV_X1 U9957 ( .A(n8331), .ZN(n8334) );
  NAND2_X1 U9958 ( .A1(n8372), .A2(n8332), .ZN(n8333) );
  NAND2_X1 U9959 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8432) );
  OAI211_X1 U9960 ( .C1(n8374), .C2(n8334), .A(n8333), .B(n8432), .ZN(n8339)
         );
  AOI211_X1 U9961 ( .C1(n8337), .C2(n8336), .A(n8377), .B(n8335), .ZN(n8338)
         );
  AOI211_X1 U9962 ( .C1(n8946), .C2(n8392), .A(n8339), .B(n8338), .ZN(n8340)
         );
  INV_X1 U9963 ( .A(n8340), .ZN(P2_U3236) );
  NAND2_X1 U9964 ( .A1(n8379), .A2(n8403), .ZN(n8344) );
  NAND2_X1 U9965 ( .A1(n8341), .A2(n8380), .ZN(n8343) );
  MUX2_X1 U9966 ( .A(n8344), .B(n8343), .S(n8342), .Z(n8351) );
  INV_X1 U9967 ( .A(n8345), .ZN(n8605) );
  NOR2_X1 U9968 ( .A1(n8346), .A2(n8383), .ZN(n8347) );
  AOI21_X1 U9969 ( .B1(n8402), .B2(n8360), .A(n8347), .ZN(n8600) );
  OAI22_X1 U9970 ( .A1(n8600), .A2(n8374), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8348), .ZN(n8349) );
  AOI21_X1 U9971 ( .B1(n8605), .B2(n8372), .A(n8349), .ZN(n8350) );
  OAI211_X1 U9972 ( .C1(n8917), .C2(n8364), .A(n8351), .B(n8350), .ZN(P2_U3237) );
  AOI21_X1 U9973 ( .B1(n8352), .B2(n4393), .A(n8377), .ZN(n8357) );
  NOR3_X1 U9974 ( .A1(n8354), .A2(n8358), .A3(n8353), .ZN(n8356) );
  OAI21_X1 U9975 ( .B1(n8357), .B2(n8356), .A(n8355), .ZN(n8363) );
  NOR2_X1 U9976 ( .A1(n8358), .A2(n8383), .ZN(n8359) );
  AOI21_X1 U9977 ( .B1(n8406), .B2(n8360), .A(n8359), .ZN(n8667) );
  NAND2_X1 U9978 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8489) );
  OAI21_X1 U9979 ( .B1(n8374), .B2(n8667), .A(n8489), .ZN(n8361) );
  AOI21_X1 U9980 ( .B1(n8672), .B2(n8372), .A(n8361), .ZN(n8362) );
  OAI211_X1 U9981 ( .C1(n8675), .C2(n8364), .A(n8363), .B(n8362), .ZN(P2_U3240) );
  XNOR2_X1 U9982 ( .A(n8365), .B(n8366), .ZN(n8378) );
  OR2_X1 U9983 ( .A1(n8367), .A2(n8385), .ZN(n8370) );
  OR2_X1 U9984 ( .A1(n8368), .A2(n8383), .ZN(n8369) );
  AND2_X1 U9985 ( .A1(n8370), .A2(n8369), .ZN(n8540) );
  INV_X1 U9986 ( .A(n8371), .ZN(n8544) );
  AOI22_X1 U9987 ( .A1(n8544), .A2(n8372), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n8373) );
  OAI21_X1 U9988 ( .B1(n8540), .B2(n8374), .A(n8373), .ZN(n8375) );
  AOI21_X1 U9989 ( .B1(n8543), .B2(n8392), .A(n8375), .ZN(n8376) );
  OAI21_X1 U9990 ( .B1(n8378), .B2(n8377), .A(n8376), .ZN(P2_U3242) );
  AOI22_X1 U9991 ( .A1(n8381), .A2(n8380), .B1(n8379), .B2(n8409), .ZN(n8395)
         );
  INV_X1 U9992 ( .A(n8382), .ZN(n8394) );
  INV_X1 U9993 ( .A(n8717), .ZN(n8390) );
  OAI22_X1 U9994 ( .A1(n8386), .A2(n8385), .B1(n8384), .B2(n8383), .ZN(n8714)
         );
  AOI22_X1 U9995 ( .A1(n8387), .A2(n8714), .B1(P2_REG3_REG_15__SCAN_IN), .B2(
        P2_U3152), .ZN(n8388) );
  OAI21_X1 U9996 ( .B1(n8390), .B2(n8389), .A(n8388), .ZN(n8391) );
  AOI21_X1 U9997 ( .B1(n8938), .B2(n8392), .A(n8391), .ZN(n8393) );
  OAI21_X1 U9998 ( .B1(n8395), .B2(n8394), .A(n8393), .ZN(P2_U3243) );
  MUX2_X1 U9999 ( .A(n8396), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8422), .Z(
        P2_U3582) );
  MUX2_X1 U10000 ( .A(n8397), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8422), .Z(
        P2_U3580) );
  MUX2_X1 U10001 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8398), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U10002 ( .A(n8399), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8422), .Z(
        P2_U3578) );
  MUX2_X1 U10003 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8400), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U10004 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8401), .S(P2_U3966), .Z(
        P2_U3576) );
  MUX2_X1 U10005 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8402), .S(P2_U3966), .Z(
        P2_U3575) );
  MUX2_X1 U10006 ( .A(n8403), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8422), .Z(
        P2_U3574) );
  MUX2_X1 U10007 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8404), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U10008 ( .A(n8405), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8422), .Z(
        P2_U3572) );
  MUX2_X1 U10009 ( .A(n8406), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8422), .Z(
        P2_U3571) );
  MUX2_X1 U10010 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8407), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U10011 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8408), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U10012 ( .A(n4621), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8422), .Z(
        P2_U3568) );
  MUX2_X1 U10013 ( .A(n8409), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8422), .Z(
        P2_U3567) );
  MUX2_X1 U10014 ( .A(n8410), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8422), .Z(
        P2_U3566) );
  MUX2_X1 U10015 ( .A(n8411), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8422), .Z(
        P2_U3565) );
  MUX2_X1 U10016 ( .A(n8412), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8422), .Z(
        P2_U3564) );
  MUX2_X1 U10017 ( .A(n8413), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8422), .Z(
        P2_U3563) );
  MUX2_X1 U10018 ( .A(n8414), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8422), .Z(
        P2_U3562) );
  MUX2_X1 U10019 ( .A(n8415), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8422), .Z(
        P2_U3561) );
  MUX2_X1 U10020 ( .A(n8416), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8422), .Z(
        P2_U3560) );
  MUX2_X1 U10021 ( .A(n8417), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8422), .Z(
        P2_U3559) );
  MUX2_X1 U10022 ( .A(n8418), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8422), .Z(
        P2_U3558) );
  MUX2_X1 U10023 ( .A(n8419), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8422), .Z(
        P2_U3557) );
  MUX2_X1 U10024 ( .A(n8420), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8422), .Z(
        P2_U3556) );
  MUX2_X1 U10025 ( .A(n8421), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8422), .Z(
        P2_U3555) );
  MUX2_X1 U10026 ( .A(n6318), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8422), .Z(
        P2_U3554) );
  MUX2_X1 U10027 ( .A(n6310), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8422), .Z(
        P2_U3553) );
  MUX2_X1 U10028 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8423), .S(P2_U3966), .Z(
        P2_U3552) );
  OAI21_X1 U10029 ( .B1(n8426), .B2(n8425), .A(n8424), .ZN(n8437) );
  OR3_X1 U10030 ( .A1(n8429), .A2(n8428), .A3(n8427), .ZN(n8430) );
  AOI21_X1 U10031 ( .B1(n8431), .B2(n8430), .A(n10261), .ZN(n8436) );
  NAND2_X1 U10032 ( .A1(n10258), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n8433) );
  OAI211_X1 U10033 ( .C1(n10260), .C2(n8434), .A(n8433), .B(n8432), .ZN(n8435)
         );
  AOI211_X1 U10034 ( .C1(n8437), .C2(n10256), .A(n8436), .B(n8435), .ZN(n8438)
         );
  INV_X1 U10035 ( .A(n8438), .ZN(P2_U3258) );
  OAI21_X1 U10036 ( .B1(n8441), .B2(n8440), .A(n8439), .ZN(n8442) );
  NAND2_X1 U10037 ( .A1(n8442), .A2(n10256), .ZN(n8452) );
  OAI21_X1 U10038 ( .B1(n8445), .B2(n8444), .A(n8443), .ZN(n8450) );
  NAND2_X1 U10039 ( .A1(n10258), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n8447) );
  OAI211_X1 U10040 ( .C1(n10260), .C2(n8448), .A(n8447), .B(n8446), .ZN(n8449)
         );
  AOI21_X1 U10041 ( .B1(n8450), .B2(n10255), .A(n8449), .ZN(n8451) );
  NAND2_X1 U10042 ( .A1(n8452), .A2(n8451), .ZN(P2_U3259) );
  XOR2_X1 U10043 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8453), .Z(n8461) );
  XNOR2_X1 U10044 ( .A(n8454), .B(P2_REG2_REG_15__SCAN_IN), .ZN(n8455) );
  NAND2_X1 U10045 ( .A1(n8455), .A2(n10256), .ZN(n8460) );
  AND2_X1 U10046 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8458) );
  NOR2_X1 U10047 ( .A1(n10260), .A2(n8456), .ZN(n8457) );
  AOI211_X1 U10048 ( .C1(P2_ADDR_REG_15__SCAN_IN), .C2(n10258), .A(n8458), .B(
        n8457), .ZN(n8459) );
  OAI211_X1 U10049 ( .C1(n10261), .C2(n8461), .A(n8460), .B(n8459), .ZN(
        P2_U3260) );
  AOI21_X1 U10050 ( .B1(n8464), .B2(n8463), .A(n8462), .ZN(n8474) );
  AOI211_X1 U10051 ( .C1(n8467), .C2(n8466), .A(n8465), .B(n10259), .ZN(n8468)
         );
  INV_X1 U10052 ( .A(n8468), .ZN(n8473) );
  NOR2_X1 U10053 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n4679), .ZN(n8471) );
  NOR2_X1 U10054 ( .A1(n10260), .A2(n8469), .ZN(n8470) );
  AOI211_X1 U10055 ( .C1(P2_ADDR_REG_16__SCAN_IN), .C2(n10258), .A(n8471), .B(
        n8470), .ZN(n8472) );
  OAI211_X1 U10056 ( .C1(n8474), .C2(n10261), .A(n8473), .B(n8472), .ZN(
        P2_U3261) );
  AOI211_X1 U10057 ( .C1(n4401), .C2(n8476), .A(n8475), .B(n10259), .ZN(n8485)
         );
  AND2_X1 U10058 ( .A1(P2_U3152), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8477) );
  AOI21_X1 U10059 ( .B1(n10258), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8477), .ZN(
        n8482) );
  OAI211_X1 U10060 ( .C1(n8480), .C2(n8479), .A(n10255), .B(n8478), .ZN(n8481)
         );
  OAI211_X1 U10061 ( .C1(n10260), .C2(n8483), .A(n8482), .B(n8481), .ZN(n8484)
         );
  OR2_X1 U10062 ( .A1(n8485), .A2(n8484), .ZN(P2_U3262) );
  OAI21_X1 U10063 ( .B1(n8488), .B2(n8487), .A(n8486), .ZN(n8493) );
  INV_X1 U10064 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8490) );
  OAI21_X1 U10065 ( .B1(n8491), .B2(n8490), .A(n8489), .ZN(n8492) );
  AOI21_X1 U10066 ( .B1(n10255), .B2(n8493), .A(n8492), .ZN(n8499) );
  OAI21_X1 U10067 ( .B1(n8496), .B2(n8495), .A(n8494), .ZN(n8497) );
  NAND2_X1 U10068 ( .A1(n10256), .A2(n8497), .ZN(n8498) );
  OAI211_X1 U10069 ( .C1(n10260), .C2(n8500), .A(n8499), .B(n8498), .ZN(
        P2_U3263) );
  INV_X1 U10070 ( .A(n8501), .ZN(n8502) );
  NAND2_X1 U10071 ( .A1(n8775), .A2(n8766), .ZN(n8507) );
  AOI21_X1 U10072 ( .B1(n10276), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8505), .ZN(
        n8506) );
  OAI211_X1 U10073 ( .C1(n5074), .C2(n8754), .A(n8507), .B(n8506), .ZN(
        P2_U3266) );
  NAND2_X1 U10074 ( .A1(n8508), .A2(n10284), .ZN(n8515) );
  INV_X1 U10075 ( .A(n8509), .ZN(n8513) );
  AOI22_X1 U10076 ( .A1(n8510), .A2(n10267), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n10276), .ZN(n8511) );
  OAI21_X1 U10077 ( .B1(n6587), .B2(n8754), .A(n8511), .ZN(n8512) );
  AOI21_X1 U10078 ( .B1(n8513), .B2(n8766), .A(n8512), .ZN(n8514) );
  OAI211_X1 U10079 ( .C1(n8516), .C2(n10276), .A(n8515), .B(n8514), .ZN(
        P2_U3268) );
  XNOR2_X1 U10080 ( .A(n8518), .B(n8517), .ZN(n8794) );
  NAND2_X1 U10081 ( .A1(n8519), .A2(n10290), .ZN(n8524) );
  AOI21_X1 U10082 ( .B1(n8535), .B2(n8521), .A(n8520), .ZN(n8523) );
  OAI21_X1 U10083 ( .B1(n8524), .B2(n8523), .A(n8522), .ZN(n8791) );
  AOI211_X1 U10084 ( .C1(n8793), .C2(n8526), .A(n10328), .B(n8525), .ZN(n8792)
         );
  NAND2_X1 U10085 ( .A1(n8792), .A2(n8766), .ZN(n8529) );
  AOI22_X1 U10086 ( .A1(n8527), .A2(n10267), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n10276), .ZN(n8528) );
  OAI211_X1 U10087 ( .C1(n8530), .C2(n8754), .A(n8529), .B(n8528), .ZN(n8531)
         );
  AOI21_X1 U10088 ( .B1(n8791), .B2(n8763), .A(n8531), .ZN(n8532) );
  OAI21_X1 U10089 ( .B1(n8794), .B2(n8769), .A(n8532), .ZN(P2_U3269) );
  INV_X1 U10090 ( .A(n8797), .ZN(n8549) );
  INV_X1 U10091 ( .A(n8535), .ZN(n8539) );
  AOI21_X1 U10092 ( .B1(n8554), .B2(n8537), .A(n8536), .ZN(n8538) );
  OAI21_X1 U10093 ( .B1(n8539), .B2(n8538), .A(n10290), .ZN(n8541) );
  NAND2_X1 U10094 ( .A1(n8541), .A2(n8540), .ZN(n8795) );
  AOI211_X1 U10095 ( .C1(n8543), .C2(n8558), .A(n10328), .B(n8542), .ZN(n8796)
         );
  NAND2_X1 U10096 ( .A1(n8796), .A2(n8766), .ZN(n8546) );
  AOI22_X1 U10097 ( .A1(n8544), .A2(n10267), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n10276), .ZN(n8545) );
  OAI211_X1 U10098 ( .C1(n8907), .C2(n8754), .A(n8546), .B(n8545), .ZN(n8547)
         );
  AOI21_X1 U10099 ( .B1(n8795), .B2(n8763), .A(n8547), .ZN(n8548) );
  OAI21_X1 U10100 ( .B1(n8549), .B2(n8769), .A(n8548), .ZN(P2_U3270) );
  NAND2_X1 U10101 ( .A1(n8569), .A2(n8568), .ZN(n8567) );
  NAND2_X1 U10102 ( .A1(n8567), .A2(n8551), .ZN(n8552) );
  XNOR2_X1 U10103 ( .A(n8552), .B(n8555), .ZN(n8804) );
  NAND2_X1 U10104 ( .A1(n4313), .A2(n8571), .ZN(n8570) );
  NAND2_X1 U10105 ( .A1(n8557), .A2(n8556), .ZN(n8800) );
  INV_X1 U10106 ( .A(n8574), .ZN(n8560) );
  INV_X1 U10107 ( .A(n8558), .ZN(n8559) );
  AOI211_X1 U10108 ( .C1(n8802), .C2(n8560), .A(n10328), .B(n8559), .ZN(n8801)
         );
  NAND2_X1 U10109 ( .A1(n8801), .A2(n8766), .ZN(n8563) );
  AOI22_X1 U10110 ( .A1(n8561), .A2(n10267), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n10276), .ZN(n8562) );
  OAI211_X1 U10111 ( .C1(n8564), .C2(n8754), .A(n8563), .B(n8562), .ZN(n8565)
         );
  AOI21_X1 U10112 ( .B1(n8800), .B2(n8763), .A(n8565), .ZN(n8566) );
  OAI21_X1 U10113 ( .B1(n8804), .B2(n8769), .A(n8566), .ZN(P2_U3271) );
  OAI21_X1 U10114 ( .B1(n8569), .B2(n8568), .A(n8567), .ZN(n8807) );
  INV_X1 U10115 ( .A(n8807), .ZN(n8581) );
  OAI211_X1 U10116 ( .C1(n4313), .C2(n8571), .A(n8570), .B(n10290), .ZN(n8573)
         );
  NAND2_X1 U10117 ( .A1(n8573), .A2(n8572), .ZN(n8805) );
  AOI211_X1 U10118 ( .C1(n8575), .C2(n5073), .A(n10328), .B(n8574), .ZN(n8806)
         );
  NAND2_X1 U10119 ( .A1(n8806), .A2(n8766), .ZN(n8578) );
  AOI22_X1 U10120 ( .A1(n8576), .A2(n10267), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n10276), .ZN(n8577) );
  OAI211_X1 U10121 ( .C1(n8912), .C2(n8754), .A(n8578), .B(n8577), .ZN(n8579)
         );
  AOI21_X1 U10122 ( .B1(n8805), .B2(n8763), .A(n8579), .ZN(n8580) );
  OAI21_X1 U10123 ( .B1(n8581), .B2(n8769), .A(n8580), .ZN(P2_U3272) );
  NAND2_X1 U10124 ( .A1(n8582), .A2(n8583), .ZN(n8584) );
  XNOR2_X1 U10125 ( .A(n8584), .B(n8587), .ZN(n8586) );
  AOI21_X1 U10126 ( .B1(n8586), .B2(n10290), .A(n8585), .ZN(n8815) );
  OR2_X1 U10127 ( .A1(n8588), .A2(n8587), .ZN(n8810) );
  NAND3_X1 U10128 ( .A1(n8811), .A2(n8810), .A3(n10284), .ZN(n8595) );
  AOI211_X1 U10129 ( .C1(n8813), .C2(n8602), .A(n10328), .B(n8589), .ZN(n8812)
         );
  INV_X1 U10130 ( .A(n8590), .ZN(n8591) );
  AOI22_X1 U10131 ( .A1(n8591), .A2(n10267), .B1(n10276), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n8592) );
  OAI21_X1 U10132 ( .B1(n5071), .B2(n8754), .A(n8592), .ZN(n8593) );
  AOI21_X1 U10133 ( .B1(n8812), .B2(n8766), .A(n8593), .ZN(n8594) );
  OAI211_X1 U10134 ( .C1(n10276), .C2(n8815), .A(n8595), .B(n8594), .ZN(
        P2_U3273) );
  XNOR2_X1 U10135 ( .A(n8597), .B(n8596), .ZN(n8819) );
  INV_X1 U10136 ( .A(n8819), .ZN(n8610) );
  OAI211_X1 U10137 ( .C1(n8599), .C2(n8598), .A(n8582), .B(n10290), .ZN(n8601)
         );
  NAND2_X1 U10138 ( .A1(n8601), .A2(n8600), .ZN(n8817) );
  INV_X1 U10139 ( .A(n8602), .ZN(n8603) );
  AOI211_X1 U10140 ( .C1(n8604), .C2(n8613), .A(n10328), .B(n8603), .ZN(n8818)
         );
  NAND2_X1 U10141 ( .A1(n8818), .A2(n8766), .ZN(n8607) );
  AOI22_X1 U10142 ( .A1(n10276), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8605), 
        .B2(n10267), .ZN(n8606) );
  OAI211_X1 U10143 ( .C1(n8917), .C2(n8754), .A(n8607), .B(n8606), .ZN(n8608)
         );
  AOI21_X1 U10144 ( .B1(n8817), .B2(n8763), .A(n8608), .ZN(n8609) );
  OAI21_X1 U10145 ( .B1(n8610), .B2(n8769), .A(n8609), .ZN(P2_U3274) );
  XNOR2_X1 U10146 ( .A(n8611), .B(n8619), .ZN(n8826) );
  INV_X1 U10147 ( .A(n8612), .ZN(n8615) );
  INV_X1 U10148 ( .A(n8613), .ZN(n8614) );
  AOI211_X1 U10149 ( .C1(n8823), .C2(n8615), .A(n10328), .B(n8614), .ZN(n8822)
         );
  AOI22_X1 U10150 ( .A1(n10276), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8616), 
        .B2(n10267), .ZN(n8617) );
  OAI21_X1 U10151 ( .B1(n8618), .B2(n8754), .A(n8617), .ZN(n8624) );
  XNOR2_X1 U10152 ( .A(n8620), .B(n8619), .ZN(n8622) );
  AOI21_X1 U10153 ( .B1(n8622), .B2(n10290), .A(n8621), .ZN(n8825) );
  NOR2_X1 U10154 ( .A1(n8825), .A2(n10276), .ZN(n8623) );
  AOI211_X1 U10155 ( .C1(n8822), .C2(n8766), .A(n8624), .B(n8623), .ZN(n8625)
         );
  OAI21_X1 U10156 ( .B1(n8826), .B2(n8769), .A(n8625), .ZN(P2_U3275) );
  XNOR2_X1 U10157 ( .A(n8626), .B(n8628), .ZN(n8829) );
  INV_X1 U10158 ( .A(n8829), .ZN(n8640) );
  NAND2_X1 U10159 ( .A1(n8629), .A2(n8628), .ZN(n8630) );
  NAND3_X1 U10160 ( .A1(n8627), .A2(n10290), .A3(n8630), .ZN(n8632) );
  NAND2_X1 U10161 ( .A1(n8632), .A2(n8631), .ZN(n8827) );
  INV_X1 U10162 ( .A(n8651), .ZN(n8633) );
  AOI211_X1 U10163 ( .C1(n8634), .C2(n8633), .A(n10328), .B(n8612), .ZN(n8828)
         );
  NAND2_X1 U10164 ( .A1(n8828), .A2(n8766), .ZN(n8637) );
  AOI22_X1 U10165 ( .A1(n10276), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8635), 
        .B2(n10267), .ZN(n8636) );
  OAI211_X1 U10166 ( .C1(n8922), .C2(n8754), .A(n8637), .B(n8636), .ZN(n8638)
         );
  AOI21_X1 U10167 ( .B1(n8827), .B2(n8763), .A(n8638), .ZN(n8639) );
  OAI21_X1 U10168 ( .B1(n8640), .B2(n8769), .A(n8639), .ZN(P2_U3276) );
  XNOR2_X1 U10169 ( .A(n8642), .B(n8641), .ZN(n8836) );
  NOR2_X1 U10170 ( .A1(n8662), .A2(n8643), .ZN(n8644) );
  NAND2_X1 U10171 ( .A1(n8682), .A2(n8644), .ZN(n8664) );
  NAND2_X1 U10172 ( .A1(n8664), .A2(n8645), .ZN(n8647) );
  XNOR2_X1 U10173 ( .A(n8647), .B(n8646), .ZN(n8649) );
  OAI21_X1 U10174 ( .B1(n8649), .B2(n8734), .A(n8648), .ZN(n8832) );
  OAI21_X1 U10175 ( .B1(n8671), .B2(n8650), .A(n8892), .ZN(n8652) );
  NOR2_X1 U10176 ( .A1(n8652), .A2(n8651), .ZN(n8833) );
  NAND2_X1 U10177 ( .A1(n8833), .A2(n8766), .ZN(n8657) );
  NAND2_X1 U10178 ( .A1(n10276), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8653) );
  OAI21_X1 U10179 ( .B1(n10279), .B2(n8654), .A(n8653), .ZN(n8655) );
  AOI21_X1 U10180 ( .B1(n8834), .B2(n10286), .A(n8655), .ZN(n8656) );
  NAND2_X1 U10181 ( .A1(n8657), .A2(n8656), .ZN(n8658) );
  AOI21_X1 U10182 ( .B1(n8832), .B2(n8763), .A(n8658), .ZN(n8659) );
  OAI21_X1 U10183 ( .B1(n8836), .B2(n8769), .A(n8659), .ZN(P2_U3277) );
  XNOR2_X1 U10184 ( .A(n8660), .B(n8662), .ZN(n8839) );
  INV_X1 U10185 ( .A(n8839), .ZN(n8678) );
  NAND2_X1 U10186 ( .A1(n8682), .A2(n8661), .ZN(n8663) );
  NAND2_X1 U10187 ( .A1(n8663), .A2(n8662), .ZN(n8665) );
  NAND2_X1 U10188 ( .A1(n8665), .A2(n8664), .ZN(n8666) );
  NAND2_X1 U10189 ( .A1(n8666), .A2(n10290), .ZN(n8668) );
  NAND2_X1 U10190 ( .A1(n8668), .A2(n8667), .ZN(n8838) );
  NAND2_X1 U10191 ( .A1(n8688), .A2(n8926), .ZN(n8669) );
  NAND2_X1 U10192 ( .A1(n8669), .A2(n8892), .ZN(n8670) );
  NOR2_X1 U10193 ( .A1(n8671), .A2(n8670), .ZN(n8837) );
  NAND2_X1 U10194 ( .A1(n8837), .A2(n8766), .ZN(n8674) );
  AOI22_X1 U10195 ( .A1(n10276), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8672), 
        .B2(n10267), .ZN(n8673) );
  OAI211_X1 U10196 ( .C1(n8675), .C2(n8754), .A(n8674), .B(n8673), .ZN(n8676)
         );
  AOI21_X1 U10197 ( .B1(n8838), .B2(n8763), .A(n8676), .ZN(n8677) );
  OAI21_X1 U10198 ( .B1(n8678), .B2(n8769), .A(n8677), .ZN(P2_U3278) );
  AOI21_X1 U10199 ( .B1(n8680), .B2(n8679), .A(n8734), .ZN(n8683) );
  AOI21_X1 U10200 ( .B1(n8683), .B2(n8682), .A(n8681), .ZN(n8846) );
  NAND2_X1 U10201 ( .A1(n8686), .A2(n8685), .ZN(n8687) );
  NAND2_X1 U10202 ( .A1(n8684), .A2(n8687), .ZN(n8844) );
  AOI21_X1 U10203 ( .B1(n8703), .B2(n8930), .A(n10328), .ZN(n8689) );
  NAND2_X1 U10204 ( .A1(n8689), .A2(n8688), .ZN(n8845) );
  AOI22_X1 U10205 ( .A1(n10276), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8690), 
        .B2(n10267), .ZN(n8692) );
  NAND2_X1 U10206 ( .A1(n8930), .A2(n10286), .ZN(n8691) );
  OAI211_X1 U10207 ( .C1(n8845), .C2(n10281), .A(n8692), .B(n8691), .ZN(n8693)
         );
  AOI21_X1 U10208 ( .B1(n8844), .B2(n10284), .A(n8693), .ZN(n8694) );
  OAI21_X1 U10209 ( .B1(n10276), .B2(n8846), .A(n8694), .ZN(P2_U3279) );
  XNOR2_X1 U10210 ( .A(n8696), .B(n8119), .ZN(n8698) );
  AOI21_X1 U10211 ( .B1(n8698), .B2(n10290), .A(n8697), .ZN(n8851) );
  NAND2_X1 U10212 ( .A1(n8699), .A2(n8700), .ZN(n8701) );
  NAND2_X1 U10213 ( .A1(n8702), .A2(n8701), .ZN(n8852) );
  INV_X1 U10214 ( .A(n8852), .ZN(n8710) );
  AOI21_X1 U10215 ( .B1(n8724), .B2(n8933), .A(n10328), .ZN(n8704) );
  NAND2_X1 U10216 ( .A1(n8704), .A2(n8703), .ZN(n8850) );
  NAND2_X1 U10217 ( .A1(n10276), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8705) );
  OAI21_X1 U10218 ( .B1(n10279), .B2(n8706), .A(n8705), .ZN(n8707) );
  AOI21_X1 U10219 ( .B1(n8933), .B2(n10286), .A(n8707), .ZN(n8708) );
  OAI21_X1 U10220 ( .B1(n8850), .B2(n10281), .A(n8708), .ZN(n8709) );
  AOI21_X1 U10221 ( .B1(n8710), .B2(n10284), .A(n8709), .ZN(n8711) );
  OAI21_X1 U10222 ( .B1(n10276), .B2(n8851), .A(n8711), .ZN(P2_U3280) );
  INV_X1 U10223 ( .A(n8721), .ZN(n8713) );
  XNOR2_X1 U10224 ( .A(n8712), .B(n8713), .ZN(n8715) );
  AOI21_X1 U10225 ( .B1(n8715), .B2(n10290), .A(n8714), .ZN(n8858) );
  INV_X1 U10226 ( .A(n8858), .ZN(n8716) );
  AOI21_X1 U10227 ( .B1(n8717), .B2(n10267), .A(n8716), .ZN(n8729) );
  NAND2_X1 U10228 ( .A1(n8719), .A2(n8718), .ZN(n8730) );
  OAI211_X1 U10229 ( .C1(n8730), .C2(n6441), .A(n8721), .B(n5205), .ZN(n8723)
         );
  NAND2_X1 U10230 ( .A1(n8723), .A2(n8722), .ZN(n8855) );
  OAI211_X1 U10231 ( .C1(n8737), .C2(n8725), .A(n8892), .B(n8724), .ZN(n8856)
         );
  AOI22_X1 U10232 ( .A1(n8938), .A2(n10286), .B1(P2_REG2_REG_15__SCAN_IN), 
        .B2(n10276), .ZN(n8726) );
  OAI21_X1 U10233 ( .B1(n8856), .B2(n10281), .A(n8726), .ZN(n8727) );
  AOI21_X1 U10234 ( .B1(n8855), .B2(n10284), .A(n8727), .ZN(n8728) );
  OAI21_X1 U10235 ( .B1(n8729), .B2(n10276), .A(n8728), .ZN(P2_U3281) );
  XNOR2_X1 U10236 ( .A(n8730), .B(n6441), .ZN(n8863) );
  INV_X1 U10237 ( .A(n8863), .ZN(n8745) );
  XNOR2_X1 U10238 ( .A(n8731), .B(n8732), .ZN(n8735) );
  OAI21_X1 U10239 ( .B1(n8735), .B2(n8734), .A(n8733), .ZN(n8861) );
  INV_X1 U10240 ( .A(n8736), .ZN(n8738) );
  AOI211_X1 U10241 ( .C1(n8739), .C2(n8738), .A(n10328), .B(n8737), .ZN(n8862)
         );
  NAND2_X1 U10242 ( .A1(n8862), .A2(n8766), .ZN(n8742) );
  AOI22_X1 U10243 ( .A1(n10276), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8740), 
        .B2(n10267), .ZN(n8741) );
  OAI211_X1 U10244 ( .C1(n8943), .C2(n8754), .A(n8742), .B(n8741), .ZN(n8743)
         );
  AOI21_X1 U10245 ( .B1(n8861), .B2(n8763), .A(n8743), .ZN(n8744) );
  OAI21_X1 U10246 ( .B1(n8745), .B2(n8769), .A(n8744), .ZN(P2_U3282) );
  XOR2_X1 U10247 ( .A(n8746), .B(n8757), .Z(n8882) );
  INV_X1 U10248 ( .A(n8882), .ZN(n8768) );
  INV_X1 U10249 ( .A(n8747), .ZN(n8750) );
  INV_X1 U10250 ( .A(n8748), .ZN(n8749) );
  AOI211_X1 U10251 ( .C1(n8751), .C2(n8750), .A(n10328), .B(n8749), .ZN(n8881)
         );
  INV_X1 U10252 ( .A(n8752), .ZN(n8753) );
  OAI22_X1 U10253 ( .A1(n8754), .A2(n8957), .B1(n8753), .B2(n10279), .ZN(n8765) );
  NAND2_X1 U10254 ( .A1(n8756), .A2(n8755), .ZN(n8758) );
  NAND2_X1 U10255 ( .A1(n8758), .A2(n8757), .ZN(n8759) );
  OAI211_X1 U10256 ( .C1(n8760), .C2(n5130), .A(n8759), .B(n10290), .ZN(n8762)
         );
  NAND2_X1 U10257 ( .A1(n8762), .A2(n8761), .ZN(n8880) );
  MUX2_X1 U10258 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n8880), .S(n8763), .Z(n8764) );
  AOI211_X1 U10259 ( .C1(n8881), .C2(n8766), .A(n8765), .B(n8764), .ZN(n8767)
         );
  OAI21_X1 U10260 ( .B1(n8769), .B2(n8768), .A(n8767), .ZN(P2_U3285) );
  INV_X1 U10261 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8771) );
  OAI21_X1 U10262 ( .B1(n8900), .B2(n8885), .A(n8772), .ZN(P2_U3551) );
  INV_X1 U10263 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8776) );
  INV_X1 U10264 ( .A(n8773), .ZN(n8774) );
  NOR2_X1 U10265 ( .A1(n8775), .A2(n8774), .ZN(n8901) );
  MUX2_X1 U10266 ( .A(n8776), .B(n8901), .S(n10352), .Z(n8777) );
  OAI21_X1 U10267 ( .B1(n5074), .B2(n8885), .A(n8777), .ZN(P2_U3550) );
  NAND2_X1 U10268 ( .A1(n4740), .A2(n10331), .ZN(n8778) );
  NOR3_X1 U10269 ( .A1(n4740), .A2(n8868), .A3(n8779), .ZN(n8787) );
  OR2_X1 U10270 ( .A1(n8780), .A2(n8868), .ZN(n8784) );
  NAND2_X1 U10271 ( .A1(n8781), .A2(n10338), .ZN(n8783) );
  OAI211_X1 U10272 ( .C1(n8785), .C2(n8784), .A(n8783), .B(n8782), .ZN(n8786)
         );
  AOI21_X1 U10273 ( .B1(n8788), .B2(n8787), .A(n8786), .ZN(n8790) );
  MUX2_X1 U10274 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8903), .S(n10352), .Z(
        P2_U3549) );
  MUX2_X1 U10275 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8904), .S(n10352), .Z(
        P2_U3547) );
  INV_X1 U10276 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8798) );
  OAI21_X1 U10277 ( .B1(n8907), .B2(n8885), .A(n8799), .ZN(P2_U3546) );
  AOI211_X1 U10278 ( .C1(n10338), .C2(n8802), .A(n8801), .B(n8800), .ZN(n8803)
         );
  OAI21_X1 U10279 ( .B1(n8804), .B2(n8868), .A(n8803), .ZN(n8908) );
  MUX2_X1 U10280 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8908), .S(n10352), .Z(
        P2_U3545) );
  INV_X1 U10281 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8808) );
  AOI211_X1 U10282 ( .C1(n8807), .C2(n10331), .A(n8806), .B(n8805), .ZN(n8909)
         );
  MUX2_X1 U10283 ( .A(n8808), .B(n8909), .S(n10352), .Z(n8809) );
  OAI21_X1 U10284 ( .B1(n8912), .B2(n8885), .A(n8809), .ZN(P2_U3544) );
  NAND3_X1 U10285 ( .A1(n8811), .A2(n8810), .A3(n10331), .ZN(n8816) );
  AOI21_X1 U10286 ( .B1(n10338), .B2(n8813), .A(n8812), .ZN(n8814) );
  NAND3_X1 U10287 ( .A1(n8816), .A2(n8815), .A3(n8814), .ZN(n8913) );
  MUX2_X1 U10288 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8913), .S(n10352), .Z(
        P2_U3543) );
  INV_X1 U10289 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8820) );
  AOI211_X1 U10290 ( .C1(n8819), .C2(n10331), .A(n8818), .B(n8817), .ZN(n8914)
         );
  MUX2_X1 U10291 ( .A(n8820), .B(n8914), .S(n10352), .Z(n8821) );
  OAI21_X1 U10292 ( .B1(n8917), .B2(n8885), .A(n8821), .ZN(P2_U3542) );
  AOI21_X1 U10293 ( .B1(n10338), .B2(n8823), .A(n8822), .ZN(n8824) );
  OAI211_X1 U10294 ( .C1(n8826), .C2(n8868), .A(n8825), .B(n8824), .ZN(n8918)
         );
  MUX2_X1 U10295 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8918), .S(n10352), .Z(
        P2_U3541) );
  INV_X1 U10296 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8830) );
  AOI211_X1 U10297 ( .C1(n8829), .C2(n10331), .A(n8828), .B(n8827), .ZN(n8919)
         );
  MUX2_X1 U10298 ( .A(n8830), .B(n8919), .S(n10352), .Z(n8831) );
  OAI21_X1 U10299 ( .B1(n8922), .B2(n8885), .A(n8831), .ZN(P2_U3540) );
  AOI211_X1 U10300 ( .C1(n10338), .C2(n8834), .A(n8833), .B(n8832), .ZN(n8835)
         );
  OAI21_X1 U10301 ( .B1(n8868), .B2(n8836), .A(n8835), .ZN(n8923) );
  MUX2_X1 U10302 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8923), .S(n10352), .Z(
        P2_U3539) );
  NOR2_X1 U10303 ( .A1(n8838), .A2(n8837), .ZN(n8841) );
  NAND2_X1 U10304 ( .A1(n8839), .A2(n10331), .ZN(n8840) );
  NAND2_X1 U10305 ( .A1(n8841), .A2(n8840), .ZN(n8924) );
  MUX2_X1 U10306 ( .A(n8924), .B(P2_REG1_REG_18__SCAN_IN), .S(n4653), .Z(n8842) );
  AOI21_X1 U10307 ( .B1(n8873), .B2(n8926), .A(n8842), .ZN(n8843) );
  INV_X1 U10308 ( .A(n8843), .ZN(P2_U3538) );
  NAND2_X1 U10309 ( .A1(n8844), .A2(n10331), .ZN(n8847) );
  NAND3_X1 U10310 ( .A1(n8847), .A2(n8846), .A3(n8845), .ZN(n8928) );
  MUX2_X1 U10311 ( .A(n8928), .B(P2_REG1_REG_17__SCAN_IN), .S(n4653), .Z(n8848) );
  AOI21_X1 U10312 ( .B1(n8873), .B2(n8930), .A(n8848), .ZN(n8849) );
  INV_X1 U10313 ( .A(n8849), .ZN(P2_U3537) );
  OAI211_X1 U10314 ( .C1(n8852), .C2(n8868), .A(n8851), .B(n8850), .ZN(n8932)
         );
  MUX2_X1 U10315 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8932), .S(n10352), .Z(
        n8854) );
  AND2_X1 U10316 ( .A1(n8933), .A2(n8873), .ZN(n8853) );
  OR2_X1 U10317 ( .A1(n8854), .A2(n8853), .ZN(P2_U3536) );
  NAND2_X1 U10318 ( .A1(n8855), .A2(n10331), .ZN(n8857) );
  NAND3_X1 U10319 ( .A1(n8858), .A2(n8857), .A3(n8856), .ZN(n8936) );
  MUX2_X1 U10320 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8936), .S(n10352), .Z(
        n8859) );
  AOI21_X1 U10321 ( .B1(n8873), .B2(n8938), .A(n8859), .ZN(n8860) );
  INV_X1 U10322 ( .A(n8860), .ZN(P2_U3535) );
  AOI211_X1 U10323 ( .C1(n10331), .C2(n8863), .A(n8862), .B(n8861), .ZN(n8940)
         );
  MUX2_X1 U10324 ( .A(n8864), .B(n8940), .S(n10352), .Z(n8865) );
  OAI21_X1 U10325 ( .B1(n8943), .B2(n8885), .A(n8865), .ZN(P2_U3534) );
  NOR2_X1 U10326 ( .A1(n8867), .A2(n8866), .ZN(n8871) );
  OR2_X1 U10327 ( .A1(n8869), .A2(n8868), .ZN(n8870) );
  NAND2_X1 U10328 ( .A1(n8871), .A2(n8870), .ZN(n8944) );
  MUX2_X1 U10329 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n8944), .S(n10352), .Z(
        n8872) );
  AOI21_X1 U10330 ( .B1(n8873), .B2(n8946), .A(n8872), .ZN(n8874) );
  INV_X1 U10331 ( .A(n8874), .ZN(P2_U3533) );
  INV_X1 U10332 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8878) );
  AOI211_X1 U10333 ( .C1(n8877), .C2(n10331), .A(n8876), .B(n8875), .ZN(n8949)
         );
  MUX2_X1 U10334 ( .A(n8878), .B(n8949), .S(n10352), .Z(n8879) );
  OAI21_X1 U10335 ( .B1(n8952), .B2(n8885), .A(n8879), .ZN(P2_U3532) );
  AOI211_X1 U10336 ( .C1(n8882), .C2(n10331), .A(n8881), .B(n8880), .ZN(n8953)
         );
  MUX2_X1 U10337 ( .A(n8883), .B(n8953), .S(n10352), .Z(n8884) );
  OAI21_X1 U10338 ( .B1(n8957), .B2(n8885), .A(n8884), .ZN(P2_U3531) );
  AOI21_X1 U10339 ( .B1(n10338), .B2(n8887), .A(n8886), .ZN(n8888) );
  OAI211_X1 U10340 ( .C1(n10342), .C2(n8890), .A(n8889), .B(n8888), .ZN(n8958)
         );
  MUX2_X1 U10341 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n8958), .S(n10352), .Z(
        P2_U3530) );
  AOI22_X1 U10342 ( .A1(n8893), .A2(n8892), .B1(n10338), .B2(n8891), .ZN(n8894) );
  OAI211_X1 U10343 ( .C1(n8896), .C2(n10342), .A(n8895), .B(n8894), .ZN(n8959)
         );
  MUX2_X1 U10344 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n8959), .S(n10352), .Z(
        P2_U3529) );
  OAI21_X1 U10345 ( .B1(n8900), .B2(n8956), .A(n8899), .ZN(P2_U3519) );
  INV_X1 U10346 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9923) );
  MUX2_X1 U10347 ( .A(n9923), .B(n8901), .S(n10345), .Z(n8902) );
  OAI21_X1 U10348 ( .B1(n5074), .B2(n8956), .A(n8902), .ZN(P2_U3518) );
  MUX2_X1 U10349 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8903), .S(n10345), .Z(
        P2_U3517) );
  MUX2_X1 U10350 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8904), .S(n10345), .Z(
        P2_U3515) );
  MUX2_X1 U10351 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8908), .S(n10345), .Z(
        P2_U3513) );
  MUX2_X1 U10352 ( .A(n8910), .B(n8909), .S(n10345), .Z(n8911) );
  OAI21_X1 U10353 ( .B1(n8912), .B2(n8956), .A(n8911), .ZN(P2_U3512) );
  MUX2_X1 U10354 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8913), .S(n10345), .Z(
        P2_U3511) );
  MUX2_X1 U10355 ( .A(n8915), .B(n8914), .S(n10345), .Z(n8916) );
  OAI21_X1 U10356 ( .B1(n8917), .B2(n8956), .A(n8916), .ZN(P2_U3510) );
  MUX2_X1 U10357 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8918), .S(n10345), .Z(
        P2_U3509) );
  MUX2_X1 U10358 ( .A(n8920), .B(n8919), .S(n10345), .Z(n8921) );
  OAI21_X1 U10359 ( .B1(n8922), .B2(n8956), .A(n8921), .ZN(P2_U3508) );
  MUX2_X1 U10360 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8923), .S(n10345), .Z(
        P2_U3507) );
  MUX2_X1 U10361 ( .A(n8924), .B(P2_REG0_REG_18__SCAN_IN), .S(n4655), .Z(n8925) );
  AOI21_X1 U10362 ( .B1(n8947), .B2(n8926), .A(n8925), .ZN(n8927) );
  INV_X1 U10363 ( .A(n8927), .ZN(P2_U3505) );
  MUX2_X1 U10364 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8928), .S(n10345), .Z(
        n8929) );
  AOI21_X1 U10365 ( .B1(n8947), .B2(n8930), .A(n8929), .ZN(n8931) );
  INV_X1 U10366 ( .A(n8931), .ZN(P2_U3502) );
  MUX2_X1 U10367 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8932), .S(n10345), .Z(
        n8935) );
  AND2_X1 U10368 ( .A1(n8933), .A2(n8947), .ZN(n8934) );
  OR2_X1 U10369 ( .A1(n8935), .A2(n8934), .ZN(P2_U3499) );
  MUX2_X1 U10370 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8936), .S(n10345), .Z(
        n8937) );
  AOI21_X1 U10371 ( .B1(n8947), .B2(n8938), .A(n8937), .ZN(n8939) );
  INV_X1 U10372 ( .A(n8939), .ZN(P2_U3496) );
  INV_X1 U10373 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8941) );
  MUX2_X1 U10374 ( .A(n8941), .B(n8940), .S(n10345), .Z(n8942) );
  OAI21_X1 U10375 ( .B1(n8943), .B2(n8956), .A(n8942), .ZN(P2_U3493) );
  MUX2_X1 U10376 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n8944), .S(n10345), .Z(
        n8945) );
  AOI21_X1 U10377 ( .B1(n8947), .B2(n8946), .A(n8945), .ZN(n8948) );
  INV_X1 U10378 ( .A(n8948), .ZN(P2_U3490) );
  INV_X1 U10379 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n8950) );
  MUX2_X1 U10380 ( .A(n8950), .B(n8949), .S(n10345), .Z(n8951) );
  OAI21_X1 U10381 ( .B1(n8952), .B2(n8956), .A(n8951), .ZN(P2_U3487) );
  INV_X1 U10382 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n8954) );
  MUX2_X1 U10383 ( .A(n8954), .B(n8953), .S(n10345), .Z(n8955) );
  OAI21_X1 U10384 ( .B1(n8957), .B2(n8956), .A(n8955), .ZN(P2_U3484) );
  MUX2_X1 U10385 ( .A(P2_REG0_REG_10__SCAN_IN), .B(n8958), .S(n10345), .Z(
        P2_U3481) );
  MUX2_X1 U10386 ( .A(P2_REG0_REG_9__SCAN_IN), .B(n8959), .S(n10345), .Z(
        P2_U3478) );
  NAND2_X1 U10387 ( .A1(n10080), .A2(n8960), .ZN(n8963) );
  NAND4_X1 U10388 ( .A1(n4310), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .A4(n8961), .ZN(n8962) );
  OAI211_X1 U10389 ( .C1(n8964), .C2(n8974), .A(n8963), .B(n8962), .ZN(
        P2_U3327) );
  INV_X1 U10390 ( .A(n8965), .ZN(n10086) );
  OAI222_X1 U10391 ( .A1(n8977), .A2(n10086), .B1(P2_U3152), .B2(n8967), .C1(
        n8966), .C2(n8974), .ZN(P2_U3329) );
  OAI222_X1 U10392 ( .A1(n8974), .A2(n8970), .B1(P2_U3152), .B2(n8969), .C1(
        n8977), .C2(n8968), .ZN(P2_U3330) );
  INV_X1 U10393 ( .A(n10090), .ZN(n8972) );
  OAI222_X1 U10394 ( .A1(n8974), .A2(n8973), .B1(n8977), .B2(n8972), .C1(n8971), .C2(P2_U3152), .ZN(P2_U3331) );
  OAI222_X1 U10395 ( .A1(n8978), .A2(P2_U3152), .B1(n8977), .B2(n8976), .C1(
        n8975), .C2(n8974), .ZN(P2_U3332) );
  MUX2_X1 U10396 ( .A(n8979), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XOR2_X1 U10397 ( .A(n8981), .B(n8980), .Z(n8982) );
  XNOR2_X1 U10398 ( .A(n8983), .B(n8982), .ZN(n8988) );
  OAI22_X1 U10399 ( .A1(n9553), .A2(n9146), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9896), .ZN(n8984) );
  AOI21_X1 U10400 ( .B1(n9590), .B2(n9150), .A(n8984), .ZN(n8985) );
  OAI21_X1 U10401 ( .B1(n9550), .B2(n9148), .A(n8985), .ZN(n8986) );
  AOI21_X1 U10402 ( .B1(n9819), .B2(n9138), .A(n8986), .ZN(n8987) );
  OAI21_X1 U10403 ( .B1(n8988), .B2(n9140), .A(n8987), .ZN(P1_U3212) );
  AOI21_X1 U10404 ( .B1(n8992), .B2(n8990), .A(n8989), .ZN(n8991) );
  AOI211_X1 U10405 ( .C1(n8993), .C2(n8992), .A(n9140), .B(n8991), .ZN(n8994)
         );
  INV_X1 U10406 ( .A(n8994), .ZN(n8997) );
  AND2_X1 U10407 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9466) );
  OAI22_X1 U10408 ( .A1(n9148), .A2(n9769), .B1(n9146), .B2(n9775), .ZN(n8995)
         );
  AOI211_X1 U10409 ( .C1(n9150), .C2(n9450), .A(n9466), .B(n8995), .ZN(n8996)
         );
  OAI211_X1 U10410 ( .C1(n9778), .C2(n9153), .A(n8997), .B(n8996), .ZN(
        P1_U3213) );
  NAND2_X1 U10411 ( .A1(n4359), .A2(n9028), .ZN(n9000) );
  XNOR2_X1 U10412 ( .A(n9000), .B(n9029), .ZN(n9005) );
  OAI22_X1 U10413 ( .A1(n9617), .A2(n9148), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9001), .ZN(n9003) );
  OAI22_X1 U10414 ( .A1(n9648), .A2(n9113), .B1(n9146), .B2(n9612), .ZN(n9002)
         );
  AOI211_X1 U10415 ( .C1(n9980), .C2(n9138), .A(n9003), .B(n9002), .ZN(n9004)
         );
  OAI21_X1 U10416 ( .B1(n9005), .B2(n9140), .A(n9004), .ZN(P1_U3214) );
  INV_X1 U10417 ( .A(n9110), .ZN(n9007) );
  NAND2_X1 U10418 ( .A1(n4335), .A2(n9006), .ZN(n9108) );
  NOR2_X1 U10419 ( .A1(n4335), .A2(n9006), .ZN(n9107) );
  AOI21_X1 U10420 ( .B1(n9007), .B2(n9108), .A(n9107), .ZN(n9011) );
  NAND2_X1 U10421 ( .A1(n9009), .A2(n9008), .ZN(n9010) );
  XNOR2_X1 U10422 ( .A(n9011), .B(n9010), .ZN(n9016) );
  NOR2_X1 U10423 ( .A1(n9934), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9521) );
  INV_X1 U10424 ( .A(n9012), .ZN(n9680) );
  OAI22_X1 U10425 ( .A1(n9647), .A2(n9148), .B1(n9146), .B2(n9680), .ZN(n9013)
         );
  AOI211_X1 U10426 ( .C1(n9150), .C2(n9714), .A(n9521), .B(n9013), .ZN(n9015)
         );
  NAND2_X1 U10427 ( .A1(n9999), .A2(n9138), .ZN(n9014) );
  OAI211_X1 U10428 ( .C1(n9016), .C2(n9140), .A(n9015), .B(n9014), .ZN(
        P1_U3217) );
  INV_X1 U10429 ( .A(n9017), .ZN(n9018) );
  NOR2_X1 U10430 ( .A1(n9019), .A2(n9018), .ZN(n9020) );
  XNOR2_X1 U10431 ( .A(n9021), .B(n9020), .ZN(n9027) );
  OAI22_X1 U10432 ( .A1(n9113), .A2(n9647), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9022), .ZN(n9025) );
  INV_X1 U10433 ( .A(n9652), .ZN(n9023) );
  OAI22_X1 U10434 ( .A1(n9648), .A2(n9148), .B1(n9146), .B2(n9023), .ZN(n9024)
         );
  AOI211_X1 U10435 ( .C1(n9991), .C2(n9138), .A(n9025), .B(n9024), .ZN(n9026)
         );
  OAI21_X1 U10436 ( .B1(n9027), .B2(n9140), .A(n9026), .ZN(P1_U3221) );
  NAND2_X1 U10437 ( .A1(n9031), .A2(n9030), .ZN(n9059) );
  OAI22_X1 U10438 ( .A1(n9617), .A2(n9113), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9034), .ZN(n9036) );
  NOR2_X1 U10439 ( .A1(n9549), .A2(n9148), .ZN(n9035) );
  AOI211_X1 U10440 ( .C1(n9584), .C2(n9134), .A(n9036), .B(n9035), .ZN(n9037)
         );
  XNOR2_X1 U10441 ( .A(n9045), .B(n9044), .ZN(n9039) );
  XNOR2_X1 U10442 ( .A(n9038), .B(n9039), .ZN(n9043) );
  NAND2_X1 U10443 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n10169)
         );
  OAI21_X1 U10444 ( .B1(n9113), .B2(n9769), .A(n10169), .ZN(n9041) );
  OAI22_X1 U10445 ( .A1(n9148), .A2(n9722), .B1(n9146), .B2(n9719), .ZN(n9040)
         );
  AOI211_X1 U10446 ( .C1(n9734), .C2(n9138), .A(n9041), .B(n9040), .ZN(n9042)
         );
  OAI21_X1 U10447 ( .B1(n9043), .B2(n9140), .A(n9042), .ZN(P1_U3224) );
  INV_X1 U10448 ( .A(n9038), .ZN(n9046) );
  OAI21_X1 U10449 ( .B1(n9046), .B2(n9045), .A(n9044), .ZN(n9047) );
  OAI21_X1 U10450 ( .B1(n9038), .B2(n9048), .A(n9047), .ZN(n9052) );
  XNOR2_X1 U10451 ( .A(n9050), .B(n9049), .ZN(n9051) );
  XNOR2_X1 U10452 ( .A(n9052), .B(n9051), .ZN(n9057) );
  AOI22_X1 U10453 ( .A1(n9150), .A2(n9750), .B1(n9134), .B2(n9709), .ZN(n9053)
         );
  NAND2_X1 U10454 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10181)
         );
  OAI211_X1 U10455 ( .C1(n9054), .C2(n9148), .A(n9053), .B(n10181), .ZN(n9055)
         );
  AOI21_X1 U10456 ( .B1(n10010), .B2(n9138), .A(n9055), .ZN(n9056) );
  OAI21_X1 U10457 ( .B1(n9057), .B2(n9140), .A(n9056), .ZN(P1_U3226) );
  NOR2_X1 U10458 ( .A1(n9567), .A2(n9148), .ZN(n9063) );
  AOI22_X1 U10459 ( .A1(n9629), .A2(n9150), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n9061) );
  OAI21_X1 U10460 ( .B1(n9146), .B2(n9602), .A(n9061), .ZN(n9062) );
  AOI211_X1 U10461 ( .C1(n9977), .C2(n9138), .A(n9063), .B(n9062), .ZN(n9064)
         );
  NAND2_X1 U10462 ( .A1(n9066), .A2(n9065), .ZN(n9068) );
  XOR2_X1 U10463 ( .A(n9068), .B(n9067), .Z(n9069) );
  NAND2_X1 U10464 ( .A1(n9069), .A2(n9145), .ZN(n9076) );
  AOI22_X1 U10465 ( .A1(n9125), .A2(n9457), .B1(n9150), .B2(n9459), .ZN(n9075)
         );
  AOI21_X1 U10466 ( .B1(n9138), .B2(n9071), .A(n9070), .ZN(n9074) );
  NAND2_X1 U10467 ( .A1(n9134), .A2(n9072), .ZN(n9073) );
  NAND4_X1 U10468 ( .A1(n9076), .A2(n9075), .A3(n9074), .A4(n9073), .ZN(
        P1_U3228) );
  INV_X1 U10469 ( .A(n9077), .ZN(n9079) );
  NAND2_X1 U10470 ( .A1(n9079), .A2(n9078), .ZN(n9080) );
  XNOR2_X1 U10471 ( .A(n9081), .B(n9080), .ZN(n9086) );
  OAI22_X1 U10472 ( .A1(n9113), .A2(n9112), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9082), .ZN(n9084) );
  OAI22_X1 U10473 ( .A1(n9220), .A2(n9148), .B1(n9146), .B2(n9660), .ZN(n9083)
         );
  AOI211_X1 U10474 ( .C1(n9994), .C2(n9138), .A(n9084), .B(n9083), .ZN(n9085)
         );
  OAI21_X1 U10475 ( .B1(n9086), .B2(n9140), .A(n9085), .ZN(P1_U3231) );
  XNOR2_X1 U10476 ( .A(n9088), .B(n9087), .ZN(n9089) );
  XNOR2_X1 U10477 ( .A(n9090), .B(n9089), .ZN(n9097) );
  OAI22_X1 U10478 ( .A1(n9220), .A2(n9113), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9091), .ZN(n9095) );
  INV_X1 U10479 ( .A(n9633), .ZN(n9092) );
  OAI22_X1 U10480 ( .A1(n9093), .A2(n9148), .B1(n9146), .B2(n9092), .ZN(n9094)
         );
  AOI211_X1 U10481 ( .C1(n9984), .C2(n9138), .A(n9095), .B(n9094), .ZN(n9096)
         );
  OAI21_X1 U10482 ( .B1(n9097), .B2(n9140), .A(n9096), .ZN(P1_U3233) );
  OAI21_X1 U10483 ( .B1(n9100), .B2(n9099), .A(n9098), .ZN(n9101) );
  NAND2_X1 U10484 ( .A1(n9101), .A2(n9145), .ZN(n9106) );
  AOI22_X1 U10485 ( .A1(n9103), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n9138), .B2(
        n9102), .ZN(n9105) );
  AOI22_X1 U10486 ( .A1(n9125), .A2(n9459), .B1(n9150), .B2(n7290), .ZN(n9104)
         );
  NAND3_X1 U10487 ( .A1(n9106), .A2(n9105), .A3(n9104), .ZN(P1_U3235) );
  INV_X1 U10488 ( .A(n9107), .ZN(n9109) );
  NAND2_X1 U10489 ( .A1(n9109), .A2(n9108), .ZN(n9111) );
  XNOR2_X1 U10490 ( .A(n9111), .B(n9110), .ZN(n9117) );
  NAND2_X1 U10491 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9492) );
  OAI21_X1 U10492 ( .B1(n9112), .B2(n9148), .A(n9492), .ZN(n9115) );
  OAI22_X1 U10493 ( .A1(n9113), .A2(n9722), .B1(n9146), .B2(n9701), .ZN(n9114)
         );
  AOI211_X1 U10494 ( .C1(n10004), .C2(n9138), .A(n9115), .B(n9114), .ZN(n9116)
         );
  OAI21_X1 U10495 ( .B1(n9117), .B2(n9140), .A(n9116), .ZN(P1_U3236) );
  XNOR2_X1 U10496 ( .A(n9119), .B(n9118), .ZN(n9120) );
  XNOR2_X1 U10497 ( .A(n4753), .B(n9120), .ZN(n9122) );
  NAND2_X1 U10498 ( .A1(n9122), .A2(n9145), .ZN(n9130) );
  AOI22_X1 U10499 ( .A1(n9150), .A2(n9457), .B1(n9123), .B2(n9138), .ZN(n9129)
         );
  AOI21_X1 U10500 ( .B1(n9125), .B2(n9455), .A(n9124), .ZN(n9128) );
  NAND2_X1 U10501 ( .A1(n9134), .A2(n9126), .ZN(n9127) );
  NAND4_X1 U10502 ( .A1(n9130), .A2(n9129), .A3(n9128), .A4(n9127), .ZN(
        P1_U3237) );
  NAND2_X1 U10503 ( .A1(n4349), .A2(n9131), .ZN(n9132) );
  XNOR2_X1 U10504 ( .A(n9133), .B(n9132), .ZN(n9141) );
  AOI22_X1 U10505 ( .A1(n9574), .A2(n9134), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9136) );
  NAND2_X1 U10506 ( .A1(n9598), .A2(n9150), .ZN(n9135) );
  OAI211_X1 U10507 ( .C1(n9566), .C2(n9148), .A(n9136), .B(n9135), .ZN(n9137)
         );
  AOI21_X1 U10508 ( .B1(n9826), .B2(n9138), .A(n9137), .ZN(n9139) );
  OAI21_X1 U10509 ( .B1(n9141), .B2(n9140), .A(n9139), .ZN(P1_U3238) );
  OAI21_X1 U10510 ( .B1(n9143), .B2(n4295), .A(n9142), .ZN(n9144) );
  OAI211_X1 U10511 ( .C1(n4361), .C2(n4295), .A(n9145), .B(n9144), .ZN(n9152)
         );
  AND2_X1 U10512 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10162) );
  OAI22_X1 U10513 ( .A1(n9148), .A2(n9147), .B1(n9146), .B2(n9756), .ZN(n9149)
         );
  AOI211_X1 U10514 ( .C1(n9150), .C2(n9797), .A(n10162), .B(n9149), .ZN(n9151)
         );
  OAI211_X1 U10515 ( .C1(n10021), .C2(n9153), .A(n9152), .B(n9151), .ZN(
        P1_U3239) );
  MUX2_X1 U10516 ( .A(n9549), .B(n9154), .S(n9267), .Z(n9245) );
  INV_X1 U10517 ( .A(n9230), .ZN(n9561) );
  NAND2_X1 U10518 ( .A1(n9246), .A2(n9395), .ZN(n9156) );
  MUX2_X1 U10519 ( .A(n9549), .B(n9154), .S(n9242), .Z(n9155) );
  NAND2_X1 U10520 ( .A1(n9156), .A2(n9155), .ZN(n9244) );
  INV_X1 U10521 ( .A(n7436), .ZN(n9157) );
  NAND2_X1 U10522 ( .A1(n9162), .A2(n9307), .ZN(n9355) );
  AOI21_X1 U10523 ( .B1(n9157), .B2(n9357), .A(n9355), .ZN(n9160) );
  NOR2_X1 U10524 ( .A1(n7468), .A2(n9158), .ZN(n9159) );
  MUX2_X1 U10525 ( .A(n9162), .B(n9161), .S(n9267), .Z(n9164) );
  NAND2_X1 U10526 ( .A1(n9164), .A2(n9163), .ZN(n9165) );
  NAND3_X1 U10527 ( .A1(n9169), .A2(n9168), .A3(n9296), .ZN(n9170) );
  NAND2_X1 U10528 ( .A1(n9170), .A2(n9175), .ZN(n9178) );
  AND2_X1 U10529 ( .A1(n9362), .A2(n9171), .ZN(n9361) );
  INV_X1 U10530 ( .A(n9172), .ZN(n9300) );
  AOI21_X1 U10531 ( .B1(n9173), .B2(n9361), .A(n9300), .ZN(n9176) );
  NAND2_X1 U10532 ( .A1(n9175), .A2(n9174), .ZN(n9312) );
  OAI21_X1 U10533 ( .B1(n9176), .B2(n9312), .A(n9296), .ZN(n9177) );
  MUX2_X1 U10534 ( .A(n9178), .B(n9177), .S(n9267), .Z(n9180) );
  NOR2_X1 U10535 ( .A1(n9180), .A2(n9179), .ZN(n9195) );
  NAND2_X1 U10536 ( .A1(n9189), .A2(n9297), .ZN(n9181) );
  MUX2_X1 U10537 ( .A(n9313), .B(n9181), .S(n9242), .Z(n9183) );
  OR3_X1 U10538 ( .A1(n9183), .A2(n9190), .A3(n9182), .ZN(n9194) );
  INV_X1 U10539 ( .A(n9184), .ZN(n9185) );
  OR2_X1 U10540 ( .A1(n9190), .A2(n9185), .ZN(n9186) );
  NAND2_X1 U10541 ( .A1(n9186), .A2(n9189), .ZN(n9315) );
  NAND2_X1 U10542 ( .A1(n9294), .A2(n9764), .ZN(n9199) );
  INV_X1 U10543 ( .A(n9187), .ZN(n9188) );
  AND2_X1 U10544 ( .A1(n9189), .A2(n9188), .ZN(n9298) );
  NOR2_X1 U10545 ( .A1(n9298), .A2(n9190), .ZN(n9191) );
  NOR2_X1 U10546 ( .A1(n9199), .A2(n9191), .ZN(n9192) );
  MUX2_X1 U10547 ( .A(n9315), .B(n9192), .S(n9267), .Z(n9193) );
  OAI21_X1 U10548 ( .B1(n9195), .B2(n9194), .A(n9193), .ZN(n9197) );
  NAND2_X1 U10549 ( .A1(n9198), .A2(n9196), .ZN(n9319) );
  AND3_X1 U10550 ( .A1(n9199), .A2(n9242), .A3(n9198), .ZN(n9200) );
  NOR2_X1 U10551 ( .A1(n9747), .A2(n9200), .ZN(n9201) );
  NAND2_X1 U10552 ( .A1(n9205), .A2(n9295), .ZN(n9203) );
  INV_X1 U10553 ( .A(n9321), .ZN(n9202) );
  MUX2_X1 U10554 ( .A(n9203), .B(n9202), .S(n9242), .Z(n9204) );
  NOR2_X1 U10555 ( .A1(n9204), .A2(n9206), .ZN(n9208) );
  INV_X1 U10556 ( .A(n9205), .ZN(n9326) );
  MUX2_X1 U10557 ( .A(n9206), .B(n9326), .S(n9242), .Z(n9207) );
  INV_X1 U10558 ( .A(n10010), .ZN(n9711) );
  INV_X1 U10559 ( .A(n9209), .ZN(n9396) );
  NAND2_X1 U10560 ( .A1(n9215), .A2(n9396), .ZN(n9327) );
  AOI21_X1 U10561 ( .B1(n9210), .B2(n9722), .A(n9327), .ZN(n9211) );
  MUX2_X1 U10562 ( .A(n9212), .B(n9211), .S(n9267), .Z(n9213) );
  AND2_X1 U10563 ( .A1(n9333), .A2(n9214), .ZN(n9216) );
  AND2_X1 U10564 ( .A1(n9293), .A2(n9215), .ZN(n9332) );
  MUX2_X1 U10565 ( .A(n9216), .B(n9332), .S(n9242), .Z(n9217) );
  MUX2_X1 U10566 ( .A(n9293), .B(n9333), .S(n9242), .Z(n9218) );
  INV_X1 U10567 ( .A(n9640), .ZN(n9642) );
  MUX2_X1 U10568 ( .A(n9334), .B(n9289), .S(n9267), .Z(n9219) );
  OR2_X1 U10569 ( .A1(n9991), .A2(n9220), .ZN(n9290) );
  NAND2_X1 U10570 ( .A1(n9336), .A2(n9290), .ZN(n9339) );
  MUX2_X1 U10571 ( .A(n9339), .B(n9292), .S(n9242), .Z(n9221) );
  INV_X1 U10572 ( .A(n9221), .ZN(n9222) );
  MUX2_X1 U10573 ( .A(n9336), .B(n9223), .S(n9267), .Z(n9227) );
  MUX2_X1 U10574 ( .A(n9629), .B(n9980), .S(n9242), .Z(n9224) );
  INV_X1 U10575 ( .A(n9224), .ZN(n9225) );
  NAND2_X1 U10576 ( .A1(n9596), .A2(n9225), .ZN(n9233) );
  NAND2_X1 U10577 ( .A1(n9596), .A2(n4328), .ZN(n9226) );
  AOI22_X1 U10578 ( .A1(n9228), .A2(n9227), .B1(n9233), .B2(n9226), .ZN(n9229)
         );
  INV_X1 U10579 ( .A(n9233), .ZN(n9232) );
  NAND2_X1 U10580 ( .A1(n9230), .A2(n9343), .ZN(n9231) );
  AOI21_X1 U10581 ( .B1(n9232), .B2(n9629), .A(n9231), .ZN(n9239) );
  NOR2_X1 U10582 ( .A1(n9233), .A2(n9615), .ZN(n9237) );
  INV_X1 U10583 ( .A(n9234), .ZN(n9235) );
  OR2_X1 U10584 ( .A1(n9236), .A2(n9235), .ZN(n9380) );
  NOR2_X1 U10585 ( .A1(n9237), .A2(n9380), .ZN(n9238) );
  NAND3_X1 U10586 ( .A1(n9819), .A2(n9566), .A3(n9242), .ZN(n9241) );
  OAI21_X1 U10587 ( .B1(n9384), .B2(n9242), .A(n9241), .ZN(n9243) );
  INV_X1 U10588 ( .A(n9243), .ZN(n9248) );
  OAI211_X1 U10589 ( .C1(n9246), .C2(n9245), .A(n4887), .B(n9244), .ZN(n9247)
         );
  MUX2_X1 U10590 ( .A(n9349), .B(n9288), .S(n9267), .Z(n9249) );
  INV_X1 U10591 ( .A(n9263), .ZN(n9445) );
  MUX2_X1 U10592 ( .A(n9250), .B(n9267), .S(n9259), .Z(n9271) );
  OR2_X1 U10593 ( .A1(n4282), .A2(n10076), .ZN(n9251) );
  NAND2_X1 U10594 ( .A1(n9254), .A2(n9253), .ZN(n9257) );
  OR2_X1 U10595 ( .A1(n4282), .A2(n10084), .ZN(n9256) );
  INV_X1 U10596 ( .A(n9444), .ZN(n9351) );
  OR2_X1 U10597 ( .A1(n9808), .A2(n9351), .ZN(n9258) );
  INV_X1 U10598 ( .A(n9266), .ZN(n9391) );
  AOI21_X1 U10599 ( .B1(n9523), .B2(n9444), .A(n9529), .ZN(n9264) );
  INV_X1 U10600 ( .A(n9264), .ZN(n9387) );
  INV_X1 U10601 ( .A(n9259), .ZN(n9541) );
  NOR3_X1 U10602 ( .A1(n9266), .A2(n9541), .A3(n9262), .ZN(n9261) );
  OAI21_X1 U10603 ( .B1(n9261), .B2(n9264), .A(n9260), .ZN(n9269) );
  NOR3_X1 U10604 ( .A1(n9264), .A2(n9263), .A3(n9262), .ZN(n9265) );
  INV_X1 U10605 ( .A(n9274), .ZN(n9272) );
  NAND3_X1 U10606 ( .A1(n5893), .A2(n9283), .A3(n9272), .ZN(n9273) );
  INV_X1 U10607 ( .A(n9437), .ZN(n9277) );
  NOR2_X1 U10608 ( .A1(n9283), .A2(n9274), .ZN(n9276) );
  INV_X1 U10609 ( .A(n9431), .ZN(n9275) );
  NAND4_X1 U10610 ( .A1(n9281), .A2(n9280), .A3(n9279), .A4(n9278), .ZN(n9282)
         );
  OAI211_X1 U10611 ( .C1(n9283), .C2(n9437), .A(n9282), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9443) );
  INV_X1 U10612 ( .A(n9284), .ZN(n9285) );
  NAND2_X1 U10613 ( .A1(n9384), .A2(n9285), .ZN(n9286) );
  NAND3_X1 U10614 ( .A1(n9288), .A2(n9287), .A3(n9286), .ZN(n9383) );
  AND2_X1 U10615 ( .A1(n9290), .A2(n5176), .ZN(n9291) );
  OR2_X1 U10616 ( .A1(n9292), .A2(n9291), .ZN(n9337) );
  OR2_X1 U10617 ( .A1(n9337), .A2(n5177), .ZN(n9375) );
  NAND2_X1 U10618 ( .A1(n9295), .A2(n9294), .ZN(n9323) );
  AND2_X1 U10619 ( .A1(n9297), .A2(n9296), .ZN(n9299) );
  OAI211_X1 U10620 ( .C1(n9313), .C2(n9299), .A(n9764), .B(n9298), .ZN(n9318)
         );
  OR3_X1 U10621 ( .A1(n9323), .A2(n9300), .A3(n9318), .ZN(n9301) );
  OR3_X1 U10622 ( .A1(n9327), .A2(n9326), .A3(n9301), .ZN(n9371) );
  AND2_X1 U10623 ( .A1(n9399), .A2(n9302), .ZN(n9303) );
  OAI21_X1 U10624 ( .B1(n9303), .B2(n9401), .A(n9398), .ZN(n9305) );
  AOI22_X1 U10625 ( .A1(n9305), .A2(n9304), .B1(n10219), .B2(n9460), .ZN(n9309) );
  INV_X1 U10626 ( .A(n9356), .ZN(n9308) );
  AND2_X1 U10627 ( .A1(n9307), .A2(n9306), .ZN(n9364) );
  OAI21_X1 U10628 ( .B1(n9309), .B2(n9308), .A(n9364), .ZN(n9310) );
  NAND3_X1 U10629 ( .A1(n9310), .A2(n5368), .A3(n9357), .ZN(n9311) );
  AND3_X1 U10630 ( .A1(n9311), .A2(n9363), .A3(n9362), .ZN(n9329) );
  NOR2_X1 U10631 ( .A1(n9313), .A2(n9312), .ZN(n9317) );
  OR2_X1 U10632 ( .A1(n9315), .A2(n9314), .ZN(n9316) );
  OAI21_X1 U10633 ( .B1(n9318), .B2(n9317), .A(n9316), .ZN(n9320) );
  NOR2_X1 U10634 ( .A1(n9320), .A2(n9319), .ZN(n9324) );
  OAI211_X1 U10635 ( .C1(n9324), .C2(n9323), .A(n9322), .B(n9321), .ZN(n9325)
         );
  INV_X1 U10636 ( .A(n9325), .ZN(n9328) );
  OR3_X1 U10637 ( .A1(n9328), .A2(n9327), .A3(n9326), .ZN(n9369) );
  OAI21_X1 U10638 ( .B1(n9371), .B2(n9329), .A(n9369), .ZN(n9330) );
  INV_X1 U10639 ( .A(n9330), .ZN(n9341) );
  INV_X1 U10640 ( .A(n9332), .ZN(n9335) );
  OAI211_X1 U10641 ( .C1(n4807), .C2(n9335), .A(n9334), .B(n9333), .ZN(n9340)
         );
  NAND2_X1 U10642 ( .A1(n9337), .A2(n9336), .ZN(n9338) );
  OAI21_X1 U10643 ( .B1(n9340), .B2(n9339), .A(n9338), .ZN(n9373) );
  OAI21_X1 U10644 ( .B1(n9375), .B2(n9341), .A(n9373), .ZN(n9344) );
  NAND2_X1 U10645 ( .A1(n9343), .A2(n9342), .ZN(n9376) );
  AOI21_X1 U10646 ( .B1(n9378), .B2(n9344), .A(n9376), .ZN(n9346) );
  INV_X1 U10647 ( .A(n9381), .ZN(n9345) );
  OAI21_X1 U10648 ( .B1(n9346), .B2(n9380), .A(n9345), .ZN(n9347) );
  NOR2_X1 U10649 ( .A1(n9557), .A2(n9347), .ZN(n9348) );
  NOR2_X1 U10650 ( .A1(n9383), .A2(n9348), .ZN(n9352) );
  NAND2_X1 U10651 ( .A1(n9350), .A2(n9349), .ZN(n9388) );
  NAND2_X1 U10652 ( .A1(n9808), .A2(n9351), .ZN(n9428) );
  OAI211_X1 U10653 ( .C1(n9352), .C2(n9388), .A(n9386), .B(n9428), .ZN(n9353)
         );
  XNOR2_X1 U10654 ( .A(n9354), .B(n5893), .ZN(n9441) );
  INV_X1 U10655 ( .A(n9355), .ZN(n9360) );
  NAND2_X1 U10656 ( .A1(n9357), .A2(n9356), .ZN(n9359) );
  AOI21_X1 U10657 ( .B1(n9360), .B2(n9359), .A(n9358), .ZN(n9368) );
  INV_X1 U10658 ( .A(n9361), .ZN(n9367) );
  NAND4_X1 U10659 ( .A1(n9365), .A2(n9364), .A3(n9363), .A4(n9362), .ZN(n9366)
         );
  OAI21_X1 U10660 ( .B1(n9368), .B2(n9367), .A(n9366), .ZN(n9370) );
  OAI21_X1 U10661 ( .B1(n9371), .B2(n9370), .A(n9369), .ZN(n9372) );
  INV_X1 U10662 ( .A(n9372), .ZN(n9374) );
  OAI21_X1 U10663 ( .B1(n9375), .B2(n9374), .A(n9373), .ZN(n9377) );
  AOI21_X1 U10664 ( .B1(n9378), .B2(n9377), .A(n9376), .ZN(n9379) );
  NOR2_X1 U10665 ( .A1(n9380), .A2(n9379), .ZN(n9382) );
  NOR2_X1 U10666 ( .A1(n9382), .A2(n9381), .ZN(n9385) );
  AOI21_X1 U10667 ( .B1(n9385), .B2(n9384), .A(n9383), .ZN(n9389) );
  OAI211_X1 U10668 ( .C1(n9389), .C2(n9388), .A(n9387), .B(n9386), .ZN(n9390)
         );
  INV_X1 U10669 ( .A(n9535), .ZN(n9429) );
  INV_X1 U10670 ( .A(n9393), .ZN(n9394) );
  INV_X1 U10671 ( .A(n9704), .ZN(n9692) );
  NAND2_X1 U10672 ( .A1(n9396), .A2(n9690), .ZN(n9712) );
  NAND2_X1 U10673 ( .A1(n9399), .A2(n9398), .ZN(n9400) );
  NOR2_X1 U10674 ( .A1(n9401), .A2(n9400), .ZN(n9405) );
  NAND4_X1 U10675 ( .A1(n9405), .A2(n9404), .A3(n9403), .A4(n9402), .ZN(n9408)
         );
  NOR3_X1 U10676 ( .A1(n9408), .A2(n9407), .A3(n9406), .ZN(n9412) );
  NAND4_X1 U10677 ( .A1(n9412), .A2(n9411), .A3(n9410), .A4(n9409), .ZN(n9414)
         );
  NOR2_X1 U10678 ( .A1(n9414), .A2(n9413), .ZN(n9416) );
  NAND4_X1 U10679 ( .A1(n9793), .A2(n4538), .A3(n9416), .A4(n9415), .ZN(n9417)
         );
  NOR2_X1 U10680 ( .A1(n9765), .A2(n9417), .ZN(n9418) );
  NAND3_X1 U10681 ( .A1(n9728), .A2(n5562), .A3(n9418), .ZN(n9419) );
  NOR2_X1 U10682 ( .A1(n9712), .A2(n9419), .ZN(n9420) );
  NAND3_X1 U10683 ( .A1(n9677), .A2(n9692), .A3(n9420), .ZN(n9421) );
  NOR2_X1 U10684 ( .A1(n9663), .A2(n9421), .ZN(n9423) );
  NAND2_X1 U10685 ( .A1(n5228), .A2(n9422), .ZN(n9627) );
  AND4_X1 U10686 ( .A1(n9616), .A2(n9423), .A3(n9642), .A4(n9627), .ZN(n9424)
         );
  NAND4_X1 U10687 ( .A1(n9563), .A2(n9596), .A3(n4272), .A4(n9424), .ZN(n9425)
         );
  NOR2_X1 U10688 ( .A1(n9425), .A2(n9557), .ZN(n9426) );
  NAND4_X1 U10689 ( .A1(n9429), .A2(n9428), .A3(n9427), .A4(n9426), .ZN(n9430)
         );
  OAI211_X1 U10690 ( .C1(n9434), .C2(n5893), .A(n9442), .B(n9436), .ZN(n9440)
         );
  NOR3_X1 U10691 ( .A1(n9436), .A2(n5893), .A3(n9435), .ZN(n9438) );
  MUX2_X1 U10692 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9444), .S(n9461), .Z(
        P1_U3585) );
  MUX2_X1 U10693 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9445), .S(n9461), .Z(
        P1_U3584) );
  MUX2_X1 U10694 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9446), .S(n9461), .Z(
        P1_U3583) );
  MUX2_X1 U10695 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9447), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10696 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9590), .S(n9461), .Z(
        P1_U3581) );
  MUX2_X1 U10697 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9598), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10698 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9589), .S(n9461), .Z(
        P1_U3579) );
  MUX2_X1 U10699 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9629), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10700 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9448), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10701 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9658), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10702 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9678), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10703 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9695), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10704 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9714), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10705 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9694), .S(n9461), .Z(
        P1_U3572) );
  MUX2_X1 U10706 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9750), .S(n9461), .Z(
        P1_U3571) );
  MUX2_X1 U10707 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9449), .S(n9461), .Z(
        P1_U3570) );
  MUX2_X1 U10708 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9797), .S(n9461), .Z(
        P1_U3569) );
  MUX2_X1 U10709 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9450), .S(n9461), .Z(
        P1_U3568) );
  MUX2_X1 U10710 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9795), .S(n9461), .Z(
        P1_U3567) );
  MUX2_X1 U10711 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9451), .S(n9461), .Z(
        P1_U3566) );
  MUX2_X1 U10712 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9452), .S(n9461), .Z(
        P1_U3565) );
  MUX2_X1 U10713 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9453), .S(n9461), .Z(
        P1_U3564) );
  MUX2_X1 U10714 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9454), .S(n9461), .Z(
        P1_U3563) );
  MUX2_X1 U10715 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9455), .S(n9461), .Z(
        P1_U3562) );
  MUX2_X1 U10716 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9456), .S(n9461), .Z(
        P1_U3561) );
  MUX2_X1 U10717 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9457), .S(n9461), .Z(
        P1_U3560) );
  MUX2_X1 U10718 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9458), .S(n9461), .Z(
        P1_U3559) );
  MUX2_X1 U10719 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9459), .S(n9461), .Z(
        P1_U3558) );
  MUX2_X1 U10720 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9460), .S(n9461), .Z(
        P1_U3557) );
  MUX2_X1 U10721 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n7290), .S(n9461), .Z(
        P1_U3556) );
  INV_X1 U10722 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9464) );
  XNOR2_X1 U10723 ( .A(n10148), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n10151) );
  INV_X1 U10724 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9483) );
  AOI22_X1 U10725 ( .A1(P1_REG1_REG_14__SCAN_IN), .A2(n9496), .B1(n9472), .B2(
        n9483), .ZN(n9465) );
  AOI21_X1 U10726 ( .B1(n4320), .B2(n9465), .A(n9482), .ZN(n9481) );
  INV_X1 U10727 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9478) );
  AOI21_X1 U10728 ( .B1(n10188), .B2(n9472), .A(n9466), .ZN(n9477) );
  OR2_X1 U10729 ( .A1(n9471), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9470) );
  NAND2_X1 U10730 ( .A1(n9471), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9469) );
  AND2_X1 U10731 ( .A1(n9470), .A2(n9469), .ZN(n10145) );
  INV_X1 U10732 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9474) );
  AND2_X1 U10733 ( .A1(n9473), .A2(n9474), .ZN(n9475) );
  OR3_X1 U10734 ( .A1(n10182), .A2(n9475), .A3(n9498), .ZN(n9476) );
  OAI211_X1 U10735 ( .C1(n9478), .C2(n10195), .A(n9477), .B(n9476), .ZN(n9479)
         );
  INV_X1 U10736 ( .A(n9479), .ZN(n9480) );
  OAI21_X1 U10737 ( .B1(n9481), .B2(n10132), .A(n9480), .ZN(P1_U3255) );
  AOI22_X1 U10738 ( .A1(n9511), .A2(n9514), .B1(P1_REG1_REG_18__SCAN_IN), .B2(
        n9513), .ZN(n9491) );
  XNOR2_X1 U10739 ( .A(n9488), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n10192) );
  INV_X1 U10740 ( .A(n10175), .ZN(n9487) );
  INV_X1 U10741 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9486) );
  XOR2_X1 U10742 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10175), .Z(n10177) );
  NAND2_X1 U10743 ( .A1(n10163), .A2(n9484), .ZN(n9485) );
  NAND2_X1 U10744 ( .A1(n10177), .A2(n10178), .ZN(n10176) );
  OAI21_X1 U10745 ( .B1(n9487), .B2(n9486), .A(n10176), .ZN(n10191) );
  NAND2_X1 U10746 ( .A1(n10192), .A2(n10191), .ZN(n10189) );
  OAI21_X1 U10747 ( .B1(n9489), .B2(n9488), .A(n10189), .ZN(n9490) );
  AOI21_X1 U10748 ( .B1(n9491), .B2(n9490), .A(n9512), .ZN(n9509) );
  NAND2_X1 U10749 ( .A1(n10188), .A2(n9511), .ZN(n9493) );
  NAND2_X1 U10750 ( .A1(n9493), .A2(n9492), .ZN(n9507) );
  INV_X1 U10751 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9494) );
  MUX2_X1 U10752 ( .A(P1_REG2_REG_18__SCAN_IN), .B(n9494), .S(n9511), .Z(n9495) );
  INV_X1 U10753 ( .A(n9495), .ZN(n9505) );
  NOR2_X1 U10754 ( .A1(n9497), .A2(n9496), .ZN(n9499) );
  NOR2_X1 U10755 ( .A1(n4330), .A2(n9500), .ZN(n9501) );
  INV_X1 U10756 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10159) );
  INV_X1 U10757 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9502) );
  MUX2_X1 U10758 ( .A(n9502), .B(P1_REG2_REG_16__SCAN_IN), .S(n10175), .Z(
        n10171) );
  NOR2_X1 U10759 ( .A1(n10172), .A2(n10171), .ZN(n10170) );
  NAND2_X1 U10760 ( .A1(n10187), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9503) );
  OAI21_X1 U10761 ( .B1(n10187), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9503), .ZN(
        n10183) );
  AOI211_X1 U10762 ( .C1(n9505), .C2(n9504), .A(n9510), .B(n10182), .ZN(n9506)
         );
  AOI211_X1 U10763 ( .C1(n10126), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n9507), .B(
        n9506), .ZN(n9508) );
  OAI21_X1 U10764 ( .B1(n9509), .B2(n10132), .A(n9508), .ZN(P1_U3259) );
  INV_X1 U10765 ( .A(n9516), .ZN(n9519) );
  NAND2_X1 U10766 ( .A1(n9529), .A2(n9528), .ZN(n9527) );
  XNOR2_X1 U10767 ( .A(n9805), .B(n9527), .ZN(n9807) );
  NAND2_X1 U10768 ( .A1(n9523), .A2(n9522), .ZN(n9810) );
  NOR2_X1 U10769 ( .A1(n10211), .A2(n9810), .ZN(n9531) );
  NOR2_X1 U10770 ( .A1(n9524), .A2(n9789), .ZN(n9525) );
  AOI211_X1 U10771 ( .C1(n10211), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9531), .B(
        n9525), .ZN(n9526) );
  OAI21_X1 U10772 ( .B1(n9807), .B2(n9762), .A(n9526), .ZN(P1_U3261) );
  OAI21_X1 U10773 ( .B1(n9529), .B2(n9528), .A(n9527), .ZN(n9811) );
  NOR2_X1 U10774 ( .A1(n9529), .A2(n9789), .ZN(n9530) );
  AOI211_X1 U10775 ( .C1(n10211), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9531), .B(
        n9530), .ZN(n9532) );
  OAI21_X1 U10776 ( .B1(n9762), .B2(n9811), .A(n9532), .ZN(P1_U3262) );
  NAND2_X1 U10777 ( .A1(n9534), .A2(n9533), .ZN(n9536) );
  XNOR2_X1 U10778 ( .A(n9536), .B(n9535), .ZN(n9546) );
  NAND2_X1 U10779 ( .A1(n9537), .A2(n10209), .ZN(n9545) );
  INV_X1 U10780 ( .A(n9538), .ZN(n9539) );
  AOI22_X1 U10781 ( .A1(n9539), .A2(n10201), .B1(P1_REG2_REG_29__SCAN_IN), 
        .B2(n10211), .ZN(n9540) );
  OAI21_X1 U10782 ( .B1(n9541), .B2(n9789), .A(n9540), .ZN(n9542) );
  AOI21_X1 U10783 ( .B1(n9543), .B2(n9802), .A(n9542), .ZN(n9544) );
  OAI211_X1 U10784 ( .C1(n9546), .C2(n9783), .A(n9545), .B(n9544), .ZN(
        P1_U3355) );
  AOI211_X1 U10785 ( .C1(n9557), .C2(n9548), .A(n9767), .B(n9547), .ZN(n9552)
         );
  OAI22_X1 U10786 ( .A1(n9550), .A2(n9770), .B1(n9549), .B2(n9772), .ZN(n9551)
         );
  NOR2_X1 U10787 ( .A1(n9552), .A2(n9551), .ZN(n9822) );
  AOI21_X1 U10788 ( .B1(n9819), .B2(n9571), .A(n4339), .ZN(n9820) );
  INV_X1 U10789 ( .A(n9553), .ZN(n9554) );
  AOI22_X1 U10790 ( .A1(n9554), .A2(n10201), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n10211), .ZN(n9555) );
  OAI21_X1 U10791 ( .B1(n5026), .B2(n9789), .A(n9555), .ZN(n9556) );
  AOI21_X1 U10792 ( .B1(n9820), .B2(n9802), .A(n9556), .ZN(n9559) );
  OR2_X1 U10793 ( .A1(n9823), .A2(n9783), .ZN(n9558) );
  OAI211_X1 U10794 ( .C1(n9822), .C2(n10211), .A(n9559), .B(n9558), .ZN(
        P1_U3264) );
  XNOR2_X1 U10795 ( .A(n9560), .B(n9563), .ZN(n9827) );
  XNOR2_X1 U10796 ( .A(n9564), .B(n9563), .ZN(n9565) );
  INV_X1 U10797 ( .A(n9582), .ZN(n9573) );
  INV_X1 U10798 ( .A(n9571), .ZN(n9572) );
  AOI211_X1 U10799 ( .C1(n9826), .C2(n9573), .A(n10239), .B(n9572), .ZN(n9825)
         );
  INV_X1 U10800 ( .A(n9825), .ZN(n9576) );
  INV_X1 U10801 ( .A(n9574), .ZN(n9575) );
  OAI22_X1 U10802 ( .A1(n9576), .A2(n5893), .B1(n9575), .B2(n9755), .ZN(n9577)
         );
  OAI21_X1 U10803 ( .B1(n9824), .B2(n9577), .A(n10209), .ZN(n9579) );
  AOI22_X1 U10804 ( .A1(n9826), .A2(n9758), .B1(n10211), .B2(
        P1_REG2_REG_26__SCAN_IN), .ZN(n9578) );
  OAI211_X1 U10805 ( .C1(n9827), .C2(n9783), .A(n9579), .B(n9578), .ZN(
        P1_U3265) );
  NOR2_X1 U10806 ( .A1(n9586), .A2(n9581), .ZN(n9583) );
  NOR2_X1 U10807 ( .A1(n9583), .A2(n9582), .ZN(n9829) );
  AOI22_X1 U10808 ( .A1(n9584), .A2(n10201), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n10211), .ZN(n9585) );
  OAI21_X1 U10809 ( .B1(n9586), .B2(n9789), .A(n9585), .ZN(n9592) );
  NOR2_X1 U10810 ( .A1(n9831), .A2(n10211), .ZN(n9591) );
  AOI211_X1 U10811 ( .C1(n9829), .C2(n9802), .A(n9592), .B(n9591), .ZN(n9593)
         );
  OAI21_X1 U10812 ( .B1(n9832), .B2(n9783), .A(n9593), .ZN(P1_U3266) );
  XOR2_X1 U10813 ( .A(n9594), .B(n9596), .Z(n9979) );
  OAI211_X1 U10814 ( .C1(n9597), .C2(n9596), .A(n9595), .B(n9799), .ZN(n9600)
         );
  AOI22_X1 U10815 ( .A1(n9598), .A2(n9796), .B1(n9794), .B2(n9629), .ZN(n9599)
         );
  NAND2_X1 U10816 ( .A1(n9600), .A2(n9599), .ZN(n9975) );
  OAI21_X1 U10817 ( .B1(n9611), .B2(n9606), .A(n10033), .ZN(n9601) );
  NOR2_X1 U10818 ( .A1(n9601), .A2(n9581), .ZN(n9976) );
  NAND2_X1 U10819 ( .A1(n9976), .A2(n9651), .ZN(n9605) );
  INV_X1 U10820 ( .A(n9602), .ZN(n9603) );
  AOI22_X1 U10821 ( .A1(n9603), .A2(n10201), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n10211), .ZN(n9604) );
  OAI211_X1 U10822 ( .C1(n9606), .C2(n9789), .A(n9605), .B(n9604), .ZN(n9607)
         );
  AOI21_X1 U10823 ( .B1(n9975), .B2(n10209), .A(n9607), .ZN(n9608) );
  OAI21_X1 U10824 ( .B1(n9783), .B2(n9979), .A(n9608), .ZN(P1_U3267) );
  XNOR2_X1 U10825 ( .A(n9609), .B(n9616), .ZN(n9983) );
  NOR2_X1 U10826 ( .A1(n9632), .A2(n9615), .ZN(n9610) );
  INV_X1 U10827 ( .A(n9612), .ZN(n9613) );
  AOI22_X1 U10828 ( .A1(n9613), .A2(n10201), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n10211), .ZN(n9614) );
  OAI21_X1 U10829 ( .B1(n9615), .B2(n9789), .A(n9614), .ZN(n9622) );
  AOI21_X1 U10830 ( .B1(n4343), .B2(n4789), .A(n9767), .ZN(n9620) );
  OAI22_X1 U10831 ( .A1(n9617), .A2(n9770), .B1(n9648), .B2(n9772), .ZN(n9618)
         );
  AOI21_X1 U10832 ( .B1(n9620), .B2(n9619), .A(n9618), .ZN(n9982) );
  NOR2_X1 U10833 ( .A1(n9982), .A2(n10211), .ZN(n9621) );
  AOI211_X1 U10834 ( .C1(n5219), .C2(n9802), .A(n9622), .B(n9621), .ZN(n9623)
         );
  OAI21_X1 U10835 ( .B1(n9983), .B2(n9783), .A(n9623), .ZN(P1_U3268) );
  XOR2_X1 U10836 ( .A(n9624), .B(n9627), .Z(n9988) );
  INV_X1 U10837 ( .A(n9643), .ZN(n9626) );
  NAND2_X1 U10838 ( .A1(n9626), .A2(n9625), .ZN(n9628) );
  XNOR2_X1 U10839 ( .A(n9628), .B(n9627), .ZN(n9630) );
  AOI222_X1 U10840 ( .A1(n9799), .A2(n9630), .B1(n9629), .B2(n9796), .C1(n9658), .C2(n9794), .ZN(n9987) );
  INV_X1 U10841 ( .A(n9987), .ZN(n9638) );
  INV_X1 U10842 ( .A(n9984), .ZN(n9636) );
  AND2_X1 U10843 ( .A1(n9650), .A2(n9984), .ZN(n9631) );
  NOR2_X1 U10844 ( .A1(n9632), .A2(n9631), .ZN(n9985) );
  NAND2_X1 U10845 ( .A1(n9985), .A2(n9802), .ZN(n9635) );
  AOI22_X1 U10846 ( .A1(n9633), .A2(n10201), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n10211), .ZN(n9634) );
  OAI211_X1 U10847 ( .C1(n9636), .C2(n9789), .A(n9635), .B(n9634), .ZN(n9637)
         );
  AOI21_X1 U10848 ( .B1(n9638), .B2(n10209), .A(n9637), .ZN(n9639) );
  OAI21_X1 U10849 ( .B1(n9988), .B2(n9783), .A(n9639), .ZN(P1_U3269) );
  XNOR2_X1 U10850 ( .A(n9641), .B(n9640), .ZN(n9993) );
  NOR2_X1 U10851 ( .A1(n9642), .A2(n5176), .ZN(n9645) );
  AOI21_X1 U10852 ( .B1(n9645), .B2(n9644), .A(n9643), .ZN(n9646) );
  OAI222_X1 U10853 ( .A1(n9770), .A2(n9648), .B1(n9772), .B2(n9647), .C1(n9767), .C2(n9646), .ZN(n9989) );
  AOI21_X1 U10854 ( .B1(n5224), .B2(n9991), .A(n10239), .ZN(n9649) );
  AND2_X1 U10855 ( .A1(n9650), .A2(n9649), .ZN(n9990) );
  NAND2_X1 U10856 ( .A1(n9990), .A2(n9651), .ZN(n9654) );
  AOI22_X1 U10857 ( .A1(n9652), .A2(n10201), .B1(n10211), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9653) );
  OAI211_X1 U10858 ( .C1(n5016), .C2(n9789), .A(n9654), .B(n9653), .ZN(n9655)
         );
  AOI21_X1 U10859 ( .B1(n9989), .B2(n10209), .A(n9655), .ZN(n9656) );
  OAI21_X1 U10860 ( .B1(n9993), .B2(n9783), .A(n9656), .ZN(P1_U3270) );
  XOR2_X1 U10861 ( .A(n9657), .B(n9663), .Z(n9659) );
  AOI222_X1 U10862 ( .A1(n9799), .A2(n9659), .B1(n9658), .B2(n9796), .C1(n9695), .C2(n9794), .ZN(n9997) );
  XOR2_X1 U10863 ( .A(n9685), .B(n9994), .Z(n9995) );
  INV_X1 U10864 ( .A(n9660), .ZN(n9661) );
  AOI22_X1 U10865 ( .A1(n10211), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9661), 
        .B2(n10201), .ZN(n9662) );
  OAI21_X1 U10866 ( .B1(n5017), .B2(n9789), .A(n9662), .ZN(n9668) );
  OR2_X1 U10867 ( .A1(n9664), .A2(n9663), .ZN(n9665) );
  NAND2_X1 U10868 ( .A1(n9666), .A2(n9665), .ZN(n9998) );
  NOR2_X1 U10869 ( .A1(n9998), .A2(n9783), .ZN(n9667) );
  AOI211_X1 U10870 ( .C1(n9995), .C2(n9802), .A(n9668), .B(n9667), .ZN(n9669)
         );
  OAI21_X1 U10871 ( .B1(n9997), .B2(n10211), .A(n9669), .ZN(P1_U3271) );
  NAND2_X1 U10872 ( .A1(n9671), .A2(n9670), .ZN(n9705) );
  NAND2_X1 U10873 ( .A1(n9705), .A2(n9704), .ZN(n10005) );
  NAND3_X1 U10874 ( .A1(n10005), .A2(n9677), .A3(n9672), .ZN(n9674) );
  NAND2_X1 U10875 ( .A1(n9674), .A2(n9673), .ZN(n10003) );
  OAI21_X1 U10876 ( .B1(n9677), .B2(n9676), .A(n9675), .ZN(n9679) );
  AOI222_X1 U10877 ( .A1(n9799), .A2(n9679), .B1(n9678), .B2(n9796), .C1(n9714), .C2(n9794), .ZN(n10002) );
  INV_X1 U10878 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9681) );
  OAI22_X1 U10879 ( .A1(n10209), .A2(n9681), .B1(n9680), .B2(n9755), .ZN(n9682) );
  AOI21_X1 U10880 ( .B1(n9999), .B2(n9758), .A(n9682), .ZN(n9687) );
  OR2_X1 U10881 ( .A1(n9699), .A2(n9683), .ZN(n9684) );
  AND2_X1 U10882 ( .A1(n9685), .A2(n9684), .ZN(n10000) );
  NAND2_X1 U10883 ( .A1(n10000), .A2(n9802), .ZN(n9686) );
  OAI211_X1 U10884 ( .C1(n10002), .C2(n10211), .A(n9687), .B(n9686), .ZN(n9688) );
  INV_X1 U10885 ( .A(n9688), .ZN(n9689) );
  OAI21_X1 U10886 ( .B1(n9783), .B2(n10003), .A(n9689), .ZN(P1_U3272) );
  INV_X1 U10887 ( .A(n9690), .ZN(n9691) );
  NOR2_X1 U10888 ( .A1(n4325), .A2(n9691), .ZN(n9693) );
  XNOR2_X1 U10889 ( .A(n9693), .B(n9692), .ZN(n9696) );
  AOI222_X1 U10890 ( .A1(n9799), .A2(n9696), .B1(n9695), .B2(n9796), .C1(n9694), .C2(n9794), .ZN(n10009) );
  NOR2_X1 U10891 ( .A1(n9697), .A2(n9700), .ZN(n9698) );
  NOR2_X1 U10892 ( .A1(n9700), .A2(n9789), .ZN(n9703) );
  OAI22_X1 U10893 ( .A1(n10209), .A2(n9494), .B1(n9701), .B2(n9755), .ZN(n9702) );
  AOI211_X1 U10894 ( .C1(n4312), .C2(n9802), .A(n9703), .B(n9702), .ZN(n9707)
         );
  OR2_X1 U10895 ( .A1(n9705), .A2(n9704), .ZN(n10006) );
  NAND3_X1 U10896 ( .A1(n10006), .A2(n10005), .A3(n9738), .ZN(n9706) );
  OAI211_X1 U10897 ( .C1(n10009), .C2(n10211), .A(n9707), .B(n9706), .ZN(
        P1_U3273) );
  XNOR2_X1 U10898 ( .A(n9708), .B(n9712), .ZN(n10014) );
  XNOR2_X1 U10899 ( .A(n9732), .B(n9711), .ZN(n10011) );
  AOI22_X1 U10900 ( .A1(n10211), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9709), 
        .B2(n10201), .ZN(n9710) );
  OAI21_X1 U10901 ( .B1(n9711), .B2(n9789), .A(n9710), .ZN(n9717) );
  XOR2_X1 U10902 ( .A(n9713), .B(n9712), .Z(n9715) );
  AOI222_X1 U10903 ( .A1(n9799), .A2(n9715), .B1(n9714), .B2(n9796), .C1(n9750), .C2(n9794), .ZN(n10013) );
  NOR2_X1 U10904 ( .A1(n10013), .A2(n10211), .ZN(n9716) );
  AOI211_X1 U10905 ( .C1(n10011), .C2(n9802), .A(n9717), .B(n9716), .ZN(n9718)
         );
  OAI21_X1 U10906 ( .B1(n9783), .B2(n10014), .A(n9718), .ZN(P1_U3274) );
  INV_X1 U10907 ( .A(n9719), .ZN(n9726) );
  INV_X1 U10908 ( .A(n9728), .ZN(n9720) );
  XNOR2_X1 U10909 ( .A(n9721), .B(n9720), .ZN(n9724) );
  OAI22_X1 U10910 ( .A1(n9722), .A2(n9770), .B1(n9769), .B2(n9772), .ZN(n9723)
         );
  AOI21_X1 U10911 ( .B1(n9724), .B2(n9799), .A(n9723), .ZN(n10020) );
  INV_X1 U10912 ( .A(n10020), .ZN(n9725) );
  AOI21_X1 U10913 ( .B1(n9726), .B2(n10201), .A(n9725), .ZN(n9740) );
  NAND2_X1 U10914 ( .A1(n9744), .A2(n9727), .ZN(n9729) );
  NAND2_X1 U10915 ( .A1(n9729), .A2(n9728), .ZN(n9730) );
  AND2_X1 U10916 ( .A1(n9731), .A2(n9730), .ZN(n10018) );
  AOI21_X1 U10917 ( .B1(n4396), .B2(n9734), .A(n10239), .ZN(n9733) );
  NAND2_X1 U10918 ( .A1(n9733), .A2(n9732), .ZN(n10015) );
  AOI22_X1 U10919 ( .A1(n9734), .A2(n9758), .B1(P1_REG2_REG_16__SCAN_IN), .B2(
        n10211), .ZN(n9735) );
  OAI21_X1 U10920 ( .B1(n10015), .B2(n9736), .A(n9735), .ZN(n9737) );
  AOI21_X1 U10921 ( .B1(n10018), .B2(n9738), .A(n9737), .ZN(n9739) );
  OAI21_X1 U10922 ( .B1(n9740), .B2(n10211), .A(n9739), .ZN(P1_U3275) );
  OR2_X1 U10923 ( .A1(n9773), .A2(n10021), .ZN(n9741) );
  NAND2_X1 U10924 ( .A1(n4396), .A2(n9741), .ZN(n10022) );
  NAND2_X1 U10925 ( .A1(n9742), .A2(n5562), .ZN(n9743) );
  AND2_X1 U10926 ( .A1(n9744), .A2(n9743), .ZN(n9754) );
  NAND2_X1 U10927 ( .A1(n9746), .A2(n9747), .ZN(n9748) );
  NAND2_X1 U10928 ( .A1(n9745), .A2(n9748), .ZN(n9749) );
  NAND2_X1 U10929 ( .A1(n9749), .A2(n9799), .ZN(n9752) );
  AOI22_X1 U10930 ( .A1(n9750), .A2(n9796), .B1(n9797), .B2(n9794), .ZN(n9751)
         );
  OAI211_X1 U10931 ( .C1(n9754), .C2(n9753), .A(n9752), .B(n9751), .ZN(n10024)
         );
  NAND2_X1 U10932 ( .A1(n10024), .A2(n10209), .ZN(n9761) );
  OAI22_X1 U10933 ( .A1(n10209), .A2(n10159), .B1(n9756), .B2(n9755), .ZN(
        n9757) );
  AOI21_X1 U10934 ( .B1(n9759), .B2(n9758), .A(n9757), .ZN(n9760) );
  OAI211_X1 U10935 ( .C1(n10022), .C2(n9762), .A(n9761), .B(n9760), .ZN(
        P1_U3276) );
  XNOR2_X1 U10936 ( .A(n9763), .B(n9765), .ZN(n10031) );
  NAND2_X1 U10937 ( .A1(n9791), .A2(n9764), .ZN(n9766) );
  XNOR2_X1 U10938 ( .A(n9766), .B(n9765), .ZN(n9768) );
  OAI222_X1 U10939 ( .A1(n9772), .A2(n9771), .B1(n9770), .B2(n9769), .C1(n9768), .C2(n9767), .ZN(n10027) );
  NAND2_X1 U10940 ( .A1(n10027), .A2(n10209), .ZN(n9782) );
  INV_X1 U10941 ( .A(n9786), .ZN(n9774) );
  AOI211_X1 U10942 ( .C1(n10029), .C2(n9774), .A(n10239), .B(n9773), .ZN(
        n10028) );
  INV_X1 U10943 ( .A(n9775), .ZN(n9776) );
  AOI22_X1 U10944 ( .A1(n10211), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9776), 
        .B2(n10201), .ZN(n9777) );
  OAI21_X1 U10945 ( .B1(n9778), .B2(n9789), .A(n9777), .ZN(n9779) );
  AOI21_X1 U10946 ( .B1(n10028), .B2(n9780), .A(n9779), .ZN(n9781) );
  OAI211_X1 U10947 ( .C1(n10031), .C2(n9783), .A(n9782), .B(n9781), .ZN(
        P1_U3277) );
  XNOR2_X1 U10948 ( .A(n9784), .B(n9785), .ZN(n10037) );
  AOI21_X1 U10949 ( .B1(n10032), .B2(n5216), .A(n9786), .ZN(n10034) );
  INV_X1 U10950 ( .A(n10032), .ZN(n9790) );
  AOI22_X1 U10951 ( .A1(n10211), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9787), 
        .B2(n10201), .ZN(n9788) );
  OAI21_X1 U10952 ( .B1(n9790), .B2(n9789), .A(n9788), .ZN(n9801) );
  OAI21_X1 U10953 ( .B1(n9793), .B2(n9792), .A(n9791), .ZN(n9798) );
  AOI222_X1 U10954 ( .A1(n9799), .A2(n9798), .B1(n9797), .B2(n9796), .C1(n9795), .C2(n9794), .ZN(n10036) );
  NOR2_X1 U10955 ( .A1(n10036), .A2(n10211), .ZN(n9800) );
  AOI211_X1 U10956 ( .C1(n10034), .C2(n9802), .A(n9801), .B(n9800), .ZN(n9803)
         );
  OAI21_X1 U10957 ( .B1(n10037), .B2(n9804), .A(n9803), .ZN(P1_U3278) );
  NAND2_X1 U10958 ( .A1(n9805), .A2(n10047), .ZN(n9806) );
  OAI211_X1 U10959 ( .C1(n9807), .C2(n10239), .A(n9810), .B(n9806), .ZN(n10052) );
  MUX2_X1 U10960 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n10052), .S(n10254), .Z(
        P1_U3554) );
  NAND2_X1 U10961 ( .A1(n9808), .A2(n10047), .ZN(n9809) );
  OAI211_X1 U10962 ( .C1(n9811), .C2(n10239), .A(n9810), .B(n9809), .ZN(n10053) );
  MUX2_X1 U10963 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n10053), .S(n10254), .Z(
        P1_U3553) );
  INV_X1 U10964 ( .A(n9812), .ZN(n9818) );
  OAI22_X1 U10965 ( .A1(n9815), .A2(n10239), .B1(n9814), .B2(n10237), .ZN(
        n9816) );
  INV_X1 U10966 ( .A(n9816), .ZN(n9817) );
  AOI22_X1 U10967 ( .A1(n9820), .A2(n10033), .B1(n9819), .B2(n10047), .ZN(
        n9821) );
  MUX2_X1 U10968 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10054), .S(n10254), .Z(
        P1_U3550) );
  MUX2_X1 U10969 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10055), .S(n10254), .Z(
        P1_U3549) );
  AOI22_X1 U10970 ( .A1(n9829), .A2(n10033), .B1(n9828), .B2(n10047), .ZN(
        n9830) );
  MUX2_X1 U10971 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10056), .S(n10254), .Z(
        n9974) );
  AOI22_X1 U10972 ( .A1(n5233), .A2(keyinput30), .B1(keyinput11), .B2(n9834), 
        .ZN(n9833) );
  OAI221_X1 U10973 ( .B1(n5233), .B2(keyinput30), .C1(n9834), .C2(keyinput11), 
        .A(n9833), .ZN(n9842) );
  AOI22_X1 U10974 ( .A1(n6160), .A2(keyinput22), .B1(n9947), .B2(keyinput7), 
        .ZN(n9835) );
  OAI221_X1 U10975 ( .B1(n6160), .B2(keyinput22), .C1(n9947), .C2(keyinput7), 
        .A(n9835), .ZN(n9841) );
  INV_X1 U10976 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n10304) );
  AOI22_X1 U10977 ( .A1(n10304), .A2(keyinput32), .B1(keyinput52), .B2(n9951), 
        .ZN(n9836) );
  OAI221_X1 U10978 ( .B1(n10304), .B2(keyinput32), .C1(n9951), .C2(keyinput52), 
        .A(n9836), .ZN(n9840) );
  AOI22_X1 U10979 ( .A1(n9838), .A2(keyinput6), .B1(keyinput48), .B2(n9938), 
        .ZN(n9837) );
  OAI221_X1 U10980 ( .B1(n9838), .B2(keyinput6), .C1(n9938), .C2(keyinput48), 
        .A(n9837), .ZN(n9839) );
  OR4_X1 U10981 ( .A1(n9842), .A2(n9841), .A3(n9840), .A4(n9839), .ZN(n9856)
         );
  AOI22_X1 U10982 ( .A1(n9844), .A2(keyinput13), .B1(keyinput42), .B2(n9962), 
        .ZN(n9843) );
  OAI221_X1 U10983 ( .B1(n9844), .B2(keyinput13), .C1(n9962), .C2(keyinput42), 
        .A(n9843), .ZN(n9855) );
  XOR2_X1 U10984 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput60), .Z(n9846) );
  XOR2_X1 U10985 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput0), .Z(n9845) );
  NOR2_X1 U10986 ( .A1(n9846), .A2(n9845), .ZN(n9848) );
  XNOR2_X1 U10987 ( .A(P1_REG3_REG_19__SCAN_IN), .B(keyinput62), .ZN(n9847) );
  OAI211_X1 U10988 ( .C1(keyinput3), .C2(n9967), .A(n9848), .B(n9847), .ZN(
        n9854) );
  XNOR2_X1 U10989 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput40), .ZN(n9852) );
  XNOR2_X1 U10990 ( .A(P2_REG3_REG_19__SCAN_IN), .B(keyinput51), .ZN(n9851) );
  XNOR2_X1 U10991 ( .A(P2_REG3_REG_5__SCAN_IN), .B(keyinput37), .ZN(n9850) );
  XNOR2_X1 U10992 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput38), .ZN(n9849) );
  NAND4_X1 U10993 ( .A1(n9852), .A2(n9851), .A3(n9850), .A4(n9849), .ZN(n9853)
         );
  NOR4_X1 U10994 ( .A1(n9856), .A2(n9855), .A3(n9854), .A4(n9853), .ZN(n9905)
         );
  AOI22_X1 U10995 ( .A1(n4736), .A2(keyinput8), .B1(keyinput15), .B2(n9858), 
        .ZN(n9857) );
  OAI221_X1 U10996 ( .B1(n4736), .B2(keyinput8), .C1(n9858), .C2(keyinput15), 
        .A(n9857), .ZN(n9867) );
  INV_X1 U10997 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9929) );
  AOI22_X1 U10998 ( .A1(n9929), .A2(keyinput14), .B1(n9930), .B2(keyinput44), 
        .ZN(n9859) );
  OAI221_X1 U10999 ( .B1(n9929), .B2(keyinput14), .C1(n9930), .C2(keyinput44), 
        .A(n9859), .ZN(n9866) );
  INV_X1 U11000 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n9861) );
  AOI22_X1 U11001 ( .A1(n9937), .A2(keyinput28), .B1(n9861), .B2(keyinput26), 
        .ZN(n9860) );
  OAI221_X1 U11002 ( .B1(n9937), .B2(keyinput28), .C1(n9861), .C2(keyinput26), 
        .A(n9860), .ZN(n9865) );
  INV_X1 U11003 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n10212) );
  AOI22_X1 U11004 ( .A1(n9863), .A2(keyinput1), .B1(n10212), .B2(keyinput46), 
        .ZN(n9862) );
  OAI221_X1 U11005 ( .B1(n9863), .B2(keyinput1), .C1(n10212), .C2(keyinput46), 
        .A(n9862), .ZN(n9864) );
  NOR4_X1 U11006 ( .A1(n9867), .A2(n9866), .A3(n9865), .A4(n9864), .ZN(n9904)
         );
  INV_X1 U11007 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10216) );
  AOI22_X1 U11008 ( .A1(n9502), .A2(keyinput58), .B1(n10216), .B2(keyinput56), 
        .ZN(n9868) );
  OAI221_X1 U11009 ( .B1(n9502), .B2(keyinput58), .C1(n10216), .C2(keyinput56), 
        .A(n9868), .ZN(n9879) );
  INV_X1 U11010 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10214) );
  INV_X1 U11011 ( .A(P1_RD_REG_SCAN_IN), .ZN(n9870) );
  AOI22_X1 U11012 ( .A1(n10214), .A2(keyinput20), .B1(keyinput63), .B2(n9870), 
        .ZN(n9869) );
  OAI221_X1 U11013 ( .B1(n10214), .B2(keyinput20), .C1(n9870), .C2(keyinput63), 
        .A(n9869), .ZN(n9878) );
  INV_X1 U11014 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n10305) );
  AOI22_X1 U11015 ( .A1(n10305), .A2(keyinput33), .B1(n6165), .B2(keyinput61), 
        .ZN(n9871) );
  OAI221_X1 U11016 ( .B1(n10305), .B2(keyinput33), .C1(n6165), .C2(keyinput61), 
        .A(n9871), .ZN(n9877) );
  XNOR2_X1 U11017 ( .A(P1_REG2_REG_1__SCAN_IN), .B(keyinput16), .ZN(n9875) );
  XNOR2_X1 U11018 ( .A(SI_3_), .B(keyinput27), .ZN(n9874) );
  XNOR2_X1 U11019 ( .A(SI_4_), .B(keyinput2), .ZN(n9873) );
  XNOR2_X1 U11020 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(keyinput4), .ZN(n9872) );
  NAND4_X1 U11021 ( .A1(n9875), .A2(n9874), .A3(n9873), .A4(n9872), .ZN(n9876)
         );
  NOR4_X1 U11022 ( .A1(n9879), .A2(n9878), .A3(n9877), .A4(n9876), .ZN(n9903)
         );
  INV_X1 U11023 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10213) );
  AOI22_X1 U11024 ( .A1(n10213), .A2(keyinput9), .B1(keyinput45), .B2(n9881), 
        .ZN(n9880) );
  OAI221_X1 U11025 ( .B1(n10213), .B2(keyinput9), .C1(n9881), .C2(keyinput45), 
        .A(n9880), .ZN(n9884) );
  INV_X1 U11026 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10157) );
  AOI22_X1 U11027 ( .A1(n6239), .A2(keyinput50), .B1(keyinput39), .B2(n10157), 
        .ZN(n9882) );
  OAI221_X1 U11028 ( .B1(n6239), .B2(keyinput50), .C1(n10157), .C2(keyinput39), 
        .A(n9882), .ZN(n9883) );
  NOR2_X1 U11029 ( .A1(n9884), .A2(n9883), .ZN(n9901) );
  INV_X1 U11030 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10228) );
  XNOR2_X1 U11031 ( .A(keyinput53), .B(n10228), .ZN(n9887) );
  XNOR2_X1 U11032 ( .A(keyinput17), .B(n9885), .ZN(n9886) );
  NOR2_X1 U11033 ( .A1(n9887), .A2(n9886), .ZN(n9900) );
  AOI22_X1 U11034 ( .A1(n9948), .A2(keyinput59), .B1(keyinput12), .B2(n9889), 
        .ZN(n9888) );
  OAI221_X1 U11035 ( .B1(n9948), .B2(keyinput59), .C1(n9889), .C2(keyinput12), 
        .A(n9888), .ZN(n9893) );
  AOI22_X1 U11036 ( .A1(n9891), .A2(keyinput57), .B1(keyinput41), .B2(n9952), 
        .ZN(n9890) );
  OAI221_X1 U11037 ( .B1(n9891), .B2(keyinput57), .C1(n9952), .C2(keyinput41), 
        .A(n9890), .ZN(n9892) );
  NOR2_X1 U11038 ( .A1(n9893), .A2(n9892), .ZN(n9899) );
  AOI22_X1 U11039 ( .A1(n9896), .A2(keyinput34), .B1(n9895), .B2(keyinput24), 
        .ZN(n9894) );
  OAI221_X1 U11040 ( .B1(n9896), .B2(keyinput34), .C1(n9895), .C2(keyinput24), 
        .A(n9894), .ZN(n9897) );
  INV_X1 U11041 ( .A(n9897), .ZN(n9898) );
  AND4_X1 U11042 ( .A1(n9901), .A2(n9900), .A3(n9899), .A4(n9898), .ZN(n9902)
         );
  AND4_X1 U11043 ( .A1(n9905), .A2(n9904), .A3(n9903), .A4(n9902), .ZN(n9972)
         );
  AOI22_X1 U11044 ( .A1(n9928), .A2(keyinput18), .B1(keyinput5), .B2(n9681), 
        .ZN(n9906) );
  OAI221_X1 U11045 ( .B1(n9928), .B2(keyinput18), .C1(n9681), .C2(keyinput5), 
        .A(n9906), .ZN(n9915) );
  INV_X1 U11046 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10215) );
  AOI22_X1 U11047 ( .A1(n9908), .A2(keyinput23), .B1(n10215), .B2(keyinput47), 
        .ZN(n9907) );
  OAI221_X1 U11048 ( .B1(n9908), .B2(keyinput23), .C1(n10215), .C2(keyinput47), 
        .A(n9907), .ZN(n9914) );
  INV_X1 U11049 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n9963) );
  INV_X1 U11050 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10223) );
  AOI22_X1 U11051 ( .A1(n9963), .A2(keyinput21), .B1(n10223), .B2(keyinput54), 
        .ZN(n9909) );
  OAI221_X1 U11052 ( .B1(n9963), .B2(keyinput21), .C1(n10223), .C2(keyinput54), 
        .A(n9909), .ZN(n9913) );
  AOI22_X1 U11053 ( .A1(n6182), .A2(keyinput49), .B1(n9911), .B2(keyinput29), 
        .ZN(n9910) );
  OAI221_X1 U11054 ( .B1(n6182), .B2(keyinput49), .C1(n9911), .C2(keyinput29), 
        .A(n9910), .ZN(n9912) );
  NOR4_X1 U11055 ( .A1(n9915), .A2(n9914), .A3(n9913), .A4(n9912), .ZN(n9971)
         );
  AOI22_X1 U11056 ( .A1(n9917), .A2(keyinput31), .B1(n5333), .B2(keyinput10), 
        .ZN(n9916) );
  OAI221_X1 U11057 ( .B1(n9917), .B2(keyinput31), .C1(n5333), .C2(keyinput10), 
        .A(n9916), .ZN(n9927) );
  INV_X1 U11058 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9919) );
  AOI22_X1 U11059 ( .A1(n8066), .A2(keyinput35), .B1(n9919), .B2(keyinput19), 
        .ZN(n9918) );
  OAI221_X1 U11060 ( .B1(n8066), .B2(keyinput35), .C1(n9919), .C2(keyinput19), 
        .A(n9918), .ZN(n9926) );
  AOI22_X1 U11061 ( .A1(n9921), .A2(keyinput25), .B1(keyinput43), .B2(n9935), 
        .ZN(n9920) );
  OAI221_X1 U11062 ( .B1(n9921), .B2(keyinput25), .C1(n9935), .C2(keyinput43), 
        .A(n9920), .ZN(n9925) );
  AOI22_X1 U11063 ( .A1(n9923), .A2(keyinput36), .B1(n6466), .B2(keyinput55), 
        .ZN(n9922) );
  OAI221_X1 U11064 ( .B1(n9923), .B2(keyinput36), .C1(n6466), .C2(keyinput55), 
        .A(n9922), .ZN(n9924) );
  NOR4_X1 U11065 ( .A1(n9927), .A2(n9926), .A3(n9925), .A4(n9924), .ZN(n9970)
         );
  NOR3_X1 U11066 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .A3(P2_REG2_REG_19__SCAN_IN), .ZN(n9933) );
  NOR4_X1 U11067 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_REG2_REG_19__SCAN_IN), 
        .A3(n9928), .A4(n6182), .ZN(n9932) );
  NOR4_X1 U11068 ( .A1(P1_REG0_REG_7__SCAN_IN), .A2(n9930), .A3(n10223), .A4(
        n9929), .ZN(n9931) );
  NAND4_X1 U11069 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9933), .A3(n9932), .A4(
        n9931), .ZN(n9961) );
  NAND4_X1 U11070 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), 
        .A3(P1_REG0_REG_5__SCAN_IN), .A4(n9934), .ZN(n9946) );
  NAND4_X1 U11071 ( .A1(SI_15_), .A2(P2_REG2_REG_2__SCAN_IN), .A3(
        P2_REG0_REG_30__SCAN_IN), .A4(n9935), .ZN(n9936) );
  NOR2_X1 U11072 ( .A1(n6160), .A2(n9936), .ZN(n9942) );
  AND4_X1 U11073 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P1_DATAO_REG_25__SCAN_IN), 
        .A3(P2_REG2_REG_1__SCAN_IN), .A4(n9937), .ZN(n9940) );
  NOR4_X1 U11074 ( .A1(P1_RD_REG_SCAN_IN), .A2(SI_23_), .A3(
        P1_REG2_REG_16__SCAN_IN), .A4(n9938), .ZN(n9939) );
  AND2_X1 U11075 ( .A1(n9940), .A2(n9939), .ZN(n9941) );
  NAND4_X1 U11076 ( .A1(n9943), .A2(P2_D_REG_21__SCAN_IN), .A3(n9942), .A4(
        n9941), .ZN(n9945) );
  NAND4_X1 U11077 ( .A1(SI_4_), .A2(SI_3_), .A3(SI_25_), .A4(
        P1_REG3_REG_27__SCAN_IN), .ZN(n9944) );
  NOR3_X1 U11078 ( .A1(n9946), .A2(n9945), .A3(n9944), .ZN(n9958) );
  NAND4_X1 U11079 ( .A1(n9948), .A2(n10228), .A3(n9947), .A4(
        P1_REG2_REG_26__SCAN_IN), .ZN(n9950) );
  NAND4_X1 U11080 ( .A1(n6293), .A2(P2_IR_REG_16__SCAN_IN), .A3(
        P2_REG3_REG_19__SCAN_IN), .A4(P1_REG2_REG_1__SCAN_IN), .ZN(n9949) );
  NOR2_X1 U11081 ( .A1(n9950), .A2(n9949), .ZN(n9956) );
  NAND4_X1 U11082 ( .A1(n9952), .A2(n9951), .A3(P1_DATAO_REG_11__SCAN_IN), 
        .A4(P2_REG3_REG_5__SCAN_IN), .ZN(n9953) );
  NOR2_X1 U11083 ( .A1(n9954), .A2(n9953), .ZN(n9955) );
  NAND4_X1 U11084 ( .A1(n9958), .A2(n9957), .A3(n9956), .A4(n9955), .ZN(n9960)
         );
  OR3_X1 U11085 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .ZN(n9959) );
  NOR3_X1 U11086 ( .A1(n9961), .A2(n9960), .A3(n9959), .ZN(n9966) );
  NOR4_X1 U11087 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(P2_REG3_REG_14__SCAN_IN), 
        .A3(n9962), .A4(n6466), .ZN(n9965) );
  NOR4_X1 U11088 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P2_B_REG_SCAN_IN), .A3(
        P1_ADDR_REG_13__SCAN_IN), .A4(n9963), .ZN(n9964) );
  AND3_X1 U11089 ( .A1(n9966), .A2(n9965), .A3(n9964), .ZN(n9968) );
  OAI21_X1 U11090 ( .B1(n9968), .B2(keyinput3), .A(n9967), .ZN(n9969) );
  NAND4_X1 U11091 ( .A1(n9972), .A2(n9971), .A3(n9970), .A4(n9969), .ZN(n9973)
         );
  XNOR2_X1 U11092 ( .A(n9974), .B(n9973), .ZN(P1_U3548) );
  AOI211_X1 U11093 ( .C1(n9977), .C2(n10047), .A(n9976), .B(n9975), .ZN(n9978)
         );
  OAI21_X1 U11094 ( .B1(n9753), .B2(n9979), .A(n9978), .ZN(n10057) );
  MUX2_X1 U11095 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10057), .S(n10254), .Z(
        P1_U3547) );
  AOI22_X1 U11096 ( .A1(n5219), .A2(n10033), .B1(n9980), .B2(n10047), .ZN(
        n9981) );
  OAI211_X1 U11097 ( .C1(n9753), .C2(n9983), .A(n9982), .B(n9981), .ZN(n10058)
         );
  MUX2_X1 U11098 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10058), .S(n10254), .Z(
        P1_U3546) );
  AOI22_X1 U11099 ( .A1(n9985), .A2(n10033), .B1(n9984), .B2(n10047), .ZN(
        n9986) );
  OAI211_X1 U11100 ( .C1(n9753), .C2(n9988), .A(n9987), .B(n9986), .ZN(n10059)
         );
  MUX2_X1 U11101 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10059), .S(n10254), .Z(
        P1_U3545) );
  AOI211_X1 U11102 ( .C1(n9991), .C2(n10047), .A(n9990), .B(n9989), .ZN(n9992)
         );
  OAI21_X1 U11103 ( .B1(n9753), .B2(n9993), .A(n9992), .ZN(n10060) );
  MUX2_X1 U11104 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10060), .S(n10254), .Z(
        P1_U3544) );
  AOI22_X1 U11105 ( .A1(n9995), .A2(n10033), .B1(n9994), .B2(n10047), .ZN(
        n9996) );
  OAI211_X1 U11106 ( .C1(n9753), .C2(n9998), .A(n9997), .B(n9996), .ZN(n10061)
         );
  MUX2_X1 U11107 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10061), .S(n10254), .Z(
        P1_U3543) );
  AOI22_X1 U11108 ( .A1(n10000), .A2(n10033), .B1(n9999), .B2(n10047), .ZN(
        n10001) );
  OAI211_X1 U11109 ( .C1(n9753), .C2(n10003), .A(n10002), .B(n10001), .ZN(
        n10062) );
  MUX2_X1 U11110 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10062), .S(n10254), .Z(
        P1_U3542) );
  AOI22_X1 U11111 ( .A1(n4312), .A2(n10033), .B1(n10004), .B2(n10047), .ZN(
        n10008) );
  NAND3_X1 U11112 ( .A1(n10006), .A2(n10005), .A3(n10234), .ZN(n10007) );
  NAND3_X1 U11113 ( .A1(n10009), .A2(n10008), .A3(n10007), .ZN(n10063) );
  MUX2_X1 U11114 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10063), .S(n10254), .Z(
        P1_U3541) );
  AOI22_X1 U11115 ( .A1(n10011), .A2(n10033), .B1(n10010), .B2(n10047), .ZN(
        n10012) );
  OAI211_X1 U11116 ( .C1(n9753), .C2(n10014), .A(n10013), .B(n10012), .ZN(
        n10064) );
  MUX2_X1 U11117 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10064), .S(n10254), .Z(
        P1_U3540) );
  OAI21_X1 U11118 ( .B1(n10016), .B2(n10237), .A(n10015), .ZN(n10017) );
  AOI21_X1 U11119 ( .B1(n10018), .B2(n10234), .A(n10017), .ZN(n10019) );
  NAND2_X1 U11120 ( .A1(n10020), .A2(n10019), .ZN(n10065) );
  MUX2_X1 U11121 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10065), .S(n10254), .Z(
        P1_U3539) );
  INV_X1 U11122 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10025) );
  OAI22_X1 U11123 ( .A1(n10022), .A2(n10239), .B1(n10021), .B2(n10237), .ZN(
        n10023) );
  NOR2_X1 U11124 ( .A1(n10024), .A2(n10023), .ZN(n10066) );
  MUX2_X1 U11125 ( .A(n10025), .B(n10066), .S(n10254), .Z(n10026) );
  INV_X1 U11126 ( .A(n10026), .ZN(P1_U3538) );
  AOI211_X1 U11127 ( .C1(n10029), .C2(n10047), .A(n10028), .B(n10027), .ZN(
        n10030) );
  OAI21_X1 U11128 ( .B1(n9753), .B2(n10031), .A(n10030), .ZN(n10069) );
  MUX2_X1 U11129 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10069), .S(n10254), .Z(
        P1_U3537) );
  AOI22_X1 U11130 ( .A1(n10034), .A2(n10033), .B1(n10032), .B2(n10047), .ZN(
        n10035) );
  OAI211_X1 U11131 ( .C1(n9753), .C2(n10037), .A(n10036), .B(n10035), .ZN(
        n10070) );
  MUX2_X1 U11132 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n10070), .S(n10254), .Z(
        P1_U3536) );
  OAI211_X1 U11133 ( .C1(n10040), .C2(n10237), .A(n10039), .B(n10038), .ZN(
        n10071) );
  MUX2_X1 U11134 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10071), .S(n10254), .Z(
        P1_U3535) );
  AOI211_X1 U11135 ( .C1(n10043), .C2(n10047), .A(n10042), .B(n10041), .ZN(
        n10044) );
  OAI21_X1 U11136 ( .B1(n9753), .B2(n10045), .A(n10044), .ZN(n10072) );
  MUX2_X1 U11137 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n10072), .S(n10254), .Z(
        P1_U3533) );
  AOI21_X1 U11138 ( .B1(n10048), .B2(n10047), .A(n10046), .ZN(n10049) );
  OAI211_X1 U11139 ( .C1(n9753), .C2(n10051), .A(n10050), .B(n10049), .ZN(
        n10073) );
  MUX2_X1 U11140 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10073), .S(n10254), .Z(
        P1_U3532) );
  MUX2_X1 U11141 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n10052), .S(n10245), .Z(
        P1_U3522) );
  MUX2_X1 U11142 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n10053), .S(n10245), .Z(
        P1_U3521) );
  MUX2_X1 U11143 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10055), .S(n10245), .Z(
        P1_U3517) );
  MUX2_X1 U11144 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10056), .S(n10245), .Z(
        P1_U3516) );
  MUX2_X1 U11145 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10057), .S(n10245), .Z(
        P1_U3515) );
  MUX2_X1 U11146 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10058), .S(n10245), .Z(
        P1_U3514) );
  MUX2_X1 U11147 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10059), .S(n10245), .Z(
        P1_U3513) );
  MUX2_X1 U11148 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10060), .S(n10245), .Z(
        P1_U3512) );
  MUX2_X1 U11149 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10061), .S(n10245), .Z(
        P1_U3511) );
  MUX2_X1 U11150 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10062), .S(n10245), .Z(
        P1_U3510) );
  MUX2_X1 U11151 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10063), .S(n10245), .Z(
        P1_U3508) );
  MUX2_X1 U11152 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10064), .S(n10245), .Z(
        P1_U3505) );
  MUX2_X1 U11153 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10065), .S(n10245), .Z(
        P1_U3502) );
  INV_X1 U11154 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10067) );
  MUX2_X1 U11155 ( .A(n10067), .B(n10066), .S(n10245), .Z(n10068) );
  INV_X1 U11156 ( .A(n10068), .ZN(P1_U3499) );
  MUX2_X1 U11157 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10069), .S(n10245), .Z(
        P1_U3496) );
  MUX2_X1 U11158 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n10070), .S(n10245), .Z(
        P1_U3493) );
  MUX2_X1 U11159 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n10071), .S(n10245), .Z(
        P1_U3490) );
  MUX2_X1 U11160 ( .A(P1_REG0_REG_10__SCAN_IN), .B(n10072), .S(n10245), .Z(
        P1_U3484) );
  MUX2_X1 U11161 ( .A(P1_REG0_REG_9__SCAN_IN), .B(n10073), .S(n10245), .Z(
        P1_U3481) );
  MUX2_X1 U11162 ( .A(n10074), .B(P1_D_REG_0__SCAN_IN), .S(n10218), .Z(
        P1_U3440) );
  INV_X1 U11163 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n10075) );
  NAND3_X1 U11164 ( .A1(n10075), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n10077) );
  OAI22_X1 U11165 ( .A1(n10078), .A2(n10077), .B1(n10076), .B2(n10094), .ZN(
        n10079) );
  AOI21_X1 U11166 ( .B1(n10080), .B2(n10089), .A(n10079), .ZN(n10081) );
  INV_X1 U11167 ( .A(n10081), .ZN(P1_U3322) );
  OAI222_X1 U11168 ( .A1(n10094), .A2(n10084), .B1(n10087), .B2(n10083), .C1(
        P1_U3084), .C2(n10082), .ZN(P1_U3323) );
  OAI222_X1 U11169 ( .A1(n10094), .A2(n10088), .B1(n10087), .B2(n10086), .C1(
        n10085), .C2(P1_U3084), .ZN(P1_U3324) );
  NAND2_X1 U11170 ( .A1(n10090), .A2(n10089), .ZN(n10092) );
  OAI211_X1 U11171 ( .C1(n10094), .C2(n10093), .A(n10092), .B(n10091), .ZN(
        P1_U3326) );
  MUX2_X1 U11172 ( .A(n10095), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  NOR2_X1 U11173 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10096) );
  AOI21_X1 U11174 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n10096), .ZN(n10359) );
  NOR2_X1 U11175 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10097) );
  AOI21_X1 U11176 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n10097), .ZN(n10362) );
  NOR2_X1 U11177 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10098) );
  AOI21_X1 U11178 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10098), .ZN(n10365) );
  NOR2_X1 U11179 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10099) );
  AOI21_X1 U11180 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n10099), .ZN(n10368) );
  NOR2_X1 U11181 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(P2_ADDR_REG_13__SCAN_IN), 
        .ZN(n10100) );
  AOI21_X1 U11182 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10100), .ZN(n10371) );
  NOR2_X1 U11183 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10107) );
  XNOR2_X1 U11184 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10398) );
  NAND2_X1 U11185 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n10105) );
  XOR2_X1 U11186 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10396) );
  NAND2_X1 U11187 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n10103) );
  XOR2_X1 U11188 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10394) );
  AOI21_X1 U11189 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10353) );
  INV_X1 U11190 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10101) );
  NAND3_X1 U11191 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10355) );
  NAND2_X1 U11192 ( .A1(n10394), .A2(n10393), .ZN(n10102) );
  NAND2_X1 U11193 ( .A1(n10103), .A2(n10102), .ZN(n10395) );
  NAND2_X1 U11194 ( .A1(n10396), .A2(n10395), .ZN(n10104) );
  NAND2_X1 U11195 ( .A1(n10105), .A2(n10104), .ZN(n10397) );
  NOR2_X1 U11196 ( .A1(n10398), .A2(n10397), .ZN(n10106) );
  NOR2_X1 U11197 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10108), .ZN(n10383) );
  NAND2_X1 U11198 ( .A1(n10110), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n10111) );
  XOR2_X1 U11199 ( .A(n10110), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10381) );
  NAND2_X1 U11200 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n10112), .ZN(n10113) );
  XOR2_X1 U11201 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n10112), .Z(n10392) );
  NAND2_X1 U11202 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n10114), .ZN(n10116) );
  XOR2_X1 U11203 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n10114), .Z(n10391) );
  NAND2_X1 U11204 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10391), .ZN(n10115) );
  NAND2_X1 U11205 ( .A1(n10116), .A2(n10115), .ZN(n10117) );
  AND2_X1 U11206 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10117), .ZN(n10118) );
  XNOR2_X1 U11207 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n10117), .ZN(n10389) );
  NAND2_X1 U11208 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n10119) );
  OAI21_X1 U11209 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n10119), .ZN(n10379) );
  NAND2_X1 U11210 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n10120) );
  OAI21_X1 U11211 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n10120), .ZN(n10376) );
  NOR2_X1 U11212 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10121) );
  AOI21_X1 U11213 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n10121), .ZN(n10373) );
  NAND2_X1 U11214 ( .A1(n10368), .A2(n10367), .ZN(n10366) );
  NAND2_X1 U11215 ( .A1(n10365), .A2(n10364), .ZN(n10363) );
  NAND2_X1 U11216 ( .A1(n10359), .A2(n10358), .ZN(n10357) );
  NOR2_X1 U11217 ( .A1(n8490), .A2(n10386), .ZN(n10122) );
  NAND2_X1 U11218 ( .A1(n8490), .A2(n10386), .ZN(n10385) );
  XOR2_X1 U11219 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .Z(n10123) );
  XNOR2_X1 U11220 ( .A(n10124), .B(n10123), .ZN(ADD_1071_U4) );
  XNOR2_X1 U11221 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11222 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  AOI22_X1 U11223 ( .A1(n10126), .A2(P1_ADDR_REG_8__SCAN_IN), .B1(n10125), 
        .B2(n10188), .ZN(n10140) );
  INV_X1 U11224 ( .A(n10127), .ZN(n10139) );
  INV_X1 U11225 ( .A(n10128), .ZN(n10129) );
  OAI211_X1 U11226 ( .C1(n10131), .C2(n10130), .A(n10129), .B(n10143), .ZN(
        n10138) );
  AOI21_X1 U11227 ( .B1(n10134), .B2(n10133), .A(n10132), .ZN(n10136) );
  NAND2_X1 U11228 ( .A1(n10136), .A2(n10135), .ZN(n10137) );
  NAND4_X1 U11229 ( .A1(n10140), .A2(n10139), .A3(n10138), .A4(n10137), .ZN(
        P1_U3249) );
  INV_X1 U11230 ( .A(n10141), .ZN(n10142) );
  OAI211_X1 U11231 ( .C1(n10145), .C2(n10144), .A(n10143), .B(n10142), .ZN(
        n10146) );
  OAI211_X1 U11232 ( .C1(n10149), .C2(n10148), .A(n10147), .B(n10146), .ZN(
        n10150) );
  INV_X1 U11233 ( .A(n10150), .ZN(n10156) );
  NOR2_X1 U11234 ( .A1(n10152), .A2(n10151), .ZN(n10153) );
  OAI21_X1 U11235 ( .B1(n10154), .B2(n10153), .A(n10190), .ZN(n10155) );
  OAI211_X1 U11236 ( .C1(n10195), .C2(n10157), .A(n10156), .B(n10155), .ZN(
        P1_U3254) );
  INV_X1 U11237 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10168) );
  AOI211_X1 U11238 ( .C1(n10160), .C2(n10159), .A(n10158), .B(n10182), .ZN(
        n10161) );
  AOI211_X1 U11239 ( .C1(n10188), .C2(n10163), .A(n10162), .B(n10161), .ZN(
        n10167) );
  OAI211_X1 U11240 ( .C1(n10165), .C2(P1_REG1_REG_15__SCAN_IN), .A(n10190), 
        .B(n10164), .ZN(n10166) );
  OAI211_X1 U11241 ( .C1(n10168), .C2(n10195), .A(n10167), .B(n10166), .ZN(
        P1_U3256) );
  INV_X1 U11242 ( .A(n10169), .ZN(n10174) );
  AOI211_X1 U11243 ( .C1(n10172), .C2(n10171), .A(n10170), .B(n10182), .ZN(
        n10173) );
  AOI211_X1 U11244 ( .C1(n10188), .C2(n10175), .A(n10174), .B(n10173), .ZN(
        n10180) );
  OAI211_X1 U11245 ( .C1(n10178), .C2(n10177), .A(n10190), .B(n10176), .ZN(
        n10179) );
  OAI211_X1 U11246 ( .C1(n4431), .C2(n10195), .A(n10180), .B(n10179), .ZN(
        P1_U3257) );
  INV_X1 U11247 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10196) );
  INV_X1 U11248 ( .A(n10181), .ZN(n10186) );
  AOI211_X1 U11249 ( .C1(n10184), .C2(n10183), .A(n4388), .B(n10182), .ZN(
        n10185) );
  AOI211_X1 U11250 ( .C1(n10188), .C2(n10187), .A(n10186), .B(n10185), .ZN(
        n10194) );
  OAI211_X1 U11251 ( .C1(n10192), .C2(n10191), .A(n10190), .B(n10189), .ZN(
        n10193) );
  OAI211_X1 U11252 ( .C1(n10196), .C2(n10195), .A(n10194), .B(n10193), .ZN(
        P1_U3258) );
  INV_X1 U11253 ( .A(n10197), .ZN(n10203) );
  AOI22_X1 U11254 ( .A1(n10201), .A2(n10200), .B1(n10199), .B2(n10198), .ZN(
        n10202) );
  OAI21_X1 U11255 ( .B1(n10203), .B2(n5893), .A(n10202), .ZN(n10206) );
  INV_X1 U11256 ( .A(n10204), .ZN(n10205) );
  AOI211_X1 U11257 ( .C1(n10208), .C2(n10207), .A(n10206), .B(n10205), .ZN(
        n10210) );
  AOI22_X1 U11258 ( .A1(n10211), .A2(n7032), .B1(n10210), .B2(n10209), .ZN(
        P1_U3286) );
  AND2_X1 U11259 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10218), .ZN(P1_U3292) );
  AND2_X1 U11260 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10218), .ZN(P1_U3293) );
  AND2_X1 U11261 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10218), .ZN(P1_U3294) );
  AND2_X1 U11262 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10218), .ZN(P1_U3295) );
  AND2_X1 U11263 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10218), .ZN(P1_U3296) );
  AND2_X1 U11264 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10218), .ZN(P1_U3297) );
  INV_X1 U11265 ( .A(n10218), .ZN(n10217) );
  NOR2_X1 U11266 ( .A1(n10217), .A2(n10212), .ZN(P1_U3298) );
  NOR2_X1 U11267 ( .A1(n10217), .A2(n10213), .ZN(P1_U3299) );
  AND2_X1 U11268 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10218), .ZN(P1_U3300) );
  AND2_X1 U11269 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10218), .ZN(P1_U3301) );
  AND2_X1 U11270 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10218), .ZN(P1_U3302) );
  AND2_X1 U11271 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10218), .ZN(P1_U3303) );
  AND2_X1 U11272 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10218), .ZN(P1_U3304) );
  AND2_X1 U11273 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10218), .ZN(P1_U3305) );
  AND2_X1 U11274 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10218), .ZN(P1_U3306) );
  AND2_X1 U11275 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10218), .ZN(P1_U3307) );
  AND2_X1 U11276 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10218), .ZN(P1_U3308) );
  AND2_X1 U11277 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10218), .ZN(P1_U3309) );
  AND2_X1 U11278 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10218), .ZN(P1_U3310) );
  NOR2_X1 U11279 ( .A1(n10217), .A2(n10214), .ZN(P1_U3311) );
  NOR2_X1 U11280 ( .A1(n10217), .A2(n10215), .ZN(P1_U3312) );
  AND2_X1 U11281 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10218), .ZN(P1_U3313) );
  AND2_X1 U11282 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10218), .ZN(P1_U3314) );
  AND2_X1 U11283 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10218), .ZN(P1_U3315) );
  AND2_X1 U11284 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10218), .ZN(P1_U3316) );
  AND2_X1 U11285 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10218), .ZN(P1_U3317) );
  AND2_X1 U11286 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10218), .ZN(P1_U3318) );
  NOR2_X1 U11287 ( .A1(n10217), .A2(n10216), .ZN(P1_U3319) );
  AND2_X1 U11288 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10218), .ZN(P1_U3320) );
  AND2_X1 U11289 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10218), .ZN(P1_U3321) );
  OAI22_X1 U11290 ( .A1(n10220), .A2(n10239), .B1(n10219), .B2(n10237), .ZN(
        n10222) );
  NOR2_X1 U11291 ( .A1(n10222), .A2(n10221), .ZN(n10246) );
  AOI22_X1 U11292 ( .A1(n10245), .A2(n10246), .B1(n10223), .B2(n10243), .ZN(
        P1_U3460) );
  OAI22_X1 U11293 ( .A1(n10225), .A2(n10239), .B1(n10224), .B2(n10237), .ZN(
        n10227) );
  NOR2_X1 U11294 ( .A1(n10227), .A2(n10226), .ZN(n10248) );
  AOI22_X1 U11295 ( .A1(n10245), .A2(n10248), .B1(n10228), .B2(n10243), .ZN(
        P1_U3466) );
  OAI22_X1 U11296 ( .A1(n10230), .A2(n10239), .B1(n10229), .B2(n10237), .ZN(
        n10232) );
  AOI211_X1 U11297 ( .C1(n10234), .C2(n10233), .A(n10232), .B(n10231), .ZN(
        n10250) );
  INV_X1 U11298 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10235) );
  AOI22_X1 U11299 ( .A1(n10245), .A2(n10250), .B1(n10235), .B2(n10243), .ZN(
        P1_U3472) );
  INV_X1 U11300 ( .A(n10236), .ZN(n10238) );
  OAI22_X1 U11301 ( .A1(n10240), .A2(n10239), .B1(n10238), .B2(n10237), .ZN(
        n10242) );
  NOR2_X1 U11302 ( .A1(n10242), .A2(n10241), .ZN(n10253) );
  INV_X1 U11303 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10244) );
  AOI22_X1 U11304 ( .A1(n10245), .A2(n10253), .B1(n10244), .B2(n10243), .ZN(
        P1_U3478) );
  AOI22_X1 U11305 ( .A1(n10254), .A2(n10246), .B1(n7017), .B2(n10251), .ZN(
        P1_U3525) );
  AOI22_X1 U11306 ( .A1(n10254), .A2(n10248), .B1(n10247), .B2(n10251), .ZN(
        P1_U3527) );
  AOI22_X1 U11307 ( .A1(n10254), .A2(n10250), .B1(n10249), .B2(n10251), .ZN(
        P1_U3529) );
  AOI22_X1 U11308 ( .A1(n10254), .A2(n10253), .B1(n10252), .B2(n10251), .ZN(
        P1_U3531) );
  AOI22_X1 U11309 ( .A1(n10256), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10255), .ZN(n10266) );
  AOI21_X1 U11310 ( .B1(n10258), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n10257), .ZN(
        n10265) );
  NOR2_X1 U11311 ( .A1(n10259), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n10263) );
  OAI21_X1 U11312 ( .B1(P2_REG1_REG_0__SCAN_IN), .B2(n10261), .A(n10260), .ZN(
        n10262) );
  OAI21_X1 U11313 ( .B1(n10263), .B2(n10262), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n10264) );
  OAI211_X1 U11314 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n10266), .A(n10265), .B(
        n10264), .ZN(P2_U3245) );
  AOI22_X1 U11315 ( .A1(n10267), .A2(n6334), .B1(P2_REG2_REG_3__SCAN_IN), .B2(
        n10276), .ZN(n10274) );
  OAI22_X1 U11316 ( .A1(n10270), .A2(n10269), .B1(n10281), .B2(n10268), .ZN(
        n10271) );
  AOI21_X1 U11317 ( .B1(n10286), .B2(n10272), .A(n10271), .ZN(n10273) );
  OAI211_X1 U11318 ( .C1(n10276), .C2(n10275), .A(n10274), .B(n10273), .ZN(
        P2_U3293) );
  AOI21_X1 U11319 ( .B1(n10285), .B2(n10313), .A(n10328), .ZN(n10278) );
  NAND2_X1 U11320 ( .A1(n10278), .A2(n10277), .ZN(n10319) );
  INV_X1 U11321 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10280) );
  OAI22_X1 U11322 ( .A1(n10281), .A2(n10319), .B1(n10280), .B2(n10279), .ZN(
        n10282) );
  INV_X1 U11323 ( .A(n10282), .ZN(n10301) );
  OAI21_X1 U11324 ( .B1(n7338), .B2(n10283), .A(n7537), .ZN(n10322) );
  NAND2_X1 U11325 ( .A1(n10284), .A2(n10322), .ZN(n10299) );
  NAND2_X1 U11326 ( .A1(n10286), .A2(n10285), .ZN(n10298) );
  INV_X1 U11327 ( .A(n10287), .ZN(n10292) );
  INV_X1 U11328 ( .A(n10288), .ZN(n10289) );
  NAND2_X1 U11329 ( .A1(n7338), .A2(n10289), .ZN(n10291) );
  OAI211_X1 U11330 ( .C1(n10293), .C2(n10292), .A(n10291), .B(n10290), .ZN(
        n10296) );
  INV_X1 U11331 ( .A(n10294), .ZN(n10295) );
  AND2_X1 U11332 ( .A1(n10296), .A2(n10295), .ZN(n10323) );
  MUX2_X1 U11333 ( .A(n10323), .B(n9858), .S(n10276), .Z(n10297) );
  AND3_X1 U11334 ( .A1(n10299), .A2(n10298), .A3(n10297), .ZN(n10300) );
  NAND2_X1 U11335 ( .A1(n10301), .A2(n10300), .ZN(P2_U3295) );
  AND2_X1 U11336 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10309), .ZN(P2_U3297) );
  AND2_X1 U11337 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10309), .ZN(P2_U3298) );
  AND2_X1 U11338 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10309), .ZN(P2_U3299) );
  AND2_X1 U11339 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10309), .ZN(P2_U3300) );
  AND2_X1 U11340 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10309), .ZN(P2_U3301) );
  AND2_X1 U11341 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10309), .ZN(P2_U3302) );
  AND2_X1 U11342 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10309), .ZN(P2_U3303) );
  AND2_X1 U11343 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10309), .ZN(P2_U3304) );
  AND2_X1 U11344 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10309), .ZN(P2_U3305) );
  AND2_X1 U11345 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10309), .ZN(P2_U3306) );
  NOR2_X1 U11346 ( .A1(n10306), .A2(n10304), .ZN(P2_U3307) );
  AND2_X1 U11347 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10309), .ZN(P2_U3308) );
  AND2_X1 U11348 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10309), .ZN(P2_U3309) );
  AND2_X1 U11349 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10309), .ZN(P2_U3310) );
  AND2_X1 U11350 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10309), .ZN(P2_U3311) );
  AND2_X1 U11351 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10309), .ZN(P2_U3312) );
  NOR2_X1 U11352 ( .A1(n10306), .A2(n10305), .ZN(P2_U3313) );
  AND2_X1 U11353 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10309), .ZN(P2_U3314) );
  AND2_X1 U11354 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10309), .ZN(P2_U3315) );
  AND2_X1 U11355 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10309), .ZN(P2_U3316) );
  AND2_X1 U11356 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10309), .ZN(P2_U3317) );
  AND2_X1 U11357 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10309), .ZN(P2_U3318) );
  AND2_X1 U11358 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10309), .ZN(P2_U3319) );
  AND2_X1 U11359 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10309), .ZN(P2_U3320) );
  AND2_X1 U11360 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10309), .ZN(P2_U3321) );
  AND2_X1 U11361 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10309), .ZN(P2_U3322) );
  AND2_X1 U11362 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10309), .ZN(P2_U3323) );
  AND2_X1 U11363 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10309), .ZN(P2_U3324) );
  AND2_X1 U11364 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10309), .ZN(P2_U3325) );
  AND2_X1 U11365 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10309), .ZN(P2_U3326) );
  AOI22_X1 U11366 ( .A1(n10312), .A2(n10308), .B1(n10307), .B2(n10309), .ZN(
        P2_U3437) );
  AOI22_X1 U11367 ( .A1(n10312), .A2(n10311), .B1(n10310), .B2(n10309), .ZN(
        P2_U3438) );
  AOI22_X1 U11368 ( .A1(n10315), .A2(n10331), .B1(n10314), .B2(n10313), .ZN(
        n10316) );
  AND2_X1 U11369 ( .A1(n10317), .A2(n10316), .ZN(n10347) );
  INV_X1 U11370 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10318) );
  AOI22_X1 U11371 ( .A1(n10345), .A2(n10347), .B1(n10318), .B2(n4655), .ZN(
        P2_U3451) );
  OAI21_X1 U11372 ( .B1(n10320), .B2(n10326), .A(n10319), .ZN(n10321) );
  AOI21_X1 U11373 ( .B1(n10322), .B2(n10331), .A(n10321), .ZN(n10324) );
  AND2_X1 U11374 ( .A1(n10324), .A2(n10323), .ZN(n10348) );
  INV_X1 U11375 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10325) );
  AOI22_X1 U11376 ( .A1(n10345), .A2(n10348), .B1(n10325), .B2(n4655), .ZN(
        P2_U3454) );
  OAI22_X1 U11377 ( .A1(n10329), .A2(n10328), .B1(n10327), .B2(n10326), .ZN(
        n10330) );
  AOI21_X1 U11378 ( .B1(n10332), .B2(n10331), .A(n10330), .ZN(n10334) );
  AND2_X1 U11379 ( .A1(n10334), .A2(n10333), .ZN(n10349) );
  INV_X1 U11380 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10335) );
  AOI22_X1 U11381 ( .A1(n10345), .A2(n10349), .B1(n10335), .B2(n4655), .ZN(
        P2_U3469) );
  AOI21_X1 U11382 ( .B1(n10338), .B2(n10337), .A(n10336), .ZN(n10339) );
  OAI211_X1 U11383 ( .C1(n10342), .C2(n10341), .A(n10340), .B(n10339), .ZN(
        n10343) );
  INV_X1 U11384 ( .A(n10343), .ZN(n10351) );
  INV_X1 U11385 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10344) );
  AOI22_X1 U11386 ( .A1(n10345), .A2(n10351), .B1(n10344), .B2(n4655), .ZN(
        P2_U3475) );
  AOI22_X1 U11387 ( .A1(n10352), .A2(n10347), .B1(n10346), .B2(n4653), .ZN(
        P2_U3520) );
  AOI22_X1 U11388 ( .A1(n10352), .A2(n10348), .B1(n6297), .B2(n4653), .ZN(
        P2_U3521) );
  AOI22_X1 U11389 ( .A1(n10352), .A2(n10349), .B1(n6211), .B2(n4653), .ZN(
        P2_U3526) );
  AOI22_X1 U11390 ( .A1(n10352), .A2(n10351), .B1(n10350), .B2(n4653), .ZN(
        P2_U3528) );
  INV_X1 U11391 ( .A(n10353), .ZN(n10354) );
  NAND2_X1 U11392 ( .A1(n10355), .A2(n10354), .ZN(n10356) );
  XNOR2_X1 U11393 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10356), .ZN(ADD_1071_U5)
         );
  XOR2_X1 U11394 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11395 ( .B1(n10359), .B2(n10358), .A(n10357), .ZN(ADD_1071_U56) );
  OAI21_X1 U11396 ( .B1(n10362), .B2(n10361), .A(n10360), .ZN(ADD_1071_U57) );
  OAI21_X1 U11397 ( .B1(n10365), .B2(n10364), .A(n10363), .ZN(ADD_1071_U58) );
  OAI21_X1 U11398 ( .B1(n10368), .B2(n10367), .A(n10366), .ZN(ADD_1071_U59) );
  OAI21_X1 U11399 ( .B1(n10371), .B2(n10370), .A(n10369), .ZN(ADD_1071_U60) );
  OAI21_X1 U11400 ( .B1(n10374), .B2(n10373), .A(n10372), .ZN(ADD_1071_U61) );
  AOI21_X1 U11401 ( .B1(n10377), .B2(n10376), .A(n10375), .ZN(ADD_1071_U62) );
  AOI21_X1 U11402 ( .B1(n10380), .B2(n10379), .A(n10378), .ZN(ADD_1071_U63) );
  XOR2_X1 U11403 ( .A(n10381), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11404 ( .A1(n10383), .A2(n10382), .ZN(n10384) );
  XOR2_X1 U11405 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10384), .Z(ADD_1071_U51) );
  OAI21_X1 U11406 ( .B1(n8490), .B2(n10386), .A(n10385), .ZN(n10387) );
  XNOR2_X1 U11407 ( .A(n10387), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11408 ( .B1(n10390), .B2(n10389), .A(n10388), .ZN(ADD_1071_U47) );
  XOR2_X1 U11409 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10391), .Z(ADD_1071_U48) );
  XOR2_X1 U11410 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10392), .Z(ADD_1071_U49) );
  XOR2_X1 U11411 ( .A(n10394), .B(n10393), .Z(ADD_1071_U54) );
  XOR2_X1 U11412 ( .A(n10395), .B(n10396), .Z(ADD_1071_U53) );
  XNOR2_X1 U11413 ( .A(n10398), .B(n10397), .ZN(ADD_1071_U52) );
  AND2_X2 U4803 ( .A1(n6932), .A2(n10314), .ZN(n7313) );
  CLKBUF_X1 U4777 ( .A(n6059), .Z(n4720) );
  CLKBUF_X1 U4796 ( .A(n6332), .Z(n6573) );
endmodule

