

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput63, keyinput62, keyinput61, keyinput60, keyinput59, keyinput58, 
        keyinput57, keyinput56, keyinput55, keyinput54, keyinput53, keyinput52, 
        keyinput51, keyinput50, keyinput49, keyinput48, keyinput47, keyinput46, 
        keyinput45, keyinput44, keyinput43, keyinput42, keyinput41, keyinput40, 
        keyinput39, keyinput38, keyinput37, keyinput36, keyinput35, keyinput34, 
        keyinput33, keyinput32, keyinput31, keyinput30, keyinput29, keyinput28, 
        keyinput27, keyinput26, keyinput25, keyinput24, keyinput23, keyinput22, 
        keyinput21, keyinput20, keyinput19, keyinput18, keyinput17, keyinput16, 
        keyinput15, keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, 
        keyinput9, keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, 
        keyinput3, keyinput2, keyinput1, keyinput0 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput63,
         keyinput62, keyinput61, keyinput60, keyinput59, keyinput58,
         keyinput57, keyinput56, keyinput55, keyinput54, keyinput53,
         keyinput52, keyinput51, keyinput50, keyinput49, keyinput48,
         keyinput47, keyinput46, keyinput45, keyinput44, keyinput43,
         keyinput42, keyinput41, keyinput40, keyinput39, keyinput38,
         keyinput37, keyinput36, keyinput35, keyinput34, keyinput33,
         keyinput32, keyinput31, keyinput30, keyinput29, keyinput28,
         keyinput27, keyinput26, keyinput25, keyinput24, keyinput23,
         keyinput22, keyinput21, keyinput20, keyinput19, keyinput18,
         keyinput17, keyinput16, keyinput15, keyinput14, keyinput13,
         keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, keyinput7,
         keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, keyinput1,
         keyinput0;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287;

  NOR2_X1 U7136 ( .A1(n13960), .A2(n13959), .ZN(n14174) );
  NAND2_X1 U7137 ( .A1(n7389), .A2(n7386), .ZN(n14187) );
  INV_X4 U7138 ( .A(n10140), .ZN(n11981) );
  INV_X1 U7140 ( .A(n7723), .ZN(n8201) );
  CLKBUF_X2 U7141 ( .A(n9417), .Z(n6399) );
  NAND2_X1 U7142 ( .A1(n6925), .A2(n6468), .ZN(n13790) );
  OR2_X1 U7143 ( .A1(n8981), .A2(n6926), .ZN(n6925) );
  NAND2_X1 U7144 ( .A1(n6969), .A2(n6972), .ZN(n9764) );
  CLKBUF_X1 U7145 ( .A(n14819), .Z(n6388) );
  AND2_X1 U7146 ( .A1(n10501), .A2(n13407), .ZN(n14819) );
  INV_X2 U7147 ( .A(n9023), .ZN(n9448) );
  INV_X1 U7148 ( .A(n12670), .ZN(n7173) );
  AND3_X1 U7149 ( .A1(n8401), .A2(n8400), .A3(n8399), .ZN(n15055) );
  INV_X1 U7150 ( .A(n12402), .ZN(n12415) );
  NOR3_X1 U7151 ( .A1(n13305), .A2(n7062), .A3(n7061), .ZN(n13267) );
  NAND2_X1 U7152 ( .A1(n13411), .A2(n13575), .ZN(n13389) );
  OR2_X1 U7153 ( .A1(n10187), .A2(n10499), .ZN(n10362) );
  AND2_X1 U7154 ( .A1(n6627), .A2(n8963), .ZN(n7603) );
  CLKBUF_X2 U7155 ( .A(n8416), .Z(n11147) );
  INV_X2 U7156 ( .A(n12586), .ZN(n12559) );
  AND2_X1 U7157 ( .A1(n12424), .A2(n12253), .ZN(n12402) );
  OR2_X1 U7158 ( .A1(n8484), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8502) );
  INV_X1 U7159 ( .A(n8637), .ZN(n12212) );
  INV_X1 U7160 ( .A(n12449), .ZN(n15047) );
  CLKBUF_X3 U7161 ( .A(n7725), .Z(n8262) );
  INV_X2 U7162 ( .A(n13390), .ZN(n10035) );
  INV_X2 U7163 ( .A(n9584), .ZN(n9276) );
  NAND2_X1 U7164 ( .A1(n11982), .A2(n14662), .ZN(n10259) );
  INV_X1 U7165 ( .A(n9036), .ZN(n9434) );
  AND2_X2 U7166 ( .A1(n8975), .A2(n14287), .ZN(n9433) );
  NOR2_X1 U7167 ( .A1(n15065), .A2(n10622), .ZN(n12259) );
  CLKBUF_X3 U7168 ( .A(n8402), .Z(n6885) );
  INV_X1 U7169 ( .A(n14646), .ZN(n10617) );
  CLKBUF_X2 U7170 ( .A(n9417), .Z(n6398) );
  AND4_X1 U7171 ( .A1(n9077), .A2(n9076), .A3(n9075), .A4(n9074), .ZN(n10612)
         );
  XNOR2_X1 U7172 ( .A(n8686), .B(n8685), .ZN(n12594) );
  INV_X1 U7173 ( .A(n14852), .ZN(n14850) );
  INV_X1 U7174 ( .A(n9419), .ZN(n9096) );
  OR2_X1 U7175 ( .A1(n12073), .A2(n12072), .ZN(n6389) );
  NAND2_X1 U7176 ( .A1(n6392), .A2(n12974), .ZN(n6390) );
  NAND2_X2 U7177 ( .A1(n6392), .A2(n12974), .ZN(n10696) );
  XNOR2_X2 U7178 ( .A(n10631), .B(n13788), .ZN(n10633) );
  AOI21_X2 U7179 ( .B1(n11289), .B2(n6718), .A(n6511), .ZN(n6717) );
  OAI21_X2 U7180 ( .B1(n14465), .B2(n6569), .A(n6567), .ZN(n12787) );
  AOI21_X2 U7182 ( .B1(n9899), .B2(P2_REG2_REG_7__SCAN_IN), .A(n9893), .ZN(
        n9910) );
  NAND2_X2 U7183 ( .A1(n14048), .A2(n14047), .ZN(n14046) );
  NOR2_X2 U7184 ( .A1(n14222), .A2(n7384), .ZN(n14048) );
  INV_X1 U7185 ( .A(n11935), .ZN(n6391) );
  XNOR2_X2 U7186 ( .A(n7222), .B(n11907), .ZN(n13760) );
  NOR4_X2 U7187 ( .A1(n9494), .A2(n9493), .A3(n13926), .A4(n9492), .ZN(n9495)
         );
  NAND2_X2 U7188 ( .A1(n7695), .A2(n6456), .ZN(n13111) );
  NAND2_X2 U7189 ( .A1(n13315), .A2(n13555), .ZN(n13305) );
  AND2_X2 U7190 ( .A1(n8180), .A2(n8179), .ZN(n13555) );
  NAND2_X4 U7191 ( .A1(n10227), .A2(n6762), .ZN(n10229) );
  XNOR2_X2 U7192 ( .A(n13907), .B(n13926), .ZN(n14164) );
  OAI21_X2 U7193 ( .B1(n12650), .B2(n12649), .A(n12248), .ZN(n12638) );
  AOI22_X2 U7194 ( .A1(n12660), .A2(n12659), .B1(n12667), .B2(n12135), .ZN(
        n12650) );
  XNOR2_X1 U7195 ( .A(n10910), .B(n12442), .ZN(n11230) );
  NOR2_X2 U7196 ( .A1(n9498), .A2(n8962), .ZN(n6627) );
  OAI22_X2 U7197 ( .A1(n12648), .A2(n12647), .B1(n12917), .B2(n12433), .ZN(
        n12637) );
  NAND2_X2 U7198 ( .A1(n7537), .A2(n7538), .ZN(n12648) );
  XNOR2_X1 U7199 ( .A(n8376), .B(n8375), .ZN(n6392) );
  CLKBUF_X2 U7200 ( .A(n9650), .Z(n6393) );
  XNOR2_X2 U7201 ( .A(n7298), .B(P3_IR_REG_26__SCAN_IN), .ZN(n11579) );
  OAI21_X2 U7202 ( .B1(n8888), .B2(P3_IR_REG_25__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7298) );
  OAI21_X2 U7203 ( .B1(n8684), .B2(n8683), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n8686) );
  NAND2_X1 U7204 ( .A1(n13972), .A2(n7396), .ZN(n7395) );
  NAND2_X1 U7205 ( .A1(n14187), .A2(n6477), .ZN(n13973) );
  AOI211_X1 U7206 ( .C1(n12597), .C2(n14993), .A(n12596), .B(n12595), .ZN(
        n12598) );
  NAND2_X1 U7207 ( .A1(n6846), .A2(n13894), .ZN(n14085) );
  AND2_X1 U7208 ( .A1(n6788), .A2(n6517), .ZN(n6968) );
  NOR2_X1 U7209 ( .A1(n12150), .A2(n6789), .ZN(n12148) );
  NOR2_X1 U7210 ( .A1(n12511), .A2(n12510), .ZN(n12531) );
  NAND2_X1 U7211 ( .A1(n14620), .A2(n11223), .ZN(n11276) );
  NAND2_X1 U7212 ( .A1(n8538), .A2(n12304), .ZN(n11600) );
  XNOR2_X1 U7213 ( .A(n8070), .B(SI_18_), .ZN(n8068) );
  NAND2_X1 U7214 ( .A1(n7022), .A2(n7021), .ZN(n8070) );
  NAND2_X1 U7215 ( .A1(n6682), .A2(n7847), .ZN(n14831) );
  INV_X1 U7216 ( .A(n9998), .ZN(n10047) );
  NAND2_X1 U7217 ( .A1(n14613), .A2(n14608), .ZN(n14125) );
  AND2_X1 U7218 ( .A1(n12270), .A2(n12266), .ZN(n15040) );
  INV_X2 U7219 ( .A(n10259), .ZN(n11985) );
  INV_X4 U7220 ( .A(n12089), .ZN(n12111) );
  INV_X1 U7221 ( .A(n13109), .ZN(n10355) );
  INV_X1 U7222 ( .A(n13108), .ZN(n10473) );
  INV_X2 U7223 ( .A(n10229), .ZN(n12089) );
  CLKBUF_X2 U7224 ( .A(n10199), .Z(n12995) );
  CLKBUF_X2 U7225 ( .A(P2_U3947), .Z(n6394) );
  INV_X2 U7226 ( .A(n9980), .ZN(n9982) );
  INV_X2 U7227 ( .A(n11983), .ZN(n11948) );
  AND2_X1 U7228 ( .A1(n8391), .A2(n8390), .ZN(n8850) );
  NAND4_X2 U7229 ( .A1(n7730), .A2(n7729), .A3(n7728), .A4(n7727), .ZN(n13110)
         );
  INV_X1 U7230 ( .A(n8312), .ZN(n9995) );
  INV_X1 U7231 ( .A(n10601), .ZN(n10023) );
  NAND2_X2 U7232 ( .A1(n9444), .A2(n11354), .ZN(n9842) );
  NAND2_X4 U7233 ( .A1(n13790), .A2(n13796), .ZN(n9584) );
  INV_X2 U7234 ( .A(n8116), .ZN(n8213) );
  OR2_X1 U7235 ( .A1(n8637), .A2(n9572), .ZN(n6787) );
  AND2_X1 U7236 ( .A1(n11856), .A2(n8365), .ZN(n8416) );
  OR2_X1 U7237 ( .A1(n12213), .A2(n9573), .ZN(n8382) );
  AND2_X1 U7238 ( .A1(n13593), .A2(n11845), .ZN(n7725) );
  INV_X2 U7239 ( .A(n7723), .ZN(n7674) );
  NAND2_X1 U7240 ( .A1(n9507), .A2(n9508), .ZN(n14297) );
  NAND2_X1 U7241 ( .A1(n8303), .A2(n7657), .ZN(n9737) );
  OR2_X1 U7242 ( .A1(n9511), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n9507) );
  AND2_X1 U7243 ( .A1(n9226), .A2(n8984), .ZN(n8987) );
  INV_X1 U7244 ( .A(n9534), .ZN(n7866) );
  NAND2_X2 U7245 ( .A1(n7650), .A2(n6897), .ZN(n9534) );
  NAND3_X1 U7246 ( .A1(n9052), .A2(n7224), .A3(n7223), .ZN(n9057) );
  INV_X4 U7247 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  OAI21_X1 U7248 ( .B1(n13548), .B2(n14846), .A(n6547), .ZN(n13549) );
  OR2_X1 U7249 ( .A1(n13955), .A2(n13954), .ZN(n14166) );
  NAND2_X1 U7250 ( .A1(n7395), .A2(n7393), .ZN(n14165) );
  OAI21_X1 U7251 ( .B1(n12613), .B2(n7534), .A(n15108), .ZN(n8945) );
  AOI21_X1 U7252 ( .B1(n13279), .B2(n14520), .A(n13278), .ZN(n13457) );
  NAND2_X1 U7253 ( .A1(n6660), .A2(n6659), .ZN(n12202) );
  XNOR2_X1 U7254 ( .A(n13179), .B(n11868), .ZN(n11864) );
  NAND2_X1 U7255 ( .A1(n14000), .A2(n6651), .ZN(n13988) );
  NAND3_X1 U7256 ( .A1(n7036), .A2(n13040), .A3(n7038), .ZN(n13039) );
  AND2_X1 U7257 ( .A1(n6786), .A2(n12691), .ZN(n6785) );
  AND2_X1 U7258 ( .A1(n7060), .A2(n6518), .ZN(n13221) );
  NAND2_X1 U7259 ( .A1(n8941), .A2(n12393), .ZN(n12391) );
  XNOR2_X1 U7260 ( .A(n8255), .B(n8254), .ZN(n13586) );
  AND2_X1 U7261 ( .A1(n7088), .A2(n7084), .ZN(n7083) );
  OAI21_X1 U7262 ( .B1(n8103), .B2(n8102), .A(n6438), .ZN(n8121) );
  NAND2_X1 U7263 ( .A1(n6589), .A2(n13194), .ZN(n13367) );
  XNOR2_X1 U7264 ( .A(n8249), .B(n8248), .ZN(n13595) );
  AOI21_X1 U7265 ( .B1(n14085), .B2(n14084), .A(n13897), .ZN(n14071) );
  NOR2_X1 U7266 ( .A1(n6481), .A2(n6968), .ZN(n12121) );
  NAND2_X1 U7267 ( .A1(n6590), .A2(n13191), .ZN(n13382) );
  NAND2_X1 U7268 ( .A1(n6572), .A2(n8875), .ZN(n12700) );
  AOI21_X1 U7269 ( .B1(n6428), .B2(n7045), .A(n7041), .ZN(n7040) );
  AOI21_X1 U7270 ( .B1(n12533), .B2(n12532), .A(n12531), .ZN(n12562) );
  NAND2_X1 U7271 ( .A1(n6883), .A2(n7192), .ZN(n12724) );
  NAND2_X1 U7272 ( .A1(n7032), .A2(n8172), .ZN(n7033) );
  XNOR2_X1 U7273 ( .A(n11998), .B(n11999), .ZN(n11997) );
  AND2_X1 U7274 ( .A1(n6588), .A2(n6592), .ZN(n13185) );
  NAND2_X1 U7275 ( .A1(n12509), .A2(n12508), .ZN(n12530) );
  NAND2_X1 U7276 ( .A1(n14508), .A2(n11803), .ZN(n11998) );
  NAND2_X1 U7277 ( .A1(n6828), .A2(n6827), .ZN(n11554) );
  NAND2_X1 U7278 ( .A1(n11544), .A2(n11543), .ZN(n11546) );
  NAND2_X1 U7279 ( .A1(n11363), .A2(n11362), .ZN(n11638) );
  NAND2_X1 U7280 ( .A1(n11600), .A2(n6469), .ZN(n12811) );
  NAND2_X1 U7281 ( .A1(n6909), .A2(n11454), .ZN(n11380) );
  NAND2_X1 U7282 ( .A1(n11378), .A2(n11377), .ZN(n11454) );
  NAND2_X1 U7283 ( .A1(n6886), .A2(n8130), .ZN(n8143) );
  NAND2_X1 U7284 ( .A1(n7095), .A2(n7091), .ZN(n11056) );
  AOI21_X1 U7285 ( .B1(n10682), .B2(P1_REG1_REG_13__SCAN_IN), .A(n10681), .ZN(
        n10683) );
  NAND2_X1 U7286 ( .A1(n10907), .A2(n10906), .ZN(n6764) );
  NAND2_X1 U7287 ( .A1(n8070), .A2(SI_18_), .ZN(n8071) );
  NAND2_X1 U7288 ( .A1(n7937), .A2(n7936), .ZN(n14696) );
  NAND2_X1 U7289 ( .A1(n8010), .A2(n6474), .ZN(n7022) );
  NAND2_X1 U7290 ( .A1(n9130), .A2(n9129), .ZN(n11348) );
  NAND2_X1 U7291 ( .A1(n7894), .A2(n7893), .ZN(n11208) );
  NAND2_X1 U7292 ( .A1(n9149), .A2(n9148), .ZN(n11312) );
  NAND2_X1 U7293 ( .A1(n6575), .A2(n6573), .ZN(n8003) );
  NAND2_X1 U7294 ( .A1(n7842), .A2(n6812), .ZN(n9581) );
  INV_X1 U7295 ( .A(n12227), .ZN(n7180) );
  NAND2_X1 U7296 ( .A1(n10533), .A2(n7197), .ZN(n11035) );
  NAND2_X1 U7297 ( .A1(n6939), .A2(n8482), .ZN(n11389) );
  INV_X2 U7298 ( .A(n14613), .ZN(n14091) );
  NAND2_X1 U7299 ( .A1(n7761), .A2(n7760), .ZN(n10499) );
  AND2_X2 U7300 ( .A1(n10663), .A2(n12822), .ZN(n12826) );
  NAND2_X1 U7301 ( .A1(n7794), .A2(n7793), .ZN(n7797) );
  NAND2_X2 U7302 ( .A1(n14009), .A2(n14638), .ZN(n14613) );
  AND2_X1 U7303 ( .A1(n12288), .A2(n12279), .ZN(n12276) );
  AND2_X1 U7304 ( .A1(n7738), .A2(n7739), .ZN(n11008) );
  INV_X1 U7305 ( .A(n10221), .ZN(n10220) );
  INV_X2 U7306 ( .A(n10199), .ZN(n12048) );
  INV_X1 U7307 ( .A(n13787), .ZN(n10636) );
  NAND4_X1 U7308 ( .A1(n7765), .A2(n7764), .A3(n7763), .A4(n7762), .ZN(n13109)
         );
  NAND4_X1 U7309 ( .A1(n9066), .A2(n9065), .A3(n9064), .A4(n9063), .ZN(n13787)
         );
  AND4_X1 U7310 ( .A1(n8406), .A2(n8405), .A3(n8404), .A4(n8403), .ZN(n15045)
         );
  AND4_X1 U7311 ( .A1(n8437), .A2(n8436), .A3(n8435), .A4(n8434), .ZN(n11116)
         );
  NAND2_X2 U7312 ( .A1(n9842), .A2(n9817), .ZN(n11983) );
  AOI21_X1 U7313 ( .B1(n7023), .B2(n6414), .A(n6540), .ZN(n7021) );
  BUF_X2 U7314 ( .A(n7768), .Z(n8298) );
  NAND2_X2 U7315 ( .A1(n9842), .A2(n9841), .ZN(n11935) );
  NAND4_X1 U7316 ( .A1(n8385), .A2(n8384), .A3(n8386), .A4(n8383), .ZN(n12449)
         );
  NAND4_X1 U7317 ( .A1(n8366), .A2(n8369), .A3(n8367), .A4(n8368), .ZN(n15065)
         );
  INV_X4 U7318 ( .A(n8242), .ZN(n7768) );
  AND2_X1 U7319 ( .A1(n9038), .A2(n9037), .ZN(n6887) );
  NAND3_X1 U7320 ( .A1(n8382), .A2(n6787), .A3(n6432), .ZN(n15074) );
  OAI21_X1 U7321 ( .B1(n7824), .B2(n7412), .A(n7863), .ZN(n7411) );
  AND2_X2 U7322 ( .A1(n8364), .A2(n12968), .ZN(n11146) );
  OR2_X1 U7323 ( .A1(n9036), .A2(n9035), .ZN(n9037) );
  NAND2_X1 U7324 ( .A1(n6964), .A2(n6965), .ZN(n11088) );
  AND3_X1 U7325 ( .A1(n8415), .A2(n8414), .A3(n8413), .ZN(n10756) );
  INV_X1 U7326 ( .A(n15055), .ZN(n6395) );
  NAND2_X1 U7327 ( .A1(n6903), .A2(n6900), .ZN(n14294) );
  NAND2_X1 U7328 ( .A1(n8975), .A2(n8976), .ZN(n9417) );
  OR2_X1 U7329 ( .A1(n11267), .A2(n11579), .ZN(n8890) );
  INV_X1 U7330 ( .A(n8365), .ZN(n12968) );
  NOR2_X1 U7331 ( .A1(n11396), .A2(n9863), .ZN(n10497) );
  XNOR2_X1 U7332 ( .A(n7668), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8286) );
  AND2_X1 U7333 ( .A1(n6774), .A2(n8888), .ZN(n11267) );
  INV_X1 U7334 ( .A(n14287), .ZN(n8976) );
  XNOR2_X1 U7335 ( .A(n8887), .B(n8356), .ZN(n11453) );
  INV_X1 U7336 ( .A(n8364), .ZN(n11856) );
  OAI21_X1 U7337 ( .B1(n6681), .B2(SI_1_), .A(n7698), .ZN(n7683) );
  INV_X1 U7338 ( .A(n8844), .ZN(n12586) );
  NAND2_X1 U7339 ( .A1(n6681), .A2(SI_1_), .ZN(n7698) );
  NAND2_X2 U7340 ( .A1(n9525), .A2(P3_U3151), .ZN(n12973) );
  XNOR2_X1 U7341 ( .A(n8376), .B(n8375), .ZN(n8844) );
  INV_X2 U7342 ( .A(n7866), .ZN(n9525) );
  NOR2_X1 U7343 ( .A1(n9081), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n7199) );
  NAND2_X1 U7344 ( .A1(n6442), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8376) );
  OR2_X1 U7345 ( .A1(n7638), .A2(n7827), .ZN(n7639) );
  NAND2_X1 U7346 ( .A1(n6680), .A2(n6679), .ZN(n6681) );
  OR2_X1 U7347 ( .A1(n8565), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n8684) );
  OAI21_X1 U7348 ( .B1(n8834), .B2(n7551), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n8377) );
  BUF_X1 U7349 ( .A(n9059), .Z(n9081) );
  NAND2_X1 U7350 ( .A1(n6770), .A2(n6491), .ZN(n6769) );
  XNOR2_X1 U7351 ( .A(n7708), .B(n7707), .ZN(n9650) );
  AND2_X1 U7352 ( .A1(n7633), .A2(n7634), .ZN(n7583) );
  AND4_X1 U7353 ( .A1(n7632), .A2(n7631), .A3(n7630), .A4(n7629), .ZN(n7633)
         );
  INV_X4 U7354 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7355 ( .A(P2_RD_REG_SCAN_IN), .ZN(n15256) );
  INV_X1 U7356 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n15212) );
  NOR2_X1 U7357 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n8960) );
  NOR3_X1 U7358 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .A3(
        P1_IR_REG_8__SCAN_IN), .ZN(n8967) );
  NOR2_X1 U7359 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n7219) );
  INV_X1 U7360 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9003) );
  NOR2_X1 U7361 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n7218) );
  NOR2_X2 U7362 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n8342) );
  NOR2_X1 U7363 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n8964) );
  INV_X1 U7364 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9052) );
  INV_X4 U7365 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7366 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n8986) );
  INV_X1 U7367 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8984) );
  INV_X1 U7368 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n7844) );
  INV_X1 U7369 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n7826) );
  NOR2_X1 U7370 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n7618) );
  INV_X1 U7371 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7646) );
  INV_X1 U7372 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n14444) );
  OAI22_X2 U7373 ( .A1(n12724), .A2(n8874), .B1(n12742), .B2(n12935), .ZN(
        n12712) );
  OAI21_X2 U7374 ( .B1(n12130), .B2(n12132), .A(n12131), .ZN(n12129) );
  INV_X1 U7375 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6396) );
  INV_X1 U7376 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6397) );
  NAND2_X2 U7377 ( .A1(n9062), .A2(n9061), .ZN(n10331) );
  AOI21_X2 U7378 ( .B1(n12141), .B2(n12140), .A(n12065), .ZN(n12150) );
  OR2_X1 U7379 ( .A1(n7706), .A2(n6396), .ZN(n7707) );
  INV_X1 U7380 ( .A(n8975), .ZN(n14284) );
  XNOR2_X2 U7381 ( .A(n8998), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9444) );
  XNOR2_X2 U7382 ( .A(n9039), .B(P1_IR_REG_1__SCAN_IN), .ZN(n9698) );
  NAND4_X2 U7383 ( .A1(n7613), .A2(n7708), .A3(n7560), .A4(n7559), .ZN(n7758)
         );
  INV_X2 U7384 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7559) );
  NOR2_X2 U7385 ( .A1(n13389), .A2(n13370), .ZN(n13371) );
  INV_X1 U7386 ( .A(n9096), .ZN(n6400) );
  NAND2_X1 U7387 ( .A1(n14284), .A2(n8976), .ZN(n9419) );
  XNOR2_X2 U7388 ( .A(n9053), .B(n9052), .ZN(n13801) );
  OR2_X1 U7389 ( .A1(n9051), .A2(n6397), .ZN(n9053) );
  XNOR2_X2 U7390 ( .A(n7296), .B(n7634), .ZN(n13600) );
  NAND2_X1 U7391 ( .A1(n11982), .A2(n14662), .ZN(n6401) );
  NAND2_X1 U7392 ( .A1(n6391), .A2(n14662), .ZN(n6402) );
  NAND2_X1 U7393 ( .A1(n8700), .A2(n8699), .ZN(n8702) );
  NOR2_X1 U7394 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n7182) );
  XNOR2_X1 U7395 ( .A(n11868), .B(n8296), .ZN(n8327) );
  INV_X1 U7396 ( .A(n11825), .ZN(n6694) );
  NAND4_X1 U7397 ( .A1(n7665), .A2(n7799), .A3(n7583), .A4(n7078), .ZN(n7651)
         );
  AND2_X1 U7398 ( .A1(n7628), .A2(n6973), .ZN(n7078) );
  OAI22_X1 U7399 ( .A1(n10635), .A2(n10140), .B1(n11935), .B2(n7255), .ZN(
        n10141) );
  NAND2_X1 U7400 ( .A1(n7421), .A2(n7424), .ZN(n8226) );
  NAND2_X1 U7401 ( .A1(n7033), .A2(n6466), .ZN(n7421) );
  AND2_X1 U7402 ( .A1(n7429), .A2(n7423), .ZN(n7422) );
  NAND2_X1 U7403 ( .A1(n8003), .A2(n6478), .ZN(n8010) );
  OR2_X1 U7404 ( .A1(n12066), .A2(n12726), .ZN(n7326) );
  AOI21_X1 U7405 ( .B1(n10912), .B2(n10911), .A(n6472), .ZN(n10913) );
  NAND2_X1 U7406 ( .A1(n10976), .A2(n9735), .ZN(n10199) );
  NOR2_X1 U7407 ( .A1(n7087), .A2(n13207), .ZN(n7086) );
  INV_X1 U7408 ( .A(n13205), .ZN(n7087) );
  AND4_X1 U7409 ( .A1(n9225), .A2(n9224), .A3(n9223), .A4(n9222), .ZN(n13764)
         );
  AOI21_X1 U7410 ( .B1(n7361), .B2(n7359), .A(n7358), .ZN(n13940) );
  NOR2_X1 U7411 ( .A1(n7363), .A2(n7360), .ZN(n7359) );
  OAI21_X1 U7412 ( .B1(n7362), .B2(n7360), .A(n6495), .ZN(n7358) );
  INV_X1 U7413 ( .A(n13988), .ZN(n7361) );
  NOR2_X1 U7414 ( .A1(n13958), .A2(n7397), .ZN(n7396) );
  NAND2_X1 U7415 ( .A1(n13909), .A2(n13908), .ZN(n14142) );
  NAND2_X1 U7416 ( .A1(n6940), .A2(n9448), .ZN(n9041) );
  INV_X1 U7417 ( .A(n9091), .ZN(n7464) );
  OAI21_X1 U7418 ( .B1(n7768), .B2(n10355), .A(n7769), .ZN(n7770) );
  NAND2_X1 U7419 ( .A1(n9078), .A2(n9079), .ZN(n6859) );
  NOR2_X1 U7420 ( .A1(n9078), .A2(n9079), .ZN(n6858) );
  INV_X1 U7421 ( .A(n9080), .ZN(n6857) );
  AOI22_X1 U7422 ( .A1(n14831), .A2(n8298), .B1(n8284), .B2(n13105), .ZN(n7858) );
  OR2_X1 U7423 ( .A1(n6862), .A2(n6865), .ZN(n6861) );
  NOR2_X1 U7424 ( .A1(n9197), .A2(n6416), .ZN(n6862) );
  AOI21_X1 U7425 ( .B1(n7591), .B2(n6409), .A(n6760), .ZN(n6759) );
  INV_X1 U7426 ( .A(n8035), .ZN(n6760) );
  AOI22_X1 U7427 ( .A1(n14511), .A2(n8284), .B1(n8298), .B2(n13101), .ZN(n8035) );
  NAND2_X1 U7428 ( .A1(n6443), .A2(n7589), .ZN(n7592) );
  AND2_X1 U7429 ( .A1(n6905), .A2(n9250), .ZN(n6907) );
  AOI21_X1 U7430 ( .B1(n9248), .B2(n9247), .A(n6906), .ZN(n6905) );
  AND2_X1 U7431 ( .A1(n8139), .A2(n8141), .ZN(n7566) );
  INV_X1 U7432 ( .A(n8191), .ZN(n7581) );
  AND2_X1 U7433 ( .A1(n9369), .A2(n6849), .ZN(n6848) );
  AOI22_X1 U7434 ( .A1(n13313), .A2(n8242), .B1(n8298), .B2(n13247), .ZN(n8170) );
  INV_X1 U7435 ( .A(n7574), .ZN(n7572) );
  AOI21_X1 U7436 ( .B1(n7580), .B2(n7579), .A(n8207), .ZN(n7578) );
  NOR2_X1 U7437 ( .A1(n12552), .A2(n12551), .ZN(n12553) );
  OR2_X1 U7438 ( .A1(n12634), .A2(n12641), .ZN(n12397) );
  INV_X1 U7439 ( .A(n7171), .ZN(n7170) );
  OAI22_X1 U7440 ( .A1(n12670), .A2(n6445), .B1(n12691), .B2(n12859), .ZN(
        n7171) );
  OR2_X1 U7441 ( .A1(n12667), .A2(n12676), .ZN(n12382) );
  OR2_X1 U7442 ( .A1(n12880), .A2(n12726), .ZN(n12350) );
  AOI21_X1 U7443 ( .B1(n11570), .B2(n12300), .A(n6408), .ZN(n7517) );
  NOR2_X1 U7444 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_16__SCAN_IN), .ZN(
        n8349) );
  NAND2_X1 U7445 ( .A1(n9547), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8460) );
  NAND2_X1 U7446 ( .A1(n9538), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8440) );
  AND2_X1 U7447 ( .A1(n12034), .A2(n13058), .ZN(n6677) );
  OR2_X1 U7448 ( .A1(n12034), .A2(n13058), .ZN(n6678) );
  INV_X1 U7449 ( .A(n13244), .ZN(n7276) );
  NOR2_X1 U7450 ( .A1(n11657), .A2(n7082), .ZN(n7081) );
  INV_X1 U7451 ( .A(n11655), .ZN(n7082) );
  OR2_X1 U7452 ( .A1(n14696), .A2(n11364), .ZN(n11361) );
  NOR2_X1 U7453 ( .A1(n13430), .A2(n6692), .ZN(n6691) );
  INV_X1 U7454 ( .A(n11827), .ZN(n6692) );
  NAND2_X1 U7455 ( .A1(n9737), .A2(n11396), .ZN(n9865) );
  NAND2_X1 U7456 ( .A1(n8286), .A2(n9737), .ZN(n9864) );
  NOR2_X1 U7457 ( .A1(n7659), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n8306) );
  AND2_X1 U7458 ( .A1(n7958), .A2(n7957), .ZN(n7974) );
  XNOR2_X1 U7459 ( .A(n14179), .B(n13962), .ZN(n13902) );
  INV_X1 U7460 ( .A(n14067), .ZN(n6815) );
  OR2_X1 U7461 ( .A1(n13887), .A2(n13686), .ZN(n13908) );
  NAND2_X1 U7462 ( .A1(n6962), .A2(n9505), .ZN(n9817) );
  AND2_X1 U7463 ( .A1(n7444), .A2(n9007), .ZN(n6962) );
  NAND2_X1 U7464 ( .A1(n11214), .A2(n7356), .ZN(n14616) );
  AND2_X1 U7465 ( .A1(n11215), .A2(n11213), .ZN(n7356) );
  AND2_X1 U7466 ( .A1(n7219), .A2(n7218), .ZN(n8966) );
  NAND2_X1 U7467 ( .A1(n7033), .A2(n8174), .ZN(n8194) );
  INV_X1 U7468 ( .A(n8021), .ZN(n7025) );
  XNOR2_X1 U7469 ( .A(n8011), .B(SI_16_), .ZN(n8021) );
  AOI21_X1 U7470 ( .B1(n6577), .B2(n6580), .A(n6574), .ZN(n6573) );
  NAND2_X1 U7471 ( .A1(n7890), .A2(n6577), .ZN(n6575) );
  AND2_X1 U7472 ( .A1(n7028), .A2(n6578), .ZN(n6577) );
  INV_X1 U7473 ( .A(n7841), .ZN(n7412) );
  NAND2_X1 U7474 ( .A1(n6840), .A2(n7820), .ZN(n6839) );
  NAND2_X1 U7475 ( .A1(n7795), .A2(SI_6_), .ZN(n7820) );
  INV_X1 U7476 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n8968) );
  AOI21_X1 U7477 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n14336), .A(n14335), .ZN(
        n14395) );
  NOR2_X1 U7478 ( .A1(n14353), .A2(n14352), .ZN(n14335) );
  INV_X1 U7479 ( .A(n7317), .ZN(n7316) );
  OAI21_X1 U7480 ( .B1(n12165), .B2(n7318), .A(n7324), .ZN(n7317) );
  NAND2_X1 U7481 ( .A1(n7320), .A2(n7322), .ZN(n7318) );
  INV_X1 U7482 ( .A(n12165), .ZN(n7319) );
  NOR2_X1 U7483 ( .A1(n10376), .A2(n6916), .ZN(n7333) );
  INV_X1 U7484 ( .A(n10370), .ZN(n6916) );
  OR2_X1 U7485 ( .A1(n11076), .A2(n7336), .ZN(n7335) );
  INV_X1 U7486 ( .A(n11374), .ZN(n7336) );
  CLKBUF_X1 U7487 ( .A(n10710), .Z(n8380) );
  NAND2_X1 U7488 ( .A1(n6600), .A2(n6599), .ZN(n6598) );
  INV_X1 U7489 ( .A(n15003), .ZN(n6599) );
  OR2_X1 U7490 ( .A1(n11696), .A2(n11697), .ZN(n7270) );
  OR2_X1 U7491 ( .A1(n12388), .A2(n12652), .ZN(n8876) );
  NAND2_X1 U7492 ( .A1(n7539), .A2(n12383), .ZN(n7538) );
  INV_X1 U7493 ( .A(n7541), .ZN(n7539) );
  INV_X1 U7494 ( .A(n12649), .ZN(n12647) );
  OR2_X1 U7495 ( .A1(n12684), .A2(n12691), .ZN(n12378) );
  OAI21_X1 U7496 ( .B1(n8698), .B2(n7545), .A(n7543), .ZN(n12704) );
  INV_X1 U7497 ( .A(n7546), .ZN(n7545) );
  AOI21_X1 U7498 ( .B1(n7546), .B2(n12362), .A(n7544), .ZN(n7543) );
  INV_X1 U7499 ( .A(n12366), .ZN(n7544) );
  AOI21_X1 U7500 ( .B1(n7193), .B2(n12756), .A(n6489), .ZN(n7192) );
  NAND2_X1 U7501 ( .A1(n6884), .A2(n7193), .ZN(n6883) );
  AOI21_X1 U7502 ( .B1(n8865), .B2(n6568), .A(n6535), .ZN(n6567) );
  INV_X1 U7503 ( .A(n8865), .ZN(n6569) );
  AND4_X1 U7504 ( .A1(n8576), .A2(n8575), .A3(n8574), .A4(n8573), .ZN(n12820)
         );
  NAND2_X1 U7505 ( .A1(n11148), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8573) );
  NAND2_X1 U7506 ( .A1(n11239), .A2(n6571), .ZN(n11568) );
  AND2_X1 U7507 ( .A1(n11570), .A2(n8859), .ZN(n6571) );
  NAND2_X1 U7508 ( .A1(n11035), .A2(n8857), .ZN(n11115) );
  NAND2_X1 U7509 ( .A1(n10530), .A2(n8854), .ZN(n10533) );
  NAND2_X1 U7510 ( .A1(n8847), .A2(n12402), .ZN(n15046) );
  INV_X1 U7511 ( .A(n12213), .ZN(n8687) );
  NAND2_X1 U7512 ( .A1(n6793), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6792) );
  OAI21_X1 U7513 ( .B1(n11849), .B2(n11848), .A(n11847), .ZN(n11853) );
  AND2_X1 U7514 ( .A1(n8363), .A2(n6793), .ZN(n8365) );
  MUX2_X1 U7515 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8362), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n8363) );
  NAND2_X1 U7516 ( .A1(n7549), .A2(n7550), .ZN(n8361) );
  NAND2_X1 U7517 ( .A1(n7149), .A2(n7150), .ZN(n8923) );
  AOI21_X1 U7518 ( .B1(n7151), .B2(n8807), .A(n6562), .ZN(n7150) );
  INV_X1 U7519 ( .A(n8765), .ZN(n7153) );
  NAND2_X1 U7520 ( .A1(n8714), .A2(n8713), .ZN(n8733) );
  NAND2_X1 U7521 ( .A1(n7120), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8713) );
  NAND2_X1 U7522 ( .A1(n8702), .A2(n8701), .ZN(n7120) );
  NAND2_X1 U7523 ( .A1(n8700), .A2(n6657), .ZN(n7119) );
  AND2_X1 U7524 ( .A1(n8699), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6657) );
  INV_X1 U7525 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8685) );
  NAND2_X1 U7526 ( .A1(n8632), .A2(n8631), .ZN(n8635) );
  INV_X1 U7527 ( .A(n7115), .ZN(n7114) );
  OAI21_X1 U7528 ( .B1(n8593), .B2(n7116), .A(n8609), .ZN(n7115) );
  INV_X1 U7529 ( .A(n8596), .ZN(n7116) );
  AND4_X1 U7530 ( .A1(n8345), .A2(n8479), .A3(n8344), .A4(n8516), .ZN(n8346)
         );
  NOR2_X1 U7531 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_8__SCAN_IN), .ZN(
        n8345) );
  AND2_X1 U7532 ( .A1(n8547), .A2(n8530), .ZN(n8545) );
  NAND2_X1 U7533 ( .A1(n9603), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8528) );
  NAND2_X1 U7534 ( .A1(n8512), .A2(n8511), .ZN(n8529) );
  NAND2_X1 U7535 ( .A1(n8473), .A2(n8472), .ZN(n7148) );
  NAND2_X1 U7536 ( .A1(n8427), .A2(n8426), .ZN(n8439) );
  AOI21_X1 U7537 ( .B1(n7052), .B2(n12051), .A(n6447), .ZN(n7051) );
  OR2_X1 U7538 ( .A1(n13021), .A2(n13024), .ZN(n13022) );
  NAND2_X1 U7539 ( .A1(n7914), .A2(n7913), .ZN(n11359) );
  NAND2_X1 U7540 ( .A1(n6746), .A2(n7555), .ZN(n7554) );
  AND2_X1 U7541 ( .A1(n8271), .A2(n7558), .ZN(n7555) );
  AOI21_X1 U7542 ( .B1(n7567), .B2(n6411), .A(n6744), .ZN(n6746) );
  AND2_X1 U7543 ( .A1(n8119), .A2(n8118), .ZN(n13239) );
  INV_X1 U7544 ( .A(n13211), .ZN(n6593) );
  NOR2_X1 U7545 ( .A1(n13254), .A2(n7285), .ZN(n7284) );
  INV_X1 U7546 ( .A(n13251), .ZN(n7285) );
  AOI21_X1 U7547 ( .B1(n7284), .B2(n7084), .A(n7283), .ZN(n7282) );
  NOR2_X1 U7548 ( .A1(n13460), .A2(n13253), .ZN(n7283) );
  INV_X1 U7549 ( .A(n13291), .ZN(n7063) );
  NAND2_X1 U7550 ( .A1(n13478), .A2(n13248), .ZN(n13309) );
  NAND2_X1 U7551 ( .A1(n6587), .A2(n13203), .ZN(n13326) );
  XNOR2_X1 U7552 ( .A(n13313), .B(n13247), .ZN(n13321) );
  NAND2_X1 U7553 ( .A1(n13371), .A2(n13567), .ZN(n13359) );
  NOR2_X1 U7554 ( .A1(n13236), .A2(n6703), .ZN(n6702) );
  INV_X1 U7555 ( .A(n13234), .ZN(n6703) );
  OAI21_X1 U7556 ( .B1(n13227), .B2(n7288), .A(n7286), .ZN(n13388) );
  INV_X1 U7557 ( .A(n7289), .ZN(n7288) );
  AOI21_X1 U7558 ( .B1(n7289), .B2(n7287), .A(n6423), .ZN(n7286) );
  NAND2_X1 U7559 ( .A1(n13227), .A2(n13226), .ZN(n7291) );
  NAND2_X1 U7560 ( .A1(n11051), .A2(n11050), .ZN(n11207) );
  AND2_X2 U7561 ( .A1(n9737), .A2(n7504), .ZN(n13390) );
  AND2_X1 U7562 ( .A1(n7505), .A2(n11396), .ZN(n7504) );
  INV_X1 U7563 ( .A(n13183), .ZN(n13261) );
  AND2_X1 U7564 ( .A1(n6582), .A2(n6581), .ZN(n14540) );
  INV_X1 U7565 ( .A(n7996), .ZN(n6581) );
  NAND2_X1 U7566 ( .A1(n10386), .A2(n7910), .ZN(n6582) );
  NAND2_X2 U7567 ( .A1(n7685), .A2(n9525), .ZN(n8277) );
  NOR2_X2 U7568 ( .A1(n7637), .A2(n7638), .ZN(n7641) );
  INV_X1 U7569 ( .A(n7636), .ZN(n7637) );
  MUX2_X1 U7570 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7635), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n7636) );
  AND4_X1 U7571 ( .A1(n7627), .A2(n7626), .A3(n7625), .A4(n7666), .ZN(n7628)
         );
  INV_X1 U7572 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7627) );
  INV_X1 U7573 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n7626) );
  NAND2_X1 U7574 ( .A1(n7615), .A2(n7614), .ZN(n7616) );
  INV_X1 U7575 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n7615) );
  INV_X1 U7576 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n7614) );
  INV_X1 U7577 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n7622) );
  NAND2_X1 U7578 ( .A1(n6713), .A2(n6908), .ZN(n13625) );
  INV_X1 U7579 ( .A(n13628), .ZN(n6908) );
  NAND2_X1 U7580 ( .A1(n13694), .A2(n6463), .ZN(n6723) );
  AOI21_X1 U7581 ( .B1(n7248), .B2(n7250), .A(n6488), .ZN(n6721) );
  INV_X2 U7582 ( .A(n9433), .ZN(n9428) );
  NOR2_X1 U7583 ( .A1(n14297), .A2(n14301), .ZN(n6706) );
  NAND2_X1 U7584 ( .A1(n9425), .A2(n9424), .ZN(n13931) );
  NAND2_X1 U7585 ( .A1(n9398), .A2(n9397), .ZN(n14171) );
  NAND2_X1 U7586 ( .A1(n13977), .A2(n13982), .ZN(n13976) );
  OR2_X1 U7587 ( .A1(n14193), .A2(n13921), .ZN(n6651) );
  NAND2_X1 U7588 ( .A1(n9279), .A2(n9278), .ZN(n14086) );
  NAND2_X1 U7589 ( .A1(n13891), .A2(n6845), .ZN(n6844) );
  AND2_X1 U7590 ( .A1(n13890), .A2(n6454), .ZN(n6845) );
  NAND2_X1 U7591 ( .A1(n11546), .A2(n7349), .ZN(n7348) );
  NOR2_X1 U7592 ( .A1(n11723), .A2(n7350), .ZN(n7349) );
  INV_X1 U7593 ( .A(n11545), .ZN(n7350) );
  XNOR2_X1 U7594 ( .A(n14562), .B(n13666), .ZN(n11550) );
  INV_X1 U7595 ( .A(n11279), .ZN(n11317) );
  XNOR2_X1 U7596 ( .A(n11312), .B(n11407), .ZN(n11020) );
  AOI21_X1 U7597 ( .B1(n10084), .B2(n10083), .A(n7598), .ZN(n10634) );
  INV_X1 U7598 ( .A(n14102), .ZN(n14135) );
  AOI21_X1 U7599 ( .B1(n13972), .B2(n13904), .A(n7360), .ZN(n13959) );
  INV_X1 U7600 ( .A(n9819), .ZN(n9809) );
  NAND2_X1 U7601 ( .A1(n9821), .A2(n9820), .ZN(n14245) );
  OR2_X1 U7602 ( .A1(n8274), .A2(n8273), .ZN(n8276) );
  NAND2_X1 U7603 ( .A1(n7825), .A2(n7824), .ZN(n7842) );
  INV_X1 U7604 ( .A(n12684), .ZN(n12859) );
  INV_X1 U7605 ( .A(n12714), .ZN(n12690) );
  NAND2_X1 U7606 ( .A1(n10037), .A2(n9740), .ZN(n10100) );
  XNOR2_X1 U7607 ( .A(n6957), .B(n13174), .ZN(n7605) );
  NAND2_X1 U7608 ( .A1(n7435), .A2(n6958), .ZN(n6957) );
  NAND2_X1 U7609 ( .A1(n9410), .A2(n9409), .ZN(n14167) );
  NAND2_X1 U7610 ( .A1(n6946), .A2(n7673), .ZN(n6731) );
  OAI21_X1 U7611 ( .B1(n7438), .B2(n7437), .A(n9069), .ZN(n9080) );
  MUX2_X1 U7612 ( .A(n9068), .B(n10514), .S(n9448), .Z(n9069) );
  OR2_X1 U7613 ( .A1(n9093), .A2(n7464), .ZN(n7463) );
  INV_X1 U7614 ( .A(n7771), .ZN(n7588) );
  INV_X1 U7615 ( .A(n7792), .ZN(n6974) );
  NAND2_X1 U7616 ( .A1(n7449), .A2(n9121), .ZN(n7448) );
  INV_X1 U7617 ( .A(n9122), .ZN(n7449) );
  OR2_X1 U7618 ( .A1(n7471), .A2(n9150), .ZN(n7469) );
  INV_X1 U7619 ( .A(n9131), .ZN(n6855) );
  NAND2_X1 U7620 ( .A1(n7840), .A2(n6459), .ZN(n7596) );
  OR2_X1 U7621 ( .A1(n7840), .A2(n6459), .ZN(n7595) );
  NAND2_X1 U7622 ( .A1(n9184), .A2(n7455), .ZN(n7454) );
  INV_X1 U7623 ( .A(n9196), .ZN(n6866) );
  NAND2_X1 U7624 ( .A1(n7904), .A2(n6461), .ZN(n7593) );
  AND2_X1 U7625 ( .A1(n7926), .A2(n6755), .ZN(n6754) );
  INV_X1 U7626 ( .A(n7924), .ZN(n6755) );
  NAND2_X1 U7627 ( .A1(n7924), .A2(n7927), .ZN(n6753) );
  INV_X1 U7628 ( .A(n9265), .ZN(n6948) );
  NOR2_X1 U7629 ( .A1(n9266), .A2(n9486), .ZN(n6949) );
  NAND2_X1 U7630 ( .A1(n7592), .A2(n6759), .ZN(n6758) );
  AND2_X1 U7631 ( .A1(n8034), .A2(n6757), .ZN(n6756) );
  NAND2_X1 U7632 ( .A1(n6759), .A2(n6761), .ZN(n6757) );
  OAI21_X1 U7633 ( .B1(n7592), .B2(n6485), .A(n6415), .ZN(n7987) );
  OAI21_X1 U7634 ( .B1(n6734), .B2(n6733), .A(n7597), .ZN(n8100) );
  NAND2_X1 U7635 ( .A1(n8084), .A2(n8086), .ZN(n7597) );
  NAND2_X1 U7636 ( .A1(n9315), .A2(n7468), .ZN(n7467) );
  INV_X1 U7637 ( .A(n9302), .ZN(n6893) );
  OAI21_X1 U7638 ( .B1(n7458), .B2(n7457), .A(n7459), .ZN(n9353) );
  NAND2_X1 U7639 ( .A1(n9339), .A2(n9341), .ZN(n7459) );
  NOR2_X1 U7640 ( .A1(n7577), .A2(n7582), .ZN(n7573) );
  NAND2_X1 U7641 ( .A1(n9387), .A2(n7451), .ZN(n7450) );
  INV_X1 U7642 ( .A(n9386), .ZN(n7451) );
  NAND2_X1 U7643 ( .A1(n9817), .A2(n7443), .ZN(n9445) );
  NAND2_X1 U7644 ( .A1(n9816), .A2(n14008), .ZN(n7443) );
  INV_X1 U7645 ( .A(n8087), .ZN(n7404) );
  NOR2_X1 U7646 ( .A1(n8088), .A2(n8069), .ZN(n7405) );
  NAND2_X1 U7647 ( .A1(n7506), .A2(n6395), .ZN(n12270) );
  INV_X1 U7648 ( .A(n8850), .ZN(n7506) );
  INV_X1 U7649 ( .A(n8169), .ZN(n6921) );
  AND2_X1 U7650 ( .A1(n7563), .A2(n7561), .ZN(n8157) );
  INV_X1 U7651 ( .A(n7573), .ZN(n7571) );
  AND2_X1 U7652 ( .A1(n7573), .A2(n7580), .ZN(n7569) );
  AOI21_X1 U7653 ( .B1(n7578), .B2(n7577), .A(n7575), .ZN(n7574) );
  INV_X1 U7654 ( .A(n8206), .ZN(n7575) );
  OR2_X1 U7655 ( .A1(n8267), .A2(n8268), .ZN(n6747) );
  INV_X1 U7656 ( .A(n7651), .ZN(n6971) );
  NOR2_X1 U7657 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n6970) );
  NOR2_X1 U7658 ( .A1(n13974), .A2(n7365), .ZN(n7364) );
  AND2_X1 U7659 ( .A1(n7366), .A2(n13994), .ZN(n7365) );
  INV_X1 U7660 ( .A(n7367), .ZN(n7366) );
  NAND2_X1 U7661 ( .A1(n6579), .A2(n7907), .ZN(n6578) );
  INV_X1 U7662 ( .A(n6835), .ZN(n6579) );
  OAI21_X1 U7663 ( .B1(n6835), .B2(n6580), .A(n7928), .ZN(n6834) );
  NAND2_X1 U7664 ( .A1(n7035), .A2(SI_3_), .ZN(n7751) );
  NOR2_X1 U7665 ( .A1(n14323), .A2(n14322), .ZN(n14325) );
  NOR2_X1 U7666 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n14383), .ZN(n14322) );
  NAND2_X1 U7667 ( .A1(n12412), .A2(n12409), .ZN(n7129) );
  AOI21_X1 U7668 ( .B1(n7510), .B2(n7508), .A(n12399), .ZN(n7507) );
  INV_X1 U7669 ( .A(n7513), .ZN(n7508) );
  NOR2_X1 U7670 ( .A1(n12628), .A2(n7514), .ZN(n7513) );
  INV_X1 U7671 ( .A(n8876), .ZN(n7514) );
  INV_X1 U7672 ( .A(n12373), .ZN(n7167) );
  NAND2_X1 U7673 ( .A1(n7173), .A2(n7175), .ZN(n7172) );
  OR2_X1 U7674 ( .A1(n12694), .A2(n12702), .ZN(n12250) );
  OR2_X1 U7675 ( .A1(n8705), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8720) );
  NAND2_X1 U7676 ( .A1(n8656), .A2(n15169), .ZN(n8672) );
  NAND2_X1 U7677 ( .A1(n8871), .A2(n8870), .ZN(n6884) );
  NAND2_X1 U7678 ( .A1(n7185), .A2(n7183), .ZN(n8871) );
  NOR2_X1 U7679 ( .A1(n8869), .A2(n7184), .ZN(n7183) );
  NOR2_X1 U7680 ( .A1(n12776), .A2(n7528), .ZN(n7527) );
  AND2_X1 U7681 ( .A1(n12788), .A2(n12334), .ZN(n7528) );
  INV_X1 U7682 ( .A(n12334), .ZN(n7525) );
  OR2_X1 U7683 ( .A1(n12439), .A2(n14493), .ZN(n12318) );
  INV_X1 U7684 ( .A(n12300), .ZN(n7518) );
  INV_X1 U7685 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8354) );
  AND2_X1 U7686 ( .A1(n8353), .A2(n8533), .ZN(n8355) );
  NAND2_X1 U7687 ( .A1(n9580), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8490) );
  NAND2_X1 U7688 ( .A1(n9523), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8426) );
  INV_X1 U7689 ( .A(n12013), .ZN(n7044) );
  INV_X1 U7690 ( .A(n7485), .ZN(n7484) );
  AND2_X1 U7691 ( .A1(n13032), .A2(n7495), .ZN(n7494) );
  NAND2_X1 U7692 ( .A1(n13024), .A2(n12007), .ZN(n7495) );
  AND2_X1 U7693 ( .A1(n8322), .A2(n13332), .ZN(n6956) );
  NAND2_X1 U7694 ( .A1(n6701), .A2(n6700), .ZN(n13241) );
  AND2_X1 U7695 ( .A1(n13355), .A2(n13238), .ZN(n6700) );
  NOR2_X1 U7696 ( .A1(n7094), .A2(n7093), .ZN(n7092) );
  INV_X1 U7697 ( .A(n10791), .ZN(n7093) );
  INV_X1 U7698 ( .A(n10789), .ZN(n7094) );
  INV_X1 U7699 ( .A(n13252), .ZN(n13253) );
  NAND2_X1 U7700 ( .A1(n6694), .A2(n11657), .ZN(n6693) );
  INV_X1 U7701 ( .A(n10052), .ZN(n10188) );
  INV_X1 U7702 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n7666) );
  AND2_X1 U7703 ( .A1(n7934), .A2(n7933), .ZN(n7958) );
  INV_X1 U7704 ( .A(n9841), .ZN(n9845) );
  INV_X1 U7705 ( .A(n7229), .ZN(n7228) );
  NOR2_X1 U7706 ( .A1(n13931), .A2(n14167), .ZN(n7209) );
  INV_X1 U7707 ( .A(n7378), .ZN(n7377) );
  OAI21_X1 U7708 ( .B1(n10828), .B2(n7379), .A(n11020), .ZN(n7378) );
  INV_X1 U7709 ( .A(n11015), .ZN(n7379) );
  INV_X1 U7710 ( .A(n13773), .ZN(n13923) );
  NAND2_X1 U7711 ( .A1(n14098), .A2(n13912), .ZN(n14100) );
  INV_X1 U7712 ( .A(n13634), .ZN(n6824) );
  INV_X1 U7713 ( .A(n14294), .ZN(n9531) );
  INV_X1 U7714 ( .A(n8193), .ZN(n7429) );
  XNOR2_X1 U7715 ( .A(n8160), .B(n8159), .ZN(n8158) );
  AND2_X1 U7716 ( .A1(n9006), .A2(n9005), .ZN(n7444) );
  NAND2_X1 U7717 ( .A1(n8995), .A2(n6934), .ZN(n9007) );
  NOR2_X1 U7718 ( .A1(n9004), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n6934) );
  INV_X1 U7719 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n7476) );
  INV_X1 U7720 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n7475) );
  INV_X1 U7721 ( .A(n7024), .ZN(n7023) );
  OAI21_X1 U7722 ( .B1(n8009), .B2(n7025), .A(n8012), .ZN(n7024) );
  NAND2_X1 U7723 ( .A1(n7867), .A2(SI_9_), .ZN(n7889) );
  OR2_X1 U7724 ( .A1(n9118), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n9127) );
  XNOR2_X1 U7725 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n14363) );
  NAND2_X1 U7726 ( .A1(n14310), .A2(n6803), .ZN(n14312) );
  NAND2_X1 U7727 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n6804), .ZN(n6803) );
  NAND2_X1 U7728 ( .A1(n6805), .A2(n14316), .ZN(n14317) );
  NAND2_X1 U7729 ( .A1(n14357), .A2(n14358), .ZN(n6805) );
  XNOR2_X1 U7730 ( .A(n14317), .B(n6982), .ZN(n14372) );
  INV_X1 U7731 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n6982) );
  AOI22_X1 U7732 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14377), .B1(n14378), .B2(
        n14320), .ZN(n14321) );
  OR2_X1 U7733 ( .A1(n14377), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n14320) );
  XOR2_X1 U7734 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(n14325), .Z(n14386) );
  AOI21_X1 U7735 ( .B1(n15184), .B2(n14343), .A(n14342), .ZN(n14399) );
  INV_X1 U7736 ( .A(n11389), .ZN(n10884) );
  NAND2_X1 U7737 ( .A1(n12092), .A2(n12091), .ZN(n6783) );
  NAND2_X1 U7738 ( .A1(n11148), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8773) );
  OR2_X1 U7739 ( .A1(n8672), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8692) );
  XNOR2_X1 U7740 ( .A(n10229), .B(n12299), .ZN(n10910) );
  AND2_X1 U7741 ( .A1(n12147), .A2(n12765), .ZN(n6789) );
  NAND2_X1 U7742 ( .A1(n8769), .A2(n8768), .ZN(n8783) );
  INV_X1 U7743 ( .A(n8770), .ZN(n8769) );
  NAND2_X1 U7744 ( .A1(n6500), .A2(n7325), .ZN(n7320) );
  NAND2_X1 U7745 ( .A1(n12178), .A2(n7326), .ZN(n7323) );
  NAND2_X1 U7746 ( .A1(n7304), .A2(n14471), .ZN(n11455) );
  INV_X1 U7747 ( .A(n11380), .ZN(n7304) );
  OR2_X1 U7748 ( .A1(n8522), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8539) );
  OR2_X1 U7749 ( .A1(n12148), .A2(n12153), .ZN(n6788) );
  NOR2_X1 U7750 ( .A1(n8906), .A2(n12958), .ZN(n10224) );
  NOR2_X1 U7751 ( .A1(n7262), .A2(n15081), .ZN(n7259) );
  INV_X1 U7752 ( .A(n6913), .ZN(n10718) );
  INV_X1 U7753 ( .A(n11463), .ZN(n11476) );
  NAND2_X1 U7754 ( .A1(n7257), .A2(n7256), .ZN(n10711) );
  OR2_X1 U7755 ( .A1(n11463), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7257) );
  AND2_X1 U7756 ( .A1(n6989), .A2(n7258), .ZN(n10712) );
  AOI21_X1 U7757 ( .B1(n7259), .B2(n10841), .A(n7262), .ZN(n7258) );
  NAND2_X1 U7758 ( .A1(n6913), .A2(n7259), .ZN(n6989) );
  NOR2_X1 U7759 ( .A1(n10712), .A2(n10711), .ZN(n11462) );
  OR2_X1 U7760 ( .A1(n11462), .A2(n7002), .ZN(n7001) );
  AND2_X1 U7761 ( .A1(n11463), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7002) );
  INV_X1 U7762 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n10378) );
  NAND2_X1 U7763 ( .A1(n14880), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7272) );
  NAND2_X1 U7764 ( .A1(n6603), .A2(n11465), .ZN(n6601) );
  NAND2_X1 U7765 ( .A1(n14853), .A2(n6603), .ZN(n6602) );
  OR2_X1 U7766 ( .A1(n14912), .A2(n14911), .ZN(n7264) );
  AND2_X1 U7767 ( .A1(n7264), .A2(n7263), .ZN(n11468) );
  NAND2_X1 U7768 ( .A1(n14919), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7263) );
  INV_X1 U7769 ( .A(n14949), .ZN(n7265) );
  OR2_X1 U7770 ( .A1(n14968), .A2(n11471), .ZN(n6600) );
  NAND2_X1 U7771 ( .A1(n11472), .A2(n11700), .ZN(n11695) );
  OAI21_X1 U7772 ( .B1(n12454), .B2(n14492), .A(n12453), .ZN(n12475) );
  NAND2_X1 U7773 ( .A1(n12456), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7267) );
  OR2_X1 U7774 ( .A1(n12474), .A2(n12485), .ZN(n6604) );
  NAND2_X1 U7775 ( .A1(n6604), .A2(n12507), .ZN(n12520) );
  NAND2_X1 U7776 ( .A1(n12637), .A2(n7513), .ZN(n7512) );
  OR2_X1 U7777 ( .A1(n12628), .A2(n12395), .ZN(n7511) );
  NAND2_X1 U7778 ( .A1(n12248), .A2(n8791), .ZN(n12649) );
  NOR2_X1 U7779 ( .A1(n12659), .A2(n7542), .ZN(n7541) );
  INV_X1 U7780 ( .A(n12378), .ZN(n7542) );
  NAND2_X1 U7781 ( .A1(n12382), .A2(n12383), .ZN(n12659) );
  NAND2_X1 U7782 ( .A1(n12671), .A2(n12670), .ZN(n12673) );
  NAND2_X1 U7783 ( .A1(n12712), .A2(n12720), .ZN(n6572) );
  NAND2_X1 U7784 ( .A1(n8698), .A2(n8697), .ZN(n7548) );
  AOI21_X1 U7785 ( .B1(n7522), .B2(n8872), .A(n7520), .ZN(n7519) );
  INV_X1 U7786 ( .A(n7522), .ZN(n7521) );
  INV_X1 U7787 ( .A(n12350), .ZN(n7520) );
  AND3_X1 U7788 ( .A1(n8696), .A2(n8695), .A3(n8694), .ZN(n12742) );
  INV_X1 U7789 ( .A(n8873), .ZN(n7194) );
  AND2_X1 U7790 ( .A1(n12350), .A2(n12355), .ZN(n12740) );
  NOR2_X1 U7791 ( .A1(n12735), .A2(n12354), .ZN(n7522) );
  INV_X1 U7792 ( .A(n12740), .ZN(n12735) );
  INV_X1 U7793 ( .A(n6884), .ZN(n12750) );
  NAND2_X1 U7794 ( .A1(n12750), .A2(n8872), .ZN(n12749) );
  NAND2_X1 U7795 ( .A1(n12757), .A2(n12756), .ZN(n12755) );
  AND2_X1 U7796 ( .A1(n12344), .A2(n12343), .ZN(n12767) );
  AND4_X1 U7797 ( .A1(n8608), .A2(n8607), .A3(n8606), .A4(n8605), .ZN(n12778)
         );
  AND2_X1 U7798 ( .A1(n12223), .A2(n12320), .ZN(n12806) );
  NAND2_X1 U7799 ( .A1(n12815), .A2(n8863), .ZN(n14465) );
  NAND2_X1 U7800 ( .A1(n11568), .A2(n7195), .ZN(n11614) );
  NOR2_X1 U7801 ( .A1(n12303), .A2(n7196), .ZN(n7195) );
  INV_X1 U7802 ( .A(n8860), .ZN(n7196) );
  NAND2_X1 U7803 ( .A1(n11566), .A2(n12297), .ZN(n11565) );
  NAND2_X1 U7804 ( .A1(n7181), .A2(n7179), .ZN(n11239) );
  AOI21_X1 U7805 ( .B1(n12226), .B2(n8858), .A(n7180), .ZN(n7179) );
  NAND2_X1 U7806 ( .A1(n12294), .A2(n12295), .ZN(n12227) );
  OR2_X1 U7807 ( .A1(n11115), .A2(n12226), .ZN(n11118) );
  AND4_X1 U7808 ( .A1(n8471), .A2(n8470), .A3(n8469), .A4(n8468), .ZN(n11231)
         );
  AND4_X1 U7809 ( .A1(n8456), .A2(n8455), .A3(n8454), .A4(n8453), .ZN(n11040)
         );
  AND2_X1 U7810 ( .A1(n8856), .A2(n8855), .ZN(n7197) );
  NAND2_X1 U7811 ( .A1(n11148), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8437) );
  NAND2_X1 U7812 ( .A1(n10393), .A2(n8853), .ZN(n10530) );
  NAND2_X1 U7813 ( .A1(n10755), .A2(n10378), .ZN(n8432) );
  AND2_X1 U7814 ( .A1(n12422), .A2(n12402), .ZN(n15067) );
  XNOR2_X1 U7815 ( .A(n8929), .B(n12222), .ZN(n8940) );
  NOR2_X1 U7816 ( .A1(n8938), .A2(n8937), .ZN(n8939) );
  AND2_X1 U7817 ( .A1(n8928), .A2(n8927), .ZN(n8957) );
  NAND2_X1 U7818 ( .A1(n8797), .A2(n8796), .ZN(n12388) );
  NAND2_X1 U7819 ( .A1(n8623), .A2(n8622), .ZN(n12337) );
  OR2_X1 U7820 ( .A1(n8637), .A2(n9562), .ZN(n8483) );
  INV_X1 U7821 ( .A(n11453), .ZN(n8907) );
  INV_X1 U7822 ( .A(n8834), .ZN(n7550) );
  AND2_X1 U7823 ( .A1(n7552), .A2(n8360), .ZN(n7549) );
  NAND2_X1 U7824 ( .A1(n8925), .A2(n8924), .ZN(n11849) );
  OR2_X1 U7825 ( .A1(n8923), .A2(n8922), .ZN(n8925) );
  INV_X1 U7826 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8360) );
  NAND2_X1 U7827 ( .A1(n6662), .A2(n8794), .ZN(n8808) );
  NAND2_X1 U7828 ( .A1(n8793), .A2(n8792), .ZN(n6662) );
  NOR2_X1 U7829 ( .A1(n8886), .A2(P3_IR_REG_22__SCAN_IN), .ZN(n8909) );
  NAND2_X1 U7830 ( .A1(n8909), .A2(n6772), .ZN(n8888) );
  AND2_X1 U7831 ( .A1(n8911), .A2(n6773), .ZN(n6772) );
  INV_X1 U7832 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n6773) );
  NAND2_X1 U7833 ( .A1(n8764), .A2(n8763), .ZN(n8765) );
  NAND2_X1 U7834 ( .A1(n6661), .A2(n8734), .ZN(n8748) );
  NAND2_X1 U7835 ( .A1(n8733), .A2(n8732), .ZN(n6661) );
  NAND2_X1 U7836 ( .A1(n8681), .A2(n8680), .ZN(n8700) );
  NAND2_X1 U7837 ( .A1(n8679), .A2(n8678), .ZN(n8681) );
  NAND2_X1 U7838 ( .A1(n6658), .A2(n7131), .ZN(n8679) );
  AOI21_X1 U7839 ( .B1(n7133), .B2(n7135), .A(n7132), .ZN(n7131) );
  NAND2_X1 U7840 ( .A1(n8635), .A2(n7133), .ZN(n6658) );
  INV_X1 U7841 ( .A(n8666), .ZN(n7132) );
  AND2_X1 U7842 ( .A1(n8650), .A2(n8633), .ZN(n8634) );
  NAND2_X1 U7843 ( .A1(n8635), .A2(n8634), .ZN(n8651) );
  AOI21_X1 U7844 ( .B1(n7114), .B2(n7116), .A(n7112), .ZN(n7111) );
  INV_X1 U7845 ( .A(n8612), .ZN(n7112) );
  NAND2_X1 U7846 ( .A1(n8580), .A2(n10060), .ZN(n8593) );
  NAND2_X1 U7847 ( .A1(n6653), .A2(n7107), .ZN(n8580) );
  AND2_X1 U7848 ( .A1(n8609), .A2(n8595), .ZN(n8596) );
  NAND2_X1 U7849 ( .A1(n8593), .A2(n6656), .ZN(n8581) );
  NAND2_X1 U7850 ( .A1(n6653), .A2(n6652), .ZN(n6656) );
  AND2_X1 U7851 ( .A1(n7107), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n6652) );
  OR2_X1 U7852 ( .A1(n8581), .A2(n10155), .ZN(n8594) );
  AND2_X1 U7853 ( .A1(n8578), .A2(n8560), .ZN(n8561) );
  AOI21_X1 U7854 ( .B1(n7139), .B2(n7141), .A(n7138), .ZN(n7137) );
  INV_X1 U7855 ( .A(n8547), .ZN(n7138) );
  NAND2_X1 U7856 ( .A1(n8550), .A2(n8549), .ZN(n8559) );
  AND2_X1 U7857 ( .A1(n8528), .A2(n8510), .ZN(n8511) );
  NAND2_X1 U7858 ( .A1(n8509), .A2(n8508), .ZN(n8512) );
  NAND2_X1 U7859 ( .A1(n8494), .A2(n8493), .ZN(n8509) );
  NOR2_X1 U7860 ( .A1(n8476), .A2(n7147), .ZN(n7146) );
  INV_X1 U7861 ( .A(n8474), .ZN(n7147) );
  NAND2_X1 U7862 ( .A1(n8461), .A2(n8460), .ZN(n8473) );
  AND2_X1 U7863 ( .A1(n8447), .A2(n8446), .ZN(n11499) );
  NAND2_X1 U7864 ( .A1(n8410), .A2(n8409), .ZN(n8425) );
  NOR2_X2 U7865 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n10710) );
  INV_X1 U7866 ( .A(n13066), .ZN(n7487) );
  AND2_X1 U7867 ( .A1(n12985), .A2(n6450), .ZN(n7485) );
  NAND2_X1 U7868 ( .A1(n13039), .A2(n7499), .ZN(n7498) );
  AND2_X1 U7869 ( .A1(n7500), .A2(n7501), .ZN(n7499) );
  INV_X1 U7870 ( .A(n13017), .ZN(n7500) );
  XNOR2_X1 U7871 ( .A(n10499), .B(n12048), .ZN(n10198) );
  OAI21_X1 U7872 ( .B1(n6671), .B2(n11997), .A(n6670), .ZN(n7496) );
  INV_X1 U7873 ( .A(n11996), .ZN(n6674) );
  INV_X1 U7874 ( .A(n6453), .ZN(n6667) );
  OAI21_X1 U7875 ( .B1(n7057), .B2(n6667), .A(n14689), .ZN(n6666) );
  NAND2_X1 U7876 ( .A1(n13004), .A2(n12033), .ZN(n12035) );
  AOI21_X1 U7877 ( .B1(n6684), .B2(n10951), .A(n6683), .ZN(n7479) );
  INV_X1 U7878 ( .A(n7481), .ZN(n6684) );
  INV_X1 U7879 ( .A(n10952), .ZN(n6683) );
  INV_X1 U7880 ( .A(n7056), .ZN(n7055) );
  OAI21_X1 U7881 ( .B1(n7058), .B2(n7057), .A(n11259), .ZN(n7056) );
  NAND2_X1 U7882 ( .A1(n7496), .A2(n7494), .ZN(n13030) );
  NAND2_X1 U7883 ( .A1(n7498), .A2(n7497), .ZN(n13084) );
  AND2_X1 U7884 ( .A1(n13085), .A2(n12044), .ZN(n7497) );
  AND4_X1 U7885 ( .A1(n8188), .A2(n8187), .A3(n8186), .A4(n8185), .ZN(n13250)
         );
  NAND2_X1 U7886 ( .A1(n6637), .A2(n6636), .ZN(n13150) );
  INV_X1 U7887 ( .A(n13138), .ZN(n6636) );
  NAND2_X1 U7888 ( .A1(n8197), .A2(n8196), .ZN(n13292) );
  NAND2_X1 U7889 ( .A1(n13601), .A2(n7910), .ZN(n8197) );
  AND2_X1 U7890 ( .A1(n13212), .A2(n13211), .ZN(n13289) );
  OR2_X1 U7891 ( .A1(n7089), .A2(n13207), .ZN(n7088) );
  AND2_X1 U7892 ( .A1(n13321), .A2(n7090), .ZN(n7089) );
  NAND2_X1 U7893 ( .A1(n6439), .A2(n13205), .ZN(n7090) );
  AOI21_X1 U7894 ( .B1(n13242), .B2(n7275), .A(n6417), .ZN(n7274) );
  NAND2_X1 U7895 ( .A1(n13349), .A2(n7275), .ZN(n7273) );
  NAND2_X1 U7896 ( .A1(n7277), .A2(n13351), .ZN(n13350) );
  NAND2_X1 U7897 ( .A1(n6584), .A2(n13200), .ZN(n13341) );
  NOR2_X1 U7898 ( .A1(n13201), .A2(n6586), .ZN(n6585) );
  NOR2_X1 U7899 ( .A1(n13399), .A2(n7290), .ZN(n7289) );
  INV_X1 U7900 ( .A(n13230), .ZN(n7290) );
  OAI21_X1 U7901 ( .B1(n6694), .B2(n6690), .A(n6688), .ZN(n13227) );
  INV_X1 U7902 ( .A(n6689), .ZN(n6688) );
  OAI21_X1 U7903 ( .B1(n11657), .B2(n6690), .A(n11828), .ZN(n6689) );
  INV_X1 U7904 ( .A(n7079), .ZN(n6592) );
  OAI21_X1 U7905 ( .B1(n11821), .B2(n7080), .A(n6493), .ZN(n7079) );
  OR2_X1 U7906 ( .A1(n13423), .A2(n13422), .ZN(n13424) );
  NOR2_X1 U7907 ( .A1(n11644), .A2(n14511), .ZN(n11667) );
  NAND2_X1 U7908 ( .A1(n11667), .A2(n14540), .ZN(n13423) );
  NAND2_X1 U7909 ( .A1(n11656), .A2(n7081), .ZN(n11822) );
  AOI21_X1 U7910 ( .B1(n11360), .B2(n7075), .A(n7074), .ZN(n7073) );
  INV_X1 U7911 ( .A(n11361), .ZN(n7074) );
  AND2_X1 U7912 ( .A1(n10792), .A2(n10791), .ZN(n7096) );
  OR2_X1 U7913 ( .A1(n10975), .A2(n10789), .ZN(n7097) );
  AND2_X1 U7914 ( .A1(n10782), .A2(n10780), .ZN(n6704) );
  OAI21_X1 U7915 ( .B1(n10476), .B2(n10544), .A(n6685), .ZN(n10540) );
  AOI21_X1 U7916 ( .B1(n10477), .B2(n6686), .A(n6484), .ZN(n6685) );
  INV_X1 U7917 ( .A(n10475), .ZN(n6686) );
  NAND2_X1 U7918 ( .A1(n10360), .A2(n10359), .ZN(n10476) );
  NAND2_X1 U7919 ( .A1(n6914), .A2(n13174), .ZN(n10976) );
  AOI21_X1 U7920 ( .B1(n13309), .B2(n6457), .A(n7280), .ZN(n13260) );
  OAI21_X1 U7921 ( .B1(n7282), .B2(n7281), .A(n6498), .ZN(n7280) );
  AND2_X1 U7922 ( .A1(n7062), .A2(n14830), .ZN(n7106) );
  NAND2_X1 U7923 ( .A1(n8163), .A2(n8162), .ZN(n13313) );
  NAND2_X1 U7924 ( .A1(n8017), .A2(n8016), .ZN(n13229) );
  AND2_X1 U7925 ( .A1(n9742), .A2(n13603), .ZN(n14820) );
  INV_X1 U7926 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8305) );
  OR2_X1 U7927 ( .A1(n8332), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n8335) );
  INV_X1 U7928 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7613) );
  INV_X1 U7929 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n7560) );
  INV_X1 U7930 ( .A(n7245), .ZN(n7244) );
  OAI21_X1 U7931 ( .B1(n7247), .B2(n7246), .A(n13723), .ZN(n7245) );
  INV_X1 U7932 ( .A(n11887), .ZN(n7246) );
  INV_X1 U7933 ( .A(n6712), .ZN(n6711) );
  OAI21_X1 U7934 ( .B1(n13750), .B2(n11975), .A(n13619), .ZN(n6712) );
  NAND2_X1 U7935 ( .A1(n10138), .A2(n10139), .ZN(n10145) );
  NOR2_X1 U7936 ( .A1(n13654), .A2(n7230), .ZN(n7229) );
  INV_X1 U7937 ( .A(n7234), .ZN(n7230) );
  AOI21_X1 U7938 ( .B1(n13760), .B2(n13761), .A(n7220), .ZN(n13683) );
  INV_X1 U7939 ( .A(n7249), .ZN(n7248) );
  OAI21_X1 U7940 ( .B1(n7250), .B2(n11288), .A(n11304), .ZN(n7249) );
  INV_X1 U7941 ( .A(n7251), .ZN(n7250) );
  NAND2_X1 U7942 ( .A1(n11683), .A2(n11682), .ZN(n11878) );
  NAND2_X1 U7943 ( .A1(n6870), .A2(n6873), .ZN(n9475) );
  INV_X1 U7944 ( .A(n6874), .ZN(n6873) );
  OAI21_X1 U7945 ( .B1(n6876), .B2(n6875), .A(n9453), .ZN(n6874) );
  INV_X1 U7946 ( .A(n9096), .ZN(n9438) );
  OR2_X1 U7947 ( .A1(n9036), .A2(n9046), .ZN(n9047) );
  OR2_X1 U7948 ( .A1(n14283), .A2(n9440), .ZN(n9442) );
  INV_X1 U7949 ( .A(n13902), .ZN(n13974) );
  NAND2_X1 U7950 ( .A1(n9365), .A2(n9364), .ZN(n13922) );
  NAND2_X1 U7951 ( .A1(n14201), .A2(n7387), .ZN(n7389) );
  NOR2_X1 U7952 ( .A1(n14001), .A2(n7391), .ZN(n7387) );
  NAND2_X1 U7953 ( .A1(n14012), .A2(n13921), .ZN(n7388) );
  XNOR2_X1 U7954 ( .A(n13922), .B(n13923), .ZN(n13994) );
  NOR2_X1 U7955 ( .A1(n13988), .A2(n13994), .ZN(n13987) );
  NOR2_X1 U7956 ( .A1(n14017), .A2(n6817), .ZN(n6814) );
  AOI21_X1 U7957 ( .B1(n14016), .B2(n13920), .A(n6648), .ZN(n14002) );
  AND2_X1 U7958 ( .A1(n14017), .A2(n13919), .ZN(n6648) );
  INV_X1 U7959 ( .A(n13901), .ZN(n14001) );
  NAND2_X1 U7960 ( .A1(n7371), .A2(n7369), .ZN(n14035) );
  NAND2_X1 U7961 ( .A1(n7370), .A2(n7373), .ZN(n7369) );
  INV_X1 U7962 ( .A(n7372), .ZN(n7370) );
  NAND2_X1 U7963 ( .A1(n6844), .A2(n6842), .ZN(n6846) );
  NOR2_X1 U7964 ( .A1(n13895), .A2(n6843), .ZN(n6842) );
  INV_X1 U7965 ( .A(n13893), .ZN(n6843) );
  AOI21_X1 U7966 ( .B1(n6404), .B2(n11553), .A(n6490), .ZN(n7392) );
  NAND2_X1 U7967 ( .A1(n7348), .A2(n6479), .ZN(n13909) );
  AND2_X1 U7968 ( .A1(n13908), .A2(n9479), .ZN(n11731) );
  AOI21_X1 U7969 ( .B1(n7343), .B2(n7346), .A(n6487), .ZN(n7341) );
  OAI21_X1 U7970 ( .B1(n11276), .B2(n13667), .A(n11275), .ZN(n11278) );
  NAND2_X1 U7971 ( .A1(n7342), .A2(n11274), .ZN(n11318) );
  NAND2_X1 U7972 ( .A1(n11273), .A2(n11272), .ZN(n7342) );
  NOR2_X1 U7973 ( .A1(n9152), .A2(n11408), .ZN(n9173) );
  NAND2_X1 U7974 ( .A1(n11019), .A2(n6476), .ZN(n11214) );
  INV_X1 U7975 ( .A(n11020), .ZN(n7357) );
  NAND2_X1 U7976 ( .A1(n6645), .A2(n6644), .ZN(n11019) );
  INV_X1 U7977 ( .A(n10828), .ZN(n6644) );
  INV_X1 U7978 ( .A(n10829), .ZN(n6645) );
  NAND2_X1 U7979 ( .A1(n6546), .A2(n6810), .ZN(n11028) );
  OAI21_X1 U7980 ( .B1(n10585), .B2(n6630), .A(n6628), .ZN(n10808) );
  INV_X1 U7981 ( .A(n6629), .ZN(n6628) );
  INV_X1 U7982 ( .A(n10516), .ZN(n6630) );
  NAND2_X1 U7983 ( .A1(n10585), .A2(n10584), .ZN(n10583) );
  INV_X1 U7984 ( .A(n14078), .ZN(n14133) );
  NAND2_X2 U7985 ( .A1(n6887), .A2(n6941), .ZN(n6940) );
  NAND2_X1 U7986 ( .A1(n9385), .A2(n9384), .ZN(n14179) );
  OR2_X1 U7987 ( .A1(n9852), .A2(n9851), .ZN(n14670) );
  NOR2_X1 U7988 ( .A1(n6424), .A2(n6561), .ZN(n7431) );
  NOR2_X1 U7989 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n7235) );
  XNOR2_X1 U7990 ( .A(n8258), .B(n8257), .ZN(n13591) );
  NAND2_X1 U7991 ( .A1(n7432), .A2(n8247), .ZN(n8258) );
  NOR2_X1 U7992 ( .A1(n8979), .A2(n9227), .ZN(n6620) );
  NAND3_X1 U7993 ( .A1(n7603), .A2(n7200), .A3(n7199), .ZN(n8982) );
  INV_X1 U7994 ( .A(n8970), .ZN(n7200) );
  INV_X1 U7995 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n6904) );
  INV_X1 U7996 ( .A(n8980), .ZN(n6902) );
  NOR2_X1 U7997 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n6901) );
  NAND2_X1 U7998 ( .A1(n9500), .A2(n6412), .ZN(n9511) );
  INV_X1 U7999 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6724) );
  NAND2_X1 U8000 ( .A1(n8997), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8998) );
  XNOR2_X1 U8001 ( .A(n8108), .B(n8107), .ZN(n11395) );
  NAND2_X1 U8002 ( .A1(n7007), .A2(SI_20_), .ZN(n8105) );
  OAI21_X1 U8003 ( .B1(n8068), .B2(n7407), .A(n8071), .ZN(n8089) );
  NAND2_X1 U8004 ( .A1(n8010), .A2(n8009), .ZN(n8022) );
  XNOR2_X1 U8005 ( .A(n7991), .B(n7990), .ZN(n10386) );
  NAND2_X1 U8006 ( .A1(n6576), .A2(n7907), .ZN(n7929) );
  NAND2_X1 U8007 ( .A1(n7890), .A2(n6835), .ZN(n6576) );
  AOI21_X1 U8008 ( .B1(n7410), .B2(n7412), .A(n7409), .ZN(n7408) );
  NAND2_X1 U8009 ( .A1(n7821), .A2(n7820), .ZN(n7825) );
  NAND2_X1 U8010 ( .A1(n7797), .A2(n7796), .ZN(n7821) );
  NOR2_X1 U8011 ( .A1(n14371), .A2(n15271), .ZN(n14374) );
  NOR2_X1 U8012 ( .A1(n14415), .A2(n14381), .ZN(n14384) );
  NOR2_X1 U8013 ( .A1(n14331), .A2(n14330), .ZN(n14355) );
  AND2_X1 U8014 ( .A1(n15202), .A2(n14356), .ZN(n14330) );
  NAND2_X1 U8015 ( .A1(n6975), .A2(n14576), .ZN(n14396) );
  OAI21_X1 U8016 ( .B1(n14578), .B2(n14577), .A(n6976), .ZN(n6975) );
  INV_X1 U8017 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n6976) );
  AOI21_X1 U8018 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n14339), .A(n14338), .ZN(
        n14349) );
  AND4_X1 U8019 ( .A1(n8630), .A2(n8629), .A3(n8628), .A4(n8627), .ZN(n12790)
         );
  AND2_X1 U8020 ( .A1(n8537), .A2(n8536), .ZN(n11604) );
  NAND2_X1 U8021 ( .A1(n8717), .A2(n8716), .ZN(n12705) );
  INV_X1 U8022 ( .A(n12438), .ZN(n14470) );
  AND2_X1 U8023 ( .A1(n8805), .A2(n8804), .ZN(n12652) );
  NAND2_X1 U8024 ( .A1(n8655), .A2(n8654), .ZN(n12348) );
  NAND2_X1 U8025 ( .A1(n10374), .A2(n10645), .ZN(n10376) );
  AND4_X1 U8026 ( .A1(n8527), .A2(n8526), .A3(n8525), .A4(n8524), .ZN(n12819)
         );
  AND2_X1 U8027 ( .A1(n7300), .A2(n7302), .ZN(n11775) );
  AND2_X1 U8028 ( .A1(n8759), .A2(n8758), .ZN(n12691) );
  NAND2_X1 U8029 ( .A1(n8727), .A2(n8726), .ZN(n12714) );
  INV_X1 U8030 ( .A(n12742), .ZN(n12713) );
  INV_X1 U8031 ( .A(n12819), .ZN(n12440) );
  NAND2_X1 U8032 ( .A1(n11148), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8507) );
  INV_X1 U8033 ( .A(n11040), .ZN(n12444) );
  INV_X1 U8034 ( .A(n15045), .ZN(n12448) );
  XNOR2_X1 U8035 ( .A(n7271), .B(n14900), .ZN(n14892) );
  AND2_X1 U8036 ( .A1(n8535), .A2(n8534), .ZN(n15009) );
  OAI211_X1 U8037 ( .C1(n7270), .C2(n6997), .A(n6995), .B(n6993), .ZN(n12452)
         );
  INV_X1 U8038 ( .A(n6998), .ZN(n6997) );
  AND2_X1 U8039 ( .A1(n6996), .A2(n6999), .ZN(n6995) );
  XNOR2_X1 U8040 ( .A(n12520), .B(n12525), .ZN(n12502) );
  OR2_X1 U8041 ( .A1(n14458), .A2(n14459), .ZN(n6992) );
  INV_X1 U8042 ( .A(n6595), .ZN(n6594) );
  OAI21_X1 U8043 ( .B1(n6429), .B2(n6596), .A(n12575), .ZN(n6595) );
  INV_X1 U8044 ( .A(n12555), .ZN(n6596) );
  NAND2_X1 U8045 ( .A1(n8813), .A2(n8812), .ZN(n12634) );
  NAND2_X1 U8046 ( .A1(n8767), .A2(n8766), .ZN(n12667) );
  NAND2_X1 U8047 ( .A1(n8752), .A2(n8751), .ZN(n12684) );
  AND3_X1 U8048 ( .A1(n8521), .A2(n8520), .A3(n8519), .ZN(n12307) );
  NAND2_X1 U8049 ( .A1(n12205), .A2(n12204), .ZN(n12832) );
  NAND2_X1 U8050 ( .A1(n8940), .A2(n8939), .ZN(n7531) );
  AOI21_X1 U8051 ( .B1(n8939), .B2(n15072), .A(n15114), .ZN(n7530) );
  NOR2_X1 U8052 ( .A1(n15117), .A2(n8956), .ZN(n7536) );
  NAND2_X1 U8053 ( .A1(n6570), .A2(n8939), .ZN(n12613) );
  OR2_X1 U8054 ( .A1(n8940), .A2(n15072), .ZN(n6570) );
  AND2_X1 U8055 ( .A1(n12607), .A2(n14490), .ZN(n7534) );
  NAND2_X1 U8056 ( .A1(n11797), .A2(n7492), .ZN(n14508) );
  NOR2_X1 U8057 ( .A1(n14506), .A2(n7493), .ZN(n7492) );
  INV_X1 U8058 ( .A(n11796), .ZN(n7493) );
  NOR2_X1 U8059 ( .A1(n6413), .A2(n13073), .ZN(n7047) );
  INV_X1 U8060 ( .A(n7052), .ZN(n7049) );
  NAND2_X1 U8061 ( .A1(n7051), .A2(n7053), .ZN(n7050) );
  NAND2_X1 U8062 ( .A1(n7054), .A2(n12997), .ZN(n7053) );
  NAND2_X1 U8063 ( .A1(n13084), .A2(n6676), .ZN(n12052) );
  OR2_X1 U8064 ( .A1(n12046), .A2(n12047), .ZN(n6676) );
  NAND3_X2 U8065 ( .A1(n7687), .A2(n6951), .A3(n7688), .ZN(n9736) );
  INV_X1 U8066 ( .A(n7498), .ZN(n13015) );
  NAND2_X1 U8067 ( .A1(n11997), .A2(n11996), .ZN(n6672) );
  INV_X1 U8068 ( .A(n13585), .ZN(n13422) );
  AND2_X1 U8069 ( .A1(n9981), .A2(n9739), .ZN(n10037) );
  NAND2_X1 U8070 ( .A1(n8091), .A2(n8090), .ZN(n13370) );
  INV_X1 U8071 ( .A(n13348), .ZN(n13491) );
  NAND2_X1 U8072 ( .A1(n7554), .A2(n7556), .ZN(n8309) );
  NOR2_X1 U8073 ( .A1(n7557), .A2(n9863), .ZN(n7553) );
  INV_X1 U8074 ( .A(n8340), .ZN(n6920) );
  NAND2_X1 U8075 ( .A1(n8262), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8165) );
  NAND2_X1 U8076 ( .A1(n8262), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8019) );
  NAND2_X1 U8077 ( .A1(n8262), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n7917) );
  NAND2_X1 U8078 ( .A1(n8262), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7897) );
  NAND2_X1 U8079 ( .A1(n8262), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7881) );
  NAND2_X1 U8080 ( .A1(n8262), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n7854) );
  NAND2_X1 U8081 ( .A1(n8262), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n7833) );
  AND2_X1 U8082 ( .A1(n6614), .A2(n6613), .ZN(n9898) );
  NAND2_X1 U8083 ( .A1(n9661), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6613) );
  NOR2_X1 U8084 ( .A1(n9907), .A2(n9906), .ZN(n9905) );
  NOR2_X1 U8085 ( .A1(n13167), .A2(n6635), .ZN(n13169) );
  INV_X1 U8086 ( .A(n6634), .ZN(n6635) );
  AND2_X1 U8087 ( .A1(n9668), .A2(n9644), .ZN(n14770) );
  AOI21_X1 U8088 ( .B1(n13445), .B2(n14806), .A(n13259), .ZN(n7294) );
  NAND2_X1 U8089 ( .A1(n7101), .A2(n6471), .ZN(n7100) );
  OAI21_X1 U8090 ( .B1(n8053), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7668) );
  AOI22_X1 U8091 ( .A1(n13260), .A2(n7017), .B1(n7015), .B2(n7014), .ZN(n7013)
         );
  NAND2_X1 U8092 ( .A1(n13258), .A2(n7016), .ZN(n7015) );
  NAND2_X1 U8093 ( .A1(n7295), .A2(n7018), .ZN(n7014) );
  NOR2_X1 U8094 ( .A1(n7295), .A2(n7019), .ZN(n7017) );
  NAND2_X1 U8095 ( .A1(n7830), .A2(n7829), .ZN(n10785) );
  AND2_X1 U8096 ( .A1(n7436), .A2(n6563), .ZN(n11868) );
  NAND2_X1 U8097 ( .A1(n13586), .A2(n7910), .ZN(n7436) );
  AOI21_X1 U8098 ( .B1(n11864), .B2(n13390), .A(n11865), .ZN(n11860) );
  AND2_X1 U8099 ( .A1(n8279), .A2(n8278), .ZN(n13545) );
  OR2_X1 U8100 ( .A1(n14283), .A2(n8277), .ZN(n8279) );
  AND2_X1 U8101 ( .A1(n7013), .A2(n7012), .ZN(n7011) );
  NOR2_X1 U8102 ( .A1(n14846), .A2(n13531), .ZN(n7012) );
  NAND2_X1 U8103 ( .A1(n7877), .A2(n7876), .ZN(n11053) );
  NAND2_X1 U8104 ( .A1(n14848), .A2(n14830), .ZN(n13584) );
  MUX2_X1 U8105 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7658), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n7660) );
  NAND2_X1 U8106 ( .A1(n9163), .A2(n9162), .ZN(n14623) );
  NAND2_X1 U8107 ( .A1(n9084), .A2(n9083), .ZN(n11004) );
  OR2_X1 U8108 ( .A1(n9604), .A2(n9440), .ZN(n9149) );
  NAND2_X1 U8109 ( .A1(n10059), .A2(n9454), .ZN(n6830) );
  INV_X1 U8110 ( .A(n13771), .ZN(n13757) );
  OR2_X1 U8111 ( .A1(n9036), .A2(n6898), .ZN(n9066) );
  INV_X1 U8112 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7648) );
  AOI21_X1 U8113 ( .B1(n13946), .B2(n14245), .A(n13945), .ZN(n14170) );
  NAND2_X1 U8114 ( .A1(n13944), .A2(n13943), .ZN(n13945) );
  NOR2_X1 U8115 ( .A1(n7394), .A2(n13905), .ZN(n7393) );
  INV_X1 U8116 ( .A(n7398), .ZN(n7394) );
  INV_X1 U8117 ( .A(n13947), .ZN(n13948) );
  INV_X1 U8118 ( .A(n14171), .ZN(n13968) );
  AOI21_X1 U8119 ( .B1(n6649), .B2(n14245), .A(n6988), .ZN(n6987) );
  INV_X1 U8120 ( .A(n13963), .ZN(n6988) );
  XNOR2_X1 U8121 ( .A(n6650), .B(n13958), .ZN(n6649) );
  NAND2_X1 U8122 ( .A1(n6979), .A2(n14421), .ZN(n14426) );
  OAI21_X1 U8123 ( .B1(n14423), .B2(n14422), .A(n6980), .ZN(n6979) );
  INV_X1 U8124 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n6980) );
  XNOR2_X1 U8125 ( .A(n14396), .B(n7159), .ZN(n14581) );
  INV_X1 U8126 ( .A(n14397), .ZN(n7159) );
  NAND2_X1 U8127 ( .A1(n14581), .A2(n14778), .ZN(n14580) );
  NAND2_X1 U8128 ( .A1(n14436), .A2(n14438), .ZN(n14441) );
  NAND2_X1 U8129 ( .A1(n14441), .A2(n14442), .ZN(n14443) );
  OAI21_X1 U8130 ( .B1(n14441), .B2(n14442), .A(n15186), .ZN(n7164) );
  NAND2_X1 U8131 ( .A1(n7768), .A2(n9736), .ZN(n7689) );
  AOI21_X1 U8132 ( .B1(n6407), .B2(n7463), .A(n7462), .ZN(n7461) );
  OAI21_X1 U8133 ( .B1(n9092), .B2(n6407), .A(n6959), .ZN(n9109) );
  NOR2_X1 U8134 ( .A1(n6960), .A2(n9108), .ZN(n6959) );
  INV_X1 U8135 ( .A(n7463), .ZN(n6960) );
  NAND2_X1 U8136 ( .A1(n9122), .A2(n7447), .ZN(n7446) );
  INV_X1 U8137 ( .A(n9121), .ZN(n7447) );
  NAND2_X1 U8138 ( .A1(n6507), .A2(n6974), .ZN(n6741) );
  NAND2_X1 U8139 ( .A1(n6856), .A2(n7470), .ZN(n9166) );
  NAND2_X1 U8140 ( .A1(n7471), .A2(n9150), .ZN(n7470) );
  NAND2_X1 U8141 ( .A1(n9131), .A2(n6854), .ZN(n6853) );
  INV_X1 U8142 ( .A(n9183), .ZN(n7455) );
  NAND2_X1 U8143 ( .A1(n6739), .A2(n6738), .ZN(n6737) );
  INV_X1 U8144 ( .A(n7888), .ZN(n6739) );
  INV_X1 U8145 ( .A(n7887), .ZN(n6738) );
  NAND2_X1 U8146 ( .A1(n7887), .A2(n7888), .ZN(n6740) );
  NAND2_X1 U8147 ( .A1(n6864), .A2(n6863), .ZN(n9242) );
  NAND2_X1 U8148 ( .A1(n6865), .A2(n9198), .ZN(n6863) );
  NAND2_X1 U8149 ( .A1(n6749), .A2(n6753), .ZN(n7950) );
  OR2_X1 U8150 ( .A1(n7925), .A2(n6754), .ZN(n6749) );
  NAND2_X1 U8151 ( .A1(n6752), .A2(n6750), .ZN(n7952) );
  AOI21_X1 U8152 ( .B1(n6754), .B2(n6753), .A(n6751), .ZN(n6750) );
  INV_X1 U8153 ( .A(n7949), .ZN(n6751) );
  AND2_X1 U8154 ( .A1(n9245), .A2(n9246), .ZN(n6906) );
  NAND2_X1 U8155 ( .A1(n9242), .A2(n9243), .ZN(n9249) );
  NAND2_X1 U8156 ( .A1(n7591), .A2(n6409), .ZN(n7590) );
  AND2_X1 U8157 ( .A1(n6947), .A2(n6869), .ZN(n6868) );
  NOR2_X1 U8158 ( .A1(n6949), .A2(n6948), .ZN(n6947) );
  NAND2_X1 U8159 ( .A1(n6758), .A2(n6756), .ZN(n8048) );
  INV_X1 U8160 ( .A(n9339), .ZN(n7460) );
  INV_X1 U8161 ( .A(n9303), .ZN(n6894) );
  INV_X1 U8162 ( .A(n9326), .ZN(n6899) );
  NAND2_X1 U8163 ( .A1(n7565), .A2(n8138), .ZN(n7564) );
  INV_X1 U8164 ( .A(n8141), .ZN(n7565) );
  AND2_X1 U8165 ( .A1(n9354), .A2(n6852), .ZN(n6851) );
  NAND2_X1 U8166 ( .A1(n6851), .A2(n6850), .ZN(n6849) );
  NOR2_X1 U8167 ( .A1(n8153), .A2(n7562), .ZN(n7561) );
  INV_X1 U8168 ( .A(n7564), .ZN(n7562) );
  INV_X1 U8169 ( .A(n8050), .ZN(n8051) );
  INV_X1 U8170 ( .A(n7953), .ZN(n7414) );
  INV_X1 U8171 ( .A(n7970), .ZN(n7417) );
  INV_X1 U8172 ( .A(n7956), .ZN(n7416) );
  INV_X1 U8173 ( .A(n8868), .ZN(n7184) );
  NAND2_X1 U8174 ( .A1(n12448), .A2(n10776), .ZN(n12272) );
  INV_X1 U8175 ( .A(n9449), .ZN(n6879) );
  NAND2_X1 U8176 ( .A1(n7453), .A2(n9386), .ZN(n7452) );
  INV_X1 U8177 ( .A(n9387), .ZN(n7453) );
  NAND2_X1 U8178 ( .A1(n9445), .A2(n8999), .ZN(n7442) );
  NAND2_X1 U8179 ( .A1(n9478), .A2(n13914), .ZN(n6626) );
  INV_X1 U8180 ( .A(n6626), .ZN(n6624) );
  INV_X1 U8181 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n15169) );
  NOR2_X1 U8182 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n8965) );
  NOR2_X1 U8183 ( .A1(n8208), .A2(n11582), .ZN(n7426) );
  INV_X1 U8184 ( .A(n7426), .ZN(n7423) );
  AOI21_X1 U8185 ( .B1(n7427), .B2(n8208), .A(n7425), .ZN(n7424) );
  NOR2_X1 U8186 ( .A1(n8192), .A2(SI_26_), .ZN(n7425) );
  INV_X1 U8187 ( .A(n8142), .ZN(n7400) );
  NAND2_X1 U8188 ( .A1(n8143), .A2(SI_22_), .ZN(n8144) );
  AND2_X1 U8189 ( .A1(n8071), .A2(n7406), .ZN(n7401) );
  INV_X1 U8190 ( .A(n8088), .ZN(n7406) );
  AND2_X1 U8191 ( .A1(n7402), .A2(n6542), .ZN(n7006) );
  INV_X1 U8192 ( .A(n8001), .ZN(n8004) );
  AND2_X1 U8193 ( .A1(n7413), .A2(n7029), .ZN(n7028) );
  NAND2_X1 U8194 ( .A1(n7030), .A2(n7932), .ZN(n7029) );
  NOR2_X1 U8195 ( .A1(n7417), .A2(n7414), .ZN(n7413) );
  INV_X1 U8196 ( .A(n7928), .ZN(n7030) );
  INV_X1 U8197 ( .A(n7026), .ZN(n6574) );
  AOI21_X1 U8198 ( .B1(n7028), .B2(n7031), .A(n7027), .ZN(n7026) );
  INV_X1 U8199 ( .A(n7415), .ZN(n7027) );
  AOI21_X1 U8200 ( .B1(n7970), .B2(n7416), .A(n6496), .ZN(n7415) );
  NAND2_X1 U8201 ( .A1(n7649), .A2(n7648), .ZN(n7650) );
  NAND3_X1 U8202 ( .A1(n14444), .A2(n7647), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n7649) );
  INV_X1 U8203 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7647) );
  NAND2_X1 U8204 ( .A1(n6801), .A2(n14313), .ZN(n14315) );
  NAND2_X1 U8205 ( .A1(n14360), .A2(n14359), .ZN(n6801) );
  INV_X1 U8206 ( .A(n12244), .ZN(n6763) );
  XNOR2_X1 U8207 ( .A(n12859), .B(n10229), .ZN(n12078) );
  INV_X1 U8208 ( .A(n10916), .ZN(n7338) );
  NAND2_X1 U8209 ( .A1(n11148), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8931) );
  AND3_X1 U8210 ( .A1(n8389), .A2(n8388), .A3(n8387), .ZN(n8391) );
  NAND2_X1 U8211 ( .A1(n14884), .A2(n6954), .ZN(n11479) );
  OR2_X1 U8212 ( .A1(n11494), .A2(n15152), .ZN(n6954) );
  INV_X1 U8213 ( .A(n14872), .ZN(n6603) );
  NAND2_X1 U8214 ( .A1(n14923), .A2(n6910), .ZN(n11482) );
  NAND2_X1 U8215 ( .A1(n14919), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n6910) );
  NAND2_X1 U8216 ( .A1(n12504), .A2(n12506), .ZN(n12524) );
  OR2_X1 U8217 ( .A1(n8828), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8879) );
  NAND2_X1 U8218 ( .A1(n8814), .A2(n12093), .ZN(n8828) );
  INV_X1 U8219 ( .A(n8815), .ZN(n8814) );
  OAI22_X1 U8220 ( .A1(n12638), .A2(n12639), .B1(n12432), .B2(n12388), .ZN(
        n12627) );
  NOR2_X1 U8221 ( .A1(n7173), .A2(n8777), .ZN(n7540) );
  NAND2_X1 U8222 ( .A1(n8719), .A2(n8718), .ZN(n8738) );
  INV_X1 U8223 ( .A(n8720), .ZN(n8719) );
  NAND2_X1 U8224 ( .A1(n11148), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8708) );
  OR2_X1 U8225 ( .A1(n8644), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8657) );
  INV_X1 U8226 ( .A(n8864), .ZN(n6568) );
  NAND2_X1 U8227 ( .A1(n8586), .A2(n11590), .ZN(n8603) );
  INV_X1 U8228 ( .A(n8587), .ZN(n8586) );
  NAND2_X1 U8229 ( .A1(n11148), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8403) );
  NAND2_X1 U8230 ( .A1(n15050), .A2(n15049), .ZN(n7198) );
  NAND2_X1 U8231 ( .A1(n8850), .A2(n15055), .ZN(n12266) );
  NAND2_X1 U8232 ( .A1(n12275), .A2(n12272), .ZN(n8852) );
  NAND2_X1 U8233 ( .A1(n10248), .A2(n12449), .ZN(n12263) );
  NAND2_X1 U8234 ( .A1(n15041), .A2(n15040), .ZN(n15043) );
  INV_X1 U8235 ( .A(n8810), .ZN(n7152) );
  NOR2_X1 U8236 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_24__SCAN_IN), .ZN(
        n6775) );
  AND2_X1 U8237 ( .A1(n7121), .A2(n11352), .ZN(n7118) );
  INV_X1 U8238 ( .A(n7134), .ZN(n7133) );
  OAI21_X1 U8239 ( .B1(n8634), .B2(n7135), .A(n8664), .ZN(n7134) );
  INV_X1 U8240 ( .A(n8650), .ZN(n7135) );
  AOI21_X1 U8241 ( .B1(n8561), .B2(n7109), .A(n7108), .ZN(n7107) );
  INV_X1 U8242 ( .A(n8578), .ZN(n7108) );
  INV_X1 U8243 ( .A(n8558), .ZN(n7109) );
  NAND2_X1 U8244 ( .A1(n8550), .A2(n6654), .ZN(n6653) );
  NOR2_X1 U8245 ( .A1(n6655), .A2(n7110), .ZN(n6654) );
  INV_X1 U8246 ( .A(n8561), .ZN(n7110) );
  INV_X1 U8247 ( .A(n8549), .ZN(n6655) );
  INV_X1 U8248 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8479) );
  INV_X1 U8249 ( .A(n7140), .ZN(n7139) );
  OAI21_X1 U8250 ( .B1(n8511), .B2(n7141), .A(n8545), .ZN(n7140) );
  INV_X1 U8251 ( .A(n8528), .ZN(n7141) );
  INV_X1 U8252 ( .A(n8490), .ZN(n7143) );
  OR2_X1 U8253 ( .A1(n8496), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n8514) );
  INV_X1 U8254 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8343) );
  NAND2_X1 U8255 ( .A1(n7572), .A2(n7571), .ZN(n7570) );
  AOI21_X1 U8256 ( .B1(n7574), .B2(n7576), .A(n7569), .ZN(n7568) );
  INV_X1 U8257 ( .A(n7578), .ZN(n7576) );
  AND2_X1 U8258 ( .A1(n6747), .A2(n6514), .ZN(n6744) );
  AND2_X1 U8259 ( .A1(n8327), .A2(n7607), .ZN(n8271) );
  NOR2_X1 U8260 ( .A1(n6617), .A2(n6616), .ZN(n6615) );
  INV_X1 U8261 ( .A(n13197), .ZN(n6586) );
  INV_X1 U8262 ( .A(n6691), .ZN(n6690) );
  INV_X1 U8263 ( .A(n11823), .ZN(n7080) );
  INV_X1 U8264 ( .A(n7077), .ZN(n7075) );
  INV_X1 U8265 ( .A(n11209), .ZN(n6698) );
  AND2_X1 U8266 ( .A1(n11210), .A2(n11197), .ZN(n7077) );
  INV_X1 U8267 ( .A(n14831), .ZN(n7068) );
  AND2_X1 U8268 ( .A1(n7066), .A2(n6435), .ZN(n11058) );
  NAND2_X1 U8269 ( .A1(n7652), .A2(n6966), .ZN(n6972) );
  NOR2_X1 U8270 ( .A1(n6971), .A2(n6970), .ZN(n6969) );
  NOR2_X1 U8271 ( .A1(n7827), .A2(n6973), .ZN(n6966) );
  INV_X1 U8272 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n7617) );
  INV_X1 U8273 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n7621) );
  AND2_X1 U8274 ( .A1(n7665), .A2(n7628), .ZN(n7653) );
  NOR2_X1 U8275 ( .A1(n7911), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n7934) );
  NOR2_X1 U8276 ( .A1(n13647), .A2(n13648), .ZN(n7243) );
  INV_X1 U8277 ( .A(n9343), .ZN(n9344) );
  NAND2_X1 U8278 ( .A1(n9344), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n9357) );
  NOR2_X1 U8279 ( .A1(n11925), .A2(n11915), .ZN(n7242) );
  OAI22_X1 U8280 ( .A1(n9449), .A2(n9450), .B1(n9451), .B2(n9452), .ZN(n6875)
         );
  INV_X1 U8281 ( .A(n6877), .ZN(n6876) );
  OAI21_X1 U8282 ( .B1(n6879), .B2(n6878), .A(n7441), .ZN(n6877) );
  INV_X1 U8283 ( .A(n9450), .ZN(n6878) );
  NAND2_X1 U8284 ( .A1(n9413), .A2(n9411), .ZN(n7441) );
  AND2_X1 U8285 ( .A1(n6872), .A2(n7439), .ZN(n6871) );
  NAND2_X1 U8286 ( .A1(n9412), .A2(n7440), .ZN(n7439) );
  INV_X1 U8287 ( .A(n6875), .ZN(n6872) );
  INV_X1 U8288 ( .A(n9411), .ZN(n7440) );
  AOI21_X1 U8289 ( .B1(n7364), .B2(n7367), .A(n6482), .ZN(n7362) );
  INV_X1 U8290 ( .A(n7364), .ZN(n7363) );
  OR2_X1 U8291 ( .A1(n14033), .A2(n13775), .ZN(n13918) );
  OR2_X1 U8292 ( .A1(n14057), .A2(n14070), .ZN(n7374) );
  NAND2_X1 U8293 ( .A1(n6625), .A2(n6622), .ZN(n14057) );
  AOI21_X1 U8294 ( .B1(n6624), .B2(n14099), .A(n6623), .ZN(n6622) );
  OR2_X1 U8295 ( .A1(n14098), .A2(n6626), .ZN(n6625) );
  INV_X1 U8296 ( .A(n13915), .ZN(n6623) );
  INV_X1 U8297 ( .A(n7381), .ZN(n6829) );
  OAI21_X1 U8298 ( .B1(n11317), .B2(n7382), .A(n11550), .ZN(n7381) );
  INV_X1 U8299 ( .A(n11280), .ZN(n7382) );
  AND2_X1 U8300 ( .A1(n11279), .A2(n7344), .ZN(n7343) );
  NAND2_X1 U8301 ( .A1(n11274), .A2(n7345), .ZN(n7344) );
  INV_X1 U8302 ( .A(n11272), .ZN(n7345) );
  INV_X1 U8303 ( .A(n11274), .ZN(n7346) );
  INV_X1 U8304 ( .A(n10080), .ZN(n10086) );
  NOR2_X1 U8305 ( .A1(n9417), .A2(n10149), .ZN(n6942) );
  AND2_X1 U8306 ( .A1(n9433), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6943) );
  INV_X1 U8307 ( .A(n7353), .ZN(n7352) );
  AOI21_X1 U8308 ( .B1(n6403), .B2(n14143), .A(n6452), .ZN(n7353) );
  NOR2_X1 U8309 ( .A1(n14237), .A2(n9486), .ZN(n7213) );
  NOR2_X1 U8310 ( .A1(n14562), .A2(n6822), .ZN(n6820) );
  NAND2_X1 U8311 ( .A1(n14618), .A2(n14617), .ZN(n14620) );
  XNOR2_X1 U8312 ( .A(n13787), .B(n6936), .ZN(n10080) );
  NAND2_X1 U8313 ( .A1(n10081), .A2(n10080), .ZN(n10512) );
  INV_X1 U8314 ( .A(n10633), .ZN(n10624) );
  INV_X1 U8315 ( .A(n8247), .ZN(n7433) );
  INV_X1 U8316 ( .A(n8248), .ZN(n7434) );
  NOR2_X1 U8317 ( .A1(n9192), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n9208) );
  XNOR2_X1 U8318 ( .A(n7955), .B(SI_12_), .ZN(n7953) );
  NAND2_X1 U8319 ( .A1(n6832), .A2(n6831), .ZN(n7954) );
  AOI21_X1 U8320 ( .B1(n6833), .B2(n6580), .A(n7031), .ZN(n6831) );
  NAND2_X1 U8321 ( .A1(n7890), .A2(n6833), .ZN(n6832) );
  INV_X1 U8322 ( .A(n6834), .ZN(n6833) );
  OR2_X1 U8323 ( .A1(n9179), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n9192) );
  NOR2_X1 U8324 ( .A1(n7908), .A2(n6836), .ZN(n6835) );
  INV_X1 U8325 ( .A(n7889), .ZN(n6836) );
  INV_X1 U8326 ( .A(n7865), .ZN(n7409) );
  INV_X1 U8327 ( .A(n7411), .ZN(n7410) );
  INV_X1 U8328 ( .A(n7820), .ZN(n6841) );
  NOR2_X1 U8329 ( .A1(n9142), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n9145) );
  OR2_X1 U8330 ( .A1(n9127), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9142) );
  NAND2_X1 U8331 ( .A1(n6499), .A2(n7820), .ZN(n6840) );
  INV_X1 U8332 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9101) );
  INV_X1 U8333 ( .A(n7034), .ZN(n7733) );
  XNOR2_X1 U8334 ( .A(n14315), .B(n14314), .ZN(n14357) );
  INV_X1 U8335 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n14314) );
  NOR2_X1 U8336 ( .A1(n14327), .A2(n14326), .ZN(n14328) );
  NOR2_X1 U8337 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n14386), .ZN(n14326) );
  INV_X1 U8338 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n6798) );
  OAI21_X1 U8339 ( .B1(n15013), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n14332), .ZN(
        n14391) );
  OR2_X1 U8340 ( .A1(n14355), .A2(n14354), .ZN(n14332) );
  NAND2_X1 U8341 ( .A1(n8691), .A2(n8690), .ZN(n8705) );
  INV_X1 U8342 ( .A(n8692), .ZN(n8691) );
  AOI21_X1 U8343 ( .B1(n12092), .B2(n12091), .A(n12110), .ZN(n7311) );
  INV_X1 U8344 ( .A(n7311), .ZN(n7309) );
  INV_X1 U8345 ( .A(n15074), .ZN(n10248) );
  NAND2_X1 U8346 ( .A1(n11148), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8801) );
  AND2_X1 U8347 ( .A1(n12088), .A2(n12087), .ZN(n12131) );
  XNOR2_X1 U8348 ( .A(n10229), .B(n10756), .ZN(n10368) );
  AND2_X1 U8349 ( .A1(n11454), .A2(n11587), .ZN(n7301) );
  NAND2_X1 U8350 ( .A1(n12129), .A2(n12088), .ZN(n12190) );
  OR2_X1 U8351 ( .A1(n8798), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8815) );
  NAND2_X1 U8352 ( .A1(n8782), .A2(n15121), .ZN(n8798) );
  INV_X1 U8353 ( .A(n8783), .ZN(n8782) );
  NAND2_X1 U8354 ( .A1(n7332), .A2(n7331), .ZN(n11814) );
  OR2_X1 U8355 ( .A1(n8603), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8625) );
  NAND2_X1 U8356 ( .A1(n8624), .A2(n15243), .ZN(n8644) );
  INV_X1 U8357 ( .A(n8625), .ZN(n8624) );
  NAND2_X1 U8358 ( .A1(n7130), .A2(n7128), .ZN(n7127) );
  AOI21_X1 U8359 ( .B1(n7129), .B2(n6455), .A(n12418), .ZN(n7128) );
  NAND2_X1 U8360 ( .A1(n12416), .A2(n12415), .ZN(n7130) );
  NAND2_X1 U8361 ( .A1(n11148), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8786) );
  OR2_X1 U8362 ( .A1(n6913), .A2(n10841), .ZN(n7260) );
  INV_X1 U8363 ( .A(n7001), .ZN(n11464) );
  INV_X1 U8364 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n10882) );
  XNOR2_X1 U8365 ( .A(n11482), .B(n11509), .ZN(n14944) );
  OR2_X1 U8366 ( .A1(n14930), .A2(n11469), .ZN(n7266) );
  OR2_X1 U8367 ( .A1(n11469), .A2(n6528), .ZN(n7000) );
  XNOR2_X1 U8368 ( .A(n11484), .B(n11520), .ZN(n14984) );
  NAND2_X1 U8369 ( .A1(n14961), .A2(n6912), .ZN(n11484) );
  OR2_X1 U8370 ( .A1(n11514), .A2(n11575), .ZN(n6912) );
  NAND2_X1 U8371 ( .A1(n6598), .A2(n6551), .ZN(n11472) );
  NAND2_X1 U8372 ( .A1(n14989), .A2(n6911), .ZN(n11701) );
  OR2_X1 U8373 ( .A1(n15009), .A2(n15115), .ZN(n6911) );
  NOR2_X1 U8374 ( .A1(n12483), .A2(n11698), .ZN(n6994) );
  NAND2_X1 U8375 ( .A1(n6998), .A2(n11698), .ZN(n6996) );
  OR2_X1 U8376 ( .A1(n12483), .A2(n7267), .ZN(n6999) );
  AND2_X1 U8377 ( .A1(n12483), .A2(n7267), .ZN(n6998) );
  XNOR2_X1 U8378 ( .A(n12524), .B(n12532), .ZN(n12505) );
  AND2_X1 U8379 ( .A1(n8845), .A2(n12586), .ZN(n10706) );
  NAND2_X1 U8380 ( .A1(n12546), .A2(n6560), .ZN(n12548) );
  XNOR2_X1 U8381 ( .A(n12548), .B(n12563), .ZN(n14451) );
  AOI21_X1 U8382 ( .B1(n7507), .B2(n7509), .A(n12394), .ZN(n6660) );
  NAND2_X1 U8383 ( .A1(n12637), .A2(n7507), .ZN(n6659) );
  INV_X1 U8384 ( .A(n7510), .ZN(n7509) );
  INV_X1 U8385 ( .A(n12391), .ZN(n6881) );
  AND2_X1 U8386 ( .A1(n7511), .A2(n12396), .ZN(n7510) );
  AND2_X1 U8387 ( .A1(n8876), .A2(n12395), .ZN(n12639) );
  AOI21_X1 U8388 ( .B1(n12700), .B2(n7168), .A(n7166), .ZN(n7165) );
  INV_X1 U8389 ( .A(n7172), .ZN(n7168) );
  OAI21_X1 U8390 ( .B1(n7172), .B2(n7167), .A(n7170), .ZN(n7166) );
  AND2_X1 U8391 ( .A1(n7169), .A2(n6445), .ZN(n12674) );
  OR2_X1 U8392 ( .A1(n7177), .A2(n7174), .ZN(n7169) );
  NOR2_X1 U8393 ( .A1(n12720), .A2(n7547), .ZN(n7546) );
  INV_X1 U8394 ( .A(n12363), .ZN(n7547) );
  AOI21_X1 U8395 ( .B1(n7527), .B2(n7525), .A(n7524), .ZN(n7523) );
  INV_X1 U8396 ( .A(n7527), .ZN(n7526) );
  INV_X1 U8397 ( .A(n12342), .ZN(n7524) );
  NAND2_X1 U8398 ( .A1(n7529), .A2(n12793), .ZN(n12792) );
  NAND2_X1 U8399 ( .A1(n8570), .A2(n8569), .ZN(n8587) );
  INV_X1 U8400 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n8569) );
  INV_X1 U8401 ( .A(n8571), .ZN(n8570) );
  AOI21_X1 U8402 ( .B1(n7517), .B2(n7518), .A(n6473), .ZN(n7515) );
  NAND2_X1 U8403 ( .A1(n8501), .A2(n10917), .ZN(n8522) );
  NAND2_X1 U8404 ( .A1(n8465), .A2(n10882), .ZN(n8484) );
  INV_X1 U8405 ( .A(n8466), .ZN(n8465) );
  NAND2_X1 U8406 ( .A1(n8431), .A2(n10650), .ZN(n8451) );
  NAND2_X1 U8407 ( .A1(n7198), .A2(n8851), .ZN(n10391) );
  INV_X1 U8408 ( .A(n15040), .ZN(n15049) );
  NAND2_X1 U8409 ( .A1(n12215), .A2(n12214), .ZN(n12600) );
  NAND2_X1 U8410 ( .A1(n8781), .A2(n8780), .ZN(n12247) );
  AND3_X1 U8411 ( .A1(n8450), .A2(n8449), .A3(n8448), .ZN(n10644) );
  NAND2_X1 U8412 ( .A1(n8891), .A2(n8890), .ZN(n6938) );
  OAI21_X1 U8413 ( .B1(n8765), .B2(n7155), .A(n7154), .ZN(n8793) );
  NAND2_X1 U8414 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n7156), .ZN(n7154) );
  AND2_X1 U8415 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n13613), .ZN(n7155) );
  NOR2_X1 U8416 ( .A1(n6775), .A2(P3_IR_REG_23__SCAN_IN), .ZN(n6771) );
  INV_X1 U8417 ( .A(n6775), .ZN(n6770) );
  OAI21_X1 U8418 ( .B1(n8748), .B2(n8747), .A(n8750), .ZN(n8761) );
  XNOR2_X1 U8419 ( .A(n8912), .B(n8911), .ZN(n10694) );
  XNOR2_X1 U8420 ( .A(n8835), .B(P3_IR_REG_21__SCAN_IN), .ZN(n12253) );
  XNOR2_X1 U8421 ( .A(n8837), .B(P3_IR_REG_20__SCAN_IN), .ZN(n8877) );
  NAND2_X1 U8422 ( .A1(n7122), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7121) );
  INV_X1 U8423 ( .A(n8701), .ZN(n7122) );
  NAND2_X1 U8424 ( .A1(n8702), .A2(n6548), .ZN(n7117) );
  AND2_X1 U8425 ( .A1(n8701), .A2(n8682), .ZN(n8699) );
  INV_X1 U8426 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8348) );
  INV_X1 U8427 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8347) );
  OR2_X1 U8428 ( .A1(n8684), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n8615) );
  AND2_X1 U8429 ( .A1(n8566), .A2(n8684), .ZN(n12454) );
  INV_X1 U8430 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8516) );
  OAI21_X1 U8431 ( .B1(n8473), .B2(n7145), .A(n7142), .ZN(n8494) );
  AOI21_X1 U8432 ( .B1(n7146), .B2(n7144), .A(n7143), .ZN(n7142) );
  INV_X1 U8433 ( .A(n7146), .ZN(n7145) );
  INV_X1 U8434 ( .A(n8472), .ZN(n7144) );
  NAND2_X1 U8435 ( .A1(n8441), .A2(n8440), .ZN(n8459) );
  AND2_X1 U8436 ( .A1(n8460), .A2(n8442), .ZN(n8458) );
  AND2_X1 U8437 ( .A1(n8426), .A2(n8411), .ZN(n8424) );
  AND2_X1 U8438 ( .A1(n8409), .A2(n8397), .ZN(n8407) );
  NAND2_X1 U8439 ( .A1(n8370), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8392) );
  NOR2_X1 U8440 ( .A1(n11138), .A2(n7059), .ZN(n7058) );
  INV_X1 U8441 ( .A(n11130), .ZN(n7059) );
  NOR2_X1 U8442 ( .A1(n12997), .A2(n12993), .ZN(n7052) );
  OR2_X1 U8443 ( .A1(n7831), .A2(n10427), .ZN(n7849) );
  XNOR2_X1 U8444 ( .A(n14831), .B(n12048), .ZN(n10950) );
  NOR2_X1 U8445 ( .A1(n10745), .A2(n7482), .ZN(n7481) );
  INV_X1 U8446 ( .A(n10742), .ZN(n7482) );
  INV_X1 U8447 ( .A(n7995), .ZN(n7779) );
  INV_X1 U8448 ( .A(n13049), .ZN(n7041) );
  NOR2_X1 U8449 ( .A1(n7939), .A2(n7938), .ZN(n7962) );
  NAND2_X1 U8450 ( .A1(n12040), .A2(n7502), .ZN(n7501) );
  INV_X1 U8451 ( .A(n12041), .ZN(n7502) );
  AND2_X1 U8452 ( .A1(n8028), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8030) );
  OR2_X1 U8453 ( .A1(n12976), .A2(n12978), .ZN(n7036) );
  NAND2_X1 U8454 ( .A1(n12039), .A2(n12038), .ZN(n7038) );
  INV_X1 U8455 ( .A(n7036), .ZN(n12977) );
  NOR2_X1 U8456 ( .A1(n7879), .A2(n7878), .ZN(n7895) );
  OR2_X1 U8457 ( .A1(n7849), .A2(n7848), .ZN(n7879) );
  NAND2_X1 U8458 ( .A1(n8092), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8111) );
  NOR2_X1 U8459 ( .A1(n8079), .A2(n8078), .ZN(n8092) );
  NAND2_X1 U8460 ( .A1(n6440), .A2(n7043), .ZN(n7042) );
  NAND2_X1 U8461 ( .A1(n7484), .A2(n12024), .ZN(n7483) );
  NOR2_X1 U8462 ( .A1(n7494), .A2(n7044), .ZN(n7043) );
  NAND2_X1 U8463 ( .A1(n6440), .A2(n12013), .ZN(n7045) );
  NOR2_X1 U8464 ( .A1(n8111), .A2(n13008), .ZN(n8133) );
  OR2_X1 U8465 ( .A1(n7915), .A2(n11261), .ZN(n7939) );
  NOR2_X1 U8466 ( .A1(n7784), .A2(n7783), .ZN(n7803) );
  OR2_X1 U8467 ( .A1(n7980), .A2(n7979), .ZN(n7997) );
  NOR2_X1 U8468 ( .A1(n7997), .A2(n11805), .ZN(n8028) );
  AND2_X1 U8469 ( .A1(n13321), .A2(n6956), .ZN(n6955) );
  AND2_X1 U8470 ( .A1(n8327), .A2(n8325), .ZN(n6958) );
  AND2_X1 U8471 ( .A1(n13174), .A2(n7505), .ZN(n8337) );
  NAND2_X1 U8472 ( .A1(n7725), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8281) );
  AND4_X1 U8473 ( .A1(n8241), .A2(n8240), .A3(n8239), .A4(n8238), .ZN(n13257)
         );
  AND4_X1 U8474 ( .A1(n8220), .A2(n8219), .A3(n8218), .A4(n8217), .ZN(n13000)
         );
  AND2_X1 U8475 ( .A1(n8064), .A2(n8063), .ZN(n13231) );
  NAND2_X1 U8476 ( .A1(n14752), .A2(n14751), .ZN(n6612) );
  INV_X1 U8477 ( .A(n6615), .ZN(n6611) );
  OAI21_X1 U8478 ( .B1(n14752), .B2(n6615), .A(n6609), .ZN(n6614) );
  AOI21_X1 U8479 ( .B1(n6610), .B2(n6611), .A(n9884), .ZN(n6609) );
  INV_X1 U8480 ( .A(n14751), .ZN(n6610) );
  NOR2_X1 U8481 ( .A1(n9905), .A2(n6631), .ZN(n9667) );
  NOR2_X1 U8482 ( .A1(n6633), .A2(n6632), .ZN(n6631) );
  NAND2_X1 U8483 ( .A1(n9667), .A2(n9666), .ZN(n10007) );
  NAND2_X1 U8484 ( .A1(n10300), .A2(n10299), .ZN(n11181) );
  NOR2_X1 U8485 ( .A1(n10287), .A2(n6647), .ZN(n10290) );
  AND2_X1 U8486 ( .A1(n10296), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6647) );
  NAND2_X1 U8487 ( .A1(n10290), .A2(n10289), .ZN(n11185) );
  NAND2_X1 U8488 ( .A1(n11181), .A2(n6950), .ZN(n14767) );
  OR2_X1 U8489 ( .A1(n11186), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6950) );
  NAND2_X1 U8490 ( .A1(n11185), .A2(n6646), .ZN(n14762) );
  OR2_X1 U8491 ( .A1(n11186), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6646) );
  NOR2_X1 U8492 ( .A1(n14762), .A2(n14763), .ZN(n14761) );
  OR2_X1 U8493 ( .A1(n11191), .A2(n11190), .ZN(n6640) );
  XNOR2_X1 U8494 ( .A(n13136), .B(n14779), .ZN(n14782) );
  AND2_X1 U8495 ( .A1(n6640), .A2(n6639), .ZN(n13136) );
  NAND2_X1 U8496 ( .A1(n13135), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6639) );
  NOR2_X1 U8497 ( .A1(n14782), .A2(n14781), .ZN(n14780) );
  OR2_X1 U8498 ( .A1(n14792), .A2(n6638), .ZN(n6637) );
  AND2_X1 U8499 ( .A1(n14801), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6638) );
  NAND2_X1 U8500 ( .A1(n6437), .A2(n6634), .ZN(n13154) );
  AOI21_X1 U8501 ( .B1(n13148), .B2(P2_REG2_REG_17__SCAN_IN), .A(n13146), .ZN(
        n13163) );
  NOR2_X1 U8502 ( .A1(n13154), .A2(n13155), .ZN(n13167) );
  NOR3_X1 U8503 ( .A1(n13305), .A2(n13446), .A3(n13292), .ZN(n7060) );
  NAND2_X1 U8504 ( .A1(n13460), .A2(n13550), .ZN(n7061) );
  AND2_X1 U8505 ( .A1(n7101), .A2(n7104), .ZN(n7099) );
  AOI21_X1 U8506 ( .B1(n7103), .B2(n13274), .A(n7102), .ZN(n7101) );
  OAI21_X1 U8507 ( .B1(n13261), .B2(n13262), .A(n14520), .ZN(n7102) );
  NAND2_X1 U8508 ( .A1(n7070), .A2(n7069), .ZN(n13334) );
  NOR2_X1 U8509 ( .A1(n8147), .A2(n12980), .ZN(n8164) );
  INV_X1 U8510 ( .A(n7070), .ZN(n13344) );
  NAND2_X1 U8511 ( .A1(n13185), .A2(n13184), .ZN(n13188) );
  NAND2_X1 U8512 ( .A1(n7071), .A2(n14546), .ZN(n11644) );
  NAND2_X1 U8513 ( .A1(n14517), .A2(n11360), .ZN(n14519) );
  OAI21_X1 U8514 ( .B1(n11207), .B2(n6696), .A(n6695), .ZN(n14533) );
  INV_X1 U8515 ( .A(n6697), .ZN(n6696) );
  AOI21_X1 U8516 ( .B1(n11055), .B2(n6697), .A(n6483), .ZN(n6695) );
  NOR2_X1 U8517 ( .A1(n11355), .A2(n6698), .ZN(n6697) );
  NAND2_X1 U8518 ( .A1(n11361), .A2(n8316), .ZN(n14532) );
  NAND2_X1 U8519 ( .A1(n11198), .A2(n7077), .ZN(n14517) );
  AOI21_X1 U8520 ( .B1(n10792), .B2(n7092), .A(n6486), .ZN(n7091) );
  NAND2_X1 U8521 ( .A1(n10972), .A2(n10783), .ZN(n11049) );
  NAND2_X1 U8522 ( .A1(n6435), .A2(n10541), .ZN(n10983) );
  NAND2_X1 U8523 ( .A1(n10541), .A2(n14813), .ZN(n10982) );
  NAND2_X1 U8524 ( .A1(n10193), .A2(n10192), .ZN(n10354) );
  NOR2_X1 U8525 ( .A1(n10000), .A2(n10107), .ZN(n10046) );
  NAND2_X1 U8526 ( .A1(n10046), .A2(n11008), .ZN(n10187) );
  NAND2_X1 U8527 ( .A1(n9996), .A2(n9997), .ZN(n9999) );
  NAND2_X1 U8528 ( .A1(n9995), .A2(n9736), .ZN(n9993) );
  NAND2_X1 U8529 ( .A1(n9979), .A2(n9980), .ZN(n9997) );
  NAND2_X1 U8530 ( .A1(n13261), .A2(n7018), .ZN(n7016) );
  NAND2_X1 U8531 ( .A1(n6583), .A2(n13213), .ZN(n13214) );
  NAND2_X1 U8532 ( .A1(n13276), .A2(n7103), .ZN(n6583) );
  AND2_X1 U8533 ( .A1(n9768), .A2(n9642), .ZN(n14522) );
  AND2_X1 U8534 ( .A1(n13329), .A2(n13328), .ZN(n13486) );
  OR2_X1 U8535 ( .A1(n13327), .A2(n13538), .ZN(n13329) );
  AND2_X1 U8536 ( .A1(n8056), .A2(n8055), .ZN(n13520) );
  NAND2_X1 U8537 ( .A1(n6693), .A2(n6691), .ZN(n13433) );
  NAND2_X1 U8538 ( .A1(n6693), .A2(n11827), .ZN(n13431) );
  INV_X1 U8539 ( .A(n14841), .ZN(n14830) );
  MUX2_X1 U8540 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7656), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n7657) );
  INV_X1 U8541 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n7503) );
  OR2_X1 U8542 ( .A1(n7974), .A2(n7827), .ZN(n7959) );
  OR2_X1 U8543 ( .A1(n7872), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n7874) );
  OR2_X1 U8544 ( .A1(n7874), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n7911) );
  NOR2_X1 U8545 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n7706) );
  INV_X2 U8546 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7708) );
  INV_X1 U8547 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8370) );
  INV_X1 U8548 ( .A(n9330), .ZN(n9331) );
  NAND2_X1 U8549 ( .A1(n9331), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n9343) );
  NAND2_X1 U8550 ( .A1(n7243), .A2(n7237), .ZN(n7236) );
  INV_X1 U8551 ( .A(n7238), .ZN(n7237) );
  NAND2_X1 U8552 ( .A1(n11938), .A2(n11937), .ZN(n7234) );
  NAND2_X1 U8553 ( .A1(n7233), .A2(n7232), .ZN(n7231) );
  INV_X1 U8554 ( .A(n13714), .ZN(n7233) );
  AND2_X1 U8555 ( .A1(n13663), .A2(n11877), .ZN(n7247) );
  INV_X1 U8556 ( .A(n13779), .ZN(n13667) );
  NOR2_X1 U8557 ( .A1(n11343), .A2(n7252), .ZN(n7251) );
  INV_X1 U8558 ( .A(n11293), .ZN(n7252) );
  NAND2_X1 U8559 ( .A1(n11289), .A2(n11288), .ZN(n7253) );
  INV_X1 U8560 ( .A(n9847), .ZN(n9848) );
  OR2_X1 U8561 ( .A1(n9185), .A2(n10281), .ZN(n9200) );
  NOR2_X1 U8562 ( .A1(n9200), .A2(n9199), .ZN(n9220) );
  AOI21_X1 U8563 ( .B1(n7227), .B2(n7228), .A(n7226), .ZN(n7225) );
  INV_X1 U8564 ( .A(n7227), .ZN(n6722) );
  INV_X1 U8565 ( .A(n13732), .ZN(n7226) );
  NOR2_X1 U8566 ( .A1(n13742), .A2(n7239), .ZN(n7238) );
  INV_X1 U8567 ( .A(n7241), .ZN(n7239) );
  NAND2_X1 U8568 ( .A1(n11924), .A2(n13692), .ZN(n7241) );
  NAND2_X1 U8569 ( .A1(n13694), .A2(n7242), .ZN(n7240) );
  NAND2_X1 U8570 ( .A1(n10855), .A2(n10854), .ZN(n10860) );
  NAND2_X1 U8571 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n9358), .ZN(n9377) );
  NAND2_X1 U8572 ( .A1(n13625), .A2(n11904), .ZN(n7222) );
  AND4_X1 U8573 ( .A1(n9239), .A2(n9238), .A3(n9237), .A4(n9236), .ZN(n13686)
         );
  AOI21_X1 U8574 ( .B1(n9709), .B2(P1_REG1_REG_7__SCAN_IN), .A(n9947), .ZN(
        n9712) );
  AOI21_X1 U8575 ( .B1(n10063), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10062), .ZN(
        n10066) );
  AOI21_X1 U8576 ( .B1(n11760), .B2(P1_REG1_REG_16__SCAN_IN), .A(n11759), .ZN(
        n11762) );
  AOI21_X1 U8577 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n13846), .A(n13845), .ZN(
        n13859) );
  OR2_X1 U8578 ( .A1(n6826), .A2(n14167), .ZN(n13947) );
  OAI21_X1 U8579 ( .B1(n7363), .B2(n13988), .A(n7362), .ZN(n6650) );
  NAND2_X1 U8580 ( .A1(n7210), .A2(n14012), .ZN(n14006) );
  NAND2_X1 U8581 ( .A1(n9338), .A2(n9337), .ZN(n14017) );
  NAND2_X1 U8582 ( .A1(n14034), .A2(n13918), .ZN(n14016) );
  NAND2_X1 U8583 ( .A1(n14035), .A2(n14036), .ZN(n14034) );
  NAND2_X1 U8584 ( .A1(n6815), .A2(n6816), .ZN(n14028) );
  INV_X1 U8585 ( .A(n13917), .ZN(n14036) );
  NAND2_X1 U8586 ( .A1(n14046), .A2(n7383), .ZN(n14027) );
  AND2_X1 U8587 ( .A1(n13899), .A2(n13916), .ZN(n7384) );
  NOR2_X1 U8588 ( .A1(n6462), .A2(n14047), .ZN(n7372) );
  NAND2_X1 U8589 ( .A1(n14057), .A2(n6427), .ZN(n7368) );
  INV_X1 U8590 ( .A(n13900), .ZN(n14047) );
  AND2_X1 U8591 ( .A1(n7374), .A2(n6427), .ZN(n14042) );
  AND2_X1 U8592 ( .A1(n9287), .A2(n9286), .ZN(n14103) );
  NAND2_X1 U8593 ( .A1(n14100), .A2(n13914), .ZN(n14076) );
  AND2_X1 U8594 ( .A1(n9271), .A2(n9270), .ZN(n9280) );
  NOR2_X1 U8595 ( .A1(n7212), .A2(n11733), .ZN(n14120) );
  OR2_X1 U8596 ( .A1(n7215), .A2(n9486), .ZN(n7212) );
  NAND2_X1 U8597 ( .A1(n7355), .A2(n7354), .ZN(n14140) );
  NAND2_X1 U8598 ( .A1(n14616), .A2(n11216), .ZN(n11273) );
  NOR2_X1 U8599 ( .A1(n14622), .A2(n14623), .ZN(n14626) );
  NAND2_X1 U8600 ( .A1(n14626), .A2(n11275), .ZN(n11324) );
  OR2_X1 U8601 ( .A1(n11028), .A2(n11312), .ZN(n14622) );
  OR2_X1 U8602 ( .A1(n9136), .A2(n8958), .ZN(n9152) );
  NAND2_X1 U8603 ( .A1(n11019), .A2(n11018), .ZN(n11021) );
  OAI21_X1 U8604 ( .B1(n6919), .B2(n7379), .A(n7377), .ZN(n11222) );
  NAND2_X1 U8605 ( .A1(n11016), .A2(n11015), .ZN(n11017) );
  CLKBUF_X1 U8606 ( .A(n10823), .Z(n6919) );
  NAND2_X1 U8607 ( .A1(n6919), .A2(n10828), .ZN(n11016) );
  AND2_X1 U8608 ( .A1(n6406), .A2(n6444), .ZN(n6811) );
  OR2_X1 U8609 ( .A1(n9112), .A2(n9111), .ZN(n9136) );
  INV_X1 U8610 ( .A(n13782), .ZN(n11309) );
  NAND2_X1 U8611 ( .A1(n10933), .A2(n10932), .ZN(n10931) );
  AND2_X1 U8612 ( .A1(n6406), .A2(n6444), .ZN(n10943) );
  NAND2_X1 U8613 ( .A1(n10808), .A2(n10807), .ZN(n10937) );
  NOR2_X1 U8614 ( .A1(n9085), .A2(n9723), .ZN(n9094) );
  AND2_X1 U8615 ( .A1(n10592), .A2(n14646), .ZN(n10594) );
  NAND2_X1 U8616 ( .A1(n10589), .A2(n10588), .ZN(n10587) );
  NAND2_X1 U8617 ( .A1(n10634), .A2(n10633), .ZN(n10632) );
  OR2_X1 U8618 ( .A1(n9853), .A2(n9822), .ZN(n14102) );
  INV_X1 U8619 ( .A(n10021), .ZN(n6932) );
  NAND2_X1 U8620 ( .A1(n9584), .A2(n7202), .ZN(n7201) );
  OAI22_X1 U8621 ( .A1(n9526), .A2(n9525), .B1(n7399), .B2(n8983), .ZN(n7202)
         );
  OR2_X1 U8622 ( .A1(n13789), .A2(n10601), .ZN(n10083) );
  NAND2_X1 U8623 ( .A1(n13928), .A2(n14245), .ZN(n14162) );
  NAND2_X1 U8624 ( .A1(n13949), .A2(n13961), .ZN(n6944) );
  AND2_X1 U8625 ( .A1(n14105), .A2(n14658), .ZN(n14257) );
  INV_X1 U8626 ( .A(n14245), .ZN(n14672) );
  NAND2_X1 U8627 ( .A1(n11214), .A2(n11213), .ZN(n14614) );
  OR2_X1 U8628 ( .A1(n9819), .A2(n9505), .ZN(n14658) );
  INV_X1 U8629 ( .A(n14662), .ZN(n14654) );
  INV_X1 U8630 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n15232) );
  AND2_X1 U8631 ( .A1(n9531), .A2(n9530), .ZN(n9814) );
  NAND2_X1 U8632 ( .A1(n14278), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8971) );
  OAI21_X1 U8633 ( .B1(n8194), .B2(n6554), .A(n6425), .ZN(n7419) );
  OR2_X1 U8634 ( .A1(n8226), .A2(n11652), .ZN(n8227) );
  XNOR2_X1 U8635 ( .A(n8226), .B(n8210), .ZN(n13598) );
  XNOR2_X1 U8636 ( .A(n8209), .B(n8195), .ZN(n13601) );
  NAND2_X1 U8637 ( .A1(n7428), .A2(n8192), .ZN(n8209) );
  NOR2_X1 U8638 ( .A1(n7474), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n7473) );
  INV_X1 U8639 ( .A(n7474), .ZN(n7472) );
  OAI21_X1 U8640 ( .B1(n8010), .B2(n7025), .A(n7023), .ZN(n8052) );
  AND2_X1 U8641 ( .A1(n9215), .A2(n9212), .ZN(n10682) );
  XNOR2_X1 U8642 ( .A(n7971), .B(n7970), .ZN(n10059) );
  NAND2_X1 U8643 ( .A1(n7418), .A2(n7956), .ZN(n7971) );
  NAND2_X1 U8644 ( .A1(n7954), .A2(n7953), .ZN(n7418) );
  XNOR2_X1 U8645 ( .A(n7954), .B(n7953), .ZN(n9891) );
  NAND2_X1 U8646 ( .A1(n7890), .A2(n7889), .ZN(n7909) );
  INV_X1 U8647 ( .A(n6840), .ZN(n7796) );
  OAI21_X1 U8648 ( .B1(P1_ADDR_REG_1__SCAN_IN), .B2(n14309), .A(n14308), .ZN(
        n14362) );
  XNOR2_X1 U8649 ( .A(n14312), .B(n6802), .ZN(n14360) );
  XNOR2_X1 U8650 ( .A(n14357), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n14370) );
  NAND2_X1 U8651 ( .A1(n15274), .A2(n14376), .ZN(n14380) );
  INV_X1 U8652 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14377) );
  NAND2_X1 U8653 ( .A1(n14319), .A2(n14318), .ZN(n14378) );
  NAND2_X1 U8654 ( .A1(n14372), .A2(n14373), .ZN(n14318) );
  XNOR2_X1 U8655 ( .A(n15232), .B(n14321), .ZN(n14383) );
  NOR2_X1 U8656 ( .A1(n15278), .A2(n14385), .ZN(n14387) );
  NAND2_X1 U8657 ( .A1(n6795), .A2(n6434), .ZN(n14393) );
  NAND2_X1 U8658 ( .A1(n6797), .A2(n6796), .ZN(n6795) );
  OAI22_X1 U8659 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n15238), .B1(n14395), 
        .B2(n14337), .ZN(n14350) );
  OAI21_X1 U8660 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n14341), .A(n14340), .ZN(
        n14346) );
  OAI21_X1 U8661 ( .B1(n14590), .B2(n6807), .A(n6806), .ZN(n14401) );
  OR2_X1 U8662 ( .A1(n14591), .A2(n15241), .ZN(n6806) );
  AND2_X1 U8663 ( .A1(n14591), .A2(n15241), .ZN(n6807) );
  NOR2_X1 U8664 ( .A1(n6779), .A2(n12187), .ZN(n6777) );
  NOR2_X1 U8665 ( .A1(n6780), .A2(n6782), .ZN(n6779) );
  NOR2_X1 U8666 ( .A1(n12092), .A2(n12091), .ZN(n6782) );
  INV_X1 U8667 ( .A(n6783), .ZN(n6780) );
  NAND2_X1 U8668 ( .A1(n6783), .A2(n7312), .ZN(n6781) );
  AND2_X1 U8669 ( .A1(n8776), .A2(n8775), .ZN(n12676) );
  NAND2_X1 U8670 ( .A1(n11077), .A2(n11076), .ZN(n11375) );
  INV_X1 U8671 ( .A(n12123), .ZN(n7313) );
  INV_X1 U8672 ( .A(n6968), .ZN(n7314) );
  NAND2_X1 U8673 ( .A1(n11454), .A2(n11455), .ZN(n11584) );
  NAND2_X1 U8674 ( .A1(n6767), .A2(n7329), .ZN(n12141) );
  AOI21_X1 U8675 ( .B1(n7330), .B2(n11778), .A(n6494), .ZN(n7329) );
  NAND2_X1 U8676 ( .A1(n11777), .A2(n7330), .ZN(n6767) );
  NAND2_X1 U8677 ( .A1(n8643), .A2(n8642), .ZN(n12769) );
  AND3_X1 U8678 ( .A1(n8676), .A2(n8675), .A3(n8674), .ZN(n12726) );
  AOI22_X1 U8679 ( .A1(n11147), .A2(P3_REG1_REG_18__SCAN_IN), .B1(n11148), 
        .B2(P3_REG0_REG_18__SCAN_IN), .ZN(n8675) );
  INV_X1 U8680 ( .A(n12433), .ZN(n12662) );
  NAND2_X1 U8681 ( .A1(n7315), .A2(n7320), .ZN(n12166) );
  NAND2_X1 U8682 ( .A1(n12179), .A2(n7321), .ZN(n7315) );
  NAND2_X1 U8683 ( .A1(n8737), .A2(n8736), .ZN(n12694) );
  INV_X1 U8684 ( .A(n11377), .ZN(n6917) );
  INV_X1 U8685 ( .A(n6788), .ZN(n12179) );
  NAND2_X1 U8686 ( .A1(n10222), .A2(n12822), .ZN(n12185) );
  NAND2_X1 U8687 ( .A1(n10238), .A2(n10219), .ZN(n12196) );
  AND2_X1 U8688 ( .A1(n11814), .A2(n11813), .ZN(n11816) );
  NAND2_X1 U8689 ( .A1(n11814), .A2(n7330), .ZN(n12062) );
  NAND2_X1 U8690 ( .A1(n7125), .A2(n7124), .ZN(n12420) );
  NAND2_X1 U8691 ( .A1(n7126), .A2(n15056), .ZN(n7124) );
  OR2_X1 U8692 ( .A1(n7126), .A2(n8949), .ZN(n7125) );
  NAND2_X1 U8693 ( .A1(n7127), .A2(n12417), .ZN(n7126) );
  OR2_X1 U8694 ( .A1(n8846), .A2(n10706), .ZN(n12422) );
  INV_X1 U8695 ( .A(n12676), .ZN(n12135) );
  NAND2_X1 U8696 ( .A1(n11148), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8649) );
  INV_X1 U8697 ( .A(n8850), .ZN(n15068) );
  INV_X1 U8698 ( .A(n12447), .ZN(n12450) );
  NAND2_X1 U8699 ( .A1(n7260), .A2(n10709), .ZN(n10897) );
  AND2_X1 U8700 ( .A1(n7260), .A2(n7259), .ZN(n10896) );
  AOI21_X1 U8701 ( .B1(n10718), .B2(n10839), .A(n10699), .ZN(n10890) );
  NOR2_X1 U8702 ( .A1(n14854), .A2(n11488), .ZN(n14853) );
  XNOR2_X1 U8703 ( .A(n7001), .B(n14863), .ZN(n14854) );
  NOR2_X1 U8704 ( .A1(n11465), .A2(n14853), .ZN(n14873) );
  INV_X1 U8705 ( .A(n7271), .ZN(n11466) );
  INV_X1 U8706 ( .A(n7264), .ZN(n14910) );
  XNOR2_X1 U8707 ( .A(n11468), .B(n11509), .ZN(n14931) );
  INV_X1 U8708 ( .A(n7266), .ZN(n14950) );
  XNOR2_X1 U8709 ( .A(n11470), .B(n11520), .ZN(n14969) );
  NAND2_X1 U8710 ( .A1(n14990), .A2(n14991), .ZN(n14989) );
  INV_X1 U8711 ( .A(n6600), .ZN(n15004) );
  INV_X1 U8712 ( .A(n6598), .ZN(n15002) );
  INV_X1 U8713 ( .A(n7268), .ZN(n12451) );
  INV_X1 U8714 ( .A(n7270), .ZN(n11699) );
  AND2_X1 U8715 ( .A1(n7268), .A2(n7267), .ZN(n12471) );
  NOR2_X1 U8716 ( .A1(n12502), .A2(n12503), .ZN(n12521) );
  NAND2_X1 U8717 ( .A1(n7005), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7004) );
  NAND2_X1 U8718 ( .A1(n12522), .A2(n7005), .ZN(n7003) );
  INV_X1 U8719 ( .A(n12523), .ZN(n7005) );
  AND2_X1 U8720 ( .A1(n10704), .A2(n10703), .ZN(n14982) );
  INV_X1 U8721 ( .A(n6992), .ZN(n14460) );
  NAND2_X1 U8722 ( .A1(n12554), .A2(n12555), .ZN(n12576) );
  NAND2_X1 U8723 ( .A1(n6992), .A2(n6429), .ZN(n12554) );
  AND2_X1 U8724 ( .A1(n10707), .A2(n10706), .ZN(n14457) );
  NAND2_X1 U8725 ( .A1(n8827), .A2(n8826), .ZN(n12620) );
  AOI21_X1 U8726 ( .B1(n12637), .B2(n8876), .A(n8806), .ZN(n12626) );
  NAND2_X1 U8727 ( .A1(n7190), .A2(n7188), .ZN(n12842) );
  INV_X1 U8728 ( .A(n7189), .ZN(n7188) );
  NAND2_X1 U8729 ( .A1(n7191), .A2(n15051), .ZN(n7190) );
  OAI22_X1 U8730 ( .A1(n12629), .A2(n15044), .B1(n15046), .B2(n12652), .ZN(
        n7189) );
  NAND2_X1 U8731 ( .A1(n12673), .A2(n12378), .ZN(n12658) );
  NAND2_X1 U8732 ( .A1(n7176), .A2(n7178), .ZN(n12688) );
  INV_X1 U8733 ( .A(n7177), .ZN(n7176) );
  NAND2_X1 U8734 ( .A1(n7548), .A2(n12363), .ZN(n12721) );
  NAND2_X1 U8735 ( .A1(n7548), .A2(n7546), .ZN(n12873) );
  NAND2_X1 U8736 ( .A1(n8704), .A2(n8703), .ZN(n12871) );
  NAND2_X1 U8737 ( .A1(n12749), .A2(n8873), .ZN(n12739) );
  NAND2_X1 U8738 ( .A1(n12755), .A2(n7522), .ZN(n12738) );
  NAND2_X1 U8739 ( .A1(n12755), .A2(n12353), .ZN(n12736) );
  NAND2_X1 U8740 ( .A1(n8671), .A2(n8670), .ZN(n12880) );
  NAND2_X1 U8741 ( .A1(n7185), .A2(n8868), .ZN(n12763) );
  NAND2_X1 U8742 ( .A1(n14465), .A2(n8864), .ZN(n12800) );
  NAND2_X1 U8743 ( .A1(n8585), .A2(n8584), .ZN(n14484) );
  NAND2_X1 U8744 ( .A1(n11600), .A2(n12311), .ZN(n12813) );
  NAND2_X1 U8745 ( .A1(n11568), .A2(n8860), .ZN(n11611) );
  NAND2_X1 U8746 ( .A1(n11565), .A2(n12300), .ZN(n11610) );
  AND2_X1 U8747 ( .A1(n11239), .A2(n8859), .ZN(n11569) );
  NAND2_X1 U8748 ( .A1(n11118), .A2(n8858), .ZN(n11240) );
  NAND2_X1 U8749 ( .A1(n10533), .A2(n8855), .ZN(n11037) );
  INV_X1 U8750 ( .A(n15034), .ZN(n12824) );
  INV_X1 U8751 ( .A(n12280), .ZN(n15035) );
  OR2_X1 U8752 ( .A1(n12594), .A2(n8877), .ZN(n15075) );
  NAND2_X1 U8753 ( .A1(n15117), .A2(n15073), .ZN(n12900) );
  INV_X1 U8754 ( .A(n12832), .ZN(n12906) );
  INV_X1 U8755 ( .A(n12620), .ZN(n12840) );
  AOI21_X1 U8756 ( .B1(n12616), .B2(n14490), .A(n12621), .ZN(n12837) );
  INV_X1 U8757 ( .A(n12634), .ZN(n12909) );
  INV_X1 U8758 ( .A(n12388), .ZN(n12913) );
  INV_X1 U8759 ( .A(n12247), .ZN(n12917) );
  OR2_X1 U8760 ( .A1(n12862), .A2(n12861), .ZN(n12922) );
  NAND2_X1 U8761 ( .A1(n8689), .A2(n8688), .ZN(n12935) );
  AND3_X1 U8762 ( .A1(n8500), .A2(n8499), .A3(n8498), .ZN(n12299) );
  AND2_X1 U8763 ( .A1(n8483), .A2(n8481), .ZN(n6939) );
  AND2_X1 U8764 ( .A1(n8905), .A2(n8904), .ZN(n12958) );
  INV_X1 U8765 ( .A(n12959), .ZN(n12957) );
  AND2_X1 U8766 ( .A1(n10694), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12959) );
  AND2_X1 U8767 ( .A1(n7549), .A2(n6791), .ZN(n6790) );
  INV_X1 U8768 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n6791) );
  AND2_X1 U8769 ( .A1(n12208), .A2(n11854), .ZN(n12203) );
  OAI21_X1 U8770 ( .B1(n8808), .B2(n8807), .A(n8810), .ZN(n8823) );
  NAND2_X1 U8771 ( .A1(n8888), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8887) );
  NAND2_X1 U8772 ( .A1(n7158), .A2(n7157), .ZN(n8778) );
  NAND2_X1 U8773 ( .A1(n8765), .A2(n13613), .ZN(n7157) );
  NAND2_X1 U8774 ( .A1(n7153), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n7158) );
  INV_X1 U8775 ( .A(n8877), .ZN(n10404) );
  INV_X1 U8776 ( .A(SI_19_), .ZN(n10156) );
  NAND2_X1 U8777 ( .A1(n8651), .A2(n8650), .ZN(n8665) );
  INV_X1 U8778 ( .A(SI_16_), .ZN(n9686) );
  OAI21_X1 U8779 ( .B1(n8594), .B2(n7116), .A(n7114), .ZN(n8613) );
  NAND2_X1 U8780 ( .A1(n8597), .A2(n8596), .ZN(n8610) );
  NAND2_X1 U8781 ( .A1(n8594), .A2(n8593), .ZN(n8597) );
  INV_X1 U8782 ( .A(SI_12_), .ZN(n9576) );
  NAND2_X1 U8783 ( .A1(n8562), .A2(n8561), .ZN(n8579) );
  NAND2_X1 U8784 ( .A1(n8559), .A2(n8558), .ZN(n8562) );
  INV_X1 U8785 ( .A(n12454), .ZN(n12456) );
  INV_X1 U8786 ( .A(SI_11_), .ZN(n9550) );
  OR2_X1 U8787 ( .A1(n8555), .A2(n8554), .ZN(n11700) );
  INV_X1 U8788 ( .A(SI_10_), .ZN(n14409) );
  NAND2_X1 U8789 ( .A1(n8529), .A2(n8528), .ZN(n8546) );
  INV_X1 U8790 ( .A(n15009), .ZN(n14414) );
  INV_X1 U8791 ( .A(n11514), .ZN(n14957) );
  NAND2_X1 U8792 ( .A1(n7148), .A2(n7146), .ZN(n8491) );
  NAND2_X1 U8793 ( .A1(n7148), .A2(n8474), .ZN(n8477) );
  INV_X1 U8794 ( .A(n11499), .ZN(n14900) );
  INV_X1 U8795 ( .A(n11489), .ZN(n14863) );
  INV_X1 U8796 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7261) );
  OR2_X1 U8797 ( .A1(n10710), .A2(n6991), .ZN(n8398) );
  OAI211_X1 U8798 ( .C1(n8379), .C2(n8378), .A(n8381), .B(n6990), .ZN(n6913)
         );
  NAND2_X1 U8799 ( .A1(n6991), .A2(n8378), .ZN(n6990) );
  OR2_X1 U8800 ( .A1(n9520), .A2(n9519), .ZN(n9641) );
  INV_X1 U8801 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10427) );
  NAND2_X1 U8802 ( .A1(n6675), .A2(n7054), .ZN(n12054) );
  INV_X1 U8803 ( .A(n12052), .ZN(n6675) );
  AND2_X1 U8804 ( .A1(n8236), .A2(n8216), .ZN(n13282) );
  NAND2_X1 U8805 ( .A1(n11131), .A2(n11130), .ZN(n11137) );
  NAND2_X1 U8806 ( .A1(n11131), .A2(n7058), .ZN(n11258) );
  NAND2_X1 U8807 ( .A1(n7478), .A2(n10117), .ZN(n10163) );
  NAND2_X1 U8808 ( .A1(n7486), .A2(n7485), .ZN(n12984) );
  AND2_X1 U8809 ( .A1(n7486), .A2(n6450), .ZN(n12986) );
  NAND2_X1 U8810 ( .A1(n7487), .A2(n12018), .ZN(n7486) );
  NAND2_X1 U8811 ( .A1(n10743), .A2(n10742), .ZN(n10744) );
  NAND2_X1 U8812 ( .A1(n6669), .A2(n6534), .ZN(n14691) );
  NAND2_X1 U8813 ( .A1(n11131), .A2(n7055), .ZN(n6669) );
  NAND2_X1 U8814 ( .A1(n7055), .A2(n7057), .ZN(n6664) );
  NAND2_X1 U8815 ( .A1(n13039), .A2(n7501), .ZN(n13016) );
  AND2_X1 U8816 ( .A1(n7489), .A2(n10200), .ZN(n7488) );
  NAND2_X1 U8817 ( .A1(n10127), .A2(n10201), .ZN(n7490) );
  NAND2_X1 U8818 ( .A1(n13022), .A2(n12007), .ZN(n13031) );
  NOR2_X1 U8819 ( .A1(n12977), .A2(n7037), .ZN(n13041) );
  INV_X1 U8820 ( .A(n7038), .ZN(n7037) );
  NAND2_X1 U8821 ( .A1(n7491), .A2(n10125), .ZN(n10203) );
  INV_X1 U8822 ( .A(n10127), .ZN(n7491) );
  INV_X1 U8823 ( .A(n11088), .ZN(n10040) );
  OAI21_X1 U8824 ( .B1(n7055), .B2(n6667), .A(n6665), .ZN(n6668) );
  INV_X1 U8825 ( .A(n6666), .ZN(n6665) );
  XNOR2_X1 U8826 ( .A(n12035), .B(n12034), .ZN(n13057) );
  NAND2_X1 U8827 ( .A1(n11258), .A2(n11257), .ZN(n11260) );
  OAI21_X1 U8828 ( .B1(n11131), .B2(n7057), .A(n7055), .ZN(n11416) );
  NAND2_X1 U8829 ( .A1(n13030), .A2(n12013), .ZN(n13066) );
  NOR2_X1 U8830 ( .A1(n13015), .A2(n12045), .ZN(n13086) );
  INV_X1 U8831 ( .A(n14540), .ZN(n11809) );
  NAND2_X1 U8832 ( .A1(n8262), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8243) );
  INV_X1 U8833 ( .A(n12999), .ZN(n13098) );
  INV_X1 U8834 ( .A(n13257), .ZN(n13217) );
  INV_X1 U8835 ( .A(n13000), .ZN(n13256) );
  NAND2_X1 U8836 ( .A1(n8262), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8202) );
  NAND2_X1 U8837 ( .A1(n8262), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n7984) );
  NAND2_X1 U8838 ( .A1(n8262), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n7943) );
  NAND2_X1 U8839 ( .A1(n7722), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7642) );
  INV_X1 U8840 ( .A(n6612), .ZN(n14754) );
  NOR2_X1 U8841 ( .A1(n9896), .A2(n6527), .ZN(n9907) );
  AOI21_X1 U8842 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n10176), .A(n10175), .ZN(
        n10179) );
  AOI21_X1 U8843 ( .B1(n11188), .B2(P2_REG1_REG_13__SCAN_IN), .A(n14761), .ZN(
        n11191) );
  INV_X1 U8844 ( .A(n6640), .ZN(n13134) );
  NOR2_X1 U8845 ( .A1(n13129), .A2(n14783), .ZN(n14798) );
  NOR2_X1 U8846 ( .A1(n14794), .A2(n14793), .ZN(n14792) );
  INV_X1 U8847 ( .A(n13150), .ZN(n13149) );
  INV_X1 U8848 ( .A(n6637), .ZN(n13139) );
  NAND2_X1 U8849 ( .A1(n13309), .A2(n7284), .ZN(n7279) );
  OR3_X1 U8850 ( .A1(n13281), .A2(n13280), .A3(n10035), .ZN(n13456) );
  OAI21_X1 U8851 ( .B1(n13309), .B2(n7084), .A(n13251), .ZN(n13288) );
  NAND2_X1 U8852 ( .A1(n7088), .A2(n7085), .ZN(n13301) );
  INV_X1 U8853 ( .A(n13555), .ZN(n13308) );
  OAI21_X1 U8854 ( .B1(n13326), .B2(n6439), .A(n13205), .ZN(n13312) );
  NAND2_X1 U8855 ( .A1(n7273), .A2(n6467), .ZN(n13478) );
  INV_X1 U8856 ( .A(n13321), .ZN(n7278) );
  NAND2_X1 U8857 ( .A1(n7273), .A2(n7274), .ZN(n13322) );
  NAND2_X1 U8858 ( .A1(n13350), .A2(n13244), .ZN(n13333) );
  AND2_X1 U8859 ( .A1(n8132), .A2(n8131), .ZN(n13348) );
  NAND2_X1 U8860 ( .A1(n13198), .A2(n13197), .ZN(n13356) );
  NAND2_X1 U8861 ( .A1(n6701), .A2(n13238), .ZN(n13358) );
  NAND2_X1 U8862 ( .A1(n13235), .A2(n13234), .ZN(n13369) );
  NAND2_X1 U8863 ( .A1(n7291), .A2(n7289), .ZN(n13398) );
  NAND2_X1 U8864 ( .A1(n7291), .A2(n13230), .ZN(n13396) );
  INV_X1 U8865 ( .A(n13520), .ZN(n13416) );
  NAND2_X1 U8866 ( .A1(n11822), .A2(n11821), .ZN(n13421) );
  NAND2_X1 U8867 ( .A1(n11656), .A2(n11655), .ZN(n11658) );
  INV_X1 U8868 ( .A(n11656), .ZN(n11639) );
  NAND2_X1 U8869 ( .A1(n6699), .A2(n11209), .ZN(n11356) );
  NAND2_X1 U8870 ( .A1(n11207), .A2(n11206), .ZN(n6699) );
  NAND2_X1 U8871 ( .A1(n7097), .A2(n7096), .ZN(n11054) );
  NAND2_X1 U8872 ( .A1(n10781), .A2(n10780), .ZN(n10970) );
  NAND2_X1 U8873 ( .A1(n10478), .A2(n10477), .ZN(n10538) );
  NAND2_X1 U8874 ( .A1(n10476), .A2(n10475), .ZN(n10478) );
  INV_X1 U8875 ( .A(n14812), .ZN(n14531) );
  OR2_X1 U8876 ( .A1(n10501), .A2(n8286), .ZN(n13413) );
  INV_X1 U8877 ( .A(n13434), .ZN(n14815) );
  INV_X1 U8878 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6930) );
  NAND2_X1 U8879 ( .A1(n6891), .A2(n14852), .ZN(n6931) );
  NAND2_X1 U8880 ( .A1(n7978), .A2(n7977), .ZN(n14511) );
  INV_X1 U8881 ( .A(n11008), .ZN(n10190) );
  OR2_X1 U8882 ( .A1(n13454), .A2(n13531), .ZN(n6923) );
  NOR2_X1 U8883 ( .A1(n13451), .A2(n7105), .ZN(n13453) );
  OR2_X1 U8884 ( .A1(n13452), .A2(n7106), .ZN(n7105) );
  NAND2_X1 U8885 ( .A1(n6705), .A2(n6892), .ZN(n13548) );
  OR2_X1 U8886 ( .A1(n13455), .A2(n13531), .ZN(n6705) );
  AND2_X1 U8887 ( .A1(n13457), .A2(n13456), .ZN(n6892) );
  INV_X1 U8888 ( .A(n13313), .ZN(n13559) );
  AND2_X1 U8889 ( .A1(n8110), .A2(n8109), .ZN(n13567) );
  INV_X1 U8890 ( .A(n13370), .ZN(n13571) );
  AND2_X1 U8891 ( .A1(n8077), .A2(n8076), .ZN(n13575) );
  AND2_X1 U8892 ( .A1(n8027), .A2(n8026), .ZN(n13585) );
  AND2_X1 U8893 ( .A1(n9770), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14827) );
  INV_X1 U8894 ( .A(n7640), .ZN(n11845) );
  INV_X1 U8895 ( .A(n7641), .ZN(n13593) );
  NAND2_X1 U8896 ( .A1(n7072), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7296) );
  XNOR2_X1 U8897 ( .A(n8331), .B(P2_IR_REG_26__SCAN_IN), .ZN(n13603) );
  OAI21_X1 U8898 ( .B1(n8335), .B2(P2_IR_REG_25__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8331) );
  AND2_X1 U8899 ( .A1(n8334), .A2(n8335), .ZN(n13610) );
  INV_X1 U8900 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10995) );
  INV_X1 U8901 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10400) );
  INV_X1 U8902 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10349) );
  INV_X1 U8903 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10387) );
  INV_X1 U8904 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n15254) );
  INV_X1 U8905 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9892) );
  INV_X1 U8906 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9719) );
  INV_X1 U8907 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9621) );
  INV_X1 U8908 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9598) );
  INV_X1 U8909 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9600) );
  INV_X1 U8910 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9578) );
  INV_X1 U8911 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9552) );
  INV_X1 U8912 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9547) );
  INV_X1 U8913 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9538) );
  INV_X1 U8914 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9523) );
  INV_X1 U8915 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9521) );
  INV_X1 U8916 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n15142) );
  NAND2_X1 U8917 ( .A1(n13748), .A2(n11976), .ZN(n13618) );
  NAND2_X1 U8918 ( .A1(n6710), .A2(n6711), .ZN(n13617) );
  OAI21_X1 U8919 ( .B1(n11878), .B2(n7246), .A(n7244), .ZN(n11896) );
  INV_X1 U8920 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n11408) );
  NAND2_X1 U8921 ( .A1(n6709), .A2(n6708), .ZN(n11989) );
  AOI21_X1 U8922 ( .B1(n6711), .B2(n11975), .A(n11980), .ZN(n6708) );
  NAND2_X1 U8923 ( .A1(n13749), .A2(n6711), .ZN(n6709) );
  XNOR2_X1 U8924 ( .A(n11987), .B(n11986), .ZN(n11988) );
  NAND2_X1 U8925 ( .A1(n7253), .A2(n11293), .ZN(n11342) );
  INV_X1 U8926 ( .A(n10145), .ZN(n10146) );
  INV_X1 U8927 ( .A(n13788), .ZN(n10260) );
  NAND2_X1 U8928 ( .A1(n7231), .A2(n7234), .ZN(n13655) );
  NAND2_X1 U8929 ( .A1(n11878), .A2(n7247), .ZN(n13662) );
  AND2_X1 U8930 ( .A1(n11878), .A2(n11877), .ZN(n13664) );
  NAND2_X1 U8931 ( .A1(n10860), .A2(n10859), .ZN(n10997) );
  AOI21_X1 U8932 ( .B1(n13694), .B2(n13693), .A(n13692), .ZN(n13696) );
  NAND2_X1 U8933 ( .A1(n7253), .A2(n7251), .ZN(n11340) );
  NAND2_X1 U8934 ( .A1(n13662), .A2(n11887), .ZN(n13724) );
  INV_X1 U8935 ( .A(n11677), .ZN(n6719) );
  NAND2_X1 U8936 ( .A1(n9182), .A2(n9181), .ZN(n11692) );
  NAND2_X1 U8937 ( .A1(n7240), .A2(n7241), .ZN(n13743) );
  NAND2_X1 U8938 ( .A1(n9855), .A2(n9854), .ZN(n13771) );
  NAND2_X1 U8939 ( .A1(n9230), .A2(n9229), .ZN(n13887) );
  NAND2_X1 U8940 ( .A1(n14638), .A2(n9838), .ZN(n13769) );
  INV_X1 U8941 ( .A(n9474), .ZN(n6889) );
  INV_X1 U8942 ( .A(n9462), .ZN(n13879) );
  NAND2_X1 U8943 ( .A1(n6926), .A2(n9227), .ZN(n6924) );
  AOI21_X1 U8944 ( .B1(n13828), .B2(P1_REG1_REG_4__SCAN_IN), .A(n13835), .ZN(
        n9722) );
  AOI21_X1 U8945 ( .B1(n9707), .B2(P1_REG1_REG_6__SCAN_IN), .A(n9915), .ZN(
        n9949) );
  XNOR2_X1 U8946 ( .A(n11432), .B(n11442), .ZN(n14595) );
  NAND2_X1 U8947 ( .A1(n14595), .A2(n14594), .ZN(n14593) );
  NAND2_X1 U8948 ( .A1(n7208), .A2(n14151), .ZN(n7204) );
  INV_X1 U8949 ( .A(n14179), .ZN(n13982) );
  NOR2_X1 U8950 ( .A1(n13987), .A2(n7367), .ZN(n13975) );
  INV_X1 U8951 ( .A(n13922), .ZN(n14183) );
  AND2_X1 U8952 ( .A1(n13994), .A2(n7388), .ZN(n7386) );
  AND2_X1 U8953 ( .A1(n7385), .A2(n7388), .ZN(n13995) );
  NAND2_X1 U8954 ( .A1(n14201), .A2(n7390), .ZN(n13999) );
  INV_X1 U8955 ( .A(n14017), .ZN(n14197) );
  NAND2_X1 U8956 ( .A1(n6844), .A2(n13893), .ZN(n14097) );
  NAND2_X1 U8957 ( .A1(n14140), .A2(n6403), .ZN(n14244) );
  AND2_X1 U8958 ( .A1(n7348), .A2(n11725), .ZN(n11726) );
  NAND2_X1 U8959 ( .A1(n11730), .A2(n6404), .ZN(n13888) );
  NAND2_X1 U8960 ( .A1(n11552), .A2(n11547), .ZN(n11730) );
  INV_X1 U8961 ( .A(n11554), .ZN(n11552) );
  NAND2_X1 U8962 ( .A1(n9219), .A2(n9218), .ZN(n13634) );
  NAND2_X1 U8963 ( .A1(n11546), .A2(n11545), .ZN(n11724) );
  NAND2_X1 U8964 ( .A1(n11316), .A2(n11317), .ZN(n7380) );
  NAND2_X1 U8965 ( .A1(n10583), .A2(n10516), .ZN(n10517) );
  OR2_X1 U8966 ( .A1(n9832), .A2(n9831), .ZN(n14638) );
  NAND2_X1 U8967 ( .A1(n6940), .A2(n14135), .ZN(n10600) );
  INV_X1 U8968 ( .A(n14148), .ZN(n14621) );
  NOR2_X1 U8969 ( .A1(n6451), .A2(n6410), .ZN(n6643) );
  NAND2_X1 U8970 ( .A1(n6607), .A2(n6605), .ZN(n14263) );
  INV_X1 U8971 ( .A(n6606), .ZN(n6605) );
  INV_X1 U8972 ( .A(n6986), .ZN(n6607) );
  OAI21_X1 U8973 ( .B1(n14174), .B2(n14658), .A(n14173), .ZN(n6606) );
  OR3_X1 U8974 ( .A1(n14233), .A2(n14232), .A3(n14231), .ZN(n14272) );
  NAND2_X1 U8975 ( .A1(n8276), .A2(n8252), .ZN(n8255) );
  NAND2_X1 U8976 ( .A1(n8276), .A2(n8275), .ZN(n14283) );
  NAND2_X1 U8977 ( .A1(n8972), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8974) );
  NAND2_X2 U8978 ( .A1(n6621), .A2(n6619), .ZN(n13796) );
  NAND2_X1 U8979 ( .A1(n8982), .A2(n6620), .ZN(n6619) );
  AOI21_X1 U8980 ( .B1(n8982), .B2(P1_IR_REG_31__SCAN_IN), .A(
        P1_IR_REG_28__SCAN_IN), .ZN(n6618) );
  NAND2_X1 U8981 ( .A1(n9507), .A2(n6888), .ZN(n6903) );
  NOR2_X1 U8982 ( .A1(n6902), .A2(n6901), .ZN(n6900) );
  NOR2_X1 U8983 ( .A1(n6904), .A2(n9227), .ZN(n6888) );
  INV_X1 U8984 ( .A(n9816), .ZN(n14304) );
  INV_X1 U8985 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10993) );
  INV_X1 U8986 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10346) );
  INV_X1 U8987 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10405) );
  INV_X1 U8988 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10350) );
  INV_X1 U8989 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9776) );
  INV_X1 U8990 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9619) );
  INV_X1 U8991 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9603) );
  OR2_X1 U8992 ( .A1(n7870), .A2(n7869), .ZN(n7871) );
  INV_X1 U8993 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9601) );
  NAND2_X1 U8994 ( .A1(n6813), .A2(n7823), .ZN(n6812) );
  INV_X1 U8995 ( .A(n7825), .ZN(n6813) );
  INV_X1 U8996 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9580) );
  INV_X1 U8997 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9574) );
  INV_X1 U8998 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9548) );
  INV_X1 U8999 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9545) );
  INV_X1 U9000 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9540) );
  INV_X1 U9001 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9543) );
  INV_X1 U9002 ( .A(n7704), .ZN(n7701) );
  NOR2_X1 U9003 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n9051) );
  XNOR2_X1 U9004 ( .A(n14370), .B(n14746), .ZN(n15272) );
  XNOR2_X1 U9005 ( .A(n7161), .B(n14374), .ZN(n15276) );
  NAND2_X1 U9006 ( .A1(n15276), .A2(n15275), .ZN(n15274) );
  XNOR2_X1 U9007 ( .A(n14380), .B(n7160), .ZN(n14416) );
  XNOR2_X1 U9008 ( .A(n14384), .B(n14382), .ZN(n15279) );
  NOR2_X1 U9009 ( .A1(n15279), .A2(n15280), .ZN(n15278) );
  XNOR2_X1 U9010 ( .A(n14387), .B(n6981), .ZN(n14420) );
  INV_X1 U9011 ( .A(n14388), .ZN(n6981) );
  NOR2_X1 U9012 ( .A1(n14393), .A2(n14392), .ZN(n14572) );
  NAND2_X1 U9013 ( .A1(n14580), .A2(n14398), .ZN(n14583) );
  NAND2_X1 U9014 ( .A1(n14583), .A2(n14584), .ZN(n14582) );
  NAND2_X1 U9015 ( .A1(n6799), .A2(n14582), .ZN(n14588) );
  OAI21_X1 U9016 ( .B1(n14583), .B2(n14584), .A(n6800), .ZN(n6799) );
  INV_X1 U9017 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n6800) );
  NAND2_X1 U9018 ( .A1(n14588), .A2(n14587), .ZN(n14586) );
  NAND2_X1 U9019 ( .A1(n14586), .A2(n6977), .ZN(n14590) );
  OAI21_X1 U9020 ( .B1(n14588), .B2(n14587), .A(n6978), .ZN(n6977) );
  NOR2_X1 U9021 ( .A1(n14401), .A2(n14402), .ZN(n14437) );
  NAND2_X1 U9022 ( .A1(n14401), .A2(n14402), .ZN(n14439) );
  NAND2_X1 U9023 ( .A1(n14439), .A2(n14440), .ZN(n14436) );
  OAI211_X1 U9024 ( .C1(n12189), .C2(n6778), .A(n6937), .B(n6776), .ZN(
        P3_U3154) );
  AND2_X1 U9025 ( .A1(n12096), .A2(n6539), .ZN(n6937) );
  NAND2_X1 U9026 ( .A1(n6781), .A2(n12192), .ZN(n6778) );
  NAND2_X1 U9027 ( .A1(n12189), .A2(n6777), .ZN(n6776) );
  NAND2_X1 U9028 ( .A1(n10371), .A2(n10370), .ZN(n10377) );
  XNOR2_X1 U9029 ( .A(n6597), .B(n12585), .ZN(n12599) );
  OAI21_X1 U9030 ( .B1(n6992), .B2(n6596), .A(n6594), .ZN(n6597) );
  NOR2_X1 U9031 ( .A1(n6531), .A2(n7536), .ZN(n7535) );
  NAND2_X1 U9032 ( .A1(n7531), .A2(n7530), .ZN(n7532) );
  NAND2_X1 U9033 ( .A1(n7534), .A2(n15117), .ZN(n7533) );
  NOR2_X1 U9034 ( .A1(n6526), .A2(n8943), .ZN(n8944) );
  NAND2_X1 U9035 ( .A1(n7050), .A2(n14692), .ZN(n7048) );
  AOI22_X1 U9036 ( .A1(n9984), .A2(n14694), .B1(n14697), .B2(n9736), .ZN(n9774) );
  NOR2_X1 U9037 ( .A1(n8309), .A2(n8301), .ZN(n8341) );
  MUX2_X1 U9038 ( .A(n13176), .B(n13175), .S(n13174), .Z(n13178) );
  OAI21_X1 U9039 ( .B1(n13449), .B2(n13434), .A(n7292), .ZN(P2_U3236) );
  NAND2_X1 U9040 ( .A1(n7013), .A2(n6405), .ZN(n13449) );
  INV_X1 U9041 ( .A(n7293), .ZN(n7292) );
  NAND2_X1 U9042 ( .A1(n7009), .A2(n6405), .ZN(n7020) );
  AND2_X1 U9043 ( .A1(n7013), .A2(n14845), .ZN(n7009) );
  OAI21_X1 U9044 ( .B1(n11860), .B2(n14846), .A(n7064), .ZN(P2_U3498) );
  INV_X1 U9045 ( .A(n7065), .ZN(n7064) );
  OAI22_X1 U9046 ( .A1(n11868), .A2(n13584), .B1(n14848), .B2(n11859), .ZN(
        n7065) );
  AOI21_X1 U9047 ( .B1(n7011), .B2(n6405), .A(n6553), .ZN(n7010) );
  AND2_X1 U9048 ( .A1(n10327), .A2(n10326), .ZN(n10335) );
  NAND2_X1 U9049 ( .A1(n13793), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7254) );
  MUX2_X1 U9050 ( .A(n13876), .B(n13875), .S(n9505), .Z(n13877) );
  NAND2_X1 U9051 ( .A1(n13971), .A2(n6608), .ZN(P1_U3266) );
  NAND2_X1 U9052 ( .A1(n6986), .A2(n14613), .ZN(n6608) );
  NAND2_X1 U9053 ( .A1(n6642), .A2(n6641), .ZN(P1_U3556) );
  NAND2_X1 U9054 ( .A1(n14685), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6641) );
  NAND2_X1 U9055 ( .A1(n14262), .A2(n14687), .ZN(n6642) );
  NAND2_X1 U9056 ( .A1(n6809), .A2(n6808), .ZN(P1_U3524) );
  NAND2_X1 U9057 ( .A1(n14678), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6808) );
  NAND2_X1 U9058 ( .A1(n14262), .A2(n14679), .ZN(n6809) );
  NOR2_X1 U9059 ( .A1(n14426), .A2(n14427), .ZN(n14425) );
  XNOR2_X1 U9060 ( .A(n6794), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  OAI21_X1 U9061 ( .B1(n14442), .B2(n14441), .A(n14443), .ZN(n6794) );
  XNOR2_X1 U9062 ( .A(n7163), .B(n7162), .ZN(SUB_1596_U4) );
  XNOR2_X1 U9063 ( .A(n14449), .B(n6566), .ZN(n7162) );
  NAND2_X1 U9064 ( .A1(n14443), .A2(n7164), .ZN(n7163) );
  CLKBUF_X3 U9065 ( .A(n8242), .Z(n8284) );
  NAND2_X4 U9066 ( .A1(n6707), .A2(n9841), .ZN(n10140) );
  AND2_X1 U9067 ( .A1(n14127), .A2(n13911), .ZN(n6403) );
  AND2_X1 U9068 ( .A1(n11732), .A2(n11729), .ZN(n6404) );
  NAND2_X1 U9069 ( .A1(n9584), .A2(n9533), .ZN(n9217) );
  OR3_X1 U9070 ( .A1(n13260), .A2(n13261), .A3(n13258), .ZN(n6405) );
  AND2_X1 U9071 ( .A1(n10592), .A2(n7203), .ZN(n6406) );
  XNOR2_X1 U9072 ( .A(n14171), .B(n13942), .ZN(n13958) );
  INV_X1 U9073 ( .A(n13958), .ZN(n7360) );
  AND2_X1 U9074 ( .A1(n9093), .A2(n7464), .ZN(n6407) );
  INV_X1 U9075 ( .A(n10076), .ZN(n7255) );
  INV_X1 U9076 ( .A(n7907), .ZN(n6580) );
  NAND2_X1 U9077 ( .A1(n8191), .A2(n8190), .ZN(n7579) );
  INV_X1 U9078 ( .A(n7579), .ZN(n7577) );
  INV_X1 U9079 ( .A(n14143), .ZN(n7354) );
  NAND2_X1 U9080 ( .A1(n7961), .A2(n7960), .ZN(n11636) );
  AND2_X1 U9081 ( .A1(n12441), .A2(n15095), .ZN(n6408) );
  AND2_X1 U9082 ( .A1(n7969), .A2(n7968), .ZN(n6409) );
  OAI21_X1 U9083 ( .B1(n12080), .B2(n12159), .A(n6784), .ZN(n12130) );
  AND2_X1 U9084 ( .A1(n14167), .A2(n14653), .ZN(n6410) );
  AND3_X1 U9085 ( .A1(n6747), .A2(n7568), .A3(n6522), .ZN(n6411) );
  INV_X1 U9086 ( .A(n11778), .ZN(n7331) );
  AND2_X1 U9087 ( .A1(n11722), .A2(n11725), .ZN(n11553) );
  NAND2_X1 U9088 ( .A1(n9313), .A2(n9312), .ZN(n14212) );
  INV_X1 U9089 ( .A(n14212), .ZN(n6818) );
  NAND2_X1 U9090 ( .A1(n8991), .A2(n8990), .ZN(n14132) );
  AND2_X1 U9091 ( .A1(n6627), .A2(n6724), .ZN(n6412) );
  AND2_X1 U9092 ( .A1(n7051), .A2(n7049), .ZN(n6413) );
  NAND2_X1 U9093 ( .A1(n6830), .A2(n9214), .ZN(n14562) );
  AND2_X1 U9094 ( .A1(n6436), .A2(n7025), .ZN(n6414) );
  AND2_X1 U9095 ( .A1(n9269), .A2(n9268), .ZN(n14110) );
  INV_X1 U9096 ( .A(n14110), .ZN(n14237) );
  AND2_X1 U9097 ( .A1(n7986), .A2(n6465), .ZN(n6415) );
  AND2_X1 U9098 ( .A1(n7456), .A2(n9183), .ZN(n6416) );
  NOR2_X1 U9099 ( .A1(n13336), .A2(n13245), .ZN(n6417) );
  AND2_X1 U9100 ( .A1(n12378), .A2(n12379), .ZN(n12670) );
  NAND2_X1 U9101 ( .A1(n6735), .A2(n6519), .ZN(n6418) );
  OR2_X1 U9102 ( .A1(n8086), .A2(n8084), .ZN(n6419) );
  INV_X1 U9103 ( .A(n13715), .ZN(n7232) );
  AND2_X1 U9104 ( .A1(n10859), .A2(n10864), .ZN(n6420) );
  AND2_X1 U9105 ( .A1(n7236), .A2(n6537), .ZN(n6421) );
  INV_X1 U9106 ( .A(n7216), .ZN(n7215) );
  NOR2_X1 U9107 ( .A1(n14132), .A2(n13887), .ZN(n7216) );
  AND2_X1 U9108 ( .A1(n7664), .A2(n7663), .ZN(n9863) );
  INV_X1 U9109 ( .A(n9863), .ZN(n7505) );
  INV_X1 U9110 ( .A(n11504), .ZN(n14919) );
  OR2_X1 U9111 ( .A1(n11733), .A2(n13887), .ZN(n6422) );
  AND2_X1 U9112 ( .A1(n13520), .A2(n13231), .ZN(n6423) );
  XNOR2_X1 U9113 ( .A(n9010), .B(n9009), .ZN(n9505) );
  INV_X1 U9114 ( .A(n13073), .ZN(n14692) );
  INV_X1 U9115 ( .A(n11348), .ZN(n6810) );
  INV_X2 U9116 ( .A(n15114), .ZN(n15117) );
  AND2_X1 U9117 ( .A1(n8257), .A2(n7433), .ZN(n6424) );
  NAND2_X1 U9118 ( .A1(n14626), .A2(n6820), .ZN(n11548) );
  INV_X1 U9119 ( .A(n11548), .ZN(n6825) );
  OR2_X1 U9120 ( .A1(n7424), .A2(SI_27_), .ZN(n6425) );
  NOR2_X1 U9121 ( .A1(n7426), .A2(SI_27_), .ZN(n6426) );
  INV_X1 U9122 ( .A(n7722), .ZN(n8116) );
  OR2_X1 U9123 ( .A1(n14080), .A2(n13899), .ZN(n6427) );
  NAND4_X1 U9124 ( .A1(n7643), .A2(n7642), .A3(n7644), .A4(n7645), .ZN(n8313)
         );
  NOR2_X1 U9125 ( .A1(n12700), .A2(n12373), .ZN(n7177) );
  AND3_X1 U9126 ( .A1(n10710), .A2(n8342), .A3(n7182), .ZN(n8445) );
  INV_X1 U9127 ( .A(n11257), .ZN(n7057) );
  INV_X1 U9128 ( .A(n12051), .ZN(n7054) );
  INV_X1 U9129 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n6991) );
  INV_X1 U9130 ( .A(n8170), .ZN(n6922) );
  AND2_X1 U9131 ( .A1(n7483), .A2(n7042), .ZN(n6428) );
  INV_X1 U9132 ( .A(n11231), .ZN(n12443) );
  OR2_X1 U9133 ( .A1(n12553), .A2(n14450), .ZN(n6429) );
  AND2_X1 U9134 ( .A1(n8364), .A2(n8365), .ZN(n8402) );
  AND2_X1 U9135 ( .A1(n7231), .A2(n7229), .ZN(n6430) );
  AND2_X1 U9136 ( .A1(n12843), .A2(n14490), .ZN(n6431) );
  OR2_X1 U9137 ( .A1(n6390), .A2(n6913), .ZN(n6432) );
  AND2_X1 U9138 ( .A1(n7240), .A2(n7238), .ZN(n6433) );
  OR2_X1 U9139 ( .A1(n14427), .A2(n6798), .ZN(n6434) );
  AND2_X1 U9140 ( .A1(n14813), .A2(n7068), .ZN(n6435) );
  INV_X1 U9141 ( .A(n13550), .ZN(n13255) );
  INV_X1 U9142 ( .A(n11657), .ZN(n11824) );
  XNOR2_X1 U9143 ( .A(n14540), .B(n13100), .ZN(n11657) );
  XNOR2_X1 U9144 ( .A(n13079), .B(n6687), .ZN(n10477) );
  INV_X1 U9145 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8375) );
  OR2_X1 U9146 ( .A1(n8051), .A2(SI_17_), .ZN(n6436) );
  INV_X1 U9147 ( .A(n13258), .ZN(n7295) );
  XNOR2_X1 U9148 ( .A(n13446), .B(n13098), .ZN(n13258) );
  OR2_X1 U9149 ( .A1(n13153), .A2(n13152), .ZN(n6437) );
  OR2_X1 U9150 ( .A1(n8100), .A2(n8101), .ZN(n6438) );
  NOR2_X1 U9151 ( .A1(n13336), .A2(n13204), .ZN(n6439) );
  AND2_X1 U9152 ( .A1(n12024), .A2(n12018), .ZN(n6440) );
  OR2_X1 U9153 ( .A1(n7904), .A2(n6461), .ZN(n6441) );
  OR2_X1 U9154 ( .A1(n8834), .A2(n8359), .ZN(n6442) );
  OR2_X1 U9155 ( .A1(n7950), .A2(n7949), .ZN(n6443) );
  AOI21_X1 U9156 ( .B1(n12035), .B2(n6678), .A(n6677), .ZN(n12037) );
  XNOR2_X1 U9157 ( .A(n6792), .B(P3_IR_REG_30__SCAN_IN), .ZN(n8364) );
  AND2_X1 U9158 ( .A1(n10848), .A2(n14646), .ZN(n6444) );
  NAND2_X1 U9159 ( .A1(n9007), .A2(n7444), .ZN(n9816) );
  NAND2_X1 U9160 ( .A1(n12694), .A2(n12435), .ZN(n6445) );
  INV_X1 U9161 ( .A(n10331), .ZN(n6936) );
  OR2_X1 U9162 ( .A1(n7710), .A2(n7709), .ZN(n10107) );
  INV_X1 U9163 ( .A(n10107), .ZN(n6896) );
  AND2_X1 U9164 ( .A1(n7512), .A2(n7510), .ZN(n6446) );
  INV_X1 U9165 ( .A(n9458), .ZN(n14151) );
  NAND2_X1 U9166 ( .A1(n9456), .A2(n9455), .ZN(n9458) );
  OAI22_X1 U9167 ( .A1(n13550), .A2(n8284), .B1(n7768), .B2(n13000), .ZN(n8222) );
  INV_X1 U9168 ( .A(n8222), .ZN(n6745) );
  AND2_X1 U9169 ( .A1(n12997), .A2(n12993), .ZN(n6447) );
  OR2_X1 U9170 ( .A1(n12629), .A2(n12840), .ZN(n6448) );
  NAND2_X1 U9171 ( .A1(n9351), .A2(n9350), .ZN(n14193) );
  INV_X1 U9172 ( .A(n14193), .ZN(n14012) );
  AOI21_X1 U9173 ( .B1(n12059), .B2(n12431), .A(n12110), .ZN(n12092) );
  INV_X1 U9174 ( .A(n12092), .ZN(n7312) );
  INV_X1 U9175 ( .A(n11570), .ZN(n12297) );
  INV_X1 U9176 ( .A(n7932), .ZN(n7031) );
  XNOR2_X1 U9177 ( .A(n12037), .B(n12036), .ZN(n12976) );
  AND2_X1 U9178 ( .A1(n10710), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7262) );
  XNOR2_X1 U9179 ( .A(n13308), .B(n13250), .ZN(n13249) );
  OR3_X1 U9180 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n6449) );
  NAND2_X1 U9181 ( .A1(n12017), .A2(n12016), .ZN(n6450) );
  INV_X1 U9182 ( .A(n9133), .ZN(n6854) );
  AND2_X1 U9183 ( .A1(n14168), .A2(n14654), .ZN(n6451) );
  AND2_X1 U9184 ( .A1(n9301), .A2(n9300), .ZN(n14218) );
  INV_X1 U9185 ( .A(n14218), .ZN(n13899) );
  AND2_X1 U9186 ( .A1(n14242), .A2(n14136), .ZN(n6452) );
  AND2_X1 U9187 ( .A1(n8212), .A2(n8211), .ZN(n13550) );
  NAND2_X1 U9188 ( .A1(n11415), .A2(n11414), .ZN(n6453) );
  NAND2_X1 U9189 ( .A1(n14242), .A2(n13892), .ZN(n6454) );
  NOR2_X1 U9190 ( .A1(n12408), .A2(n12415), .ZN(n6455) );
  AND3_X1 U9191 ( .A1(n7696), .A2(n7694), .A3(n7697), .ZN(n6456) );
  AND2_X1 U9192 ( .A1(n13274), .A2(n7284), .ZN(n6457) );
  AND2_X1 U9193 ( .A1(n12814), .A2(n8862), .ZN(n6458) );
  AND2_X1 U9194 ( .A1(n8233), .A2(n8232), .ZN(n13265) );
  INV_X1 U9195 ( .A(n13265), .ZN(n7062) );
  XNOR2_X1 U9196 ( .A(n8398), .B(n7261), .ZN(n11463) );
  NAND2_X1 U9197 ( .A1(n8342), .A2(n8380), .ZN(n8422) );
  NAND2_X1 U9198 ( .A1(n7708), .A2(n7706), .ZN(n7736) );
  OR2_X1 U9199 ( .A1(n7969), .A2(n7968), .ZN(n7591) );
  INV_X1 U9200 ( .A(n7591), .ZN(n6761) );
  AND2_X1 U9201 ( .A1(n7838), .A2(n7837), .ZN(n6459) );
  OR2_X1 U9202 ( .A1(n12694), .A2(n12435), .ZN(n6460) );
  AND2_X1 U9203 ( .A1(n7902), .A2(n7901), .ZN(n6461) );
  AND2_X1 U9204 ( .A1(n14070), .A2(n6427), .ZN(n6462) );
  AND2_X1 U9205 ( .A1(n7243), .A2(n7242), .ZN(n6463) );
  NOR2_X1 U9206 ( .A1(n12521), .A2(n12522), .ZN(n6464) );
  NOR2_X1 U9207 ( .A1(n12740), .A2(n7194), .ZN(n7193) );
  OR2_X1 U9208 ( .A1(n8035), .A2(n7590), .ZN(n6465) );
  INV_X1 U9209 ( .A(n6826), .ZN(n13964) );
  OR2_X1 U9210 ( .A1(n13976), .A2(n14171), .ZN(n6826) );
  AND2_X1 U9211 ( .A1(n8174), .A2(n7422), .ZN(n6466) );
  AND2_X1 U9212 ( .A1(n7278), .A2(n7274), .ZN(n6467) );
  AND2_X1 U9213 ( .A1(n8982), .A2(n6924), .ZN(n6468) );
  AND2_X1 U9214 ( .A1(n12817), .A2(n12311), .ZN(n6469) );
  AND2_X1 U9215 ( .A1(n8260), .A2(n8259), .ZN(n13225) );
  INV_X1 U9216 ( .A(n13225), .ZN(n13446) );
  AND2_X1 U9217 ( .A1(n7368), .A2(n7372), .ZN(n6470) );
  OR2_X1 U9218 ( .A1(n13261), .A2(n13274), .ZN(n6471) );
  NOR2_X1 U9219 ( .A1(n13246), .A2(n7276), .ZN(n7275) );
  AND2_X1 U9220 ( .A1(n10910), .A2(n12442), .ZN(n6472) );
  AND2_X1 U9221 ( .A1(n12306), .A2(n12307), .ZN(n6473) );
  AND2_X1 U9222 ( .A1(n7023), .A2(n6436), .ZN(n6474) );
  NAND2_X1 U9223 ( .A1(n8987), .A2(n7473), .ZN(n9001) );
  NOR2_X1 U9224 ( .A1(n8300), .A2(n8299), .ZN(n6475) );
  INV_X1 U9225 ( .A(n7557), .ZN(n7556) );
  OAI21_X1 U9226 ( .B1(n8295), .B2(n7604), .A(n6475), .ZN(n7557) );
  AND2_X1 U9227 ( .A1(n7357), .A2(n11018), .ZN(n6476) );
  OR2_X1 U9228 ( .A1(n13923), .A2(n14183), .ZN(n6477) );
  AND2_X1 U9229 ( .A1(n8002), .A2(n8007), .ZN(n6478) );
  INV_X1 U9230 ( .A(n7391), .ZN(n7390) );
  AND2_X1 U9231 ( .A1(n11725), .A2(n11731), .ZN(n6479) );
  AND2_X1 U9232 ( .A1(n12673), .A2(n7541), .ZN(n6480) );
  INV_X1 U9233 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9227) );
  AND2_X1 U9234 ( .A1(n11815), .A2(n11813), .ZN(n7330) );
  INV_X1 U9235 ( .A(n10128), .ZN(n10125) );
  XNOR2_X1 U9236 ( .A(n10198), .B(n10197), .ZN(n10128) );
  NAND2_X1 U9237 ( .A1(n7313), .A2(n7316), .ZN(n6481) );
  NOR2_X1 U9238 ( .A1(n13982), .A2(n13962), .ZN(n6482) );
  NOR2_X1 U9239 ( .A1(n11359), .A2(n14523), .ZN(n6483) );
  NOR2_X1 U9240 ( .A1(n13079), .A2(n13107), .ZN(n6484) );
  INV_X1 U9241 ( .A(n7019), .ZN(n7018) );
  NOR2_X1 U9242 ( .A1(n13265), .A2(n13257), .ZN(n7019) );
  OR2_X1 U9243 ( .A1(n8035), .A2(n6761), .ZN(n6485) );
  NOR2_X1 U9244 ( .A1(n11053), .A2(n11052), .ZN(n6486) );
  NOR2_X1 U9245 ( .A1(n13661), .A2(n11882), .ZN(n6487) );
  NOR2_X1 U9246 ( .A1(n11400), .A2(n11399), .ZN(n6488) );
  NOR2_X1 U9247 ( .A1(n12880), .A2(n12752), .ZN(n6489) );
  NOR2_X1 U9248 ( .A1(n13887), .A2(n14134), .ZN(n6490) );
  INV_X1 U9249 ( .A(n13292), .ZN(n13460) );
  INV_X1 U9250 ( .A(n7322), .ZN(n7321) );
  NAND2_X1 U9251 ( .A1(n7325), .A2(n7326), .ZN(n7322) );
  NAND2_X1 U9252 ( .A1(n8996), .A2(n8997), .ZN(n11354) );
  INV_X1 U9253 ( .A(n7175), .ZN(n7174) );
  AND2_X1 U9254 ( .A1(n6460), .A2(n7178), .ZN(n7175) );
  NAND2_X1 U9255 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_24__SCAN_IN), 
        .ZN(n6491) );
  OR2_X1 U9256 ( .A1(n9401), .A2(n9402), .ZN(n6492) );
  NAND2_X1 U9257 ( .A1(n13585), .A2(n13099), .ZN(n6493) );
  AND2_X1 U9258 ( .A1(n12061), .A2(n12437), .ZN(n6494) );
  NAND2_X1 U9259 ( .A1(n14171), .A2(n13924), .ZN(n6495) );
  AND2_X1 U9260 ( .A1(n14303), .A2(n9584), .ZN(n14206) );
  INV_X1 U9261 ( .A(n14206), .ZN(n14033) );
  INV_X1 U9262 ( .A(n6817), .ZN(n6816) );
  NAND2_X1 U9263 ( .A1(n14033), .A2(n6818), .ZN(n6817) );
  INV_X1 U9264 ( .A(n6822), .ZN(n6821) );
  NAND2_X1 U9265 ( .A1(n11275), .A2(n6823), .ZN(n6822) );
  INV_X1 U9266 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n6926) );
  INV_X1 U9267 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8911) );
  AND2_X1 U9268 ( .A1(n7972), .A2(n9596), .ZN(n6496) );
  AND2_X1 U9269 ( .A1(n14033), .A2(n14043), .ZN(n6497) );
  NAND2_X1 U9270 ( .A1(n13241), .A2(n13240), .ZN(n13349) );
  INV_X1 U9271 ( .A(n13349), .ZN(n7277) );
  NAND2_X1 U9272 ( .A1(n13255), .A2(n13256), .ZN(n6498) );
  AOI21_X1 U9273 ( .B1(n7229), .B2(n13715), .A(n13733), .ZN(n7227) );
  OR2_X1 U9274 ( .A1(n12620), .A2(n12629), .ZN(n8941) );
  OR2_X1 U9275 ( .A1(n7795), .A2(SI_6_), .ZN(n6499) );
  INV_X1 U9276 ( .A(n9478), .ZN(n14084) );
  AND2_X1 U9277 ( .A1(n9291), .A2(n13915), .ZN(n9478) );
  INV_X1 U9278 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8979) );
  NAND2_X1 U9279 ( .A1(n7323), .A2(n12103), .ZN(n6500) );
  INV_X1 U9280 ( .A(n7208), .ZN(n7207) );
  NAND2_X1 U9281 ( .A1(n14156), .A2(n7209), .ZN(n7208) );
  INV_X1 U9282 ( .A(n9352), .ZN(n6852) );
  INV_X1 U9283 ( .A(n13882), .ZN(n14156) );
  NAND2_X1 U9284 ( .A1(n9442), .A2(n9441), .ZN(n13882) );
  INV_X1 U9285 ( .A(n9184), .ZN(n7456) );
  OR2_X1 U9286 ( .A1(n13949), .A2(n13961), .ZN(n6501) );
  AND2_X1 U9287 ( .A1(n11587), .A2(n12439), .ZN(n6502) );
  AND2_X1 U9288 ( .A1(n11585), .A2(n12801), .ZN(n6503) );
  AND2_X1 U9289 ( .A1(n12290), .A2(n12289), .ZN(n12226) );
  INV_X1 U9290 ( .A(n11215), .ZN(n14617) );
  OR2_X1 U9291 ( .A1(n7861), .A2(n7860), .ZN(n6504) );
  OR2_X1 U9292 ( .A1(n11476), .A2(n10713), .ZN(n6505) );
  OR2_X1 U9293 ( .A1(n13447), .A2(n14846), .ZN(n6506) );
  AND2_X1 U9294 ( .A1(n7791), .A2(n7790), .ZN(n6507) );
  NOR2_X1 U9295 ( .A1(n9479), .A2(n9459), .ZN(n6508) );
  NOR2_X1 U9296 ( .A1(n14562), .A2(n13777), .ZN(n6509) );
  NOR2_X1 U9297 ( .A1(n11312), .A2(n13781), .ZN(n6510) );
  NOR2_X1 U9298 ( .A1(n11681), .A2(n11680), .ZN(n6511) );
  AND2_X1 U9299 ( .A1(n11553), .A2(n13777), .ZN(n6512) );
  AND2_X1 U9300 ( .A1(n7373), .A2(n6427), .ZN(n6513) );
  AND2_X1 U9301 ( .A1(n6748), .A2(n6745), .ZN(n6514) );
  NOR2_X1 U9302 ( .A1(n14590), .A2(n14591), .ZN(n6515) );
  AND2_X1 U9303 ( .A1(n6967), .A2(n12080), .ZN(n6516) );
  AND2_X1 U9304 ( .A1(n7319), .A2(n7320), .ZN(n6517) );
  INV_X1 U9305 ( .A(n7281), .ZN(n13274) );
  XNOR2_X1 U9306 ( .A(n13550), .B(n13000), .ZN(n7281) );
  INV_X1 U9307 ( .A(n7552), .ZN(n7551) );
  NOR2_X1 U9308 ( .A1(n8359), .A2(P3_IR_REG_27__SCAN_IN), .ZN(n7552) );
  AND2_X1 U9309 ( .A1(n13265), .A2(n13550), .ZN(n6518) );
  AND2_X1 U9310 ( .A1(n6441), .A2(n6737), .ZN(n6519) );
  NAND2_X1 U9311 ( .A1(n12634), .A2(n12641), .ZN(n12396) );
  AND2_X1 U9312 ( .A1(n7207), .A2(n9458), .ZN(n6520) );
  INV_X1 U9313 ( .A(n7104), .ZN(n7103) );
  NAND2_X1 U9314 ( .A1(n13261), .A2(n13262), .ZN(n7104) );
  NAND2_X1 U9315 ( .A1(n9476), .A2(n9460), .ZN(n6521) );
  OR2_X1 U9316 ( .A1(n6748), .A2(n6745), .ZN(n6522) );
  NAND2_X1 U9317 ( .A1(n9340), .A2(n7460), .ZN(n6523) );
  AND2_X1 U9318 ( .A1(n8354), .A2(n7339), .ZN(n6524) );
  INV_X1 U9319 ( .A(n9151), .ZN(n7471) );
  AND2_X1 U9320 ( .A1(n8189), .A2(n7581), .ZN(n7580) );
  NAND2_X1 U9321 ( .A1(n9352), .A2(n9355), .ZN(n6850) );
  INV_X1 U9322 ( .A(n7604), .ZN(n7558) );
  INV_X1 U9323 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6973) );
  INV_X1 U9324 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n8973) );
  NAND2_X1 U9325 ( .A1(n7770), .A2(n7588), .ZN(n7587) );
  NAND2_X1 U9326 ( .A1(n6706), .A2(n9531), .ZN(n9841) );
  AND2_X1 U9327 ( .A1(n9133), .A2(n6855), .ZN(n6525) );
  OR2_X1 U9328 ( .A1(n12253), .A2(n10404), .ZN(n12244) );
  INV_X1 U9329 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n7339) );
  INV_X1 U9330 ( .A(n7726), .ZN(n8246) );
  NAND2_X1 U9331 ( .A1(n8146), .A2(n8145), .ZN(n13336) );
  INV_X1 U9332 ( .A(n13336), .ZN(n7069) );
  AND2_X1 U9333 ( .A1(n7297), .A2(n11579), .ZN(n8892) );
  NAND2_X1 U9334 ( .A1(n8987), .A2(n8986), .ZN(n8992) );
  AND2_X1 U9335 ( .A1(n9022), .A2(n9021), .ZN(n14242) );
  INV_X1 U9336 ( .A(n14242), .ZN(n9486) );
  NAND2_X1 U9337 ( .A1(n11596), .A2(n6458), .ZN(n12815) );
  NOR2_X1 U9338 ( .A1(n8957), .A2(n12955), .ZN(n6526) );
  NAND2_X1 U9339 ( .A1(n11278), .A2(n11277), .ZN(n11316) );
  AND2_X1 U9340 ( .A1(n9899), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6527) );
  OAI21_X1 U9341 ( .B1(n7496), .B2(n7045), .A(n6428), .ZN(n13051) );
  AND2_X1 U9342 ( .A1(n14957), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n6528) );
  NAND2_X1 U9343 ( .A1(n12792), .A2(n12334), .ZN(n12780) );
  NAND2_X1 U9344 ( .A1(n7380), .A2(n11280), .ZN(n11551) );
  OR2_X1 U9345 ( .A1(n12909), .A2(n12955), .ZN(n6529) );
  INV_X1 U9346 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8356) );
  NAND2_X1 U9347 ( .A1(n6815), .A2(n6814), .ZN(n6819) );
  NOR2_X1 U9348 ( .A1(n11733), .A2(n7215), .ZN(n6530) );
  INV_X1 U9349 ( .A(n7351), .ZN(n14098) );
  NAND2_X1 U9350 ( .A1(n11797), .A2(n11796), .ZN(n14505) );
  NOR2_X1 U9351 ( .A1(n8957), .A2(n12900), .ZN(n6531) );
  AND2_X1 U9352 ( .A1(n11730), .A2(n11729), .ZN(n6532) );
  AND2_X1 U9353 ( .A1(n12749), .A2(n7193), .ZN(n6533) );
  AND2_X1 U9354 ( .A1(n6664), .A2(n6453), .ZN(n6534) );
  INV_X1 U9355 ( .A(n7211), .ZN(n14049) );
  NOR2_X1 U9356 ( .A1(n14067), .A2(n14212), .ZN(n7211) );
  AND2_X1 U9357 ( .A1(n14484), .A2(n12438), .ZN(n6535) );
  INV_X1 U9358 ( .A(n8069), .ZN(n7407) );
  OR2_X1 U9359 ( .A1(n13550), .A2(n13541), .ZN(n6536) );
  NAND2_X1 U9360 ( .A1(n11933), .A2(n11934), .ZN(n6537) );
  INV_X1 U9361 ( .A(n6819), .ZN(n7210) );
  INV_X1 U9362 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7399) );
  AND2_X1 U9363 ( .A1(n6723), .A2(n7236), .ZN(n6538) );
  OR2_X1 U9364 ( .A1(n12909), .A2(n12201), .ZN(n6539) );
  AND2_X1 U9365 ( .A1(n8051), .A2(SI_17_), .ZN(n6540) );
  OR2_X1 U9366 ( .A1(n13550), .A2(n13584), .ZN(n6541) );
  NAND2_X1 U9367 ( .A1(n8745), .A2(n8744), .ZN(n12435) );
  INV_X1 U9368 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6616) );
  AND2_X1 U9369 ( .A1(n7609), .A2(n7606), .ZN(n6542) );
  INV_X1 U9370 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10060) );
  OR2_X1 U9371 ( .A1(n7265), .A2(n6528), .ZN(n6543) );
  AND2_X1 U9372 ( .A1(n14140), .A2(n13911), .ZN(n6544) );
  INV_X1 U9373 ( .A(n14132), .ZN(n7217) );
  AND2_X1 U9374 ( .A1(n8916), .A2(n8915), .ZN(n15110) );
  INV_X1 U9375 ( .A(n13226), .ZN(n7287) );
  INV_X1 U9376 ( .A(n9505), .ZN(n14008) );
  NAND2_X1 U9377 ( .A1(n7490), .A2(n7488), .ZN(n10411) );
  NAND2_X1 U9378 ( .A1(n9195), .A2(n9194), .ZN(n13661) );
  INV_X1 U9379 ( .A(n13661), .ZN(n6823) );
  AND2_X1 U9380 ( .A1(n10743), .A2(n7481), .ZN(n6545) );
  INV_X1 U9381 ( .A(n12187), .ZN(n12192) );
  AND2_X1 U9382 ( .A1(n6811), .A2(n10925), .ZN(n6546) );
  INV_X1 U9383 ( .A(n11698), .ZN(n7269) );
  OR2_X1 U9384 ( .A1(n14848), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6547) );
  INV_X1 U9385 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6632) );
  AND2_X1 U9386 ( .A1(n8701), .A2(n7123), .ZN(n6548) );
  NAND2_X1 U9387 ( .A1(n11596), .A2(n8862), .ZN(n6549) );
  NAND2_X1 U9388 ( .A1(n14626), .A2(n6821), .ZN(n6550) );
  NAND2_X1 U9389 ( .A1(n6825), .A2(n6824), .ZN(n11733) );
  OR2_X1 U9390 ( .A1(n15009), .A2(n11606), .ZN(n6551) );
  INV_X1 U9391 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7160) );
  AND2_X1 U9392 ( .A1(n7097), .A2(n10791), .ZN(n6552) );
  NOR2_X1 U9393 ( .A1(n14848), .A2(n15187), .ZN(n6553) );
  NAND2_X1 U9394 ( .A1(n7429), .A2(n6426), .ZN(n6554) );
  INV_X1 U9395 ( .A(n7071), .ZN(n14535) );
  NOR2_X1 U9396 ( .A1(n14534), .A2(n14696), .ZN(n7071) );
  NAND2_X1 U9397 ( .A1(n8192), .A2(SI_26_), .ZN(n7427) );
  AND2_X1 U9398 ( .A1(n7434), .A2(n8257), .ZN(n6555) );
  AND2_X1 U9399 ( .A1(n11198), .A2(n11197), .ZN(n6556) );
  AND2_X1 U9400 ( .A1(n10411), .A2(n10410), .ZN(n6557) );
  AND2_X1 U9401 ( .A1(n7266), .A2(n7265), .ZN(n6558) );
  INV_X1 U9402 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11352) );
  INV_X1 U9403 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7123) );
  OR2_X1 U9404 ( .A1(n8992), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n6559) );
  AND2_X1 U9405 ( .A1(n8950), .A2(n12245), .ZN(n15072) );
  INV_X1 U9406 ( .A(n15072), .ZN(n15051) );
  INV_X1 U9407 ( .A(n11053), .ZN(n7067) );
  AND2_X2 U9408 ( .A1(n10031), .A2(n10566), .ZN(n14687) );
  AND2_X2 U9409 ( .A1(n10031), .A2(n9815), .ZN(n14679) );
  NAND2_X1 U9410 ( .A1(n9105), .A2(n9104), .ZN(n14652) );
  INV_X1 U9411 ( .A(n10951), .ZN(n7480) );
  OR2_X1 U9412 ( .A1(n12547), .A2(n15253), .ZN(n6560) );
  AND2_X1 U9413 ( .A1(n8250), .A2(n15242), .ZN(n6561) );
  AND2_X1 U9414 ( .A1(n14834), .A2(n10976), .ZN(n13531) );
  AND2_X1 U9415 ( .A1(n8824), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6562) );
  NAND2_X1 U9416 ( .A1(n8256), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n6563) );
  NOR2_X1 U9417 ( .A1(n8822), .A2(n7152), .ZN(n7151) );
  INV_X1 U9418 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7156) );
  INV_X1 U9419 ( .A(n9663), .ZN(n6633) );
  INV_X1 U9420 ( .A(n9659), .ZN(n6617) );
  INV_X1 U9421 ( .A(n8286), .ZN(n13174) );
  AND2_X1 U9422 ( .A1(n10497), .A2(n9737), .ZN(n9734) );
  INV_X1 U9423 ( .A(n9734), .ZN(n6915) );
  AND2_X1 U9424 ( .A1(n12594), .A2(n10404), .ZN(n12419) );
  NOR2_X1 U9425 ( .A1(n14873), .A2(n14872), .ZN(n6564) );
  AND2_X1 U9426 ( .A1(n6612), .A2(n6611), .ZN(n6565) );
  INV_X1 U9427 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n6978) );
  INV_X1 U9428 ( .A(n9698), .ZN(n7347) );
  INV_X1 U9429 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n6802) );
  XOR2_X1 U9430 ( .A(n7646), .B(n14445), .Z(n6566) );
  INV_X1 U9431 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n14311) );
  INV_X1 U9432 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6804) );
  INV_X1 U9433 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6898) );
  INV_X1 U9434 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n14309) );
  OAI21_X1 U9435 ( .B1(n13448), .B2(n6388), .A(n7294), .ZN(n7293) );
  OR2_X1 U9436 ( .A1(n14819), .A2(n10498), .ZN(n13434) );
  OAI22_X1 U9437 ( .A1(n12840), .A2(n12955), .B1(n15108), .B2(n8917), .ZN(
        n8918) );
  XNOR2_X1 U9438 ( .A(n12553), .B(n14450), .ZN(n14458) );
  OR2_X1 U9439 ( .A1(n14212), .A2(n14062), .ZN(n7383) );
  NAND2_X1 U9440 ( .A1(n6818), .A2(n14062), .ZN(n7373) );
  NAND2_X1 U9441 ( .A1(n12787), .A2(n12788), .ZN(n8867) );
  INV_X1 U9442 ( .A(n8852), .ZN(n12225) );
  NAND3_X1 U9443 ( .A1(n8533), .A2(n8353), .A3(n8354), .ZN(n8834) );
  OR2_X2 U9444 ( .A1(n13273), .A2(n13274), .ZN(n13276) );
  NAND2_X1 U9445 ( .A1(n13198), .A2(n6585), .ZN(n6584) );
  NAND2_X1 U9446 ( .A1(n13341), .A2(n13242), .ZN(n6587) );
  NAND3_X1 U9447 ( .A1(n11656), .A2(n7081), .A3(n11823), .ZN(n6588) );
  NAND2_X1 U9448 ( .A1(n13382), .A2(n13192), .ZN(n6589) );
  NAND2_X1 U9449 ( .A1(n13401), .A2(n13189), .ZN(n6590) );
  NAND2_X1 U9450 ( .A1(n10470), .A2(n10469), .ZN(n10472) );
  NAND2_X1 U9451 ( .A1(n6591), .A2(n10356), .ZN(n10470) );
  NAND2_X1 U9452 ( .A1(n10354), .A2(n10353), .ZN(n6591) );
  OR2_X2 U9453 ( .A1(n11640), .A2(n11663), .ZN(n11656) );
  XNOR2_X1 U9454 ( .A(n13110), .B(n11008), .ZN(n10052) );
  AOI21_X2 U9455 ( .B1(n13290), .B2(n13212), .A(n6593), .ZN(n13273) );
  OAI21_X2 U9456 ( .B1(n11198), .B2(n7076), .A(n7073), .ZN(n11363) );
  NAND2_X2 U9457 ( .A1(n11056), .A2(n11055), .ZN(n11198) );
  NAND2_X2 U9458 ( .A1(n7685), .A2(n8983), .ZN(n7995) );
  NAND2_X2 U9459 ( .A1(n13600), .A2(n9764), .ZN(n7685) );
  NAND3_X1 U9460 ( .A1(n6602), .A2(n6601), .A3(n7272), .ZN(n7271) );
  NOR2_X1 U9461 ( .A1(n14891), .A2(n11467), .ZN(n14912) );
  INV_X1 U9462 ( .A(n6604), .ZN(n12501) );
  NOR2_X1 U9463 ( .A1(n12473), .A2(n12472), .ZN(n12474) );
  INV_X1 U9464 ( .A(n6614), .ZN(n9883) );
  INV_X1 U9465 ( .A(n6618), .ZN(n6621) );
  NAND2_X1 U9466 ( .A1(n9500), .A2(n6627), .ZN(n9509) );
  OAI21_X1 U9467 ( .B1(n6630), .B2(n10584), .A(n10799), .ZN(n6629) );
  NAND2_X1 U9468 ( .A1(n13153), .A2(n13152), .ZN(n6634) );
  NAND3_X1 U9469 ( .A1(n14170), .A2(n14169), .A3(n6643), .ZN(n14262) );
  NAND2_X2 U9470 ( .A1(n12397), .A2(n12396), .ZN(n12628) );
  NAND2_X1 U9471 ( .A1(n7113), .A2(n7111), .ZN(n8632) );
  NAND2_X1 U9472 ( .A1(n8761), .A2(n8760), .ZN(n8764) );
  NAND3_X1 U9473 ( .A1(n6668), .A2(n14688), .A3(n6663), .ZN(n11792) );
  NAND3_X1 U9474 ( .A1(n11131), .A2(n7055), .A3(n14689), .ZN(n6663) );
  AOI21_X1 U9475 ( .B1(n12001), .B2(n6674), .A(n6673), .ZN(n6670) );
  INV_X1 U9476 ( .A(n12001), .ZN(n6671) );
  NAND2_X1 U9477 ( .A1(n6672), .A2(n12001), .ZN(n13021) );
  INV_X1 U9478 ( .A(n12007), .ZN(n6673) );
  NAND2_X1 U9479 ( .A1(n9534), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6680) );
  NAND3_X1 U9480 ( .A1(n7650), .A2(P2_DATAO_REG_1__SCAN_IN), .A3(n6897), .ZN(
        n6679) );
  INV_X1 U9481 ( .A(n7683), .ZN(n7680) );
  XNOR2_X1 U9482 ( .A(n10949), .B(n10950), .ZN(n10745) );
  NAND2_X1 U9483 ( .A1(n9599), .A2(n7910), .ZN(n6682) );
  INV_X1 U9484 ( .A(n10477), .ZN(n10544) );
  INV_X1 U9485 ( .A(n13107), .ZN(n6687) );
  NAND2_X1 U9486 ( .A1(n13235), .A2(n6702), .ZN(n6701) );
  NAND2_X1 U9487 ( .A1(n10781), .A2(n6704), .ZN(n10972) );
  XNOR2_X1 U9488 ( .A(n9995), .B(n9736), .ZN(n9980) );
  NAND2_X1 U9489 ( .A1(n13749), .A2(n13750), .ZN(n13748) );
  OR2_X2 U9490 ( .A1(n13749), .A2(n11975), .ZN(n6710) );
  INV_X1 U9491 ( .A(n13627), .ZN(n6713) );
  NAND2_X1 U9492 ( .A1(n6715), .A2(n6714), .ZN(n10261) );
  INV_X1 U9493 ( .A(n10142), .ZN(n6714) );
  INV_X1 U9494 ( .A(n6716), .ZN(n6715) );
  XNOR2_X1 U9495 ( .A(n10141), .B(n11983), .ZN(n6716) );
  NAND2_X1 U9496 ( .A1(n6716), .A2(n10142), .ZN(n10143) );
  OAI21_X1 U9497 ( .B1(n6721), .B2(n6719), .A(n6717), .ZN(n11685) );
  AND2_X1 U9498 ( .A1(n7248), .A2(n11677), .ZN(n6718) );
  NAND2_X1 U9499 ( .A1(n6720), .A2(n6721), .ZN(n11678) );
  NAND2_X1 U9500 ( .A1(n11289), .A2(n7248), .ZN(n6720) );
  OAI21_X1 U9501 ( .B1(n11289), .B2(n7250), .A(n7248), .ZN(n11401) );
  OAI21_X2 U9502 ( .B1(n13714), .B2(n6722), .A(n7225), .ZN(n13731) );
  AND2_X2 U9503 ( .A1(n6723), .A2(n6421), .ZN(n13714) );
  NAND2_X2 U9504 ( .A1(n10611), .A2(n10610), .ZN(n10858) );
  NAND2_X1 U9505 ( .A1(n10327), .A2(n6725), .ZN(n10611) );
  AND2_X1 U9506 ( .A1(n10334), .A2(n10326), .ZN(n6725) );
  XNOR2_X2 U9507 ( .A(n10858), .B(n10856), .ZN(n10855) );
  NAND2_X1 U9508 ( .A1(n6729), .A2(n6726), .ZN(n7716) );
  NAND2_X1 U9509 ( .A1(n6728), .A2(n6727), .ZN(n6726) );
  INV_X1 U9510 ( .A(n6732), .ZN(n6727) );
  INV_X1 U9511 ( .A(n6731), .ZN(n6728) );
  NAND2_X1 U9512 ( .A1(n6730), .A2(n7693), .ZN(n6729) );
  NAND2_X1 U9513 ( .A1(n6732), .A2(n6731), .ZN(n6730) );
  NAND2_X1 U9514 ( .A1(n7690), .A2(n7689), .ZN(n6732) );
  AOI21_X1 U9515 ( .B1(n8067), .B2(n8066), .A(n8065), .ZN(n6733) );
  OAI21_X1 U9516 ( .B1(n8067), .B2(n8066), .A(n6419), .ZN(n6734) );
  INV_X1 U9517 ( .A(n7859), .ZN(n6736) );
  NAND3_X1 U9518 ( .A1(n6736), .A2(n6504), .A3(n6740), .ZN(n6735) );
  NAND3_X1 U9519 ( .A1(n6743), .A2(n6742), .A3(n6741), .ZN(n7814) );
  NAND3_X1 U9520 ( .A1(n7585), .A2(n6974), .A3(n7587), .ZN(n6742) );
  NAND3_X1 U9521 ( .A1(n7585), .A2(n6507), .A3(n7587), .ZN(n6743) );
  INV_X1 U9522 ( .A(n8221), .ZN(n6748) );
  NAND2_X1 U9523 ( .A1(n7925), .A2(n6753), .ZN(n6752) );
  NAND3_X1 U9524 ( .A1(n8891), .A2(n8890), .A3(n6763), .ZN(n6762) );
  NAND3_X1 U9525 ( .A1(n6764), .A2(n7337), .A3(n11374), .ZN(n7334) );
  NAND2_X1 U9526 ( .A1(n6764), .A2(n10913), .ZN(n10915) );
  NAND2_X1 U9527 ( .A1(n6764), .A2(n7337), .ZN(n11077) );
  NAND2_X1 U9528 ( .A1(n6765), .A2(n12702), .ZN(n7328) );
  INV_X1 U9529 ( .A(n12172), .ZN(n6765) );
  NAND2_X1 U9530 ( .A1(n6766), .A2(n6389), .ZN(n12172) );
  OR2_X1 U9531 ( .A1(n12075), .A2(n12074), .ZN(n6766) );
  OAI22_X2 U9532 ( .A1(n11775), .A2(n11774), .B1(n14470), .B2(n11773), .ZN(
        n11777) );
  NAND2_X1 U9533 ( .A1(n6768), .A2(n6769), .ZN(n6774) );
  NAND2_X1 U9534 ( .A1(n8909), .A2(n6771), .ZN(n6768) );
  NAND3_X1 U9535 ( .A1(n6967), .A2(n12080), .A3(n12691), .ZN(n12097) );
  NAND3_X1 U9536 ( .A1(n6967), .A2(n12080), .A3(n6785), .ZN(n6784) );
  INV_X1 U9537 ( .A(n12159), .ZN(n6786) );
  NAND2_X1 U9538 ( .A1(n7550), .A2(n6790), .ZN(n6793) );
  NAND2_X1 U9539 ( .A1(n14427), .A2(n6798), .ZN(n6796) );
  INV_X1 U9540 ( .A(n14426), .ZN(n6797) );
  XNOR2_X1 U9541 ( .A(n14372), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n14375) );
  OAI21_X2 U9542 ( .B1(n9581), .B2(n9440), .A(n9120), .ZN(n11178) );
  NAND2_X1 U9543 ( .A1(n6404), .A2(n11554), .ZN(n6985) );
  NAND2_X1 U9544 ( .A1(n6829), .A2(n11316), .ZN(n6827) );
  AOI21_X1 U9545 ( .B1(n6829), .B2(n7382), .A(n6509), .ZN(n6828) );
  NAND2_X2 U9546 ( .A1(n13973), .A2(n13974), .ZN(n13972) );
  AOI21_X2 U9547 ( .B1(n14027), .B2(n13917), .A(n6497), .ZN(n14024) );
  NAND3_X1 U9548 ( .A1(n6838), .A2(n7408), .A3(n6837), .ZN(n7870) );
  NAND3_X1 U9549 ( .A1(n7410), .A2(n6839), .A3(n6841), .ZN(n6837) );
  NAND3_X1 U9550 ( .A1(n7797), .A2(n6839), .A3(n7410), .ZN(n6838) );
  NAND2_X1 U9551 ( .A1(n13891), .A2(n13890), .ZN(n14118) );
  NAND2_X1 U9552 ( .A1(n9353), .A2(n6850), .ZN(n6847) );
  OAI21_X1 U9553 ( .B1(n9353), .B2(n6851), .A(n6850), .ZN(n9368) );
  NAND2_X1 U9554 ( .A1(n6847), .A2(n6848), .ZN(n9367) );
  OAI211_X1 U9555 ( .C1(n9132), .C2(n6525), .A(n6853), .B(n7469), .ZN(n6856)
         );
  OAI21_X1 U9556 ( .B1(n6857), .B2(n6858), .A(n6859), .ZN(n9092) );
  NAND2_X1 U9557 ( .A1(n9092), .A2(n7463), .ZN(n6860) );
  NAND2_X1 U9558 ( .A1(n7461), .A2(n6860), .ZN(n9107) );
  NAND2_X1 U9559 ( .A1(n6983), .A2(n6861), .ZN(n6864) );
  AOI21_X1 U9560 ( .B1(n6416), .B2(n9197), .A(n6866), .ZN(n6865) );
  NAND3_X1 U9561 ( .A1(n7603), .A2(n9226), .A3(n7235), .ZN(n8972) );
  NAND4_X1 U9562 ( .A1(n7603), .A2(n9226), .A3(n7235), .A4(n8973), .ZN(n14278)
         );
  NAND2_X1 U9563 ( .A1(n6868), .A2(n6867), .ZN(n9288) );
  NAND3_X1 U9564 ( .A1(n9251), .A2(n6907), .A3(n9258), .ZN(n6867) );
  NAND2_X1 U9565 ( .A1(n9258), .A2(n6508), .ZN(n6869) );
  NAND3_X1 U9566 ( .A1(n9403), .A2(n6492), .A3(n6871), .ZN(n6870) );
  AOI21_X1 U9567 ( .B1(n6895), .B2(n6894), .A(n6893), .ZN(n7466) );
  OAI21_X1 U9568 ( .B1(n9288), .B2(n13894), .A(n9275), .ZN(n9290) );
  OAI21_X1 U9569 ( .B1(n9459), .B2(n7612), .A(n9033), .ZN(n9040) );
  NAND2_X1 U9570 ( .A1(n9166), .A2(n9167), .ZN(n9165) );
  OAI211_X1 U9571 ( .C1(n14164), .C2(n14257), .A(n14163), .B(n14162), .ZN(
        n14261) );
  NAND3_X1 U9572 ( .A1(n8921), .A2(n6880), .A3(n15051), .ZN(n8885) );
  NAND2_X1 U9573 ( .A1(n6882), .A2(n6881), .ZN(n6880) );
  INV_X1 U9574 ( .A(n8878), .ZN(n6882) );
  NAND2_X2 U9575 ( .A1(n12263), .A2(n12262), .ZN(n15063) );
  NAND2_X1 U9576 ( .A1(n15047), .A2(n15074), .ZN(n12262) );
  NAND2_X1 U9577 ( .A1(n7006), .A2(n7403), .ZN(n6886) );
  NAND2_X2 U9578 ( .A1(n14024), .A2(n14023), .ZN(n14201) );
  NAND2_X1 U9579 ( .A1(n10822), .A2(n10821), .ZN(n10823) );
  INV_X1 U9580 ( .A(n6940), .ZN(n10635) );
  NAND2_X1 U9581 ( .A1(n10307), .A2(n10306), .ZN(n10371) );
  OR2_X1 U9582 ( .A1(n8140), .A2(n7566), .ZN(n7563) );
  OAI21_X1 U9583 ( .B1(n8157), .B2(n8156), .A(n8155), .ZN(n8171) );
  OAI21_X1 U9584 ( .B1(n8049), .B2(n8048), .A(n8047), .ZN(n8067) );
  NAND2_X1 U9585 ( .A1(n10045), .A2(n10052), .ZN(n10185) );
  NAND2_X1 U9586 ( .A1(n9999), .A2(n9998), .ZN(n10044) );
  INV_X1 U9587 ( .A(n9304), .ZN(n6895) );
  OAI21_X1 U9588 ( .B1(n6890), .B2(n6889), .A(n7601), .ZN(n9503) );
  INV_X1 U9589 ( .A(n9475), .ZN(n6890) );
  INV_X1 U9590 ( .A(n13548), .ZN(n6891) );
  XNOR2_X1 U9591 ( .A(n13111), .B(n6896), .ZN(n9998) );
  OAI21_X1 U9592 ( .B1(n9327), .B2(n9328), .A(n6523), .ZN(n7457) );
  NAND2_X1 U9593 ( .A1(n6933), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n6897) );
  AOI21_X1 U9594 ( .B1(n8330), .B2(n8329), .A(n6920), .ZN(n6927) );
  NAND2_X1 U9595 ( .A1(n13289), .A2(n6955), .ZN(n8323) );
  AND2_X1 U9596 ( .A1(n8326), .A2(n13258), .ZN(n7435) );
  NAND2_X1 U9597 ( .A1(n10144), .A2(n10145), .ZN(n10262) );
  NAND2_X1 U9598 ( .A1(n13683), .A2(n13684), .ZN(n13694) );
  NAND2_X1 U9599 ( .A1(n13674), .A2(n13675), .ZN(n13673) );
  NAND2_X1 U9600 ( .A1(n9032), .A2(n9459), .ZN(n9033) );
  NAND2_X1 U9601 ( .A1(n9305), .A2(n7467), .ZN(n7465) );
  AOI21_X1 U9602 ( .B1(n9327), .B2(n9328), .A(n6899), .ZN(n7458) );
  AND2_X1 U9603 ( .A1(n9844), .A2(n9843), .ZN(n9850) );
  INV_X1 U9604 ( .A(n8194), .ZN(n7420) );
  OAI22_X1 U9605 ( .A1(n7466), .A2(n7465), .B1(n7468), .B2(n9315), .ZN(n9327)
         );
  AOI21_X1 U9606 ( .B1(n7599), .B2(n10076), .A(n9042), .ZN(n9043) );
  NAND2_X1 U9607 ( .A1(n8987), .A2(n7472), .ZN(n9008) );
  NAND3_X1 U9608 ( .A1(n8967), .A2(n8966), .A3(n6963), .ZN(n8970) );
  NAND2_X1 U9609 ( .A1(n13704), .A2(n13705), .ZN(n13703) );
  INV_X1 U9610 ( .A(n11685), .ZN(n11683) );
  NAND2_X1 U9611 ( .A1(n6935), .A2(n7452), .ZN(n9401) );
  NAND2_X1 U9612 ( .A1(n7445), .A2(n7448), .ZN(n9132) );
  NAND2_X1 U9613 ( .A1(n13637), .A2(n11961), .ZN(n13704) );
  NAND2_X1 U9614 ( .A1(n11168), .A2(n11167), .ZN(n11289) );
  NAND2_X1 U9615 ( .A1(n13731), .A2(n11956), .ZN(n13638) );
  NOR2_X1 U9616 ( .A1(n12121), .A2(n12071), .ZN(n12073) );
  NAND2_X1 U9617 ( .A1(n6918), .A2(n6917), .ZN(n6909) );
  XNOR2_X1 U9618 ( .A(n11477), .B(n11489), .ZN(n14867) );
  NAND2_X1 U9619 ( .A1(n14886), .A2(n14885), .ZN(n14884) );
  NAND2_X1 U9620 ( .A1(n11792), .A2(n11791), .ZN(n11797) );
  OAI21_X2 U9621 ( .B1(n7480), .B2(n10743), .A(n7479), .ZN(n11131) );
  NAND2_X1 U9622 ( .A1(n10124), .A2(n10122), .ZN(n10162) );
  NAND2_X1 U9623 ( .A1(n12054), .A2(n12053), .ZN(n12058) );
  NAND2_X1 U9624 ( .A1(n7477), .A2(n10123), .ZN(n10160) );
  OAI21_X1 U9625 ( .B1(n9737), .B2(n10497), .A(n6915), .ZN(n6914) );
  AOI21_X1 U9626 ( .B1(n8171), .B2(n6922), .A(n6921), .ZN(n6953) );
  NAND2_X1 U9627 ( .A1(n7721), .A2(n7720), .ZN(n7745) );
  AOI21_X1 U9628 ( .B1(n10040), .B2(n8242), .A(n7671), .ZN(n7669) );
  AOI21_X1 U9629 ( .B1(n7861), .B2(n7860), .A(n7858), .ZN(n7859) );
  NAND2_X1 U9630 ( .A1(n12263), .A2(n12259), .ZN(n10231) );
  XNOR2_X1 U9631 ( .A(n10229), .B(n15074), .ZN(n10228) );
  XNOR2_X1 U9632 ( .A(n11267), .B(n8936), .ZN(n7299) );
  INV_X1 U9633 ( .A(n11378), .ZN(n6918) );
  NAND2_X1 U9634 ( .A1(n7334), .A2(n7335), .ZN(n11378) );
  NAND2_X1 U9635 ( .A1(n9481), .A2(n6932), .ZN(n10078) );
  NAND2_X1 U9636 ( .A1(n7299), .A2(n11453), .ZN(n7297) );
  NAND2_X1 U9637 ( .A1(n13388), .A2(n13232), .ZN(n13235) );
  NAND2_X1 U9638 ( .A1(n12908), .A2(n6529), .ZN(P3_U3454) );
  NAND2_X1 U9639 ( .A1(n7516), .A2(n7515), .ZN(n11602) );
  NAND2_X1 U9640 ( .A1(n7512), .A2(n7511), .ZN(n12625) );
  NAND2_X1 U9641 ( .A1(n12907), .A2(n15108), .ZN(n7187) );
  OAI21_X2 U9642 ( .B1(n12757), .B2(n7521), .A(n7519), .ZN(n12728) );
  NAND2_X1 U9643 ( .A1(n13453), .A2(n6923), .ZN(n13547) );
  NAND2_X1 U9644 ( .A1(n8228), .A2(n8227), .ZN(n8249) );
  INV_X1 U9645 ( .A(n7419), .ZN(n8225) );
  AOI21_X1 U9646 ( .B1(n9043), .B2(n9044), .A(n10624), .ZN(n7438) );
  NAND2_X1 U9647 ( .A1(n7554), .A2(n7553), .ZN(n8330) );
  NAND2_X1 U9648 ( .A1(n13549), .A2(n6541), .ZN(P2_U3494) );
  NAND2_X1 U9649 ( .A1(n13458), .A2(n6536), .ZN(P2_U3526) );
  OAI21_X1 U9650 ( .B1(n6928), .B2(n8341), .A(n6927), .ZN(P2_U3328) );
  NAND2_X1 U9651 ( .A1(n8308), .A2(n11768), .ZN(n6928) );
  NAND2_X1 U9652 ( .A1(n6931), .A2(n6929), .ZN(n13458) );
  NAND2_X1 U9653 ( .A1(n14850), .A2(n6930), .ZN(n6929) );
  NAND2_X1 U9654 ( .A1(n11666), .A2(n11665), .ZN(n11825) );
  NAND2_X1 U9655 ( .A1(n7279), .A2(n7282), .ZN(n13272) );
  NAND2_X1 U9656 ( .A1(n10540), .A2(n10539), .ZN(n10781) );
  AOI21_X1 U9657 ( .B1(n14533), .B2(n14532), .A(n11357), .ZN(n11633) );
  NAND2_X1 U9658 ( .A1(n10805), .A2(n10810), .ZN(n10822) );
  XNOR2_X2 U9659 ( .A(n6940), .B(n10076), .ZN(n10026) );
  NAND2_X1 U9660 ( .A1(n13940), .A2(n6501), .ZN(n6945) );
  XNOR2_X1 U9661 ( .A(n8173), .B(SI_24_), .ZN(n8175) );
  NAND3_X1 U9662 ( .A1(n15256), .A2(n7646), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n6933) );
  NAND3_X1 U9663 ( .A1(n9373), .A2(n9372), .A3(n7450), .ZN(n6935) );
  AND2_X1 U9664 ( .A1(n8965), .A2(n8964), .ZN(n6963) );
  OAI21_X1 U9665 ( .B1(n14174), .B2(n14105), .A(n6987), .ZN(n6986) );
  NAND2_X1 U9666 ( .A1(n7401), .A2(n8068), .ZN(n7403) );
  NAND2_X1 U9667 ( .A1(n6945), .A2(n6944), .ZN(n13927) );
  AND2_X1 U9668 ( .A1(n10233), .A2(n10230), .ZN(n10253) );
  NAND2_X1 U9669 ( .A1(n10371), .A2(n7333), .ZN(n10646) );
  INV_X1 U9670 ( .A(n8355), .ZN(n8836) );
  NAND2_X1 U9671 ( .A1(n10823), .A2(n7377), .ZN(n7376) );
  NAND2_X1 U9672 ( .A1(n10625), .A2(n10624), .ZN(n10623) );
  NOR2_X1 U9674 ( .A1(n6943), .A2(n6942), .ZN(n6941) );
  NAND2_X1 U9675 ( .A1(n10803), .A2(n10802), .ZN(n10933) );
  NAND2_X1 U9676 ( .A1(n6985), .A2(n7392), .ZN(n14131) );
  NAND2_X1 U9677 ( .A1(n10646), .A2(n10645), .ZN(n10647) );
  NAND2_X2 U9678 ( .A1(n9734), .A2(n8286), .ZN(n8242) );
  NAND2_X1 U9679 ( .A1(n7660), .A2(n7659), .ZN(n11396) );
  INV_X1 U9680 ( .A(n8121), .ZN(n8122) );
  AOI22_X1 U9681 ( .A1(n8284), .A2(n10190), .B1(n13110), .B2(n7768), .ZN(n7742) );
  NAND2_X1 U9682 ( .A1(n7745), .A2(n7746), .ZN(n7744) );
  INV_X1 U9683 ( .A(n9108), .ZN(n7462) );
  NAND2_X1 U9684 ( .A1(n7752), .A2(n7751), .ZN(n7756) );
  NAND2_X1 U9685 ( .A1(n7773), .A2(n7772), .ZN(n7777) );
  AND2_X1 U9686 ( .A1(n8100), .A2(n8101), .ZN(n8103) );
  NAND2_X1 U9687 ( .A1(n7734), .A2(n7733), .ZN(n7752) );
  NAND2_X1 U9688 ( .A1(n7669), .A2(n7670), .ZN(n6946) );
  NAND2_X2 U9689 ( .A1(n9584), .A2(n8983), .ZN(n9440) );
  AOI21_X2 U9690 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n9663), .A(n9908), .ZN(
        n9636) );
  AOI21_X2 U9691 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n10176), .A(n10167), .ZN(
        n10171) );
  AOI21_X2 U9692 ( .B1(n9659), .B2(P2_REG2_REG_5__SCAN_IN), .A(n14747), .ZN(
        n9882) );
  AOI21_X2 U9693 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n11188), .A(n14766), .ZN(
        n13125) );
  NOR2_X2 U9694 ( .A1(n13127), .A2(n13126), .ZN(n13128) );
  NAND2_X2 U9695 ( .A1(n12077), .A2(n12076), .ZN(n12080) );
  INV_X1 U9696 ( .A(n11360), .ZN(n7076) );
  NAND3_X1 U9697 ( .A1(n7020), .A2(n13447), .A3(n13448), .ZN(n13546) );
  NAND2_X1 U9698 ( .A1(n8154), .A2(n8153), .ZN(n8155) );
  OR2_X1 U9699 ( .A1(n8277), .A2(n9526), .ZN(n6951) );
  OAI21_X1 U9700 ( .B1(n6953), .B2(n6952), .A(n7570), .ZN(n7567) );
  NOR2_X1 U9701 ( .A1(n8171), .A2(n6922), .ZN(n6952) );
  NAND2_X1 U9702 ( .A1(n8075), .A2(n7559), .ZN(n6964) );
  NAND2_X1 U9703 ( .A1(n11475), .A2(n6505), .ZN(n11477) );
  AOI21_X1 U9704 ( .B1(n7377), .B2(n7379), .A(n6510), .ZN(n7375) );
  NAND2_X1 U9705 ( .A1(n7842), .A2(n7841), .ZN(n7864) );
  NAND2_X1 U9706 ( .A1(n7376), .A2(n7375), .ZN(n14618) );
  AND2_X1 U9707 ( .A1(n7665), .A2(n7799), .ZN(n8023) );
  NOR2_X4 U9708 ( .A1(n7758), .A2(n7616), .ZN(n7799) );
  NAND2_X1 U9709 ( .A1(n7655), .A2(n7654), .ZN(n7659) );
  NAND2_X1 U9710 ( .A1(n13615), .A2(n7685), .ZN(n6965) );
  INV_X4 U9711 ( .A(n7866), .ZN(n9533) );
  NAND2_X1 U9712 ( .A1(n7420), .A2(n7429), .ZN(n7428) );
  OAI21_X1 U9713 ( .B1(n9503), .B2(n9504), .A(n9502), .ZN(n9517) );
  NAND2_X1 U9714 ( .A1(n6961), .A2(n9240), .ZN(n9241) );
  NAND2_X1 U9715 ( .A1(n9249), .A2(n6512), .ZN(n6961) );
  NOR2_X2 U9716 ( .A1(n8970), .A2(n9059), .ZN(n9226) );
  OAI21_X1 U9717 ( .B1(n9475), .B2(n6521), .A(n7600), .ZN(n9504) );
  NAND2_X1 U9718 ( .A1(n7952), .A2(n7951), .ZN(n7589) );
  AOI22_X1 U9719 ( .A1(n8125), .A2(n8124), .B1(n8122), .B2(n8123), .ZN(n8140)
         );
  NAND3_X1 U9720 ( .A1(n7750), .A2(n7586), .A3(n7749), .ZN(n7585) );
  NAND2_X1 U9721 ( .A1(n10872), .A2(n10871), .ZN(n11168) );
  NAND2_X1 U9722 ( .A1(n12079), .A2(n12078), .ZN(n6967) );
  AND2_X1 U9723 ( .A1(n10913), .A2(n7338), .ZN(n7337) );
  NAND2_X2 U9724 ( .A1(n12190), .A2(n12191), .ZN(n12189) );
  NAND2_X1 U9725 ( .A1(n8309), .A2(n7602), .ZN(n8308) );
  INV_X1 U9726 ( .A(n14375), .ZN(n7161) );
  NOR2_X1 U9727 ( .A1(n14780), .A2(n13137), .ZN(n14794) );
  XNOR2_X2 U9728 ( .A(n7686), .B(P2_IR_REG_1__SCAN_IN), .ZN(n9652) );
  NAND3_X1 U9729 ( .A1(n9171), .A2(n9170), .A3(n7454), .ZN(n6983) );
  NAND2_X1 U9730 ( .A1(n6984), .A2(n9292), .ZN(n9304) );
  NAND3_X1 U9731 ( .A1(n9290), .A2(n9289), .A3(n9478), .ZN(n6984) );
  OAI21_X2 U9732 ( .B1(n8158), .B2(n10991), .A(n8161), .ZN(n8173) );
  INV_X1 U9733 ( .A(n13249), .ZN(n7084) );
  NAND2_X1 U9734 ( .A1(n7270), .A2(n6994), .ZN(n6993) );
  NAND2_X1 U9735 ( .A1(n7270), .A2(n7269), .ZN(n7268) );
  NOR2_X1 U9736 ( .A1(n12452), .A2(n12805), .ZN(n12472) );
  OAI21_X1 U9737 ( .B1(n14930), .B2(n7000), .A(n6543), .ZN(n11470) );
  OAI21_X1 U9738 ( .B1(n12502), .B2(n7004), .A(n7003), .ZN(n12552) );
  NAND2_X1 U9739 ( .A1(n7403), .A2(n7402), .ZN(n7008) );
  INV_X1 U9740 ( .A(n7008), .ZN(n7007) );
  XNOR2_X1 U9741 ( .A(n7008), .B(SI_20_), .ZN(n8104) );
  OAI211_X1 U9742 ( .C1(n13448), .C2(n14846), .A(n7010), .B(n6506), .ZN(
        P2_U3496) );
  INV_X1 U9743 ( .A(n8175), .ZN(n7032) );
  OAI21_X1 U9744 ( .B1(n7035), .B2(SI_3_), .A(n7751), .ZN(n7034) );
  MUX2_X1 U9745 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n7866), .Z(n7035) );
  NAND3_X1 U9746 ( .A1(n10411), .A2(n13076), .A3(n10410), .ZN(n13075) );
  OAI211_X1 U9747 ( .C1(n6557), .C2(n13076), .A(n13075), .B(n14692), .ZN(
        n13083) );
  NAND2_X1 U9748 ( .A1(n7496), .A2(n6428), .ZN(n7039) );
  NAND2_X1 U9749 ( .A1(n7039), .A2(n7040), .ZN(n12029) );
  NAND2_X1 U9750 ( .A1(n12052), .A2(n7047), .ZN(n7046) );
  OAI211_X1 U9751 ( .C1(n12052), .C2(n7048), .A(n7046), .B(n13003), .ZN(
        P2_U3192) );
  NOR2_X2 U9752 ( .A1(n13305), .A2(n13292), .ZN(n13291) );
  NOR2_X2 U9753 ( .A1(n7063), .A2(n13255), .ZN(n13281) );
  NAND3_X1 U9754 ( .A1(n7066), .A2(n6435), .A3(n11159), .ZN(n11201) );
  AND2_X2 U9755 ( .A1(n10541), .A2(n7067), .ZN(n7066) );
  NOR2_X2 U9756 ( .A1(n13359), .A2(n13491), .ZN(n7070) );
  NAND4_X1 U9757 ( .A1(n7665), .A2(n7799), .A3(n7628), .A4(n7633), .ZN(n7072)
         );
  NOR2_X2 U9758 ( .A1(n7624), .A2(n7623), .ZN(n7665) );
  NOR2_X2 U9759 ( .A1(n10362), .A2(n11100), .ZN(n10481) );
  NAND2_X1 U9760 ( .A1(n7779), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7688) );
  NAND2_X1 U9761 ( .A1(n8262), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n7786) );
  NAND3_X1 U9762 ( .A1(n7653), .A2(n7583), .A3(n7799), .ZN(n7652) );
  NAND2_X1 U9763 ( .A1(n13326), .A2(n7086), .ZN(n7085) );
  NAND2_X1 U9764 ( .A1(n7085), .A2(n7083), .ZN(n13210) );
  NAND2_X1 U9765 ( .A1(n10975), .A2(n7096), .ZN(n7095) );
  OAI211_X1 U9766 ( .C1(n13273), .C2(n7100), .A(n7098), .B(n13264), .ZN(n13451) );
  NAND2_X1 U9767 ( .A1(n13273), .A2(n7099), .ZN(n7098) );
  NAND2_X1 U9768 ( .A1(n8594), .A2(n7114), .ZN(n7113) );
  NAND3_X1 U9769 ( .A1(n7119), .A2(n7121), .A3(n7117), .ZN(n8712) );
  NAND3_X1 U9770 ( .A1(n7119), .A2(n7118), .A3(n7117), .ZN(n8714) );
  NAND2_X1 U9771 ( .A1(n8512), .A2(n7139), .ZN(n7136) );
  NAND2_X1 U9772 ( .A1(n7136), .A2(n7137), .ZN(n8550) );
  NAND2_X1 U9773 ( .A1(n8808), .A2(n7151), .ZN(n7149) );
  INV_X1 U9774 ( .A(n7165), .ZN(n12660) );
  OR2_X1 U9775 ( .A1(n12705), .A2(n12714), .ZN(n7178) );
  NAND2_X1 U9776 ( .A1(n11115), .A2(n8858), .ZN(n7181) );
  NAND2_X1 U9777 ( .A1(n8867), .A2(n8866), .ZN(n12775) );
  NAND2_X1 U9778 ( .A1(n12775), .A2(n12776), .ZN(n7185) );
  NAND2_X1 U9779 ( .A1(n7187), .A2(n7186), .ZN(n12908) );
  OR2_X1 U9780 ( .A1(n15108), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n7186) );
  NOR2_X2 U9781 ( .A1(n12842), .A2(n6431), .ZN(n12907) );
  XNOR2_X1 U9782 ( .A(n12627), .B(n12628), .ZN(n7191) );
  NAND3_X1 U9783 ( .A1(n7198), .A2(n8852), .A3(n8851), .ZN(n10393) );
  OAI21_X2 U9784 ( .B1(n9584), .B2(n7347), .A(n7201), .ZN(n10076) );
  NAND2_X1 U9785 ( .A1(n6444), .A2(n10592), .ZN(n10944) );
  INV_X1 U9786 ( .A(n14652), .ZN(n7203) );
  AND2_X1 U9787 ( .A1(n13964), .A2(n7209), .ZN(n13930) );
  NAND2_X1 U9788 ( .A1(n13964), .A2(n7207), .ZN(n14152) );
  NAND3_X1 U9789 ( .A1(n7206), .A2(n7205), .A3(n7204), .ZN(n14149) );
  OR2_X1 U9790 ( .A1(n13964), .A2(n9458), .ZN(n7205) );
  NAND2_X1 U9791 ( .A1(n13964), .A2(n6520), .ZN(n7206) );
  INV_X1 U9792 ( .A(n11733), .ZN(n7214) );
  NAND3_X1 U9793 ( .A1(n7216), .A2(n7214), .A3(n7213), .ZN(n14109) );
  NOR2_X1 U9794 ( .A1(n7222), .A2(n7221), .ZN(n7220) );
  INV_X1 U9795 ( .A(n11907), .ZN(n7221) );
  INV_X1 U9796 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7224) );
  INV_X1 U9797 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n7223) );
  NAND2_X1 U9798 ( .A1(n10860), .A2(n6420), .ZN(n10872) );
  NAND2_X1 U9799 ( .A1(n7603), .A2(n9500), .ZN(n8980) );
  NAND2_X1 U9800 ( .A1(n10635), .A2(n7255), .ZN(n10077) );
  NAND2_X1 U9801 ( .A1(n10076), .A2(n10635), .ZN(n10084) );
  AND2_X1 U9802 ( .A1(n6940), .A2(n7255), .ZN(n7598) );
  OAI21_X1 U9803 ( .B1(n10635), .B2(n13793), .A(n7254), .ZN(P1_U3561) );
  NAND2_X1 U9804 ( .A1(n11463), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7256) );
  NAND4_X1 U9805 ( .A1(n7799), .A2(n7665), .A3(n7628), .A4(n7503), .ZN(n7663)
         );
  INV_X2 U9806 ( .A(n9736), .ZN(n10565) );
  NAND2_X1 U9807 ( .A1(n10186), .A2(n10352), .ZN(n10358) );
  NAND2_X1 U9808 ( .A1(n10185), .A2(n10184), .ZN(n10186) );
  NAND2_X1 U9809 ( .A1(n11635), .A2(n11634), .ZN(n11664) );
  OR2_X1 U9810 ( .A1(n6401), .A2(n10150), .ZN(n9843) );
  NAND4_X1 U9811 ( .A1(n9027), .A2(n9025), .A3(n9026), .A4(n9028), .ZN(n13789)
         );
  NAND2_X1 U9812 ( .A1(n10261), .A2(n10143), .ZN(n10147) );
  NOR2_X2 U9813 ( .A1(n13313), .A2(n13334), .ZN(n13315) );
  AND2_X2 U9814 ( .A1(n10486), .A2(n10481), .ZN(n10541) );
  NOR2_X2 U9815 ( .A1(n13424), .A2(n13229), .ZN(n13410) );
  NAND2_X1 U9817 ( .A1(n9850), .A2(n10136), .ZN(n10139) );
  NAND3_X1 U9818 ( .A1(n7297), .A2(n8889), .A3(n11579), .ZN(n8891) );
  NAND2_X1 U9819 ( .A1(n7301), .A2(n11380), .ZN(n7300) );
  AOI21_X1 U9820 ( .B1(n11454), .B2(n6502), .A(n7303), .ZN(n7302) );
  AND2_X1 U9821 ( .A1(n6503), .A2(n11587), .ZN(n7303) );
  OAI211_X1 U9822 ( .C1(n12189), .C2(n7310), .A(n7307), .B(n7305), .ZN(n12120)
         );
  OAI22_X1 U9823 ( .A1(n7306), .A2(n7309), .B1(n12112), .B2(n7311), .ZN(n7305)
         );
  NOR2_X1 U9824 ( .A1(n12092), .A2(n12112), .ZN(n7306) );
  NAND2_X1 U9825 ( .A1(n12189), .A2(n7308), .ZN(n7307) );
  NOR2_X1 U9826 ( .A1(n12112), .A2(n7309), .ZN(n7308) );
  NAND2_X1 U9827 ( .A1(n12092), .A2(n12112), .ZN(n7310) );
  NAND2_X1 U9828 ( .A1(n7314), .A2(n7316), .ZN(n12122) );
  OAI21_X1 U9829 ( .B1(n12179), .B2(n12178), .A(n7326), .ZN(n12104) );
  OR2_X1 U9830 ( .A1(n12068), .A2(n12727), .ZN(n7324) );
  NAND2_X1 U9831 ( .A1(n12067), .A2(n12713), .ZN(n7325) );
  NAND2_X1 U9832 ( .A1(n7328), .A2(n6389), .ZN(n12077) );
  AND2_X1 U9833 ( .A1(n7328), .A2(n7327), .ZN(n12177) );
  NAND2_X1 U9834 ( .A1(n12172), .A2(n12435), .ZN(n7327) );
  INV_X1 U9835 ( .A(n11777), .ZN(n7332) );
  NAND2_X1 U9836 ( .A1(n8355), .A2(n6524), .ZN(n8886) );
  NAND2_X1 U9837 ( .A1(n11273), .A2(n7343), .ZN(n7340) );
  NAND2_X1 U9838 ( .A1(n7340), .A2(n7341), .ZN(n11544) );
  INV_X2 U9839 ( .A(n9217), .ZN(n9277) );
  AOI21_X1 U9840 ( .B1(n14142), .B2(n6403), .A(n7352), .ZN(n7351) );
  INV_X1 U9841 ( .A(n14142), .ZN(n7355) );
  AND2_X1 U9842 ( .A1(n13922), .A2(n13923), .ZN(n7367) );
  NAND2_X1 U9843 ( .A1(n14057), .A2(n6513), .ZN(n7371) );
  INV_X1 U9844 ( .A(n7374), .ZN(n14060) );
  CLKBUF_X1 U9845 ( .A(n7389), .Z(n7385) );
  INV_X1 U9846 ( .A(n7385), .ZN(n13998) );
  NOR2_X1 U9847 ( .A1(n14197), .A2(n13919), .ZN(n7391) );
  AND2_X1 U9848 ( .A1(n7395), .A2(n7398), .ZN(n13955) );
  INV_X1 U9849 ( .A(n7395), .ZN(n13960) );
  INV_X1 U9850 ( .A(n13904), .ZN(n7397) );
  NAND2_X1 U9851 ( .A1(n13968), .A2(n13924), .ZN(n7398) );
  OAI21_X2 U9852 ( .B1(n9324), .B2(n7400), .A(n8144), .ZN(n8160) );
  XNOR2_X2 U9853 ( .A(n8143), .B(SI_22_), .ZN(n9324) );
  AOI21_X2 U9854 ( .B1(n8071), .B2(n7405), .A(n7404), .ZN(n7402) );
  NAND2_X1 U9855 ( .A1(n7430), .A2(n7431), .ZN(n8274) );
  NAND3_X1 U9856 ( .A1(n8228), .A2(n8227), .A3(n6555), .ZN(n7430) );
  NAND3_X1 U9857 ( .A1(n8228), .A2(n8227), .A3(n7434), .ZN(n7432) );
  NAND2_X1 U9858 ( .A1(n9067), .A2(n10086), .ZN(n7437) );
  OAI21_X2 U9859 ( .B1(n9445), .B2(n11354), .A(n7442), .ZN(n9023) );
  NAND3_X1 U9860 ( .A1(n9110), .A2(n7446), .A3(n9109), .ZN(n7445) );
  INV_X1 U9861 ( .A(n9314), .ZN(n7468) );
  NAND3_X1 U9862 ( .A1(n8986), .A2(n7476), .A3(n7475), .ZN(n7474) );
  INV_X1 U9863 ( .A(n10163), .ZN(n7477) );
  NAND2_X1 U9864 ( .A1(n10113), .A2(n10112), .ZN(n7478) );
  NAND2_X1 U9865 ( .A1(n10128), .A2(n10201), .ZN(n7489) );
  NAND2_X1 U9866 ( .A1(n7653), .A2(n7799), .ZN(n7661) );
  INV_X1 U9867 ( .A(n8306), .ZN(n8303) );
  NAND2_X1 U9868 ( .A1(n11566), .A2(n7517), .ZN(n7516) );
  OAI21_X1 U9869 ( .B1(n12791), .B2(n7526), .A(n7523), .ZN(n12768) );
  INV_X1 U9870 ( .A(n12791), .ZN(n7529) );
  NAND3_X1 U9871 ( .A1(n7533), .A2(n7535), .A3(n7532), .ZN(P3_U3488) );
  NAND2_X1 U9872 ( .A1(n12671), .A2(n7540), .ZN(n7537) );
  NAND3_X1 U9873 ( .A1(n8380), .A2(n8342), .A3(n8343), .ZN(n8443) );
  NAND2_X1 U9874 ( .A1(n7563), .A2(n7564), .ZN(n8154) );
  INV_X1 U9875 ( .A(n8207), .ZN(n7582) );
  NAND2_X1 U9876 ( .A1(n7771), .A2(n7584), .ZN(n7586) );
  INV_X1 U9877 ( .A(n7770), .ZN(n7584) );
  NAND2_X1 U9878 ( .A1(n6418), .A2(n7593), .ZN(n7925) );
  NAND2_X1 U9879 ( .A1(n7594), .A2(n7596), .ZN(n7861) );
  NAND3_X1 U9880 ( .A1(n7819), .A2(n7595), .A3(n7818), .ZN(n7594) );
  NAND2_X2 U9881 ( .A1(n14284), .A2(n14287), .ZN(n9036) );
  NAND2_X1 U9882 ( .A1(n8969), .A2(n8968), .ZN(n9059) );
  INV_X1 U9883 ( .A(n9057), .ZN(n8969) );
  INV_X1 U9884 ( .A(n9444), .ZN(n8999) );
  NAND2_X1 U9885 ( .A1(n8306), .A2(n8305), .ZN(n8332) );
  NAND2_X1 U9886 ( .A1(n10106), .A2(n10105), .ZN(n10113) );
  NAND2_X1 U9887 ( .A1(n7726), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7675) );
  INV_X1 U9888 ( .A(n12077), .ZN(n12079) );
  AOI21_X1 U9889 ( .B1(n12052), .B2(n12051), .A(n13073), .ZN(n12053) );
  AND2_X1 U9890 ( .A1(n12738), .A2(n12737), .ZN(n12882) );
  NAND4_X2 U9891 ( .A1(n9050), .A2(n9049), .A3(n9048), .A4(n9047), .ZN(n13788)
         );
  OAI222_X1 U9892 ( .A1(P3_U3151), .A2(n12974), .B1(n12973), .B2(n12972), .C1(
        n14410), .C2(n12971), .ZN(P3_U3267) );
  AND2_X1 U9893 ( .A1(n9459), .A2(n10635), .ZN(n7599) );
  AND3_X1 U9894 ( .A1(n9467), .A2(n9466), .A3(n9465), .ZN(n7600) );
  NAND2_X1 U9895 ( .A1(n9497), .A2(n9496), .ZN(n7601) );
  OR2_X1 U9896 ( .A1(n8302), .A2(n13174), .ZN(n7602) );
  INV_X1 U9897 ( .A(P3_U3897), .ZN(n12447) );
  INV_X1 U9898 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9000) );
  INV_X1 U9899 ( .A(n14080), .ZN(n13916) );
  AND2_X1 U9900 ( .A1(n8294), .A2(n8293), .ZN(n7604) );
  OR2_X1 U9901 ( .A1(n8128), .A2(SI_21_), .ZN(n7606) );
  AND2_X1 U9902 ( .A1(n8270), .A2(n8269), .ZN(n7607) );
  AND4_X1 U9903 ( .A1(n11553), .A2(n13908), .A3(n9459), .A4(n14562), .ZN(n7608) );
  OR2_X1 U9904 ( .A1(n8126), .A2(SI_20_), .ZN(n7609) );
  NOR2_X1 U9905 ( .A1(n14120), .A2(n14119), .ZN(n7610) );
  INV_X1 U9906 ( .A(n12756), .ZN(n8872) );
  INV_X1 U9907 ( .A(n14819), .ZN(n13438) );
  OR3_X1 U9908 ( .A1(n9826), .A2(n14078), .A3(n14290), .ZN(n7611) );
  AND2_X1 U9909 ( .A1(n9031), .A2(n9480), .ZN(n7612) );
  NOR2_X1 U9910 ( .A1(n9041), .A2(n10076), .ZN(n9042) );
  OAI21_X1 U9911 ( .B1(n6896), .B2(n8284), .A(n7713), .ZN(n7714) );
  AND2_X1 U9912 ( .A1(n13908), .A2(n11722), .ZN(n9240) );
  OAI21_X1 U9913 ( .B1(n11358), .B2(n8284), .A(n7923), .ZN(n7924) );
  OAI21_X1 U9914 ( .B1(n7768), .B2(n11364), .A(n7948), .ZN(n7951) );
  OR2_X1 U9915 ( .A1(n8043), .A2(n8042), .ZN(n8046) );
  AND2_X1 U9916 ( .A1(n8046), .A2(n8045), .ZN(n8047) );
  OAI22_X1 U9917 ( .A1(n13567), .A2(n8284), .B1(n7768), .B2(n13239), .ZN(n8120) );
  INV_X1 U9918 ( .A(n8152), .ZN(n8156) );
  INV_X1 U9919 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8351) );
  INV_X1 U9920 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8344) );
  INV_X1 U9921 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n7620) );
  NOR2_X1 U9922 ( .A1(n8683), .A2(n8352), .ZN(n8353) );
  INV_X1 U9923 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n7625) );
  INV_X1 U9924 ( .A(n8657), .ZN(n8656) );
  INV_X1 U9925 ( .A(n12276), .ZN(n8856) );
  INV_X1 U9926 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n11590) );
  INV_X1 U9927 ( .A(n12038), .ZN(n12036) );
  INV_X1 U9928 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7783) );
  INV_X1 U9929 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7848) );
  OAI21_X1 U9930 ( .B1(n11935), .B2(n10601), .A(n9846), .ZN(n9847) );
  INV_X1 U9931 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n9199) );
  INV_X1 U9932 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9723) );
  INV_X1 U9933 ( .A(n7905), .ZN(n7906) );
  NAND2_X1 U9934 ( .A1(n10647), .A2(n10648), .ZN(n10907) );
  NOR2_X1 U9935 ( .A1(n12629), .A2(n15046), .ZN(n8937) );
  INV_X1 U9936 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8553) );
  NAND2_X1 U9937 ( .A1(n9601), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8508) );
  INV_X1 U9938 ( .A(n10162), .ZN(n10123) );
  AND2_X1 U9939 ( .A1(n8261), .A2(n8237), .ZN(n12998) );
  OR2_X1 U9940 ( .A1(n8058), .A2(n8057), .ZN(n8079) );
  NOR2_X1 U9941 ( .A1(n9737), .A2(n11396), .ZN(n9768) );
  INV_X1 U9942 ( .A(n11686), .ZN(n11682) );
  INV_X1 U9943 ( .A(n9357), .ZN(n9358) );
  OR2_X1 U9944 ( .A1(n9232), .A2(n9231), .ZN(n9234) );
  INV_X1 U9945 ( .A(n11354), .ZN(n9461) );
  OR2_X1 U9946 ( .A1(n9293), .A2(n13717), .ZN(n9306) );
  INV_X1 U9947 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n15243) );
  NOR2_X1 U9948 ( .A1(n14351), .A2(n14350), .ZN(n14338) );
  INV_X1 U9949 ( .A(n12442), .ZN(n11612) );
  INV_X1 U9950 ( .A(n10693), .ZN(n10240) );
  NAND2_X1 U9951 ( .A1(n10211), .A2(n12959), .ZN(n10693) );
  INV_X1 U9952 ( .A(n11146), .ZN(n8932) );
  INV_X1 U9953 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n10650) );
  INV_X1 U9954 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n10917) );
  INV_X1 U9955 ( .A(n12435), .ZN(n12702) );
  INV_X1 U9956 ( .A(n12349), .ZN(n12765) );
  OR2_X1 U9957 ( .A1(n12602), .A2(n12601), .ZN(n12901) );
  INV_X1 U9958 ( .A(n10696), .ZN(n8846) );
  INV_X1 U9959 ( .A(n10644), .ZN(n11251) );
  INV_X1 U9960 ( .A(n14490), .ZN(n14494) );
  INV_X1 U9961 ( .A(n15067), .ZN(n15044) );
  AND2_X1 U9962 ( .A1(n8631), .A2(n8611), .ZN(n8612) );
  AND2_X1 U9963 ( .A1(n8558), .A2(n8548), .ZN(n8549) );
  AND2_X1 U9964 ( .A1(n8508), .A2(n8492), .ZN(n8493) );
  AND2_X1 U9965 ( .A1(n8440), .A2(n8428), .ZN(n8438) );
  INV_X1 U9966 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7938) );
  INV_X1 U9967 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n11261) );
  INV_X1 U9968 ( .A(n14694), .ZN(n13091) );
  NAND2_X1 U9969 ( .A1(n8030), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8058) );
  INV_X1 U9970 ( .A(n13067), .ZN(n14524) );
  OR3_X1 U9971 ( .A1(n13412), .A2(n13411), .A3(n10035), .ZN(n13518) );
  NAND2_X1 U9972 ( .A1(n9280), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9293) );
  INV_X1 U9973 ( .A(n13781), .ZN(n11407) );
  INV_X1 U9974 ( .A(n13777), .ZN(n13666) );
  INV_X1 U9975 ( .A(n13783), .ZN(n11344) );
  NAND2_X1 U9976 ( .A1(n10336), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13763) );
  NOR2_X1 U9977 ( .A1(n9306), .A2(n13656), .ZN(n9316) );
  NOR2_X1 U9978 ( .A1(n9234), .A2(n11428), .ZN(n9271) );
  INV_X1 U9979 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n10281) );
  INV_X1 U9980 ( .A(n13898), .ZN(n14070) );
  OR2_X1 U9981 ( .A1(n9853), .A2(n13796), .ZN(n14078) );
  INV_X1 U9982 ( .A(n14670), .ZN(n14653) );
  INV_X1 U9983 ( .A(n13887), .ZN(n11906) );
  OR2_X1 U9984 ( .A1(n10590), .A2(n14008), .ZN(n14105) );
  AND2_X1 U9985 ( .A1(n9808), .A2(n9834), .ZN(n10569) );
  INV_X1 U9986 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9009) );
  XNOR2_X1 U9987 ( .A(n7972), .B(SI_13_), .ZN(n7970) );
  XNOR2_X1 U9988 ( .A(n7930), .B(n9550), .ZN(n7928) );
  INV_X1 U9989 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n14358) );
  INV_X1 U9990 ( .A(n12181), .ZN(n12198) );
  AND2_X1 U9991 ( .A1(n8711), .A2(n8710), .ZN(n12727) );
  AND2_X1 U9992 ( .A1(n10707), .A2(n12559), .ZN(n14993) );
  INV_X1 U9993 ( .A(n15046), .ZN(n15066) );
  INV_X1 U9994 ( .A(n12820), .ZN(n12801) );
  INV_X1 U9995 ( .A(n10664), .ZN(n12822) );
  INV_X1 U9996 ( .A(n12829), .ZN(n14476) );
  AND2_X1 U9997 ( .A1(n8948), .A2(n8947), .ZN(n10661) );
  OR2_X1 U9998 ( .A1(n15106), .A2(n15099), .ZN(n14490) );
  NAND2_X1 U9999 ( .A1(n8841), .A2(n12258), .ZN(n15100) );
  XNOR2_X1 U10000 ( .A(n8833), .B(P3_IR_REG_22__SCAN_IN), .ZN(n12424) );
  OR2_X1 U10001 ( .A1(n8639), .A2(P3_IR_REG_16__SCAN_IN), .ZN(n8668) );
  AND2_X1 U10002 ( .A1(n9641), .A2(n9640), .ZN(n9646) );
  AND4_X1 U10003 ( .A1(n8266), .A2(n8265), .A3(n8264), .A4(n8263), .ZN(n12999)
         );
  AND4_X1 U10004 ( .A1(n8137), .A2(n8136), .A3(n8135), .A4(n8134), .ZN(n13243)
         );
  NAND4_X2 U10005 ( .A1(n7678), .A2(n7677), .A3(n7676), .A4(n7675), .ZN(n8312)
         );
  INV_X1 U10006 ( .A(n14770), .ZN(n14795) );
  INV_X1 U10007 ( .A(n14774), .ZN(n14802) );
  XNOR2_X1 U10008 ( .A(n13214), .B(n7295), .ZN(n13220) );
  INV_X1 U10009 ( .A(n13407), .ZN(n14808) );
  INV_X1 U10010 ( .A(n13413), .ZN(n14806) );
  NAND2_X1 U10011 ( .A1(n14827), .A2(n9762), .ZN(n13407) );
  INV_X1 U10012 ( .A(n14520), .ZN(n13538) );
  INV_X1 U10013 ( .A(n13541), .ZN(n11748) );
  OR2_X1 U10014 ( .A1(n9868), .A2(n9867), .ZN(n14520) );
  INV_X1 U10015 ( .A(n13531), .ZN(n14845) );
  AND2_X1 U10016 ( .A1(n9520), .A2(n9638), .ZN(n9770) );
  INV_X1 U10017 ( .A(n13763), .ZN(n13711) );
  AND2_X1 U10018 ( .A1(n10569), .A2(n9833), .ZN(n13753) );
  AND2_X1 U10019 ( .A1(n9299), .A2(n9298), .ZN(n14080) );
  AND2_X1 U10020 ( .A1(n9675), .A2(n9822), .ZN(n13873) );
  XOR2_X1 U10021 ( .A(n13941), .B(n13931), .Z(n13926) );
  INV_X1 U10022 ( .A(n13920), .ZN(n14023) );
  OR2_X1 U10023 ( .A1(n14662), .A2(n9505), .ZN(n9832) );
  AND2_X1 U10024 ( .A1(n10573), .A2(n10572), .ZN(n14146) );
  AOI21_X1 U10025 ( .B1(n9814), .B2(n9813), .A(n9812), .ZN(n10566) );
  INV_X1 U10026 ( .A(n14257), .ZN(n14677) );
  AND3_X1 U10027 ( .A1(n10569), .A2(n9832), .A3(n10567), .ZN(n10031) );
  NAND2_X1 U10028 ( .A1(n8908), .A2(n11579), .ZN(n10211) );
  AND2_X1 U10029 ( .A1(n10243), .A2(n10242), .ZN(n12187) );
  AND2_X1 U10030 ( .A1(n11153), .A2(n11152), .ZN(n12602) );
  NAND2_X1 U10031 ( .A1(n8790), .A2(n8789), .ZN(n12433) );
  INV_X1 U10032 ( .A(n12790), .ZN(n12437) );
  INV_X1 U10033 ( .A(n14457), .ZN(n15005) );
  NAND2_X1 U10034 ( .A1(n15036), .A2(n15015), .ZN(n12829) );
  NAND2_X1 U10035 ( .A1(n10661), .A2(n8955), .ZN(n15114) );
  INV_X1 U10036 ( .A(n12600), .ZN(n12903) );
  INV_X2 U10037 ( .A(n15110), .ZN(n15108) );
  OR2_X1 U10038 ( .A1(n15110), .A2(n15100), .ZN(n12955) );
  INV_X1 U10039 ( .A(n12253), .ZN(n12258) );
  INV_X1 U10040 ( .A(SI_13_), .ZN(n9596) );
  INV_X1 U10041 ( .A(n11494), .ZN(n14880) );
  NAND2_X1 U10042 ( .A1(n10129), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14701) );
  INV_X1 U10043 ( .A(n14697), .ZN(n13096) );
  NAND2_X1 U10044 ( .A1(n9760), .A2(n9759), .ZN(n13073) );
  INV_X1 U10045 ( .A(n13231), .ZN(n13190) );
  NAND2_X1 U10046 ( .A1(n14702), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14774) );
  INV_X1 U10047 ( .A(n14719), .ZN(n14805) );
  OR2_X1 U10048 ( .A1(n14819), .A2(n10500), .ZN(n14812) );
  NAND2_X1 U10049 ( .A1(n14852), .A2(n14830), .ZN(n13541) );
  AND2_X2 U10050 ( .A1(n9862), .A2(n9861), .ZN(n14852) );
  NAND2_X1 U10051 ( .A1(n10496), .A2(n10436), .ZN(n14846) );
  INV_X2 U10052 ( .A(n14846), .ZN(n14848) );
  OR2_X1 U10053 ( .A1(n14824), .A2(n14820), .ZN(n14821) );
  INV_X1 U10054 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10155) );
  NAND2_X1 U10055 ( .A1(n7611), .A2(n9515), .ZN(n9516) );
  OAI21_X1 U10056 ( .B1(n14050), .B2(n6399), .A(n9311), .ZN(n14062) );
  INV_X1 U10057 ( .A(n13873), .ZN(n14600) );
  INV_X1 U10058 ( .A(n14687), .ZN(n14685) );
  INV_X1 U10059 ( .A(n14679), .ZN(n14678) );
  AND2_X1 U10060 ( .A1(n9582), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9532) );
  INV_X1 U10061 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10385) );
  INV_X1 U10062 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9977) );
  NOR2_X2 U10063 ( .A1(n10211), .A2(n12957), .ZN(P3_U3897) );
  NOR2_X1 U10064 ( .A1(n9641), .A2(P2_U3088), .ZN(P2_U3947) );
  INV_X1 U10065 ( .A(n13793), .ZN(P1_U4016) );
  NOR2_X1 U10066 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), 
        .ZN(n7619) );
  NAND4_X1 U10067 ( .A1(n7619), .A2(n7618), .A3(n7617), .A4(n7826), .ZN(n7624)
         );
  NAND4_X1 U10068 ( .A1(n7622), .A2(n7621), .A3(n7620), .A4(n7844), .ZN(n7623)
         );
  NOR2_X1 U10069 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), 
        .ZN(n7632) );
  NOR2_X1 U10070 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), 
        .ZN(n7631) );
  NOR2_X1 U10071 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), 
        .ZN(n7630) );
  INV_X1 U10072 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n7629) );
  INV_X1 U10073 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7634) );
  NAND2_X1 U10074 ( .A1(n7651), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7635) );
  NOR2_X2 U10075 ( .A1(n7651), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n7638) );
  XNOR2_X2 U10076 ( .A(n7639), .B(P2_IR_REG_30__SCAN_IN), .ZN(n7640) );
  AND2_X2 U10077 ( .A1(n13593), .A2(n7640), .ZN(n7726) );
  NAND2_X1 U10078 ( .A1(n7726), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7645) );
  NAND2_X2 U10079 ( .A1(n7640), .A2(n7641), .ZN(n7723) );
  NAND2_X1 U10080 ( .A1(n7674), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7644) );
  NAND2_X1 U10081 ( .A1(n7725), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n7643) );
  AND2_X2 U10082 ( .A1(n7641), .A2(n11845), .ZN(n7722) );
  NAND2_X1 U10083 ( .A1(n9533), .A2(SI_0_), .ZN(n8373) );
  XNOR2_X1 U10084 ( .A(n8373), .B(n8370), .ZN(n13615) );
  NAND2_X1 U10085 ( .A1(n8313), .A2(n11088), .ZN(n7670) );
  INV_X1 U10086 ( .A(n7663), .ZN(n7655) );
  INV_X1 U10087 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n7654) );
  NAND2_X1 U10088 ( .A1(n7659), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7656) );
  NAND2_X1 U10089 ( .A1(n7663), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7658) );
  NAND2_X1 U10090 ( .A1(n7661), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7662) );
  MUX2_X1 U10091 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7662), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n7664) );
  NAND2_X1 U10092 ( .A1(n8023), .A2(n7666), .ZN(n8014) );
  INV_X1 U10093 ( .A(n8014), .ZN(n7667) );
  NAND2_X1 U10094 ( .A1(n7667), .A2(n7625), .ZN(n8053) );
  AND2_X1 U10095 ( .A1(n9864), .A2(n10497), .ZN(n7671) );
  NAND2_X1 U10096 ( .A1(n10040), .A2(n7671), .ZN(n7672) );
  NAND3_X1 U10097 ( .A1(n7672), .A2(n8313), .A3(n8242), .ZN(n7673) );
  NAND2_X1 U10098 ( .A1(n7722), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7678) );
  NAND2_X1 U10099 ( .A1(n7674), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n7677) );
  NAND2_X1 U10100 ( .A1(n7725), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7676) );
  NAND2_X1 U10101 ( .A1(n8312), .A2(n8242), .ZN(n7690) );
  INV_X1 U10102 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8371) );
  MUX2_X1 U10103 ( .A(n8371), .B(n8370), .S(n9534), .Z(n7679) );
  INV_X1 U10104 ( .A(SI_0_), .ZN(n9029) );
  NOR2_X1 U10105 ( .A1(n7679), .A2(n9029), .ZN(n7681) );
  NAND2_X1 U10106 ( .A1(n7680), .A2(n7681), .ZN(n7699) );
  INV_X1 U10107 ( .A(n7681), .ZN(n7682) );
  NAND2_X1 U10108 ( .A1(n7683), .A2(n7682), .ZN(n7684) );
  NAND2_X1 U10109 ( .A1(n7699), .A2(n7684), .ZN(n9526) );
  INV_X4 U10110 ( .A(n7685), .ZN(n8075) );
  NAND2_X1 U10111 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n7686) );
  NAND2_X1 U10112 ( .A1(n8075), .A2(n9652), .ZN(n7687) );
  NAND2_X1 U10113 ( .A1(n8242), .A2(n9736), .ZN(n7692) );
  NAND2_X1 U10114 ( .A1(n8312), .A2(n7768), .ZN(n7691) );
  NAND2_X1 U10115 ( .A1(n7692), .A2(n7691), .ZN(n7693) );
  NAND2_X1 U10116 ( .A1(n7722), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7697) );
  NAND2_X1 U10117 ( .A1(n7674), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7696) );
  NAND2_X1 U10118 ( .A1(n8262), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n7695) );
  NAND2_X1 U10119 ( .A1(n7726), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7694) );
  NAND2_X1 U10120 ( .A1(n13111), .A2(n7768), .ZN(n7712) );
  NAND2_X1 U10121 ( .A1(n7699), .A2(n7698), .ZN(n7704) );
  MUX2_X1 U10122 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n9534), .Z(n7700) );
  NAND2_X1 U10123 ( .A1(n7700), .A2(SI_2_), .ZN(n7731) );
  OAI21_X1 U10124 ( .B1(n7700), .B2(SI_2_), .A(n7731), .ZN(n7702) );
  NAND2_X1 U10125 ( .A1(n7701), .A2(n7702), .ZN(n7705) );
  INV_X1 U10126 ( .A(n7702), .ZN(n7703) );
  NAND2_X1 U10127 ( .A1(n7704), .A2(n7703), .ZN(n7732) );
  NAND2_X1 U10128 ( .A1(n7705), .A2(n7732), .ZN(n9544) );
  NOR2_X1 U10129 ( .A1(n9544), .A2(n8277), .ZN(n7710) );
  OAI22_X1 U10130 ( .A1(n7995), .A2(n9521), .B1(n7685), .B2(n6393), .ZN(n7709)
         );
  NAND2_X1 U10131 ( .A1(n8242), .A2(n10107), .ZN(n7711) );
  NAND2_X1 U10132 ( .A1(n7712), .A2(n7711), .ZN(n7717) );
  NAND2_X1 U10133 ( .A1(n7716), .A2(n7717), .ZN(n7715) );
  NAND2_X1 U10134 ( .A1(n13111), .A2(n8284), .ZN(n7713) );
  NAND2_X1 U10135 ( .A1(n7715), .A2(n7714), .ZN(n7721) );
  INV_X1 U10136 ( .A(n7716), .ZN(n7719) );
  INV_X1 U10137 ( .A(n7717), .ZN(n7718) );
  NAND2_X1 U10138 ( .A1(n7719), .A2(n7718), .ZN(n7720) );
  NAND2_X1 U10139 ( .A1(n8213), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7730) );
  INV_X1 U10140 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7724) );
  NAND2_X1 U10141 ( .A1(n8201), .A2(n7724), .ZN(n7729) );
  NAND2_X1 U10142 ( .A1(n8262), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n7728) );
  INV_X2 U10143 ( .A(n8246), .ZN(n8280) );
  NAND2_X1 U10144 ( .A1(n8280), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7727) );
  NAND2_X1 U10145 ( .A1(n13110), .A2(n8284), .ZN(n7741) );
  NAND2_X1 U10146 ( .A1(n7732), .A2(n7731), .ZN(n7734) );
  OR2_X1 U10147 ( .A1(n7734), .A2(n7733), .ZN(n7735) );
  AND2_X1 U10148 ( .A1(n7752), .A2(n7735), .ZN(n9522) );
  INV_X2 U10149 ( .A(n8277), .ZN(n7910) );
  NAND2_X1 U10150 ( .A1(n9522), .A2(n7910), .ZN(n7739) );
  INV_X2 U10151 ( .A(n7995), .ZN(n8256) );
  NAND2_X1 U10152 ( .A1(n7736), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7737) );
  XNOR2_X1 U10153 ( .A(n7737), .B(P2_IR_REG_3__SCAN_IN), .ZN(n13116) );
  AOI22_X1 U10154 ( .A1(n8256), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n8075), .B2(
        n13116), .ZN(n7738) );
  NAND2_X1 U10155 ( .A1(n10190), .A2(n8298), .ZN(n7740) );
  NAND2_X1 U10156 ( .A1(n7741), .A2(n7740), .ZN(n7746) );
  INV_X1 U10157 ( .A(n7742), .ZN(n7743) );
  NAND2_X1 U10158 ( .A1(n7744), .A2(n7743), .ZN(n7750) );
  INV_X1 U10159 ( .A(n7745), .ZN(n7748) );
  INV_X1 U10160 ( .A(n7746), .ZN(n7747) );
  NAND2_X1 U10161 ( .A1(n7748), .A2(n7747), .ZN(n7749) );
  MUX2_X1 U10162 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n9525), .Z(n7753) );
  NAND2_X1 U10163 ( .A1(n7753), .A2(SI_4_), .ZN(n7772) );
  OAI21_X1 U10164 ( .B1(n7753), .B2(SI_4_), .A(n7772), .ZN(n7754) );
  INV_X1 U10165 ( .A(n7754), .ZN(n7755) );
  NAND2_X1 U10166 ( .A1(n7756), .A2(n7755), .ZN(n7773) );
  OR2_X1 U10167 ( .A1(n7756), .A2(n7755), .ZN(n7757) );
  AND2_X1 U10168 ( .A1(n7773), .A2(n7757), .ZN(n9537) );
  NAND2_X1 U10169 ( .A1(n9537), .A2(n7910), .ZN(n7761) );
  NAND2_X1 U10170 ( .A1(n7758), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7759) );
  XNOR2_X1 U10171 ( .A(n7759), .B(P2_IR_REG_4__SCAN_IN), .ZN(n14739) );
  AOI22_X1 U10172 ( .A1(n8256), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n8075), .B2(
        n14739), .ZN(n7760) );
  NAND2_X1 U10173 ( .A1(n10499), .A2(n8284), .ZN(n7767) );
  NAND2_X1 U10174 ( .A1(n8280), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7765) );
  NAND2_X1 U10175 ( .A1(n8213), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7764) );
  NAND2_X1 U10176 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7784) );
  OAI21_X1 U10177 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n7784), .ZN(n10130) );
  INV_X1 U10178 ( .A(n10130), .ZN(n10502) );
  NAND2_X1 U10179 ( .A1(n8201), .A2(n10502), .ZN(n7763) );
  NAND2_X1 U10180 ( .A1(n8262), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n7762) );
  NAND2_X1 U10181 ( .A1(n13109), .A2(n7768), .ZN(n7766) );
  NAND2_X1 U10182 ( .A1(n7767), .A2(n7766), .ZN(n7771) );
  NAND2_X1 U10183 ( .A1(n10499), .A2(n7768), .ZN(n7769) );
  MUX2_X1 U10184 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n9533), .Z(n7774) );
  NAND2_X1 U10185 ( .A1(n7774), .A2(SI_5_), .ZN(n7793) );
  OAI21_X1 U10186 ( .B1(n7774), .B2(SI_5_), .A(n7793), .ZN(n7775) );
  INV_X1 U10187 ( .A(n7775), .ZN(n7776) );
  NAND2_X1 U10188 ( .A1(n7777), .A2(n7776), .ZN(n7794) );
  OR2_X1 U10189 ( .A1(n7777), .A2(n7776), .ZN(n7778) );
  NAND2_X1 U10190 ( .A1(n7794), .A2(n7778), .ZN(n9549) );
  OR2_X1 U10191 ( .A1(n9549), .A2(n8277), .ZN(n7782) );
  OAI21_X1 U10192 ( .B1(n7758), .B2(P2_IR_REG_4__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7780) );
  XNOR2_X1 U10193 ( .A(n7780), .B(P2_IR_REG_5__SCAN_IN), .ZN(n9659) );
  AOI22_X1 U10194 ( .A1(n8256), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8075), .B2(
        n9659), .ZN(n7781) );
  NAND2_X1 U10195 ( .A1(n7782), .A2(n7781), .ZN(n11100) );
  NAND2_X1 U10196 ( .A1(n11100), .A2(n8298), .ZN(n7791) );
  NAND2_X1 U10197 ( .A1(n8280), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7789) );
  NAND2_X1 U10198 ( .A1(n8213), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7788) );
  AND2_X1 U10199 ( .A1(n7784), .A2(n7783), .ZN(n7785) );
  NOR2_X1 U10200 ( .A1(n7803), .A2(n7785), .ZN(n11094) );
  NAND2_X1 U10201 ( .A1(n8201), .A2(n11094), .ZN(n7787) );
  NAND4_X1 U10202 ( .A1(n7789), .A2(n7788), .A3(n7787), .A4(n7786), .ZN(n13108) );
  NAND2_X1 U10203 ( .A1(n13108), .A2(n8284), .ZN(n7790) );
  AOI22_X1 U10204 ( .A1(n11100), .A2(n8284), .B1(n8298), .B2(n13108), .ZN(
        n7792) );
  MUX2_X1 U10205 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n9533), .Z(n7795) );
  OR2_X1 U10206 ( .A1(n7797), .A2(n7796), .ZN(n7798) );
  NAND2_X1 U10207 ( .A1(n7821), .A2(n7798), .ZN(n9575) );
  OR2_X1 U10208 ( .A1(n9575), .A2(n8277), .ZN(n7802) );
  OR2_X1 U10209 ( .A1(n7799), .A2(n7827), .ZN(n7800) );
  XNOR2_X1 U10210 ( .A(n7800), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9661) );
  AOI22_X1 U10211 ( .A1(n8256), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8075), .B2(
        n9661), .ZN(n7801) );
  NAND2_X1 U10212 ( .A1(n7802), .A2(n7801), .ZN(n13079) );
  NAND2_X1 U10213 ( .A1(n13079), .A2(n8284), .ZN(n7810) );
  NAND2_X1 U10214 ( .A1(n8280), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7808) );
  NAND2_X1 U10215 ( .A1(n8213), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7807) );
  NAND2_X1 U10216 ( .A1(n7803), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7831) );
  OR2_X1 U10217 ( .A1(n7803), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7804) );
  AND2_X1 U10218 ( .A1(n7831), .A2(n7804), .ZN(n13078) );
  NAND2_X1 U10219 ( .A1(n8201), .A2(n13078), .ZN(n7806) );
  NAND2_X1 U10220 ( .A1(n8262), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n7805) );
  NAND4_X1 U10221 ( .A1(n7808), .A2(n7807), .A3(n7806), .A4(n7805), .ZN(n13107) );
  NAND2_X1 U10222 ( .A1(n13107), .A2(n8298), .ZN(n7809) );
  NAND2_X1 U10223 ( .A1(n7810), .A2(n7809), .ZN(n7815) );
  NAND2_X1 U10224 ( .A1(n7814), .A2(n7815), .ZN(n7813) );
  NAND2_X1 U10225 ( .A1(n13079), .A2(n8298), .ZN(n7811) );
  OAI21_X1 U10226 ( .B1(n7768), .B2(n6687), .A(n7811), .ZN(n7812) );
  NAND2_X1 U10227 ( .A1(n7813), .A2(n7812), .ZN(n7819) );
  INV_X1 U10228 ( .A(n7814), .ZN(n7817) );
  INV_X1 U10229 ( .A(n7815), .ZN(n7816) );
  NAND2_X1 U10230 ( .A1(n7817), .A2(n7816), .ZN(n7818) );
  MUX2_X1 U10231 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n9533), .Z(n7822) );
  NAND2_X1 U10232 ( .A1(n7822), .A2(SI_7_), .ZN(n7841) );
  OAI21_X1 U10233 ( .B1(n7822), .B2(SI_7_), .A(n7841), .ZN(n7823) );
  INV_X1 U10234 ( .A(n7823), .ZN(n7824) );
  OR2_X1 U10235 ( .A1(n9581), .A2(n8277), .ZN(n7830) );
  AND2_X1 U10236 ( .A1(n7799), .A2(n7826), .ZN(n7845) );
  INV_X1 U10237 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n7827) );
  OR2_X1 U10238 ( .A1(n7845), .A2(n7827), .ZN(n7828) );
  XNOR2_X1 U10239 ( .A(n7828), .B(P2_IR_REG_7__SCAN_IN), .ZN(n9899) );
  AOI22_X1 U10240 ( .A1(n8256), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8075), .B2(
        n9899), .ZN(n7829) );
  NAND2_X1 U10241 ( .A1(n10785), .A2(n8298), .ZN(n7838) );
  NAND2_X1 U10242 ( .A1(n8280), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7836) );
  NAND2_X1 U10243 ( .A1(n8213), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7835) );
  NAND2_X1 U10244 ( .A1(n7831), .A2(n10427), .ZN(n7832) );
  AND2_X1 U10245 ( .A1(n7849), .A2(n7832), .ZN(n14809) );
  NAND2_X1 U10246 ( .A1(n8201), .A2(n14809), .ZN(n7834) );
  NAND4_X1 U10247 ( .A1(n7836), .A2(n7835), .A3(n7834), .A4(n7833), .ZN(n13106) );
  NAND2_X1 U10248 ( .A1(n13106), .A2(n8284), .ZN(n7837) );
  INV_X1 U10249 ( .A(n13106), .ZN(n10784) );
  NAND2_X1 U10250 ( .A1(n10785), .A2(n8284), .ZN(n7839) );
  OAI21_X1 U10251 ( .B1(n10784), .B2(n8284), .A(n7839), .ZN(n7840) );
  MUX2_X1 U10252 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n9533), .Z(n7843) );
  NAND2_X1 U10253 ( .A1(n7843), .A2(SI_8_), .ZN(n7865) );
  OAI21_X1 U10254 ( .B1(SI_8_), .B2(n7843), .A(n7865), .ZN(n7862) );
  XNOR2_X1 U10255 ( .A(n7864), .B(n7862), .ZN(n9599) );
  NAND2_X1 U10256 ( .A1(n7845), .A2(n7844), .ZN(n7872) );
  NAND2_X1 U10257 ( .A1(n7872), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7846) );
  XNOR2_X1 U10258 ( .A(n7846), .B(P2_IR_REG_8__SCAN_IN), .ZN(n9663) );
  AOI22_X1 U10259 ( .A1(n8256), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8075), .B2(
        n9663), .ZN(n7847) );
  NAND2_X1 U10260 ( .A1(n14831), .A2(n8284), .ZN(n7857) );
  NAND2_X1 U10261 ( .A1(n8213), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7855) );
  NAND2_X1 U10262 ( .A1(n7849), .A2(n7848), .ZN(n7850) );
  NAND2_X1 U10263 ( .A1(n7879), .A2(n7850), .ZN(n10980) );
  INV_X1 U10264 ( .A(n10980), .ZN(n7851) );
  NAND2_X1 U10265 ( .A1(n8201), .A2(n7851), .ZN(n7853) );
  NAND2_X1 U10266 ( .A1(n8280), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7852) );
  NAND4_X1 U10267 ( .A1(n7855), .A2(n7854), .A3(n7853), .A4(n7852), .ZN(n13105) );
  NAND2_X1 U10268 ( .A1(n13105), .A2(n8298), .ZN(n7856) );
  NAND2_X1 U10269 ( .A1(n7857), .A2(n7856), .ZN(n7860) );
  INV_X1 U10270 ( .A(n7862), .ZN(n7863) );
  MUX2_X1 U10271 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n9525), .Z(n7867) );
  OAI21_X1 U10272 ( .B1(n7867), .B2(SI_9_), .A(n7889), .ZN(n7868) );
  INV_X1 U10273 ( .A(n7868), .ZN(n7869) );
  NAND2_X1 U10274 ( .A1(n7870), .A2(n7869), .ZN(n7890) );
  NAND2_X1 U10275 ( .A1(n7890), .A2(n7871), .ZN(n9604) );
  OR2_X1 U10276 ( .A1(n9604), .A2(n8277), .ZN(n7877) );
  NAND2_X1 U10277 ( .A1(n7874), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7873) );
  MUX2_X1 U10278 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7873), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n7875) );
  NAND2_X1 U10279 ( .A1(n7875), .A2(n7911), .ZN(n9664) );
  INV_X1 U10280 ( .A(n9664), .ZN(n10013) );
  AOI22_X1 U10281 ( .A1(n8256), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n10013), 
        .B2(n8075), .ZN(n7876) );
  NAND2_X1 U10282 ( .A1(n11053), .A2(n8298), .ZN(n7886) );
  NAND2_X1 U10283 ( .A1(n8213), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7884) );
  NAND2_X1 U10284 ( .A1(n8280), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7883) );
  INV_X1 U10285 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7878) );
  AND2_X1 U10286 ( .A1(n7879), .A2(n7878), .ZN(n7880) );
  NOR2_X1 U10287 ( .A1(n7895), .A2(n7880), .ZN(n10958) );
  NAND2_X1 U10288 ( .A1(n8201), .A2(n10958), .ZN(n7882) );
  NAND4_X1 U10289 ( .A1(n7884), .A2(n7883), .A3(n7882), .A4(n7881), .ZN(n13104) );
  NAND2_X1 U10290 ( .A1(n13104), .A2(n8284), .ZN(n7885) );
  NAND2_X1 U10291 ( .A1(n7886), .A2(n7885), .ZN(n7888) );
  AOI22_X1 U10292 ( .A1(n11053), .A2(n8284), .B1(n8298), .B2(n13104), .ZN(
        n7887) );
  MUX2_X1 U10293 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n9533), .Z(n7905) );
  XNOR2_X1 U10294 ( .A(n7905), .B(SI_10_), .ZN(n7891) );
  XNOR2_X1 U10295 ( .A(n7909), .B(n7891), .ZN(n9618) );
  NAND2_X1 U10296 ( .A1(n9618), .A2(n7910), .ZN(n7894) );
  NAND2_X1 U10297 ( .A1(n7911), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7892) );
  XNOR2_X1 U10298 ( .A(n7892), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10176) );
  AOI22_X1 U10299 ( .A1(n8256), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n10176), 
        .B2(n8075), .ZN(n7893) );
  NAND2_X1 U10300 ( .A1(n11208), .A2(n8284), .ZN(n7902) );
  NAND2_X1 U10301 ( .A1(n8280), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7900) );
  NAND2_X1 U10302 ( .A1(n8213), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7899) );
  OR2_X1 U10303 ( .A1(n7895), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7896) );
  NAND2_X1 U10304 ( .A1(n7895), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7915) );
  AND2_X1 U10305 ( .A1(n7896), .A2(n7915), .ZN(n11143) );
  NAND2_X1 U10306 ( .A1(n8201), .A2(n11143), .ZN(n7898) );
  NAND4_X1 U10307 ( .A1(n7900), .A2(n7899), .A3(n7898), .A4(n7897), .ZN(n13103) );
  NAND2_X1 U10308 ( .A1(n13103), .A2(n8298), .ZN(n7901) );
  INV_X1 U10309 ( .A(n13103), .ZN(n11196) );
  NAND2_X1 U10310 ( .A1(n11208), .A2(n8298), .ZN(n7903) );
  OAI21_X1 U10311 ( .B1(n8298), .B2(n11196), .A(n7903), .ZN(n7904) );
  NOR2_X1 U10312 ( .A1(n7906), .A2(n14409), .ZN(n7908) );
  NAND2_X1 U10313 ( .A1(n7906), .A2(n14409), .ZN(n7907) );
  MUX2_X1 U10314 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n9525), .Z(n7930) );
  XNOR2_X1 U10315 ( .A(n7929), .B(n7928), .ZN(n9718) );
  NAND2_X1 U10316 ( .A1(n9718), .A2(n7910), .ZN(n7914) );
  OR2_X1 U10317 ( .A1(n7934), .A2(n7827), .ZN(n7912) );
  XNOR2_X1 U10318 ( .A(n7912), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10296) );
  AOI22_X1 U10319 ( .A1(n10296), .A2(n8075), .B1(n8256), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n7913) );
  NAND2_X1 U10320 ( .A1(n11359), .A2(n8298), .ZN(n7922) );
  NAND2_X1 U10321 ( .A1(n8280), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7920) );
  NAND2_X1 U10322 ( .A1(n8213), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7919) );
  NAND2_X1 U10323 ( .A1(n7915), .A2(n11261), .ZN(n7916) );
  AND2_X1 U10324 ( .A1(n7939), .A2(n7916), .ZN(n11264) );
  NAND2_X1 U10325 ( .A1(n7674), .A2(n11264), .ZN(n7918) );
  NAND4_X1 U10326 ( .A1(n7920), .A2(n7919), .A3(n7918), .A4(n7917), .ZN(n14523) );
  NAND2_X1 U10327 ( .A1(n14523), .A2(n8284), .ZN(n7921) );
  NAND2_X1 U10328 ( .A1(n7922), .A2(n7921), .ZN(n7926) );
  INV_X1 U10329 ( .A(n14523), .ZN(n11358) );
  NAND2_X1 U10330 ( .A1(n11359), .A2(n8284), .ZN(n7923) );
  INV_X1 U10331 ( .A(n7926), .ZN(n7927) );
  INV_X1 U10332 ( .A(n7930), .ZN(n7931) );
  NAND2_X1 U10333 ( .A1(n7931), .A2(n9550), .ZN(n7932) );
  MUX2_X1 U10334 ( .A(n9977), .B(n9892), .S(n9533), .Z(n7955) );
  NAND2_X1 U10335 ( .A1(n9891), .A2(n7910), .ZN(n7937) );
  INV_X1 U10336 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n7933) );
  OR2_X1 U10337 ( .A1(n7958), .A2(n7827), .ZN(n7935) );
  XNOR2_X1 U10338 ( .A(n7935), .B(P2_IR_REG_12__SCAN_IN), .ZN(n11186) );
  AOI22_X1 U10339 ( .A1(n11186), .A2(n8075), .B1(n8256), .B2(
        P1_DATAO_REG_12__SCAN_IN), .ZN(n7936) );
  NAND2_X1 U10340 ( .A1(n14696), .A2(n8284), .ZN(n7947) );
  NAND2_X1 U10341 ( .A1(n8213), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7945) );
  INV_X1 U10342 ( .A(n7962), .ZN(n7941) );
  NAND2_X1 U10343 ( .A1(n7939), .A2(n7938), .ZN(n7940) );
  NAND2_X1 U10344 ( .A1(n7941), .A2(n7940), .ZN(n14700) );
  INV_X1 U10345 ( .A(n14700), .ZN(n14530) );
  NAND2_X1 U10346 ( .A1(n8201), .A2(n14530), .ZN(n7944) );
  NAND2_X1 U10347 ( .A1(n8280), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7942) );
  NAND4_X1 U10348 ( .A1(n7945), .A2(n7944), .A3(n7943), .A4(n7942), .ZN(n13102) );
  NAND2_X1 U10349 ( .A1(n13102), .A2(n8298), .ZN(n7946) );
  NAND2_X1 U10350 ( .A1(n7947), .A2(n7946), .ZN(n7949) );
  INV_X1 U10351 ( .A(n13102), .ZN(n11364) );
  NAND2_X1 U10352 ( .A1(n14696), .A2(n8298), .ZN(n7948) );
  NAND2_X1 U10353 ( .A1(n7955), .A2(n9576), .ZN(n7956) );
  MUX2_X1 U10354 ( .A(n10060), .B(n10155), .S(n9525), .Z(n7972) );
  NAND2_X1 U10355 ( .A1(n10059), .A2(n7910), .ZN(n7961) );
  INV_X1 U10356 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n7957) );
  XNOR2_X1 U10357 ( .A(n7959), .B(P2_IR_REG_13__SCAN_IN), .ZN(n11188) );
  AOI22_X1 U10358 ( .A1(n11188), .A2(n8075), .B1(n8256), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n7960) );
  NAND2_X1 U10359 ( .A1(n8213), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7967) );
  NAND2_X1 U10360 ( .A1(n7962), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7980) );
  OR2_X1 U10361 ( .A1(n7962), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7963) );
  AND2_X1 U10362 ( .A1(n7980), .A2(n7963), .ZN(n11421) );
  NAND2_X1 U10363 ( .A1(n7674), .A2(n11421), .ZN(n7966) );
  NAND2_X1 U10364 ( .A1(n8262), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n7965) );
  NAND2_X1 U10365 ( .A1(n8280), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7964) );
  NAND4_X1 U10366 ( .A1(n7967), .A2(n7966), .A3(n7965), .A4(n7964), .ZN(n14525) );
  AOI22_X1 U10367 ( .A1(n11636), .A2(n7768), .B1(n8284), .B2(n14525), .ZN(
        n7968) );
  INV_X1 U10368 ( .A(n11636), .ZN(n14546) );
  INV_X1 U10369 ( .A(n14525), .ZN(n11641) );
  OAI22_X1 U10370 ( .A1(n14546), .A2(n8298), .B1(n11641), .B2(n8284), .ZN(
        n7969) );
  XNOR2_X1 U10371 ( .A(n8003), .B(SI_14_), .ZN(n7989) );
  MUX2_X1 U10372 ( .A(n10350), .B(n15254), .S(n9525), .Z(n8001) );
  XNOR2_X1 U10373 ( .A(n7989), .B(n8001), .ZN(n10344) );
  NAND2_X1 U10374 ( .A1(n10344), .A2(n7910), .ZN(n7978) );
  INV_X1 U10375 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n7973) );
  NAND2_X1 U10376 ( .A1(n7974), .A2(n7973), .ZN(n7992) );
  NAND2_X1 U10377 ( .A1(n7992), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7975) );
  XNOR2_X1 U10378 ( .A(n7975), .B(P2_IR_REG_14__SCAN_IN), .ZN(n13135) );
  NOR2_X1 U10379 ( .A1(n7995), .A2(n15254), .ZN(n7976) );
  AOI21_X1 U10380 ( .B1(n13135), .B2(n8075), .A(n7976), .ZN(n7977) );
  INV_X1 U10381 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7979) );
  NAND2_X1 U10382 ( .A1(n7980), .A2(n7979), .ZN(n7981) );
  NAND2_X1 U10383 ( .A1(n7997), .A2(n7981), .ZN(n14514) );
  INV_X1 U10384 ( .A(n14514), .ZN(n11645) );
  NAND2_X1 U10385 ( .A1(n11645), .A2(n8201), .ZN(n7985) );
  NAND2_X1 U10386 ( .A1(n8213), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7983) );
  NAND2_X1 U10387 ( .A1(n8280), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7982) );
  NAND4_X1 U10388 ( .A1(n7985), .A2(n7984), .A3(n7983), .A4(n7982), .ZN(n13101) );
  INV_X1 U10389 ( .A(n14511), .ZN(n11745) );
  INV_X1 U10390 ( .A(n13101), .ZN(n11654) );
  OAI22_X1 U10391 ( .A1(n11745), .A2(n8284), .B1(n7768), .B2(n11654), .ZN(
        n7986) );
  INV_X1 U10392 ( .A(n7987), .ZN(n8049) );
  INV_X1 U10393 ( .A(SI_14_), .ZN(n9616) );
  AND2_X1 U10394 ( .A1(n8003), .A2(n9616), .ZN(n7988) );
  AOI21_X1 U10395 ( .B1(n7989), .B2(n8001), .A(n7988), .ZN(n7991) );
  MUX2_X1 U10396 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n9525), .Z(n8005) );
  XNOR2_X1 U10397 ( .A(n8005), .B(SI_15_), .ZN(n7990) );
  OAI21_X1 U10398 ( .B1(n7992), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7994) );
  INV_X1 U10399 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n7993) );
  XNOR2_X1 U10400 ( .A(n7994), .B(n7993), .ZN(n14779) );
  OAI22_X1 U10401 ( .A1(n14779), .A2(n7685), .B1(n7995), .B2(n10387), .ZN(
        n7996) );
  INV_X1 U10402 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n11805) );
  AND2_X1 U10403 ( .A1(n7997), .A2(n11805), .ZN(n7998) );
  OR2_X1 U10404 ( .A1(n7998), .A2(n8028), .ZN(n11804) );
  AOI22_X1 U10405 ( .A1(n8213), .A2(P2_REG1_REG_15__SCAN_IN), .B1(n8280), .B2(
        P2_REG2_REG_15__SCAN_IN), .ZN(n8000) );
  NAND2_X1 U10406 ( .A1(n8262), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n7999) );
  OAI211_X1 U10407 ( .C1(n11804), .C2(n7723), .A(n8000), .B(n7999), .ZN(n13100) );
  AOI22_X1 U10408 ( .A1(n11809), .A2(n8284), .B1(n8298), .B2(n13100), .ZN(
        n8036) );
  INV_X1 U10409 ( .A(n13100), .ZN(n11826) );
  OAI22_X1 U10410 ( .A1(n14540), .A2(n8284), .B1(n7768), .B2(n11826), .ZN(
        n8037) );
  NAND2_X1 U10411 ( .A1(n8005), .A2(SI_15_), .ZN(n8007) );
  NAND2_X1 U10412 ( .A1(n8004), .A2(SI_14_), .ZN(n8002) );
  NOR2_X1 U10413 ( .A1(n8004), .A2(SI_14_), .ZN(n8008) );
  INV_X1 U10414 ( .A(SI_15_), .ZN(n9622) );
  INV_X1 U10415 ( .A(n8005), .ZN(n8006) );
  AOI22_X1 U10416 ( .A1(n8008), .A2(n8007), .B1(n9622), .B2(n8006), .ZN(n8009)
         );
  MUX2_X1 U10417 ( .A(n10346), .B(n10349), .S(n9533), .Z(n8011) );
  NAND2_X1 U10418 ( .A1(n8011), .A2(n9686), .ZN(n8012) );
  MUX2_X1 U10419 ( .A(n10385), .B(n10400), .S(n9533), .Z(n8050) );
  XNOR2_X1 U10420 ( .A(n8050), .B(SI_17_), .ZN(n8013) );
  XNOR2_X1 U10421 ( .A(n8052), .B(n8013), .ZN(n10384) );
  NAND2_X1 U10422 ( .A1(n10384), .A2(n7910), .ZN(n8017) );
  NAND2_X1 U10423 ( .A1(n8014), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8015) );
  XNOR2_X1 U10424 ( .A(n8015), .B(P2_IR_REG_17__SCAN_IN), .ZN(n13148) );
  AOI22_X1 U10425 ( .A1(n8256), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8075), 
        .B2(n13148), .ZN(n8016) );
  OR2_X1 U10426 ( .A1(n8030), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8018) );
  NAND2_X1 U10427 ( .A1(n8058), .A2(n8018), .ZN(n13034) );
  AOI22_X1 U10428 ( .A1(n8213), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n8280), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n8020) );
  OAI211_X1 U10429 ( .C1(n13034), .C2(n7723), .A(n8020), .B(n8019), .ZN(n13228) );
  AOI22_X1 U10430 ( .A1(n13229), .A2(n7768), .B1(n8284), .B2(n13228), .ZN(
        n8044) );
  INV_X1 U10431 ( .A(n13229), .ZN(n13580) );
  INV_X1 U10432 ( .A(n13228), .ZN(n13186) );
  OAI22_X1 U10433 ( .A1(n13580), .A2(n7768), .B1(n13186), .B2(n8284), .ZN(
        n8033) );
  XNOR2_X1 U10434 ( .A(n8022), .B(n8021), .ZN(n10345) );
  NAND2_X1 U10435 ( .A1(n10345), .A2(n7910), .ZN(n8027) );
  INV_X1 U10436 ( .A(n8023), .ZN(n8024) );
  NAND2_X1 U10437 ( .A1(n8024), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8025) );
  XNOR2_X1 U10438 ( .A(n8025), .B(P2_IR_REG_16__SCAN_IN), .ZN(n14801) );
  AOI22_X1 U10439 ( .A1(n8256), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8075), 
        .B2(n14801), .ZN(n8026) );
  NOR2_X1 U10440 ( .A1(n8028), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8029) );
  OR2_X1 U10441 ( .A1(n8030), .A2(n8029), .ZN(n13426) );
  AOI22_X1 U10442 ( .A1(n8213), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n8262), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n8032) );
  NAND2_X1 U10443 ( .A1(n8280), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8031) );
  OAI211_X1 U10444 ( .C1(n13426), .C2(n7723), .A(n8032), .B(n8031), .ZN(n13099) );
  AOI22_X1 U10445 ( .A1(n13422), .A2(n7768), .B1(n8284), .B2(n13099), .ZN(
        n8039) );
  INV_X1 U10446 ( .A(n13099), .ZN(n11830) );
  OAI22_X1 U10447 ( .A1(n13585), .A2(n7768), .B1(n11830), .B2(n8284), .ZN(
        n8038) );
  OAI22_X1 U10448 ( .A1(n8044), .A2(n8033), .B1(n8039), .B2(n8038), .ZN(n8042)
         );
  AOI21_X1 U10449 ( .B1(n8036), .B2(n8037), .A(n8042), .ZN(n8034) );
  INV_X1 U10450 ( .A(n8036), .ZN(n8041) );
  INV_X1 U10451 ( .A(n8037), .ZN(n8040) );
  AOI22_X1 U10452 ( .A1(n8041), .A2(n8040), .B1(n8039), .B2(n8038), .ZN(n8043)
         );
  OAI21_X1 U10453 ( .B1(n13228), .B2(n13229), .A(n8044), .ZN(n8045) );
  MUX2_X1 U10454 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n9533), .Z(n8069) );
  XNOR2_X1 U10455 ( .A(n8068), .B(n8069), .ZN(n10760) );
  NAND2_X1 U10456 ( .A1(n10760), .A2(n7910), .ZN(n8056) );
  NAND2_X1 U10457 ( .A1(n8053), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8054) );
  XNOR2_X1 U10458 ( .A(n8054), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13152) );
  AOI22_X1 U10459 ( .A1(n8256), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8075), 
        .B2(n13152), .ZN(n8055) );
  INV_X1 U10460 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8057) );
  NAND2_X1 U10461 ( .A1(n8058), .A2(n8057), .ZN(n8059) );
  NAND2_X1 U10462 ( .A1(n8079), .A2(n8059), .ZN(n13408) );
  OR2_X1 U10463 ( .A1(n13408), .A2(n7723), .ZN(n8064) );
  INV_X1 U10464 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n13409) );
  NAND2_X1 U10465 ( .A1(n8262), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8061) );
  NAND2_X1 U10466 ( .A1(n8213), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8060) );
  OAI211_X1 U10467 ( .C1(n8246), .C2(n13409), .A(n8061), .B(n8060), .ZN(n8062)
         );
  INV_X1 U10468 ( .A(n8062), .ZN(n8063) );
  OAI22_X1 U10469 ( .A1(n13520), .A2(n7768), .B1(n13231), .B2(n8284), .ZN(
        n8066) );
  AOI22_X1 U10470 ( .A1(n13416), .A2(n7768), .B1(n8284), .B2(n13190), .ZN(
        n8065) );
  MUX2_X1 U10471 ( .A(n10993), .B(n10995), .S(n9525), .Z(n8072) );
  NAND2_X1 U10472 ( .A1(n8072), .A2(n10156), .ZN(n8087) );
  INV_X1 U10473 ( .A(n8072), .ZN(n8073) );
  NAND2_X1 U10474 ( .A1(n8073), .A2(SI_19_), .ZN(n8074) );
  NAND2_X1 U10475 ( .A1(n8087), .A2(n8074), .ZN(n8088) );
  XNOR2_X1 U10476 ( .A(n8089), .B(n8088), .ZN(n10992) );
  NAND2_X1 U10477 ( .A1(n10992), .A2(n7910), .ZN(n8077) );
  AOI22_X1 U10478 ( .A1(n8256), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8286), 
        .B2(n8075), .ZN(n8076) );
  INV_X1 U10479 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8078) );
  AND2_X1 U10480 ( .A1(n8079), .A2(n8078), .ZN(n8080) );
  NOR2_X1 U10481 ( .A1(n8080), .A2(n8092), .ZN(n13391) );
  INV_X1 U10482 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13168) );
  NAND2_X1 U10483 ( .A1(n8262), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8082) );
  NAND2_X1 U10484 ( .A1(n8280), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8081) );
  OAI211_X1 U10485 ( .C1(n8116), .C2(n13168), .A(n8082), .B(n8081), .ZN(n8083)
         );
  AOI21_X1 U10486 ( .B1(n13391), .B2(n8201), .A(n8083), .ZN(n13233) );
  OAI22_X1 U10487 ( .A1(n13575), .A2(n8284), .B1(n7768), .B2(n13233), .ZN(
        n8085) );
  INV_X1 U10488 ( .A(n8085), .ZN(n8084) );
  OAI22_X1 U10489 ( .A1(n13575), .A2(n7768), .B1(n13233), .B2(n8284), .ZN(
        n8086) );
  MUX2_X1 U10490 ( .A(n11352), .B(n7123), .S(n9525), .Z(n8127) );
  XNOR2_X1 U10491 ( .A(n8104), .B(n8127), .ZN(n11331) );
  NAND2_X1 U10492 ( .A1(n11331), .A2(n7910), .ZN(n8091) );
  NAND2_X1 U10493 ( .A1(n8256), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8090) );
  OR2_X1 U10494 ( .A1(n8092), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8093) );
  NAND2_X1 U10495 ( .A1(n8111), .A2(n8093), .ZN(n13375) );
  OR2_X1 U10496 ( .A1(n13375), .A2(n7723), .ZN(n8098) );
  INV_X1 U10497 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n13508) );
  NAND2_X1 U10498 ( .A1(n8280), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8095) );
  NAND2_X1 U10499 ( .A1(n8262), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8094) );
  OAI211_X1 U10500 ( .C1(n8116), .C2(n13508), .A(n8095), .B(n8094), .ZN(n8096)
         );
  INV_X1 U10501 ( .A(n8096), .ZN(n8097) );
  NAND2_X1 U10502 ( .A1(n8098), .A2(n8097), .ZN(n13237) );
  AOI22_X1 U10503 ( .A1(n13370), .A2(n8284), .B1(n8298), .B2(n13237), .ZN(
        n8099) );
  AOI22_X1 U10504 ( .A1(n13370), .A2(n7768), .B1(n8284), .B2(n13237), .ZN(
        n8102) );
  INV_X1 U10505 ( .A(n8099), .ZN(n8101) );
  INV_X1 U10506 ( .A(n8127), .ZN(n8126) );
  NAND2_X1 U10507 ( .A1(n8104), .A2(n8126), .ZN(n8106) );
  INV_X1 U10508 ( .A(SI_20_), .ZN(n10402) );
  NAND2_X1 U10509 ( .A1(n8106), .A2(n8105), .ZN(n8108) );
  MUX2_X1 U10510 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9533), .Z(n8128) );
  XNOR2_X1 U10511 ( .A(n8128), .B(SI_21_), .ZN(n8107) );
  NAND2_X1 U10512 ( .A1(n11395), .A2(n7910), .ZN(n8110) );
  NAND2_X1 U10513 ( .A1(n8256), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8109) );
  INV_X1 U10514 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13008) );
  NAND2_X1 U10515 ( .A1(n8111), .A2(n13008), .ZN(n8113) );
  INV_X1 U10516 ( .A(n8133), .ZN(n8112) );
  NAND2_X1 U10517 ( .A1(n8113), .A2(n8112), .ZN(n13360) );
  OR2_X1 U10518 ( .A1(n13360), .A2(n7723), .ZN(n8119) );
  INV_X1 U10519 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n15201) );
  NAND2_X1 U10520 ( .A1(n8280), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8115) );
  NAND2_X1 U10521 ( .A1(n8262), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8114) );
  OAI211_X1 U10522 ( .C1(n8116), .C2(n15201), .A(n8115), .B(n8114), .ZN(n8117)
         );
  INV_X1 U10523 ( .A(n8117), .ZN(n8118) );
  NAND2_X1 U10524 ( .A1(n8121), .A2(n8120), .ZN(n8125) );
  OAI22_X1 U10525 ( .A1(n13567), .A2(n7768), .B1(n13239), .B2(n8284), .ZN(
        n8124) );
  INV_X1 U10526 ( .A(n8120), .ZN(n8123) );
  NOR2_X1 U10527 ( .A1(n8127), .A2(n10402), .ZN(n8129) );
  AOI22_X1 U10528 ( .A1(n8129), .A2(n7606), .B1(n8128), .B2(SI_21_), .ZN(n8130) );
  MUX2_X1 U10529 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n9533), .Z(n8142) );
  XNOR2_X1 U10530 ( .A(n9324), .B(n8142), .ZN(n11541) );
  NAND2_X1 U10531 ( .A1(n11541), .A2(n7910), .ZN(n8132) );
  NAND2_X1 U10532 ( .A1(n8256), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8131) );
  NAND2_X1 U10533 ( .A1(n8280), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8137) );
  NAND2_X1 U10534 ( .A1(n8213), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8136) );
  NAND2_X1 U10535 ( .A1(n8133), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8147) );
  OAI21_X1 U10536 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(n8133), .A(n8147), .ZN(
        n13061) );
  INV_X1 U10537 ( .A(n13061), .ZN(n13346) );
  NAND2_X1 U10538 ( .A1(n8201), .A2(n13346), .ZN(n8135) );
  NAND2_X1 U10539 ( .A1(n8262), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8134) );
  OAI22_X1 U10540 ( .A1(n13348), .A2(n7768), .B1(n13243), .B2(n8284), .ZN(
        n8138) );
  INV_X1 U10541 ( .A(n8138), .ZN(n8139) );
  OAI22_X1 U10542 ( .A1(n13348), .A2(n8284), .B1(n7768), .B2(n13243), .ZN(
        n8141) );
  MUX2_X1 U10543 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n9525), .Z(n8159) );
  XNOR2_X1 U10544 ( .A(n8158), .B(SI_23_), .ZN(n11767) );
  NAND2_X1 U10545 ( .A1(n11767), .A2(n7910), .ZN(n8146) );
  NAND2_X1 U10546 ( .A1(n8256), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8145) );
  NAND2_X1 U10547 ( .A1(n8213), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8151) );
  NAND2_X1 U10548 ( .A1(n7726), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8150) );
  INV_X1 U10549 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n12980) );
  AOI21_X1 U10550 ( .B1(n12980), .B2(n8147), .A(n8164), .ZN(n13331) );
  NAND2_X1 U10551 ( .A1(n8201), .A2(n13331), .ZN(n8149) );
  NAND2_X1 U10552 ( .A1(n8262), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8148) );
  NAND4_X1 U10553 ( .A1(n8151), .A2(n8150), .A3(n8149), .A4(n8148), .ZN(n13245) );
  AOI22_X1 U10554 ( .A1(n13336), .A2(n7768), .B1(n8284), .B2(n13245), .ZN(
        n8153) );
  INV_X1 U10555 ( .A(n13245), .ZN(n13204) );
  OAI22_X1 U10556 ( .A1(n7069), .A2(n7768), .B1(n13204), .B2(n8284), .ZN(n8152) );
  NAND2_X1 U10557 ( .A1(n8160), .A2(n8159), .ZN(n8161) );
  MUX2_X1 U10558 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n9533), .Z(n8172) );
  XNOR2_X1 U10559 ( .A(n8175), .B(n8172), .ZN(n13609) );
  NAND2_X1 U10560 ( .A1(n13609), .A2(n7910), .ZN(n8163) );
  NAND2_X1 U10561 ( .A1(n8256), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8162) );
  NAND2_X1 U10562 ( .A1(n8213), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8168) );
  NAND2_X1 U10563 ( .A1(n8280), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8167) );
  NAND2_X1 U10564 ( .A1(n8164), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n8182) );
  OAI21_X1 U10565 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(n8164), .A(n8182), .ZN(
        n13045) );
  INV_X1 U10566 ( .A(n13045), .ZN(n13317) );
  NAND2_X1 U10567 ( .A1(n7674), .A2(n13317), .ZN(n8166) );
  NAND4_X1 U10568 ( .A1(n8168), .A2(n8167), .A3(n8166), .A4(n8165), .ZN(n13247) );
  INV_X1 U10569 ( .A(n13247), .ZN(n13206) );
  OAI22_X1 U10570 ( .A1(n13559), .A2(n8284), .B1(n7768), .B2(n13206), .ZN(
        n8169) );
  NAND2_X1 U10571 ( .A1(n8173), .A2(SI_24_), .ZN(n8174) );
  INV_X1 U10572 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n14295) );
  INV_X1 U10573 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13608) );
  MUX2_X1 U10574 ( .A(n14295), .B(n13608), .S(n9525), .Z(n8176) );
  INV_X1 U10575 ( .A(SI_25_), .ZN(n11452) );
  NAND2_X1 U10576 ( .A1(n8176), .A2(n11452), .ZN(n8192) );
  INV_X1 U10577 ( .A(n8176), .ZN(n8177) );
  NAND2_X1 U10578 ( .A1(n8177), .A2(SI_25_), .ZN(n8178) );
  NAND2_X1 U10579 ( .A1(n8192), .A2(n8178), .ZN(n8193) );
  XNOR2_X1 U10580 ( .A(n8194), .B(n8193), .ZN(n13606) );
  NAND2_X1 U10581 ( .A1(n13606), .A2(n7910), .ZN(n8180) );
  NAND2_X1 U10582 ( .A1(n8256), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8179) );
  NAND2_X1 U10583 ( .A1(n8213), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8188) );
  NAND2_X1 U10584 ( .A1(n8262), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8187) );
  INV_X1 U10585 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8181) );
  NAND2_X1 U10586 ( .A1(n8181), .A2(n8182), .ZN(n8184) );
  INV_X1 U10587 ( .A(n8182), .ZN(n8183) );
  NAND2_X1 U10588 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(n8183), .ZN(n8199) );
  AND2_X1 U10589 ( .A1(n8184), .A2(n8199), .ZN(n13302) );
  NAND2_X1 U10590 ( .A1(n8201), .A2(n13302), .ZN(n8186) );
  NAND2_X1 U10591 ( .A1(n7726), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8185) );
  OAI22_X1 U10592 ( .A1(n13555), .A2(n8284), .B1(n7768), .B2(n13250), .ZN(
        n8189) );
  OAI22_X1 U10593 ( .A1(n13555), .A2(n7768), .B1(n13250), .B2(n8284), .ZN(
        n8191) );
  INV_X1 U10594 ( .A(n8189), .ZN(n8190) );
  INV_X1 U10595 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14292) );
  INV_X1 U10596 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8809) );
  MUX2_X1 U10597 ( .A(n14292), .B(n8809), .S(n9525), .Z(n8208) );
  XNOR2_X1 U10598 ( .A(n8208), .B(SI_26_), .ZN(n8195) );
  NAND2_X1 U10599 ( .A1(n8256), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8196) );
  NAND2_X1 U10600 ( .A1(n7726), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8205) );
  NAND2_X1 U10601 ( .A1(n8213), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8204) );
  INV_X1 U10602 ( .A(n8199), .ZN(n8198) );
  NAND2_X1 U10603 ( .A1(n8198), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n8215) );
  INV_X1 U10604 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n13090) );
  NAND2_X1 U10605 ( .A1(n8199), .A2(n13090), .ZN(n8200) );
  AND2_X1 U10606 ( .A1(n8215), .A2(n8200), .ZN(n13293) );
  NAND2_X1 U10607 ( .A1(n8201), .A2(n13293), .ZN(n8203) );
  NAND4_X1 U10608 ( .A1(n8205), .A2(n8204), .A3(n8203), .A4(n8202), .ZN(n13252) );
  AOI22_X1 U10609 ( .A1(n13292), .A2(n8284), .B1(n8298), .B2(n13252), .ZN(
        n8207) );
  OAI22_X1 U10610 ( .A1(n13460), .A2(n8284), .B1(n7768), .B2(n13253), .ZN(
        n8206) );
  INV_X1 U10611 ( .A(SI_26_), .ZN(n11582) );
  INV_X1 U10612 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8824) );
  INV_X1 U10613 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13599) );
  MUX2_X1 U10614 ( .A(n8824), .B(n13599), .S(n9533), .Z(n8223) );
  XNOR2_X1 U10615 ( .A(n8223), .B(SI_27_), .ZN(n8210) );
  NAND2_X1 U10616 ( .A1(n13598), .A2(n7910), .ZN(n8212) );
  NAND2_X1 U10617 ( .A1(n8256), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8211) );
  NAND2_X1 U10618 ( .A1(n7726), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8220) );
  NAND2_X1 U10619 ( .A1(n8213), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8219) );
  INV_X1 U10620 ( .A(n8215), .ZN(n8214) );
  NAND2_X1 U10621 ( .A1(n8214), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8236) );
  INV_X1 U10622 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n12055) );
  NAND2_X1 U10623 ( .A1(n8215), .A2(n12055), .ZN(n8216) );
  NAND2_X1 U10624 ( .A1(n7674), .A2(n13282), .ZN(n8218) );
  NAND2_X1 U10625 ( .A1(n8262), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8217) );
  AOI22_X1 U10626 ( .A1(n13255), .A2(n8242), .B1(n8298), .B2(n13256), .ZN(
        n8221) );
  INV_X1 U10627 ( .A(SI_27_), .ZN(n11652) );
  INV_X1 U10628 ( .A(n8223), .ZN(n8224) );
  NAND2_X1 U10629 ( .A1(n8225), .A2(n8224), .ZN(n8228) );
  INV_X1 U10630 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n11869) );
  INV_X1 U10631 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n15244) );
  MUX2_X1 U10632 ( .A(n11869), .B(n15244), .S(n9533), .Z(n8229) );
  INV_X1 U10633 ( .A(SI_28_), .ZN(n12972) );
  NAND2_X1 U10634 ( .A1(n8229), .A2(n12972), .ZN(n8247) );
  INV_X1 U10635 ( .A(n8229), .ZN(n8230) );
  NAND2_X1 U10636 ( .A1(n8230), .A2(SI_28_), .ZN(n8231) );
  NAND2_X1 U10637 ( .A1(n8247), .A2(n8231), .ZN(n8248) );
  NAND2_X1 U10638 ( .A1(n13595), .A2(n7910), .ZN(n8233) );
  NAND2_X1 U10639 ( .A1(n8256), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8232) );
  NAND2_X1 U10640 ( .A1(n7726), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8241) );
  NAND2_X1 U10641 ( .A1(n7722), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8240) );
  INV_X1 U10642 ( .A(n8236), .ZN(n8234) );
  NAND2_X1 U10643 ( .A1(n8234), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8261) );
  INV_X1 U10644 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8235) );
  NAND2_X1 U10645 ( .A1(n8236), .A2(n8235), .ZN(n8237) );
  NAND2_X1 U10646 ( .A1(n8201), .A2(n12998), .ZN(n8239) );
  NAND2_X1 U10647 ( .A1(n8262), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8238) );
  AOI22_X1 U10648 ( .A1(n7062), .A2(n8298), .B1(n8242), .B2(n13217), .ZN(n8267) );
  OAI22_X1 U10649 ( .A1(n13265), .A2(n7768), .B1(n13257), .B2(n8242), .ZN(
        n8268) );
  INV_X1 U10650 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8245) );
  NAND2_X1 U10651 ( .A1(n7722), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8244) );
  OAI211_X1 U10652 ( .C1(n8246), .C2(n8245), .A(n8244), .B(n8243), .ZN(n13097)
         );
  INV_X1 U10653 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14285) );
  INV_X1 U10654 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13592) );
  MUX2_X1 U10655 ( .A(n14285), .B(n13592), .S(n9525), .Z(n8250) );
  XNOR2_X1 U10656 ( .A(n8250), .B(SI_29_), .ZN(n8257) );
  INV_X1 U10657 ( .A(SI_29_), .ZN(n15242) );
  MUX2_X1 U10658 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n9533), .Z(n8251) );
  NAND2_X1 U10659 ( .A1(n8251), .A2(SI_30_), .ZN(n8252) );
  OAI21_X1 U10660 ( .B1(SI_30_), .B2(n8251), .A(n8252), .ZN(n8273) );
  MUX2_X1 U10661 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9525), .Z(n8253) );
  XNOR2_X1 U10662 ( .A(n8253), .B(SI_31_), .ZN(n8254) );
  NAND2_X1 U10663 ( .A1(n13591), .A2(n7910), .ZN(n8260) );
  NAND2_X1 U10664 ( .A1(n8256), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8259) );
  NAND2_X1 U10665 ( .A1(n7726), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8266) );
  NAND2_X1 U10666 ( .A1(n7722), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8265) );
  INV_X1 U10667 ( .A(n8261), .ZN(n13223) );
  NAND2_X1 U10668 ( .A1(n8201), .A2(n13223), .ZN(n8264) );
  NAND2_X1 U10669 ( .A1(n8262), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8263) );
  OAI22_X1 U10670 ( .A1(n13225), .A2(n7768), .B1(n12999), .B2(n8284), .ZN(
        n8289) );
  AOI22_X1 U10671 ( .A1(n13446), .A2(n8298), .B1(n8284), .B2(n13098), .ZN(
        n8290) );
  NAND2_X1 U10672 ( .A1(n8289), .A2(n8290), .ZN(n8270) );
  NAND2_X1 U10673 ( .A1(n8268), .A2(n8267), .ZN(n8269) );
  INV_X1 U10674 ( .A(n13097), .ZN(n8296) );
  MUX2_X1 U10675 ( .A(n7768), .B(n13097), .S(n11868), .Z(n8272) );
  OAI21_X1 U10676 ( .B1(n8296), .B2(n8242), .A(n8272), .ZN(n8292) );
  NAND2_X1 U10677 ( .A1(n8274), .A2(n8273), .ZN(n8275) );
  NAND2_X1 U10678 ( .A1(n8256), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8278) );
  NAND2_X1 U10679 ( .A1(n7722), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8283) );
  NAND2_X1 U10680 ( .A1(n8280), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8282) );
  AND3_X1 U10681 ( .A1(n8283), .A2(n8282), .A3(n8281), .ZN(n8285) );
  OAI22_X1 U10682 ( .A1(n13545), .A2(n7768), .B1(n8285), .B2(n8284), .ZN(n8293) );
  INV_X1 U10683 ( .A(n13545), .ZN(n8324) );
  INV_X1 U10684 ( .A(n8285), .ZN(n13215) );
  NOR2_X1 U10685 ( .A1(n13174), .A2(n9737), .ZN(n9868) );
  AOI211_X1 U10686 ( .C1(n9868), .C2(n7505), .A(n11396), .B(n8337), .ZN(n8287)
         );
  OAI21_X1 U10687 ( .B1(n8296), .B2(n7768), .A(n8287), .ZN(n8288) );
  AOI22_X1 U10688 ( .A1(n8324), .A2(n8298), .B1(n13215), .B2(n8288), .ZN(n8294) );
  OAI22_X1 U10689 ( .A1(n8293), .A2(n8294), .B1(n8290), .B2(n8289), .ZN(n8291)
         );
  NAND2_X1 U10690 ( .A1(n8292), .A2(n8291), .ZN(n8295) );
  INV_X1 U10691 ( .A(n11868), .ZN(n8297) );
  NOR3_X1 U10692 ( .A1(n8297), .A2(n8296), .A3(n8242), .ZN(n8300) );
  NOR3_X1 U10693 ( .A1(n11868), .A2(n8298), .A3(n13097), .ZN(n8299) );
  INV_X1 U10694 ( .A(n8337), .ZN(n9769) );
  OAI211_X1 U10695 ( .C1(n8286), .C2(n11396), .A(n6915), .B(n9769), .ZN(n8301)
         );
  MUX2_X1 U10696 ( .A(n11396), .B(n9737), .S(n7505), .Z(n8302) );
  NAND2_X1 U10697 ( .A1(n8303), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8304) );
  MUX2_X1 U10698 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8304), .S(
        P2_IR_REG_23__SCAN_IN), .Z(n8307) );
  NAND2_X1 U10699 ( .A1(n8307), .A2(n8332), .ZN(n9638) );
  INV_X1 U10700 ( .A(n9638), .ZN(n9519) );
  AND2_X1 U10701 ( .A1(n9519), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11768) );
  NAND2_X1 U10702 ( .A1(n13265), .A2(n13217), .ZN(n13213) );
  OAI21_X1 U10703 ( .B1(n13265), .B2(n13217), .A(n13213), .ZN(n13183) );
  OR2_X1 U10704 ( .A1(n13292), .A2(n13253), .ZN(n13212) );
  NAND2_X1 U10705 ( .A1(n13292), .A2(n13253), .ZN(n13211) );
  XNOR2_X1 U10706 ( .A(n13491), .B(n13243), .ZN(n13351) );
  INV_X1 U10707 ( .A(n13567), .ZN(n8310) );
  XNOR2_X1 U10708 ( .A(n8310), .B(n13239), .ZN(n13355) );
  INV_X1 U10709 ( .A(n13237), .ZN(n13196) );
  XNOR2_X1 U10710 ( .A(n13370), .B(n13196), .ZN(n13368) );
  INV_X1 U10711 ( .A(n13575), .ZN(n8311) );
  INV_X1 U10712 ( .A(n13233), .ZN(n13193) );
  XNOR2_X1 U10713 ( .A(n8311), .B(n13193), .ZN(n13386) );
  XNOR2_X1 U10714 ( .A(n13229), .B(n13186), .ZN(n13226) );
  XNOR2_X1 U10715 ( .A(n13422), .B(n13099), .ZN(n13430) );
  INV_X1 U10716 ( .A(n13105), .ZN(n10790) );
  XNOR2_X1 U10717 ( .A(n14831), .B(n10790), .ZN(n10782) );
  XNOR2_X1 U10718 ( .A(n11208), .B(n11196), .ZN(n11206) );
  XNOR2_X1 U10719 ( .A(n11053), .B(n13104), .ZN(n10792) );
  XNOR2_X1 U10720 ( .A(n11100), .B(n10473), .ZN(n10359) );
  XNOR2_X1 U10721 ( .A(n10355), .B(n10499), .ZN(n10352) );
  INV_X1 U10722 ( .A(n8313), .ZN(n9738) );
  NAND2_X1 U10723 ( .A1(n8313), .A2(n10040), .ZN(n9979) );
  OAI21_X1 U10724 ( .B1(n8313), .B2(n10040), .A(n9979), .ZN(n11092) );
  NAND4_X1 U10725 ( .A1(n10047), .A2(n9982), .A3(n9863), .A4(n11092), .ZN(
        n8314) );
  NOR4_X1 U10726 ( .A1(n10359), .A2(n10352), .A3(n10052), .A4(n8314), .ZN(
        n8315) );
  XNOR2_X1 U10727 ( .A(n10785), .B(n13106), .ZN(n10548) );
  NAND4_X1 U10728 ( .A1(n10792), .A2(n8315), .A3(n10548), .A4(n10544), .ZN(
        n8317) );
  NAND2_X1 U10729 ( .A1(n14696), .A2(n11364), .ZN(n8316) );
  NOR4_X1 U10730 ( .A1(n10782), .A2(n11206), .A3(n8317), .A4(n14532), .ZN(
        n8318) );
  XNOR2_X1 U10731 ( .A(n11636), .B(n14525), .ZN(n11362) );
  XNOR2_X1 U10732 ( .A(n11359), .B(n14523), .ZN(n11210) );
  NAND4_X1 U10733 ( .A1(n13430), .A2(n8318), .A3(n11362), .A4(n11210), .ZN(
        n8319) );
  XNOR2_X1 U10734 ( .A(n14511), .B(n11654), .ZN(n11663) );
  NOR3_X1 U10735 ( .A1(n13226), .A2(n8319), .A3(n11663), .ZN(n8320) );
  XNOR2_X1 U10736 ( .A(n13416), .B(n13190), .ZN(n13399) );
  NAND4_X1 U10737 ( .A1(n13386), .A2(n8320), .A3(n13399), .A4(n11824), .ZN(
        n8321) );
  NOR4_X1 U10738 ( .A1(n13351), .A2(n13355), .A3(n13368), .A4(n8321), .ZN(
        n8322) );
  XNOR2_X1 U10739 ( .A(n13336), .B(n13245), .ZN(n13332) );
  NOR4_X1 U10740 ( .A1(n13183), .A2(n13249), .A3(n13274), .A4(n8323), .ZN(
        n8326) );
  XNOR2_X1 U10741 ( .A(n8324), .B(n13215), .ZN(n8325) );
  INV_X1 U10742 ( .A(n11396), .ZN(n8328) );
  INV_X1 U10743 ( .A(n11768), .ZN(n8339) );
  NOR3_X1 U10744 ( .A1(n7605), .A2(n8328), .A3(n8339), .ZN(n8329) );
  INV_X1 U10745 ( .A(n9737), .ZN(n11540) );
  NAND2_X1 U10746 ( .A1(n8332), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8333) );
  MUX2_X1 U10747 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8333), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n8334) );
  NAND2_X1 U10748 ( .A1(n8335), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8336) );
  XNOR2_X1 U10749 ( .A(n8336), .B(P2_IR_REG_25__SCAN_IN), .ZN(n9743) );
  NAND3_X1 U10750 ( .A1(n13603), .A2(n13610), .A3(n9743), .ZN(n9520) );
  INV_X1 U10751 ( .A(n13600), .ZN(n9644) );
  INV_X1 U10752 ( .A(n9764), .ZN(n9642) );
  NAND4_X1 U10753 ( .A1(n14827), .A2(n8337), .A3(n9644), .A4(n14522), .ZN(
        n8338) );
  OAI211_X1 U10754 ( .C1(n11540), .C2(n8339), .A(n8338), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8340) );
  AND2_X2 U10755 ( .A1(n8445), .A2(n8346), .ZN(n8533) );
  NOR2_X1 U10756 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), 
        .ZN(n8350) );
  NAND4_X1 U10757 ( .A1(n8350), .A2(n8349), .A3(n8348), .A4(n8347), .ZN(n8683)
         );
  NAND3_X1 U10758 ( .A1(n8553), .A2(n8351), .A3(n8685), .ZN(n8352) );
  NOR2_X1 U10759 ( .A1(P3_IR_REG_26__SCAN_IN), .A2(P3_IR_REG_24__SCAN_IN), 
        .ZN(n8358) );
  NOR2_X1 U10760 ( .A1(P3_IR_REG_23__SCAN_IN), .A2(P3_IR_REG_22__SCAN_IN), 
        .ZN(n8357) );
  NAND4_X1 U10761 ( .A1(n8358), .A2(n8357), .A3(n8356), .A4(n7339), .ZN(n8359)
         );
  NAND2_X1 U10762 ( .A1(n8361), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8362) );
  NAND2_X1 U10763 ( .A1(n8402), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8369) );
  NAND2_X1 U10764 ( .A1(n8416), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8368) );
  NAND2_X1 U10765 ( .A1(n11146), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8367) );
  AND2_X4 U10766 ( .A1(n11856), .A2(n12968), .ZN(n11148) );
  NAND2_X1 U10767 ( .A1(n11148), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8366) );
  NAND2_X1 U10768 ( .A1(n8371), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8372) );
  AND2_X1 U10769 ( .A1(n8392), .A2(n8372), .ZN(n8374) );
  OAI21_X1 U10770 ( .B1(n9533), .B2(n8374), .A(n8373), .ZN(n12975) );
  XNOR2_X2 U10771 ( .A(n8377), .B(n8360), .ZN(n12974) );
  MUX2_X1 U10772 ( .A(P3_IR_REG_0__SCAN_IN), .B(n12975), .S(n10696), .Z(n10665) );
  INV_X1 U10773 ( .A(n10665), .ZN(n10622) );
  NAND2_X1 U10774 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n8379) );
  INV_X1 U10775 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n8378) );
  INV_X1 U10776 ( .A(n8380), .ZN(n8381) );
  NAND2_X4 U10777 ( .A1(n10696), .A2(n9533), .ZN(n12213) );
  INV_X1 U10778 ( .A(SI_1_), .ZN(n9573) );
  NAND2_X2 U10779 ( .A1(n6390), .A2(n8983), .ZN(n8637) );
  XNOR2_X1 U10780 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8394) );
  XNOR2_X1 U10781 ( .A(n8394), .B(n8392), .ZN(n9572) );
  NAND2_X1 U10782 ( .A1(n11148), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8385) );
  NAND2_X1 U10783 ( .A1(n8402), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8384) );
  NAND2_X1 U10784 ( .A1(n8416), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8383) );
  NAND2_X1 U10785 ( .A1(n11146), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n8386) );
  NAND2_X1 U10786 ( .A1(n10231), .A2(n12262), .ZN(n15041) );
  NAND2_X1 U10787 ( .A1(n11148), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8389) );
  NAND2_X1 U10788 ( .A1(n8416), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8388) );
  NAND2_X1 U10789 ( .A1(n8402), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8387) );
  NAND2_X1 U10790 ( .A1(n11146), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8390) );
  OR2_X1 U10791 ( .A1(n12213), .A2(SI_2_), .ZN(n8401) );
  INV_X1 U10792 ( .A(n8392), .ZN(n8393) );
  NAND2_X1 U10793 ( .A1(n8394), .A2(n8393), .ZN(n8396) );
  NAND2_X1 U10794 ( .A1(n15142), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8395) );
  NAND2_X1 U10795 ( .A1(n8396), .A2(n8395), .ZN(n8408) );
  NAND2_X1 U10796 ( .A1(n9521), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8409) );
  NAND2_X1 U10797 ( .A1(n9543), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8397) );
  XNOR2_X1 U10798 ( .A(n8408), .B(n8407), .ZN(n9569) );
  OR2_X1 U10799 ( .A1(n8637), .A2(n9569), .ZN(n8400) );
  OR2_X1 U10800 ( .A1(n10696), .A2(n11476), .ZN(n8399) );
  NAND2_X1 U10801 ( .A1(n15043), .A2(n12266), .ZN(n10389) );
  INV_X2 U10802 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n10755) );
  NAND2_X1 U10803 ( .A1(n8402), .A2(n10755), .ZN(n8406) );
  NAND2_X1 U10804 ( .A1(n8416), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8405) );
  NAND2_X1 U10805 ( .A1(n11146), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n8404) );
  OR2_X1 U10806 ( .A1(n12213), .A2(SI_3_), .ZN(n8415) );
  NAND2_X1 U10807 ( .A1(n8408), .A2(n8407), .ZN(n8410) );
  NAND2_X1 U10808 ( .A1(n9540), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8411) );
  XNOR2_X1 U10809 ( .A(n8425), .B(n8424), .ZN(n9553) );
  OR2_X1 U10810 ( .A1(n8637), .A2(n9553), .ZN(n8414) );
  NAND2_X1 U10811 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n6449), .ZN(n8412) );
  XNOR2_X1 U10812 ( .A(n8412), .B(P3_IR_REG_3__SCAN_IN), .ZN(n11489) );
  OR2_X1 U10813 ( .A1(n6390), .A2(n11489), .ZN(n8413) );
  NAND2_X1 U10814 ( .A1(n15045), .A2(n10756), .ZN(n12275) );
  INV_X1 U10815 ( .A(n10756), .ZN(n10776) );
  NAND2_X1 U10816 ( .A1(n10389), .A2(n12225), .ZN(n10388) );
  NAND2_X1 U10817 ( .A1(n10388), .A2(n12275), .ZN(n10528) );
  NAND2_X1 U10818 ( .A1(n11148), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8421) );
  NAND2_X1 U10819 ( .A1(n11147), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8420) );
  NAND2_X1 U10820 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8417) );
  NAND2_X1 U10821 ( .A1(n8432), .A2(n8417), .ZN(n15033) );
  NAND2_X1 U10822 ( .A1(n8402), .A2(n15033), .ZN(n8419) );
  NAND2_X1 U10823 ( .A1(n11146), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8418) );
  NAND4_X1 U10824 ( .A1(n8421), .A2(n8420), .A3(n8419), .A4(n8418), .ZN(n12446) );
  NAND2_X1 U10825 ( .A1(n8422), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8423) );
  XNOR2_X1 U10826 ( .A(n8423), .B(P3_IR_REG_4__SCAN_IN), .ZN(n11494) );
  NAND2_X1 U10827 ( .A1(n8425), .A2(n8424), .ZN(n8427) );
  NAND2_X1 U10828 ( .A1(n9545), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8428) );
  XNOR2_X1 U10829 ( .A(n8439), .B(n8438), .ZN(n9559) );
  OR2_X1 U10830 ( .A1(n8637), .A2(n9559), .ZN(n8430) );
  OR2_X1 U10831 ( .A1(n12213), .A2(SI_4_), .ZN(n8429) );
  OAI211_X1 U10832 ( .C1(n11494), .C2(n10696), .A(n8430), .B(n8429), .ZN(
        n12280) );
  XNOR2_X1 U10833 ( .A(n12280), .B(n12446), .ZN(n8854) );
  INV_X1 U10834 ( .A(n8854), .ZN(n12274) );
  NAND2_X1 U10835 ( .A1(n10528), .A2(n12274), .ZN(n10527) );
  INV_X1 U10836 ( .A(n12446), .ZN(n11039) );
  NAND2_X1 U10837 ( .A1(n11039), .A2(n15035), .ZN(n12281) );
  NAND2_X1 U10838 ( .A1(n10527), .A2(n12281), .ZN(n11034) );
  NAND2_X1 U10839 ( .A1(n11147), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8436) );
  INV_X1 U10840 ( .A(n8432), .ZN(n8431) );
  NAND2_X1 U10841 ( .A1(n8432), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n8433) );
  NAND2_X1 U10842 ( .A1(n8451), .A2(n8433), .ZN(n10643) );
  NAND2_X1 U10843 ( .A1(n6885), .A2(n10643), .ZN(n8435) );
  NAND2_X1 U10844 ( .A1(n11146), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8434) );
  OR2_X1 U10845 ( .A1(n12213), .A2(SI_5_), .ZN(n8450) );
  NAND2_X1 U10846 ( .A1(n8439), .A2(n8438), .ZN(n8441) );
  NAND2_X1 U10847 ( .A1(n9548), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8442) );
  XNOR2_X1 U10848 ( .A(n8459), .B(n8458), .ZN(n9556) );
  OR2_X1 U10849 ( .A1(n8637), .A2(n9556), .ZN(n8449) );
  NAND2_X1 U10850 ( .A1(n8443), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8444) );
  MUX2_X1 U10851 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8444), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n8447) );
  INV_X1 U10852 ( .A(n8445), .ZN(n8446) );
  OR2_X1 U10853 ( .A1(n10696), .A2(n11499), .ZN(n8448) );
  NAND2_X1 U10854 ( .A1(n11116), .A2(n10644), .ZN(n12288) );
  INV_X1 U10855 ( .A(n11116), .ZN(n12445) );
  NAND2_X1 U10856 ( .A1(n12445), .A2(n11251), .ZN(n12279) );
  NAND2_X1 U10857 ( .A1(n11034), .A2(n12276), .ZN(n11033) );
  NAND2_X1 U10858 ( .A1(n11033), .A2(n12288), .ZN(n11113) );
  NAND2_X1 U10859 ( .A1(n11148), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8456) );
  NAND2_X1 U10860 ( .A1(n11147), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8455) );
  OR2_X2 U10861 ( .A1(n8451), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8466) );
  NAND2_X1 U10862 ( .A1(n8451), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8452) );
  NAND2_X1 U10863 ( .A1(n8466), .A2(n8452), .ZN(n15026) );
  NAND2_X1 U10864 ( .A1(n8402), .A2(n15026), .ZN(n8454) );
  NAND2_X1 U10865 ( .A1(n11146), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8453) );
  OR2_X1 U10866 ( .A1(n8445), .A2(n6991), .ZN(n8457) );
  XNOR2_X1 U10867 ( .A(n8457), .B(P3_IR_REG_6__SCAN_IN), .ZN(n11504) );
  NAND2_X1 U10868 ( .A1(n8459), .A2(n8458), .ZN(n8461) );
  XNOR2_X1 U10869 ( .A(n9552), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n8462) );
  XNOR2_X1 U10870 ( .A(n8473), .B(n8462), .ZN(n9536) );
  OR2_X1 U10871 ( .A1(n8637), .A2(n9536), .ZN(n8464) );
  INV_X1 U10872 ( .A(SI_6_), .ZN(n9535) );
  OR2_X1 U10873 ( .A1(n12213), .A2(n9535), .ZN(n8463) );
  OAI211_X1 U10874 ( .C1(n6390), .C2(n14919), .A(n8464), .B(n8463), .ZN(n15025) );
  NAND2_X1 U10875 ( .A1(n11040), .A2(n15025), .ZN(n12290) );
  INV_X1 U10876 ( .A(n15025), .ZN(n11123) );
  NAND2_X1 U10877 ( .A1(n12444), .A2(n11123), .ZN(n12289) );
  NAND2_X1 U10878 ( .A1(n11113), .A2(n12226), .ZN(n11112) );
  NAND2_X1 U10879 ( .A1(n11112), .A2(n12290), .ZN(n11238) );
  NAND2_X1 U10880 ( .A1(n8416), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8471) );
  NAND2_X1 U10881 ( .A1(n11148), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8470) );
  NAND2_X1 U10882 ( .A1(n8466), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8467) );
  NAND2_X1 U10883 ( .A1(n8484), .A2(n8467), .ZN(n11387) );
  NAND2_X1 U10884 ( .A1(n8402), .A2(n11387), .ZN(n8469) );
  NAND2_X1 U10885 ( .A1(n11146), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8468) );
  NAND2_X1 U10886 ( .A1(n9574), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8472) );
  NAND2_X1 U10887 ( .A1(n9552), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8474) );
  NAND2_X1 U10888 ( .A1(n9578), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8475) );
  NAND2_X1 U10889 ( .A1(n8490), .A2(n8475), .ZN(n8476) );
  NAND2_X1 U10890 ( .A1(n8477), .A2(n8476), .ZN(n8478) );
  AND2_X1 U10891 ( .A1(n8478), .A2(n8491), .ZN(n9562) );
  OR2_X1 U10892 ( .A1(n12213), .A2(SI_7_), .ZN(n8482) );
  NAND2_X1 U10893 ( .A1(n8445), .A2(n8479), .ZN(n8496) );
  NAND2_X1 U10894 ( .A1(n8496), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8480) );
  XNOR2_X1 U10895 ( .A(n8480), .B(P3_IR_REG_7__SCAN_IN), .ZN(n11509) );
  OR2_X1 U10896 ( .A1(n10696), .A2(n11509), .ZN(n8481) );
  NAND2_X1 U10897 ( .A1(n11231), .A2(n10884), .ZN(n12294) );
  NAND2_X1 U10898 ( .A1(n12443), .A2(n11389), .ZN(n12295) );
  NAND2_X1 U10899 ( .A1(n11238), .A2(n7180), .ZN(n11237) );
  NAND2_X1 U10900 ( .A1(n11237), .A2(n12294), .ZN(n11566) );
  NAND2_X1 U10901 ( .A1(n11148), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8489) );
  NAND2_X1 U10902 ( .A1(n11147), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8488) );
  NAND2_X1 U10903 ( .A1(n8484), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8485) );
  NAND2_X1 U10904 ( .A1(n8502), .A2(n8485), .ZN(n15019) );
  NAND2_X1 U10905 ( .A1(n8402), .A2(n15019), .ZN(n8487) );
  NAND2_X1 U10906 ( .A1(n11146), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8486) );
  NAND4_X1 U10907 ( .A1(n8489), .A2(n8488), .A3(n8487), .A4(n8486), .ZN(n12442) );
  NAND2_X1 U10908 ( .A1(n9600), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8492) );
  OR2_X1 U10909 ( .A1(n8494), .A2(n8493), .ZN(n8495) );
  NAND2_X1 U10910 ( .A1(n8509), .A2(n8495), .ZN(n9568) );
  OR2_X1 U10911 ( .A1(n8637), .A2(n9568), .ZN(n8500) );
  INV_X1 U10912 ( .A(SI_8_), .ZN(n9567) );
  OR2_X1 U10913 ( .A1(n12213), .A2(n9567), .ZN(n8499) );
  NAND2_X1 U10914 ( .A1(n8514), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8497) );
  XNOR2_X1 U10915 ( .A(n8497), .B(P3_IR_REG_8__SCAN_IN), .ZN(n11514) );
  OR2_X1 U10916 ( .A1(n6390), .A2(n14957), .ZN(n8498) );
  XNOR2_X1 U10917 ( .A(n12442), .B(n12299), .ZN(n11570) );
  INV_X1 U10918 ( .A(n12299), .ZN(n15018) );
  NAND2_X1 U10919 ( .A1(n11612), .A2(n15018), .ZN(n12300) );
  NAND2_X1 U10920 ( .A1(n11147), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8506) );
  INV_X1 U10921 ( .A(n8502), .ZN(n8501) );
  NAND2_X1 U10922 ( .A1(n8502), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n8503) );
  NAND2_X1 U10923 ( .A1(n8522), .A2(n8503), .ZN(n11616) );
  NAND2_X1 U10924 ( .A1(n8402), .A2(n11616), .ZN(n8505) );
  NAND2_X1 U10925 ( .A1(n11146), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8504) );
  NAND4_X1 U10926 ( .A1(n8507), .A2(n8506), .A3(n8505), .A4(n8504), .ZN(n12441) );
  NAND2_X1 U10927 ( .A1(n9598), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8510) );
  OR2_X1 U10928 ( .A1(n8512), .A2(n8511), .ZN(n8513) );
  NAND2_X1 U10929 ( .A1(n8529), .A2(n8513), .ZN(n9566) );
  NAND2_X1 U10930 ( .A1(n12212), .A2(n9566), .ZN(n8521) );
  OR2_X1 U10931 ( .A1(n12213), .A2(SI_9_), .ZN(n8520) );
  NOR2_X1 U10932 ( .A1(n8514), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n8517) );
  OR2_X1 U10933 ( .A1(n8517), .A2(n6991), .ZN(n8515) );
  MUX2_X1 U10934 ( .A(n8515), .B(P3_IR_REG_31__SCAN_IN), .S(n8516), .Z(n8518)
         );
  NAND2_X1 U10935 ( .A1(n8517), .A2(n8516), .ZN(n8531) );
  NAND2_X1 U10936 ( .A1(n8518), .A2(n8531), .ZN(n14978) );
  INV_X1 U10937 ( .A(n14978), .ZN(n11520) );
  OR2_X1 U10938 ( .A1(n10696), .A2(n11520), .ZN(n8519) );
  INV_X1 U10939 ( .A(n12307), .ZN(n15095) );
  INV_X1 U10940 ( .A(n12441), .ZN(n12306) );
  INV_X1 U10941 ( .A(n11602), .ZN(n8538) );
  NAND2_X1 U10942 ( .A1(n11148), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8527) );
  NAND2_X1 U10943 ( .A1(n11147), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8526) );
  NAND2_X1 U10944 ( .A1(n8522), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8523) );
  NAND2_X1 U10945 ( .A1(n8539), .A2(n8523), .ZN(n11603) );
  NAND2_X1 U10946 ( .A1(n6885), .A2(n11603), .ZN(n8525) );
  NAND2_X1 U10947 ( .A1(n11146), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8524) );
  NAND2_X1 U10948 ( .A1(n9619), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8547) );
  NAND2_X1 U10949 ( .A1(n9621), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8530) );
  XNOR2_X1 U10950 ( .A(n8546), .B(n8545), .ZN(n14411) );
  NAND2_X1 U10951 ( .A1(n14411), .A2(n12212), .ZN(n8537) );
  NAND2_X1 U10952 ( .A1(n8531), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8532) );
  MUX2_X1 U10953 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8532), .S(
        P3_IR_REG_10__SCAN_IN), .Z(n8535) );
  INV_X1 U10954 ( .A(n8533), .ZN(n8534) );
  AOI22_X1 U10955 ( .A1(n8687), .A2(n14409), .B1(n8846), .B2(n14414), .ZN(
        n8536) );
  NAND2_X1 U10956 ( .A1(n12819), .A2(n11604), .ZN(n12310) );
  INV_X1 U10957 ( .A(n11604), .ZN(n15101) );
  NAND2_X1 U10958 ( .A1(n12440), .A2(n15101), .ZN(n12311) );
  NAND2_X1 U10959 ( .A1(n12310), .A2(n12311), .ZN(n12313) );
  NAND2_X1 U10960 ( .A1(n11148), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8544) );
  NAND2_X1 U10961 ( .A1(n11147), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8543) );
  OR2_X2 U10962 ( .A1(n8539), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8571) );
  NAND2_X1 U10963 ( .A1(n8539), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8540) );
  NAND2_X1 U10964 ( .A1(n8571), .A2(n8540), .ZN(n12821) );
  NAND2_X1 U10965 ( .A1(n6885), .A2(n12821), .ZN(n8542) );
  NAND2_X1 U10966 ( .A1(n11146), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8541) );
  NAND4_X1 U10967 ( .A1(n8544), .A2(n8543), .A3(n8542), .A4(n8541), .ZN(n12439) );
  NAND2_X1 U10968 ( .A1(n9776), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8558) );
  NAND2_X1 U10969 ( .A1(n9719), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8548) );
  OR2_X1 U10970 ( .A1(n8550), .A2(n8549), .ZN(n8551) );
  NAND2_X1 U10971 ( .A1(n8559), .A2(n8551), .ZN(n9551) );
  NAND2_X1 U10972 ( .A1(n9551), .A2(n12212), .ZN(n8557) );
  NOR2_X1 U10973 ( .A1(n8533), .A2(n6991), .ZN(n8552) );
  MUX2_X1 U10974 ( .A(n6991), .B(n8552), .S(P3_IR_REG_11__SCAN_IN), .Z(n8555)
         );
  NAND2_X1 U10975 ( .A1(n8533), .A2(n8553), .ZN(n8565) );
  INV_X1 U10976 ( .A(n8565), .ZN(n8554) );
  AOI22_X1 U10977 ( .A1(n8687), .A2(n9550), .B1(n8846), .B2(n11700), .ZN(n8556) );
  NAND2_X1 U10978 ( .A1(n8557), .A2(n8556), .ZN(n14493) );
  NAND2_X1 U10979 ( .A1(n14493), .A2(n12439), .ZN(n12323) );
  NAND2_X1 U10980 ( .A1(n12318), .A2(n12323), .ZN(n12814) );
  NAND2_X1 U10981 ( .A1(n12811), .A2(n12318), .ZN(n14475) );
  NAND2_X1 U10982 ( .A1(n9977), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8578) );
  NAND2_X1 U10983 ( .A1(n9892), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n8560) );
  OR2_X1 U10984 ( .A1(n8562), .A2(n8561), .ZN(n8563) );
  NAND2_X1 U10985 ( .A1(n8579), .A2(n8563), .ZN(n9577) );
  OR2_X1 U10986 ( .A1(n9577), .A2(n8637), .ZN(n8568) );
  NAND2_X1 U10987 ( .A1(n8565), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8564) );
  MUX2_X1 U10988 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8564), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n8566) );
  AOI22_X1 U10989 ( .A1(n8687), .A2(SI_12_), .B1(n8846), .B2(n12454), .ZN(
        n8567) );
  NAND2_X1 U10990 ( .A1(n8568), .A2(n8567), .ZN(n14486) );
  NAND2_X1 U10991 ( .A1(n8571), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8572) );
  NAND2_X1 U10992 ( .A1(n8587), .A2(n8572), .ZN(n14477) );
  NAND2_X1 U10993 ( .A1(n6885), .A2(n14477), .ZN(n8576) );
  NAND2_X1 U10994 ( .A1(n11147), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8575) );
  NAND2_X1 U10995 ( .A1(n11146), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8574) );
  OR2_X1 U10996 ( .A1(n14486), .A2(n12820), .ZN(n12324) );
  NAND2_X1 U10997 ( .A1(n14486), .A2(n12820), .ZN(n12326) );
  NAND2_X1 U10998 ( .A1(n12324), .A2(n12326), .ZN(n14466) );
  INV_X1 U10999 ( .A(n14466), .ZN(n14474) );
  NAND2_X1 U11000 ( .A1(n14475), .A2(n14474), .ZN(n8577) );
  NAND2_X1 U11001 ( .A1(n8577), .A2(n12326), .ZN(n12807) );
  NAND2_X1 U11002 ( .A1(n8581), .A2(n10155), .ZN(n8582) );
  NAND2_X1 U11003 ( .A1(n8594), .A2(n8582), .ZN(n9597) );
  OR2_X1 U11004 ( .A1(n9597), .A2(n8637), .ZN(n8585) );
  NAND2_X1 U11005 ( .A1(n8684), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8583) );
  XNOR2_X1 U11006 ( .A(n8583), .B(P3_IR_REG_13__SCAN_IN), .ZN(n12483) );
  AOI22_X1 U11007 ( .A1(n8687), .A2(SI_13_), .B1(n8846), .B2(n12483), .ZN(
        n8584) );
  NAND2_X1 U11008 ( .A1(n11148), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8592) );
  NAND2_X1 U11009 ( .A1(n11147), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8591) );
  NAND2_X1 U11010 ( .A1(n8587), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8588) );
  NAND2_X1 U11011 ( .A1(n8603), .A2(n8588), .ZN(n11589) );
  NAND2_X1 U11012 ( .A1(n6885), .A2(n11589), .ZN(n8590) );
  NAND2_X1 U11013 ( .A1(n11146), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n8589) );
  NAND4_X1 U11014 ( .A1(n8592), .A2(n8591), .A3(n8590), .A4(n8589), .ZN(n12438) );
  AND2_X1 U11015 ( .A1(n14484), .A2(n14470), .ZN(n12328) );
  OR2_X1 U11016 ( .A1(n14484), .A2(n14470), .ZN(n12320) );
  OAI21_X1 U11017 ( .B1(n12807), .B2(n12328), .A(n12320), .ZN(n12791) );
  NAND2_X1 U11018 ( .A1(n10350), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8609) );
  NAND2_X1 U11019 ( .A1(n15254), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8595) );
  OR2_X1 U11020 ( .A1(n8597), .A2(n8596), .ZN(n8598) );
  NAND2_X1 U11021 ( .A1(n8610), .A2(n8598), .ZN(n9617) );
  OR2_X1 U11022 ( .A1(n9617), .A2(n8637), .ZN(n8602) );
  NAND2_X1 U11023 ( .A1(n8615), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8600) );
  INV_X1 U11024 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8599) );
  XNOR2_X1 U11025 ( .A(n8600), .B(n8599), .ZN(n12495) );
  INV_X1 U11026 ( .A(n12495), .ZN(n12479) );
  AOI22_X1 U11027 ( .A1(n8687), .A2(SI_14_), .B1(n8846), .B2(n12479), .ZN(
        n8601) );
  NAND2_X1 U11028 ( .A1(n8602), .A2(n8601), .ZN(n12794) );
  NAND2_X1 U11029 ( .A1(n11148), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8608) );
  NAND2_X1 U11030 ( .A1(n11147), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8607) );
  NAND2_X1 U11031 ( .A1(n8603), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8604) );
  NAND2_X1 U11032 ( .A1(n8625), .A2(n8604), .ZN(n12795) );
  NAND2_X1 U11033 ( .A1(n6885), .A2(n12795), .ZN(n8606) );
  NAND2_X1 U11034 ( .A1(n11146), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8605) );
  OR2_X1 U11035 ( .A1(n12794), .A2(n12778), .ZN(n12333) );
  NAND2_X1 U11036 ( .A1(n12794), .A2(n12778), .ZN(n12334) );
  NAND2_X1 U11037 ( .A1(n12333), .A2(n12334), .ZN(n12788) );
  NAND2_X1 U11038 ( .A1(n10405), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8631) );
  NAND2_X1 U11039 ( .A1(n10387), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8611) );
  OR2_X1 U11040 ( .A1(n8613), .A2(n8612), .ZN(n8614) );
  NAND2_X1 U11041 ( .A1(n8632), .A2(n8614), .ZN(n9623) );
  OR2_X1 U11042 ( .A1(n9623), .A2(n8637), .ZN(n8623) );
  NOR2_X1 U11043 ( .A1(n8615), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n8619) );
  NOR2_X1 U11044 ( .A1(n8619), .A2(n6991), .ZN(n8616) );
  MUX2_X1 U11045 ( .A(n6991), .B(n8616), .S(P3_IR_REG_15__SCAN_IN), .Z(n8617)
         );
  INV_X1 U11046 ( .A(n8617), .ZN(n8620) );
  INV_X1 U11047 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8618) );
  NAND2_X1 U11048 ( .A1(n8619), .A2(n8618), .ZN(n8639) );
  NAND2_X1 U11049 ( .A1(n8620), .A2(n8639), .ZN(n12525) );
  OAI22_X1 U11050 ( .A1(n12213), .A2(n9622), .B1(n12525), .B2(n6390), .ZN(
        n8621) );
  INV_X1 U11051 ( .A(n8621), .ZN(n8622) );
  NAND2_X1 U11052 ( .A1(n11148), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8630) );
  NAND2_X1 U11053 ( .A1(n11147), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8629) );
  NAND2_X1 U11054 ( .A1(n8625), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8626) );
  NAND2_X1 U11055 ( .A1(n8644), .A2(n8626), .ZN(n12782) );
  NAND2_X1 U11056 ( .A1(n6885), .A2(n12782), .ZN(n8628) );
  NAND2_X1 U11057 ( .A1(n11146), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8627) );
  XNOR2_X1 U11058 ( .A(n12337), .B(n12790), .ZN(n12776) );
  INV_X1 U11059 ( .A(n12776), .ZN(n12781) );
  NAND2_X1 U11060 ( .A1(n12337), .A2(n12790), .ZN(n12342) );
  NAND2_X1 U11061 ( .A1(n10346), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8650) );
  NAND2_X1 U11062 ( .A1(n10349), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8633) );
  OR2_X1 U11063 ( .A1(n8635), .A2(n8634), .ZN(n8636) );
  NAND2_X1 U11064 ( .A1(n8651), .A2(n8636), .ZN(n9687) );
  OR2_X1 U11065 ( .A1(n9687), .A2(n8637), .ZN(n8643) );
  NAND2_X1 U11066 ( .A1(n8639), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8638) );
  MUX2_X1 U11067 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8638), .S(
        P3_IR_REG_16__SCAN_IN), .Z(n8640) );
  NAND2_X1 U11068 ( .A1(n8640), .A2(n8668), .ZN(n12550) );
  OAI22_X1 U11069 ( .A1(n12213), .A2(n9686), .B1(n12550), .B2(n10696), .ZN(
        n8641) );
  INV_X1 U11070 ( .A(n8641), .ZN(n8642) );
  NAND2_X1 U11071 ( .A1(n11147), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8648) );
  NAND2_X1 U11072 ( .A1(n8644), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8645) );
  NAND2_X1 U11073 ( .A1(n8657), .A2(n8645), .ZN(n12770) );
  NAND2_X1 U11074 ( .A1(n6885), .A2(n12770), .ZN(n8647) );
  NAND2_X1 U11075 ( .A1(n11146), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8646) );
  NAND4_X1 U11076 ( .A1(n8649), .A2(n8648), .A3(n8647), .A4(n8646), .ZN(n12751) );
  INV_X1 U11077 ( .A(n12751), .ZN(n12779) );
  OR2_X1 U11078 ( .A1(n12769), .A2(n12779), .ZN(n12344) );
  NAND2_X1 U11079 ( .A1(n12769), .A2(n12779), .ZN(n12343) );
  NAND2_X1 U11080 ( .A1(n12768), .A2(n12767), .ZN(n12766) );
  NAND2_X1 U11081 ( .A1(n12766), .A2(n12343), .ZN(n12757) );
  NAND2_X1 U11082 ( .A1(n10385), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8666) );
  NAND2_X1 U11083 ( .A1(n10400), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8652) );
  NAND2_X1 U11084 ( .A1(n8666), .A2(n8652), .ZN(n8663) );
  XNOR2_X1 U11085 ( .A(n8665), .B(n8663), .ZN(n9990) );
  NAND2_X1 U11086 ( .A1(n9990), .A2(n12212), .ZN(n8655) );
  NAND2_X1 U11087 ( .A1(n8668), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8653) );
  XNOR2_X1 U11088 ( .A(n8653), .B(P3_IR_REG_17__SCAN_IN), .ZN(n14450) );
  AOI22_X1 U11089 ( .A1(SI_17_), .A2(n8687), .B1(n14450), .B2(n8846), .ZN(
        n8654) );
  NAND2_X1 U11090 ( .A1(n8657), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8658) );
  NAND2_X1 U11091 ( .A1(n8672), .A2(n8658), .ZN(n12758) );
  NAND2_X1 U11092 ( .A1(n12758), .A2(n6885), .ZN(n8662) );
  NAND2_X1 U11093 ( .A1(n11148), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8661) );
  NAND2_X1 U11094 ( .A1(n11147), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8660) );
  NAND2_X1 U11095 ( .A1(n11146), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8659) );
  NAND4_X1 U11096 ( .A1(n8662), .A2(n8661), .A3(n8660), .A4(n8659), .ZN(n12349) );
  XNOR2_X1 U11097 ( .A(n12348), .B(n12349), .ZN(n12756) );
  NAND2_X1 U11098 ( .A1(n12348), .A2(n12765), .ZN(n12353) );
  INV_X1 U11099 ( .A(n8663), .ZN(n8664) );
  INV_X1 U11100 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10761) );
  NAND2_X1 U11101 ( .A1(n10761), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8680) );
  INV_X1 U11102 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10763) );
  NAND2_X1 U11103 ( .A1(n10763), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8667) );
  NAND2_X1 U11104 ( .A1(n8680), .A2(n8667), .ZN(n8677) );
  XNOR2_X1 U11105 ( .A(n8679), .B(n8677), .ZN(n10073) );
  NAND2_X1 U11106 ( .A1(n10073), .A2(n12212), .ZN(n8671) );
  OAI21_X1 U11107 ( .B1(n8668), .B2(P3_IR_REG_17__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8669) );
  XNOR2_X1 U11108 ( .A(n8669), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12582) );
  AOI22_X1 U11109 ( .A1(n12582), .A2(n8846), .B1(n8687), .B2(SI_18_), .ZN(
        n8670) );
  NAND2_X1 U11110 ( .A1(n8672), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8673) );
  NAND2_X1 U11111 ( .A1(n8692), .A2(n8673), .ZN(n12180) );
  NAND2_X1 U11112 ( .A1(n12180), .A2(n6885), .ZN(n8676) );
  NAND2_X1 U11113 ( .A1(n11146), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8674) );
  NAND2_X1 U11114 ( .A1(n12880), .A2(n12726), .ZN(n12355) );
  INV_X1 U11115 ( .A(n12728), .ZN(n8698) );
  INV_X1 U11116 ( .A(n8677), .ZN(n8678) );
  NAND2_X1 U11117 ( .A1(n10993), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8701) );
  NAND2_X1 U11118 ( .A1(n10995), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8682) );
  XNOR2_X1 U11119 ( .A(n8700), .B(n8699), .ZN(n10157) );
  NAND2_X1 U11120 ( .A1(n10157), .A2(n12212), .ZN(n8689) );
  AOI22_X1 U11121 ( .A1(n8687), .A2(n10156), .B1(n8846), .B2(n12594), .ZN(
        n8688) );
  INV_X1 U11122 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n8690) );
  NAND2_X1 U11123 ( .A1(n8692), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8693) );
  NAND2_X1 U11124 ( .A1(n8705), .A2(n8693), .ZN(n12730) );
  NAND2_X1 U11125 ( .A1(n12730), .A2(n6885), .ZN(n8696) );
  AOI22_X1 U11126 ( .A1(n11147), .A2(P3_REG1_REG_19__SCAN_IN), .B1(n11148), 
        .B2(P3_REG0_REG_19__SCAN_IN), .ZN(n8695) );
  NAND2_X1 U11127 ( .A1(n11146), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n8694) );
  AND2_X1 U11128 ( .A1(n12935), .A2(n12713), .ZN(n12362) );
  INV_X1 U11129 ( .A(n12362), .ZN(n8697) );
  OR2_X1 U11130 ( .A1(n12935), .A2(n12713), .ZN(n12363) );
  XNOR2_X1 U11131 ( .A(n8712), .B(n11352), .ZN(n10401) );
  NAND2_X1 U11132 ( .A1(n10401), .A2(n12212), .ZN(n8704) );
  OR2_X1 U11133 ( .A1(n12213), .A2(n10402), .ZN(n8703) );
  NAND2_X1 U11134 ( .A1(n8705), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8706) );
  NAND2_X1 U11135 ( .A1(n8720), .A2(n8706), .ZN(n12716) );
  NAND2_X1 U11136 ( .A1(n12716), .A2(n6885), .ZN(n8711) );
  INV_X1 U11137 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n12718) );
  NAND2_X1 U11138 ( .A1(n11147), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n8707) );
  OAI211_X1 U11139 ( .C1(n12718), .C2(n8932), .A(n8708), .B(n8707), .ZN(n8709)
         );
  INV_X1 U11140 ( .A(n8709), .ZN(n8710) );
  XNOR2_X1 U11141 ( .A(n12871), .B(n12727), .ZN(n12720) );
  OR2_X1 U11142 ( .A1(n12871), .A2(n12727), .ZN(n12366) );
  INV_X1 U11143 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11563) );
  NAND2_X1 U11144 ( .A1(n11563), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8734) );
  INV_X1 U11145 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11397) );
  NAND2_X1 U11146 ( .A1(n11397), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8715) );
  NAND2_X1 U11147 ( .A1(n8734), .A2(n8715), .ZN(n8731) );
  XNOR2_X1 U11148 ( .A(n8733), .B(n8731), .ZN(n10669) );
  NAND2_X1 U11149 ( .A1(n10669), .A2(n12212), .ZN(n8717) );
  INV_X1 U11150 ( .A(SI_21_), .ZN(n10670) );
  OR2_X1 U11151 ( .A1(n12213), .A2(n10670), .ZN(n8716) );
  INV_X1 U11152 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n8718) );
  NAND2_X1 U11153 ( .A1(n8720), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8721) );
  NAND2_X1 U11154 ( .A1(n8738), .A2(n8721), .ZN(n12706) );
  NAND2_X1 U11155 ( .A1(n12706), .A2(n6885), .ZN(n8727) );
  INV_X1 U11156 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n8724) );
  NAND2_X1 U11157 ( .A1(n11148), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8723) );
  NAND2_X1 U11158 ( .A1(n11147), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8722) );
  OAI211_X1 U11159 ( .C1(n8724), .C2(n8932), .A(n8723), .B(n8722), .ZN(n8725)
         );
  INV_X1 U11160 ( .A(n8725), .ZN(n8726) );
  NAND2_X1 U11161 ( .A1(n12705), .A2(n12690), .ZN(n8728) );
  NAND2_X1 U11162 ( .A1(n12704), .A2(n8728), .ZN(n8730) );
  OR2_X1 U11163 ( .A1(n12705), .A2(n12690), .ZN(n8729) );
  NAND2_X1 U11164 ( .A1(n8730), .A2(n8729), .ZN(n12693) );
  INV_X1 U11165 ( .A(n8731), .ZN(n8732) );
  INV_X1 U11166 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8749) );
  XNOR2_X1 U11167 ( .A(n8749), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n8747) );
  XNOR2_X1 U11168 ( .A(n8748), .B(n8747), .ZN(n10672) );
  NAND2_X1 U11169 ( .A1(n10672), .A2(n12212), .ZN(n8737) );
  INV_X1 U11170 ( .A(SI_22_), .ZN(n8735) );
  OR2_X1 U11171 ( .A1(n12213), .A2(n8735), .ZN(n8736) );
  OR2_X2 U11172 ( .A1(n8738), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8753) );
  NAND2_X1 U11173 ( .A1(n8738), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8739) );
  NAND2_X1 U11174 ( .A1(n8753), .A2(n8739), .ZN(n12695) );
  NAND2_X1 U11175 ( .A1(n12695), .A2(n6885), .ZN(n8745) );
  INV_X1 U11176 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n8742) );
  NAND2_X1 U11177 ( .A1(n11148), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8741) );
  NAND2_X1 U11178 ( .A1(n11147), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8740) );
  OAI211_X1 U11179 ( .C1(n8742), .C2(n8932), .A(n8741), .B(n8740), .ZN(n8743)
         );
  INV_X1 U11180 ( .A(n8743), .ZN(n8744) );
  NAND2_X1 U11181 ( .A1(n12694), .A2(n12702), .ZN(n12251) );
  NAND2_X1 U11182 ( .A1(n12693), .A2(n12251), .ZN(n8746) );
  NAND2_X1 U11183 ( .A1(n8746), .A2(n12250), .ZN(n12671) );
  NAND2_X1 U11184 ( .A1(n8749), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8750) );
  XNOR2_X1 U11185 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n8760) );
  XNOR2_X1 U11186 ( .A(n8761), .B(n8760), .ZN(n10989) );
  NAND2_X1 U11187 ( .A1(n10989), .A2(n12212), .ZN(n8752) );
  INV_X1 U11188 ( .A(SI_23_), .ZN(n10991) );
  OR2_X1 U11189 ( .A1(n12213), .A2(n10991), .ZN(n8751) );
  OR2_X2 U11190 ( .A1(n8753), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8770) );
  NAND2_X1 U11191 ( .A1(n8753), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8754) );
  NAND2_X1 U11192 ( .A1(n8770), .A2(n8754), .ZN(n12680) );
  NAND2_X1 U11193 ( .A1(n12680), .A2(n6885), .ZN(n8759) );
  INV_X1 U11194 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n12681) );
  NAND2_X1 U11195 ( .A1(n11148), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8756) );
  NAND2_X1 U11196 ( .A1(n11147), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8755) );
  OAI211_X1 U11197 ( .C1(n12681), .C2(n8932), .A(n8756), .B(n8755), .ZN(n8757)
         );
  INV_X1 U11198 ( .A(n8757), .ZN(n8758) );
  NAND2_X1 U11199 ( .A1(n12684), .A2(n12691), .ZN(n12379) );
  INV_X1 U11200 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8762) );
  NAND2_X1 U11201 ( .A1(n8762), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8763) );
  INV_X1 U11202 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n13613) );
  XNOR2_X1 U11203 ( .A(n8778), .B(n7156), .ZN(n11268) );
  NAND2_X1 U11204 ( .A1(n11268), .A2(n12212), .ZN(n8767) );
  INV_X1 U11205 ( .A(SI_24_), .ZN(n11269) );
  OR2_X1 U11206 ( .A1(n12213), .A2(n11269), .ZN(n8766) );
  INV_X1 U11207 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n8768) );
  NAND2_X1 U11208 ( .A1(n8770), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8771) );
  NAND2_X1 U11209 ( .A1(n8783), .A2(n8771), .ZN(n12663) );
  NAND2_X1 U11210 ( .A1(n12663), .A2(n6885), .ZN(n8776) );
  INV_X1 U11211 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n12664) );
  NAND2_X1 U11212 ( .A1(n11147), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8772) );
  OAI211_X1 U11213 ( .C1(n12664), .C2(n8932), .A(n8773), .B(n8772), .ZN(n8774)
         );
  INV_X1 U11214 ( .A(n8774), .ZN(n8775) );
  NAND2_X1 U11215 ( .A1(n12667), .A2(n12676), .ZN(n12383) );
  INV_X1 U11216 ( .A(n12383), .ZN(n8777) );
  XNOR2_X1 U11217 ( .A(n13608), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n8779) );
  XNOR2_X1 U11218 ( .A(n8793), .B(n8779), .ZN(n11450) );
  NAND2_X1 U11219 ( .A1(n11450), .A2(n12212), .ZN(n8781) );
  OR2_X1 U11220 ( .A1(n12213), .A2(n11452), .ZN(n8780) );
  INV_X1 U11221 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n15121) );
  NAND2_X1 U11222 ( .A1(n8783), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8784) );
  NAND2_X1 U11223 ( .A1(n8798), .A2(n8784), .ZN(n12653) );
  NAND2_X1 U11224 ( .A1(n12653), .A2(n6885), .ZN(n8790) );
  INV_X1 U11225 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n8787) );
  NAND2_X1 U11226 ( .A1(n11147), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8785) );
  OAI211_X1 U11227 ( .C1(n8787), .C2(n8932), .A(n8786), .B(n8785), .ZN(n8788)
         );
  INV_X1 U11228 ( .A(n8788), .ZN(n8789) );
  NAND2_X1 U11229 ( .A1(n12247), .A2(n12433), .ZN(n12248) );
  OR2_X1 U11230 ( .A1(n12247), .A2(n12433), .ZN(n8791) );
  NAND2_X1 U11231 ( .A1(n13608), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8792) );
  NAND2_X1 U11232 ( .A1(n14295), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8794) );
  XNOR2_X1 U11233 ( .A(n8809), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n8795) );
  XNOR2_X1 U11234 ( .A(n8808), .B(n8795), .ZN(n11580) );
  NAND2_X1 U11235 ( .A1(n11580), .A2(n12212), .ZN(n8797) );
  OR2_X1 U11236 ( .A1(n12213), .A2(n11582), .ZN(n8796) );
  NAND2_X1 U11237 ( .A1(n8798), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8799) );
  NAND2_X1 U11238 ( .A1(n8815), .A2(n8799), .ZN(n12642) );
  NAND2_X1 U11239 ( .A1(n12642), .A2(n6885), .ZN(n8805) );
  INV_X1 U11240 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n8802) );
  NAND2_X1 U11241 ( .A1(n11147), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8800) );
  OAI211_X1 U11242 ( .C1(n8802), .C2(n8932), .A(n8801), .B(n8800), .ZN(n8803)
         );
  INV_X1 U11243 ( .A(n8803), .ZN(n8804) );
  NAND2_X1 U11244 ( .A1(n12388), .A2(n12652), .ZN(n12395) );
  INV_X1 U11245 ( .A(n12395), .ZN(n8806) );
  AND2_X1 U11246 ( .A1(n14292), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8807) );
  NAND2_X1 U11247 ( .A1(n8809), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8810) );
  XNOR2_X1 U11248 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n8811) );
  XNOR2_X1 U11249 ( .A(n8823), .B(n8811), .ZN(n11651) );
  NAND2_X1 U11250 ( .A1(n11651), .A2(n12212), .ZN(n8813) );
  OR2_X1 U11251 ( .A1(n12213), .A2(n11652), .ZN(n8812) );
  INV_X1 U11252 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n12093) );
  NAND2_X1 U11253 ( .A1(n8815), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8816) );
  NAND2_X1 U11254 ( .A1(n8828), .A2(n8816), .ZN(n12630) );
  NAND2_X1 U11255 ( .A1(n12630), .A2(n6885), .ZN(n8821) );
  INV_X1 U11256 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n12631) );
  NAND2_X1 U11257 ( .A1(n11148), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8818) );
  NAND2_X1 U11258 ( .A1(n11147), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8817) );
  OAI211_X1 U11259 ( .C1(n12631), .C2(n8932), .A(n8818), .B(n8817), .ZN(n8819)
         );
  INV_X1 U11260 ( .A(n8819), .ZN(n8820) );
  AND2_X2 U11261 ( .A1(n8821), .A2(n8820), .ZN(n12641) );
  AND2_X1 U11262 ( .A1(n13599), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8822) );
  XNOR2_X1 U11263 ( .A(n15244), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n8825) );
  XNOR2_X1 U11264 ( .A(n8923), .B(n8825), .ZN(n12970) );
  NAND2_X1 U11265 ( .A1(n12970), .A2(n12212), .ZN(n8827) );
  OR2_X1 U11266 ( .A1(n12213), .A2(n12972), .ZN(n8826) );
  NAND2_X1 U11267 ( .A1(n8828), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8829) );
  NAND2_X1 U11268 ( .A1(n8879), .A2(n8829), .ZN(n12115) );
  INV_X1 U11269 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n12617) );
  NAND2_X1 U11270 ( .A1(n8416), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8831) );
  NAND2_X1 U11271 ( .A1(n11148), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8830) );
  OAI211_X1 U11272 ( .C1(n12617), .C2(n8932), .A(n8831), .B(n8830), .ZN(n8832)
         );
  AOI21_X2 U11273 ( .B1(n12115), .B2(n6885), .A(n8832), .ZN(n12629) );
  NAND2_X1 U11274 ( .A1(n12620), .A2(n12629), .ZN(n12393) );
  XNOR2_X1 U11275 ( .A(n6446), .B(n12391), .ZN(n12616) );
  NAND2_X1 U11276 ( .A1(n8886), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8833) );
  NAND2_X1 U11277 ( .A1(n8834), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8835) );
  NAND2_X1 U11278 ( .A1(n8836), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8837) );
  NOR2_X1 U11279 ( .A1(n12253), .A2(n8877), .ZN(n8951) );
  INV_X1 U11280 ( .A(n8951), .ZN(n8838) );
  XNOR2_X1 U11281 ( .A(n12424), .B(n8838), .ZN(n8840) );
  NAND2_X1 U11282 ( .A1(n12594), .A2(n12258), .ZN(n8839) );
  NAND2_X1 U11283 ( .A1(n8840), .A2(n8839), .ZN(n10239) );
  INV_X1 U11284 ( .A(n12424), .ZN(n8841) );
  NAND3_X1 U11285 ( .A1(n10239), .A2(n12419), .A3(n15100), .ZN(n8843) );
  AND3_X1 U11286 ( .A1(n12424), .A2(n12594), .A3(n8877), .ZN(n10656) );
  INV_X1 U11287 ( .A(n10656), .ZN(n8842) );
  NAND2_X1 U11288 ( .A1(n8843), .A2(n8842), .ZN(n15106) );
  NOR2_X1 U11289 ( .A1(n15075), .A2(n12424), .ZN(n15099) );
  INV_X1 U11290 ( .A(n12974), .ZN(n8845) );
  INV_X1 U11291 ( .A(n12422), .ZN(n8847) );
  NAND2_X1 U11292 ( .A1(n15065), .A2(n10665), .ZN(n10252) );
  NAND2_X1 U11293 ( .A1(n15063), .A2(n10252), .ZN(n8849) );
  NAND2_X1 U11294 ( .A1(n15047), .A2(n10248), .ZN(n8848) );
  NAND2_X1 U11295 ( .A1(n8849), .A2(n8848), .ZN(n15050) );
  NAND2_X1 U11296 ( .A1(n8850), .A2(n6395), .ZN(n8851) );
  NAND2_X1 U11297 ( .A1(n12448), .A2(n10756), .ZN(n8853) );
  NAND2_X1 U11298 ( .A1(n12446), .A2(n15035), .ZN(n8855) );
  NAND2_X1 U11299 ( .A1(n11116), .A2(n11251), .ZN(n8857) );
  NAND2_X1 U11300 ( .A1(n12444), .A2(n15025), .ZN(n8858) );
  NAND2_X1 U11301 ( .A1(n12443), .A2(n10884), .ZN(n8859) );
  NAND2_X1 U11302 ( .A1(n11612), .A2(n12299), .ZN(n8860) );
  XNOR2_X1 U11303 ( .A(n12441), .B(n12307), .ZN(n12303) );
  NAND2_X1 U11304 ( .A1(n12441), .A2(n12307), .ZN(n8861) );
  NAND2_X1 U11305 ( .A1(n11614), .A2(n8861), .ZN(n11597) );
  NAND2_X1 U11306 ( .A1(n11597), .A2(n12313), .ZN(n11596) );
  NAND2_X1 U11307 ( .A1(n11604), .A2(n12440), .ZN(n8862) );
  INV_X1 U11308 ( .A(n12439), .ZN(n14471) );
  NAND2_X1 U11309 ( .A1(n14493), .A2(n14471), .ZN(n14467) );
  AND2_X1 U11310 ( .A1(n14466), .A2(n14467), .ZN(n8863) );
  NAND2_X1 U11311 ( .A1(n14486), .A2(n12801), .ZN(n8864) );
  OR2_X1 U11312 ( .A1(n14484), .A2(n12438), .ZN(n8865) );
  INV_X1 U11313 ( .A(n12778), .ZN(n12802) );
  NAND2_X1 U11314 ( .A1(n12794), .A2(n12802), .ZN(n8866) );
  NAND2_X1 U11315 ( .A1(n12337), .A2(n12437), .ZN(n8868) );
  AND2_X1 U11316 ( .A1(n12769), .A2(n12751), .ZN(n8869) );
  OR2_X1 U11317 ( .A1(n12769), .A2(n12751), .ZN(n8870) );
  NAND2_X1 U11318 ( .A1(n12348), .A2(n12349), .ZN(n8873) );
  INV_X1 U11319 ( .A(n12726), .ZN(n12752) );
  AND2_X1 U11320 ( .A1(n12935), .A2(n12742), .ZN(n8874) );
  INV_X1 U11321 ( .A(n12727), .ZN(n12436) );
  NAND2_X1 U11322 ( .A1(n12871), .A2(n12436), .ZN(n8875) );
  AND2_X1 U11323 ( .A1(n12705), .A2(n12714), .ZN(n12373) );
  INV_X1 U11324 ( .A(n12652), .ZN(n12432) );
  AOI22_X1 U11325 ( .A1(n12627), .A2(n12628), .B1(n12641), .B2(n12909), .ZN(
        n8878) );
  NAND2_X1 U11326 ( .A1(n8878), .A2(n12391), .ZN(n8921) );
  INV_X1 U11327 ( .A(n12594), .ZN(n12219) );
  NAND2_X1 U11328 ( .A1(n12219), .A2(n12424), .ZN(n8950) );
  NAND2_X1 U11329 ( .A1(n12253), .A2(n8877), .ZN(n12245) );
  INV_X1 U11330 ( .A(n8879), .ZN(n12603) );
  NAND2_X1 U11331 ( .A1(n12603), .A2(n6885), .ZN(n11153) );
  INV_X1 U11332 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n12611) );
  NAND2_X1 U11333 ( .A1(n11147), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8881) );
  NAND2_X1 U11334 ( .A1(n11148), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8880) );
  OAI211_X1 U11335 ( .C1(n8932), .C2(n12611), .A(n8881), .B(n8880), .ZN(n8882)
         );
  INV_X1 U11336 ( .A(n8882), .ZN(n8883) );
  NAND2_X1 U11337 ( .A1(n11153), .A2(n8883), .ZN(n12430) );
  NAND2_X1 U11338 ( .A1(n12430), .A2(n15067), .ZN(n8884) );
  OAI211_X1 U11339 ( .C1(n12641), .C2(n15046), .A(n8885), .B(n8884), .ZN(
        n12621) );
  INV_X1 U11340 ( .A(P3_B_REG_SCAN_IN), .ZN(n8936) );
  INV_X1 U11341 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n8889) );
  NOR4_X1 U11342 ( .A1(P3_D_REG_20__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_27__SCAN_IN), .ZN(n8901) );
  OR4_X1 U11343 ( .A1(P3_D_REG_22__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_17__SCAN_IN), .A4(P3_D_REG_25__SCAN_IN), .ZN(n8898) );
  NOR4_X1 U11344 ( .A1(P3_D_REG_26__SCAN_IN), .A2(P3_D_REG_9__SCAN_IN), .A3(
        P3_D_REG_16__SCAN_IN), .A4(P3_D_REG_15__SCAN_IN), .ZN(n8896) );
  NOR4_X1 U11345 ( .A1(P3_D_REG_12__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_11__SCAN_IN), .ZN(n8895) );
  NOR4_X1 U11346 ( .A1(P3_D_REG_6__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8894) );
  NOR4_X1 U11347 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_13__SCAN_IN), .A3(
        P3_D_REG_28__SCAN_IN), .A4(P3_D_REG_23__SCAN_IN), .ZN(n8893) );
  NAND4_X1 U11348 ( .A1(n8896), .A2(n8895), .A3(n8894), .A4(n8893), .ZN(n8897)
         );
  NOR4_X1 U11349 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        n8898), .A4(n8897), .ZN(n8900) );
  NOR4_X1 U11350 ( .A1(P3_D_REG_24__SCAN_IN), .A2(P3_D_REG_29__SCAN_IN), .A3(
        P3_D_REG_10__SCAN_IN), .A4(P3_D_REG_31__SCAN_IN), .ZN(n8899) );
  NAND3_X1 U11351 ( .A1(n8901), .A2(n8900), .A3(n8899), .ZN(n8902) );
  NAND2_X1 U11352 ( .A1(n8892), .A2(n8902), .ZN(n8946) );
  NAND2_X1 U11353 ( .A1(n6938), .A2(n8946), .ZN(n8906) );
  INV_X1 U11354 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n8903) );
  NAND2_X1 U11355 ( .A1(n8892), .A2(n8903), .ZN(n8905) );
  OR2_X1 U11356 ( .A1(n11579), .A2(n8907), .ZN(n8904) );
  AND2_X1 U11357 ( .A1(n8907), .A2(n11267), .ZN(n8908) );
  INV_X1 U11358 ( .A(n8909), .ZN(n8910) );
  NAND2_X1 U11359 ( .A1(n8910), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8912) );
  AND2_X1 U11360 ( .A1(n10224), .A2(n10240), .ZN(n10238) );
  NAND2_X1 U11361 ( .A1(n10238), .A2(n10239), .ZN(n8916) );
  INV_X1 U11362 ( .A(n6938), .ZN(n12960) );
  AND3_X1 U11363 ( .A1(n12960), .A2(n12958), .A3(n8946), .ZN(n10241) );
  OR2_X1 U11364 ( .A1(n8950), .A2(n12244), .ZN(n10236) );
  NAND2_X1 U11365 ( .A1(n12402), .A2(n12419), .ZN(n8913) );
  OR2_X1 U11366 ( .A1(n10693), .A2(n8913), .ZN(n12423) );
  OAI21_X1 U11367 ( .B1(n10693), .B2(n10236), .A(n12423), .ZN(n8914) );
  NAND2_X1 U11368 ( .A1(n10241), .A2(n8914), .ZN(n8915) );
  OR2_X1 U11369 ( .A1(n12837), .A2(n15110), .ZN(n8920) );
  INV_X1 U11370 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n8917) );
  INV_X1 U11371 ( .A(n8918), .ZN(n8919) );
  NAND2_X1 U11372 ( .A1(n8920), .A2(n8919), .ZN(P3_U3455) );
  NAND2_X1 U11373 ( .A1(n8921), .A2(n6448), .ZN(n8929) );
  AND2_X1 U11374 ( .A1(n11869), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8922) );
  NAND2_X1 U11375 ( .A1(n15244), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8924) );
  NAND2_X1 U11376 ( .A1(n14285), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n11847) );
  NAND2_X1 U11377 ( .A1(n13592), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8926) );
  AND2_X1 U11378 ( .A1(n11847), .A2(n8926), .ZN(n11846) );
  XNOR2_X1 U11379 ( .A(n11849), .B(n11846), .ZN(n12967) );
  NAND2_X1 U11380 ( .A1(n12967), .A2(n12212), .ZN(n8928) );
  OR2_X1 U11381 ( .A1(n12213), .A2(n15242), .ZN(n8927) );
  NAND2_X1 U11382 ( .A1(n8957), .A2(n12430), .ZN(n12411) );
  INV_X1 U11383 ( .A(n8957), .ZN(n12608) );
  INV_X1 U11384 ( .A(n12430), .ZN(n12116) );
  NAND2_X1 U11385 ( .A1(n12608), .A2(n12116), .ZN(n12206) );
  NAND2_X1 U11386 ( .A1(n12411), .A2(n12206), .ZN(n12222) );
  INV_X1 U11387 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n8933) );
  NAND2_X1 U11388 ( .A1(n8416), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8930) );
  OAI211_X1 U11389 ( .C1(n8933), .C2(n8932), .A(n8931), .B(n8930), .ZN(n8934)
         );
  INV_X1 U11390 ( .A(n8934), .ZN(n8935) );
  AND2_X1 U11391 ( .A1(n11153), .A2(n8935), .ZN(n12216) );
  OAI21_X1 U11392 ( .B1(n12974), .B2(n8936), .A(n15067), .ZN(n12601) );
  NOR2_X1 U11393 ( .A1(n12216), .A2(n12601), .ZN(n8938) );
  INV_X1 U11394 ( .A(n8941), .ZN(n12399) );
  XOR2_X1 U11395 ( .A(n12222), .B(n12202), .Z(n12607) );
  INV_X1 U11396 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n8942) );
  NOR2_X1 U11397 ( .A1(n15108), .A2(n8942), .ZN(n8943) );
  NAND2_X1 U11398 ( .A1(n8945), .A2(n8944), .ZN(P3_U3456) );
  INV_X1 U11399 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n8956) );
  XNOR2_X1 U11400 ( .A(n6938), .B(n12958), .ZN(n8948) );
  AND2_X1 U11401 ( .A1(n8946), .A2(n10240), .ZN(n8947) );
  MUX2_X1 U11402 ( .A(n10656), .B(n12419), .S(n12402), .Z(n10658) );
  INV_X1 U11403 ( .A(n12419), .ZN(n8949) );
  OAI211_X1 U11404 ( .C1(n12424), .C2(n8951), .A(n8950), .B(n8949), .ZN(n8952)
         );
  AND2_X1 U11405 ( .A1(n8952), .A2(n12415), .ZN(n8954) );
  INV_X1 U11406 ( .A(n12958), .ZN(n8953) );
  MUX2_X1 U11407 ( .A(n10658), .B(n8954), .S(n8953), .Z(n8955) );
  INV_X1 U11408 ( .A(n15100), .ZN(n15073) );
  NAND2_X1 U11409 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9085) );
  NAND2_X1 U11410 ( .A1(n9094), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9112) );
  INV_X1 U11411 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n9111) );
  NAND2_X1 U11412 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .ZN(n8958) );
  NAND2_X1 U11413 ( .A1(n9173), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9185) );
  NAND2_X1 U11414 ( .A1(n9220), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9232) );
  INV_X1 U11415 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9231) );
  INV_X1 U11416 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n11428) );
  AND2_X1 U11417 ( .A1(n9234), .A2(n11428), .ZN(n8959) );
  OR2_X1 U11418 ( .A1(n8959), .A2(n9271), .ZN(n14137) );
  NOR2_X1 U11419 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n8961) );
  NAND4_X1 U11420 ( .A1(n8961), .A2(n8960), .A3(n8994), .A4(n9003), .ZN(n9498)
         );
  NAND3_X1 U11421 ( .A1(n15212), .A2(n8986), .A3(n8984), .ZN(n8962) );
  NOR3_X1 U11422 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), 
        .A3(P1_IR_REG_25__SCAN_IN), .ZN(n8963) );
  XNOR2_X2 U11423 ( .A(n8974), .B(n8973), .ZN(n14287) );
  AOI22_X1 U11424 ( .A1(n9433), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9434), .B2(
        P1_REG0_REG_16__SCAN_IN), .ZN(n8978) );
  NAND2_X1 U11425 ( .A1(n9096), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8977) );
  OAI211_X1 U11426 ( .C1(n14137), .C2(n6398), .A(n8978), .B(n8977), .ZN(n13889) );
  NAND2_X1 U11427 ( .A1(n8980), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8981) );
  INV_X1 U11428 ( .A(n9533), .ZN(n8983) );
  INV_X4 U11429 ( .A(n9440), .ZN(n9454) );
  NAND2_X1 U11430 ( .A1(n10345), .A2(n9454), .ZN(n8991) );
  NOR2_X1 U11431 ( .A1(n8987), .A2(n9227), .ZN(n8985) );
  MUX2_X1 U11432 ( .A(n9227), .B(n8985), .S(P1_IR_REG_16__SCAN_IN), .Z(n8989)
         );
  INV_X1 U11433 ( .A(n8992), .ZN(n8988) );
  OR2_X1 U11434 ( .A1(n8989), .A2(n8988), .ZN(n11444) );
  INV_X1 U11435 ( .A(n11444), .ZN(n11760) );
  AOI22_X1 U11436 ( .A1(n9277), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9276), 
        .B2(n11760), .ZN(n8990) );
  NAND2_X1 U11437 ( .A1(n9001), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8993) );
  MUX2_X1 U11438 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8993), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n8996) );
  INV_X1 U11439 ( .A(n9001), .ZN(n8995) );
  INV_X1 U11440 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8994) );
  NAND2_X1 U11441 ( .A1(n8995), .A2(n8994), .ZN(n8997) );
  NAND2_X1 U11442 ( .A1(n8994), .A2(n9000), .ZN(n9004) );
  NAND3_X1 U11443 ( .A1(n9001), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_IR_REG_22__SCAN_IN), .ZN(n9006) );
  XNOR2_X1 U11444 ( .A(P1_IR_REG_31__SCAN_IN), .B(P1_IR_REG_22__SCAN_IN), .ZN(
        n9002) );
  OAI21_X1 U11445 ( .B1(n9004), .B2(n9003), .A(n9002), .ZN(n9005) );
  NAND2_X1 U11446 ( .A1(n9008), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9010) );
  MUX2_X1 U11447 ( .A(n13889), .B(n14132), .S(n9448), .Z(n9263) );
  OR2_X1 U11448 ( .A1(n14132), .A2(n9448), .ZN(n9253) );
  INV_X1 U11449 ( .A(n9253), .ZN(n9019) );
  INV_X1 U11450 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9011) );
  XNOR2_X1 U11451 ( .A(n9271), .B(n9011), .ZN(n14121) );
  INV_X1 U11452 ( .A(n6399), .ZN(n9282) );
  NAND2_X1 U11453 ( .A1(n14121), .A2(n9282), .ZN(n9017) );
  INV_X1 U11454 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9014) );
  NAND2_X1 U11455 ( .A1(n9434), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n9013) );
  INV_X1 U11456 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n11754) );
  OR2_X1 U11457 ( .A1(n9428), .A2(n11754), .ZN(n9012) );
  OAI211_X1 U11458 ( .C1(n9014), .C2(n6400), .A(n9013), .B(n9012), .ZN(n9015)
         );
  INV_X1 U11459 ( .A(n9015), .ZN(n9016) );
  NAND2_X1 U11460 ( .A1(n9017), .A2(n9016), .ZN(n14136) );
  NAND2_X1 U11461 ( .A1(n9459), .A2(n14136), .ZN(n9255) );
  INV_X1 U11462 ( .A(n9255), .ZN(n9018) );
  AOI21_X1 U11463 ( .B1(n9263), .B2(n9019), .A(n9018), .ZN(n9266) );
  NAND2_X1 U11464 ( .A1(n10384), .A2(n9454), .ZN(n9022) );
  NAND2_X1 U11465 ( .A1(n8992), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9020) );
  XNOR2_X1 U11466 ( .A(n9020), .B(P1_IR_REG_17__SCAN_IN), .ZN(n13846) );
  AOI22_X1 U11467 ( .A1(n9277), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9276), 
        .B2(n13846), .ZN(n9021) );
  NAND2_X1 U11468 ( .A1(n9433), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9028) );
  INV_X1 U11469 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10599) );
  OR2_X1 U11470 ( .A1(n6399), .A2(n10599), .ZN(n9027) );
  INV_X1 U11471 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9591) );
  OR2_X1 U11472 ( .A1(n9419), .A2(n9591), .ZN(n9026) );
  INV_X1 U11473 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9024) );
  OR2_X1 U11474 ( .A1(n9036), .A2(n9024), .ZN(n9025) );
  NOR2_X1 U11475 ( .A1(n9525), .A2(n9029), .ZN(n9030) );
  XNOR2_X1 U11476 ( .A(n9030), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n14305) );
  MUX2_X1 U11477 ( .A(n7224), .B(n14305), .S(n9584), .Z(n10601) );
  NAND2_X1 U11478 ( .A1(n10083), .A2(n9842), .ZN(n9031) );
  NAND2_X1 U11479 ( .A1(n13789), .A2(n10601), .ZN(n9480) );
  INV_X1 U11480 ( .A(n10083), .ZN(n9032) );
  INV_X1 U11481 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10149) );
  INV_X1 U11482 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9034) );
  OR2_X1 U11483 ( .A1(n9419), .A2(n9034), .ZN(n9038) );
  INV_X1 U11484 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9035) );
  NAND2_X1 U11485 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9039) );
  NAND2_X1 U11486 ( .A1(n9040), .A2(n10026), .ZN(n9044) );
  NAND2_X1 U11487 ( .A1(n9433), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9050) );
  INV_X1 U11488 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n13798) );
  OR2_X1 U11489 ( .A1(n6398), .A2(n13798), .ZN(n9049) );
  INV_X1 U11490 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9045) );
  OR2_X1 U11491 ( .A1(n9419), .A2(n9045), .ZN(n9048) );
  INV_X1 U11492 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9046) );
  NOR2_X1 U11493 ( .A1(n9544), .A2(n9440), .ZN(n9055) );
  OAI22_X1 U11494 ( .A1(n9217), .A2(n9543), .B1(n9584), .B2(n13801), .ZN(n9054) );
  OR2_X1 U11495 ( .A1(n9055), .A2(n9054), .ZN(n10631) );
  NAND2_X1 U11496 ( .A1(n10260), .A2(n10631), .ZN(n10085) );
  INV_X1 U11497 ( .A(n10631), .ZN(n14640) );
  NAND2_X1 U11498 ( .A1(n13788), .A2(n14640), .ZN(n9056) );
  MUX2_X1 U11499 ( .A(n10085), .B(n9056), .S(n9448), .Z(n9067) );
  NAND2_X1 U11500 ( .A1(n9522), .A2(n9454), .ZN(n9062) );
  NAND2_X1 U11501 ( .A1(n9057), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9058) );
  MUX2_X1 U11502 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9058), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n9060) );
  AND2_X1 U11503 ( .A1(n9060), .A2(n9081), .ZN(n13821) );
  AOI22_X1 U11504 ( .A1(n9277), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n9276), .B2(
        n13821), .ZN(n9061) );
  INV_X1 U11505 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n9688) );
  OR2_X1 U11506 ( .A1(n9428), .A2(n9688), .ZN(n9065) );
  INV_X1 U11507 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9702) );
  OR2_X1 U11508 ( .A1(n9419), .A2(n9702), .ZN(n9064) );
  OR2_X1 U11509 ( .A1(n6398), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9063) );
  NAND2_X1 U11510 ( .A1(n6936), .A2(n13787), .ZN(n9068) );
  NAND2_X1 U11511 ( .A1(n10636), .A2(n10331), .ZN(n10514) );
  NAND2_X1 U11512 ( .A1(n9537), .A2(n9454), .ZN(n9072) );
  NAND2_X1 U11513 ( .A1(n9081), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9070) );
  XNOR2_X1 U11514 ( .A(n9070), .B(P1_IR_REG_4__SCAN_IN), .ZN(n13828) );
  AOI22_X1 U11515 ( .A1(n9277), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n9276), .B2(
        n13828), .ZN(n9071) );
  AND2_X2 U11516 ( .A1(n9072), .A2(n9071), .ZN(n14646) );
  NAND2_X1 U11517 ( .A1(n9096), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9077) );
  OR2_X1 U11518 ( .A1(n9428), .A2(n15240), .ZN(n9076) );
  OAI21_X1 U11519 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n9085), .ZN(n10614) );
  OR2_X1 U11520 ( .A1(n6399), .A2(n10614), .ZN(n9075) );
  INV_X1 U11521 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9073) );
  OR2_X1 U11522 ( .A1(n9036), .A2(n9073), .ZN(n9074) );
  MUX2_X1 U11523 ( .A(n14646), .B(n10612), .S(n9448), .Z(n9079) );
  INV_X1 U11524 ( .A(n10612), .ZN(n13786) );
  MUX2_X1 U11525 ( .A(n13786), .B(n10617), .S(n9448), .Z(n9078) );
  OR2_X1 U11526 ( .A1(n9549), .A2(n9440), .ZN(n9084) );
  NOR2_X1 U11527 ( .A1(n9081), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n9102) );
  OR2_X1 U11528 ( .A1(n9102), .A2(n9227), .ZN(n9082) );
  XNOR2_X1 U11529 ( .A(n9082), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9705) );
  AOI22_X1 U11530 ( .A1(n9277), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n9276), .B2(
        n9705), .ZN(n9083) );
  NAND2_X1 U11531 ( .A1(n9434), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9090) );
  INV_X1 U11532 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10847) );
  OR2_X1 U11533 ( .A1(n9428), .A2(n10847), .ZN(n9089) );
  AND2_X1 U11534 ( .A1(n9085), .A2(n9723), .ZN(n9086) );
  OR2_X1 U11535 ( .A1(n9086), .A2(n9094), .ZN(n11002) );
  OR2_X1 U11536 ( .A1(n6398), .A2(n11002), .ZN(n9088) );
  INV_X1 U11537 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9704) );
  OR2_X1 U11538 ( .A1(n6400), .A2(n9704), .ZN(n9087) );
  NAND4_X1 U11539 ( .A1(n9090), .A2(n9089), .A3(n9088), .A4(n9087), .ZN(n13785) );
  MUX2_X1 U11540 ( .A(n11004), .B(n13785), .S(n9459), .Z(n9093) );
  MUX2_X1 U11541 ( .A(n13785), .B(n11004), .S(n9459), .Z(n9091) );
  NAND2_X1 U11542 ( .A1(n9434), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n9100) );
  INV_X1 U11543 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10942) );
  OR2_X1 U11544 ( .A1(n9428), .A2(n10942), .ZN(n9099) );
  OR2_X1 U11545 ( .A1(n9094), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9095) );
  NAND2_X1 U11546 ( .A1(n9112), .A2(n9095), .ZN(n10945) );
  OR2_X1 U11547 ( .A1(n6398), .A2(n10945), .ZN(n9098) );
  INV_X1 U11548 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9706) );
  OR2_X1 U11549 ( .A1(n9438), .A2(n9706), .ZN(n9097) );
  NAND4_X1 U11550 ( .A1(n9100), .A2(n9099), .A3(n9098), .A4(n9097), .ZN(n13784) );
  OR2_X1 U11551 ( .A1(n9575), .A2(n9440), .ZN(n9105) );
  NAND2_X1 U11552 ( .A1(n9102), .A2(n9101), .ZN(n9118) );
  NAND2_X1 U11553 ( .A1(n9118), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9103) );
  XNOR2_X1 U11554 ( .A(n9103), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9707) );
  AOI22_X1 U11555 ( .A1(n9277), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n9276), .B2(
        n9707), .ZN(n9104) );
  MUX2_X1 U11556 ( .A(n13784), .B(n14652), .S(n9459), .Z(n9108) );
  MUX2_X1 U11557 ( .A(n14652), .B(n13784), .S(n9459), .Z(n9106) );
  NAND2_X1 U11558 ( .A1(n9107), .A2(n9106), .ZN(n9110) );
  NAND2_X1 U11559 ( .A1(n9434), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n9117) );
  INV_X1 U11560 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10924) );
  OR2_X1 U11561 ( .A1(n9428), .A2(n10924), .ZN(n9116) );
  NAND2_X1 U11562 ( .A1(n9112), .A2(n9111), .ZN(n9113) );
  NAND2_X1 U11563 ( .A1(n9136), .A2(n9113), .ZN(n11174) );
  OR2_X1 U11564 ( .A1(n6399), .A2(n11174), .ZN(n9115) );
  INV_X1 U11565 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9708) );
  OR2_X1 U11566 ( .A1(n9438), .A2(n9708), .ZN(n9114) );
  NAND4_X1 U11567 ( .A1(n9117), .A2(n9116), .A3(n9115), .A4(n9114), .ZN(n13783) );
  NAND2_X1 U11568 ( .A1(n9127), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9119) );
  XNOR2_X1 U11569 ( .A(n9119), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9709) );
  AOI22_X1 U11570 ( .A1(n9277), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n9276), .B2(
        n9709), .ZN(n9120) );
  MUX2_X1 U11571 ( .A(n13783), .B(n11178), .S(n9448), .Z(n9122) );
  MUX2_X1 U11572 ( .A(n13783), .B(n11178), .S(n9459), .Z(n9121) );
  NAND2_X1 U11573 ( .A1(n9434), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n9126) );
  INV_X1 U11574 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9783) );
  OR2_X1 U11575 ( .A1(n9428), .A2(n9783), .ZN(n9125) );
  INV_X1 U11576 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n9135) );
  XNOR2_X1 U11577 ( .A(n9136), .B(n9135), .ZN(n10824) );
  OR2_X1 U11578 ( .A1(n6399), .A2(n10824), .ZN(n9124) );
  INV_X1 U11579 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9710) );
  OR2_X1 U11580 ( .A1(n9438), .A2(n9710), .ZN(n9123) );
  NAND4_X1 U11581 ( .A1(n9126), .A2(n9125), .A3(n9124), .A4(n9123), .ZN(n13782) );
  NAND2_X1 U11582 ( .A1(n9599), .A2(n9454), .ZN(n9130) );
  NAND2_X1 U11583 ( .A1(n9142), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9128) );
  XNOR2_X1 U11584 ( .A(n9128), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9780) );
  AOI22_X1 U11585 ( .A1(n9277), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n9276), .B2(
        n9780), .ZN(n9129) );
  MUX2_X1 U11586 ( .A(n13782), .B(n11348), .S(n9459), .Z(n9133) );
  MUX2_X1 U11587 ( .A(n13782), .B(n11348), .S(n9448), .Z(n9131) );
  NAND2_X1 U11588 ( .A1(n9434), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n9141) );
  INV_X1 U11589 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n11026) );
  OR2_X1 U11590 ( .A1(n9428), .A2(n11026), .ZN(n9140) );
  INV_X1 U11591 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n9134) );
  OAI21_X1 U11592 ( .B1(n9136), .B2(n9135), .A(n9134), .ZN(n9137) );
  NAND2_X1 U11593 ( .A1(n9137), .A2(n9152), .ZN(n11308) );
  OR2_X1 U11594 ( .A1(n6399), .A2(n11308), .ZN(n9139) );
  INV_X1 U11595 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9778) );
  OR2_X1 U11596 ( .A1(n9438), .A2(n9778), .ZN(n9138) );
  NAND4_X1 U11597 ( .A1(n9141), .A2(n9140), .A3(n9139), .A4(n9138), .ZN(n13781) );
  NOR2_X1 U11598 ( .A1(n9145), .A2(n9227), .ZN(n9143) );
  MUX2_X1 U11599 ( .A(n9227), .B(n9143), .S(P1_IR_REG_9__SCAN_IN), .Z(n9147)
         );
  INV_X1 U11600 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9144) );
  NAND2_X1 U11601 ( .A1(n9145), .A2(n9144), .ZN(n9179) );
  INV_X1 U11602 ( .A(n9179), .ZN(n9146) );
  NOR2_X1 U11603 ( .A1(n9147), .A2(n9146), .ZN(n9966) );
  INV_X1 U11604 ( .A(n9217), .ZN(n9213) );
  AOI22_X1 U11605 ( .A1(n9966), .A2(n9276), .B1(n9213), .B2(
        P2_DATAO_REG_9__SCAN_IN), .ZN(n9148) );
  MUX2_X1 U11606 ( .A(n13781), .B(n11312), .S(n9448), .Z(n9151) );
  MUX2_X1 U11607 ( .A(n13781), .B(n11312), .S(n9459), .Z(n9150) );
  NAND2_X1 U11608 ( .A1(n9096), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9160) );
  INV_X1 U11609 ( .A(n9173), .ZN(n9154) );
  NAND2_X1 U11610 ( .A1(n9152), .A2(n11408), .ZN(n9153) );
  NAND2_X1 U11611 ( .A1(n9154), .A2(n9153), .ZN(n14637) );
  OR2_X1 U11612 ( .A1(n6398), .A2(n14637), .ZN(n9159) );
  INV_X1 U11613 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n9155) );
  OR2_X1 U11614 ( .A1(n9428), .A2(n9155), .ZN(n9158) );
  INV_X1 U11615 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9156) );
  OR2_X1 U11616 ( .A1(n9036), .A2(n9156), .ZN(n9157) );
  NAND4_X1 U11617 ( .A1(n9160), .A2(n9159), .A3(n9158), .A4(n9157), .ZN(n13780) );
  NAND2_X1 U11618 ( .A1(n9618), .A2(n9454), .ZN(n9163) );
  NAND2_X1 U11619 ( .A1(n9179), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9161) );
  XNOR2_X1 U11620 ( .A(n9161), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10063) );
  AOI22_X1 U11621 ( .A1(n10063), .A2(n9276), .B1(n9213), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n9162) );
  MUX2_X1 U11622 ( .A(n13780), .B(n14623), .S(n9459), .Z(n9167) );
  MUX2_X1 U11623 ( .A(n13780), .B(n14623), .S(n9448), .Z(n9164) );
  NAND2_X1 U11624 ( .A1(n9165), .A2(n9164), .ZN(n9171) );
  INV_X1 U11625 ( .A(n9166), .ZN(n9169) );
  INV_X1 U11626 ( .A(n9167), .ZN(n9168) );
  NAND2_X1 U11627 ( .A1(n9169), .A2(n9168), .ZN(n9170) );
  NAND2_X1 U11628 ( .A1(n9434), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n9178) );
  INV_X1 U11629 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9172) );
  OR2_X1 U11630 ( .A1(n9428), .A2(n9172), .ZN(n9177) );
  OR2_X1 U11631 ( .A1(n9173), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9174) );
  NAND2_X1 U11632 ( .A1(n9185), .A2(n9174), .ZN(n11690) );
  OR2_X1 U11633 ( .A1(n6399), .A2(n11690), .ZN(n9176) );
  INV_X1 U11634 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10064) );
  OR2_X1 U11635 ( .A1(n9438), .A2(n10064), .ZN(n9175) );
  NAND4_X1 U11636 ( .A1(n9178), .A2(n9177), .A3(n9176), .A4(n9175), .ZN(n13779) );
  NAND2_X1 U11637 ( .A1(n9718), .A2(n9454), .ZN(n9182) );
  NAND2_X1 U11638 ( .A1(n9192), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9180) );
  XNOR2_X1 U11639 ( .A(n9180), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10277) );
  AOI22_X1 U11640 ( .A1(n10277), .A2(n9276), .B1(n9213), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n9181) );
  MUX2_X1 U11641 ( .A(n13779), .B(n11692), .S(n9448), .Z(n9184) );
  MUX2_X1 U11642 ( .A(n13779), .B(n11692), .S(n9459), .Z(n9183) );
  NAND2_X1 U11643 ( .A1(n9434), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n9191) );
  INV_X1 U11644 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11326) );
  OR2_X1 U11645 ( .A1(n9428), .A2(n11326), .ZN(n9190) );
  NAND2_X1 U11646 ( .A1(n9185), .A2(n10281), .ZN(n9186) );
  NAND2_X1 U11647 ( .A1(n9200), .A2(n9186), .ZN(n13665) );
  OR2_X1 U11648 ( .A1(n6398), .A2(n13665), .ZN(n9189) );
  INV_X1 U11649 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9187) );
  OR2_X1 U11650 ( .A1(n9438), .A2(n9187), .ZN(n9188) );
  NAND4_X1 U11651 ( .A1(n9191), .A2(n9190), .A3(n9189), .A4(n9188), .ZN(n13778) );
  NAND2_X1 U11652 ( .A1(n9891), .A2(n9454), .ZN(n9195) );
  OR2_X1 U11653 ( .A1(n9208), .A2(n9227), .ZN(n9193) );
  XNOR2_X1 U11654 ( .A(n9193), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10459) );
  AOI22_X1 U11655 ( .A1(n10459), .A2(n9276), .B1(n9213), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n9194) );
  MUX2_X1 U11656 ( .A(n13778), .B(n13661), .S(n9459), .Z(n9197) );
  MUX2_X1 U11657 ( .A(n13778), .B(n13661), .S(n9448), .Z(n9196) );
  INV_X1 U11658 ( .A(n9197), .ZN(n9198) );
  NAND2_X1 U11659 ( .A1(n9434), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n9206) );
  INV_X1 U11660 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11284) );
  OR2_X1 U11661 ( .A1(n9428), .A2(n11284), .ZN(n9205) );
  INV_X1 U11662 ( .A(n9220), .ZN(n9202) );
  NAND2_X1 U11663 ( .A1(n9200), .A2(n9199), .ZN(n9201) );
  NAND2_X1 U11664 ( .A1(n9202), .A2(n9201), .ZN(n13727) );
  OR2_X1 U11665 ( .A1(n6398), .A2(n13727), .ZN(n9204) );
  INV_X1 U11666 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10460) );
  OR2_X1 U11667 ( .A1(n6400), .A2(n10460), .ZN(n9203) );
  NAND4_X1 U11668 ( .A1(n9206), .A2(n9205), .A3(n9204), .A4(n9203), .ZN(n13777) );
  INV_X1 U11669 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9207) );
  NAND2_X1 U11670 ( .A1(n9208), .A2(n9207), .ZN(n9209) );
  NAND2_X1 U11671 ( .A1(n9209), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9211) );
  INV_X1 U11672 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9210) );
  NAND2_X1 U11673 ( .A1(n9211), .A2(n9210), .ZN(n9215) );
  OR2_X1 U11674 ( .A1(n9211), .A2(n9210), .ZN(n9212) );
  AOI22_X1 U11675 ( .A1(n10682), .A2(n9276), .B1(n9213), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n9214) );
  MUX2_X1 U11676 ( .A(n13777), .B(n14562), .S(n9448), .Z(n9243) );
  NAND2_X1 U11677 ( .A1(n10344), .A2(n9454), .ZN(n9219) );
  NAND2_X1 U11678 ( .A1(n9215), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9216) );
  XNOR2_X1 U11679 ( .A(n9216), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11438) );
  AOI22_X1 U11680 ( .A1(n11438), .A2(n9276), .B1(n9213), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n9218) );
  NAND2_X1 U11681 ( .A1(n9434), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n9225) );
  OR2_X1 U11682 ( .A1(n9220), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9221) );
  NAND2_X1 U11683 ( .A1(n9232), .A2(n9221), .ZN(n13632) );
  OR2_X1 U11684 ( .A1(n13632), .A2(n6399), .ZN(n9224) );
  INV_X1 U11685 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11624) );
  OR2_X1 U11686 ( .A1(n9428), .A2(n11624), .ZN(n9223) );
  INV_X1 U11687 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10680) );
  OR2_X1 U11688 ( .A1(n9438), .A2(n10680), .ZN(n9222) );
  OR2_X1 U11689 ( .A1(n13634), .A2(n13764), .ZN(n11722) );
  NAND2_X1 U11690 ( .A1(n13634), .A2(n13764), .ZN(n11725) );
  NAND2_X1 U11691 ( .A1(n10386), .A2(n9454), .ZN(n9230) );
  OR2_X1 U11692 ( .A1(n9500), .A2(n9227), .ZN(n9228) );
  XNOR2_X1 U11693 ( .A(n9228), .B(P1_IR_REG_15__SCAN_IN), .ZN(n11442) );
  AOI22_X1 U11694 ( .A1(n9277), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n9276), 
        .B2(n11442), .ZN(n9229) );
  NAND2_X1 U11695 ( .A1(n9232), .A2(n9231), .ZN(n9233) );
  AND2_X1 U11696 ( .A1(n9234), .A2(n9233), .ZN(n11734) );
  NAND2_X1 U11697 ( .A1(n11734), .A2(n9282), .ZN(n9239) );
  INV_X1 U11698 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n11735) );
  OR2_X1 U11699 ( .A1(n9428), .A2(n11735), .ZN(n9238) );
  INV_X1 U11700 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9235) );
  OR2_X1 U11701 ( .A1(n9036), .A2(n9235), .ZN(n9237) );
  INV_X1 U11702 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14594) );
  OR2_X1 U11703 ( .A1(n6400), .A2(n14594), .ZN(n9236) );
  NAND2_X1 U11704 ( .A1(n9241), .A2(n9448), .ZN(n9251) );
  INV_X1 U11705 ( .A(n9242), .ZN(n9248) );
  INV_X1 U11706 ( .A(n9243), .ZN(n9244) );
  AND3_X1 U11707 ( .A1(n11553), .A2(n13908), .A3(n9244), .ZN(n9247) );
  INV_X1 U11708 ( .A(n13686), .ZN(n14134) );
  AOI21_X1 U11709 ( .B1(n11725), .B2(n14134), .A(n9448), .ZN(n9246) );
  OAI21_X1 U11710 ( .B1(n14134), .B2(n11725), .A(n11906), .ZN(n9245) );
  NAND2_X1 U11711 ( .A1(n9249), .A2(n7608), .ZN(n9250) );
  NAND2_X1 U11712 ( .A1(n13887), .A2(n13686), .ZN(n9479) );
  NAND2_X1 U11713 ( .A1(n9263), .A2(n14136), .ZN(n9252) );
  INV_X1 U11714 ( .A(n13889), .ZN(n13910) );
  NAND2_X1 U11715 ( .A1(n13910), .A2(n9448), .ZN(n9259) );
  AOI21_X1 U11716 ( .B1(n9252), .B2(n9259), .A(n14242), .ZN(n9257) );
  INV_X1 U11717 ( .A(n14136), .ZN(n13892) );
  NAND2_X1 U11718 ( .A1(n9263), .A2(n13892), .ZN(n9254) );
  AOI21_X1 U11719 ( .B1(n9254), .B2(n9253), .A(n9486), .ZN(n9256) );
  OAI22_X1 U11720 ( .A1(n14132), .A2(n9255), .B1(n14136), .B2(n9259), .ZN(
        n9262) );
  OR3_X1 U11721 ( .A1(n9257), .A2(n9256), .A3(n9262), .ZN(n9258) );
  INV_X1 U11722 ( .A(n9259), .ZN(n9260) );
  NAND2_X1 U11723 ( .A1(n9263), .A2(n9260), .ZN(n9261) );
  OAI21_X1 U11724 ( .B1(n9459), .B2(n14136), .A(n9261), .ZN(n9264) );
  AOI22_X1 U11725 ( .A1(n9264), .A2(n9486), .B1(n9263), .B2(n9262), .ZN(n9265)
         );
  NAND2_X1 U11726 ( .A1(n10760), .A2(n9454), .ZN(n9269) );
  NAND2_X1 U11727 ( .A1(n6559), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9267) );
  XNOR2_X1 U11728 ( .A(n9267), .B(P1_IR_REG_18__SCAN_IN), .ZN(n13865) );
  AOI22_X1 U11729 ( .A1(n9277), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9276), 
        .B2(n13865), .ZN(n9268) );
  AND2_X1 U11730 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_17__SCAN_IN), 
        .ZN(n9270) );
  AOI21_X1 U11731 ( .B1(n9271), .B2(P1_REG3_REG_17__SCAN_IN), .A(
        P1_REG3_REG_18__SCAN_IN), .ZN(n9272) );
  OR2_X1 U11732 ( .A1(n9280), .A2(n9272), .ZN(n14107) );
  AOI22_X1 U11733 ( .A1(n9433), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9434), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n9274) );
  INV_X1 U11734 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n13848) );
  OR2_X1 U11735 ( .A1(n9438), .A2(n13848), .ZN(n9273) );
  OAI211_X1 U11736 ( .C1(n14107), .C2(n6398), .A(n9274), .B(n9273), .ZN(n13913) );
  OR2_X1 U11737 ( .A1(n14237), .A2(n13913), .ZN(n13894) );
  INV_X1 U11738 ( .A(n13913), .ZN(n14079) );
  MUX2_X1 U11739 ( .A(n14079), .B(n14110), .S(n9459), .Z(n9275) );
  NAND2_X1 U11740 ( .A1(n10992), .A2(n9454), .ZN(n9279) );
  AOI22_X1 U11741 ( .A1(n9277), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14008), 
        .B2(n9276), .ZN(n9278) );
  OR2_X1 U11742 ( .A1(n9280), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9281) );
  AND2_X1 U11743 ( .A1(n9293), .A2(n9281), .ZN(n14090) );
  NAND2_X1 U11744 ( .A1(n14090), .A2(n9282), .ZN(n9287) );
  INV_X1 U11745 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n13862) );
  NAND2_X1 U11746 ( .A1(n9433), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n9284) );
  NAND2_X1 U11747 ( .A1(n9434), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n9283) );
  OAI211_X1 U11748 ( .C1(n9438), .C2(n13862), .A(n9284), .B(n9283), .ZN(n9285)
         );
  INV_X1 U11749 ( .A(n9285), .ZN(n9286) );
  OR2_X1 U11750 ( .A1(n14086), .A2(n14103), .ZN(n9291) );
  NAND2_X1 U11751 ( .A1(n14086), .A2(n14103), .ZN(n13915) );
  AND2_X1 U11752 ( .A1(n14237), .A2(n13913), .ZN(n13895) );
  NAND2_X1 U11753 ( .A1(n9288), .A2(n13895), .ZN(n9289) );
  MUX2_X1 U11754 ( .A(n13915), .B(n9291), .S(n9448), .Z(n9292) );
  INV_X1 U11755 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13717) );
  NAND2_X1 U11756 ( .A1(n9293), .A2(n13717), .ZN(n9294) );
  NAND2_X1 U11757 ( .A1(n9306), .A2(n9294), .ZN(n14056) );
  OR2_X1 U11758 ( .A1(n14056), .A2(n6398), .ZN(n9299) );
  INV_X1 U11759 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n15155) );
  NAND2_X1 U11760 ( .A1(n9433), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n9296) );
  NAND2_X1 U11761 ( .A1(n9096), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n9295) );
  OAI211_X1 U11762 ( .C1(n9036), .C2(n15155), .A(n9296), .B(n9295), .ZN(n9297)
         );
  INV_X1 U11763 ( .A(n9297), .ZN(n9298) );
  NAND2_X1 U11764 ( .A1(n11331), .A2(n9454), .ZN(n9301) );
  NAND2_X1 U11765 ( .A1(n9213), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9300) );
  MUX2_X1 U11766 ( .A(n14080), .B(n14218), .S(n9448), .Z(n9303) );
  MUX2_X1 U11767 ( .A(n13916), .B(n13899), .S(n9459), .Z(n9302) );
  NAND2_X1 U11768 ( .A1(n9304), .A2(n9303), .ZN(n9305) );
  INV_X1 U11769 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n13656) );
  AND2_X1 U11770 ( .A1(n9306), .A2(n13656), .ZN(n9307) );
  OR2_X1 U11771 ( .A1(n9316), .A2(n9307), .ZN(n14050) );
  INV_X1 U11772 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n15190) );
  NAND2_X1 U11773 ( .A1(n9434), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n9309) );
  NAND2_X1 U11774 ( .A1(n9433), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9308) );
  OAI211_X1 U11775 ( .C1(n15190), .C2(n6400), .A(n9309), .B(n9308), .ZN(n9310)
         );
  INV_X1 U11776 ( .A(n9310), .ZN(n9311) );
  NAND2_X1 U11777 ( .A1(n11395), .A2(n9454), .ZN(n9313) );
  NAND2_X1 U11778 ( .A1(n9213), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9312) );
  MUX2_X1 U11779 ( .A(n14062), .B(n14212), .S(n9459), .Z(n9315) );
  MUX2_X1 U11780 ( .A(n14062), .B(n14212), .S(n9448), .Z(n9314) );
  OR2_X1 U11781 ( .A1(n9316), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9317) );
  NAND2_X1 U11782 ( .A1(n9316), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9330) );
  NAND2_X1 U11783 ( .A1(n9317), .A2(n9330), .ZN(n14030) );
  OR2_X1 U11784 ( .A1(n14030), .A2(n6399), .ZN(n9323) );
  INV_X1 U11785 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9320) );
  NAND2_X1 U11786 ( .A1(n9434), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n9319) );
  NAND2_X1 U11787 ( .A1(n9433), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9318) );
  OAI211_X1 U11788 ( .C1(n9320), .C2(n9438), .A(n9319), .B(n9318), .ZN(n9321)
         );
  INV_X1 U11789 ( .A(n9321), .ZN(n9322) );
  NAND2_X1 U11790 ( .A1(n9323), .A2(n9322), .ZN(n13775) );
  OR2_X1 U11791 ( .A1(n9324), .A2(n9533), .ZN(n9325) );
  XNOR2_X1 U11792 ( .A(n9325), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14303) );
  MUX2_X1 U11793 ( .A(n13775), .B(n14206), .S(n9448), .Z(n9328) );
  MUX2_X1 U11794 ( .A(n13775), .B(n14206), .S(n9459), .Z(n9326) );
  NAND2_X1 U11795 ( .A1(n9096), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n9336) );
  INV_X1 U11796 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9329) );
  OR2_X1 U11797 ( .A1(n9428), .A2(n9329), .ZN(n9335) );
  OAI21_X1 U11798 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n9331), .A(n9343), .ZN(
        n14018) );
  OR2_X1 U11799 ( .A1(n6399), .A2(n14018), .ZN(n9334) );
  INV_X1 U11800 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9332) );
  OR2_X1 U11801 ( .A1(n9036), .A2(n9332), .ZN(n9333) );
  NAND4_X1 U11802 ( .A1(n9336), .A2(n9335), .A3(n9334), .A4(n9333), .ZN(n14037) );
  NAND2_X1 U11803 ( .A1(n11767), .A2(n9454), .ZN(n9338) );
  NAND2_X1 U11804 ( .A1(n9213), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9337) );
  MUX2_X1 U11805 ( .A(n14037), .B(n14017), .S(n9459), .Z(n9340) );
  MUX2_X1 U11806 ( .A(n14037), .B(n14017), .S(n9448), .Z(n9339) );
  INV_X1 U11807 ( .A(n9340), .ZN(n9341) );
  NAND2_X1 U11808 ( .A1(n9434), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n9349) );
  INV_X1 U11809 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9342) );
  OR2_X1 U11810 ( .A1(n9428), .A2(n9342), .ZN(n9348) );
  OAI21_X1 U11811 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n9344), .A(n9357), .ZN(
        n13707) );
  OR2_X1 U11812 ( .A1(n6399), .A2(n13707), .ZN(n9347) );
  INV_X1 U11813 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9345) );
  OR2_X1 U11814 ( .A1(n6400), .A2(n9345), .ZN(n9346) );
  NAND4_X1 U11815 ( .A1(n9349), .A2(n9348), .A3(n9347), .A4(n9346), .ZN(n13774) );
  NAND2_X1 U11816 ( .A1(n13609), .A2(n9454), .ZN(n9351) );
  NAND2_X1 U11817 ( .A1(n9213), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n9350) );
  MUX2_X1 U11818 ( .A(n13774), .B(n14193), .S(n9448), .Z(n9354) );
  MUX2_X1 U11819 ( .A(n13774), .B(n14193), .S(n9023), .Z(n9352) );
  INV_X1 U11820 ( .A(n9354), .ZN(n9355) );
  NAND2_X1 U11821 ( .A1(n9434), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n9363) );
  INV_X1 U11822 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9356) );
  OR2_X1 U11823 ( .A1(n9428), .A2(n9356), .ZN(n9362) );
  OAI21_X1 U11824 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n9358), .A(n9377), .ZN(
        n13989) );
  OR2_X1 U11825 ( .A1(n6398), .A2(n13989), .ZN(n9361) );
  INV_X1 U11826 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9359) );
  OR2_X1 U11827 ( .A1(n6400), .A2(n9359), .ZN(n9360) );
  NAND4_X1 U11828 ( .A1(n9363), .A2(n9362), .A3(n9361), .A4(n9360), .ZN(n13773) );
  NAND2_X1 U11829 ( .A1(n13606), .A2(n9454), .ZN(n9365) );
  NAND2_X1 U11830 ( .A1(n9213), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9364) );
  MUX2_X1 U11831 ( .A(n13773), .B(n13922), .S(n9459), .Z(n9369) );
  MUX2_X1 U11832 ( .A(n13773), .B(n13922), .S(n9448), .Z(n9366) );
  NAND2_X1 U11833 ( .A1(n9367), .A2(n9366), .ZN(n9373) );
  INV_X1 U11834 ( .A(n9368), .ZN(n9371) );
  INV_X1 U11835 ( .A(n9369), .ZN(n9370) );
  NAND2_X1 U11836 ( .A1(n9371), .A2(n9370), .ZN(n9372) );
  NAND2_X1 U11837 ( .A1(n9433), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n9383) );
  INV_X1 U11838 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9374) );
  OR2_X1 U11839 ( .A1(n9036), .A2(n9374), .ZN(n9382) );
  INV_X1 U11840 ( .A(n9377), .ZN(n9375) );
  NAND2_X1 U11841 ( .A1(n9375), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n9390) );
  INV_X1 U11842 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9376) );
  NAND2_X1 U11843 ( .A1(n9377), .A2(n9376), .ZN(n9378) );
  NAND2_X1 U11844 ( .A1(n9390), .A2(n9378), .ZN(n13978) );
  OR2_X1 U11845 ( .A1(n6398), .A2(n13978), .ZN(n9381) );
  INV_X1 U11846 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9379) );
  OR2_X1 U11847 ( .A1(n9438), .A2(n9379), .ZN(n9380) );
  NAND4_X1 U11848 ( .A1(n9383), .A2(n9382), .A3(n9381), .A4(n9380), .ZN(n13962) );
  NAND2_X1 U11849 ( .A1(n13601), .A2(n9454), .ZN(n9385) );
  NAND2_X1 U11850 ( .A1(n9213), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9384) );
  MUX2_X1 U11851 ( .A(n13962), .B(n14179), .S(n9448), .Z(n9387) );
  MUX2_X1 U11852 ( .A(n13962), .B(n14179), .S(n9459), .Z(n9386) );
  NAND2_X1 U11853 ( .A1(n9433), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n9396) );
  INV_X1 U11854 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n15246) );
  OR2_X1 U11855 ( .A1(n9036), .A2(n15246), .ZN(n9395) );
  INV_X1 U11856 ( .A(n9390), .ZN(n9388) );
  NAND2_X1 U11857 ( .A1(n9388), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n9415) );
  INV_X1 U11858 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9389) );
  NAND2_X1 U11859 ( .A1(n9390), .A2(n9389), .ZN(n9391) );
  NAND2_X1 U11860 ( .A1(n9415), .A2(n9391), .ZN(n13965) );
  OR2_X1 U11861 ( .A1(n6399), .A2(n13965), .ZN(n9394) );
  INV_X1 U11862 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9392) );
  OR2_X1 U11863 ( .A1(n6400), .A2(n9392), .ZN(n9393) );
  NAND4_X1 U11864 ( .A1(n9396), .A2(n9395), .A3(n9394), .A4(n9393), .ZN(n13942) );
  NAND2_X1 U11865 ( .A1(n13598), .A2(n9454), .ZN(n9398) );
  NAND2_X1 U11866 ( .A1(n9213), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9397) );
  MUX2_X1 U11867 ( .A(n13942), .B(n14171), .S(n9459), .Z(n9402) );
  NAND2_X1 U11868 ( .A1(n9401), .A2(n9402), .ZN(n9400) );
  MUX2_X1 U11869 ( .A(n13942), .B(n14171), .S(n9448), .Z(n9399) );
  NAND2_X1 U11870 ( .A1(n9400), .A2(n9399), .ZN(n9403) );
  NAND2_X1 U11871 ( .A1(n9434), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n9408) );
  INV_X1 U11872 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n13951) );
  OR2_X1 U11873 ( .A1(n9428), .A2(n13951), .ZN(n9407) );
  INV_X1 U11874 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n11990) );
  XNOR2_X1 U11875 ( .A(n9415), .B(n11990), .ZN(n13950) );
  OR2_X1 U11876 ( .A1(n6398), .A2(n13950), .ZN(n9406) );
  INV_X1 U11877 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9404) );
  OR2_X1 U11878 ( .A1(n9438), .A2(n9404), .ZN(n9405) );
  NAND4_X1 U11879 ( .A1(n9408), .A2(n9407), .A3(n9406), .A4(n9405), .ZN(n13961) );
  NAND2_X1 U11880 ( .A1(n13595), .A2(n9454), .ZN(n9410) );
  NAND2_X1 U11881 ( .A1(n9213), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9409) );
  MUX2_X1 U11882 ( .A(n13961), .B(n14167), .S(n9448), .Z(n9412) );
  MUX2_X1 U11883 ( .A(n13961), .B(n14167), .S(n9023), .Z(n9411) );
  INV_X1 U11884 ( .A(n9412), .ZN(n9413) );
  NAND2_X1 U11885 ( .A1(n9434), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n9423) );
  INV_X1 U11886 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9414) );
  OR2_X1 U11887 ( .A1(n9428), .A2(n9414), .ZN(n9422) );
  INV_X1 U11888 ( .A(n9415), .ZN(n9416) );
  NAND2_X1 U11889 ( .A1(n9416), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n13934) );
  OR2_X1 U11890 ( .A1(n6398), .A2(n13934), .ZN(n9421) );
  INV_X1 U11891 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n9418) );
  OR2_X1 U11892 ( .A1(n6400), .A2(n9418), .ZN(n9420) );
  NAND4_X1 U11893 ( .A1(n9423), .A2(n9422), .A3(n9421), .A4(n9420), .ZN(n13941) );
  NAND2_X1 U11894 ( .A1(n13591), .A2(n9454), .ZN(n9425) );
  NAND2_X1 U11895 ( .A1(n9213), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n9424) );
  MUX2_X1 U11896 ( .A(n13941), .B(n13931), .S(n9023), .Z(n9450) );
  INV_X1 U11897 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9426) );
  OR2_X1 U11898 ( .A1(n9438), .A2(n9426), .ZN(n9432) );
  INV_X1 U11899 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9427) );
  OR2_X1 U11900 ( .A1(n9428), .A2(n9427), .ZN(n9431) );
  INV_X1 U11901 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9429) );
  OR2_X1 U11902 ( .A1(n9036), .A2(n9429), .ZN(n9430) );
  AND3_X1 U11903 ( .A1(n9432), .A2(n9431), .A3(n9430), .ZN(n9462) );
  INV_X1 U11904 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9437) );
  NAND2_X1 U11905 ( .A1(n9433), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9436) );
  NAND2_X1 U11906 ( .A1(n9434), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n9435) );
  OAI211_X1 U11907 ( .C1(n6400), .C2(n9437), .A(n9436), .B(n9435), .ZN(n13933)
         );
  OAI21_X1 U11908 ( .B1(n13879), .B2(n11354), .A(n13933), .ZN(n9439) );
  INV_X1 U11909 ( .A(n9439), .ZN(n9443) );
  NAND2_X1 U11910 ( .A1(n9213), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n9441) );
  MUX2_X1 U11911 ( .A(n9443), .B(n13882), .S(n9023), .Z(n9451) );
  INV_X1 U11912 ( .A(n9445), .ZN(n9446) );
  OAI22_X1 U11913 ( .A1(n9448), .A2(n9462), .B1(n9444), .B2(n9446), .ZN(n9447)
         );
  AOI22_X1 U11914 ( .A1(n13882), .A2(n9448), .B1(n13933), .B2(n9447), .ZN(
        n9452) );
  INV_X1 U11915 ( .A(n13941), .ZN(n11991) );
  INV_X1 U11916 ( .A(n13931), .ZN(n14159) );
  MUX2_X1 U11917 ( .A(n11991), .B(n14159), .S(n9448), .Z(n9449) );
  NAND2_X1 U11918 ( .A1(n9452), .A2(n9451), .ZN(n9453) );
  NAND2_X1 U11919 ( .A1(n13586), .A2(n9454), .ZN(n9456) );
  NAND2_X1 U11920 ( .A1(n9213), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n9455) );
  XNOR2_X1 U11921 ( .A(n9458), .B(n13879), .ZN(n9476) );
  OR2_X1 U11922 ( .A1(n9842), .A2(n9505), .ZN(n10570) );
  NAND2_X1 U11923 ( .A1(n9444), .A2(n14304), .ZN(n9853) );
  NAND2_X1 U11924 ( .A1(n11354), .A2(n9816), .ZN(n9819) );
  NAND2_X1 U11925 ( .A1(n9853), .A2(n9819), .ZN(n9457) );
  AND2_X1 U11926 ( .A1(n10570), .A2(n9457), .ZN(n9460) );
  NAND2_X1 U11927 ( .A1(n9458), .A2(n9459), .ZN(n9470) );
  INV_X1 U11928 ( .A(n9460), .ZN(n9463) );
  OR3_X1 U11929 ( .A1(n9470), .A2(n13879), .A3(n9463), .ZN(n9467) );
  NAND2_X1 U11930 ( .A1(n8999), .A2(n9461), .ZN(n9837) );
  AND2_X1 U11931 ( .A1(n9463), .A2(n9837), .ZN(n9469) );
  NAND4_X1 U11932 ( .A1(n9470), .A2(n9462), .A3(n9469), .A4(n9458), .ZN(n9466)
         );
  OR2_X1 U11933 ( .A1(n9458), .A2(n9023), .ZN(n9468) );
  XNOR2_X1 U11934 ( .A(n9468), .B(n9463), .ZN(n9464) );
  NAND4_X1 U11935 ( .A1(n9464), .A2(n14151), .A3(n9837), .A4(n13879), .ZN(
        n9465) );
  INV_X1 U11936 ( .A(n9468), .ZN(n9473) );
  INV_X1 U11937 ( .A(n9469), .ZN(n9472) );
  NOR2_X1 U11938 ( .A1(n9470), .A2(n13879), .ZN(n9471) );
  AOI211_X1 U11939 ( .C1(n9473), .C2(n13879), .A(n9472), .B(n9471), .ZN(n9474)
         );
  INV_X1 U11940 ( .A(n9476), .ZN(n9494) );
  XOR2_X1 U11941 ( .A(n13933), .B(n13882), .Z(n9493) );
  NAND2_X1 U11942 ( .A1(n14167), .A2(n13961), .ZN(n13906) );
  OAI21_X1 U11943 ( .B1(n14167), .B2(n13961), .A(n13906), .ZN(n13905) );
  XOR2_X1 U11944 ( .A(n13774), .B(n14193), .Z(n13901) );
  NAND2_X1 U11945 ( .A1(n14033), .A2(n13775), .ZN(n9477) );
  NAND2_X1 U11946 ( .A1(n13918), .A2(n9477), .ZN(n13917) );
  XNOR2_X1 U11947 ( .A(n14237), .B(n14079), .ZN(n14099) );
  INV_X1 U11948 ( .A(n11553), .ZN(n11547) );
  XNOR2_X1 U11949 ( .A(n14132), .B(n13910), .ZN(n14143) );
  XNOR2_X1 U11950 ( .A(n11692), .B(n13779), .ZN(n11224) );
  XNOR2_X1 U11951 ( .A(n11348), .B(n11309), .ZN(n10828) );
  XNOR2_X1 U11952 ( .A(n11178), .B(n11344), .ZN(n10810) );
  XNOR2_X1 U11953 ( .A(n14652), .B(n13784), .ZN(n10936) );
  INV_X1 U11954 ( .A(n10026), .ZN(n9481) );
  NAND2_X1 U11955 ( .A1(n10083), .A2(n9480), .ZN(n10604) );
  NOR4_X1 U11956 ( .A1(n10080), .A2(n10624), .A3(n9481), .A4(n10604), .ZN(
        n9482) );
  XNOR2_X1 U11957 ( .A(n11004), .B(n13785), .ZN(n10799) );
  XNOR2_X1 U11958 ( .A(n10617), .B(n13786), .ZN(n10584) );
  NAND4_X1 U11959 ( .A1(n10936), .A2(n9482), .A3(n10799), .A4(n10584), .ZN(
        n9483) );
  NOR4_X1 U11960 ( .A1(n11020), .A2(n10828), .A3(n10810), .A4(n9483), .ZN(
        n9484) );
  XNOR2_X1 U11961 ( .A(n13661), .B(n13778), .ZN(n11279) );
  XNOR2_X1 U11962 ( .A(n14623), .B(n13780), .ZN(n11215) );
  NAND4_X1 U11963 ( .A1(n11224), .A2(n9484), .A3(n11279), .A4(n11215), .ZN(
        n9485) );
  NOR4_X1 U11964 ( .A1(n11547), .A2(n11550), .A3(n14143), .A4(n9485), .ZN(
        n9487) );
  XNOR2_X1 U11965 ( .A(n9486), .B(n14136), .ZN(n14127) );
  NAND3_X1 U11966 ( .A1(n11731), .A2(n9487), .A3(n14127), .ZN(n9488) );
  NOR4_X1 U11967 ( .A1(n13917), .A2(n14099), .A3(n14084), .A4(n9488), .ZN(
        n9489) );
  XNOR2_X1 U11968 ( .A(n14017), .B(n14037), .ZN(n13920) );
  XNOR2_X1 U11969 ( .A(n14212), .B(n14062), .ZN(n13900) );
  XNOR2_X1 U11970 ( .A(n13899), .B(n13916), .ZN(n13898) );
  NAND4_X1 U11971 ( .A1(n9489), .A2(n13920), .A3(n13900), .A4(n13898), .ZN(
        n9490) );
  NOR3_X1 U11972 ( .A1(n13901), .A2(n13994), .A3(n9490), .ZN(n9491) );
  NAND4_X1 U11973 ( .A1(n13905), .A2(n9491), .A3(n13958), .A4(n13902), .ZN(
        n9492) );
  XOR2_X1 U11974 ( .A(n9495), .B(n14008), .Z(n9497) );
  INV_X1 U11975 ( .A(n9837), .ZN(n9496) );
  OAI21_X1 U11976 ( .B1(n8992), .B2(n9498), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9499) );
  MUX2_X1 U11977 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9499), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n9501) );
  NAND2_X1 U11978 ( .A1(n9501), .A2(n9509), .ZN(n9582) );
  OR2_X1 U11979 ( .A1(n9582), .A2(P1_U3086), .ZN(n11770) );
  INV_X1 U11980 ( .A(n11770), .ZN(n9502) );
  AND2_X1 U11981 ( .A1(n11354), .A2(n9505), .ZN(n9851) );
  OR2_X1 U11982 ( .A1(n9853), .A2(n9851), .ZN(n9808) );
  NAND2_X1 U11983 ( .A1(n9511), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9506) );
  MUX2_X1 U11984 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9506), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n9508) );
  NAND2_X1 U11985 ( .A1(n9509), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9510) );
  MUX2_X1 U11986 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9510), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n9512) );
  NAND2_X1 U11987 ( .A1(n9512), .A2(n9511), .ZN(n14301) );
  AND2_X1 U11988 ( .A1(n9841), .A2(n9582), .ZN(n9513) );
  NAND2_X1 U11989 ( .A1(n9808), .A2(n9513), .ZN(n9826) );
  INV_X1 U11990 ( .A(n13790), .ZN(n13878) );
  NAND2_X1 U11991 ( .A1(n13878), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14290) );
  OAI21_X1 U11992 ( .B1(n14304), .B2(n11770), .A(P1_B_REG_SCAN_IN), .ZN(n9514)
         );
  INV_X1 U11993 ( .A(n9514), .ZN(n9515) );
  NAND2_X1 U11994 ( .A1(n9517), .A2(n9516), .ZN(P1_U3242) );
  INV_X1 U11995 ( .A(n9532), .ZN(n9518) );
  OR2_X2 U11996 ( .A1(n9841), .A2(n9518), .ZN(n13793) );
  AND2_X1 U11997 ( .A1(n9533), .A2(P2_U3088), .ZN(n13594) );
  INV_X2 U11998 ( .A(n13594), .ZN(n13605) );
  INV_X1 U11999 ( .A(n9652), .ZN(n14703) );
  NOR2_X1 U12000 ( .A1(n9533), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13602) );
  INV_X2 U12001 ( .A(n13602), .ZN(n13614) );
  OAI222_X1 U12002 ( .A1(n13605), .A2(n9526), .B1(n14703), .B2(P2_U3088), .C1(
        n15142), .C2(n13614), .ZN(P2_U3326) );
  OAI222_X1 U12003 ( .A1(n13605), .A2(n9544), .B1(n6393), .B2(P2_U3088), .C1(
        n9521), .C2(n13614), .ZN(P2_U3325) );
  INV_X1 U12004 ( .A(n9522), .ZN(n9541) );
  INV_X1 U12005 ( .A(n13116), .ZN(n9524) );
  OAI222_X1 U12006 ( .A1(n13605), .A2(n9541), .B1(n9524), .B2(P2_U3088), .C1(
        n9523), .C2(n13614), .ZN(P2_U3324) );
  AND2_X1 U12007 ( .A1(n9533), .A2(P1_U3086), .ZN(n14288) );
  INV_X2 U12008 ( .A(n14288), .ZN(n14298) );
  NOR2_X1 U12009 ( .A1(n9533), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14280) );
  INV_X2 U12010 ( .A(n14280), .ZN(n14300) );
  OAI222_X1 U12011 ( .A1(n14298), .A2(n7399), .B1(n14300), .B2(n9526), .C1(
        P1_U3086), .C2(n7347), .ZN(P1_U3354) );
  AND2_X1 U12012 ( .A1(n14301), .A2(P1_B_REG_SCAN_IN), .ZN(n9529) );
  INV_X1 U12013 ( .A(n14301), .ZN(n9528) );
  INV_X1 U12014 ( .A(P1_B_REG_SCAN_IN), .ZN(n9527) );
  AOI22_X1 U12015 ( .A1(n14297), .A2(n9529), .B1(n9528), .B2(n9527), .ZN(n9530) );
  NAND2_X1 U12016 ( .A1(n9841), .A2(n9532), .ZN(n9831) );
  OR2_X1 U12017 ( .A1(n9814), .A2(n9831), .ZN(n15229) );
  INV_X1 U12018 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9811) );
  AND2_X1 U12019 ( .A1(n14294), .A2(n14297), .ZN(n9810) );
  AOI22_X1 U12020 ( .A1(n15229), .A2(n9811), .B1(n9532), .B2(n9810), .ZN(
        P1_U3446) );
  INV_X1 U12021 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9813) );
  AND2_X1 U12022 ( .A1(n14294), .A2(n14301), .ZN(n9812) );
  AOI22_X1 U12023 ( .A1(n15229), .A2(n9813), .B1(n9532), .B2(n9812), .ZN(
        P1_U3445) );
  NOR2_X1 U12024 ( .A1(n9533), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12961) );
  INV_X2 U12025 ( .A(n12961), .ZN(n14410) );
  OAI222_X1 U12026 ( .A1(n14919), .A2(P3_U3151), .B1(n14410), .B2(n9536), .C1(
        n9535), .C2(n12973), .ZN(P3_U3289) );
  INV_X1 U12027 ( .A(n9537), .ZN(n9546) );
  INV_X1 U12028 ( .A(n14739), .ZN(n9539) );
  OAI222_X1 U12029 ( .A1(n13605), .A2(n9546), .B1(n9539), .B2(P2_U3088), .C1(
        n9538), .C2(n13614), .ZN(P2_U3323) );
  INV_X1 U12030 ( .A(n13821), .ZN(n9542) );
  OAI222_X1 U12031 ( .A1(P1_U3086), .A2(n9542), .B1(n14300), .B2(n9541), .C1(
        n9540), .C2(n14298), .ZN(P1_U3352) );
  OAI222_X1 U12032 ( .A1(P1_U3086), .A2(n13801), .B1(n14300), .B2(n9544), .C1(
        n9543), .C2(n14298), .ZN(P1_U3353) );
  INV_X1 U12033 ( .A(n13828), .ZN(n9694) );
  OAI222_X1 U12034 ( .A1(P1_U3086), .A2(n9694), .B1(n14300), .B2(n9546), .C1(
        n9545), .C2(n14298), .ZN(P1_U3351) );
  OAI222_X1 U12035 ( .A1(n13605), .A2(n9549), .B1(n6617), .B2(P2_U3088), .C1(
        n9547), .C2(n13614), .ZN(P2_U3322) );
  INV_X1 U12036 ( .A(n9705), .ZN(n9725) );
  OAI222_X1 U12037 ( .A1(P1_U3086), .A2(n9725), .B1(n14300), .B2(n9549), .C1(
        n9548), .C2(n14298), .ZN(P1_U3350) );
  OAI222_X1 U12038 ( .A1(n14410), .A2(n9551), .B1(n12973), .B2(n9550), .C1(
        n11700), .C2(P3_U3151), .ZN(P3_U3284) );
  INV_X1 U12039 ( .A(n9661), .ZN(n9887) );
  OAI222_X1 U12040 ( .A1(n13605), .A2(n9575), .B1(n9887), .B2(P2_U3088), .C1(
        n9552), .C2(n13614), .ZN(P2_U3321) );
  INV_X1 U12041 ( .A(n9553), .ZN(n9555) );
  INV_X1 U12042 ( .A(SI_3_), .ZN(n9554) );
  OAI222_X1 U12043 ( .A1(n14410), .A2(n9555), .B1(n12973), .B2(n9554), .C1(
        n14863), .C2(P3_U3151), .ZN(P3_U3292) );
  INV_X1 U12044 ( .A(n9556), .ZN(n9558) );
  INV_X1 U12045 ( .A(SI_5_), .ZN(n9557) );
  OAI222_X1 U12046 ( .A1(n14410), .A2(n9558), .B1(n12973), .B2(n9557), .C1(
        n14900), .C2(P3_U3151), .ZN(P3_U3290) );
  INV_X1 U12047 ( .A(n9559), .ZN(n9561) );
  INV_X1 U12048 ( .A(SI_4_), .ZN(n9560) );
  OAI222_X1 U12049 ( .A1(n14410), .A2(n9561), .B1(n12973), .B2(n9560), .C1(
        n14880), .C2(P3_U3151), .ZN(P3_U3291) );
  INV_X1 U12050 ( .A(n9562), .ZN(n9564) );
  INV_X1 U12051 ( .A(SI_7_), .ZN(n9563) );
  INV_X1 U12052 ( .A(n11509), .ZN(n14939) );
  OAI222_X1 U12053 ( .A1(n14410), .A2(n9564), .B1(n12973), .B2(n9563), .C1(
        n14939), .C2(P3_U3151), .ZN(P3_U3288) );
  INV_X1 U12054 ( .A(SI_9_), .ZN(n9565) );
  OAI222_X1 U12055 ( .A1(n14410), .A2(n9566), .B1(n12973), .B2(n9565), .C1(
        n14978), .C2(P3_U3151), .ZN(P3_U3286) );
  OAI222_X1 U12056 ( .A1(n14410), .A2(n9568), .B1(n12973), .B2(n9567), .C1(
        n14957), .C2(P3_U3151), .ZN(P3_U3287) );
  INV_X1 U12057 ( .A(n9569), .ZN(n9571) );
  INV_X1 U12058 ( .A(SI_2_), .ZN(n9570) );
  OAI222_X1 U12059 ( .A1(n14410), .A2(n9571), .B1(n12973), .B2(n9570), .C1(
        n11463), .C2(P3_U3151), .ZN(P3_U3293) );
  OAI222_X1 U12060 ( .A1(P3_U3151), .A2(n6913), .B1(n12973), .B2(n9573), .C1(
        n14410), .C2(n9572), .ZN(P3_U3294) );
  INV_X1 U12061 ( .A(n9707), .ZN(n9924) );
  OAI222_X1 U12062 ( .A1(P1_U3086), .A2(n9924), .B1(n14300), .B2(n9575), .C1(
        n9574), .C2(n14298), .ZN(P1_U3349) );
  OAI222_X1 U12063 ( .A1(n14410), .A2(n9577), .B1(n12456), .B2(P3_U3151), .C1(
        n9576), .C2(n12973), .ZN(P3_U3283) );
  INV_X1 U12064 ( .A(n9899), .ZN(n9579) );
  OAI222_X1 U12065 ( .A1(n13605), .A2(n9581), .B1(n9579), .B2(P2_U3088), .C1(
        n9578), .C2(n13614), .ZN(P2_U3320) );
  INV_X1 U12066 ( .A(n9709), .ZN(n9958) );
  OAI222_X1 U12067 ( .A1(P1_U3086), .A2(n9958), .B1(n14300), .B2(n9581), .C1(
        n9580), .C2(n14298), .ZN(P1_U3348) );
  INV_X1 U12068 ( .A(n9582), .ZN(n9583) );
  OR2_X1 U12069 ( .A1(n9853), .A2(n9583), .ZN(n9585) );
  NAND2_X1 U12070 ( .A1(n9585), .A2(n9584), .ZN(n9586) );
  NAND2_X1 U12071 ( .A1(n9831), .A2(n11770), .ZN(n9587) );
  NAND2_X1 U12072 ( .A1(n9586), .A2(n9587), .ZN(n14607) );
  INV_X1 U12073 ( .A(n14607), .ZN(n13817) );
  NOR2_X1 U12074 ( .A1(n13817), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U12075 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9595) );
  INV_X1 U12076 ( .A(n9586), .ZN(n9588) );
  AND2_X1 U12077 ( .A1(n9588), .A2(n9587), .ZN(n9678) );
  INV_X1 U12078 ( .A(n13796), .ZN(n9822) );
  INV_X1 U12079 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9589) );
  NAND2_X1 U12080 ( .A1(n13878), .A2(n9589), .ZN(n9590) );
  NAND2_X1 U12081 ( .A1(n9822), .A2(n9590), .ZN(n13794) );
  AOI21_X1 U12082 ( .B1(n13790), .B2(n9591), .A(n13794), .ZN(n9592) );
  XNOR2_X1 U12083 ( .A(n9592), .B(n7224), .ZN(n9593) );
  AOI22_X1 U12084 ( .A1(n9678), .A2(n9593), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n9594) );
  OAI21_X1 U12085 ( .B1(n14607), .B2(n9595), .A(n9594), .ZN(P1_U3243) );
  INV_X1 U12086 ( .A(n12483), .ZN(n12476) );
  OAI222_X1 U12087 ( .A1(n14410), .A2(n9597), .B1(n12476), .B2(P3_U3151), .C1(
        n9596), .C2(n12973), .ZN(P3_U3282) );
  OAI222_X1 U12088 ( .A1(n13605), .A2(n9604), .B1(n9664), .B2(P2_U3088), .C1(
        n9598), .C2(n13614), .ZN(P2_U3318) );
  INV_X1 U12089 ( .A(n9599), .ZN(n9602) );
  OAI222_X1 U12090 ( .A1(n13614), .A2(n9600), .B1(n13605), .B2(n9602), .C1(
        P2_U3088), .C2(n6633), .ZN(P2_U3319) );
  INV_X1 U12091 ( .A(n9780), .ZN(n9784) );
  OAI222_X1 U12092 ( .A1(n9784), .A2(P1_U3086), .B1(n14300), .B2(n9602), .C1(
        n9601), .C2(n14298), .ZN(P1_U3347) );
  INV_X1 U12093 ( .A(n9966), .ZN(n9792) );
  OAI222_X1 U12094 ( .A1(P1_U3086), .A2(n9792), .B1(n14300), .B2(n9604), .C1(
        n9603), .C2(n14298), .ZN(P1_U3346) );
  NOR2_X2 U12095 ( .A1(n8892), .A2(n12957), .ZN(n9928) );
  INV_X1 U12096 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n9605) );
  NOR2_X1 U12097 ( .A1(n9928), .A2(n9605), .ZN(P3_U3249) );
  INV_X1 U12098 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n9606) );
  NOR2_X1 U12099 ( .A1(n9928), .A2(n9606), .ZN(P3_U3247) );
  INV_X1 U12100 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n9607) );
  NOR2_X1 U12101 ( .A1(n9928), .A2(n9607), .ZN(P3_U3251) );
  INV_X1 U12102 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n9608) );
  NOR2_X1 U12103 ( .A1(n9928), .A2(n9608), .ZN(P3_U3248) );
  INV_X1 U12104 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n9609) );
  NOR2_X1 U12105 ( .A1(n9928), .A2(n9609), .ZN(P3_U3259) );
  INV_X1 U12106 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n9610) );
  NOR2_X1 U12107 ( .A1(n9928), .A2(n9610), .ZN(P3_U3258) );
  INV_X1 U12108 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n9611) );
  NOR2_X1 U12109 ( .A1(n9928), .A2(n9611), .ZN(P3_U3252) );
  INV_X1 U12110 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n9612) );
  NOR2_X1 U12111 ( .A1(n9928), .A2(n9612), .ZN(P3_U3261) );
  INV_X1 U12112 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n9613) );
  NOR2_X1 U12113 ( .A1(n9928), .A2(n9613), .ZN(P3_U3253) );
  INV_X1 U12114 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n9614) );
  NOR2_X1 U12115 ( .A1(n9928), .A2(n9614), .ZN(P3_U3246) );
  INV_X1 U12116 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n9615) );
  NOR2_X1 U12117 ( .A1(n9928), .A2(n9615), .ZN(P3_U3250) );
  INV_X1 U12118 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n15170) );
  NOR2_X1 U12119 ( .A1(n9928), .A2(n15170), .ZN(P3_U3260) );
  OAI222_X1 U12120 ( .A1(n14410), .A2(n9617), .B1(n12973), .B2(n9616), .C1(
        n12495), .C2(P3_U3151), .ZN(P3_U3281) );
  INV_X1 U12121 ( .A(n10063), .ZN(n9973) );
  INV_X1 U12122 ( .A(n9618), .ZN(n9620) );
  OAI222_X1 U12123 ( .A1(n9973), .A2(P1_U3086), .B1(n14300), .B2(n9620), .C1(
        n9619), .C2(n14298), .ZN(P1_U3345) );
  INV_X1 U12124 ( .A(n10176), .ZN(n10017) );
  OAI222_X1 U12125 ( .A1(n13614), .A2(n9621), .B1(n13605), .B2(n9620), .C1(
        P2_U3088), .C2(n10017), .ZN(P2_U3317) );
  OAI222_X1 U12126 ( .A1(n14410), .A2(n9623), .B1(n12973), .B2(n9622), .C1(
        n12525), .C2(P3_U3151), .ZN(P3_U3280) );
  XNOR2_X1 U12127 ( .A(n9664), .B(P2_REG2_REG_9__SCAN_IN), .ZN(n9637) );
  INV_X1 U12128 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9624) );
  MUX2_X1 U12129 ( .A(n9624), .B(P2_REG2_REG_2__SCAN_IN), .S(n6393), .Z(n14725) );
  INV_X1 U12130 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n15247) );
  MUX2_X1 U12131 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n15247), .S(n9652), .Z(
        n14708) );
  AND2_X1 U12132 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n14707) );
  NAND2_X1 U12133 ( .A1(n14708), .A2(n14707), .ZN(n14706) );
  NAND2_X1 U12134 ( .A1(n9652), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9625) );
  NAND2_X1 U12135 ( .A1(n14706), .A2(n9625), .ZN(n14724) );
  NAND2_X1 U12136 ( .A1(n14725), .A2(n14724), .ZN(n14723) );
  INV_X1 U12137 ( .A(n6393), .ZN(n14726) );
  NAND2_X1 U12138 ( .A1(n14726), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n9626) );
  NAND2_X1 U12139 ( .A1(n14723), .A2(n9626), .ZN(n13118) );
  INV_X1 U12140 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9627) );
  MUX2_X1 U12141 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n9627), .S(n13116), .Z(
        n13119) );
  NAND2_X1 U12142 ( .A1(n13118), .A2(n13119), .ZN(n13117) );
  NAND2_X1 U12143 ( .A1(n13116), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9628) );
  NAND2_X1 U12144 ( .A1(n13117), .A2(n9628), .ZN(n14737) );
  INV_X1 U12145 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9629) );
  MUX2_X1 U12146 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n9629), .S(n14739), .Z(
        n14738) );
  NAND2_X1 U12147 ( .A1(n14737), .A2(n14738), .ZN(n14736) );
  NAND2_X1 U12148 ( .A1(n14739), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9630) );
  NAND2_X1 U12149 ( .A1(n14736), .A2(n9630), .ZN(n14749) );
  INV_X1 U12150 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n9631) );
  MUX2_X1 U12151 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n9631), .S(n9659), .Z(n14750) );
  AND2_X1 U12152 ( .A1(n14749), .A2(n14750), .ZN(n14747) );
  INV_X1 U12153 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n9632) );
  MUX2_X1 U12154 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n9632), .S(n9661), .Z(n9633)
         );
  INV_X1 U12155 ( .A(n9633), .ZN(n9881) );
  NOR2_X1 U12156 ( .A1(n9882), .A2(n9881), .ZN(n9880) );
  AOI21_X1 U12157 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n9661), .A(n9880), .ZN(
        n9895) );
  INV_X1 U12158 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9634) );
  MUX2_X1 U12159 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n9634), .S(n9899), .Z(n9635)
         );
  INV_X1 U12160 ( .A(n9635), .ZN(n9894) );
  NOR2_X1 U12161 ( .A1(n9895), .A2(n9894), .ZN(n9893) );
  XNOR2_X1 U12162 ( .A(n9663), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n9909) );
  NOR2_X1 U12163 ( .A1(n9910), .A2(n9909), .ZN(n9908) );
  NAND2_X1 U12164 ( .A1(n9636), .A2(n9637), .ZN(n10012) );
  OAI21_X1 U12165 ( .B1(n9637), .B2(n9636), .A(n10012), .ZN(n9649) );
  NAND2_X1 U12166 ( .A1(n9768), .A2(n9638), .ZN(n9639) );
  NAND2_X1 U12167 ( .A1(n9639), .A2(n7685), .ZN(n9640) );
  INV_X1 U12168 ( .A(n9646), .ZN(n9645) );
  NAND2_X1 U12169 ( .A1(n9642), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13596) );
  INV_X1 U12170 ( .A(n13596), .ZN(n9643) );
  AND2_X1 U12171 ( .A1(n9645), .A2(n9643), .ZN(n9668) );
  AND2_X1 U12172 ( .A1(n9645), .A2(n9764), .ZN(n14702) );
  NAND2_X1 U12173 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n10955) );
  AND2_X1 U12174 ( .A1(n9646), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14719) );
  NAND2_X1 U12175 ( .A1(n14719), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n9647) );
  OAI211_X1 U12176 ( .C1(n14774), .C2(n9664), .A(n10955), .B(n9647), .ZN(n9648) );
  AOI21_X1 U12177 ( .B1(n9649), .B2(n14770), .A(n9648), .ZN(n9671) );
  INV_X1 U12178 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10003) );
  MUX2_X1 U12179 ( .A(n10003), .B(P2_REG1_REG_2__SCAN_IN), .S(n6393), .Z(
        n14722) );
  INV_X1 U12180 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9987) );
  MUX2_X1 U12181 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n9987), .S(n9652), .Z(n14710) );
  AND2_X1 U12182 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n9651) );
  NAND2_X1 U12183 ( .A1(n14710), .A2(n9651), .ZN(n14711) );
  NAND2_X1 U12184 ( .A1(n9652), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9653) );
  NAND2_X1 U12185 ( .A1(n14711), .A2(n9653), .ZN(n14721) );
  NAND2_X1 U12186 ( .A1(n14722), .A2(n14721), .ZN(n14720) );
  NAND2_X1 U12187 ( .A1(n14726), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9654) );
  NAND2_X1 U12188 ( .A1(n14720), .A2(n9654), .ZN(n13113) );
  INV_X1 U12189 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9655) );
  MUX2_X1 U12190 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n9655), .S(n13116), .Z(
        n13114) );
  NAND2_X1 U12191 ( .A1(n13113), .A2(n13114), .ZN(n13112) );
  NAND2_X1 U12192 ( .A1(n13116), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9656) );
  NAND2_X1 U12193 ( .A1(n13112), .A2(n9656), .ZN(n14734) );
  INV_X1 U12194 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9657) );
  MUX2_X1 U12195 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n9657), .S(n14739), .Z(
        n14735) );
  NAND2_X1 U12196 ( .A1(n14734), .A2(n14735), .ZN(n14733) );
  NAND2_X1 U12197 ( .A1(n14739), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9658) );
  NAND2_X1 U12198 ( .A1(n14733), .A2(n9658), .ZN(n14752) );
  MUX2_X1 U12199 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6616), .S(n9659), .Z(n14751) );
  INV_X1 U12200 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9660) );
  MUX2_X1 U12201 ( .A(n9660), .B(P2_REG1_REG_6__SCAN_IN), .S(n9661), .Z(n9884)
         );
  INV_X1 U12202 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9662) );
  MUX2_X1 U12203 ( .A(n9662), .B(P2_REG1_REG_7__SCAN_IN), .S(n9899), .Z(n9897)
         );
  NOR2_X1 U12204 ( .A1(n9898), .A2(n9897), .ZN(n9896) );
  MUX2_X1 U12205 ( .A(n6632), .B(P2_REG1_REG_8__SCAN_IN), .S(n9663), .Z(n9906)
         );
  INV_X1 U12206 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9665) );
  MUX2_X1 U12207 ( .A(n9665), .B(P2_REG1_REG_9__SCAN_IN), .S(n9664), .Z(n9666)
         );
  OAI21_X1 U12208 ( .B1(n9667), .B2(n9666), .A(n10007), .ZN(n9669) );
  NAND2_X1 U12209 ( .A1(n9668), .A2(n13600), .ZN(n14791) );
  INV_X1 U12210 ( .A(n14791), .ZN(n14765) );
  NAND2_X1 U12211 ( .A1(n9669), .A2(n14765), .ZN(n9670) );
  NAND2_X1 U12212 ( .A1(n9671), .A2(n9670), .ZN(P2_U3223) );
  AND2_X1 U12213 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9673) );
  INV_X1 U12214 ( .A(n9673), .ZN(n13792) );
  MUX2_X1 U12215 ( .A(n9672), .B(P1_REG2_REG_1__SCAN_IN), .S(n9698), .Z(n9677)
         );
  INV_X1 U12216 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9672) );
  MUX2_X1 U12217 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n9672), .S(n9698), .Z(n9674)
         );
  NAND2_X1 U12218 ( .A1(n9674), .A2(n9673), .ZN(n13803) );
  INV_X1 U12219 ( .A(n13803), .ZN(n9676) );
  NAND2_X1 U12220 ( .A1(n9678), .A2(n13878), .ZN(n13869) );
  INV_X1 U12221 ( .A(n13869), .ZN(n9675) );
  AOI211_X1 U12222 ( .C1(n13792), .C2(n9677), .A(n9676), .B(n14600), .ZN(n9685) );
  NAND2_X1 U12223 ( .A1(n9678), .A2(n13796), .ZN(n14598) );
  MUX2_X1 U12224 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9034), .S(n9698), .Z(n9681)
         );
  AND2_X1 U12225 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9680) );
  INV_X1 U12226 ( .A(n9678), .ZN(n9679) );
  NOR2_X2 U12227 ( .A1(n9679), .A2(n13878), .ZN(n14604) );
  NAND2_X1 U12228 ( .A1(n9681), .A2(n9680), .ZN(n9700) );
  OAI211_X1 U12229 ( .C1(n9681), .C2(n9680), .A(n14604), .B(n9700), .ZN(n9683)
         );
  AOI22_X1 U12230 ( .A1(n13817), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9682) );
  OAI211_X1 U12231 ( .C1(n14598), .C2(n7347), .A(n9683), .B(n9682), .ZN(n9684)
         );
  OR2_X1 U12232 ( .A1(n9685), .A2(n9684), .ZN(P1_U3244) );
  OAI222_X1 U12233 ( .A1(n14410), .A2(n9687), .B1(n12550), .B2(P3_U3151), .C1(
        n9686), .C2(n12973), .ZN(P3_U3279) );
  MUX2_X1 U12234 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n9688), .S(n13821), .Z(n9693) );
  INV_X1 U12235 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9689) );
  MUX2_X1 U12236 ( .A(n9689), .B(P1_REG2_REG_2__SCAN_IN), .S(n13801), .Z(n9691) );
  NAND2_X1 U12237 ( .A1(n9698), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n13802) );
  NAND2_X1 U12238 ( .A1(n13803), .A2(n13802), .ZN(n9690) );
  NAND2_X1 U12239 ( .A1(n9691), .A2(n9690), .ZN(n13813) );
  INV_X1 U12240 ( .A(n13801), .ZN(n13800) );
  NAND2_X1 U12241 ( .A1(n13800), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n13812) );
  NAND2_X1 U12242 ( .A1(n13813), .A2(n13812), .ZN(n9692) );
  NAND2_X1 U12243 ( .A1(n9693), .A2(n9692), .ZN(n13832) );
  NAND2_X1 U12244 ( .A1(n13821), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n13831) );
  INV_X1 U12245 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n15240) );
  MUX2_X1 U12246 ( .A(n15240), .B(P1_REG2_REG_4__SCAN_IN), .S(n13828), .Z(
        n13830) );
  AOI21_X1 U12247 ( .B1(n13832), .B2(n13831), .A(n13830), .ZN(n13829) );
  NOR2_X1 U12248 ( .A1(n9694), .A2(n15240), .ZN(n9726) );
  MUX2_X1 U12249 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10847), .S(n9705), .Z(n9727) );
  OAI21_X1 U12250 ( .B1(n13829), .B2(n9726), .A(n9727), .ZN(n9920) );
  NAND2_X1 U12251 ( .A1(n9705), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9919) );
  MUX2_X1 U12252 ( .A(n10942), .B(P1_REG2_REG_6__SCAN_IN), .S(n9707), .Z(n9918) );
  AOI21_X1 U12253 ( .B1(n9920), .B2(n9919), .A(n9918), .ZN(n9953) );
  NOR2_X1 U12254 ( .A1(n9924), .A2(n10942), .ZN(n9952) );
  MUX2_X1 U12255 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10924), .S(n9709), .Z(n9951) );
  OAI21_X1 U12256 ( .B1(n9953), .B2(n9952), .A(n9951), .ZN(n9950) );
  NAND2_X1 U12257 ( .A1(n9709), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9696) );
  MUX2_X1 U12258 ( .A(n9783), .B(P1_REG2_REG_8__SCAN_IN), .S(n9780), .Z(n9695)
         );
  AOI21_X1 U12259 ( .B1(n9950), .B2(n9696), .A(n9695), .ZN(n9787) );
  NAND3_X1 U12260 ( .A1(n9950), .A2(n9696), .A3(n9695), .ZN(n9697) );
  NAND2_X1 U12261 ( .A1(n13873), .A2(n9697), .ZN(n9717) );
  MUX2_X1 U12262 ( .A(n9045), .B(P1_REG1_REG_2__SCAN_IN), .S(n13801), .Z(
        n13808) );
  NAND2_X1 U12263 ( .A1(n9698), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9699) );
  NAND2_X1 U12264 ( .A1(n9700), .A2(n9699), .ZN(n13807) );
  NAND2_X1 U12265 ( .A1(n13808), .A2(n13807), .ZN(n13806) );
  NAND2_X1 U12266 ( .A1(n13800), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9701) );
  NAND2_X1 U12267 ( .A1(n13806), .A2(n9701), .ZN(n13819) );
  XNOR2_X1 U12268 ( .A(n13821), .B(n9702), .ZN(n13820) );
  NAND2_X1 U12269 ( .A1(n13819), .A2(n13820), .ZN(n13818) );
  NAND2_X1 U12270 ( .A1(n13821), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9703) );
  NAND2_X1 U12271 ( .A1(n13818), .A2(n9703), .ZN(n13837) );
  XNOR2_X1 U12272 ( .A(n13828), .B(n14681), .ZN(n13838) );
  AND2_X1 U12273 ( .A1(n13837), .A2(n13838), .ZN(n13835) );
  MUX2_X1 U12274 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n9704), .S(n9705), .Z(n9721)
         );
  NAND2_X1 U12275 ( .A1(n9722), .A2(n9721), .ZN(n9720) );
  OAI21_X1 U12276 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n9705), .A(n9720), .ZN(
        n9916) );
  MUX2_X1 U12277 ( .A(n9706), .B(P1_REG1_REG_6__SCAN_IN), .S(n9707), .Z(n9917)
         );
  NOR2_X1 U12278 ( .A1(n9916), .A2(n9917), .ZN(n9915) );
  MUX2_X1 U12279 ( .A(n9708), .B(P1_REG1_REG_7__SCAN_IN), .S(n9709), .Z(n9948)
         );
  NOR2_X1 U12280 ( .A1(n9949), .A2(n9948), .ZN(n9947) );
  MUX2_X1 U12281 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n9710), .S(n9780), .Z(n9711)
         );
  NAND2_X1 U12282 ( .A1(n9712), .A2(n9711), .ZN(n9779) );
  OAI21_X1 U12283 ( .B1(n9712), .B2(n9711), .A(n9779), .ZN(n9713) );
  NAND2_X1 U12284 ( .A1(n9713), .A2(n14604), .ZN(n9716) );
  AND2_X1 U12285 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n11346) );
  NOR2_X1 U12286 ( .A1(n14598), .A2(n9784), .ZN(n9714) );
  AOI211_X1 U12287 ( .C1(n13817), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n11346), .B(
        n9714), .ZN(n9715) );
  OAI211_X1 U12288 ( .C1(n9787), .C2(n9717), .A(n9716), .B(n9715), .ZN(
        P1_U3251) );
  INV_X1 U12289 ( .A(n9718), .ZN(n9777) );
  INV_X1 U12290 ( .A(n10296), .ZN(n10174) );
  OAI222_X1 U12291 ( .A1(n13605), .A2(n9777), .B1(n10174), .B2(P2_U3088), .C1(
        n9719), .C2(n13614), .ZN(P2_U3316) );
  OAI21_X1 U12292 ( .B1(n9722), .B2(n9721), .A(n9720), .ZN(n9732) );
  NOR2_X1 U12293 ( .A1(n9723), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10999) );
  AOI21_X1 U12294 ( .B1(n13817), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n10999), .ZN(
        n9724) );
  OAI21_X1 U12295 ( .B1(n14598), .B2(n9725), .A(n9724), .ZN(n9731) );
  INV_X1 U12296 ( .A(n9920), .ZN(n9729) );
  NOR3_X1 U12297 ( .A1(n13829), .A2(n9727), .A3(n9726), .ZN(n9728) );
  NOR3_X1 U12298 ( .A1(n14600), .A2(n9729), .A3(n9728), .ZN(n9730) );
  AOI211_X1 U12299 ( .C1(n14604), .C2(n9732), .A(n9731), .B(n9730), .ZN(n9733)
         );
  INV_X1 U12300 ( .A(n9733), .ZN(P1_U3248) );
  INV_X1 U12301 ( .A(n10497), .ZN(n9735) );
  XNOR2_X1 U12302 ( .A(n10199), .B(n9736), .ZN(n10102) );
  NAND2_X1 U12303 ( .A1(n8312), .A2(n10035), .ZN(n10103) );
  XNOR2_X1 U12304 ( .A(n10102), .B(n10103), .ZN(n10101) );
  NAND2_X1 U12305 ( .A1(n9738), .A2(n10040), .ZN(n9981) );
  NAND2_X1 U12306 ( .A1(n10040), .A2(n13390), .ZN(n9739) );
  NAND2_X1 U12307 ( .A1(n10199), .A2(n11088), .ZN(n9740) );
  XOR2_X1 U12308 ( .A(n10101), .B(n10100), .Z(n9775) );
  INV_X1 U12309 ( .A(P2_B_REG_SCAN_IN), .ZN(n11857) );
  XNOR2_X1 U12310 ( .A(n13610), .B(n11857), .ZN(n9741) );
  INV_X1 U12311 ( .A(n9743), .ZN(n13607) );
  NAND2_X1 U12312 ( .A1(n9741), .A2(n13607), .ZN(n9742) );
  INV_X1 U12313 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14825) );
  NAND2_X1 U12314 ( .A1(n14820), .A2(n14825), .ZN(n9745) );
  OR2_X1 U12315 ( .A1(n13603), .A2(n9743), .ZN(n9744) );
  NAND2_X1 U12316 ( .A1(n9745), .A2(n9744), .ZN(n14826) );
  INV_X1 U12317 ( .A(n14826), .ZN(n9756) );
  NOR2_X1 U12318 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n9749) );
  NOR4_X1 U12319 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n9748) );
  NOR4_X1 U12320 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n9747) );
  NOR4_X1 U12321 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n9746) );
  NAND4_X1 U12322 ( .A1(n9749), .A2(n9748), .A3(n9747), .A4(n9746), .ZN(n9755)
         );
  NOR4_X1 U12323 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n9753) );
  NOR4_X1 U12324 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n9752) );
  NOR4_X1 U12325 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9751) );
  NOR4_X1 U12326 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n9750) );
  NAND4_X1 U12327 ( .A1(n9753), .A2(n9752), .A3(n9751), .A4(n9750), .ZN(n9754)
         );
  OAI21_X1 U12328 ( .B1(n9755), .B2(n9754), .A(n14820), .ZN(n9858) );
  NAND2_X1 U12329 ( .A1(n9756), .A2(n9858), .ZN(n10494) );
  INV_X1 U12330 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14823) );
  NOR2_X1 U12331 ( .A1(n13603), .A2(n13610), .ZN(n9757) );
  AOI21_X1 U12332 ( .B1(n14820), .B2(n14823), .A(n9757), .ZN(n10433) );
  NAND2_X1 U12333 ( .A1(n10433), .A2(n14827), .ZN(n14822) );
  OR2_X1 U12334 ( .A1(n10494), .A2(n14822), .ZN(n9763) );
  INV_X1 U12335 ( .A(n9763), .ZN(n9760) );
  INV_X1 U12336 ( .A(n9865), .ZN(n9761) );
  NAND2_X1 U12337 ( .A1(n9769), .A2(n9761), .ZN(n14841) );
  INV_X1 U12338 ( .A(n9768), .ZN(n9758) );
  AND2_X1 U12339 ( .A1(n14841), .A2(n9758), .ZN(n9759) );
  NAND2_X1 U12340 ( .A1(n9761), .A2(n9863), .ZN(n10500) );
  NAND2_X1 U12341 ( .A1(n13390), .A2(n8286), .ZN(n9859) );
  INV_X1 U12342 ( .A(n9859), .ZN(n9762) );
  OAI21_X2 U12343 ( .B1(n9763), .B2(n10500), .A(n13407), .ZN(n14697) );
  NOR2_X2 U12344 ( .A1(n9763), .A2(n9769), .ZN(n14694) );
  NAND2_X1 U12345 ( .A1(n8313), .A2(n14522), .ZN(n9766) );
  NAND2_X1 U12346 ( .A1(n9768), .A2(n9764), .ZN(n13067) );
  NAND2_X1 U12347 ( .A1(n13111), .A2(n14524), .ZN(n9765) );
  NAND2_X1 U12348 ( .A1(n9766), .A2(n9765), .ZN(n9984) );
  INV_X1 U12349 ( .A(n10433), .ZN(n9767) );
  OAI21_X1 U12350 ( .B1(n10494), .B2(n9767), .A(n9859), .ZN(n9772) );
  NAND2_X1 U12351 ( .A1(n9769), .A2(n9768), .ZN(n9860) );
  AND2_X1 U12352 ( .A1(n9770), .A2(n9860), .ZN(n9771) );
  NAND2_X1 U12353 ( .A1(n9772), .A2(n9771), .ZN(n10129) );
  OR2_X1 U12354 ( .A1(n10129), .A2(P2_U3088), .ZN(n10109) );
  NAND2_X1 U12355 ( .A1(n10109), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n9773) );
  OAI211_X1 U12356 ( .C1(n9775), .C2(n13073), .A(n9774), .B(n9773), .ZN(
        P2_U3194) );
  INV_X1 U12357 ( .A(n10277), .ZN(n10273) );
  OAI222_X1 U12358 ( .A1(P1_U3086), .A2(n10273), .B1(n14300), .B2(n9777), .C1(
        n9776), .C2(n14298), .ZN(P1_U3344) );
  MUX2_X1 U12359 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n9778), .S(n9966), .Z(n9782)
         );
  OAI21_X1 U12360 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n9780), .A(n9779), .ZN(
        n9781) );
  NAND2_X1 U12361 ( .A1(n9781), .A2(n9782), .ZN(n9963) );
  OAI21_X1 U12362 ( .B1(n9782), .B2(n9781), .A(n9963), .ZN(n9795) );
  NOR2_X1 U12363 ( .A1(n9784), .A2(n9783), .ZN(n9786) );
  MUX2_X1 U12364 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n11026), .S(n9966), .Z(n9785) );
  OAI21_X1 U12365 ( .B1(n9787), .B2(n9786), .A(n9785), .ZN(n9969) );
  INV_X1 U12366 ( .A(n9969), .ZN(n9789) );
  NOR3_X1 U12367 ( .A1(n9787), .A2(n9786), .A3(n9785), .ZN(n9788) );
  NOR3_X1 U12368 ( .A1(n14600), .A2(n9789), .A3(n9788), .ZN(n9794) );
  NAND2_X1 U12369 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n11307) );
  INV_X1 U12370 ( .A(n11307), .ZN(n9790) );
  AOI21_X1 U12371 ( .B1(n13817), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n9790), .ZN(
        n9791) );
  OAI21_X1 U12372 ( .B1(n14598), .B2(n9792), .A(n9791), .ZN(n9793) );
  AOI211_X1 U12373 ( .C1(n9795), .C2(n14604), .A(n9794), .B(n9793), .ZN(n9796)
         );
  INV_X1 U12374 ( .A(n9796), .ZN(P1_U3252) );
  NOR2_X1 U12375 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .ZN(
        n9800) );
  NOR4_X1 U12376 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n9799) );
  NOR4_X1 U12377 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n9798) );
  NOR4_X1 U12378 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n9797) );
  NAND4_X1 U12379 ( .A1(n9800), .A2(n9799), .A3(n9798), .A4(n9797), .ZN(n9806)
         );
  NOR4_X1 U12380 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n9804) );
  NOR4_X1 U12381 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n9803) );
  NOR4_X1 U12382 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9802) );
  NOR4_X1 U12383 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n9801) );
  NAND4_X1 U12384 ( .A1(n9804), .A2(n9803), .A3(n9802), .A4(n9801), .ZN(n9805)
         );
  OAI21_X1 U12385 ( .B1(n9806), .B2(n9805), .A(n9814), .ZN(n9827) );
  INV_X1 U12386 ( .A(n9831), .ZN(n9807) );
  AND2_X1 U12387 ( .A1(n9827), .A2(n9807), .ZN(n9834) );
  NAND2_X2 U12388 ( .A1(n9809), .A2(n8999), .ZN(n14662) );
  AOI21_X1 U12389 ( .B1(n9814), .B2(n9811), .A(n9810), .ZN(n9825) );
  INV_X1 U12390 ( .A(n9825), .ZN(n10567) );
  INV_X1 U12391 ( .A(n10566), .ZN(n9815) );
  NAND2_X1 U12392 ( .A1(n8999), .A2(n9816), .ZN(n9852) );
  OR2_X1 U12393 ( .A1(n9842), .A2(n9817), .ZN(n9818) );
  NAND2_X1 U12394 ( .A1(n11983), .A2(n9818), .ZN(n10590) );
  OR2_X1 U12395 ( .A1(n11354), .A2(n8999), .ZN(n9821) );
  NAND2_X1 U12396 ( .A1(n14304), .A2(n14008), .ZN(n9820) );
  OAI21_X1 U12397 ( .B1(n14677), .B2(n14245), .A(n10604), .ZN(n9823) );
  OAI211_X1 U12398 ( .C1(n9852), .C2(n10601), .A(n9823), .B(n10600), .ZN(
        n14258) );
  NAND2_X1 U12399 ( .A1(n14258), .A2(n14679), .ZN(n9824) );
  OAI21_X1 U12400 ( .B1(n14679), .B2(n9024), .A(n9824), .ZN(P1_U3459) );
  AND2_X1 U12401 ( .A1(n10566), .A2(n9825), .ZN(n9833) );
  NAND2_X1 U12402 ( .A1(n13753), .A2(n14135), .ZN(n13766) );
  INV_X1 U12403 ( .A(n9826), .ZN(n9830) );
  NAND2_X1 U12404 ( .A1(n9833), .A2(n9827), .ZN(n9828) );
  NAND2_X1 U12405 ( .A1(n9832), .A2(n9828), .ZN(n9829) );
  NAND2_X1 U12406 ( .A1(n9830), .A2(n9829), .ZN(n10336) );
  NOR2_X1 U12407 ( .A1(n10336), .A2(P1_U3086), .ZN(n10265) );
  INV_X1 U12408 ( .A(n10265), .ZN(n9839) );
  INV_X1 U12409 ( .A(n9833), .ZN(n9836) );
  INV_X1 U12410 ( .A(n9834), .ZN(n9835) );
  NOR2_X1 U12411 ( .A1(n9836), .A2(n9835), .ZN(n9855) );
  NOR2_X1 U12412 ( .A1(n9837), .A2(n14304), .ZN(n14608) );
  NAND2_X1 U12413 ( .A1(n9855), .A2(n14608), .ZN(n9838) );
  AOI22_X1 U12414 ( .A1(n9839), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n10023), .B2(
        n13769), .ZN(n9857) );
  OAI22_X1 U12415 ( .A1(n10140), .A2(n10601), .B1(n9841), .B2(n7224), .ZN(
        n9840) );
  INV_X1 U12416 ( .A(n9840), .ZN(n9844) );
  INV_X4 U12417 ( .A(n11935), .ZN(n11982) );
  INV_X1 U12418 ( .A(n13789), .ZN(n10150) );
  OR2_X1 U12419 ( .A1(n10140), .A2(n10150), .ZN(n9849) );
  NAND2_X1 U12420 ( .A1(n9845), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9846) );
  NAND2_X1 U12421 ( .A1(n9849), .A2(n9848), .ZN(n10136) );
  OAI21_X1 U12422 ( .B1(n9850), .B2(n10136), .A(n10139), .ZN(n13791) );
  AND2_X1 U12423 ( .A1(n14670), .A2(n9853), .ZN(n9854) );
  NAND2_X1 U12424 ( .A1(n13791), .A2(n13757), .ZN(n9856) );
  OAI211_X1 U12425 ( .C1(n10635), .C2(n13766), .A(n9857), .B(n9856), .ZN(
        P1_U3232) );
  NAND3_X1 U12426 ( .A1(n14826), .A2(n9859), .A3(n9858), .ZN(n10435) );
  INV_X1 U12427 ( .A(n9860), .ZN(n10432) );
  NOR2_X1 U12428 ( .A1(n10435), .A2(n10432), .ZN(n9862) );
  INV_X1 U12429 ( .A(n14822), .ZN(n9861) );
  INV_X1 U12430 ( .A(n11092), .ZN(n9869) );
  NOR2_X1 U12431 ( .A1(n9864), .A2(n9863), .ZN(n13516) );
  NAND2_X1 U12432 ( .A1(n8312), .A2(n14524), .ZN(n11087) );
  OAI21_X1 U12433 ( .B1(n9865), .B2(n11088), .A(n11087), .ZN(n9866) );
  AOI21_X1 U12434 ( .B1(n9869), .B2(n13516), .A(n9866), .ZN(n9871) );
  INV_X1 U12435 ( .A(n10976), .ZN(n13402) );
  NOR2_X1 U12436 ( .A1(n7505), .A2(n11396), .ZN(n9867) );
  OAI21_X1 U12437 ( .B1(n13402), .B2(n14520), .A(n9869), .ZN(n9870) );
  AND2_X1 U12438 ( .A1(n9871), .A2(n9870), .ZN(n14829) );
  NAND2_X1 U12439 ( .A1(n14850), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9872) );
  OAI21_X1 U12440 ( .B1(n14850), .B2(n14829), .A(n9872), .ZN(P2_U3499) );
  INV_X1 U12441 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9873) );
  NAND2_X1 U12442 ( .A1(n14770), .A2(n9873), .ZN(n9874) );
  OAI211_X1 U12443 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n14791), .A(n9874), .B(
        n14774), .ZN(n9875) );
  INV_X1 U12444 ( .A(n9875), .ZN(n9877) );
  AOI22_X1 U12445 ( .A1(n14765), .A2(P2_REG1_REG_0__SCAN_IN), .B1(n14770), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n9876) );
  MUX2_X1 U12446 ( .A(n9877), .B(n9876), .S(n7559), .Z(n9879) );
  AOI22_X1 U12447 ( .A1(n14719), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n9878) );
  NAND2_X1 U12448 ( .A1(n9879), .A2(n9878), .ZN(P2_U3214) );
  AOI211_X1 U12449 ( .C1(n9882), .C2(n9881), .A(n9880), .B(n14795), .ZN(n9890)
         );
  AOI211_X1 U12450 ( .C1(n6565), .C2(n9884), .A(n9883), .B(n14791), .ZN(n9889)
         );
  NAND2_X1 U12451 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n9886) );
  NAND2_X1 U12452 ( .A1(n14719), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9885) );
  OAI211_X1 U12453 ( .C1(n14774), .C2(n9887), .A(n9886), .B(n9885), .ZN(n9888)
         );
  OR3_X1 U12454 ( .A1(n9890), .A2(n9889), .A3(n9888), .ZN(P2_U3220) );
  INV_X1 U12455 ( .A(n9891), .ZN(n9978) );
  INV_X1 U12456 ( .A(n11186), .ZN(n10292) );
  OAI222_X1 U12457 ( .A1(n13605), .A2(n9978), .B1(n10292), .B2(P2_U3088), .C1(
        n9892), .C2(n13614), .ZN(P2_U3315) );
  AOI211_X1 U12458 ( .C1(n9895), .C2(n9894), .A(n14795), .B(n9893), .ZN(n9904)
         );
  AOI211_X1 U12459 ( .C1(n9898), .C2(n9897), .A(n14791), .B(n9896), .ZN(n9903)
         );
  INV_X1 U12460 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n14382) );
  NAND2_X1 U12461 ( .A1(n14802), .A2(n9899), .ZN(n9901) );
  NAND2_X1 U12462 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n9900) );
  OAI211_X1 U12463 ( .C1(n14805), .C2(n14382), .A(n9901), .B(n9900), .ZN(n9902) );
  OR3_X1 U12464 ( .A1(n9904), .A2(n9903), .A3(n9902), .ZN(P2_U3221) );
  AOI211_X1 U12465 ( .C1(n9907), .C2(n9906), .A(n14791), .B(n9905), .ZN(n9914)
         );
  AOI211_X1 U12466 ( .C1(n9910), .C2(n9909), .A(n14795), .B(n9908), .ZN(n9913)
         );
  NAND2_X1 U12467 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n10750) );
  NAND2_X1 U12468 ( .A1(n14719), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n9911) );
  OAI211_X1 U12469 ( .C1(n14774), .C2(n6633), .A(n10750), .B(n9911), .ZN(n9912) );
  OR3_X1 U12470 ( .A1(n9914), .A2(n9913), .A3(n9912), .ZN(P2_U3222) );
  INV_X1 U12471 ( .A(n14604), .ZN(n13847) );
  AOI211_X1 U12472 ( .C1(n9917), .C2(n9916), .A(n9915), .B(n13847), .ZN(n9927)
         );
  AND3_X1 U12473 ( .A1(n9920), .A2(n9919), .A3(n9918), .ZN(n9921) );
  NOR3_X1 U12474 ( .A1(n14600), .A2(n9953), .A3(n9921), .ZN(n9926) );
  INV_X1 U12475 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n10875) );
  NOR2_X1 U12476 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10875), .ZN(n9922) );
  AOI21_X1 U12477 ( .B1(n13817), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n9922), .ZN(
        n9923) );
  OAI21_X1 U12478 ( .B1(n14598), .B2(n9924), .A(n9923), .ZN(n9925) );
  OR3_X1 U12479 ( .A1(n9927), .A2(n9926), .A3(n9925), .ZN(P1_U3249) );
  CLKBUF_X1 U12480 ( .A(n9928), .Z(n9946) );
  INV_X1 U12481 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n15141) );
  NOR2_X1 U12482 ( .A1(n9946), .A2(n15141), .ZN(P3_U3243) );
  INV_X1 U12483 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n9929) );
  NOR2_X1 U12484 ( .A1(n9946), .A2(n9929), .ZN(P3_U3240) );
  INV_X1 U12485 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n9930) );
  NOR2_X1 U12486 ( .A1(n9946), .A2(n9930), .ZN(P3_U3241) );
  INV_X1 U12487 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n9931) );
  NOR2_X1 U12488 ( .A1(n9946), .A2(n9931), .ZN(P3_U3242) );
  INV_X1 U12489 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n9932) );
  NOR2_X1 U12490 ( .A1(n9946), .A2(n9932), .ZN(P3_U3239) );
  INV_X1 U12491 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n9933) );
  NOR2_X1 U12492 ( .A1(n9946), .A2(n9933), .ZN(P3_U3262) );
  INV_X1 U12493 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n9934) );
  NOR2_X1 U12494 ( .A1(n9946), .A2(n9934), .ZN(P3_U3237) );
  INV_X1 U12495 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n9935) );
  NOR2_X1 U12496 ( .A1(n9946), .A2(n9935), .ZN(P3_U3255) );
  INV_X1 U12497 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n9936) );
  NOR2_X1 U12498 ( .A1(n9946), .A2(n9936), .ZN(P3_U3256) );
  INV_X1 U12499 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n9937) );
  NOR2_X1 U12500 ( .A1(n9946), .A2(n9937), .ZN(P3_U3254) );
  INV_X1 U12501 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n9938) );
  NOR2_X1 U12502 ( .A1(n9946), .A2(n9938), .ZN(P3_U3235) );
  INV_X1 U12503 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n9939) );
  NOR2_X1 U12504 ( .A1(n9946), .A2(n9939), .ZN(P3_U3245) );
  INV_X1 U12505 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n9940) );
  NOR2_X1 U12506 ( .A1(n9946), .A2(n9940), .ZN(P3_U3257) );
  INV_X1 U12507 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n9941) );
  NOR2_X1 U12508 ( .A1(n9946), .A2(n9941), .ZN(P3_U3244) );
  INV_X1 U12509 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n9942) );
  NOR2_X1 U12510 ( .A1(n9946), .A2(n9942), .ZN(P3_U3263) );
  INV_X1 U12511 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n9943) );
  NOR2_X1 U12512 ( .A1(n9946), .A2(n9943), .ZN(P3_U3236) );
  INV_X1 U12513 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n9944) );
  NOR2_X1 U12514 ( .A1(n9946), .A2(n9944), .ZN(P3_U3238) );
  INV_X1 U12515 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n9945) );
  NOR2_X1 U12516 ( .A1(n9946), .A2(n9945), .ZN(P3_U3234) );
  AOI211_X1 U12517 ( .C1(n9949), .C2(n9948), .A(n13847), .B(n9947), .ZN(n9961)
         );
  INV_X1 U12518 ( .A(n9950), .ZN(n9955) );
  NOR3_X1 U12519 ( .A1(n9953), .A2(n9952), .A3(n9951), .ZN(n9954) );
  NOR3_X1 U12520 ( .A1(n14600), .A2(n9955), .A3(n9954), .ZN(n9960) );
  NAND2_X1 U12521 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n11173) );
  INV_X1 U12522 ( .A(n11173), .ZN(n9956) );
  AOI21_X1 U12523 ( .B1(n13817), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n9956), .ZN(
        n9957) );
  OAI21_X1 U12524 ( .B1(n14598), .B2(n9958), .A(n9957), .ZN(n9959) );
  OR3_X1 U12525 ( .A1(n9961), .A2(n9960), .A3(n9959), .ZN(P1_U3250) );
  INV_X1 U12526 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9962) );
  MUX2_X1 U12527 ( .A(n9962), .B(P1_REG1_REG_10__SCAN_IN), .S(n10063), .Z(
        n9965) );
  OAI21_X1 U12528 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9966), .A(n9963), .ZN(
        n9964) );
  NOR2_X1 U12529 ( .A1(n9964), .A2(n9965), .ZN(n10062) );
  AOI211_X1 U12530 ( .C1(n9965), .C2(n9964), .A(n13847), .B(n10062), .ZN(n9976) );
  NAND2_X1 U12531 ( .A1(n9966), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9968) );
  MUX2_X1 U12532 ( .A(n9155), .B(P1_REG2_REG_10__SCAN_IN), .S(n10063), .Z(
        n9967) );
  AOI21_X1 U12533 ( .B1(n9969), .B2(n9968), .A(n9967), .ZN(n10061) );
  AND3_X1 U12534 ( .A1(n9969), .A2(n9968), .A3(n9967), .ZN(n9970) );
  NOR3_X1 U12535 ( .A1(n10061), .A2(n9970), .A3(n14600), .ZN(n9975) );
  NOR2_X1 U12536 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11408), .ZN(n9971) );
  AOI21_X1 U12537 ( .B1(n13817), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n9971), .ZN(
        n9972) );
  OAI21_X1 U12538 ( .B1(n14598), .B2(n9973), .A(n9972), .ZN(n9974) );
  OR3_X1 U12539 ( .A1(n9976), .A2(n9975), .A3(n9974), .ZN(P1_U3253) );
  INV_X1 U12540 ( .A(n10459), .ZN(n10282) );
  OAI222_X1 U12541 ( .A1(P1_U3086), .A2(n10282), .B1(n14300), .B2(n9978), .C1(
        n9977), .C2(n14298), .ZN(P1_U3343) );
  OAI21_X1 U12542 ( .B1(n9980), .B2(n9979), .A(n9997), .ZN(n10562) );
  INV_X1 U12543 ( .A(n10562), .ZN(n9986) );
  INV_X1 U12544 ( .A(n13516), .ZN(n14834) );
  INV_X1 U12545 ( .A(n9981), .ZN(n9983) );
  NAND2_X1 U12546 ( .A1(n9983), .A2(n9982), .ZN(n9994) );
  OAI21_X1 U12547 ( .B1(n9983), .B2(n9982), .A(n9994), .ZN(n9985) );
  AOI21_X1 U12548 ( .B1(n9985), .B2(n14520), .A(n9984), .ZN(n10559) );
  NAND2_X1 U12549 ( .A1(n10565), .A2(n11088), .ZN(n10000) );
  OAI211_X1 U12550 ( .C1(n10565), .C2(n11088), .A(n13390), .B(n10000), .ZN(
        n10558) );
  OAI211_X1 U12551 ( .C1(n9986), .C2(n13531), .A(n10559), .B(n10558), .ZN(
        n10492) );
  OAI22_X1 U12552 ( .A1(n13541), .A2(n10565), .B1(n14852), .B2(n9987), .ZN(
        n9988) );
  AOI21_X1 U12553 ( .B1(n14852), .B2(n10492), .A(n9988), .ZN(n9989) );
  INV_X1 U12554 ( .A(n9989), .ZN(P2_U3500) );
  INV_X1 U12555 ( .A(n14450), .ZN(n12563) );
  INV_X1 U12556 ( .A(n9990), .ZN(n9992) );
  INV_X1 U12557 ( .A(SI_17_), .ZN(n9991) );
  OAI222_X1 U12558 ( .A1(n12563), .A2(P3_U3151), .B1(n14410), .B2(n9992), .C1(
        n9991), .C2(n12973), .ZN(P3_U3278) );
  NAND2_X1 U12559 ( .A1(n9994), .A2(n9993), .ZN(n10048) );
  XNOR2_X1 U12560 ( .A(n10048), .B(n9998), .ZN(n10771) );
  NAND2_X1 U12561 ( .A1(n9995), .A2(n10565), .ZN(n9996) );
  OAI21_X1 U12562 ( .B1(n9999), .B2(n9998), .A(n10044), .ZN(n10767) );
  AOI22_X1 U12563 ( .A1(n14522), .A2(n8312), .B1(n13110), .B2(n14524), .ZN(
        n10768) );
  INV_X1 U12564 ( .A(n10768), .ZN(n10001) );
  AOI211_X1 U12565 ( .C1(n10107), .C2(n10000), .A(n10035), .B(n10046), .ZN(
        n10764) );
  AOI211_X1 U12566 ( .C1(n14845), .C2(n10767), .A(n10001), .B(n10764), .ZN(
        n10002) );
  OAI21_X1 U12567 ( .B1(n13538), .B2(n10771), .A(n10002), .ZN(n10467) );
  OAI22_X1 U12568 ( .A1(n13541), .A2(n6896), .B1(n14852), .B2(n10003), .ZN(
        n10004) );
  AOI21_X1 U12569 ( .B1(n10467), .B2(n14852), .A(n10004), .ZN(n10005) );
  INV_X1 U12570 ( .A(n10005), .ZN(P2_U3501) );
  INV_X1 U12571 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10006) );
  MUX2_X1 U12572 ( .A(n10006), .B(P2_REG1_REG_10__SCAN_IN), .S(n10176), .Z(
        n10009) );
  OAI21_X1 U12573 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n10013), .A(n10007), .ZN(
        n10008) );
  NOR2_X1 U12574 ( .A1(n10008), .A2(n10009), .ZN(n10175) );
  AOI211_X1 U12575 ( .C1(n10009), .C2(n10008), .A(n14791), .B(n10175), .ZN(
        n10020) );
  INV_X1 U12576 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10010) );
  MUX2_X1 U12577 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n10010), .S(n10176), .Z(
        n10011) );
  INV_X1 U12578 ( .A(n10011), .ZN(n10015) );
  OAI21_X1 U12579 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n10013), .A(n10012), .ZN(
        n10014) );
  NOR2_X1 U12580 ( .A1(n10014), .A2(n10015), .ZN(n10167) );
  AOI211_X1 U12581 ( .C1(n10015), .C2(n10014), .A(n14795), .B(n10167), .ZN(
        n10019) );
  NAND2_X1 U12582 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n11140)
         );
  NAND2_X1 U12583 ( .A1(n14719), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n10016) );
  OAI211_X1 U12584 ( .C1(n14774), .C2(n10017), .A(n11140), .B(n10016), .ZN(
        n10018) );
  OR3_X1 U12585 ( .A1(n10020), .A2(n10019), .A3(n10018), .ZN(P2_U3224) );
  INV_X1 U12586 ( .A(n14658), .ZN(n14645) );
  AND2_X1 U12587 ( .A1(n13789), .A2(n10023), .ZN(n10021) );
  NAND2_X1 U12588 ( .A1(n10026), .A2(n10021), .ZN(n10022) );
  NAND2_X1 U12589 ( .A1(n10078), .A2(n10022), .ZN(n10581) );
  NAND2_X1 U12590 ( .A1(n7255), .A2(n10601), .ZN(n10626) );
  NAND2_X1 U12591 ( .A1(n10023), .A2(n10076), .ZN(n10024) );
  NAND2_X1 U12592 ( .A1(n10626), .A2(n10024), .ZN(n10574) );
  OAI22_X1 U12593 ( .A1(n10574), .A2(n14662), .B1(n14670), .B2(n7255), .ZN(
        n10030) );
  XNOR2_X1 U12594 ( .A(n10635), .B(n10574), .ZN(n10025) );
  MUX2_X1 U12595 ( .A(n10026), .B(n10025), .S(n10150), .Z(n10029) );
  AOI22_X1 U12596 ( .A1(n14133), .A2(n13789), .B1(n14135), .B2(n13788), .ZN(
        n10028) );
  INV_X1 U12597 ( .A(n14105), .ZN(n11323) );
  NAND2_X1 U12598 ( .A1(n10581), .A2(n11323), .ZN(n10027) );
  OAI211_X1 U12599 ( .C1(n10029), .C2(n14672), .A(n10028), .B(n10027), .ZN(
        n10578) );
  AOI211_X1 U12600 ( .C1(n14645), .C2(n10581), .A(n10030), .B(n10578), .ZN(
        n10034) );
  NAND2_X1 U12601 ( .A1(n14685), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10032) );
  OAI21_X1 U12602 ( .B1(n10034), .B2(n14685), .A(n10032), .ZN(P1_U3529) );
  NAND2_X1 U12603 ( .A1(n14678), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n10033) );
  OAI21_X1 U12604 ( .B1(n10034), .B2(n14678), .A(n10033), .ZN(P1_U3462) );
  INV_X1 U12605 ( .A(n10109), .ZN(n10042) );
  INV_X1 U12606 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n11086) );
  NAND3_X1 U12607 ( .A1(n8313), .A2(n11088), .A3(n10035), .ZN(n10036) );
  AOI21_X1 U12608 ( .B1(n10037), .B2(n10036), .A(n13073), .ZN(n10039) );
  NOR2_X1 U12609 ( .A1(n13091), .A2(n11087), .ZN(n10038) );
  AOI211_X1 U12610 ( .C1(n10040), .C2(n14697), .A(n10039), .B(n10038), .ZN(
        n10041) );
  OAI21_X1 U12611 ( .B1(n10042), .B2(n11086), .A(n10041), .ZN(P2_U3204) );
  INV_X1 U12612 ( .A(n13111), .ZN(n10049) );
  NAND2_X1 U12613 ( .A1(n10049), .A2(n6896), .ZN(n10043) );
  NAND2_X1 U12614 ( .A1(n10044), .A2(n10043), .ZN(n10045) );
  OAI21_X1 U12615 ( .B1(n10045), .B2(n10052), .A(n10185), .ZN(n11013) );
  OAI211_X1 U12616 ( .C1(n10046), .C2(n11008), .A(n13390), .B(n10187), .ZN(
        n11007) );
  INV_X1 U12617 ( .A(n11007), .ZN(n10057) );
  NAND2_X1 U12618 ( .A1(n10048), .A2(n10047), .ZN(n10051) );
  NAND2_X1 U12619 ( .A1(n10049), .A2(n10107), .ZN(n10050) );
  NAND2_X1 U12620 ( .A1(n10051), .A2(n10050), .ZN(n10189) );
  XNOR2_X1 U12621 ( .A(n10189), .B(n10188), .ZN(n10055) );
  NAND2_X1 U12622 ( .A1(n13111), .A2(n14522), .ZN(n10054) );
  NAND2_X1 U12623 ( .A1(n13109), .A2(n14524), .ZN(n10053) );
  NAND2_X1 U12624 ( .A1(n10054), .A2(n10053), .ZN(n10158) );
  AOI21_X1 U12625 ( .B1(n10055), .B2(n14520), .A(n10158), .ZN(n11009) );
  INV_X1 U12626 ( .A(n11009), .ZN(n10056) );
  AOI211_X1 U12627 ( .C1(n14845), .C2(n11013), .A(n10057), .B(n10056), .ZN(
        n10448) );
  AOI22_X1 U12628 ( .A1(n11748), .A2(n10190), .B1(n14850), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n10058) );
  OAI21_X1 U12629 ( .B1(n10448), .B2(n14850), .A(n10058), .ZN(P2_U3502) );
  INV_X1 U12630 ( .A(n10682), .ZN(n10457) );
  INV_X1 U12631 ( .A(n10059), .ZN(n10154) );
  OAI222_X1 U12632 ( .A1(P1_U3086), .A2(n10457), .B1(n14300), .B2(n10154), 
        .C1(n10060), .C2(n14298), .ZN(P1_U3342) );
  AOI21_X1 U12633 ( .B1(n10063), .B2(P1_REG2_REG_10__SCAN_IN), .A(n10061), 
        .ZN(n10271) );
  MUX2_X1 U12634 ( .A(n9172), .B(P1_REG2_REG_11__SCAN_IN), .S(n10277), .Z(
        n10270) );
  XNOR2_X1 U12635 ( .A(n10271), .B(n10270), .ZN(n10072) );
  MUX2_X1 U12636 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10064), .S(n10277), .Z(
        n10065) );
  NAND2_X1 U12637 ( .A1(n10066), .A2(n10065), .ZN(n10276) );
  OAI21_X1 U12638 ( .B1(n10066), .B2(n10065), .A(n10276), .ZN(n10067) );
  NAND2_X1 U12639 ( .A1(n10067), .A2(n14604), .ZN(n10071) );
  NAND2_X1 U12640 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n11689)
         );
  INV_X1 U12641 ( .A(n11689), .ZN(n10069) );
  NOR2_X1 U12642 ( .A1(n14598), .A2(n10273), .ZN(n10068) );
  AOI211_X1 U12643 ( .C1(n13817), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n10069), 
        .B(n10068), .ZN(n10070) );
  OAI211_X1 U12644 ( .C1(n14600), .C2(n10072), .A(n10071), .B(n10070), .ZN(
        P1_U3254) );
  INV_X1 U12645 ( .A(n12582), .ZN(n12577) );
  INV_X1 U12646 ( .A(n10073), .ZN(n10075) );
  INV_X1 U12647 ( .A(SI_18_), .ZN(n10074) );
  OAI222_X1 U12648 ( .A1(n12577), .A2(P3_U3151), .B1(n14410), .B2(n10075), 
        .C1(n10074), .C2(n12973), .ZN(P3_U3277) );
  NAND2_X1 U12649 ( .A1(n10078), .A2(n10077), .ZN(n10625) );
  OR2_X1 U12650 ( .A1(n10631), .A2(n13788), .ZN(n10079) );
  NAND2_X1 U12651 ( .A1(n10623), .A2(n10079), .ZN(n10081) );
  OR2_X1 U12652 ( .A1(n10081), .A2(n10080), .ZN(n10082) );
  NAND2_X1 U12653 ( .A1(n10512), .A2(n10082), .ZN(n11838) );
  INV_X1 U12654 ( .A(n11838), .ZN(n10096) );
  NAND2_X1 U12655 ( .A1(n11838), .A2(n11323), .ZN(n10092) );
  NAND2_X1 U12656 ( .A1(n10632), .A2(n10085), .ZN(n10087) );
  NAND2_X1 U12657 ( .A1(n10087), .A2(n10086), .ZN(n10515) );
  OAI21_X1 U12658 ( .B1(n10087), .B2(n10086), .A(n10515), .ZN(n10090) );
  OR2_X1 U12659 ( .A1(n14102), .A2(n10612), .ZN(n10088) );
  OAI21_X1 U12660 ( .B1(n10260), .B2(n14078), .A(n10088), .ZN(n10089) );
  AOI21_X1 U12661 ( .B1(n10090), .B2(n14245), .A(n10089), .ZN(n10091) );
  NAND2_X1 U12662 ( .A1(n10092), .A2(n10091), .ZN(n11836) );
  INV_X1 U12663 ( .A(n11836), .ZN(n10095) );
  OR2_X1 U12664 ( .A1(n10631), .A2(n10626), .ZN(n10627) );
  NOR2_X1 U12665 ( .A1(n10627), .A2(n10331), .ZN(n10592) );
  AND2_X1 U12666 ( .A1(n10627), .A2(n10331), .ZN(n10093) );
  NOR2_X1 U12667 ( .A1(n10592), .A2(n10093), .ZN(n11840) );
  AOI22_X1 U12668 ( .A1(n11840), .A2(n14654), .B1(n14653), .B2(n10331), .ZN(
        n10094) );
  OAI211_X1 U12669 ( .C1(n10096), .C2(n14658), .A(n10095), .B(n10094), .ZN(
        n10098) );
  NAND2_X1 U12670 ( .A1(n10098), .A2(n14687), .ZN(n10097) );
  OAI21_X1 U12671 ( .B1(n14687), .B2(n9702), .A(n10097), .ZN(P1_U3531) );
  NAND2_X1 U12672 ( .A1(n10098), .A2(n14679), .ZN(n10099) );
  OAI21_X1 U12673 ( .B1(n14679), .B2(n6898), .A(n10099), .ZN(P1_U3468) );
  NAND2_X1 U12674 ( .A1(n10101), .A2(n10100), .ZN(n10106) );
  INV_X1 U12675 ( .A(n10102), .ZN(n10104) );
  NAND2_X1 U12676 ( .A1(n10104), .A2(n10103), .ZN(n10105) );
  XNOR2_X1 U12677 ( .A(n10199), .B(n10107), .ZN(n10114) );
  NAND2_X1 U12678 ( .A1(n13111), .A2(n10035), .ZN(n10115) );
  XNOR2_X1 U12679 ( .A(n10114), .B(n10115), .ZN(n10112) );
  XOR2_X1 U12680 ( .A(n10113), .B(n10112), .Z(n10111) );
  OAI22_X1 U12681 ( .A1(n6896), .A2(n13096), .B1(n13091), .B2(n10768), .ZN(
        n10108) );
  AOI21_X1 U12682 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n10109), .A(n10108), .ZN(
        n10110) );
  OAI21_X1 U12683 ( .B1(n10111), .B2(n13073), .A(n10110), .ZN(P2_U3209) );
  NAND2_X1 U12684 ( .A1(n13109), .A2(n10035), .ZN(n10197) );
  INV_X1 U12685 ( .A(n10114), .ZN(n10116) );
  NAND2_X1 U12686 ( .A1(n10116), .A2(n10115), .ZN(n10117) );
  XNOR2_X1 U12687 ( .A(n12048), .B(n10190), .ZN(n10121) );
  INV_X1 U12688 ( .A(n10121), .ZN(n10119) );
  NAND2_X1 U12689 ( .A1(n13110), .A2(n10035), .ZN(n10120) );
  INV_X1 U12690 ( .A(n10120), .ZN(n10118) );
  NAND2_X1 U12691 ( .A1(n10119), .A2(n10118), .ZN(n10124) );
  NAND2_X1 U12692 ( .A1(n10121), .A2(n10120), .ZN(n10122) );
  NAND2_X1 U12693 ( .A1(n10160), .A2(n10124), .ZN(n10127) );
  INV_X1 U12694 ( .A(n10203), .ZN(n10126) );
  AOI21_X1 U12695 ( .B1(n10128), .B2(n10127), .A(n10126), .ZN(n10135) );
  NOR2_X1 U12696 ( .A1(n14701), .A2(n10130), .ZN(n10133) );
  AOI22_X1 U12697 ( .A1(n14522), .A2(n13110), .B1(n13108), .B2(n14524), .ZN(
        n10194) );
  INV_X1 U12698 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10131) );
  OAI22_X1 U12699 ( .A1(n13091), .A2(n10194), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10131), .ZN(n10132) );
  AOI211_X1 U12700 ( .C1(n10499), .C2(n14697), .A(n10133), .B(n10132), .ZN(
        n10134) );
  OAI21_X1 U12701 ( .B1(n10135), .B2(n13073), .A(n10134), .ZN(P2_U3202) );
  INV_X1 U12702 ( .A(n10136), .ZN(n10137) );
  NAND2_X1 U12703 ( .A1(n10137), .A2(n11983), .ZN(n10138) );
  OAI22_X1 U12704 ( .A1(n6402), .A2(n10635), .B1(n7255), .B2(n10140), .ZN(
        n10142) );
  INV_X1 U12705 ( .A(n10147), .ZN(n10144) );
  NAND2_X1 U12706 ( .A1(n10147), .A2(n10146), .ZN(n10148) );
  AOI21_X1 U12707 ( .B1(n10262), .B2(n10148), .A(n13771), .ZN(n10153) );
  INV_X1 U12708 ( .A(n13769), .ZN(n13741) );
  OAI22_X1 U12709 ( .A1(n10265), .A2(n10149), .B1(n13741), .B2(n7255), .ZN(
        n10152) );
  NAND2_X1 U12710 ( .A1(n13753), .A2(n14133), .ZN(n13765) );
  OAI22_X1 U12711 ( .A1(n10150), .A2(n13765), .B1(n13766), .B2(n10260), .ZN(
        n10151) );
  OR3_X1 U12712 ( .A1(n10153), .A2(n10152), .A3(n10151), .ZN(P1_U3222) );
  INV_X1 U12713 ( .A(n11188), .ZN(n14773) );
  OAI222_X1 U12714 ( .A1(n13614), .A2(n10155), .B1(n14773), .B2(P2_U3088), 
        .C1(n13605), .C2(n10154), .ZN(P2_U3314) );
  OAI222_X1 U12715 ( .A1(n12594), .A2(P3_U3151), .B1(n14410), .B2(n10157), 
        .C1(n10156), .C2(n12973), .ZN(P3_U3276) );
  INV_X1 U12716 ( .A(n14701), .ZN(n13093) );
  AOI22_X1 U12717 ( .A1(n14694), .A2(n10158), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10159) );
  OAI21_X1 U12718 ( .B1(n13096), .B2(n11008), .A(n10159), .ZN(n10165) );
  INV_X1 U12719 ( .A(n10160), .ZN(n10161) );
  AOI211_X1 U12720 ( .C1(n10163), .C2(n10162), .A(n13073), .B(n10161), .ZN(
        n10164) );
  AOI211_X1 U12721 ( .C1(n13093), .C2(n7724), .A(n10165), .B(n10164), .ZN(
        n10166) );
  INV_X1 U12722 ( .A(n10166), .ZN(P2_U3190) );
  INV_X1 U12723 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10168) );
  MUX2_X1 U12724 ( .A(n10168), .B(P2_REG2_REG_11__SCAN_IN), .S(n10296), .Z(
        n10169) );
  INV_X1 U12725 ( .A(n10169), .ZN(n10170) );
  NAND2_X1 U12726 ( .A1(n10171), .A2(n10170), .ZN(n10295) );
  OAI21_X1 U12727 ( .B1(n10171), .B2(n10170), .A(n10295), .ZN(n10182) );
  NAND2_X1 U12728 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n10173)
         );
  NAND2_X1 U12729 ( .A1(n14719), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n10172) );
  OAI211_X1 U12730 ( .C1(n14774), .C2(n10174), .A(n10173), .B(n10172), .ZN(
        n10181) );
  INV_X1 U12731 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10177) );
  MUX2_X1 U12732 ( .A(n10177), .B(P2_REG1_REG_11__SCAN_IN), .S(n10296), .Z(
        n10178) );
  NOR2_X1 U12733 ( .A1(n10179), .A2(n10178), .ZN(n10287) );
  AOI211_X1 U12734 ( .C1(n10179), .C2(n10178), .A(n14791), .B(n10287), .ZN(
        n10180) );
  AOI211_X1 U12735 ( .C1(n14770), .C2(n10182), .A(n10181), .B(n10180), .ZN(
        n10183) );
  INV_X1 U12736 ( .A(n10183), .ZN(P2_U3225) );
  INV_X1 U12737 ( .A(n13110), .ZN(n10191) );
  NAND2_X1 U12738 ( .A1(n10191), .A2(n11008), .ZN(n10184) );
  OAI21_X1 U12739 ( .B1(n10186), .B2(n10352), .A(n10358), .ZN(n10509) );
  INV_X1 U12740 ( .A(n10362), .ZN(n10364) );
  AOI211_X1 U12741 ( .C1(n10499), .C2(n10187), .A(n10035), .B(n10364), .ZN(
        n10503) );
  NAND2_X1 U12742 ( .A1(n10189), .A2(n10188), .ZN(n10193) );
  NAND2_X1 U12743 ( .A1(n10191), .A2(n10190), .ZN(n10192) );
  XNOR2_X1 U12744 ( .A(n10354), .B(n10352), .ZN(n10195) );
  OAI21_X1 U12745 ( .B1(n10195), .B2(n13538), .A(n10194), .ZN(n10506) );
  AOI211_X1 U12746 ( .C1(n14845), .C2(n10509), .A(n10503), .B(n10506), .ZN(
        n10440) );
  AOI22_X1 U12747 ( .A1(n11748), .A2(n10499), .B1(n14850), .B2(
        P2_REG1_REG_4__SCAN_IN), .ZN(n10196) );
  OAI21_X1 U12748 ( .B1(n10440), .B2(n14850), .A(n10196), .ZN(P2_U3503) );
  NAND2_X1 U12749 ( .A1(n10198), .A2(n10197), .ZN(n10201) );
  XNOR2_X1 U12750 ( .A(n11100), .B(n12995), .ZN(n10407) );
  NAND2_X1 U12751 ( .A1(n13108), .A2(n10035), .ZN(n10408) );
  XNOR2_X1 U12752 ( .A(n10407), .B(n10408), .ZN(n10200) );
  INV_X1 U12753 ( .A(n10200), .ZN(n10202) );
  NAND3_X1 U12754 ( .A1(n10203), .A2(n10202), .A3(n10201), .ZN(n10204) );
  AOI21_X1 U12755 ( .B1(n10411), .B2(n10204), .A(n13073), .ZN(n10210) );
  INV_X1 U12756 ( .A(n11100), .ZN(n10474) );
  NAND2_X1 U12757 ( .A1(n13093), .A2(n11094), .ZN(n10208) );
  NAND2_X1 U12758 ( .A1(n13109), .A2(n14522), .ZN(n10206) );
  NAND2_X1 U12759 ( .A1(n13107), .A2(n14524), .ZN(n10205) );
  AND2_X1 U12760 ( .A1(n10206), .A2(n10205), .ZN(n10365) );
  INV_X1 U12761 ( .A(n10365), .ZN(n11097) );
  AOI22_X1 U12762 ( .A1(n14694), .A2(n11097), .B1(P2_REG3_REG_5__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10207) );
  OAI211_X1 U12763 ( .C1(n13096), .C2(n10474), .A(n10208), .B(n10207), .ZN(
        n10209) );
  OR2_X1 U12764 ( .A1(n10210), .A2(n10209), .ZN(P2_U3199) );
  INV_X1 U12765 ( .A(n10239), .ZN(n10215) );
  OR2_X1 U12766 ( .A1(n10224), .A2(n10236), .ZN(n10214) );
  OAI211_X1 U12767 ( .C1(n12419), .C2(n12415), .A(n10211), .B(n10694), .ZN(
        n10212) );
  INV_X1 U12768 ( .A(n10212), .ZN(n10213) );
  OAI211_X1 U12769 ( .C1(n10241), .C2(n10215), .A(n10214), .B(n10213), .ZN(
        n10216) );
  NAND2_X1 U12770 ( .A1(n10216), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10218) );
  OR2_X1 U12771 ( .A1(n10224), .A2(n12423), .ZN(n10217) );
  AND2_X1 U12772 ( .A1(n10218), .A2(n10217), .ZN(n12181) );
  NOR2_X1 U12773 ( .A1(n12198), .A2(P3_U3151), .ZN(n10314) );
  INV_X1 U12774 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n10705) );
  AND2_X1 U12775 ( .A1(n15067), .A2(n12419), .ZN(n10219) );
  INV_X1 U12776 ( .A(n12196), .ZN(n10738) );
  OR2_X1 U12777 ( .A1(n10693), .A2(n15100), .ZN(n10221) );
  NAND2_X1 U12778 ( .A1(n10241), .A2(n10220), .ZN(n10222) );
  NOR2_X2 U12779 ( .A1(n10221), .A2(n15075), .ZN(n10664) );
  INV_X1 U12780 ( .A(n12185), .ZN(n12201) );
  NOR2_X1 U12781 ( .A1(n12423), .A2(n12422), .ZN(n10223) );
  NAND2_X1 U12782 ( .A1(n10224), .A2(n10223), .ZN(n12114) );
  OAI22_X1 U12783 ( .A1(n12201), .A2(n6395), .B1(n15047), .B2(n12114), .ZN(
        n10225) );
  AOI21_X1 U12784 ( .B1(n10738), .B2(n12448), .A(n10225), .ZN(n10246) );
  AND2_X1 U12785 ( .A1(n12253), .A2(n10404), .ZN(n10226) );
  NOR2_X1 U12786 ( .A1(n12419), .A2(n10226), .ZN(n10227) );
  XNOR2_X1 U12787 ( .A(n10229), .B(n15055), .ZN(n10304) );
  XNOR2_X1 U12788 ( .A(n10304), .B(n15068), .ZN(n10235) );
  NAND2_X1 U12789 ( .A1(n10228), .A2(n15047), .ZN(n10233) );
  NAND3_X1 U12790 ( .A1(n12089), .A2(n12449), .A3(n15074), .ZN(n10230) );
  INV_X1 U12791 ( .A(n10252), .ZN(n15062) );
  AOI21_X1 U12792 ( .B1(n10231), .B2(n10229), .A(n15062), .ZN(n10232) );
  NAND2_X1 U12793 ( .A1(n10253), .A2(n10232), .ZN(n10251) );
  NAND2_X1 U12794 ( .A1(n10251), .A2(n10233), .ZN(n10234) );
  NAND2_X1 U12795 ( .A1(n10234), .A2(n10235), .ZN(n10307) );
  OAI21_X1 U12796 ( .B1(n10235), .B2(n10234), .A(n10307), .ZN(n10244) );
  INV_X1 U12797 ( .A(n10236), .ZN(n10237) );
  NAND2_X1 U12798 ( .A1(n10238), .A2(n10237), .ZN(n10243) );
  AND2_X1 U12799 ( .A1(n10239), .A2(n15100), .ZN(n10318) );
  NAND3_X1 U12800 ( .A1(n10241), .A2(n10240), .A3(n10318), .ZN(n10242) );
  NAND2_X1 U12801 ( .A1(n10244), .A2(n12192), .ZN(n10245) );
  OAI211_X1 U12802 ( .C1(n10314), .C2(n10705), .A(n10246), .B(n10245), .ZN(
        P3_U3177) );
  INV_X1 U12803 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10257) );
  INV_X1 U12804 ( .A(n15065), .ZN(n10247) );
  OAI22_X1 U12805 ( .A1(n12201), .A2(n10248), .B1(n10247), .B2(n12114), .ZN(
        n10249) );
  AOI21_X1 U12806 ( .B1(n10738), .B2(n15068), .A(n10249), .ZN(n10256) );
  INV_X1 U12807 ( .A(n12259), .ZN(n15064) );
  NAND3_X1 U12808 ( .A1(n15064), .A2(n10229), .A3(n15063), .ZN(n10250) );
  OAI211_X1 U12809 ( .C1(n10253), .C2(n10252), .A(n10251), .B(n10250), .ZN(
        n10254) );
  NAND2_X1 U12810 ( .A1(n10254), .A2(n12192), .ZN(n10255) );
  OAI211_X1 U12811 ( .C1(n10314), .C2(n10257), .A(n10256), .B(n10255), .ZN(
        P3_U3162) );
  OAI22_X1 U12812 ( .A1(n10260), .A2(n10140), .B1(n11935), .B2(n14640), .ZN(
        n10258) );
  XNOR2_X1 U12813 ( .A(n10258), .B(n11948), .ZN(n10323) );
  OAI22_X1 U12814 ( .A1(n6402), .A2(n10260), .B1(n14640), .B2(n10140), .ZN(
        n10324) );
  XNOR2_X1 U12815 ( .A(n10323), .B(n10324), .ZN(n10264) );
  NAND2_X1 U12816 ( .A1(n10262), .A2(n10261), .ZN(n10263) );
  NAND2_X1 U12817 ( .A1(n10263), .A2(n10264), .ZN(n10327) );
  OAI21_X1 U12818 ( .B1(n10264), .B2(n10263), .A(n10327), .ZN(n10268) );
  OAI22_X1 U12819 ( .A1(n10265), .A2(n13798), .B1(n13741), .B2(n14640), .ZN(
        n10267) );
  OAI22_X1 U12820 ( .A1(n10635), .A2(n13765), .B1(n13766), .B2(n10636), .ZN(
        n10266) );
  AOI211_X1 U12821 ( .C1(n10268), .C2(n13757), .A(n10267), .B(n10266), .ZN(
        n10269) );
  INV_X1 U12822 ( .A(n10269), .ZN(P1_U3237) );
  AOI22_X1 U12823 ( .A1(n10459), .A2(n11326), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n10282), .ZN(n10275) );
  OR2_X1 U12824 ( .A1(n10271), .A2(n10270), .ZN(n10272) );
  OAI21_X1 U12825 ( .B1(n10273), .B2(n9172), .A(n10272), .ZN(n10274) );
  NOR2_X1 U12826 ( .A1(n10275), .A2(n10274), .ZN(n10449) );
  AOI21_X1 U12827 ( .B1(n10275), .B2(n10274), .A(n10449), .ZN(n10286) );
  AOI22_X1 U12828 ( .A1(n10459), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n9187), 
        .B2(n10282), .ZN(n10279) );
  OAI21_X1 U12829 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n10277), .A(n10276), 
        .ZN(n10278) );
  NAND2_X1 U12830 ( .A1(n10279), .A2(n10278), .ZN(n10458) );
  OAI21_X1 U12831 ( .B1(n10279), .B2(n10278), .A(n10458), .ZN(n10280) );
  NAND2_X1 U12832 ( .A1(n10280), .A2(n14604), .ZN(n10285) );
  NOR2_X1 U12833 ( .A1(n10281), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13669) );
  NOR2_X1 U12834 ( .A1(n14598), .A2(n10282), .ZN(n10283) );
  AOI211_X1 U12835 ( .C1(n13817), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n13669), 
        .B(n10283), .ZN(n10284) );
  OAI211_X1 U12836 ( .C1(n10286), .C2(n14600), .A(n10285), .B(n10284), .ZN(
        P1_U3255) );
  INV_X1 U12837 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10288) );
  MUX2_X1 U12838 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n10288), .S(n11186), .Z(
        n10289) );
  OAI21_X1 U12839 ( .B1(n10290), .B2(n10289), .A(n11185), .ZN(n10294) );
  NAND2_X1 U12840 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n14698)
         );
  NAND2_X1 U12841 ( .A1(n14719), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n10291) );
  OAI211_X1 U12842 ( .C1(n14774), .C2(n10292), .A(n14698), .B(n10291), .ZN(
        n10293) );
  AOI21_X1 U12843 ( .B1(n10294), .B2(n14765), .A(n10293), .ZN(n10303) );
  OAI21_X1 U12844 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n10296), .A(n10295), 
        .ZN(n10300) );
  INV_X1 U12845 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n10297) );
  MUX2_X1 U12846 ( .A(n10297), .B(P2_REG2_REG_12__SCAN_IN), .S(n11186), .Z(
        n10298) );
  INV_X1 U12847 ( .A(n10298), .ZN(n10299) );
  OAI21_X1 U12848 ( .B1(n10300), .B2(n10299), .A(n11181), .ZN(n10301) );
  NAND2_X1 U12849 ( .A1(n10301), .A2(n14770), .ZN(n10302) );
  NAND2_X1 U12850 ( .A1(n10303), .A2(n10302), .ZN(P2_U3226) );
  NAND2_X1 U12851 ( .A1(n10304), .A2(n8850), .ZN(n10305) );
  AND2_X1 U12852 ( .A1(n10307), .A2(n10305), .ZN(n10309) );
  XNOR2_X1 U12853 ( .A(n10368), .B(n12448), .ZN(n10308) );
  AND2_X1 U12854 ( .A1(n10308), .A2(n10305), .ZN(n10306) );
  OAI211_X1 U12855 ( .C1(n10309), .C2(n10308), .A(n12192), .B(n10371), .ZN(
        n10313) );
  INV_X1 U12856 ( .A(n12114), .ZN(n12194) );
  NOR2_X1 U12857 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10755), .ZN(n14865) );
  AOI21_X1 U12858 ( .B1(n12194), .B2(n15068), .A(n14865), .ZN(n10310) );
  OAI21_X1 U12859 ( .B1(n12201), .B2(n10776), .A(n10310), .ZN(n10311) );
  AOI21_X1 U12860 ( .B1(n10738), .B2(n12446), .A(n10311), .ZN(n10312) );
  OAI211_X1 U12861 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12181), .A(n10313), .B(
        n10312), .ZN(P3_U3158) );
  AND2_X1 U12862 ( .A1(n15065), .A2(n10622), .ZN(n12252) );
  NOR2_X1 U12863 ( .A1(n12252), .A2(n12259), .ZN(n12224) );
  INV_X1 U12864 ( .A(n10314), .ZN(n10315) );
  NAND2_X1 U12865 ( .A1(n10315), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10317) );
  AOI22_X1 U12866 ( .A1(n10738), .A2(n12449), .B1(n10665), .B2(n12185), .ZN(
        n10316) );
  OAI211_X1 U12867 ( .C1(n12224), .C2(n12187), .A(n10317), .B(n10316), .ZN(
        P3_U3172) );
  NOR2_X1 U12868 ( .A1(n10318), .A2(n15051), .ZN(n10319) );
  OAI22_X1 U12869 ( .A1(n12224), .A2(n10319), .B1(n15047), .B2(n15044), .ZN(
        n10666) );
  INV_X1 U12870 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10320) );
  NOR2_X1 U12871 ( .A1(n15108), .A2(n10320), .ZN(n10321) );
  AOI21_X1 U12872 ( .B1(n15108), .B2(n10666), .A(n10321), .ZN(n10322) );
  OAI21_X1 U12873 ( .B1(n10622), .B2(n12955), .A(n10322), .ZN(P3_U3390) );
  INV_X1 U12874 ( .A(n10323), .ZN(n10325) );
  OR2_X1 U12875 ( .A1(n10325), .A2(n10324), .ZN(n10326) );
  NAND2_X1 U12876 ( .A1(n11982), .A2(n10331), .ZN(n10329) );
  OR2_X1 U12877 ( .A1(n10140), .A2(n10636), .ZN(n10328) );
  NAND2_X1 U12878 ( .A1(n10329), .A2(n10328), .ZN(n10330) );
  XNOR2_X1 U12879 ( .A(n10330), .B(n11948), .ZN(n10607) );
  OR2_X1 U12880 ( .A1(n6402), .A2(n10636), .ZN(n10333) );
  NAND2_X1 U12881 ( .A1(n11981), .A2(n10331), .ZN(n10332) );
  NAND2_X1 U12882 ( .A1(n10333), .A2(n10332), .ZN(n10608) );
  XNOR2_X1 U12883 ( .A(n10607), .B(n10608), .ZN(n10334) );
  OAI211_X1 U12884 ( .C1(n10335), .C2(n10334), .A(n10611), .B(n13757), .ZN(
        n10341) );
  INV_X1 U12885 ( .A(n13765), .ZN(n10339) );
  OAI22_X1 U12886 ( .A1(n6936), .A2(n13741), .B1(n13766), .B2(n10612), .ZN(
        n10338) );
  MUX2_X1 U12887 ( .A(n13711), .B(P1_U3086), .S(P1_REG3_REG_3__SCAN_IN), .Z(
        n10337) );
  AOI211_X1 U12888 ( .C1(n10339), .C2(n13788), .A(n10338), .B(n10337), .ZN(
        n10340) );
  NAND2_X1 U12889 ( .A1(n10341), .A2(n10340), .ZN(P1_U3218) );
  INV_X1 U12890 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n15211) );
  NAND2_X1 U12891 ( .A1(n12349), .A2(n12450), .ZN(n10342) );
  OAI21_X1 U12892 ( .B1(n12450), .B2(n15211), .A(n10342), .ZN(P3_U3508) );
  INV_X1 U12893 ( .A(P3_DATAO_REG_12__SCAN_IN), .ZN(n15199) );
  NAND2_X1 U12894 ( .A1(n12801), .A2(n12450), .ZN(n10343) );
  OAI21_X1 U12895 ( .B1(n12450), .B2(n15199), .A(n10343), .ZN(P3_U3503) );
  INV_X1 U12896 ( .A(n10344), .ZN(n10351) );
  INV_X1 U12897 ( .A(n13135), .ZN(n13124) );
  OAI222_X1 U12898 ( .A1(n13605), .A2(n10351), .B1(n13124), .B2(P2_U3088), 
        .C1(n15254), .C2(n13614), .ZN(P2_U3313) );
  INV_X1 U12899 ( .A(n10345), .ZN(n10347) );
  OAI222_X1 U12900 ( .A1(P1_U3086), .A2(n11444), .B1(n14300), .B2(n10347), 
        .C1(n10346), .C2(n14298), .ZN(P1_U3339) );
  INV_X1 U12901 ( .A(n14801), .ZN(n10348) );
  OAI222_X1 U12902 ( .A1(n13614), .A2(n10349), .B1(n10348), .B2(P2_U3088), 
        .C1(n13605), .C2(n10347), .ZN(P2_U3311) );
  INV_X1 U12903 ( .A(n11438), .ZN(n10687) );
  OAI222_X1 U12904 ( .A1(P1_U3086), .A2(n10687), .B1(n14300), .B2(n10351), 
        .C1(n10350), .C2(n14298), .ZN(P1_U3341) );
  INV_X1 U12905 ( .A(n10352), .ZN(n10353) );
  NAND2_X1 U12906 ( .A1(n10499), .A2(n10355), .ZN(n10356) );
  INV_X1 U12907 ( .A(n10359), .ZN(n10469) );
  XNOR2_X1 U12908 ( .A(n10470), .B(n10469), .ZN(n11101) );
  OR2_X1 U12909 ( .A1(n10499), .A2(n13109), .ZN(n10357) );
  NAND2_X1 U12910 ( .A1(n10358), .A2(n10357), .ZN(n10360) );
  OAI21_X1 U12911 ( .B1(n10360), .B2(n10359), .A(n10476), .ZN(n10361) );
  INV_X1 U12912 ( .A(n10361), .ZN(n11104) );
  INV_X1 U12913 ( .A(n10481), .ZN(n10363) );
  OAI211_X1 U12914 ( .C1(n10474), .C2(n10364), .A(n10363), .B(n13390), .ZN(
        n11096) );
  OAI211_X1 U12915 ( .C1(n11104), .C2(n13531), .A(n10365), .B(n11096), .ZN(
        n10366) );
  AOI21_X1 U12916 ( .B1(n14520), .B2(n11101), .A(n10366), .ZN(n10444) );
  AOI22_X1 U12917 ( .A1(n11748), .A2(n11100), .B1(n14850), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n10367) );
  OAI21_X1 U12918 ( .B1(n10444), .B2(n14850), .A(n10367), .ZN(P2_U3504) );
  INV_X1 U12919 ( .A(n10368), .ZN(n10369) );
  NAND2_X1 U12920 ( .A1(n10369), .A2(n12448), .ZN(n10370) );
  XNOR2_X1 U12921 ( .A(n10229), .B(n15035), .ZN(n10372) );
  NAND2_X1 U12922 ( .A1(n10372), .A2(n11039), .ZN(n10645) );
  INV_X1 U12923 ( .A(n10372), .ZN(n10373) );
  NAND2_X1 U12924 ( .A1(n10373), .A2(n12446), .ZN(n10374) );
  INV_X1 U12925 ( .A(n10646), .ZN(n10375) );
  AOI21_X1 U12926 ( .B1(n10377), .B2(n10376), .A(n10375), .ZN(n10383) );
  NOR2_X1 U12927 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10378), .ZN(n14883) );
  NOR2_X1 U12928 ( .A1(n12114), .A2(n15045), .ZN(n10379) );
  AOI211_X1 U12929 ( .C1(n15035), .C2(n12185), .A(n14883), .B(n10379), .ZN(
        n10380) );
  OAI21_X1 U12930 ( .B1(n11116), .B2(n12196), .A(n10380), .ZN(n10381) );
  AOI21_X1 U12931 ( .B1(n15033), .B2(n12198), .A(n10381), .ZN(n10382) );
  OAI21_X1 U12932 ( .B1(n10383), .B2(n12187), .A(n10382), .ZN(P3_U3170) );
  INV_X1 U12933 ( .A(n13846), .ZN(n13854) );
  INV_X1 U12934 ( .A(n10384), .ZN(n10399) );
  OAI222_X1 U12935 ( .A1(P1_U3086), .A2(n13854), .B1(n14300), .B2(n10399), 
        .C1(n10385), .C2(n14298), .ZN(P1_U3338) );
  INV_X1 U12936 ( .A(n10386), .ZN(n10406) );
  OAI222_X1 U12937 ( .A1(n13605), .A2(n10406), .B1(n14779), .B2(P2_U3088), 
        .C1(n10387), .C2(n13614), .ZN(P2_U3312) );
  OAI21_X1 U12938 ( .B1(n10389), .B2(n12225), .A(n10388), .ZN(n10390) );
  INV_X1 U12939 ( .A(n10390), .ZN(n10759) );
  NAND2_X1 U12940 ( .A1(n10391), .A2(n12225), .ZN(n10392) );
  NAND3_X1 U12941 ( .A1(n10393), .A2(n15051), .A3(n10392), .ZN(n10395) );
  AOI22_X1 U12942 ( .A1(n15068), .A2(n15066), .B1(n15067), .B2(n12446), .ZN(
        n10394) );
  AND2_X1 U12943 ( .A1(n10395), .A2(n10394), .ZN(n10754) );
  OAI21_X1 U12944 ( .B1(n10759), .B2(n14494), .A(n10754), .ZN(n10778) );
  INV_X1 U12945 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n10396) );
  OAI22_X1 U12946 ( .A1(n10776), .A2(n12955), .B1(n15108), .B2(n10396), .ZN(
        n10397) );
  AOI21_X1 U12947 ( .B1(n15108), .B2(n10778), .A(n10397), .ZN(n10398) );
  INV_X1 U12948 ( .A(n10398), .ZN(P3_U3399) );
  INV_X1 U12949 ( .A(n13148), .ZN(n13145) );
  OAI222_X1 U12950 ( .A1(n13614), .A2(n10400), .B1(n13145), .B2(P2_U3088), 
        .C1(n13605), .C2(n10399), .ZN(P2_U3310) );
  INV_X1 U12951 ( .A(n10401), .ZN(n10403) );
  OAI222_X1 U12952 ( .A1(n10404), .A2(P3_U3151), .B1(n14410), .B2(n10403), 
        .C1(n10402), .C2(n12973), .ZN(P3_U3275) );
  INV_X1 U12953 ( .A(n11442), .ZN(n14599) );
  OAI222_X1 U12954 ( .A1(P1_U3086), .A2(n14599), .B1(n14300), .B2(n10406), 
        .C1(n10405), .C2(n14298), .ZN(P1_U3340) );
  INV_X1 U12955 ( .A(n10785), .ZN(n14813) );
  INV_X1 U12956 ( .A(n10407), .ZN(n10409) );
  NAND2_X1 U12957 ( .A1(n10409), .A2(n10408), .ZN(n10410) );
  XNOR2_X1 U12958 ( .A(n13079), .B(n12995), .ZN(n10412) );
  AND2_X1 U12959 ( .A1(n13107), .A2(n10035), .ZN(n10413) );
  NAND2_X1 U12960 ( .A1(n10412), .A2(n10413), .ZN(n10417) );
  INV_X1 U12961 ( .A(n10412), .ZN(n10415) );
  INV_X1 U12962 ( .A(n10413), .ZN(n10414) );
  NAND2_X1 U12963 ( .A1(n10415), .A2(n10414), .ZN(n10416) );
  AND2_X1 U12964 ( .A1(n10417), .A2(n10416), .ZN(n13076) );
  NAND2_X1 U12965 ( .A1(n13075), .A2(n10417), .ZN(n10424) );
  XNOR2_X1 U12966 ( .A(n10785), .B(n12995), .ZN(n10418) );
  AND2_X1 U12967 ( .A1(n13106), .A2(n10035), .ZN(n10419) );
  NAND2_X1 U12968 ( .A1(n10418), .A2(n10419), .ZN(n10742) );
  INV_X1 U12969 ( .A(n10418), .ZN(n10421) );
  INV_X1 U12970 ( .A(n10419), .ZN(n10420) );
  NAND2_X1 U12971 ( .A1(n10421), .A2(n10420), .ZN(n10422) );
  AND2_X1 U12972 ( .A1(n10742), .A2(n10422), .ZN(n10423) );
  NAND2_X1 U12973 ( .A1(n10424), .A2(n10423), .ZN(n10743) );
  OAI211_X1 U12974 ( .C1(n10424), .C2(n10423), .A(n10743), .B(n14692), .ZN(
        n10431) );
  NAND2_X1 U12975 ( .A1(n13107), .A2(n14522), .ZN(n10426) );
  NAND2_X1 U12976 ( .A1(n13105), .A2(n14524), .ZN(n10425) );
  NAND2_X1 U12977 ( .A1(n10426), .A2(n10425), .ZN(n10549) );
  INV_X1 U12978 ( .A(n10549), .ZN(n10428) );
  OAI22_X1 U12979 ( .A1(n13091), .A2(n10428), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10427), .ZN(n10429) );
  AOI21_X1 U12980 ( .B1(n14809), .B2(n13093), .A(n10429), .ZN(n10430) );
  OAI211_X1 U12981 ( .C1(n14813), .C2(n13096), .A(n10431), .B(n10430), .ZN(
        P2_U3185) );
  NOR2_X1 U12982 ( .A1(n10433), .A2(n10432), .ZN(n10434) );
  AND2_X1 U12983 ( .A1(n10434), .A2(n14827), .ZN(n10496) );
  INV_X1 U12984 ( .A(n10435), .ZN(n10436) );
  INV_X1 U12985 ( .A(n13584), .ZN(n10967) );
  INV_X1 U12986 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10437) );
  NOR2_X1 U12987 ( .A1(n14848), .A2(n10437), .ZN(n10438) );
  AOI21_X1 U12988 ( .B1(n10967), .B2(n10499), .A(n10438), .ZN(n10439) );
  OAI21_X1 U12989 ( .B1(n10440), .B2(n14846), .A(n10439), .ZN(P2_U3442) );
  INV_X1 U12990 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10441) );
  OAI22_X1 U12991 ( .A1(n13584), .A2(n10474), .B1(n14848), .B2(n10441), .ZN(
        n10442) );
  INV_X1 U12992 ( .A(n10442), .ZN(n10443) );
  OAI21_X1 U12993 ( .B1(n10444), .B2(n14846), .A(n10443), .ZN(P2_U3445) );
  INV_X1 U12994 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10445) );
  OAI22_X1 U12995 ( .A1(n13584), .A2(n11008), .B1(n14848), .B2(n10445), .ZN(
        n10446) );
  INV_X1 U12996 ( .A(n10446), .ZN(n10447) );
  OAI21_X1 U12997 ( .B1(n10448), .B2(n14846), .A(n10447), .ZN(P2_U3439) );
  NOR2_X1 U12998 ( .A1(n10459), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n10450) );
  NOR2_X1 U12999 ( .A1(n10450), .A2(n10449), .ZN(n10453) );
  MUX2_X1 U13000 ( .A(n11284), .B(P1_REG2_REG_13__SCAN_IN), .S(n10682), .Z(
        n10451) );
  INV_X1 U13001 ( .A(n10451), .ZN(n10452) );
  NAND2_X1 U13002 ( .A1(n10452), .A2(n10453), .ZN(n10675) );
  OAI211_X1 U13003 ( .C1(n10453), .C2(n10452), .A(n13873), .B(n10675), .ZN(
        n10456) );
  NAND2_X1 U13004 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n13726)
         );
  INV_X1 U13005 ( .A(n13726), .ZN(n10454) );
  AOI21_X1 U13006 ( .B1(n13817), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10454), 
        .ZN(n10455) );
  OAI211_X1 U13007 ( .C1(n14598), .C2(n10457), .A(n10456), .B(n10455), .ZN(
        n10464) );
  OAI21_X1 U13008 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n10459), .A(n10458), 
        .ZN(n10462) );
  MUX2_X1 U13009 ( .A(n10460), .B(P1_REG1_REG_13__SCAN_IN), .S(n10682), .Z(
        n10461) );
  NOR2_X1 U13010 ( .A1(n10462), .A2(n10461), .ZN(n10681) );
  AOI211_X1 U13011 ( .C1(n10462), .C2(n10461), .A(n10681), .B(n13847), .ZN(
        n10463) );
  OR2_X1 U13012 ( .A1(n10464), .A2(n10463), .ZN(P1_U3256) );
  INV_X1 U13013 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10465) );
  OAI22_X1 U13014 ( .A1(n13584), .A2(n6896), .B1(n14848), .B2(n10465), .ZN(
        n10466) );
  AOI21_X1 U13015 ( .B1(n10467), .B2(n14848), .A(n10466), .ZN(n10468) );
  INV_X1 U13016 ( .A(n10468), .ZN(P2_U3436) );
  NAND2_X1 U13017 ( .A1(n11100), .A2(n10473), .ZN(n10471) );
  NAND2_X1 U13018 ( .A1(n10472), .A2(n10471), .ZN(n10545) );
  XNOR2_X1 U13019 ( .A(n10545), .B(n10544), .ZN(n11065) );
  NAND2_X1 U13020 ( .A1(n10474), .A2(n10473), .ZN(n10475) );
  OAI21_X1 U13021 ( .B1(n10478), .B2(n10477), .A(n10538), .ZN(n11071) );
  INV_X1 U13022 ( .A(n11071), .ZN(n10482) );
  NAND2_X1 U13023 ( .A1(n13108), .A2(n14522), .ZN(n10480) );
  NAND2_X1 U13024 ( .A1(n13106), .A2(n14524), .ZN(n10479) );
  AND2_X1 U13025 ( .A1(n10480), .A2(n10479), .ZN(n11066) );
  INV_X1 U13026 ( .A(n13079), .ZN(n10486) );
  INV_X1 U13027 ( .A(n10541), .ZN(n10543) );
  OAI211_X1 U13028 ( .C1(n10486), .C2(n10481), .A(n10543), .B(n13390), .ZN(
        n11068) );
  OAI211_X1 U13029 ( .C1(n10482), .C2(n13531), .A(n11066), .B(n11068), .ZN(
        n10483) );
  AOI21_X1 U13030 ( .B1(n14520), .B2(n11065), .A(n10483), .ZN(n10489) );
  AOI22_X1 U13031 ( .A1(n11748), .A2(n13079), .B1(n14850), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n10484) );
  OAI21_X1 U13032 ( .B1(n10489), .B2(n14850), .A(n10484), .ZN(P2_U3505) );
  INV_X1 U13033 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10485) );
  OAI22_X1 U13034 ( .A1(n13584), .A2(n10486), .B1(n14848), .B2(n10485), .ZN(
        n10487) );
  INV_X1 U13035 ( .A(n10487), .ZN(n10488) );
  OAI21_X1 U13036 ( .B1(n10489), .B2(n14846), .A(n10488), .ZN(P2_U3448) );
  INV_X1 U13037 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10490) );
  OAI22_X1 U13038 ( .A1(n13584), .A2(n10565), .B1(n14848), .B2(n10490), .ZN(
        n10491) );
  AOI21_X1 U13039 ( .B1(n14848), .B2(n10492), .A(n10491), .ZN(n10493) );
  INV_X1 U13040 ( .A(n10493), .ZN(P2_U3433) );
  INV_X1 U13041 ( .A(n10494), .ZN(n10495) );
  NAND2_X1 U13042 ( .A1(n10496), .A2(n10495), .ZN(n10501) );
  NAND2_X1 U13043 ( .A1(n10497), .A2(n8286), .ZN(n10973) );
  AND2_X1 U13044 ( .A1(n10976), .A2(n10973), .ZN(n10498) );
  INV_X1 U13045 ( .A(n10499), .ZN(n10505) );
  AOI22_X1 U13046 ( .A1(n10503), .A2(n14806), .B1(n10502), .B2(n14808), .ZN(
        n10504) );
  OAI21_X1 U13047 ( .B1(n10505), .B2(n14812), .A(n10504), .ZN(n10508) );
  MUX2_X1 U13048 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n10506), .S(n13438), .Z(
        n10507) );
  AOI211_X1 U13049 ( .C1(n14815), .C2(n10509), .A(n10508), .B(n10507), .ZN(
        n10510) );
  INV_X1 U13050 ( .A(n10510), .ZN(P2_U3261) );
  NAND2_X1 U13051 ( .A1(n6936), .A2(n10636), .ZN(n10511) );
  NAND2_X1 U13052 ( .A1(n10512), .A2(n10511), .ZN(n10589) );
  INV_X1 U13053 ( .A(n10584), .ZN(n10588) );
  NAND2_X1 U13054 ( .A1(n14646), .A2(n10612), .ZN(n10513) );
  NAND2_X1 U13055 ( .A1(n10587), .A2(n10513), .ZN(n10801) );
  XNOR2_X1 U13056 ( .A(n10801), .B(n10799), .ZN(n10853) );
  NAND2_X1 U13057 ( .A1(n10515), .A2(n10514), .ZN(n10585) );
  NAND2_X1 U13058 ( .A1(n10617), .A2(n10612), .ZN(n10516) );
  OAI21_X1 U13059 ( .B1(n10517), .B2(n10799), .A(n10808), .ZN(n10519) );
  INV_X1 U13060 ( .A(n13784), .ZN(n11175) );
  OAI22_X1 U13061 ( .A1(n11175), .A2(n14102), .B1(n10612), .B2(n14078), .ZN(
        n11000) );
  NOR2_X1 U13062 ( .A1(n10853), .A2(n14105), .ZN(n10518) );
  AOI211_X1 U13063 ( .C1(n14245), .C2(n10519), .A(n11000), .B(n10518), .ZN(
        n10846) );
  INV_X1 U13064 ( .A(n10594), .ZN(n10521) );
  INV_X1 U13065 ( .A(n11004), .ZN(n10848) );
  INV_X1 U13066 ( .A(n10944), .ZN(n10520) );
  AOI21_X1 U13067 ( .B1(n11004), .B2(n10521), .A(n10520), .ZN(n10850) );
  AOI22_X1 U13068 ( .A1(n10850), .A2(n14654), .B1(n14653), .B2(n11004), .ZN(
        n10522) );
  OAI211_X1 U13069 ( .C1(n14658), .C2(n10853), .A(n10846), .B(n10522), .ZN(
        n10524) );
  NAND2_X1 U13070 ( .A1(n10524), .A2(n14687), .ZN(n10523) );
  OAI21_X1 U13071 ( .B1(n14687), .B2(n9704), .A(n10523), .ZN(P1_U3533) );
  INV_X1 U13072 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10526) );
  NAND2_X1 U13073 ( .A1(n10524), .A2(n14679), .ZN(n10525) );
  OAI21_X1 U13074 ( .B1(n14679), .B2(n10526), .A(n10525), .ZN(P1_U3474) );
  OAI21_X1 U13075 ( .B1(n10528), .B2(n12274), .A(n10527), .ZN(n10529) );
  INV_X1 U13076 ( .A(n10529), .ZN(n15031) );
  INV_X1 U13077 ( .A(n10530), .ZN(n10531) );
  AOI21_X1 U13078 ( .B1(n10531), .B2(n12274), .A(n15072), .ZN(n10534) );
  OAI22_X1 U13079 ( .A1(n15045), .A2(n15046), .B1(n11116), .B2(n15044), .ZN(
        n10532) );
  AOI21_X1 U13080 ( .B1(n10534), .B2(n10533), .A(n10532), .ZN(n15030) );
  OAI21_X1 U13081 ( .B1(n14494), .B2(n15031), .A(n15030), .ZN(n10773) );
  INV_X1 U13082 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n10535) );
  OAI22_X1 U13083 ( .A1(n12280), .A2(n12955), .B1(n15108), .B2(n10535), .ZN(
        n10536) );
  AOI21_X1 U13084 ( .B1(n10773), .B2(n15108), .A(n10536), .ZN(n10537) );
  INV_X1 U13085 ( .A(n10537), .ZN(P3_U3402) );
  INV_X1 U13086 ( .A(n10548), .ZN(n10539) );
  OAI21_X1 U13087 ( .B1(n10540), .B2(n10539), .A(n10781), .ZN(n14816) );
  INV_X1 U13088 ( .A(n10982), .ZN(n10542) );
  AOI211_X1 U13089 ( .C1(n10785), .C2(n10543), .A(n10035), .B(n10542), .ZN(
        n14807) );
  NAND2_X1 U13090 ( .A1(n10545), .A2(n10544), .ZN(n10547) );
  NAND2_X1 U13091 ( .A1(n13079), .A2(n6687), .ZN(n10546) );
  NAND2_X1 U13092 ( .A1(n10547), .A2(n10546), .ZN(n10788) );
  XNOR2_X1 U13093 ( .A(n10788), .B(n10548), .ZN(n10550) );
  AOI21_X1 U13094 ( .B1(n10550), .B2(n14520), .A(n10549), .ZN(n14818) );
  INV_X1 U13095 ( .A(n14818), .ZN(n10551) );
  AOI211_X1 U13096 ( .C1(n14845), .C2(n14816), .A(n14807), .B(n10551), .ZN(
        n10556) );
  INV_X1 U13097 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10552) );
  OAI22_X1 U13098 ( .A1(n13584), .A2(n14813), .B1(n14848), .B2(n10552), .ZN(
        n10553) );
  INV_X1 U13099 ( .A(n10553), .ZN(n10554) );
  OAI21_X1 U13100 ( .B1(n10556), .B2(n14846), .A(n10554), .ZN(P2_U3451) );
  AOI22_X1 U13101 ( .A1(n11748), .A2(n10785), .B1(n14850), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n10555) );
  OAI21_X1 U13102 ( .B1(n10556), .B2(n14850), .A(n10555), .ZN(P2_U3506) );
  INV_X1 U13103 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10557) );
  OAI22_X1 U13104 ( .A1(n13413), .A2(n10558), .B1(n10557), .B2(n13407), .ZN(
        n10561) );
  NOR2_X1 U13105 ( .A1(n6388), .A2(n10559), .ZN(n10560) );
  AOI211_X1 U13106 ( .C1(n6388), .C2(P2_REG2_REG_1__SCAN_IN), .A(n10561), .B(
        n10560), .ZN(n10564) );
  NAND2_X1 U13107 ( .A1(n14815), .A2(n10562), .ZN(n10563) );
  OAI211_X1 U13108 ( .C1(n10565), .C2(n14812), .A(n10564), .B(n10563), .ZN(
        P2_U3264) );
  NOR2_X1 U13109 ( .A1(n10567), .A2(n10566), .ZN(n10568) );
  NAND2_X1 U13110 ( .A1(n10569), .A2(n10568), .ZN(n14009) );
  INV_X1 U13111 ( .A(n10570), .ZN(n10571) );
  NAND2_X1 U13112 ( .A1(n14613), .A2(n10571), .ZN(n14117) );
  INV_X1 U13113 ( .A(n14117), .ZN(n11837) );
  INV_X1 U13114 ( .A(n14009), .ZN(n10573) );
  NOR2_X1 U13115 ( .A1(n14662), .A2(n14008), .ZN(n10572) );
  INV_X1 U13116 ( .A(n10574), .ZN(n10575) );
  NAND2_X1 U13117 ( .A1(n14146), .A2(n10575), .ZN(n10577) );
  INV_X1 U13118 ( .A(n14638), .ZN(n14089) );
  NAND2_X1 U13119 ( .A1(n14089), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n10576) );
  OAI211_X1 U13120 ( .C1(n14125), .C2(n7255), .A(n10577), .B(n10576), .ZN(
        n10580) );
  MUX2_X1 U13121 ( .A(n10578), .B(P1_REG2_REG_1__SCAN_IN), .S(n14091), .Z(
        n10579) );
  AOI211_X1 U13122 ( .C1(n11837), .C2(n10581), .A(n10580), .B(n10579), .ZN(
        n10582) );
  INV_X1 U13123 ( .A(n10582), .ZN(P1_U3292) );
  OAI21_X1 U13124 ( .B1(n10585), .B2(n10584), .A(n10583), .ZN(n10586) );
  AOI222_X1 U13125 ( .A1(n14245), .A2(n10586), .B1(n13785), .B2(n14135), .C1(
        n13787), .C2(n14133), .ZN(n14648) );
  MUX2_X1 U13126 ( .A(n15240), .B(n14648), .S(n14613), .Z(n10598) );
  OAI21_X1 U13127 ( .B1(n10589), .B2(n10588), .A(n10587), .ZN(n14651) );
  INV_X1 U13128 ( .A(n10590), .ZN(n10591) );
  NAND2_X1 U13129 ( .A1(n14613), .A2(n10591), .ZN(n14148) );
  INV_X1 U13130 ( .A(n14146), .ZN(n14111) );
  NOR2_X1 U13131 ( .A1(n10592), .A2(n14646), .ZN(n10593) );
  OR2_X1 U13132 ( .A1(n10594), .A2(n10593), .ZN(n14647) );
  NOR2_X1 U13133 ( .A1(n14111), .A2(n14647), .ZN(n10596) );
  OAI22_X1 U13134 ( .A1(n14125), .A2(n14646), .B1(n10614), .B2(n14638), .ZN(
        n10595) );
  AOI211_X1 U13135 ( .C1(n14651), .C2(n14621), .A(n10596), .B(n10595), .ZN(
        n10597) );
  NAND2_X1 U13136 ( .A1(n10598), .A2(n10597), .ZN(P1_U3289) );
  OAI22_X1 U13137 ( .A1(n14091), .A2(n10600), .B1(n10599), .B2(n14638), .ZN(
        n10603) );
  AOI21_X1 U13138 ( .B1(n14111), .B2(n14125), .A(n10601), .ZN(n10602) );
  AOI211_X1 U13139 ( .C1(n14091), .C2(P1_REG2_REG_0__SCAN_IN), .A(n10603), .B(
        n10602), .ZN(n10606) );
  AND2_X1 U13140 ( .A1(n14613), .A2(n14245), .ZN(n14128) );
  OAI21_X1 U13141 ( .B1(n14621), .B2(n14128), .A(n10604), .ZN(n10605) );
  NAND2_X1 U13142 ( .A1(n10606), .A2(n10605), .ZN(P1_U3293) );
  INV_X1 U13143 ( .A(n10607), .ZN(n10609) );
  NAND2_X1 U13144 ( .A1(n10609), .A2(n10608), .ZN(n10610) );
  AOI22_X1 U13145 ( .A1(n10617), .A2(n11981), .B1(n11985), .B2(n13786), .ZN(
        n10856) );
  OAI22_X1 U13146 ( .A1(n14646), .A2(n11935), .B1(n10612), .B2(n10140), .ZN(
        n10613) );
  XNOR2_X1 U13147 ( .A(n10613), .B(n11983), .ZN(n10854) );
  XNOR2_X1 U13148 ( .A(n10855), .B(n10854), .ZN(n10619) );
  NAND2_X1 U13149 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n13826) );
  OAI21_X1 U13150 ( .B1(n13763), .B2(n10614), .A(n13826), .ZN(n10616) );
  INV_X1 U13151 ( .A(n13785), .ZN(n10938) );
  OAI22_X1 U13152 ( .A1(n10636), .A2(n13765), .B1(n13766), .B2(n10938), .ZN(
        n10615) );
  AOI211_X1 U13153 ( .C1(n10617), .C2(n13769), .A(n10616), .B(n10615), .ZN(
        n10618) );
  OAI21_X1 U13154 ( .B1(n10619), .B2(n13771), .A(n10618), .ZN(P1_U3230) );
  INV_X1 U13155 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10698) );
  NOR2_X1 U13156 ( .A1(n15117), .A2(n10698), .ZN(n10620) );
  AOI21_X1 U13157 ( .B1(n15117), .B2(n10666), .A(n10620), .ZN(n10621) );
  OAI21_X1 U13158 ( .B1(n10622), .B2(n12900), .A(n10621), .ZN(P3_U3459) );
  OAI21_X1 U13159 ( .B1(n10625), .B2(n10624), .A(n10623), .ZN(n14644) );
  INV_X1 U13160 ( .A(n14644), .ZN(n10642) );
  INV_X1 U13161 ( .A(n14125), .ZN(n14114) );
  NOR2_X1 U13162 ( .A1(n14613), .A2(n9689), .ZN(n10630) );
  INV_X1 U13163 ( .A(n10626), .ZN(n10628) );
  OAI21_X1 U13164 ( .B1(n10628), .B2(n14640), .A(n10627), .ZN(n14641) );
  OAI22_X1 U13165 ( .A1(n14111), .A2(n14641), .B1(n13798), .B2(n14638), .ZN(
        n10629) );
  AOI211_X1 U13166 ( .C1(n14114), .C2(n10631), .A(n10630), .B(n10629), .ZN(
        n10641) );
  OAI21_X1 U13167 ( .B1(n10634), .B2(n10633), .A(n10632), .ZN(n10638) );
  OAI22_X1 U13168 ( .A1(n10636), .A2(n14102), .B1(n10635), .B2(n14078), .ZN(
        n10637) );
  AOI21_X1 U13169 ( .B1(n10638), .B2(n14245), .A(n10637), .ZN(n10639) );
  OAI21_X1 U13170 ( .B1(n10642), .B2(n14105), .A(n10639), .ZN(n14642) );
  NAND2_X1 U13171 ( .A1(n14642), .A2(n14613), .ZN(n10640) );
  OAI211_X1 U13172 ( .C1(n10642), .C2(n14117), .A(n10641), .B(n10640), .ZN(
        P1_U3291) );
  INV_X1 U13173 ( .A(n10643), .ZN(n11250) );
  XNOR2_X1 U13174 ( .A(n12111), .B(n10644), .ZN(n10733) );
  XNOR2_X1 U13175 ( .A(n10733), .B(n12445), .ZN(n10648) );
  OAI21_X1 U13176 ( .B1(n10648), .B2(n10647), .A(n10907), .ZN(n10649) );
  NAND2_X1 U13177 ( .A1(n10649), .A2(n12192), .ZN(n10654) );
  NOR2_X1 U13178 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10650), .ZN(n14903) );
  AOI21_X1 U13179 ( .B1(n12194), .B2(n12446), .A(n14903), .ZN(n10651) );
  OAI21_X1 U13180 ( .B1(n12201), .B2(n11251), .A(n10651), .ZN(n10652) );
  AOI21_X1 U13181 ( .B1(n10738), .B2(n12444), .A(n10652), .ZN(n10653) );
  OAI211_X1 U13182 ( .C1(n11250), .C2(n12181), .A(n10654), .B(n10653), .ZN(
        P3_U3167) );
  INV_X1 U13183 ( .A(P3_DATAO_REG_24__SCAN_IN), .ZN(n15217) );
  NAND2_X1 U13184 ( .A1(n12135), .A2(n12450), .ZN(n10655) );
  OAI21_X1 U13185 ( .B1(n12450), .B2(n15217), .A(n10655), .ZN(P3_U3515) );
  INV_X1 U13186 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10708) );
  OAI21_X1 U13187 ( .B1(n12402), .B2(n10656), .A(n12958), .ZN(n10657) );
  OAI21_X1 U13188 ( .B1(n12958), .B2(n10658), .A(n10657), .ZN(n10659) );
  INV_X1 U13189 ( .A(n10659), .ZN(n10660) );
  NAND2_X1 U13190 ( .A1(n10661), .A2(n10660), .ZN(n10663) );
  INV_X2 U13191 ( .A(n12826), .ZN(n15036) );
  INV_X1 U13192 ( .A(n15075), .ZN(n15056) );
  OR2_X1 U13193 ( .A1(n15100), .A2(n15056), .ZN(n10662) );
  NOR2_X2 U13194 ( .A1(n10663), .A2(n10662), .ZN(n15034) );
  AOI22_X1 U13195 ( .A1(n15034), .A2(n10665), .B1(n10664), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n10668) );
  NAND2_X1 U13196 ( .A1(n10666), .A2(n15036), .ZN(n10667) );
  OAI211_X1 U13197 ( .C1(n10708), .C2(n15036), .A(n10668), .B(n10667), .ZN(
        P3_U3233) );
  INV_X1 U13198 ( .A(n10669), .ZN(n10671) );
  OAI222_X1 U13199 ( .A1(n12258), .A2(P3_U3151), .B1(n14410), .B2(n10671), 
        .C1(n10670), .C2(n12973), .ZN(P3_U3274) );
  INV_X1 U13200 ( .A(n10672), .ZN(n10674) );
  OAI22_X1 U13201 ( .A1(n12424), .A2(P3_U3151), .B1(SI_22_), .B2(n12973), .ZN(
        n10673) );
  AOI21_X1 U13202 ( .B1(n10674), .B2(n12961), .A(n10673), .ZN(P3_U3273) );
  NAND2_X1 U13203 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n10682), .ZN(n10676) );
  NAND2_X1 U13204 ( .A1(n10676), .A2(n10675), .ZN(n10679) );
  MUX2_X1 U13205 ( .A(n11624), .B(P1_REG2_REG_14__SCAN_IN), .S(n11438), .Z(
        n10677) );
  INV_X1 U13206 ( .A(n10677), .ZN(n10678) );
  NAND2_X1 U13207 ( .A1(n10678), .A2(n10679), .ZN(n11439) );
  OAI211_X1 U13208 ( .C1(n10679), .C2(n10678), .A(n13873), .B(n11439), .ZN(
        n10691) );
  XNOR2_X1 U13209 ( .A(n11438), .B(n10680), .ZN(n10684) );
  NAND2_X1 U13210 ( .A1(n10684), .A2(n10683), .ZN(n11431) );
  OAI21_X1 U13211 ( .B1(n10684), .B2(n10683), .A(n11431), .ZN(n10689) );
  NAND2_X1 U13212 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n13631)
         );
  INV_X1 U13213 ( .A(n13631), .ZN(n10685) );
  AOI21_X1 U13214 ( .B1(n13817), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n10685), 
        .ZN(n10686) );
  OAI21_X1 U13215 ( .B1(n14598), .B2(n10687), .A(n10686), .ZN(n10688) );
  AOI21_X1 U13216 ( .B1(n10689), .B2(n14604), .A(n10688), .ZN(n10690) );
  NAND2_X1 U13217 ( .A1(n10691), .A2(n10690), .ZN(P1_U3257) );
  INV_X1 U13218 ( .A(n10694), .ZN(n10692) );
  NAND2_X1 U13219 ( .A1(n10692), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12427) );
  NAND2_X1 U13220 ( .A1(n10693), .A2(n12427), .ZN(n10704) );
  NAND2_X1 U13221 ( .A1(n10694), .A2(n12402), .ZN(n10695) );
  AND2_X1 U13222 ( .A1(n10696), .A2(n10695), .ZN(n10702) );
  AND2_X1 U13223 ( .A1(n10704), .A2(n10702), .ZN(n10707) );
  INV_X1 U13224 ( .A(n10707), .ZN(n10697) );
  MUX2_X1 U13225 ( .A(n12447), .B(n10697), .S(n12974), .Z(n14977) );
  INV_X1 U13226 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10713) );
  MUX2_X1 U13227 ( .A(n10713), .B(P3_REG1_REG_2__SCAN_IN), .S(n11476), .Z(
        n10701) );
  OR2_X1 U13228 ( .A1(n10698), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10839) );
  NOR2_X1 U13229 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10839), .ZN(n10699) );
  NAND2_X1 U13230 ( .A1(P3_REG1_REG_1__SCAN_IN), .A2(n10890), .ZN(n10889) );
  OAI21_X1 U13231 ( .B1(P3_IR_REG_1__SCAN_IN), .B2(n10839), .A(n10889), .ZN(
        n10700) );
  NAND2_X1 U13232 ( .A1(n10701), .A2(n10700), .ZN(n11475) );
  OAI21_X1 U13233 ( .B1(n10701), .B2(n10700), .A(n11475), .ZN(n10731) );
  INV_X1 U13234 ( .A(n10702), .ZN(n10703) );
  INV_X1 U13235 ( .A(n14982), .ZN(n15014) );
  OAI22_X1 U13236 ( .A1(n15014), .A2(n14311), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10705), .ZN(n10730) );
  INV_X1 U13237 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n15081) );
  NOR2_X1 U13238 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n10708), .ZN(n10841) );
  NAND2_X1 U13239 ( .A1(n8380), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10709) );
  INV_X1 U13240 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n15061) );
  AOI21_X1 U13241 ( .B1(n10712), .B2(n10711), .A(n11462), .ZN(n10728) );
  MUX2_X1 U13242 ( .A(n15061), .B(n10713), .S(n8844), .Z(n10714) );
  NAND2_X1 U13243 ( .A1(n10714), .A2(n11476), .ZN(n14855) );
  INV_X1 U13244 ( .A(n10714), .ZN(n10715) );
  NAND2_X1 U13245 ( .A1(n10715), .A2(n11463), .ZN(n10716) );
  AND2_X1 U13246 ( .A1(n14855), .A2(n10716), .ZN(n10724) );
  INV_X1 U13247 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10717) );
  MUX2_X1 U13248 ( .A(n15081), .B(n10717), .S(n8844), .Z(n10720) );
  NAND2_X1 U13249 ( .A1(n10720), .A2(n10718), .ZN(n10723) );
  INV_X1 U13250 ( .A(n10723), .ZN(n10719) );
  NOR2_X1 U13251 ( .A1(n10724), .A2(n10719), .ZN(n10726) );
  INV_X1 U13252 ( .A(n10720), .ZN(n10721) );
  NAND2_X1 U13253 ( .A1(n10721), .A2(n6913), .ZN(n10722) );
  AND2_X1 U13254 ( .A1(n10723), .A2(n10722), .ZN(n10892) );
  MUX2_X1 U13255 ( .A(n10708), .B(n10698), .S(n8844), .Z(n10836) );
  AND2_X1 U13256 ( .A1(n10836), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10893) );
  NAND2_X1 U13257 ( .A1(n10892), .A2(n10893), .ZN(n10891) );
  NAND2_X1 U13258 ( .A1(n10891), .A2(n10723), .ZN(n10725) );
  NAND2_X1 U13259 ( .A1(n10725), .A2(n10724), .ZN(n11487) );
  INV_X1 U13260 ( .A(n11487), .ZN(n14858) );
  AOI21_X1 U13261 ( .B1(n10726), .B2(n10891), .A(n14858), .ZN(n10727) );
  NAND2_X1 U13262 ( .A1(n12450), .A2(n12974), .ZN(n14999) );
  OAI22_X1 U13263 ( .A1(n15005), .A2(n10728), .B1(n10727), .B2(n14999), .ZN(
        n10729) );
  AOI211_X1 U13264 ( .C1(n14993), .C2(n10731), .A(n10730), .B(n10729), .ZN(
        n10732) );
  OAI21_X1 U13265 ( .B1(n11463), .B2(n14977), .A(n10732), .ZN(P3_U3184) );
  INV_X1 U13266 ( .A(n15026), .ZN(n10741) );
  NAND2_X1 U13267 ( .A1(n10733), .A2(n11116), .ZN(n10903) );
  AND2_X1 U13268 ( .A1(n10907), .A2(n10903), .ZN(n10735) );
  XNOR2_X1 U13269 ( .A(n12111), .B(n11123), .ZN(n10904) );
  XNOR2_X1 U13270 ( .A(n10904), .B(n11040), .ZN(n10734) );
  NAND2_X1 U13271 ( .A1(n10735), .A2(n10734), .ZN(n10881) );
  OAI211_X1 U13272 ( .C1(n10735), .C2(n10734), .A(n10881), .B(n12192), .ZN(
        n10740) );
  AND2_X1 U13273 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n14922) );
  AOI21_X1 U13274 ( .B1(n12194), .B2(n12445), .A(n14922), .ZN(n10736) );
  OAI21_X1 U13275 ( .B1(n12201), .B2(n11123), .A(n10736), .ZN(n10737) );
  AOI21_X1 U13276 ( .B1(n10738), .B2(n12443), .A(n10737), .ZN(n10739) );
  OAI211_X1 U13277 ( .C1(n10741), .C2(n12181), .A(n10740), .B(n10739), .ZN(
        P3_U3179) );
  NAND2_X1 U13278 ( .A1(n13105), .A2(n10035), .ZN(n10949) );
  AOI21_X1 U13279 ( .B1(n10745), .B2(n10744), .A(n6545), .ZN(n10753) );
  NAND2_X1 U13280 ( .A1(n13106), .A2(n14522), .ZN(n10747) );
  NAND2_X1 U13281 ( .A1(n13104), .A2(n14524), .ZN(n10746) );
  AND2_X1 U13282 ( .A1(n10747), .A2(n10746), .ZN(n10977) );
  INV_X1 U13283 ( .A(n10977), .ZN(n10748) );
  NAND2_X1 U13284 ( .A1(n14694), .A2(n10748), .ZN(n10749) );
  OAI211_X1 U13285 ( .C1(n14701), .C2(n10980), .A(n10750), .B(n10749), .ZN(
        n10751) );
  AOI21_X1 U13286 ( .B1(n14831), .B2(n14697), .A(n10751), .ZN(n10752) );
  OAI21_X1 U13287 ( .B1(n10753), .B2(n13073), .A(n10752), .ZN(P2_U3193) );
  NOR2_X1 U13288 ( .A1(n15075), .A2(n12258), .ZN(n15076) );
  OR2_X1 U13289 ( .A1(n15106), .A2(n15076), .ZN(n15015) );
  INV_X1 U13290 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n11488) );
  MUX2_X1 U13291 ( .A(n10754), .B(n11488), .S(n12826), .Z(n10758) );
  AOI22_X1 U13292 ( .A1(n15034), .A2(n10756), .B1(n10664), .B2(n10755), .ZN(
        n10757) );
  OAI211_X1 U13293 ( .C1(n10759), .C2(n12829), .A(n10758), .B(n10757), .ZN(
        P3_U3230) );
  INV_X1 U13294 ( .A(n13865), .ZN(n13858) );
  INV_X1 U13295 ( .A(n10760), .ZN(n10762) );
  OAI222_X1 U13296 ( .A1(n13858), .A2(P1_U3086), .B1(n14300), .B2(n10762), 
        .C1(n10761), .C2(n14298), .ZN(P1_U3337) );
  INV_X1 U13297 ( .A(n13152), .ZN(n13162) );
  OAI222_X1 U13298 ( .A1(n13614), .A2(n10763), .B1(n13605), .B2(n10762), .C1(
        P2_U3088), .C2(n13162), .ZN(P2_U3309) );
  OR2_X1 U13299 ( .A1(n14819), .A2(n13538), .ZN(n13440) );
  AOI22_X1 U13300 ( .A1(n14806), .A2(n10764), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n14808), .ZN(n10765) );
  OAI21_X1 U13301 ( .B1(n6896), .B2(n14812), .A(n10765), .ZN(n10766) );
  AOI21_X1 U13302 ( .B1(n14815), .B2(n10767), .A(n10766), .ZN(n10770) );
  MUX2_X1 U13303 ( .A(n10768), .B(n9624), .S(n6388), .Z(n10769) );
  OAI211_X1 U13304 ( .C1(n10771), .C2(n13440), .A(n10770), .B(n10769), .ZN(
        P2_U3263) );
  INV_X1 U13305 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15152) );
  OAI22_X1 U13306 ( .A1(n12900), .A2(n12280), .B1(n15117), .B2(n15152), .ZN(
        n10772) );
  AOI21_X1 U13307 ( .B1(n10773), .B2(n15117), .A(n10772), .ZN(n10774) );
  INV_X1 U13308 ( .A(n10774), .ZN(P3_U3463) );
  INV_X1 U13309 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10775) );
  OAI22_X1 U13310 ( .A1(n12900), .A2(n10776), .B1(n15117), .B2(n10775), .ZN(
        n10777) );
  AOI21_X1 U13311 ( .B1(n10778), .B2(n15117), .A(n10777), .ZN(n10779) );
  INV_X1 U13312 ( .A(n10779), .ZN(P3_U3462) );
  OR2_X1 U13313 ( .A1(n10785), .A2(n13106), .ZN(n10780) );
  INV_X1 U13314 ( .A(n10782), .ZN(n10974) );
  NAND2_X1 U13315 ( .A1(n14831), .A2(n13105), .ZN(n10783) );
  XNOR2_X1 U13316 ( .A(n11049), .B(n10792), .ZN(n10963) );
  INV_X1 U13317 ( .A(n10963), .ZN(n10798) );
  AND2_X1 U13318 ( .A1(n10785), .A2(n10784), .ZN(n10787) );
  OR2_X1 U13319 ( .A1(n10785), .A2(n10784), .ZN(n10786) );
  OAI21_X2 U13320 ( .B1(n10788), .B2(n10787), .A(n10786), .ZN(n10975) );
  NOR2_X1 U13321 ( .A1(n14831), .A2(n10790), .ZN(n10789) );
  NAND2_X1 U13322 ( .A1(n14831), .A2(n10790), .ZN(n10791) );
  INV_X1 U13323 ( .A(n10792), .ZN(n11048) );
  OAI211_X1 U13324 ( .C1(n6552), .C2(n10792), .A(n14520), .B(n11054), .ZN(
        n10793) );
  AOI22_X1 U13325 ( .A1(n14522), .A2(n13105), .B1(n13103), .B2(n14524), .ZN(
        n10956) );
  NAND2_X1 U13326 ( .A1(n10793), .A2(n10956), .ZN(n10961) );
  AOI211_X1 U13327 ( .C1(n11053), .C2(n10983), .A(n10035), .B(n11058), .ZN(
        n10962) );
  NAND2_X1 U13328 ( .A1(n10962), .A2(n14806), .ZN(n10795) );
  AOI22_X1 U13329 ( .A1(n14819), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n10958), 
        .B2(n14808), .ZN(n10794) );
  OAI211_X1 U13330 ( .C1(n7067), .C2(n14812), .A(n10795), .B(n10794), .ZN(
        n10796) );
  AOI21_X1 U13331 ( .B1(n10961), .B2(n13438), .A(n10796), .ZN(n10797) );
  OAI21_X1 U13332 ( .B1(n10798), .B2(n13434), .A(n10797), .ZN(P2_U3256) );
  INV_X1 U13333 ( .A(n10799), .ZN(n10800) );
  NAND2_X1 U13334 ( .A1(n10801), .A2(n10800), .ZN(n10803) );
  NAND2_X1 U13335 ( .A1(n10848), .A2(n10938), .ZN(n10802) );
  INV_X1 U13336 ( .A(n10936), .ZN(n10932) );
  OR2_X1 U13337 ( .A1(n14652), .A2(n13784), .ZN(n10804) );
  NAND2_X1 U13338 ( .A1(n10931), .A2(n10804), .ZN(n10805) );
  OAI21_X1 U13339 ( .B1(n10805), .B2(n10810), .A(n10822), .ZN(n10806) );
  INV_X1 U13340 ( .A(n10806), .ZN(n10930) );
  NAND2_X1 U13341 ( .A1(n11004), .A2(n10938), .ZN(n10807) );
  NAND2_X1 U13342 ( .A1(n10937), .A2(n10936), .ZN(n10935) );
  NAND2_X1 U13343 ( .A1(n14652), .A2(n11175), .ZN(n10809) );
  NAND2_X1 U13344 ( .A1(n10935), .A2(n10809), .ZN(n10812) );
  INV_X1 U13345 ( .A(n10810), .ZN(n10811) );
  NAND2_X1 U13346 ( .A1(n10812), .A2(n10811), .ZN(n10827) );
  OAI21_X1 U13347 ( .B1(n10812), .B2(n10811), .A(n10827), .ZN(n10815) );
  OAI22_X1 U13348 ( .A1(n11309), .A2(n14102), .B1(n11175), .B2(n14078), .ZN(
        n10814) );
  NOR2_X1 U13349 ( .A1(n10930), .A2(n14105), .ZN(n10813) );
  AOI211_X1 U13350 ( .C1(n14245), .C2(n10815), .A(n10814), .B(n10813), .ZN(
        n10923) );
  INV_X1 U13351 ( .A(n10943), .ZN(n10816) );
  INV_X1 U13352 ( .A(n11178), .ZN(n10925) );
  AOI21_X1 U13353 ( .B1(n11178), .B2(n10816), .A(n6546), .ZN(n10927) );
  AOI22_X1 U13354 ( .A1(n10927), .A2(n14654), .B1(n14653), .B2(n11178), .ZN(
        n10817) );
  OAI211_X1 U13355 ( .C1(n10930), .C2(n14658), .A(n10923), .B(n10817), .ZN(
        n10819) );
  NAND2_X1 U13356 ( .A1(n10819), .A2(n14687), .ZN(n10818) );
  OAI21_X1 U13357 ( .B1(n14687), .B2(n9708), .A(n10818), .ZN(P1_U3535) );
  INV_X1 U13358 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n15245) );
  NAND2_X1 U13359 ( .A1(n10819), .A2(n14679), .ZN(n10820) );
  OAI21_X1 U13360 ( .B1(n14679), .B2(n15245), .A(n10820), .ZN(P1_U3480) );
  OR2_X1 U13361 ( .A1(n11178), .A2(n13783), .ZN(n10821) );
  OAI21_X1 U13362 ( .B1(n6919), .B2(n10828), .A(n11016), .ZN(n14666) );
  OAI21_X1 U13363 ( .B1(n6810), .B2(n6546), .A(n11028), .ZN(n14663) );
  INV_X1 U13364 ( .A(n10824), .ZN(n11347) );
  AOI22_X1 U13365 ( .A1(n11348), .A2(n14114), .B1(n11347), .B2(n14089), .ZN(
        n10825) );
  OAI21_X1 U13366 ( .B1(n14663), .B2(n14111), .A(n10825), .ZN(n10834) );
  NAND2_X1 U13367 ( .A1(n11178), .A2(n11344), .ZN(n10826) );
  NAND2_X1 U13368 ( .A1(n10827), .A2(n10826), .ZN(n10829) );
  NAND2_X1 U13369 ( .A1(n10829), .A2(n10828), .ZN(n10830) );
  NAND3_X1 U13370 ( .A1(n11019), .A2(n14245), .A3(n10830), .ZN(n10832) );
  AOI22_X1 U13371 ( .A1(n14133), .A2(n13783), .B1(n14135), .B2(n13781), .ZN(
        n10831) );
  NAND2_X1 U13372 ( .A1(n10832), .A2(n10831), .ZN(n14664) );
  MUX2_X1 U13373 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n14664), .S(n14613), .Z(
        n10833) );
  AOI211_X1 U13374 ( .C1(n14621), .C2(n14666), .A(n10834), .B(n10833), .ZN(
        n10835) );
  INV_X1 U13375 ( .A(n10835), .ZN(P1_U3285) );
  INV_X1 U13376 ( .A(n14999), .ZN(n14859) );
  NOR3_X1 U13377 ( .A1(n14457), .A2(n14993), .A3(n14859), .ZN(n10845) );
  INV_X1 U13378 ( .A(n10893), .ZN(n10844) );
  OR2_X1 U13379 ( .A1(n14999), .A2(n10836), .ZN(n10837) );
  MUX2_X1 U13380 ( .A(n10837), .B(n14977), .S(P3_IR_REG_0__SCAN_IN), .Z(n10843) );
  INV_X1 U13381 ( .A(n14993), .ZN(n12572) );
  AOI22_X1 U13382 ( .A1(n14982), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n10838) );
  OAI21_X1 U13383 ( .B1(n12572), .B2(n10839), .A(n10838), .ZN(n10840) );
  AOI21_X1 U13384 ( .B1(n14457), .B2(n10841), .A(n10840), .ZN(n10842) );
  OAI211_X1 U13385 ( .C1(n10845), .C2(n10844), .A(n10843), .B(n10842), .ZN(
        P3_U3182) );
  MUX2_X1 U13386 ( .A(n10847), .B(n10846), .S(n14613), .Z(n10852) );
  OAI22_X1 U13387 ( .A1(n14125), .A2(n10848), .B1(n11002), .B2(n14638), .ZN(
        n10849) );
  AOI21_X1 U13388 ( .B1(n10850), .B2(n14146), .A(n10849), .ZN(n10851) );
  OAI211_X1 U13389 ( .C1(n10853), .C2(n14117), .A(n10852), .B(n10851), .ZN(
        P1_U3288) );
  INV_X1 U13390 ( .A(n10856), .ZN(n10857) );
  NAND2_X1 U13391 ( .A1(n10858), .A2(n10857), .ZN(n10859) );
  NAND2_X1 U13392 ( .A1(n11004), .A2(n11982), .ZN(n10862) );
  OR2_X1 U13393 ( .A1(n10140), .A2(n10938), .ZN(n10861) );
  NAND2_X1 U13394 ( .A1(n10862), .A2(n10861), .ZN(n10863) );
  XNOR2_X1 U13395 ( .A(n10863), .B(n11948), .ZN(n10870) );
  AOI22_X1 U13396 ( .A1(n11004), .A2(n11981), .B1(n11985), .B2(n13785), .ZN(
        n10869) );
  XNOR2_X1 U13397 ( .A(n10870), .B(n10869), .ZN(n10998) );
  INV_X1 U13398 ( .A(n10998), .ZN(n10864) );
  NAND2_X1 U13399 ( .A1(n14652), .A2(n6391), .ZN(n10866) );
  OR2_X1 U13400 ( .A1(n10140), .A2(n11175), .ZN(n10865) );
  NAND2_X1 U13401 ( .A1(n10866), .A2(n10865), .ZN(n10867) );
  XNOR2_X1 U13402 ( .A(n10867), .B(n11983), .ZN(n11164) );
  NOR2_X1 U13403 ( .A1(n10259), .A2(n11175), .ZN(n10868) );
  AOI21_X1 U13404 ( .B1(n14652), .B2(n11981), .A(n10868), .ZN(n11165) );
  XNOR2_X1 U13405 ( .A(n11164), .B(n11165), .ZN(n10873) );
  NAND2_X1 U13406 ( .A1(n10870), .A2(n10869), .ZN(n10874) );
  AND2_X1 U13407 ( .A1(n10873), .A2(n10874), .ZN(n10871) );
  NAND2_X1 U13408 ( .A1(n11168), .A2(n13757), .ZN(n10880) );
  AOI21_X1 U13409 ( .B1(n10872), .B2(n10874), .A(n10873), .ZN(n10879) );
  OAI22_X1 U13410 ( .A1(n13763), .A2(n10945), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10875), .ZN(n10877) );
  OAI22_X1 U13411 ( .A1(n10938), .A2(n13765), .B1(n13766), .B2(n11344), .ZN(
        n10876) );
  AOI211_X1 U13412 ( .C1(n14652), .C2(n13769), .A(n10877), .B(n10876), .ZN(
        n10878) );
  OAI21_X1 U13413 ( .B1(n10880), .B2(n10879), .A(n10878), .ZN(P1_U3239) );
  NAND2_X1 U13414 ( .A1(n10904), .A2(n12444), .ZN(n10908) );
  NAND2_X1 U13415 ( .A1(n10881), .A2(n10908), .ZN(n11228) );
  XNOR2_X1 U13416 ( .A(n7180), .B(n12111), .ZN(n10909) );
  XNOR2_X1 U13417 ( .A(n11228), .B(n10909), .ZN(n10888) );
  NOR2_X1 U13418 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10882), .ZN(n14942) );
  NOR2_X1 U13419 ( .A1(n12114), .A2(n11040), .ZN(n10883) );
  AOI211_X1 U13420 ( .C1(n10884), .C2(n12185), .A(n14942), .B(n10883), .ZN(
        n10885) );
  OAI21_X1 U13421 ( .B1(n11612), .B2(n12196), .A(n10885), .ZN(n10886) );
  AOI21_X1 U13422 ( .B1(n11387), .B2(n12198), .A(n10886), .ZN(n10887) );
  OAI21_X1 U13423 ( .B1(n10888), .B2(n12187), .A(n10887), .ZN(P3_U3153) );
  OAI21_X1 U13424 ( .B1(n10890), .B2(P3_REG1_REG_1__SCAN_IN), .A(n10889), .ZN(
        n10901) );
  OAI21_X1 U13425 ( .B1(n10893), .B2(n10892), .A(n10891), .ZN(n10894) );
  AOI22_X1 U13426 ( .A1(n14859), .A2(n10894), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(P3_U3151), .ZN(n10895) );
  OAI21_X1 U13427 ( .B1(n15014), .B2(n14309), .A(n10895), .ZN(n10900) );
  AOI21_X1 U13428 ( .B1(n10897), .B2(n15081), .A(n10896), .ZN(n10898) );
  NOR2_X1 U13429 ( .A1(n15005), .A2(n10898), .ZN(n10899) );
  AOI211_X1 U13430 ( .C1(n14993), .C2(n10901), .A(n10900), .B(n10899), .ZN(
        n10902) );
  OAI21_X1 U13431 ( .B1(n6913), .B2(n14977), .A(n10902), .ZN(P3_U3183) );
  XNOR2_X1 U13432 ( .A(n12111), .B(n12307), .ZN(n11074) );
  XNOR2_X1 U13433 ( .A(n11074), .B(n12306), .ZN(n10916) );
  OAI211_X1 U13434 ( .C1(n10904), .C2(n12444), .A(n10909), .B(n10903), .ZN(
        n10905) );
  NOR2_X1 U13435 ( .A1(n11230), .A2(n10905), .ZN(n10906) );
  OAI21_X1 U13436 ( .B1(n11230), .B2(n10908), .A(n10909), .ZN(n10912) );
  INV_X1 U13437 ( .A(n10909), .ZN(n11227) );
  OAI21_X1 U13438 ( .B1(n11230), .B2(n11231), .A(n11227), .ZN(n10911) );
  INV_X1 U13439 ( .A(n11077), .ZN(n10914) );
  AOI21_X1 U13440 ( .B1(n10916), .B2(n10915), .A(n10914), .ZN(n10922) );
  NOR2_X1 U13441 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10917), .ZN(n14981) );
  NOR2_X1 U13442 ( .A1(n12114), .A2(n11612), .ZN(n10918) );
  AOI211_X1 U13443 ( .C1(n12307), .C2(n12185), .A(n14981), .B(n10918), .ZN(
        n10919) );
  OAI21_X1 U13444 ( .B1(n12819), .B2(n12196), .A(n10919), .ZN(n10920) );
  AOI21_X1 U13445 ( .B1(n11616), .B2(n12198), .A(n10920), .ZN(n10921) );
  OAI21_X1 U13446 ( .B1(n10922), .B2(n12187), .A(n10921), .ZN(P3_U3171) );
  MUX2_X1 U13447 ( .A(n10924), .B(n10923), .S(n14613), .Z(n10929) );
  OAI22_X1 U13448 ( .A1(n10925), .A2(n14125), .B1(n11174), .B2(n14638), .ZN(
        n10926) );
  AOI21_X1 U13449 ( .B1(n10927), .B2(n14146), .A(n10926), .ZN(n10928) );
  OAI211_X1 U13450 ( .C1(n10930), .C2(n14117), .A(n10929), .B(n10928), .ZN(
        P1_U3286) );
  OAI21_X1 U13451 ( .B1(n10933), .B2(n10932), .A(n10931), .ZN(n10934) );
  INV_X1 U13452 ( .A(n10934), .ZN(n14659) );
  OAI21_X1 U13453 ( .B1(n10937), .B2(n10936), .A(n10935), .ZN(n10941) );
  OAI22_X1 U13454 ( .A1(n11344), .A2(n14102), .B1(n10938), .B2(n14078), .ZN(
        n10940) );
  NOR2_X1 U13455 ( .A1(n14659), .A2(n14105), .ZN(n10939) );
  AOI211_X1 U13456 ( .C1(n14245), .C2(n10941), .A(n10940), .B(n10939), .ZN(
        n14657) );
  MUX2_X1 U13457 ( .A(n10942), .B(n14657), .S(n14613), .Z(n10948) );
  AOI21_X1 U13458 ( .B1(n14652), .B2(n10944), .A(n10943), .ZN(n14655) );
  OAI22_X1 U13459 ( .A1(n7203), .A2(n14125), .B1(n10945), .B2(n14638), .ZN(
        n10946) );
  AOI21_X1 U13460 ( .B1(n14655), .B2(n14146), .A(n10946), .ZN(n10947) );
  OAI211_X1 U13461 ( .C1(n14659), .C2(n14117), .A(n10948), .B(n10947), .ZN(
        P1_U3287) );
  NAND2_X1 U13462 ( .A1(n10950), .A2(n10949), .ZN(n10951) );
  XNOR2_X1 U13463 ( .A(n11053), .B(n12995), .ZN(n11127) );
  NAND2_X1 U13464 ( .A1(n13104), .A2(n10035), .ZN(n11128) );
  XNOR2_X1 U13465 ( .A(n11127), .B(n11128), .ZN(n10952) );
  NOR3_X1 U13466 ( .A1(n6545), .A2(n7480), .A3(n10952), .ZN(n10954) );
  INV_X1 U13467 ( .A(n11131), .ZN(n10953) );
  OAI21_X1 U13468 ( .B1(n10954), .B2(n10953), .A(n14692), .ZN(n10960) );
  OAI21_X1 U13469 ( .B1(n13091), .B2(n10956), .A(n10955), .ZN(n10957) );
  AOI21_X1 U13470 ( .B1(n10958), .B2(n13093), .A(n10957), .ZN(n10959) );
  OAI211_X1 U13471 ( .C1(n7067), .C2(n13096), .A(n10960), .B(n10959), .ZN(
        P2_U3203) );
  AOI211_X1 U13472 ( .C1(n14845), .C2(n10963), .A(n10962), .B(n10961), .ZN(
        n10969) );
  AOI22_X1 U13473 ( .A1(n11053), .A2(n11748), .B1(n14850), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n10964) );
  OAI21_X1 U13474 ( .B1(n10969), .B2(n14850), .A(n10964), .ZN(P2_U3508) );
  INV_X1 U13475 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10965) );
  NOR2_X1 U13476 ( .A1(n14848), .A2(n10965), .ZN(n10966) );
  AOI21_X1 U13477 ( .B1(n11053), .B2(n10967), .A(n10966), .ZN(n10968) );
  OAI21_X1 U13478 ( .B1(n10969), .B2(n14846), .A(n10968), .ZN(P2_U3457) );
  NAND2_X1 U13479 ( .A1(n10970), .A2(n10974), .ZN(n10971) );
  NAND2_X1 U13480 ( .A1(n10972), .A2(n10971), .ZN(n14835) );
  OR2_X1 U13481 ( .A1(n6388), .A2(n10973), .ZN(n13419) );
  XNOR2_X1 U13482 ( .A(n10975), .B(n10974), .ZN(n10979) );
  OR2_X1 U13483 ( .A1(n14835), .A2(n10976), .ZN(n10978) );
  OAI211_X1 U13484 ( .C1(n13538), .C2(n10979), .A(n10978), .B(n10977), .ZN(
        n14837) );
  NAND2_X1 U13485 ( .A1(n14837), .A2(n13438), .ZN(n10988) );
  INV_X1 U13486 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10981) );
  OAI22_X1 U13487 ( .A1(n13438), .A2(n10981), .B1(n10980), .B2(n13407), .ZN(
        n10986) );
  AOI21_X1 U13488 ( .B1(n14831), .B2(n10982), .A(n10035), .ZN(n10984) );
  NAND2_X1 U13489 ( .A1(n10984), .A2(n10983), .ZN(n14833) );
  NOR2_X1 U13490 ( .A1(n14833), .A2(n13413), .ZN(n10985) );
  AOI211_X1 U13491 ( .C1(n14531), .C2(n14831), .A(n10986), .B(n10985), .ZN(
        n10987) );
  OAI211_X1 U13492 ( .C1(n14835), .C2(n13419), .A(n10988), .B(n10987), .ZN(
        P2_U3257) );
  NAND2_X1 U13493 ( .A1(n10989), .A2(n12961), .ZN(n10990) );
  OAI211_X1 U13494 ( .C1(n10991), .C2(n12973), .A(n10990), .B(n12427), .ZN(
        P3_U3272) );
  INV_X1 U13495 ( .A(n10992), .ZN(n10994) );
  OAI222_X1 U13496 ( .A1(P1_U3086), .A2(n9505), .B1(n14300), .B2(n10994), .C1(
        n10993), .C2(n14298), .ZN(P1_U3336) );
  OAI222_X1 U13497 ( .A1(n13614), .A2(n10995), .B1(n13605), .B2(n10994), .C1(
        P2_U3088), .C2(n13174), .ZN(P2_U3308) );
  INV_X1 U13498 ( .A(n10872), .ZN(n10996) );
  AOI21_X1 U13499 ( .B1(n10998), .B2(n10997), .A(n10996), .ZN(n11006) );
  AOI21_X1 U13500 ( .B1(n11000), .B2(n13753), .A(n10999), .ZN(n11001) );
  OAI21_X1 U13501 ( .B1(n11002), .B2(n13763), .A(n11001), .ZN(n11003) );
  AOI21_X1 U13502 ( .B1(n11004), .B2(n13769), .A(n11003), .ZN(n11005) );
  OAI21_X1 U13503 ( .B1(n11006), .B2(n13771), .A(n11005), .ZN(P1_U3227) );
  OAI22_X1 U13504 ( .A1(n14812), .A2(n11008), .B1(n11007), .B2(n13413), .ZN(
        n11012) );
  OAI21_X1 U13505 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(n13407), .A(n11009), .ZN(
        n11010) );
  MUX2_X1 U13506 ( .A(n11010), .B(P2_REG2_REG_3__SCAN_IN), .S(n14819), .Z(
        n11011) );
  AOI211_X1 U13507 ( .C1(n14815), .C2(n11013), .A(n11012), .B(n11011), .ZN(
        n11014) );
  INV_X1 U13508 ( .A(n11014), .ZN(P2_U3262) );
  OR2_X1 U13509 ( .A1(n11348), .A2(n13782), .ZN(n11015) );
  OAI21_X1 U13510 ( .B1(n11017), .B2(n11020), .A(n11222), .ZN(n11025) );
  INV_X1 U13511 ( .A(n11025), .ZN(n11108) );
  INV_X1 U13512 ( .A(n13780), .ZN(n11405) );
  OAI22_X1 U13513 ( .A1(n11405), .A2(n14102), .B1(n11309), .B2(n14078), .ZN(
        n11024) );
  OR2_X1 U13514 ( .A1(n11348), .A2(n11309), .ZN(n11018) );
  NAND2_X1 U13515 ( .A1(n11021), .A2(n11020), .ZN(n11022) );
  AOI21_X1 U13516 ( .B1(n11214), .B2(n11022), .A(n14672), .ZN(n11023) );
  AOI211_X1 U13517 ( .C1(n11323), .C2(n11025), .A(n11024), .B(n11023), .ZN(
        n11107) );
  MUX2_X1 U13518 ( .A(n11026), .B(n11107), .S(n14613), .Z(n11032) );
  INV_X1 U13519 ( .A(n14622), .ZN(n11027) );
  AOI21_X1 U13520 ( .B1(n11312), .B2(n11028), .A(n11027), .ZN(n11105) );
  INV_X1 U13521 ( .A(n11312), .ZN(n11029) );
  OAI22_X1 U13522 ( .A1(n11029), .A2(n14125), .B1(n11308), .B2(n14638), .ZN(
        n11030) );
  AOI21_X1 U13523 ( .B1(n11105), .B2(n14146), .A(n11030), .ZN(n11031) );
  OAI211_X1 U13524 ( .C1(n11108), .C2(n14117), .A(n11032), .B(n11031), .ZN(
        P1_U3284) );
  OAI21_X1 U13525 ( .B1(n11034), .B2(n12276), .A(n11033), .ZN(n11255) );
  INV_X1 U13526 ( .A(n11035), .ZN(n11036) );
  AOI21_X1 U13527 ( .B1(n12276), .B2(n11037), .A(n11036), .ZN(n11038) );
  OAI222_X1 U13528 ( .A1(n15044), .A2(n11040), .B1(n15046), .B2(n11039), .C1(
        n15072), .C2(n11038), .ZN(n11252) );
  AOI21_X1 U13529 ( .B1(n14490), .B2(n11255), .A(n11252), .ZN(n11047) );
  INV_X1 U13530 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n11041) );
  OAI22_X1 U13531 ( .A1(n11251), .A2(n12955), .B1(n15108), .B2(n11041), .ZN(
        n11042) );
  INV_X1 U13532 ( .A(n11042), .ZN(n11043) );
  OAI21_X1 U13533 ( .B1(n11047), .B2(n15110), .A(n11043), .ZN(P3_U3405) );
  INV_X1 U13534 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n11044) );
  OAI22_X1 U13535 ( .A1(n12900), .A2(n11251), .B1(n15117), .B2(n11044), .ZN(
        n11045) );
  INV_X1 U13536 ( .A(n11045), .ZN(n11046) );
  OAI21_X1 U13537 ( .B1(n11047), .B2(n15114), .A(n11046), .ZN(P3_U3464) );
  NAND2_X1 U13538 ( .A1(n11049), .A2(n11048), .ZN(n11051) );
  NAND2_X1 U13539 ( .A1(n11053), .A2(n13104), .ZN(n11050) );
  INV_X1 U13540 ( .A(n11206), .ZN(n11055) );
  XNOR2_X1 U13541 ( .A(n11207), .B(n11055), .ZN(n11157) );
  INV_X1 U13542 ( .A(n11157), .ZN(n11064) );
  INV_X1 U13543 ( .A(n13104), .ZN(n11052) );
  OAI211_X1 U13544 ( .C1(n11056), .C2(n11055), .A(n11198), .B(n14520), .ZN(
        n11057) );
  AOI22_X1 U13545 ( .A1(n14522), .A2(n13104), .B1(n14523), .B2(n14524), .ZN(
        n11141) );
  NAND2_X1 U13546 ( .A1(n11057), .A2(n11141), .ZN(n11155) );
  INV_X1 U13547 ( .A(n11208), .ZN(n11159) );
  INV_X1 U13548 ( .A(n11058), .ZN(n11059) );
  INV_X1 U13549 ( .A(n11201), .ZN(n11202) );
  AOI211_X1 U13550 ( .C1(n11208), .C2(n11059), .A(n10035), .B(n11202), .ZN(
        n11156) );
  NAND2_X1 U13551 ( .A1(n11156), .A2(n14806), .ZN(n11061) );
  AOI22_X1 U13552 ( .A1(n14819), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n11143), 
        .B2(n14808), .ZN(n11060) );
  OAI211_X1 U13553 ( .C1(n11159), .C2(n14812), .A(n11061), .B(n11060), .ZN(
        n11062) );
  AOI21_X1 U13554 ( .B1(n13438), .B2(n11155), .A(n11062), .ZN(n11063) );
  OAI21_X1 U13555 ( .B1(n13434), .B2(n11064), .A(n11063), .ZN(P2_U3255) );
  INV_X1 U13556 ( .A(n11065), .ZN(n11073) );
  INV_X1 U13557 ( .A(n11066), .ZN(n13077) );
  MUX2_X1 U13558 ( .A(n13077), .B(P2_REG2_REG_6__SCAN_IN), .S(n14819), .Z(
        n11070) );
  AOI22_X1 U13559 ( .A1(n14531), .A2(n13079), .B1(n14808), .B2(n13078), .ZN(
        n11067) );
  OAI21_X1 U13560 ( .B1(n13413), .B2(n11068), .A(n11067), .ZN(n11069) );
  AOI211_X1 U13561 ( .C1(n14815), .C2(n11071), .A(n11070), .B(n11069), .ZN(
        n11072) );
  OAI21_X1 U13562 ( .B1(n11073), .B2(n13440), .A(n11072), .ZN(P2_U3259) );
  INV_X1 U13563 ( .A(n11603), .ZN(n11084) );
  NAND2_X1 U13564 ( .A1(n11074), .A2(n12306), .ZN(n11075) );
  AND2_X1 U13565 ( .A1(n11077), .A2(n11075), .ZN(n11079) );
  XNOR2_X1 U13566 ( .A(n12111), .B(n11604), .ZN(n11372) );
  XNOR2_X1 U13567 ( .A(n11372), .B(n12440), .ZN(n11078) );
  AND2_X1 U13568 ( .A1(n11078), .A2(n11075), .ZN(n11076) );
  OAI211_X1 U13569 ( .C1(n11079), .C2(n11078), .A(n12192), .B(n11375), .ZN(
        n11083) );
  AND2_X1 U13570 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n14992) );
  AOI21_X1 U13571 ( .B1(n12194), .B2(n12441), .A(n14992), .ZN(n11080) );
  OAI21_X1 U13572 ( .B1(n14471), .B2(n12196), .A(n11080), .ZN(n11081) );
  AOI21_X1 U13573 ( .B1(n11604), .B2(n12185), .A(n11081), .ZN(n11082) );
  OAI211_X1 U13574 ( .C1(n11084), .C2(n12181), .A(n11083), .B(n11082), .ZN(
        P3_U3157) );
  NAND2_X1 U13575 ( .A1(n12447), .A2(P3_DATAO_REG_28__SCAN_IN), .ZN(n11085) );
  OAI21_X1 U13576 ( .B1(n12629), .B2(n12447), .A(n11085), .ZN(P3_U3519) );
  INV_X1 U13577 ( .A(n13440), .ZN(n13299) );
  NOR2_X1 U13578 ( .A1(n14815), .A2(n13299), .ZN(n11093) );
  OAI22_X1 U13579 ( .A1(n6388), .A2(n11087), .B1(n11086), .B2(n13407), .ZN(
        n11090) );
  NOR2_X1 U13580 ( .A1(n13413), .A2(n10035), .ZN(n11863) );
  INV_X1 U13581 ( .A(n11863), .ZN(n11669) );
  AOI21_X1 U13582 ( .B1(n11669), .B2(n14812), .A(n11088), .ZN(n11089) );
  AOI211_X1 U13583 ( .C1(n6388), .C2(P2_REG2_REG_0__SCAN_IN), .A(n11090), .B(
        n11089), .ZN(n11091) );
  OAI21_X1 U13584 ( .B1(n11093), .B2(n11092), .A(n11091), .ZN(P2_U3265) );
  INV_X1 U13585 ( .A(n11094), .ZN(n11095) );
  OAI22_X1 U13586 ( .A1(n13413), .A2(n11096), .B1(n11095), .B2(n13407), .ZN(
        n11099) );
  MUX2_X1 U13587 ( .A(n11097), .B(P2_REG2_REG_5__SCAN_IN), .S(n14819), .Z(
        n11098) );
  AOI211_X1 U13588 ( .C1(n14531), .C2(n11100), .A(n11099), .B(n11098), .ZN(
        n11103) );
  NAND2_X1 U13589 ( .A1(n11101), .A2(n13299), .ZN(n11102) );
  OAI211_X1 U13590 ( .C1(n11104), .C2(n13434), .A(n11103), .B(n11102), .ZN(
        P2_U3260) );
  AOI22_X1 U13591 ( .A1(n11105), .A2(n14654), .B1(n14653), .B2(n11312), .ZN(
        n11106) );
  OAI211_X1 U13592 ( .C1(n11108), .C2(n14658), .A(n11107), .B(n11106), .ZN(
        n11110) );
  NAND2_X1 U13593 ( .A1(n11110), .A2(n14687), .ZN(n11109) );
  OAI21_X1 U13594 ( .B1(n14687), .B2(n9778), .A(n11109), .ZN(P1_U3537) );
  INV_X1 U13595 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n15177) );
  NAND2_X1 U13596 ( .A1(n11110), .A2(n14679), .ZN(n11111) );
  OAI21_X1 U13597 ( .B1(n14679), .B2(n15177), .A(n11111), .ZN(P1_U3486) );
  OAI21_X1 U13598 ( .B1(n11113), .B2(n12226), .A(n11112), .ZN(n11114) );
  INV_X1 U13599 ( .A(n11114), .ZN(n15024) );
  AOI21_X1 U13600 ( .B1(n11115), .B2(n12226), .A(n15072), .ZN(n11119) );
  OAI22_X1 U13601 ( .A1(n11231), .A2(n15044), .B1(n11116), .B2(n15046), .ZN(
        n11117) );
  AOI21_X1 U13602 ( .B1(n11119), .B2(n11118), .A(n11117), .ZN(n15023) );
  OAI21_X1 U13603 ( .B1(n15024), .B2(n14494), .A(n15023), .ZN(n11125) );
  INV_X1 U13604 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n11120) );
  OAI22_X1 U13605 ( .A1(n11123), .A2(n12955), .B1(n15108), .B2(n11120), .ZN(
        n11121) );
  AOI21_X1 U13606 ( .B1(n11125), .B2(n15108), .A(n11121), .ZN(n11122) );
  INV_X1 U13607 ( .A(n11122), .ZN(P3_U3408) );
  INV_X1 U13608 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n11481) );
  OAI22_X1 U13609 ( .A1(n12900), .A2(n11123), .B1(n15117), .B2(n11481), .ZN(
        n11124) );
  AOI21_X1 U13610 ( .B1(n11125), .B2(n15117), .A(n11124), .ZN(n11126) );
  INV_X1 U13611 ( .A(n11126), .ZN(P3_U3465) );
  INV_X1 U13612 ( .A(n11127), .ZN(n11129) );
  NAND2_X1 U13613 ( .A1(n11129), .A2(n11128), .ZN(n11130) );
  XNOR2_X1 U13614 ( .A(n11208), .B(n12995), .ZN(n11132) );
  AND2_X1 U13615 ( .A1(n13103), .A2(n10035), .ZN(n11133) );
  NAND2_X1 U13616 ( .A1(n11132), .A2(n11133), .ZN(n11257) );
  INV_X1 U13617 ( .A(n11132), .ZN(n11135) );
  INV_X1 U13618 ( .A(n11133), .ZN(n11134) );
  NAND2_X1 U13619 ( .A1(n11135), .A2(n11134), .ZN(n11136) );
  NAND2_X1 U13620 ( .A1(n11257), .A2(n11136), .ZN(n11138) );
  AOI21_X1 U13621 ( .B1(n11137), .B2(n11138), .A(n13073), .ZN(n11139) );
  NAND2_X1 U13622 ( .A1(n11139), .A2(n11258), .ZN(n11145) );
  OAI21_X1 U13623 ( .B1(n13091), .B2(n11141), .A(n11140), .ZN(n11142) );
  AOI21_X1 U13624 ( .B1(n11143), .B2(n13093), .A(n11142), .ZN(n11144) );
  OAI211_X1 U13625 ( .C1(n11159), .C2(n13096), .A(n11145), .B(n11144), .ZN(
        P2_U3189) );
  NAND2_X1 U13626 ( .A1(n11146), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n11151) );
  NAND2_X1 U13627 ( .A1(n11147), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n11150) );
  NAND2_X1 U13628 ( .A1(n11148), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n11149) );
  AND3_X1 U13629 ( .A1(n11151), .A2(n11150), .A3(n11149), .ZN(n11152) );
  NAND2_X1 U13630 ( .A1(n12447), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(n11154) );
  OAI21_X1 U13631 ( .B1(n12602), .B2(n12447), .A(n11154), .ZN(P3_U3522) );
  AOI211_X1 U13632 ( .C1(n11157), .C2(n14845), .A(n11156), .B(n11155), .ZN(
        n11163) );
  INV_X1 U13633 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n11158) );
  OAI22_X1 U13634 ( .A1(n11159), .A2(n13584), .B1(n14848), .B2(n11158), .ZN(
        n11160) );
  INV_X1 U13635 ( .A(n11160), .ZN(n11161) );
  OAI21_X1 U13636 ( .B1(n11163), .B2(n14846), .A(n11161), .ZN(P2_U3460) );
  AOI22_X1 U13637 ( .A1(n11208), .A2(n11748), .B1(n14850), .B2(
        P2_REG1_REG_10__SCAN_IN), .ZN(n11162) );
  OAI21_X1 U13638 ( .B1(n11163), .B2(n14850), .A(n11162), .ZN(P2_U3509) );
  INV_X1 U13639 ( .A(n11164), .ZN(n11166) );
  OR2_X1 U13640 ( .A1(n11166), .A2(n11165), .ZN(n11167) );
  NAND2_X1 U13641 ( .A1(n11178), .A2(n11982), .ZN(n11170) );
  OR2_X1 U13642 ( .A1(n10140), .A2(n11344), .ZN(n11169) );
  NAND2_X1 U13643 ( .A1(n11170), .A2(n11169), .ZN(n11171) );
  XNOR2_X1 U13644 ( .A(n11171), .B(n11983), .ZN(n11290) );
  NOR2_X1 U13645 ( .A1(n10259), .A2(n11344), .ZN(n11172) );
  AOI21_X1 U13646 ( .B1(n11178), .B2(n11981), .A(n11172), .ZN(n11291) );
  XNOR2_X1 U13647 ( .A(n11290), .B(n11291), .ZN(n11288) );
  XNOR2_X1 U13648 ( .A(n11289), .B(n11288), .ZN(n11180) );
  OAI21_X1 U13649 ( .B1(n13763), .B2(n11174), .A(n11173), .ZN(n11177) );
  OAI22_X1 U13650 ( .A1(n11175), .A2(n13765), .B1(n13766), .B2(n11309), .ZN(
        n11176) );
  AOI211_X1 U13651 ( .C1(n11178), .C2(n13769), .A(n11177), .B(n11176), .ZN(
        n11179) );
  OAI21_X1 U13652 ( .B1(n11180), .B2(n13771), .A(n11179), .ZN(P1_U3213) );
  INV_X1 U13653 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11182) );
  MUX2_X1 U13654 ( .A(n11182), .B(P2_REG2_REG_13__SCAN_IN), .S(n11188), .Z(
        n14768) );
  NOR2_X1 U13655 ( .A1(n14767), .A2(n14768), .ZN(n14766) );
  XNOR2_X1 U13656 ( .A(n13124), .B(n13125), .ZN(n11184) );
  INV_X1 U13657 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n11183) );
  NOR2_X1 U13658 ( .A1(n11183), .A2(n11184), .ZN(n13126) );
  AOI211_X1 U13659 ( .C1(n11184), .C2(n11183), .A(n13126), .B(n14795), .ZN(
        n11195) );
  INV_X1 U13660 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11187) );
  MUX2_X1 U13661 ( .A(n11187), .B(P2_REG1_REG_13__SCAN_IN), .S(n11188), .Z(
        n14763) );
  INV_X1 U13662 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n11189) );
  MUX2_X1 U13663 ( .A(n11189), .B(P2_REG1_REG_14__SCAN_IN), .S(n13135), .Z(
        n11190) );
  AOI211_X1 U13664 ( .C1(n11191), .C2(n11190), .A(n13134), .B(n14791), .ZN(
        n11194) );
  NAND2_X1 U13665 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14512)
         );
  NAND2_X1 U13666 ( .A1(n14719), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n11192) );
  OAI211_X1 U13667 ( .C1(n14774), .C2(n13124), .A(n14512), .B(n11192), .ZN(
        n11193) );
  OR3_X1 U13668 ( .A1(n11195), .A2(n11194), .A3(n11193), .ZN(P2_U3228) );
  OR2_X1 U13669 ( .A1(n11208), .A2(n11196), .ZN(n11197) );
  OAI21_X1 U13670 ( .B1(n6556), .B2(n11210), .A(n14517), .ZN(n11200) );
  AOI22_X1 U13671 ( .A1(n14522), .A2(n13103), .B1(n13102), .B2(n14524), .ZN(
        n11262) );
  INV_X1 U13672 ( .A(n11262), .ZN(n11199) );
  AOI21_X1 U13673 ( .B1(n11200), .B2(n14520), .A(n11199), .ZN(n14840) );
  INV_X1 U13674 ( .A(n11359), .ZN(n14842) );
  OR2_X2 U13675 ( .A1(n11201), .A2(n11359), .ZN(n14534) );
  OAI211_X1 U13676 ( .C1(n11202), .C2(n14842), .A(n13390), .B(n14534), .ZN(
        n14839) );
  INV_X1 U13677 ( .A(n14839), .ZN(n11205) );
  AOI22_X1 U13678 ( .A1(n6388), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n11264), 
        .B2(n14808), .ZN(n11203) );
  OAI21_X1 U13679 ( .B1(n14842), .B2(n14812), .A(n11203), .ZN(n11204) );
  AOI21_X1 U13680 ( .B1(n11205), .B2(n14806), .A(n11204), .ZN(n11212) );
  NAND2_X1 U13681 ( .A1(n11208), .A2(n13103), .ZN(n11209) );
  XNOR2_X1 U13682 ( .A(n11356), .B(n11210), .ZN(n14844) );
  NAND2_X1 U13683 ( .A1(n14844), .A2(n14815), .ZN(n11211) );
  OAI211_X1 U13684 ( .C1(n14840), .C2(n6388), .A(n11212), .B(n11211), .ZN(
        P2_U3254) );
  NAND2_X1 U13685 ( .A1(n11312), .A2(n11407), .ZN(n11213) );
  OR2_X1 U13686 ( .A1(n14623), .A2(n11405), .ZN(n11216) );
  XOR2_X1 U13687 ( .A(n11224), .B(n11273), .Z(n11217) );
  INV_X1 U13688 ( .A(n13778), .ZN(n11882) );
  OAI22_X1 U13689 ( .A1(n11882), .A2(n14102), .B1(n11405), .B2(n14078), .ZN(
        n11687) );
  AOI21_X1 U13690 ( .B1(n11217), .B2(n14245), .A(n11687), .ZN(n11334) );
  INV_X1 U13691 ( .A(n14626), .ZN(n11219) );
  INV_X1 U13692 ( .A(n11692), .ZN(n11275) );
  INV_X1 U13693 ( .A(n11324), .ZN(n11218) );
  AOI21_X1 U13694 ( .B1(n11692), .B2(n11219), .A(n11218), .ZN(n11332) );
  NOR2_X1 U13695 ( .A1(n11275), .A2(n14125), .ZN(n11221) );
  OAI22_X1 U13696 ( .A1(n14613), .A2(n9172), .B1(n11690), .B2(n14638), .ZN(
        n11220) );
  AOI211_X1 U13697 ( .C1(n11332), .C2(n14146), .A(n11221), .B(n11220), .ZN(
        n11226) );
  OR2_X1 U13698 ( .A1(n14623), .A2(n13780), .ZN(n11223) );
  XNOR2_X1 U13699 ( .A(n11276), .B(n11224), .ZN(n11335) );
  OR2_X1 U13700 ( .A1(n11335), .A2(n14148), .ZN(n11225) );
  OAI211_X1 U13701 ( .C1(n11334), .C2(n14091), .A(n11226), .B(n11225), .ZN(
        P1_U3282) );
  MUX2_X1 U13702 ( .A(n11228), .B(n12443), .S(n11227), .Z(n11229) );
  XOR2_X1 U13703 ( .A(n11230), .B(n11229), .Z(n11236) );
  AND2_X1 U13704 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n14960) );
  NOR2_X1 U13705 ( .A1(n12114), .A2(n11231), .ZN(n11232) );
  AOI211_X1 U13706 ( .C1(n15018), .C2(n12185), .A(n14960), .B(n11232), .ZN(
        n11233) );
  OAI21_X1 U13707 ( .B1(n12306), .B2(n12196), .A(n11233), .ZN(n11234) );
  AOI21_X1 U13708 ( .B1(n15019), .B2(n12198), .A(n11234), .ZN(n11235) );
  OAI21_X1 U13709 ( .B1(n11236), .B2(n12187), .A(n11235), .ZN(P3_U3161) );
  OAI21_X1 U13710 ( .B1(n11238), .B2(n7180), .A(n11237), .ZN(n11393) );
  OAI211_X1 U13711 ( .C1(n11240), .C2(n12227), .A(n11239), .B(n15051), .ZN(
        n11242) );
  AOI22_X1 U13712 ( .A1(n12444), .A2(n15066), .B1(n15067), .B2(n12442), .ZN(
        n11241) );
  NAND2_X1 U13713 ( .A1(n11242), .A2(n11241), .ZN(n11390) );
  AOI21_X1 U13714 ( .B1(n14490), .B2(n11393), .A(n11390), .ZN(n11249) );
  INV_X1 U13715 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n11243) );
  OAI22_X1 U13716 ( .A1(n11389), .A2(n12955), .B1(n15108), .B2(n11243), .ZN(
        n11244) );
  INV_X1 U13717 ( .A(n11244), .ZN(n11245) );
  OAI21_X1 U13718 ( .B1(n11249), .B2(n15110), .A(n11245), .ZN(P3_U3411) );
  INV_X1 U13719 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n11246) );
  OAI22_X1 U13720 ( .A1(n12900), .A2(n11389), .B1(n15117), .B2(n11246), .ZN(
        n11247) );
  INV_X1 U13721 ( .A(n11247), .ZN(n11248) );
  OAI21_X1 U13722 ( .B1(n11249), .B2(n15114), .A(n11248), .ZN(P3_U3466) );
  OAI22_X1 U13723 ( .A1(n12824), .A2(n11251), .B1(n11250), .B2(n12822), .ZN(
        n11254) );
  MUX2_X1 U13724 ( .A(P3_REG2_REG_5__SCAN_IN), .B(n11252), .S(n15036), .Z(
        n11253) );
  AOI211_X1 U13725 ( .C1(n14476), .C2(n11255), .A(n11254), .B(n11253), .ZN(
        n11256) );
  INV_X1 U13726 ( .A(n11256), .ZN(P3_U3228) );
  XNOR2_X1 U13727 ( .A(n11359), .B(n12995), .ZN(n11415) );
  NAND2_X1 U13728 ( .A1(n14523), .A2(n10035), .ZN(n11413) );
  XNOR2_X1 U13729 ( .A(n11415), .B(n11413), .ZN(n11259) );
  OAI211_X1 U13730 ( .C1(n11260), .C2(n11259), .A(n11416), .B(n14692), .ZN(
        n11266) );
  OAI22_X1 U13731 ( .A1(n13091), .A2(n11262), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11261), .ZN(n11263) );
  AOI21_X1 U13732 ( .B1(n11264), .B2(n13093), .A(n11263), .ZN(n11265) );
  OAI211_X1 U13733 ( .C1(n14842), .C2(n13096), .A(n11266), .B(n11265), .ZN(
        P2_U3208) );
  INV_X1 U13734 ( .A(n11267), .ZN(n11271) );
  INV_X1 U13735 ( .A(n11268), .ZN(n11270) );
  OAI222_X1 U13736 ( .A1(P3_U3151), .A2(n11271), .B1(n14410), .B2(n11270), 
        .C1(n11269), .C2(n12973), .ZN(P3_U3271) );
  NAND2_X1 U13737 ( .A1(n11692), .A2(n13667), .ZN(n11272) );
  OR2_X1 U13738 ( .A1(n11692), .A2(n13667), .ZN(n11274) );
  INV_X1 U13739 ( .A(n11550), .ZN(n11543) );
  XNOR2_X1 U13740 ( .A(n11544), .B(n11543), .ZN(n14566) );
  INV_X1 U13741 ( .A(n14128), .ZN(n14633) );
  NAND2_X1 U13742 ( .A1(n11276), .A2(n13667), .ZN(n11277) );
  OR2_X1 U13743 ( .A1(n13661), .A2(n13778), .ZN(n11280) );
  XNOR2_X1 U13744 ( .A(n11551), .B(n11550), .ZN(n14568) );
  NAND2_X1 U13745 ( .A1(n14568), .A2(n14621), .ZN(n11287) );
  AOI21_X1 U13746 ( .B1(n14562), .B2(n6550), .A(n6825), .ZN(n14563) );
  NAND2_X1 U13747 ( .A1(n14562), .A2(n14114), .ZN(n11283) );
  OAI22_X1 U13748 ( .A1(n13764), .A2(n14102), .B1(n11882), .B2(n14078), .ZN(
        n14561) );
  INV_X1 U13749 ( .A(n13727), .ZN(n11281) );
  AOI22_X1 U13750 ( .A1(n14613), .A2(n14561), .B1(n14089), .B2(n11281), .ZN(
        n11282) );
  OAI211_X1 U13751 ( .C1(n14613), .C2(n11284), .A(n11283), .B(n11282), .ZN(
        n11285) );
  AOI21_X1 U13752 ( .B1(n14563), .B2(n14146), .A(n11285), .ZN(n11286) );
  OAI211_X1 U13753 ( .C1(n14566), .C2(n14633), .A(n11287), .B(n11286), .ZN(
        P1_U3280) );
  INV_X1 U13754 ( .A(n11290), .ZN(n11292) );
  OR2_X1 U13755 ( .A1(n11292), .A2(n11291), .ZN(n11293) );
  NAND2_X1 U13756 ( .A1(n11348), .A2(n11982), .ZN(n11295) );
  OR2_X1 U13757 ( .A1(n10140), .A2(n11309), .ZN(n11294) );
  NAND2_X1 U13758 ( .A1(n11295), .A2(n11294), .ZN(n11296) );
  XNOR2_X1 U13759 ( .A(n11296), .B(n11948), .ZN(n11303) );
  NOR2_X1 U13760 ( .A1(n10259), .A2(n11309), .ZN(n11297) );
  AOI21_X1 U13761 ( .B1(n11348), .B2(n11981), .A(n11297), .ZN(n11302) );
  XNOR2_X1 U13762 ( .A(n11303), .B(n11302), .ZN(n11343) );
  NAND2_X1 U13763 ( .A1(n11312), .A2(n11982), .ZN(n11299) );
  OR2_X1 U13764 ( .A1(n10140), .A2(n11407), .ZN(n11298) );
  NAND2_X1 U13765 ( .A1(n11299), .A2(n11298), .ZN(n11300) );
  XNOR2_X1 U13766 ( .A(n11300), .B(n11983), .ZN(n11398) );
  NOR2_X1 U13767 ( .A1(n10259), .A2(n11407), .ZN(n11301) );
  AOI21_X1 U13768 ( .B1(n11312), .B2(n11981), .A(n11301), .ZN(n11399) );
  XNOR2_X1 U13769 ( .A(n11398), .B(n11399), .ZN(n11305) );
  NAND2_X1 U13770 ( .A1(n11303), .A2(n11302), .ZN(n11306) );
  AND2_X1 U13771 ( .A1(n11305), .A2(n11306), .ZN(n11304) );
  NAND2_X1 U13772 ( .A1(n11401), .A2(n13757), .ZN(n11315) );
  AOI21_X1 U13773 ( .B1(n11340), .B2(n11306), .A(n11305), .ZN(n11314) );
  OAI21_X1 U13774 ( .B1(n13763), .B2(n11308), .A(n11307), .ZN(n11311) );
  OAI22_X1 U13775 ( .A1(n11309), .A2(n13765), .B1(n13766), .B2(n11405), .ZN(
        n11310) );
  AOI211_X1 U13776 ( .C1(n11312), .C2(n13769), .A(n11311), .B(n11310), .ZN(
        n11313) );
  OAI21_X1 U13777 ( .B1(n11315), .B2(n11314), .A(n11313), .ZN(P1_U3231) );
  XNOR2_X1 U13778 ( .A(n11316), .B(n11317), .ZN(n14431) );
  XNOR2_X1 U13779 ( .A(n11318), .B(n11317), .ZN(n11319) );
  NAND2_X1 U13780 ( .A1(n11319), .A2(n14245), .ZN(n11321) );
  AOI22_X1 U13781 ( .A1(n14133), .A2(n13779), .B1(n14135), .B2(n13777), .ZN(
        n11320) );
  NAND2_X1 U13782 ( .A1(n11321), .A2(n11320), .ZN(n11322) );
  AOI21_X1 U13783 ( .B1(n14431), .B2(n11323), .A(n11322), .ZN(n14433) );
  NAND2_X1 U13784 ( .A1(n13661), .A2(n11324), .ZN(n11325) );
  NAND2_X1 U13785 ( .A1(n6550), .A2(n11325), .ZN(n14429) );
  OAI22_X1 U13786 ( .A1(n14613), .A2(n11326), .B1(n13665), .B2(n14638), .ZN(
        n11327) );
  AOI21_X1 U13787 ( .B1(n13661), .B2(n14114), .A(n11327), .ZN(n11328) );
  OAI21_X1 U13788 ( .B1(n14429), .B2(n14111), .A(n11328), .ZN(n11329) );
  AOI21_X1 U13789 ( .B1(n14431), .B2(n11837), .A(n11329), .ZN(n11330) );
  OAI21_X1 U13790 ( .B1(n14433), .B2(n14091), .A(n11330), .ZN(P1_U3281) );
  INV_X1 U13791 ( .A(n11331), .ZN(n11353) );
  OAI222_X1 U13792 ( .A1(n13605), .A2(n11353), .B1(n7505), .B2(P2_U3088), .C1(
        n7123), .C2(n13614), .ZN(P2_U3307) );
  AOI22_X1 U13793 ( .A1(n11332), .A2(n14654), .B1(n14653), .B2(n11692), .ZN(
        n11333) );
  OAI211_X1 U13794 ( .C1(n14257), .C2(n11335), .A(n11334), .B(n11333), .ZN(
        n11337) );
  NAND2_X1 U13795 ( .A1(n11337), .A2(n14687), .ZN(n11336) );
  OAI21_X1 U13796 ( .B1(n14687), .B2(n10064), .A(n11336), .ZN(P1_U3539) );
  INV_X1 U13797 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n11339) );
  NAND2_X1 U13798 ( .A1(n11337), .A2(n14679), .ZN(n11338) );
  OAI21_X1 U13799 ( .B1(n14679), .B2(n11339), .A(n11338), .ZN(P1_U3492) );
  INV_X1 U13800 ( .A(n11340), .ZN(n11341) );
  AOI21_X1 U13801 ( .B1(n11343), .B2(n11342), .A(n11341), .ZN(n11351) );
  OAI22_X1 U13802 ( .A1(n11344), .A2(n13765), .B1(n13766), .B2(n11407), .ZN(
        n11345) );
  AOI211_X1 U13803 ( .C1(n13711), .C2(n11347), .A(n11346), .B(n11345), .ZN(
        n11350) );
  NAND2_X1 U13804 ( .A1(n11348), .A2(n13769), .ZN(n11349) );
  OAI211_X1 U13805 ( .C1(n11351), .C2(n13771), .A(n11350), .B(n11349), .ZN(
        P1_U3221) );
  OAI222_X1 U13806 ( .A1(n11354), .A2(P1_U3086), .B1(n14300), .B2(n11353), 
        .C1(n11352), .C2(n14298), .ZN(P1_U3335) );
  AND2_X1 U13807 ( .A1(n11359), .A2(n14523), .ZN(n11355) );
  NOR2_X1 U13808 ( .A1(n14696), .A2(n13102), .ZN(n11357) );
  XNOR2_X1 U13809 ( .A(n11633), .B(n11362), .ZN(n14549) );
  INV_X1 U13810 ( .A(n14549), .ZN(n11371) );
  AND2_X1 U13811 ( .A1(n11359), .A2(n11358), .ZN(n14515) );
  NOR2_X1 U13812 ( .A1(n14532), .A2(n14515), .ZN(n11360) );
  OAI211_X1 U13813 ( .C1(n11363), .C2(n11362), .A(n11638), .B(n14520), .ZN(
        n11366) );
  INV_X1 U13814 ( .A(n14522), .ZN(n13059) );
  OAI22_X1 U13815 ( .A1(n11654), .A2(n13067), .B1(n11364), .B2(n13059), .ZN(
        n11422) );
  INV_X1 U13816 ( .A(n11422), .ZN(n11365) );
  NAND2_X1 U13817 ( .A1(n11366), .A2(n11365), .ZN(n14547) );
  OAI211_X1 U13818 ( .C1(n14546), .C2(n7071), .A(n13390), .B(n11644), .ZN(
        n14545) );
  AOI22_X1 U13819 ( .A1(n6388), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n11421), 
        .B2(n14808), .ZN(n11368) );
  NAND2_X1 U13820 ( .A1(n11636), .A2(n14531), .ZN(n11367) );
  OAI211_X1 U13821 ( .C1(n14545), .C2(n13413), .A(n11368), .B(n11367), .ZN(
        n11369) );
  AOI21_X1 U13822 ( .B1(n14547), .B2(n13438), .A(n11369), .ZN(n11370) );
  OAI21_X1 U13823 ( .B1(n11371), .B2(n13434), .A(n11370), .ZN(P2_U3252) );
  INV_X1 U13824 ( .A(n11372), .ZN(n11373) );
  NAND2_X1 U13825 ( .A1(n11373), .A2(n12440), .ZN(n11374) );
  INV_X1 U13826 ( .A(n14493), .ZN(n11376) );
  XNOR2_X1 U13827 ( .A(n12111), .B(n11376), .ZN(n11377) );
  INV_X1 U13828 ( .A(n11455), .ZN(n11379) );
  AOI21_X1 U13829 ( .B1(n12439), .B2(n11380), .A(n11379), .ZN(n11386) );
  INV_X1 U13830 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11381) );
  NOR2_X1 U13831 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11381), .ZN(n11533) );
  NOR2_X1 U13832 ( .A1(n12196), .A2(n12820), .ZN(n11382) );
  AOI211_X1 U13833 ( .C1(n12194), .C2(n12440), .A(n11533), .B(n11382), .ZN(
        n11383) );
  OAI21_X1 U13834 ( .B1(n12201), .B2(n14493), .A(n11383), .ZN(n11384) );
  AOI21_X1 U13835 ( .B1(n12821), .B2(n12198), .A(n11384), .ZN(n11385) );
  OAI21_X1 U13836 ( .B1(n11386), .B2(n12187), .A(n11385), .ZN(P3_U3176) );
  INV_X1 U13837 ( .A(n11387), .ZN(n11388) );
  OAI22_X1 U13838 ( .A1(n12824), .A2(n11389), .B1(n11388), .B2(n12822), .ZN(
        n11392) );
  MUX2_X1 U13839 ( .A(n11390), .B(P3_REG2_REG_7__SCAN_IN), .S(n12826), .Z(
        n11391) );
  AOI211_X1 U13840 ( .C1(n14476), .C2(n11393), .A(n11392), .B(n11391), .ZN(
        n11394) );
  INV_X1 U13841 ( .A(n11394), .ZN(P3_U3226) );
  INV_X1 U13842 ( .A(n11395), .ZN(n11564) );
  OAI222_X1 U13843 ( .A1(n13614), .A2(n11397), .B1(n13605), .B2(n11564), .C1(
        P2_U3088), .C2(n11396), .ZN(P2_U3306) );
  INV_X1 U13844 ( .A(n11398), .ZN(n11400) );
  NAND2_X1 U13845 ( .A1(n14623), .A2(n11982), .ZN(n11403) );
  OR2_X1 U13846 ( .A1(n10140), .A2(n11405), .ZN(n11402) );
  NAND2_X1 U13847 ( .A1(n11403), .A2(n11402), .ZN(n11404) );
  XNOR2_X1 U13848 ( .A(n11404), .B(n11983), .ZN(n11679) );
  NOR2_X1 U13849 ( .A1(n10259), .A2(n11405), .ZN(n11406) );
  AOI21_X1 U13850 ( .B1(n14623), .B2(n11981), .A(n11406), .ZN(n11680) );
  XNOR2_X1 U13851 ( .A(n11679), .B(n11680), .ZN(n11677) );
  XNOR2_X1 U13852 ( .A(n11678), .B(n11677), .ZN(n11412) );
  NOR2_X1 U13853 ( .A1(n13763), .A2(n14637), .ZN(n11410) );
  NOR2_X1 U13854 ( .A1(n11407), .A2(n14078), .ZN(n14609) );
  NOR2_X1 U13855 ( .A1(n13667), .A2(n14102), .ZN(n14627) );
  NOR2_X1 U13856 ( .A1(n14609), .A2(n14627), .ZN(n14668) );
  INV_X1 U13857 ( .A(n13753), .ZN(n13709) );
  OAI22_X1 U13858 ( .A1(n14668), .A2(n13709), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11408), .ZN(n11409) );
  AOI211_X1 U13859 ( .C1(n14623), .C2(n13769), .A(n11410), .B(n11409), .ZN(
        n11411) );
  OAI21_X1 U13860 ( .B1(n11412), .B2(n13771), .A(n11411), .ZN(P1_U3217) );
  INV_X1 U13861 ( .A(n11413), .ZN(n11414) );
  XNOR2_X1 U13862 ( .A(n14696), .B(n12048), .ZN(n11417) );
  NAND2_X1 U13863 ( .A1(n13102), .A2(n10035), .ZN(n11418) );
  NAND2_X1 U13864 ( .A1(n11417), .A2(n11418), .ZN(n14689) );
  INV_X1 U13865 ( .A(n11417), .ZN(n11420) );
  INV_X1 U13866 ( .A(n11418), .ZN(n11419) );
  NAND2_X1 U13867 ( .A1(n11420), .A2(n11419), .ZN(n14688) );
  XNOR2_X1 U13868 ( .A(n11636), .B(n12995), .ZN(n11795) );
  NAND2_X1 U13869 ( .A1(n14525), .A2(n10035), .ZN(n11793) );
  XNOR2_X1 U13870 ( .A(n11795), .B(n11793), .ZN(n11791) );
  XNOR2_X1 U13871 ( .A(n11792), .B(n11791), .ZN(n11427) );
  INV_X1 U13872 ( .A(n11421), .ZN(n11424) );
  AOI22_X1 U13873 ( .A1(n14694), .A2(n11422), .B1(P2_REG3_REG_13__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11423) );
  OAI21_X1 U13874 ( .B1(n11424), .B2(n14701), .A(n11423), .ZN(n11425) );
  AOI21_X1 U13875 ( .B1(n11636), .B2(n14697), .A(n11425), .ZN(n11426) );
  OAI21_X1 U13876 ( .B1(n11427), .B2(n13073), .A(n11426), .ZN(P2_U3206) );
  INV_X1 U13877 ( .A(n14598), .ZN(n13852) );
  INV_X1 U13878 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n11430) );
  NOR2_X1 U13879 ( .A1(n11428), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13688) );
  INV_X1 U13880 ( .A(n13688), .ZN(n11429) );
  OAI21_X1 U13881 ( .B1(n14607), .B2(n11430), .A(n11429), .ZN(n11437) );
  OAI21_X1 U13882 ( .B1(n11438), .B2(P1_REG1_REG_14__SCAN_IN), .A(n11431), 
        .ZN(n11432) );
  NAND2_X1 U13883 ( .A1(n14599), .A2(n11432), .ZN(n11433) );
  NAND2_X1 U13884 ( .A1(n11433), .A2(n14593), .ZN(n11435) );
  XNOR2_X1 U13885 ( .A(n11760), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n11434) );
  NOR2_X1 U13886 ( .A1(n11434), .A2(n11435), .ZN(n11759) );
  AOI211_X1 U13887 ( .C1(n11435), .C2(n11434), .A(n11759), .B(n13847), .ZN(
        n11436) );
  AOI211_X1 U13888 ( .C1(n13852), .C2(n11760), .A(n11437), .B(n11436), .ZN(
        n11449) );
  NAND2_X1 U13889 ( .A1(n11438), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11440) );
  NAND2_X1 U13890 ( .A1(n11440), .A2(n11439), .ZN(n11441) );
  NOR2_X1 U13891 ( .A1(n11442), .A2(n11441), .ZN(n11443) );
  XNOR2_X1 U13892 ( .A(n11442), .B(n11441), .ZN(n14597) );
  NOR2_X1 U13893 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14597), .ZN(n14596) );
  NOR2_X1 U13894 ( .A1(n11443), .A2(n14596), .ZN(n11447) );
  INV_X1 U13895 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11445) );
  NOR2_X1 U13896 ( .A1(n11444), .A2(n11445), .ZN(n11751) );
  AOI21_X1 U13897 ( .B1(n11445), .B2(n11444), .A(n11751), .ZN(n11446) );
  NAND2_X1 U13898 ( .A1(n11446), .A2(n11447), .ZN(n11752) );
  OAI211_X1 U13899 ( .C1(n11447), .C2(n11446), .A(n13873), .B(n11752), .ZN(
        n11448) );
  NAND2_X1 U13900 ( .A1(n11449), .A2(n11448), .ZN(P1_U3259) );
  INV_X1 U13901 ( .A(n11450), .ZN(n11451) );
  OAI222_X1 U13902 ( .A1(n11453), .A2(P3_U3151), .B1(n12973), .B2(n11452), 
        .C1(n14410), .C2(n11451), .ZN(P3_U3270) );
  XNOR2_X1 U13903 ( .A(n12089), .B(n14486), .ZN(n11585) );
  XNOR2_X1 U13904 ( .A(n11585), .B(n12801), .ZN(n11456) );
  XNOR2_X1 U13905 ( .A(n11584), .B(n11456), .ZN(n11461) );
  NAND2_X1 U13906 ( .A1(n12198), .A2(n14477), .ZN(n11458) );
  AND2_X1 U13907 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n11715) );
  AOI21_X1 U13908 ( .B1(n12194), .B2(n12439), .A(n11715), .ZN(n11457) );
  OAI211_X1 U13909 ( .C1(n14470), .C2(n12196), .A(n11458), .B(n11457), .ZN(
        n11459) );
  AOI21_X1 U13910 ( .B1(n14486), .B2(n12185), .A(n11459), .ZN(n11460) );
  OAI21_X1 U13911 ( .B1(n11461), .B2(n12187), .A(n11460), .ZN(P3_U3164) );
  NOR2_X1 U13912 ( .A1(n11489), .A2(n11464), .ZN(n11465) );
  INV_X1 U13913 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n15039) );
  AOI22_X1 U13914 ( .A1(P3_REG2_REG_4__SCAN_IN), .A2(n11494), .B1(n14880), 
        .B2(n15039), .ZN(n14872) );
  NOR2_X1 U13915 ( .A1(n11499), .A2(n11466), .ZN(n11467) );
  INV_X1 U13916 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n14893) );
  NOR2_X1 U13917 ( .A1(n14893), .A2(n14892), .ZN(n14891) );
  INV_X1 U13918 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n15029) );
  AOI22_X1 U13919 ( .A1(P3_REG2_REG_6__SCAN_IN), .A2(n11504), .B1(n14919), 
        .B2(n15029), .ZN(n14911) );
  NOR2_X1 U13920 ( .A1(n11509), .A2(n11468), .ZN(n11469) );
  INV_X1 U13921 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n14932) );
  NOR2_X1 U13922 ( .A1(n14932), .A2(n14931), .ZN(n14930) );
  INV_X1 U13923 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n15022) );
  AOI22_X1 U13924 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n11514), .B1(n14957), 
        .B2(n15022), .ZN(n14949) );
  NOR2_X1 U13925 ( .A1(n11520), .A2(n11470), .ZN(n11471) );
  INV_X1 U13926 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n14970) );
  NOR2_X1 U13927 ( .A1(n14970), .A2(n14969), .ZN(n14968) );
  INV_X1 U13928 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11606) );
  AOI22_X1 U13929 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n15009), .B1(n14414), 
        .B2(n11606), .ZN(n15003) );
  OAI21_X1 U13930 ( .B1(n11472), .B2(n11700), .A(n11695), .ZN(n11474) );
  INV_X1 U13931 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11473) );
  NOR2_X1 U13932 ( .A1(n11473), .A2(n11474), .ZN(n11696) );
  AOI21_X1 U13933 ( .B1(n11474), .B2(n11473), .A(n11696), .ZN(n11539) );
  INV_X1 U13934 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n15115) );
  AOI22_X1 U13935 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n14414), .B1(n15009), 
        .B2(n15115), .ZN(n14991) );
  INV_X1 U13936 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n11575) );
  AOI22_X1 U13937 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n14957), .B1(n11514), 
        .B2(n11575), .ZN(n14962) );
  AOI22_X1 U13938 ( .A1(P3_REG1_REG_6__SCAN_IN), .A2(n14919), .B1(n11504), 
        .B2(n11481), .ZN(n14924) );
  AOI22_X1 U13939 ( .A1(P3_REG1_REG_4__SCAN_IN), .A2(n14880), .B1(n11494), 
        .B2(n15152), .ZN(n14885) );
  NAND2_X1 U13940 ( .A1(n14863), .A2(n11477), .ZN(n11478) );
  NAND2_X1 U13941 ( .A1(P3_REG1_REG_3__SCAN_IN), .A2(n14867), .ZN(n14866) );
  NAND2_X1 U13942 ( .A1(n11478), .A2(n14866), .ZN(n14886) );
  NAND2_X1 U13943 ( .A1(n14900), .A2(n11479), .ZN(n11480) );
  XNOR2_X1 U13944 ( .A(n11499), .B(n11479), .ZN(n14905) );
  NAND2_X1 U13945 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(n14905), .ZN(n14904) );
  NAND2_X1 U13946 ( .A1(n11480), .A2(n14904), .ZN(n14925) );
  NAND2_X1 U13947 ( .A1(n14924), .A2(n14925), .ZN(n14923) );
  NAND2_X1 U13948 ( .A1(n14939), .A2(n11482), .ZN(n11483) );
  NAND2_X1 U13949 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n14944), .ZN(n14943) );
  NAND2_X1 U13950 ( .A1(n11483), .A2(n14943), .ZN(n14963) );
  NAND2_X1 U13951 ( .A1(n14962), .A2(n14963), .ZN(n14961) );
  NAND2_X1 U13952 ( .A1(n14978), .A2(n11484), .ZN(n11485) );
  NAND2_X1 U13953 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n14984), .ZN(n14983) );
  NAND2_X1 U13954 ( .A1(n11485), .A2(n14983), .ZN(n14990) );
  INV_X1 U13955 ( .A(n11700), .ZN(n11707) );
  XNOR2_X1 U13956 ( .A(n11701), .B(n11707), .ZN(n11486) );
  NAND2_X1 U13957 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n11486), .ZN(n11702) );
  OAI21_X1 U13958 ( .B1(n11486), .B2(P3_REG1_REG_11__SCAN_IN), .A(n11702), 
        .ZN(n11537) );
  NAND2_X1 U13959 ( .A1(n11487), .A2(n14855), .ZN(n11493) );
  MUX2_X1 U13960 ( .A(n11488), .B(n10775), .S(n12559), .Z(n11490) );
  NAND2_X1 U13961 ( .A1(n11490), .A2(n11489), .ZN(n14874) );
  INV_X1 U13962 ( .A(n11490), .ZN(n11491) );
  NAND2_X1 U13963 ( .A1(n11491), .A2(n14863), .ZN(n11492) );
  AND2_X1 U13964 ( .A1(n14874), .A2(n11492), .ZN(n14856) );
  NAND2_X1 U13965 ( .A1(n11493), .A2(n14856), .ZN(n14878) );
  NAND2_X1 U13966 ( .A1(n14878), .A2(n14874), .ZN(n11498) );
  MUX2_X1 U13967 ( .A(n15039), .B(n15152), .S(n12559), .Z(n11495) );
  NAND2_X1 U13968 ( .A1(n11495), .A2(n11494), .ZN(n14894) );
  INV_X1 U13969 ( .A(n11495), .ZN(n11496) );
  NAND2_X1 U13970 ( .A1(n11496), .A2(n14880), .ZN(n11497) );
  AND2_X1 U13971 ( .A1(n14894), .A2(n11497), .ZN(n14876) );
  NAND2_X1 U13972 ( .A1(n11498), .A2(n14876), .ZN(n14898) );
  NAND2_X1 U13973 ( .A1(n14898), .A2(n14894), .ZN(n11503) );
  MUX2_X1 U13974 ( .A(n14893), .B(n11044), .S(n12559), .Z(n11500) );
  NAND2_X1 U13975 ( .A1(n11500), .A2(n11499), .ZN(n14913) );
  INV_X1 U13976 ( .A(n11500), .ZN(n11501) );
  NAND2_X1 U13977 ( .A1(n11501), .A2(n14900), .ZN(n11502) );
  AND2_X1 U13978 ( .A1(n14913), .A2(n11502), .ZN(n14896) );
  NAND2_X1 U13979 ( .A1(n11503), .A2(n14896), .ZN(n14917) );
  NAND2_X1 U13980 ( .A1(n14917), .A2(n14913), .ZN(n11508) );
  MUX2_X1 U13981 ( .A(n15029), .B(n11481), .S(n12559), .Z(n11505) );
  NAND2_X1 U13982 ( .A1(n11505), .A2(n11504), .ZN(n14933) );
  INV_X1 U13983 ( .A(n11505), .ZN(n11506) );
  NAND2_X1 U13984 ( .A1(n11506), .A2(n14919), .ZN(n11507) );
  AND2_X1 U13985 ( .A1(n14933), .A2(n11507), .ZN(n14915) );
  NAND2_X1 U13986 ( .A1(n11508), .A2(n14915), .ZN(n14937) );
  NAND2_X1 U13987 ( .A1(n14937), .A2(n14933), .ZN(n11513) );
  MUX2_X1 U13988 ( .A(n14932), .B(n11246), .S(n12559), .Z(n11510) );
  NAND2_X1 U13989 ( .A1(n11510), .A2(n11509), .ZN(n14951) );
  INV_X1 U13990 ( .A(n11510), .ZN(n11511) );
  NAND2_X1 U13991 ( .A1(n11511), .A2(n14939), .ZN(n11512) );
  AND2_X1 U13992 ( .A1(n14951), .A2(n11512), .ZN(n14935) );
  NAND2_X1 U13993 ( .A1(n11513), .A2(n14935), .ZN(n14955) );
  NAND2_X1 U13994 ( .A1(n14955), .A2(n14951), .ZN(n11518) );
  MUX2_X1 U13995 ( .A(n15022), .B(n11575), .S(n12559), .Z(n11515) );
  NAND2_X1 U13996 ( .A1(n11515), .A2(n11514), .ZN(n14971) );
  INV_X1 U13997 ( .A(n11515), .ZN(n11516) );
  NAND2_X1 U13998 ( .A1(n11516), .A2(n14957), .ZN(n11517) );
  AND2_X1 U13999 ( .A1(n14971), .A2(n11517), .ZN(n14953) );
  NAND2_X1 U14000 ( .A1(n11518), .A2(n14953), .ZN(n14975) );
  NAND2_X1 U14001 ( .A1(n14975), .A2(n14971), .ZN(n11524) );
  INV_X1 U14002 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11519) );
  MUX2_X1 U14003 ( .A(n14970), .B(n11519), .S(n12559), .Z(n11521) );
  NAND2_X1 U14004 ( .A1(n11521), .A2(n11520), .ZN(n14997) );
  INV_X1 U14005 ( .A(n11521), .ZN(n11522) );
  NAND2_X1 U14006 ( .A1(n11522), .A2(n14978), .ZN(n11523) );
  AND2_X1 U14007 ( .A1(n14997), .A2(n11523), .ZN(n14973) );
  NAND2_X1 U14008 ( .A1(n11524), .A2(n14973), .ZN(n14998) );
  NAND2_X1 U14009 ( .A1(n14998), .A2(n14997), .ZN(n11528) );
  MUX2_X1 U14010 ( .A(n11606), .B(n15115), .S(n12559), .Z(n11525) );
  NAND2_X1 U14011 ( .A1(n11525), .A2(n15009), .ZN(n11529) );
  INV_X1 U14012 ( .A(n11525), .ZN(n11526) );
  NAND2_X1 U14013 ( .A1(n11526), .A2(n14414), .ZN(n11527) );
  AND2_X1 U14014 ( .A1(n11529), .A2(n11527), .ZN(n14995) );
  NAND2_X1 U14015 ( .A1(n11528), .A2(n14995), .ZN(n15001) );
  NAND2_X1 U14016 ( .A1(n15001), .A2(n11529), .ZN(n11531) );
  MUX2_X1 U14017 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12559), .Z(n11706) );
  XNOR2_X1 U14018 ( .A(n11706), .B(n11707), .ZN(n11530) );
  NAND2_X1 U14019 ( .A1(n11531), .A2(n11530), .ZN(n11712) );
  OAI21_X1 U14020 ( .B1(n11531), .B2(n11530), .A(n11712), .ZN(n11532) );
  NAND2_X1 U14021 ( .A1(n11532), .A2(n14859), .ZN(n11535) );
  AOI21_X1 U14022 ( .B1(n14982), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n11533), 
        .ZN(n11534) );
  OAI211_X1 U14023 ( .C1(n14977), .C2(n11700), .A(n11535), .B(n11534), .ZN(
        n11536) );
  AOI21_X1 U14024 ( .B1(n11537), .B2(n14993), .A(n11536), .ZN(n11538) );
  OAI21_X1 U14025 ( .B1(n11539), .B2(n15005), .A(n11538), .ZN(P3_U3193) );
  AOI222_X1 U14026 ( .A1(n11541), .A2(n13594), .B1(P1_DATAO_REG_22__SCAN_IN), 
        .B2(n13602), .C1(P2_STATE_REG_SCAN_IN), .C2(n11540), .ZN(n11542) );
  INV_X1 U14027 ( .A(n11542), .ZN(P2_U3305) );
  OR2_X1 U14028 ( .A1(n14562), .A2(n13666), .ZN(n11545) );
  XNOR2_X1 U14029 ( .A(n11724), .B(n11547), .ZN(n11621) );
  NAND2_X1 U14030 ( .A1(n13634), .A2(n11548), .ZN(n11549) );
  NAND2_X1 U14031 ( .A1(n11733), .A2(n11549), .ZN(n11625) );
  NAND2_X1 U14032 ( .A1(n11554), .A2(n11553), .ZN(n11628) );
  NAND3_X1 U14033 ( .A1(n11730), .A2(n11628), .A3(n14677), .ZN(n11558) );
  OR2_X1 U14034 ( .A1(n14102), .A2(n13686), .ZN(n11556) );
  OR2_X1 U14035 ( .A1(n14078), .A2(n13666), .ZN(n11555) );
  NAND2_X1 U14036 ( .A1(n11556), .A2(n11555), .ZN(n13629) );
  AOI21_X1 U14037 ( .B1(n13634), .B2(n14653), .A(n13629), .ZN(n11557) );
  OAI211_X1 U14038 ( .C1(n14662), .C2(n11625), .A(n11558), .B(n11557), .ZN(
        n11559) );
  AOI21_X1 U14039 ( .B1(n14245), .B2(n11621), .A(n11559), .ZN(n11562) );
  NAND2_X1 U14040 ( .A1(n14678), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n11560) );
  OAI21_X1 U14041 ( .B1(n11562), .B2(n14678), .A(n11560), .ZN(P1_U3501) );
  NAND2_X1 U14042 ( .A1(n14685), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n11561) );
  OAI21_X1 U14043 ( .B1(n11562), .B2(n14685), .A(n11561), .ZN(P1_U3542) );
  OAI222_X1 U14044 ( .A1(P1_U3086), .A2(n8999), .B1(n14300), .B2(n11564), .C1(
        n11563), .C2(n14298), .ZN(P1_U3334) );
  OAI21_X1 U14045 ( .B1(n11566), .B2(n12297), .A(n11565), .ZN(n11567) );
  INV_X1 U14046 ( .A(n11567), .ZN(n15017) );
  OAI21_X1 U14047 ( .B1(n11570), .B2(n11569), .A(n11568), .ZN(n11571) );
  AOI222_X1 U14048 ( .A1(n15051), .A2(n11571), .B1(n12443), .B2(n15066), .C1(
        n12441), .C2(n15067), .ZN(n15016) );
  OAI21_X1 U14049 ( .B1(n14494), .B2(n15017), .A(n15016), .ZN(n11577) );
  INV_X1 U14050 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n11572) );
  OAI22_X1 U14051 ( .A1(n12299), .A2(n12955), .B1(n15108), .B2(n11572), .ZN(
        n11573) );
  AOI21_X1 U14052 ( .B1(n11577), .B2(n15108), .A(n11573), .ZN(n11574) );
  INV_X1 U14053 ( .A(n11574), .ZN(P3_U3414) );
  OAI22_X1 U14054 ( .A1(n12900), .A2(n12299), .B1(n15117), .B2(n11575), .ZN(
        n11576) );
  AOI21_X1 U14055 ( .B1(n11577), .B2(n15117), .A(n11576), .ZN(n11578) );
  INV_X1 U14056 ( .A(n11578), .ZN(P3_U3467) );
  INV_X1 U14057 ( .A(n11579), .ZN(n11583) );
  INV_X1 U14058 ( .A(n11580), .ZN(n11581) );
  OAI222_X1 U14059 ( .A1(n11583), .A2(P3_U3151), .B1(n12973), .B2(n11582), 
        .C1(n14410), .C2(n11581), .ZN(P3_U3269) );
  INV_X1 U14060 ( .A(n11585), .ZN(n11586) );
  NAND2_X1 U14061 ( .A1(n11586), .A2(n12820), .ZN(n11587) );
  XNOR2_X1 U14062 ( .A(n14484), .B(n12111), .ZN(n11773) );
  XNOR2_X1 U14063 ( .A(n11773), .B(n14470), .ZN(n11588) );
  XNOR2_X1 U14064 ( .A(n11775), .B(n11588), .ZN(n11595) );
  INV_X1 U14065 ( .A(n11589), .ZN(n12804) );
  NOR2_X1 U14066 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11590), .ZN(n12464) );
  NOR2_X1 U14067 ( .A1(n12196), .A2(n12778), .ZN(n11591) );
  AOI211_X1 U14068 ( .C1(n12194), .C2(n12801), .A(n12464), .B(n11591), .ZN(
        n11592) );
  OAI21_X1 U14069 ( .B1(n12804), .B2(n12181), .A(n11592), .ZN(n11593) );
  AOI21_X1 U14070 ( .B1(n14484), .B2(n12185), .A(n11593), .ZN(n11594) );
  OAI21_X1 U14071 ( .B1(n11595), .B2(n12187), .A(n11594), .ZN(P3_U3174) );
  OAI211_X1 U14072 ( .C1(n11597), .C2(n12313), .A(n11596), .B(n15051), .ZN(
        n11599) );
  AOI22_X1 U14073 ( .A1(n15067), .A2(n12439), .B1(n12441), .B2(n15066), .ZN(
        n11598) );
  NAND2_X1 U14074 ( .A1(n11599), .A2(n11598), .ZN(n15105) );
  INV_X1 U14075 ( .A(n15105), .ZN(n11609) );
  INV_X1 U14076 ( .A(n11600), .ZN(n11601) );
  AOI21_X1 U14077 ( .B1(n12313), .B2(n11602), .A(n11601), .ZN(n15107) );
  AOI22_X1 U14078 ( .A1(n15034), .A2(n11604), .B1(n10664), .B2(n11603), .ZN(
        n11605) );
  OAI21_X1 U14079 ( .B1(n11606), .B2(n15036), .A(n11605), .ZN(n11607) );
  AOI21_X1 U14080 ( .B1(n15107), .B2(n14476), .A(n11607), .ZN(n11608) );
  OAI21_X1 U14081 ( .B1(n12826), .B2(n11609), .A(n11608), .ZN(P3_U3223) );
  XNOR2_X1 U14082 ( .A(n11610), .B(n12303), .ZN(n15097) );
  AOI21_X1 U14083 ( .B1(n11611), .B2(n12303), .A(n15072), .ZN(n11615) );
  OAI22_X1 U14084 ( .A1(n11612), .A2(n15046), .B1(n12819), .B2(n15044), .ZN(
        n11613) );
  AOI21_X1 U14085 ( .B1(n11615), .B2(n11614), .A(n11613), .ZN(n15094) );
  AOI22_X1 U14086 ( .A1(n15034), .A2(n12307), .B1(n10664), .B2(n11616), .ZN(
        n11618) );
  OR2_X1 U14087 ( .A1(n15036), .A2(n14970), .ZN(n11617) );
  OAI211_X1 U14088 ( .C1(n15094), .C2(n12826), .A(n11618), .B(n11617), .ZN(
        n11619) );
  AOI21_X1 U14089 ( .B1(n14476), .B2(n15097), .A(n11619), .ZN(n11620) );
  INV_X1 U14090 ( .A(n11620), .ZN(P3_U3224) );
  INV_X1 U14091 ( .A(n11621), .ZN(n11631) );
  INV_X1 U14092 ( .A(n13632), .ZN(n11622) );
  AOI22_X1 U14093 ( .A1(n14613), .A2(n13629), .B1(n14089), .B2(n11622), .ZN(
        n11623) );
  OAI21_X1 U14094 ( .B1(n11624), .B2(n14613), .A(n11623), .ZN(n11627) );
  NOR2_X1 U14095 ( .A1(n11625), .A2(n14111), .ZN(n11626) );
  AOI211_X1 U14096 ( .C1(n14114), .C2(n13634), .A(n11627), .B(n11626), .ZN(
        n11630) );
  NAND3_X1 U14097 ( .A1(n11730), .A2(n11628), .A3(n14621), .ZN(n11629) );
  OAI211_X1 U14098 ( .C1(n11631), .C2(n14633), .A(n11630), .B(n11629), .ZN(
        P1_U3279) );
  OR2_X1 U14099 ( .A1(n11636), .A2(n14525), .ZN(n11632) );
  NAND2_X1 U14100 ( .A1(n11633), .A2(n11632), .ZN(n11635) );
  NAND2_X1 U14101 ( .A1(n11636), .A2(n14525), .ZN(n11634) );
  XOR2_X1 U14102 ( .A(n11664), .B(n11663), .Z(n11743) );
  INV_X1 U14103 ( .A(n11743), .ZN(n11650) );
  OR2_X1 U14104 ( .A1(n11636), .A2(n11641), .ZN(n11637) );
  NAND2_X1 U14105 ( .A1(n11638), .A2(n11637), .ZN(n11640) );
  AOI21_X1 U14106 ( .B1(n11663), .B2(n11640), .A(n11639), .ZN(n11643) );
  OAI22_X1 U14107 ( .A1(n11826), .A2(n13067), .B1(n11641), .B2(n13059), .ZN(
        n14510) );
  INV_X1 U14108 ( .A(n14510), .ZN(n11642) );
  OAI21_X1 U14109 ( .B1(n11643), .B2(n13538), .A(n11642), .ZN(n11741) );
  AOI211_X1 U14110 ( .C1(n14511), .C2(n11644), .A(n10035), .B(n11667), .ZN(
        n11742) );
  NAND2_X1 U14111 ( .A1(n11742), .A2(n14806), .ZN(n11647) );
  AOI22_X1 U14112 ( .A1(n14819), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n11645), 
        .B2(n14808), .ZN(n11646) );
  OAI211_X1 U14113 ( .C1(n11745), .C2(n14812), .A(n11647), .B(n11646), .ZN(
        n11648) );
  AOI21_X1 U14114 ( .B1(n11741), .B2(n13438), .A(n11648), .ZN(n11649) );
  OAI21_X1 U14115 ( .B1(n11650), .B2(n13434), .A(n11649), .ZN(P2_U3251) );
  INV_X1 U14116 ( .A(n11651), .ZN(n11653) );
  OAI222_X1 U14117 ( .A1(n8844), .A2(P3_U3151), .B1(n14410), .B2(n11653), .C1(
        n11652), .C2(n12973), .ZN(P3_U3268) );
  INV_X1 U14118 ( .A(n11804), .ZN(n11662) );
  NAND2_X1 U14119 ( .A1(n14511), .A2(n11654), .ZN(n11655) );
  NAND2_X1 U14120 ( .A1(n11658), .A2(n11657), .ZN(n11659) );
  NAND3_X1 U14121 ( .A1(n11822), .A2(n14520), .A3(n11659), .ZN(n11661) );
  AND2_X1 U14122 ( .A1(n13101), .A2(n14522), .ZN(n11660) );
  AOI21_X1 U14123 ( .B1(n13099), .B2(n14524), .A(n11660), .ZN(n11806) );
  NAND2_X1 U14124 ( .A1(n11661), .A2(n11806), .ZN(n14542) );
  AOI21_X1 U14125 ( .B1(n11662), .B2(n14808), .A(n14542), .ZN(n11672) );
  NAND2_X1 U14126 ( .A1(n11664), .A2(n11663), .ZN(n11666) );
  NAND2_X1 U14127 ( .A1(n14511), .A2(n13101), .ZN(n11665) );
  XNOR2_X1 U14128 ( .A(n11825), .B(n11824), .ZN(n14544) );
  OAI21_X1 U14129 ( .B1(n14540), .B2(n11667), .A(n13423), .ZN(n14541) );
  AOI22_X1 U14130 ( .A1(n11809), .A2(n14531), .B1(P2_REG2_REG_15__SCAN_IN), 
        .B2(n14819), .ZN(n11668) );
  OAI21_X1 U14131 ( .B1(n14541), .B2(n11669), .A(n11668), .ZN(n11670) );
  AOI21_X1 U14132 ( .B1(n14544), .B2(n14815), .A(n11670), .ZN(n11671) );
  OAI21_X1 U14133 ( .B1(n11672), .B2(n6388), .A(n11671), .ZN(P2_U3250) );
  NAND2_X1 U14134 ( .A1(n11692), .A2(n6391), .ZN(n11674) );
  OR2_X1 U14135 ( .A1(n10140), .A2(n13667), .ZN(n11673) );
  NAND2_X1 U14136 ( .A1(n11674), .A2(n11673), .ZN(n11675) );
  XNOR2_X1 U14137 ( .A(n11675), .B(n11948), .ZN(n11876) );
  NOR2_X1 U14138 ( .A1(n10259), .A2(n13667), .ZN(n11676) );
  AOI21_X1 U14139 ( .B1(n11692), .B2(n11981), .A(n11676), .ZN(n11875) );
  XNOR2_X1 U14140 ( .A(n11876), .B(n11875), .ZN(n11686) );
  INV_X1 U14141 ( .A(n11679), .ZN(n11681) );
  INV_X1 U14142 ( .A(n11878), .ZN(n11684) );
  AOI21_X1 U14143 ( .B1(n11686), .B2(n11685), .A(n11684), .ZN(n11694) );
  NAND2_X1 U14144 ( .A1(n11687), .A2(n13753), .ZN(n11688) );
  OAI211_X1 U14145 ( .C1(n13763), .C2(n11690), .A(n11689), .B(n11688), .ZN(
        n11691) );
  AOI21_X1 U14146 ( .B1(n11692), .B2(n13769), .A(n11691), .ZN(n11693) );
  OAI21_X1 U14147 ( .B1(n11694), .B2(n13771), .A(n11693), .ZN(P1_U3236) );
  INV_X1 U14148 ( .A(n11695), .ZN(n11697) );
  INV_X1 U14149 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n14479) );
  AOI22_X1 U14150 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n12454), .B1(n12456), 
        .B2(n14479), .ZN(n11698) );
  AOI21_X1 U14151 ( .B1(n11699), .B2(n11698), .A(n12451), .ZN(n11721) );
  INV_X1 U14152 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14492) );
  AOI22_X1 U14153 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n12456), .B1(n12454), 
        .B2(n14492), .ZN(n11705) );
  NAND2_X1 U14154 ( .A1(n11701), .A2(n11700), .ZN(n11703) );
  NAND2_X1 U14155 ( .A1(n11703), .A2(n11702), .ZN(n11704) );
  NAND2_X1 U14156 ( .A1(n11705), .A2(n11704), .ZN(n12453) );
  OAI21_X1 U14157 ( .B1(n11705), .B2(n11704), .A(n12453), .ZN(n11719) );
  MUX2_X1 U14158 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12559), .Z(n12457) );
  XNOR2_X1 U14159 ( .A(n12457), .B(n12454), .ZN(n11710) );
  INV_X1 U14160 ( .A(n11706), .ZN(n11708) );
  NAND2_X1 U14161 ( .A1(n11708), .A2(n11707), .ZN(n11711) );
  AND2_X1 U14162 ( .A1(n11710), .A2(n11711), .ZN(n11709) );
  NAND2_X1 U14163 ( .A1(n11712), .A2(n11709), .ZN(n12461) );
  INV_X1 U14164 ( .A(n12461), .ZN(n11714) );
  AOI21_X1 U14165 ( .B1(n11712), .B2(n11711), .A(n11710), .ZN(n11713) );
  NOR3_X1 U14166 ( .A1(n11714), .A2(n11713), .A3(n14999), .ZN(n11718) );
  AOI21_X1 U14167 ( .B1(n14982), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n11715), 
        .ZN(n11716) );
  OAI21_X1 U14168 ( .B1(n14977), .B2(n12456), .A(n11716), .ZN(n11717) );
  AOI211_X1 U14169 ( .C1(n11719), .C2(n14993), .A(n11718), .B(n11717), .ZN(
        n11720) );
  OAI21_X1 U14170 ( .B1(n11721), .B2(n15005), .A(n11720), .ZN(P3_U3194) );
  INV_X1 U14171 ( .A(n11722), .ZN(n11723) );
  OAI211_X1 U14172 ( .C1(n11726), .C2(n11731), .A(n13909), .B(n14245), .ZN(
        n11728) );
  INV_X1 U14173 ( .A(n13764), .ZN(n13776) );
  AOI22_X1 U14174 ( .A1(n14133), .A2(n13776), .B1(n13889), .B2(n14135), .ZN(
        n11727) );
  NAND2_X1 U14175 ( .A1(n11728), .A2(n11727), .ZN(n11785) );
  INV_X1 U14176 ( .A(n11785), .ZN(n11740) );
  NAND2_X1 U14177 ( .A1(n13634), .A2(n13776), .ZN(n11729) );
  INV_X1 U14178 ( .A(n11731), .ZN(n11732) );
  OAI21_X1 U14179 ( .B1(n6532), .B2(n11732), .A(n13888), .ZN(n11787) );
  OAI21_X1 U14180 ( .B1(n11906), .B2(n7214), .A(n6422), .ZN(n11784) );
  INV_X1 U14181 ( .A(n11734), .ZN(n13762) );
  OAI22_X1 U14182 ( .A1(n14613), .A2(n11735), .B1(n13762), .B2(n14638), .ZN(
        n11736) );
  AOI21_X1 U14183 ( .B1(n13887), .B2(n14114), .A(n11736), .ZN(n11737) );
  OAI21_X1 U14184 ( .B1(n11784), .B2(n14111), .A(n11737), .ZN(n11738) );
  AOI21_X1 U14185 ( .B1(n11787), .B2(n14621), .A(n11738), .ZN(n11739) );
  OAI21_X1 U14186 ( .B1(n14091), .B2(n11740), .A(n11739), .ZN(P1_U3278) );
  AOI211_X1 U14187 ( .C1(n14845), .C2(n11743), .A(n11742), .B(n11741), .ZN(
        n11750) );
  INV_X1 U14188 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n11744) );
  OAI22_X1 U14189 ( .A1(n11745), .A2(n13584), .B1(n14848), .B2(n11744), .ZN(
        n11746) );
  INV_X1 U14190 ( .A(n11746), .ZN(n11747) );
  OAI21_X1 U14191 ( .B1(n11750), .B2(n14846), .A(n11747), .ZN(P2_U3472) );
  AOI22_X1 U14192 ( .A1(n14511), .A2(n11748), .B1(n14850), .B2(
        P2_REG1_REG_14__SCAN_IN), .ZN(n11749) );
  OAI21_X1 U14193 ( .B1(n11750), .B2(n14850), .A(n11749), .ZN(P2_U3513) );
  INV_X1 U14194 ( .A(n11751), .ZN(n11753) );
  NAND2_X1 U14195 ( .A1(n11753), .A2(n11752), .ZN(n11757) );
  NOR2_X1 U14196 ( .A1(n13854), .A2(n11754), .ZN(n11755) );
  AOI21_X1 U14197 ( .B1(n11754), .B2(n13854), .A(n11755), .ZN(n11756) );
  NAND2_X1 U14198 ( .A1(n11756), .A2(n11757), .ZN(n13853) );
  OAI211_X1 U14199 ( .C1(n11757), .C2(n11756), .A(n13873), .B(n13853), .ZN(
        n11766) );
  INV_X1 U14200 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n11758) );
  NAND2_X1 U14201 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13699)
         );
  OAI21_X1 U14202 ( .B1(n14607), .B2(n11758), .A(n13699), .ZN(n11764) );
  XNOR2_X1 U14203 ( .A(n13846), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n11761) );
  NOR2_X1 U14204 ( .A1(n11762), .A2(n11761), .ZN(n13845) );
  AOI211_X1 U14205 ( .C1(n11762), .C2(n11761), .A(n13845), .B(n13847), .ZN(
        n11763) );
  AOI211_X1 U14206 ( .C1(n13852), .C2(n13846), .A(n11764), .B(n11763), .ZN(
        n11765) );
  NAND2_X1 U14207 ( .A1(n11766), .A2(n11765), .ZN(P1_U3260) );
  INV_X1 U14208 ( .A(n11767), .ZN(n11772) );
  AOI21_X1 U14209 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n13602), .A(n11768), 
        .ZN(n11769) );
  OAI21_X1 U14210 ( .B1(n11772), .B2(n13605), .A(n11769), .ZN(P2_U3304) );
  NAND2_X1 U14211 ( .A1(n14288), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n11771) );
  OAI211_X1 U14212 ( .C1(n11772), .C2(n14300), .A(n11771), .B(n11770), .ZN(
        P1_U3332) );
  XNOR2_X1 U14213 ( .A(n12794), .B(n12111), .ZN(n11812) );
  XNOR2_X1 U14214 ( .A(n11812), .B(n12778), .ZN(n11778) );
  AND2_X1 U14215 ( .A1(n11773), .A2(n14470), .ZN(n11774) );
  INV_X1 U14216 ( .A(n11814), .ZN(n11776) );
  AOI21_X1 U14217 ( .B1(n11778), .B2(n11777), .A(n11776), .ZN(n11783) );
  NAND2_X1 U14218 ( .A1(n12198), .A2(n12795), .ZN(n11780) );
  AND2_X1 U14219 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n12493) );
  AOI21_X1 U14220 ( .B1(n12194), .B2(n12438), .A(n12493), .ZN(n11779) );
  OAI211_X1 U14221 ( .C1(n12790), .C2(n12196), .A(n11780), .B(n11779), .ZN(
        n11781) );
  AOI21_X1 U14222 ( .B1(n12794), .B2(n12185), .A(n11781), .ZN(n11782) );
  OAI21_X1 U14223 ( .B1(n11783), .B2(n12187), .A(n11782), .ZN(P3_U3155) );
  OAI22_X1 U14224 ( .A1(n11784), .A2(n14662), .B1(n11906), .B2(n14670), .ZN(
        n11786) );
  AOI211_X1 U14225 ( .C1(n11787), .C2(n14677), .A(n11786), .B(n11785), .ZN(
        n11790) );
  NAND2_X1 U14226 ( .A1(n14678), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n11788) );
  OAI21_X1 U14227 ( .B1(n11790), .B2(n14678), .A(n11788), .ZN(P1_U3504) );
  NAND2_X1 U14228 ( .A1(n14685), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n11789) );
  OAI21_X1 U14229 ( .B1(n11790), .B2(n14685), .A(n11789), .ZN(P1_U3543) );
  INV_X1 U14230 ( .A(n11793), .ZN(n11794) );
  NAND2_X1 U14231 ( .A1(n11795), .A2(n11794), .ZN(n11796) );
  XNOR2_X1 U14232 ( .A(n14511), .B(n12048), .ZN(n11798) );
  NAND2_X1 U14233 ( .A1(n13101), .A2(n10035), .ZN(n11799) );
  NAND2_X1 U14234 ( .A1(n11798), .A2(n11799), .ZN(n11803) );
  INV_X1 U14235 ( .A(n11798), .ZN(n11801) );
  INV_X1 U14236 ( .A(n11799), .ZN(n11800) );
  NAND2_X1 U14237 ( .A1(n11801), .A2(n11800), .ZN(n11802) );
  NAND2_X1 U14238 ( .A1(n11803), .A2(n11802), .ZN(n14506) );
  XNOR2_X1 U14239 ( .A(n14540), .B(n12048), .ZN(n11999) );
  AND2_X1 U14240 ( .A1(n13100), .A2(n10035), .ZN(n11996) );
  XNOR2_X1 U14241 ( .A(n11997), .B(n11996), .ZN(n11811) );
  NOR2_X1 U14242 ( .A1(n14701), .A2(n11804), .ZN(n11808) );
  OAI22_X1 U14243 ( .A1(n13091), .A2(n11806), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11805), .ZN(n11807) );
  AOI211_X1 U14244 ( .C1(n11809), .C2(n14697), .A(n11808), .B(n11807), .ZN(
        n11810) );
  OAI21_X1 U14245 ( .B1(n11811), .B2(n13073), .A(n11810), .ZN(P2_U3213) );
  INV_X1 U14246 ( .A(n12337), .ZN(n12951) );
  NAND2_X1 U14247 ( .A1(n11812), .A2(n12778), .ZN(n11813) );
  XNOR2_X1 U14248 ( .A(n12337), .B(n12111), .ZN(n12060) );
  XNOR2_X1 U14249 ( .A(n12060), .B(n12437), .ZN(n11815) );
  OAI211_X1 U14250 ( .C1(n11816), .C2(n11815), .A(n12062), .B(n12192), .ZN(
        n11820) );
  NOR2_X1 U14251 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15243), .ZN(n12513) );
  AOI21_X1 U14252 ( .B1(n12194), .B2(n12802), .A(n12513), .ZN(n11817) );
  OAI21_X1 U14253 ( .B1(n12779), .B2(n12196), .A(n11817), .ZN(n11818) );
  AOI21_X1 U14254 ( .B1(n12198), .B2(n12782), .A(n11818), .ZN(n11819) );
  OAI211_X1 U14255 ( .C1(n12951), .C2(n12201), .A(n11820), .B(n11819), .ZN(
        P3_U3181) );
  NAND2_X1 U14256 ( .A1(n14540), .A2(n13100), .ZN(n11821) );
  OR2_X1 U14257 ( .A1(n13585), .A2(n13099), .ZN(n11823) );
  XNOR2_X1 U14258 ( .A(n13185), .B(n13226), .ZN(n13528) );
  NAND2_X1 U14259 ( .A1(n14540), .A2(n11826), .ZN(n11827) );
  OR2_X1 U14260 ( .A1(n13585), .A2(n11830), .ZN(n11828) );
  XNOR2_X1 U14261 ( .A(n13227), .B(n7287), .ZN(n13523) );
  AND2_X1 U14262 ( .A1(n13424), .A2(n13229), .ZN(n11829) );
  OR3_X1 U14263 ( .A1(n13410), .A2(n11829), .A3(n10035), .ZN(n13525) );
  OAI22_X1 U14264 ( .A1(n13231), .A2(n13067), .B1(n11830), .B2(n13059), .ZN(
        n13036) );
  INV_X1 U14265 ( .A(n13036), .ZN(n13524) );
  OAI22_X1 U14266 ( .A1(n14819), .A2(n13524), .B1(n13034), .B2(n13407), .ZN(
        n11832) );
  NOR2_X1 U14267 ( .A1(n13580), .A2(n14812), .ZN(n11831) );
  AOI211_X1 U14268 ( .C1(n14819), .C2(P2_REG2_REG_17__SCAN_IN), .A(n11832), 
        .B(n11831), .ZN(n11833) );
  OAI21_X1 U14269 ( .B1(n13525), .B2(n13413), .A(n11833), .ZN(n11834) );
  AOI21_X1 U14270 ( .B1(n13523), .B2(n14815), .A(n11834), .ZN(n11835) );
  OAI21_X1 U14271 ( .B1(n13440), .B2(n13528), .A(n11835), .ZN(P2_U3248) );
  MUX2_X1 U14272 ( .A(n11836), .B(P1_REG2_REG_3__SCAN_IN), .S(n14091), .Z(
        n11844) );
  NAND2_X1 U14273 ( .A1(n11838), .A2(n11837), .ZN(n11842) );
  INV_X1 U14274 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n11839) );
  AOI22_X1 U14275 ( .A1(n14146), .A2(n11840), .B1(n14089), .B2(n11839), .ZN(
        n11841) );
  OAI211_X1 U14276 ( .C1(n6936), .C2(n14125), .A(n11842), .B(n11841), .ZN(
        n11843) );
  OR2_X1 U14277 ( .A1(n11844), .A2(n11843), .ZN(P1_U3290) );
  INV_X1 U14278 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n11850) );
  OAI222_X1 U14279 ( .A1(n13605), .A2(n14283), .B1(n11845), .B2(P2_U3088), 
        .C1(n11850), .C2(n13614), .ZN(P2_U3297) );
  INV_X1 U14280 ( .A(SI_30_), .ZN(n15123) );
  INV_X1 U14281 ( .A(n11846), .ZN(n11848) );
  INV_X1 U14282 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14282) );
  NAND2_X1 U14283 ( .A1(n14282), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12207) );
  NAND2_X1 U14284 ( .A1(n11850), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n11851) );
  AND2_X1 U14285 ( .A1(n12207), .A2(n11851), .ZN(n11852) );
  NAND2_X1 U14286 ( .A1(n11853), .A2(n11852), .ZN(n12208) );
  OR2_X1 U14287 ( .A1(n11853), .A2(n11852), .ZN(n11854) );
  INV_X1 U14288 ( .A(n12203), .ZN(n11855) );
  OAI222_X1 U14289 ( .A1(P3_U3151), .A2(n11856), .B1(n12973), .B2(n15123), 
        .C1(n14410), .C2(n11855), .ZN(P3_U3265) );
  INV_X1 U14290 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n11859) );
  AND2_X2 U14291 ( .A1(n13410), .A2(n13520), .ZN(n13411) );
  NAND2_X1 U14292 ( .A1(n13221), .A2(n13545), .ZN(n13179) );
  NOR2_X1 U14293 ( .A1(n13600), .A2(n11857), .ZN(n11858) );
  NOR2_X1 U14294 ( .A1(n13067), .A2(n11858), .ZN(n13216) );
  AND2_X1 U14295 ( .A1(n13097), .A2(n13216), .ZN(n11865) );
  INV_X1 U14296 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n11861) );
  MUX2_X1 U14297 ( .A(n11861), .B(n11860), .S(n14852), .Z(n11862) );
  OAI21_X1 U14298 ( .B1(n11868), .B2(n13541), .A(n11862), .ZN(P2_U3530) );
  NAND2_X1 U14299 ( .A1(n11864), .A2(n11863), .ZN(n11867) );
  INV_X1 U14300 ( .A(n11865), .ZN(n13441) );
  NOR2_X1 U14301 ( .A1(n6388), .A2(n13441), .ZN(n13181) );
  AOI21_X1 U14302 ( .B1(n6388), .B2(P2_REG2_REG_31__SCAN_IN), .A(n13181), .ZN(
        n11866) );
  OAI211_X1 U14303 ( .C1(n11868), .C2(n14812), .A(n11867), .B(n11866), .ZN(
        P2_U3234) );
  INV_X1 U14304 ( .A(n13595), .ZN(n11870) );
  OAI222_X1 U14305 ( .A1(n13796), .A2(P1_U3086), .B1(n14300), .B2(n11870), 
        .C1(n11869), .C2(n14298), .ZN(P1_U3327) );
  NOR2_X1 U14306 ( .A1(n14103), .A2(n10259), .ZN(n11871) );
  AOI21_X1 U14307 ( .B1(n14086), .B2(n11981), .A(n11871), .ZN(n11931) );
  INV_X1 U14308 ( .A(n11931), .ZN(n11934) );
  NAND2_X1 U14309 ( .A1(n14086), .A2(n11982), .ZN(n11873) );
  INV_X1 U14310 ( .A(n14103), .ZN(n13896) );
  NAND2_X1 U14311 ( .A1(n13896), .A2(n11981), .ZN(n11872) );
  NAND2_X1 U14312 ( .A1(n11873), .A2(n11872), .ZN(n11874) );
  XNOR2_X1 U14313 ( .A(n11874), .B(n11948), .ZN(n11932) );
  INV_X1 U14314 ( .A(n11932), .ZN(n11933) );
  NAND2_X1 U14315 ( .A1(n11876), .A2(n11875), .ZN(n11877) );
  NAND2_X1 U14316 ( .A1(n13661), .A2(n11982), .ZN(n11880) );
  OR2_X1 U14317 ( .A1(n10140), .A2(n11882), .ZN(n11879) );
  NAND2_X1 U14318 ( .A1(n11880), .A2(n11879), .ZN(n11881) );
  XNOR2_X1 U14319 ( .A(n11881), .B(n11983), .ZN(n11884) );
  NOR2_X1 U14320 ( .A1(n10259), .A2(n11882), .ZN(n11883) );
  AOI21_X1 U14321 ( .B1(n13661), .B2(n11981), .A(n11883), .ZN(n11885) );
  XNOR2_X1 U14322 ( .A(n11884), .B(n11885), .ZN(n13663) );
  INV_X1 U14323 ( .A(n11884), .ZN(n11886) );
  OR2_X1 U14324 ( .A1(n11886), .A2(n11885), .ZN(n11887) );
  NAND2_X1 U14325 ( .A1(n14562), .A2(n11982), .ZN(n11889) );
  OR2_X1 U14326 ( .A1(n10140), .A2(n13666), .ZN(n11888) );
  NAND2_X1 U14327 ( .A1(n11889), .A2(n11888), .ZN(n11890) );
  XNOR2_X1 U14328 ( .A(n11890), .B(n11983), .ZN(n11892) );
  NOR2_X1 U14329 ( .A1(n10259), .A2(n13666), .ZN(n11891) );
  AOI21_X1 U14330 ( .B1(n14562), .B2(n11981), .A(n11891), .ZN(n11893) );
  XNOR2_X1 U14331 ( .A(n11892), .B(n11893), .ZN(n13723) );
  INV_X1 U14332 ( .A(n11892), .ZN(n11894) );
  OR2_X1 U14333 ( .A1(n11894), .A2(n11893), .ZN(n11895) );
  NAND2_X1 U14334 ( .A1(n11896), .A2(n11895), .ZN(n13627) );
  NAND2_X1 U14335 ( .A1(n13634), .A2(n11982), .ZN(n11898) );
  OR2_X1 U14336 ( .A1(n13764), .A2(n10140), .ZN(n11897) );
  NAND2_X1 U14337 ( .A1(n11898), .A2(n11897), .ZN(n11899) );
  XNOR2_X1 U14338 ( .A(n11899), .B(n11948), .ZN(n11902) );
  NOR2_X1 U14339 ( .A1(n10259), .A2(n13764), .ZN(n11900) );
  AOI21_X1 U14340 ( .B1(n13634), .B2(n11981), .A(n11900), .ZN(n11901) );
  NAND2_X1 U14341 ( .A1(n11902), .A2(n11901), .ZN(n11904) );
  OR2_X1 U14342 ( .A1(n11902), .A2(n11901), .ZN(n11903) );
  NAND2_X1 U14343 ( .A1(n11904), .A2(n11903), .ZN(n13628) );
  OAI22_X1 U14344 ( .A1(n11906), .A2(n11935), .B1(n13686), .B2(n10140), .ZN(
        n11905) );
  XNOR2_X1 U14345 ( .A(n11905), .B(n11983), .ZN(n11907) );
  OAI22_X1 U14346 ( .A1(n11906), .A2(n10140), .B1(n13686), .B2(n10259), .ZN(
        n13761) );
  NAND2_X1 U14347 ( .A1(n14132), .A2(n6391), .ZN(n11909) );
  NAND2_X1 U14348 ( .A1(n13889), .A2(n11981), .ZN(n11908) );
  NAND2_X1 U14349 ( .A1(n11909), .A2(n11908), .ZN(n11910) );
  XNOR2_X1 U14350 ( .A(n11910), .B(n11983), .ZN(n11914) );
  NAND2_X1 U14351 ( .A1(n14132), .A2(n11981), .ZN(n11912) );
  NAND2_X1 U14352 ( .A1(n11985), .A2(n13889), .ZN(n11911) );
  NAND2_X1 U14353 ( .A1(n11912), .A2(n11911), .ZN(n11913) );
  NOR2_X1 U14354 ( .A1(n11914), .A2(n11913), .ZN(n11915) );
  AOI21_X1 U14355 ( .B1(n11914), .B2(n11913), .A(n11915), .ZN(n13684) );
  INV_X1 U14356 ( .A(n11915), .ZN(n13693) );
  OAI22_X1 U14357 ( .A1(n14242), .A2(n11935), .B1(n13892), .B2(n10140), .ZN(
        n11916) );
  XNOR2_X1 U14358 ( .A(n11916), .B(n11948), .ZN(n11919) );
  OR2_X1 U14359 ( .A1(n14242), .A2(n10140), .ZN(n11918) );
  NAND2_X1 U14360 ( .A1(n11985), .A2(n14136), .ZN(n11917) );
  AND2_X1 U14361 ( .A1(n11918), .A2(n11917), .ZN(n11920) );
  NAND2_X1 U14362 ( .A1(n11919), .A2(n11920), .ZN(n11924) );
  INV_X1 U14363 ( .A(n11919), .ZN(n11922) );
  INV_X1 U14364 ( .A(n11920), .ZN(n11921) );
  NAND2_X1 U14365 ( .A1(n11922), .A2(n11921), .ZN(n11923) );
  NAND2_X1 U14366 ( .A1(n11924), .A2(n11923), .ZN(n13692) );
  INV_X1 U14367 ( .A(n11924), .ZN(n11925) );
  OAI22_X1 U14368 ( .A1(n14110), .A2(n11935), .B1(n14079), .B2(n10140), .ZN(
        n11926) );
  XNOR2_X1 U14369 ( .A(n11926), .B(n11983), .ZN(n11930) );
  OR2_X1 U14370 ( .A1(n14110), .A2(n10140), .ZN(n11928) );
  NAND2_X1 U14371 ( .A1(n13913), .A2(n11985), .ZN(n11927) );
  NAND2_X1 U14372 ( .A1(n11928), .A2(n11927), .ZN(n11929) );
  XNOR2_X1 U14373 ( .A(n11930), .B(n11929), .ZN(n13742) );
  NOR2_X1 U14374 ( .A1(n11930), .A2(n11929), .ZN(n13648) );
  XNOR2_X1 U14375 ( .A(n11932), .B(n11931), .ZN(n13647) );
  OAI22_X1 U14376 ( .A1(n14218), .A2(n11935), .B1(n14080), .B2(n10140), .ZN(
        n11936) );
  XNOR2_X1 U14377 ( .A(n11936), .B(n11983), .ZN(n11938) );
  OAI22_X1 U14378 ( .A1(n14218), .A2(n10140), .B1(n14080), .B2(n10259), .ZN(
        n11937) );
  XNOR2_X1 U14379 ( .A(n11938), .B(n11937), .ZN(n13715) );
  NAND2_X1 U14380 ( .A1(n14212), .A2(n6391), .ZN(n11940) );
  NAND2_X1 U14381 ( .A1(n14062), .A2(n11981), .ZN(n11939) );
  NAND2_X1 U14382 ( .A1(n11940), .A2(n11939), .ZN(n11941) );
  XNOR2_X1 U14383 ( .A(n11941), .B(n11948), .ZN(n11944) );
  AND2_X1 U14384 ( .A1(n14062), .A2(n11985), .ZN(n11942) );
  AOI21_X1 U14385 ( .B1(n14212), .B2(n11981), .A(n11942), .ZN(n11943) );
  NAND2_X1 U14386 ( .A1(n11944), .A2(n11943), .ZN(n11945) );
  OAI21_X1 U14387 ( .B1(n11944), .B2(n11943), .A(n11945), .ZN(n13654) );
  INV_X1 U14388 ( .A(n11945), .ZN(n13733) );
  NAND2_X1 U14389 ( .A1(n14206), .A2(n11982), .ZN(n11947) );
  NAND2_X1 U14390 ( .A1(n13775), .A2(n11981), .ZN(n11946) );
  NAND2_X1 U14391 ( .A1(n11947), .A2(n11946), .ZN(n11949) );
  XNOR2_X1 U14392 ( .A(n11949), .B(n11948), .ZN(n11951) );
  AND2_X1 U14393 ( .A1(n13775), .A2(n11985), .ZN(n11950) );
  AOI21_X1 U14394 ( .B1(n14206), .B2(n11981), .A(n11950), .ZN(n11952) );
  NAND2_X1 U14395 ( .A1(n11951), .A2(n11952), .ZN(n11956) );
  INV_X1 U14396 ( .A(n11951), .ZN(n11954) );
  INV_X1 U14397 ( .A(n11952), .ZN(n11953) );
  NAND2_X1 U14398 ( .A1(n11954), .A2(n11953), .ZN(n11955) );
  AND2_X1 U14399 ( .A1(n11956), .A2(n11955), .ZN(n13732) );
  AOI22_X1 U14400 ( .A1(n14017), .A2(n6391), .B1(n11981), .B2(n14037), .ZN(
        n11957) );
  XOR2_X1 U14401 ( .A(n11983), .B(n11957), .Z(n11959) );
  INV_X1 U14402 ( .A(n14037), .ZN(n13919) );
  OAI22_X1 U14403 ( .A1(n14197), .A2(n10140), .B1(n13919), .B2(n10259), .ZN(
        n11958) );
  NOR2_X1 U14404 ( .A1(n11959), .A2(n11958), .ZN(n11960) );
  AOI21_X1 U14405 ( .B1(n11959), .B2(n11958), .A(n11960), .ZN(n13639) );
  NAND2_X1 U14406 ( .A1(n13638), .A2(n13639), .ZN(n13637) );
  INV_X1 U14407 ( .A(n11960), .ZN(n11961) );
  AOI22_X1 U14408 ( .A1(n14193), .A2(n11982), .B1(n11981), .B2(n13774), .ZN(
        n11962) );
  XOR2_X1 U14409 ( .A(n11983), .B(n11962), .Z(n11964) );
  INV_X1 U14410 ( .A(n13774), .ZN(n13921) );
  OAI22_X1 U14411 ( .A1(n14012), .A2(n10140), .B1(n13921), .B2(n10259), .ZN(
        n11963) );
  NOR2_X1 U14412 ( .A1(n11964), .A2(n11963), .ZN(n11965) );
  AOI21_X1 U14413 ( .B1(n11964), .B2(n11963), .A(n11965), .ZN(n13705) );
  INV_X1 U14414 ( .A(n11965), .ZN(n11966) );
  NAND2_X1 U14415 ( .A1(n13703), .A2(n11966), .ZN(n13674) );
  AOI22_X1 U14416 ( .A1(n13922), .A2(n11982), .B1(n11981), .B2(n13773), .ZN(
        n11967) );
  XOR2_X1 U14417 ( .A(n11983), .B(n11967), .Z(n11969) );
  OAI22_X1 U14418 ( .A1(n14183), .A2(n10140), .B1(n13923), .B2(n10259), .ZN(
        n11968) );
  NOR2_X1 U14419 ( .A1(n11969), .A2(n11968), .ZN(n11970) );
  AOI21_X1 U14420 ( .B1(n11969), .B2(n11968), .A(n11970), .ZN(n13675) );
  INV_X1 U14421 ( .A(n11970), .ZN(n11971) );
  NAND2_X1 U14422 ( .A1(n13673), .A2(n11971), .ZN(n13749) );
  AOI22_X1 U14423 ( .A1(n14179), .A2(n6391), .B1(n11981), .B2(n13962), .ZN(
        n11972) );
  XOR2_X1 U14424 ( .A(n11983), .B(n11972), .Z(n11974) );
  INV_X1 U14425 ( .A(n13962), .ZN(n13903) );
  OAI22_X1 U14426 ( .A1(n13982), .A2(n10140), .B1(n13903), .B2(n10259), .ZN(
        n11973) );
  NOR2_X1 U14427 ( .A1(n11974), .A2(n11973), .ZN(n11975) );
  AOI21_X1 U14428 ( .B1(n11974), .B2(n11973), .A(n11975), .ZN(n13750) );
  INV_X1 U14429 ( .A(n11975), .ZN(n11976) );
  AOI22_X1 U14430 ( .A1(n14171), .A2(n6391), .B1(n11981), .B2(n13942), .ZN(
        n11977) );
  XOR2_X1 U14431 ( .A(n11983), .B(n11977), .Z(n11979) );
  INV_X1 U14432 ( .A(n13942), .ZN(n13924) );
  OAI22_X1 U14433 ( .A1(n13968), .A2(n10140), .B1(n13924), .B2(n10259), .ZN(
        n11978) );
  NOR2_X1 U14434 ( .A1(n11979), .A2(n11978), .ZN(n11980) );
  AOI21_X1 U14435 ( .B1(n11979), .B2(n11978), .A(n11980), .ZN(n13619) );
  AOI22_X1 U14436 ( .A1(n14167), .A2(n11982), .B1(n11981), .B2(n13961), .ZN(
        n11984) );
  XNOR2_X1 U14437 ( .A(n11984), .B(n11983), .ZN(n11987) );
  AOI22_X1 U14438 ( .A1(n14167), .A2(n11981), .B1(n11985), .B2(n13961), .ZN(
        n11986) );
  XNOR2_X1 U14439 ( .A(n11989), .B(n11988), .ZN(n11995) );
  OAI22_X1 U14440 ( .A1(n13763), .A2(n13950), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11990), .ZN(n11993) );
  OAI22_X1 U14441 ( .A1(n13924), .A2(n13765), .B1(n13766), .B2(n11991), .ZN(
        n11992) );
  AOI211_X1 U14442 ( .C1(n14167), .C2(n13769), .A(n11993), .B(n11992), .ZN(
        n11994) );
  OAI21_X1 U14443 ( .B1(n11995), .B2(n13771), .A(n11994), .ZN(P1_U3220) );
  NOR2_X1 U14444 ( .A1(n13253), .A2(n13390), .ZN(n12047) );
  XNOR2_X1 U14445 ( .A(n13292), .B(n12995), .ZN(n12046) );
  NOR2_X1 U14446 ( .A1(n13206), .A2(n13390), .ZN(n12041) );
  XNOR2_X1 U14447 ( .A(n13559), .B(n12995), .ZN(n12040) );
  INV_X1 U14448 ( .A(n11998), .ZN(n12000) );
  NAND2_X1 U14449 ( .A1(n12000), .A2(n11999), .ZN(n12001) );
  XNOR2_X1 U14450 ( .A(n13585), .B(n12995), .ZN(n12002) );
  NAND2_X1 U14451 ( .A1(n13099), .A2(n10035), .ZN(n12003) );
  NAND2_X1 U14452 ( .A1(n12002), .A2(n12003), .ZN(n12007) );
  INV_X1 U14453 ( .A(n12002), .ZN(n12005) );
  INV_X1 U14454 ( .A(n12003), .ZN(n12004) );
  NAND2_X1 U14455 ( .A1(n12005), .A2(n12004), .ZN(n12006) );
  NAND2_X1 U14456 ( .A1(n12007), .A2(n12006), .ZN(n13024) );
  XNOR2_X1 U14457 ( .A(n13229), .B(n12048), .ZN(n12008) );
  NAND2_X1 U14458 ( .A1(n13228), .A2(n10035), .ZN(n12009) );
  NAND2_X1 U14459 ( .A1(n12008), .A2(n12009), .ZN(n12013) );
  INV_X1 U14460 ( .A(n12008), .ZN(n12011) );
  INV_X1 U14461 ( .A(n12009), .ZN(n12010) );
  NAND2_X1 U14462 ( .A1(n12011), .A2(n12010), .ZN(n12012) );
  AND2_X1 U14463 ( .A1(n12013), .A2(n12012), .ZN(n13032) );
  XNOR2_X1 U14464 ( .A(n13520), .B(n12995), .ZN(n12014) );
  NAND2_X1 U14465 ( .A1(n13190), .A2(n10035), .ZN(n12015) );
  XNOR2_X1 U14466 ( .A(n12014), .B(n12015), .ZN(n13065) );
  INV_X1 U14467 ( .A(n13065), .ZN(n12018) );
  INV_X1 U14468 ( .A(n12014), .ZN(n12017) );
  INV_X1 U14469 ( .A(n12015), .ZN(n12016) );
  XNOR2_X1 U14470 ( .A(n13575), .B(n12995), .ZN(n12019) );
  OR2_X1 U14471 ( .A1(n13233), .A2(n13390), .ZN(n12020) );
  NAND2_X1 U14472 ( .A1(n12019), .A2(n12020), .ZN(n12024) );
  INV_X1 U14473 ( .A(n12019), .ZN(n12022) );
  INV_X1 U14474 ( .A(n12020), .ZN(n12021) );
  NAND2_X1 U14475 ( .A1(n12022), .A2(n12021), .ZN(n12023) );
  AND2_X1 U14476 ( .A1(n12024), .A2(n12023), .ZN(n12985) );
  XNOR2_X1 U14477 ( .A(n13370), .B(n12048), .ZN(n12025) );
  NAND2_X1 U14478 ( .A1(n13237), .A2(n10035), .ZN(n12026) );
  NAND2_X1 U14479 ( .A1(n12025), .A2(n12026), .ZN(n13049) );
  INV_X1 U14480 ( .A(n12025), .ZN(n12028) );
  INV_X1 U14481 ( .A(n12026), .ZN(n12027) );
  NAND2_X1 U14482 ( .A1(n12028), .A2(n12027), .ZN(n13050) );
  NAND2_X1 U14483 ( .A1(n12029), .A2(n13050), .ZN(n13006) );
  XNOR2_X1 U14484 ( .A(n13567), .B(n12995), .ZN(n12030) );
  NOR2_X1 U14485 ( .A1(n13239), .A2(n13390), .ZN(n12031) );
  XNOR2_X1 U14486 ( .A(n12030), .B(n12031), .ZN(n13005) );
  NAND2_X1 U14487 ( .A1(n13006), .A2(n13005), .ZN(n13004) );
  INV_X1 U14488 ( .A(n12030), .ZN(n12032) );
  NAND2_X1 U14489 ( .A1(n12032), .A2(n12031), .ZN(n12033) );
  XNOR2_X1 U14490 ( .A(n13491), .B(n12995), .ZN(n12034) );
  NOR2_X1 U14491 ( .A1(n13243), .A2(n13390), .ZN(n13058) );
  INV_X1 U14492 ( .A(n12037), .ZN(n12039) );
  XNOR2_X1 U14493 ( .A(n13336), .B(n12995), .ZN(n12038) );
  NAND2_X1 U14494 ( .A1(n13245), .A2(n10035), .ZN(n12978) );
  XNOR2_X1 U14495 ( .A(n12040), .B(n12041), .ZN(n13040) );
  XNOR2_X1 U14496 ( .A(n13555), .B(n12048), .ZN(n12043) );
  NOR2_X1 U14497 ( .A1(n13250), .A2(n13390), .ZN(n12042) );
  NAND2_X1 U14498 ( .A1(n12043), .A2(n12042), .ZN(n12044) );
  OAI21_X1 U14499 ( .B1(n12043), .B2(n12042), .A(n12044), .ZN(n13017) );
  INV_X1 U14500 ( .A(n12044), .ZN(n12045) );
  XOR2_X1 U14501 ( .A(n12047), .B(n12046), .Z(n13085) );
  XNOR2_X1 U14502 ( .A(n13550), .B(n12048), .ZN(n12050) );
  NOR2_X1 U14503 ( .A1(n13000), .A2(n13390), .ZN(n12049) );
  NAND2_X1 U14504 ( .A1(n12050), .A2(n12049), .ZN(n12992) );
  OAI21_X1 U14505 ( .B1(n12050), .B2(n12049), .A(n12992), .ZN(n12051) );
  AOI22_X1 U14506 ( .A1(n13217), .A2(n14524), .B1(n14522), .B2(n13252), .ZN(
        n13277) );
  OAI22_X1 U14507 ( .A1(n13091), .A2(n13277), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12055), .ZN(n12056) );
  AOI21_X1 U14508 ( .B1(n13282), .B2(n13093), .A(n12056), .ZN(n12057) );
  OAI211_X1 U14509 ( .C1(n13550), .C2(n13096), .A(n12058), .B(n12057), .ZN(
        P2_U3186) );
  XNOR2_X1 U14510 ( .A(n12089), .B(n12634), .ZN(n12059) );
  INV_X1 U14511 ( .A(n12641), .ZN(n12431) );
  NOR2_X1 U14512 ( .A1(n12059), .A2(n12431), .ZN(n12110) );
  XNOR2_X1 U14513 ( .A(n12348), .B(n10229), .ZN(n12147) );
  INV_X1 U14514 ( .A(n12060), .ZN(n12061) );
  XNOR2_X1 U14515 ( .A(n12769), .B(n10229), .ZN(n12063) );
  XNOR2_X1 U14516 ( .A(n12063), .B(n12751), .ZN(n12140) );
  INV_X1 U14517 ( .A(n12063), .ZN(n12064) );
  AND2_X1 U14518 ( .A1(n12064), .A2(n12751), .ZN(n12065) );
  NOR2_X1 U14519 ( .A1(n12147), .A2(n12765), .ZN(n12153) );
  XNOR2_X1 U14520 ( .A(n12880), .B(n12111), .ZN(n12066) );
  XNOR2_X1 U14521 ( .A(n12066), .B(n12726), .ZN(n12178) );
  XNOR2_X1 U14522 ( .A(n12935), .B(n10229), .ZN(n12067) );
  XNOR2_X1 U14523 ( .A(n12067), .B(n12742), .ZN(n12103) );
  XNOR2_X1 U14524 ( .A(n12871), .B(n12111), .ZN(n12068) );
  XNOR2_X1 U14525 ( .A(n12068), .B(n12727), .ZN(n12165) );
  XNOR2_X1 U14526 ( .A(n12705), .B(n10229), .ZN(n12069) );
  NAND2_X1 U14527 ( .A1(n12069), .A2(n12690), .ZN(n12070) );
  OAI21_X1 U14528 ( .B1(n12069), .B2(n12690), .A(n12070), .ZN(n12123) );
  INV_X1 U14529 ( .A(n12070), .ZN(n12071) );
  INV_X1 U14530 ( .A(n12073), .ZN(n12075) );
  XOR2_X1 U14531 ( .A(n12111), .B(n12694), .Z(n12072) );
  INV_X1 U14532 ( .A(n12072), .ZN(n12074) );
  INV_X1 U14533 ( .A(n12078), .ZN(n12076) );
  XNOR2_X1 U14534 ( .A(n12667), .B(n12111), .ZN(n12081) );
  NAND2_X1 U14535 ( .A1(n12081), .A2(n12676), .ZN(n12084) );
  INV_X1 U14536 ( .A(n12081), .ZN(n12082) );
  NAND2_X1 U14537 ( .A1(n12082), .A2(n12135), .ZN(n12083) );
  NAND2_X1 U14538 ( .A1(n12084), .A2(n12083), .ZN(n12159) );
  INV_X1 U14539 ( .A(n12084), .ZN(n12132) );
  XNOR2_X1 U14540 ( .A(n12247), .B(n10229), .ZN(n12085) );
  NAND2_X1 U14541 ( .A1(n12085), .A2(n12662), .ZN(n12088) );
  INV_X1 U14542 ( .A(n12085), .ZN(n12086) );
  NAND2_X1 U14543 ( .A1(n12086), .A2(n12433), .ZN(n12087) );
  XNOR2_X1 U14544 ( .A(n12089), .B(n12388), .ZN(n12090) );
  NOR2_X1 U14545 ( .A1(n12090), .A2(n12432), .ZN(n12091) );
  AOI21_X1 U14546 ( .B1(n12090), .B2(n12432), .A(n12091), .ZN(n12191) );
  OAI22_X1 U14547 ( .A1(n12652), .A2(n12114), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12093), .ZN(n12095) );
  NOR2_X1 U14548 ( .A1(n12629), .A2(n12196), .ZN(n12094) );
  AOI211_X1 U14549 ( .C1(n12630), .C2(n12198), .A(n12095), .B(n12094), .ZN(
        n12096) );
  OAI21_X1 U14550 ( .B1(n12691), .B2(n6516), .A(n12097), .ZN(n12098) );
  NAND2_X1 U14551 ( .A1(n12098), .A2(n12192), .ZN(n12102) );
  AOI22_X1 U14552 ( .A1(n12435), .A2(n12194), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12099) );
  OAI21_X1 U14553 ( .B1(n12676), .B2(n12196), .A(n12099), .ZN(n12100) );
  AOI21_X1 U14554 ( .B1(n12680), .B2(n12198), .A(n12100), .ZN(n12101) );
  OAI211_X1 U14555 ( .C1(n12859), .C2(n12201), .A(n12102), .B(n12101), .ZN(
        P3_U3156) );
  XNOR2_X1 U14556 ( .A(n12104), .B(n12103), .ZN(n12109) );
  NAND2_X1 U14557 ( .A1(n12194), .A2(n12752), .ZN(n12105) );
  NAND2_X1 U14558 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12593)
         );
  OAI211_X1 U14559 ( .C1(n12196), .C2(n12727), .A(n12105), .B(n12593), .ZN(
        n12107) );
  NOR2_X1 U14560 ( .A1(n12935), .A2(n12201), .ZN(n12106) );
  AOI211_X1 U14561 ( .C1(n12730), .C2(n12198), .A(n12107), .B(n12106), .ZN(
        n12108) );
  OAI21_X1 U14562 ( .B1(n12109), .B2(n12187), .A(n12108), .ZN(P3_U3159) );
  XNOR2_X1 U14563 ( .A(n12391), .B(n12111), .ZN(n12112) );
  INV_X1 U14564 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n12113) );
  OAI22_X1 U14565 ( .A1(n12641), .A2(n12114), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12113), .ZN(n12118) );
  INV_X1 U14566 ( .A(n12115), .ZN(n12618) );
  OAI22_X1 U14567 ( .A1(n12116), .A2(n12196), .B1(n12618), .B2(n12181), .ZN(
        n12117) );
  AOI211_X1 U14568 ( .C1(n12620), .C2(n12185), .A(n12118), .B(n12117), .ZN(
        n12119) );
  OAI21_X1 U14569 ( .B1(n12120), .B2(n12187), .A(n12119), .ZN(P3_U3160) );
  AOI21_X1 U14570 ( .B1(n12123), .B2(n12122), .A(n12121), .ZN(n12128) );
  NAND2_X1 U14571 ( .A1(n12198), .A2(n12706), .ZN(n12125) );
  AOI22_X1 U14572 ( .A1(n12194), .A2(n12436), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12124) );
  OAI211_X1 U14573 ( .C1(n12702), .C2(n12196), .A(n12125), .B(n12124), .ZN(
        n12126) );
  AOI21_X1 U14574 ( .B1(n12705), .B2(n12185), .A(n12126), .ZN(n12127) );
  OAI21_X1 U14575 ( .B1(n12128), .B2(n12187), .A(n12127), .ZN(P3_U3163) );
  INV_X1 U14576 ( .A(n12129), .ZN(n12134) );
  NOR3_X1 U14577 ( .A1(n12130), .A2(n12132), .A3(n12131), .ZN(n12133) );
  OAI21_X1 U14578 ( .B1(n12134), .B2(n12133), .A(n12192), .ZN(n12139) );
  AOI22_X1 U14579 ( .A1(n12135), .A2(n12194), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12136) );
  OAI21_X1 U14580 ( .B1(n12652), .B2(n12196), .A(n12136), .ZN(n12137) );
  AOI21_X1 U14581 ( .B1(n12653), .B2(n12198), .A(n12137), .ZN(n12138) );
  OAI211_X1 U14582 ( .C1(n12917), .C2(n12201), .A(n12139), .B(n12138), .ZN(
        P3_U3165) );
  XNOR2_X1 U14583 ( .A(n12141), .B(n12140), .ZN(n12146) );
  NAND2_X1 U14584 ( .A1(n12198), .A2(n12770), .ZN(n12143) );
  AND2_X1 U14585 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12539) );
  AOI21_X1 U14586 ( .B1(n12194), .B2(n12437), .A(n12539), .ZN(n12142) );
  OAI211_X1 U14587 ( .C1(n12765), .C2(n12196), .A(n12143), .B(n12142), .ZN(
        n12144) );
  AOI21_X1 U14588 ( .B1(n12769), .B2(n12185), .A(n12144), .ZN(n12145) );
  OAI21_X1 U14589 ( .B1(n12146), .B2(n12187), .A(n12145), .ZN(P3_U3166) );
  INV_X1 U14590 ( .A(n12150), .ZN(n12152) );
  XNOR2_X1 U14591 ( .A(n12147), .B(n12765), .ZN(n12149) );
  AOI21_X1 U14592 ( .B1(n12150), .B2(n12149), .A(n12148), .ZN(n12151) );
  AOI21_X1 U14593 ( .B1(n12153), .B2(n12152), .A(n12151), .ZN(n12158) );
  NAND2_X1 U14594 ( .A1(n12198), .A2(n12758), .ZN(n12155) );
  AOI22_X1 U14595 ( .A1(n12194), .A2(n12751), .B1(P3_REG3_REG_17__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12154) );
  OAI211_X1 U14596 ( .C1(n12726), .C2(n12196), .A(n12155), .B(n12154), .ZN(
        n12156) );
  AOI21_X1 U14597 ( .B1(n12348), .B2(n12185), .A(n12156), .ZN(n12157) );
  OAI21_X1 U14598 ( .B1(n12158), .B2(n12187), .A(n12157), .ZN(P3_U3168) );
  INV_X1 U14599 ( .A(n12667), .ZN(n12921) );
  AND3_X1 U14600 ( .A1(n12097), .A2(n12080), .A3(n12159), .ZN(n12160) );
  OAI21_X1 U14601 ( .B1(n12130), .B2(n12160), .A(n12192), .ZN(n12164) );
  INV_X1 U14602 ( .A(n12691), .ZN(n12434) );
  AOI22_X1 U14603 ( .A1(n12434), .A2(n12194), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12161) );
  OAI21_X1 U14604 ( .B1(n12662), .B2(n12196), .A(n12161), .ZN(n12162) );
  AOI21_X1 U14605 ( .B1(n12663), .B2(n12198), .A(n12162), .ZN(n12163) );
  OAI211_X1 U14606 ( .C1(n12921), .C2(n12201), .A(n12164), .B(n12163), .ZN(
        P3_U3169) );
  XNOR2_X1 U14607 ( .A(n12166), .B(n12165), .ZN(n12171) );
  NAND2_X1 U14608 ( .A1(n12198), .A2(n12716), .ZN(n12168) );
  AOI22_X1 U14609 ( .A1(n12194), .A2(n12713), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12167) );
  OAI211_X1 U14610 ( .C1(n12690), .C2(n12196), .A(n12168), .B(n12167), .ZN(
        n12169) );
  AOI21_X1 U14611 ( .B1(n12871), .B2(n12185), .A(n12169), .ZN(n12170) );
  OAI21_X1 U14612 ( .B1(n12171), .B2(n12187), .A(n12170), .ZN(P3_U3173) );
  NAND2_X1 U14613 ( .A1(n12198), .A2(n12695), .ZN(n12174) );
  AOI22_X1 U14614 ( .A1(n12194), .A2(n12714), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12173) );
  OAI211_X1 U14615 ( .C1(n12691), .C2(n12196), .A(n12174), .B(n12173), .ZN(
        n12175) );
  AOI21_X1 U14616 ( .B1(n12694), .B2(n12185), .A(n12175), .ZN(n12176) );
  OAI21_X1 U14617 ( .B1(n12177), .B2(n12187), .A(n12176), .ZN(P3_U3175) );
  XNOR2_X1 U14618 ( .A(n12179), .B(n12178), .ZN(n12188) );
  INV_X1 U14619 ( .A(n12180), .ZN(n12743) );
  NOR2_X1 U14620 ( .A1(n12181), .A2(n12743), .ZN(n12184) );
  NAND2_X1 U14621 ( .A1(n12194), .A2(n12349), .ZN(n12182) );
  NAND2_X1 U14622 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12557)
         );
  OAI211_X1 U14623 ( .C1(n12196), .C2(n12742), .A(n12182), .B(n12557), .ZN(
        n12183) );
  AOI211_X1 U14624 ( .C1(n12880), .C2(n12185), .A(n12184), .B(n12183), .ZN(
        n12186) );
  OAI21_X1 U14625 ( .B1(n12188), .B2(n12187), .A(n12186), .ZN(P3_U3178) );
  OAI21_X1 U14626 ( .B1(n12191), .B2(n12190), .A(n12189), .ZN(n12193) );
  NAND2_X1 U14627 ( .A1(n12193), .A2(n12192), .ZN(n12200) );
  AOI22_X1 U14628 ( .A1(n12433), .A2(n12194), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12195) );
  OAI21_X1 U14629 ( .B1(n12641), .B2(n12196), .A(n12195), .ZN(n12197) );
  AOI21_X1 U14630 ( .B1(n12642), .B2(n12198), .A(n12197), .ZN(n12199) );
  OAI211_X1 U14631 ( .C1(n12913), .C2(n12201), .A(n12200), .B(n12199), .ZN(
        P3_U3180) );
  NAND2_X1 U14632 ( .A1(n12202), .A2(n12411), .ZN(n12218) );
  NAND2_X1 U14633 ( .A1(n12203), .A2(n12212), .ZN(n12205) );
  OR2_X1 U14634 ( .A1(n12213), .A2(n15123), .ZN(n12204) );
  NAND2_X1 U14635 ( .A1(n12832), .A2(n12216), .ZN(n12413) );
  NAND2_X1 U14636 ( .A1(n12413), .A2(n12206), .ZN(n12407) );
  NAND2_X1 U14637 ( .A1(n12208), .A2(n12207), .ZN(n12211) );
  INV_X1 U14638 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n12209) );
  XNOR2_X1 U14639 ( .A(n12209), .B(P2_DATAO_REG_31__SCAN_IN), .ZN(n12210) );
  XNOR2_X1 U14640 ( .A(n12211), .B(n12210), .ZN(n12962) );
  NAND2_X1 U14641 ( .A1(n12962), .A2(n12212), .ZN(n12215) );
  INV_X1 U14642 ( .A(SI_31_), .ZN(n12966) );
  OR2_X1 U14643 ( .A1(n12213), .A2(n12966), .ZN(n12214) );
  NOR2_X1 U14644 ( .A1(n12600), .A2(n12602), .ZN(n12418) );
  AOI211_X1 U14645 ( .C1(n12602), .C2(n12832), .A(n12407), .B(n12418), .ZN(
        n12217) );
  NAND2_X1 U14646 ( .A1(n12600), .A2(n12602), .ZN(n12417) );
  INV_X1 U14647 ( .A(n12216), .ZN(n12429) );
  NAND2_X1 U14648 ( .A1(n12906), .A2(n12429), .ZN(n12410) );
  NAND2_X1 U14649 ( .A1(n12417), .A2(n12410), .ZN(n12221) );
  AOI22_X1 U14650 ( .A1(n12218), .A2(n12217), .B1(n12600), .B2(n12221), .ZN(
        n12220) );
  XNOR2_X1 U14651 ( .A(n12220), .B(n12219), .ZN(n12246) );
  INV_X1 U14652 ( .A(n12221), .ZN(n12241) );
  INV_X1 U14653 ( .A(n12222), .ZN(n12405) );
  INV_X1 U14654 ( .A(n12413), .ZN(n12238) );
  INV_X1 U14655 ( .A(n12659), .ZN(n12236) );
  XNOR2_X1 U14656 ( .A(n12705), .B(n12690), .ZN(n12703) );
  NAND2_X1 U14657 ( .A1(n12250), .A2(n12251), .ZN(n12692) );
  INV_X1 U14658 ( .A(n12720), .ZN(n12711) );
  XNOR2_X1 U14659 ( .A(n12935), .B(n12742), .ZN(n12729) );
  INV_X1 U14660 ( .A(n12788), .ZN(n12793) );
  INV_X1 U14661 ( .A(n12328), .ZN(n12223) );
  NAND4_X1 U14662 ( .A1(n12226), .A2(n12276), .A3(n12225), .A4(n12224), .ZN(
        n12228) );
  NOR4_X1 U14663 ( .A1(n12228), .A2(n15049), .A3(n15063), .A4(n12227), .ZN(
        n12229) );
  NAND4_X1 U14664 ( .A1(n12229), .A2(n12274), .A3(n12303), .A4(n12297), .ZN(
        n12230) );
  NOR4_X1 U14665 ( .A1(n12230), .A2(n12313), .A3(n12814), .A4(n14466), .ZN(
        n12231) );
  NAND4_X1 U14666 ( .A1(n12767), .A2(n12793), .A3(n12806), .A4(n12231), .ZN(
        n12232) );
  NOR3_X1 U14667 ( .A1(n12232), .A2(n12776), .A3(n12735), .ZN(n12233) );
  NAND4_X1 U14668 ( .A1(n12711), .A2(n12729), .A3(n12233), .A4(n12756), .ZN(
        n12234) );
  NOR4_X1 U14669 ( .A1(n7173), .A2(n12703), .A3(n12692), .A4(n12234), .ZN(
        n12235) );
  NAND4_X1 U14670 ( .A1(n12639), .A2(n12236), .A3(n12235), .A4(n12649), .ZN(
        n12237) );
  NOR4_X1 U14671 ( .A1(n12238), .A2(n12391), .A3(n12628), .A4(n12237), .ZN(
        n12240) );
  INV_X1 U14672 ( .A(n12418), .ZN(n12239) );
  NAND4_X1 U14673 ( .A1(n12241), .A2(n12405), .A3(n12240), .A4(n12239), .ZN(
        n12242) );
  XNOR2_X1 U14674 ( .A(n12242), .B(n12594), .ZN(n12243) );
  OAI22_X1 U14675 ( .A1(n12246), .A2(n12245), .B1(n12244), .B2(n12243), .ZN(
        n12421) );
  MUX2_X1 U14676 ( .A(n12433), .B(n12247), .S(n12415), .Z(n12249) );
  NAND2_X1 U14677 ( .A1(n12249), .A2(n12248), .ZN(n12387) );
  MUX2_X1 U14678 ( .A(n12251), .B(n12250), .S(n12402), .Z(n12377) );
  INV_X1 U14679 ( .A(n12252), .ZN(n12254) );
  NAND2_X1 U14680 ( .A1(n12254), .A2(n12424), .ZN(n12257) );
  NAND2_X1 U14681 ( .A1(n12254), .A2(n12253), .ZN(n12255) );
  NAND3_X1 U14682 ( .A1(n12262), .A2(n12415), .A3(n12255), .ZN(n12256) );
  OAI21_X1 U14683 ( .B1(n15063), .B2(n12257), .A(n12256), .ZN(n12261) );
  NAND2_X1 U14684 ( .A1(n12259), .A2(n12258), .ZN(n12260) );
  NAND2_X1 U14685 ( .A1(n12261), .A2(n12260), .ZN(n12265) );
  MUX2_X1 U14686 ( .A(n12263), .B(n12262), .S(n12402), .Z(n12264) );
  NAND3_X1 U14687 ( .A1(n12265), .A2(n15040), .A3(n12264), .ZN(n12269) );
  NAND2_X1 U14688 ( .A1(n12275), .A2(n12266), .ZN(n12267) );
  NAND2_X1 U14689 ( .A1(n12267), .A2(n12415), .ZN(n12268) );
  NAND2_X1 U14690 ( .A1(n12269), .A2(n12268), .ZN(n12273) );
  AOI21_X1 U14691 ( .B1(n12272), .B2(n12270), .A(n12415), .ZN(n12271) );
  AOI21_X1 U14692 ( .B1(n12273), .B2(n12272), .A(n12271), .ZN(n12278) );
  OAI21_X1 U14693 ( .B1(n12415), .B2(n12275), .A(n12274), .ZN(n12277) );
  OAI21_X1 U14694 ( .B1(n12278), .B2(n12277), .A(n12276), .ZN(n12287) );
  NAND2_X1 U14695 ( .A1(n12289), .A2(n12279), .ZN(n12282) );
  NAND2_X1 U14696 ( .A1(n12282), .A2(n12415), .ZN(n12286) );
  AND2_X1 U14697 ( .A1(n12446), .A2(n12280), .ZN(n12284) );
  NOR2_X1 U14698 ( .A1(n12282), .A2(n12281), .ZN(n12283) );
  MUX2_X1 U14699 ( .A(n12284), .B(n12283), .S(n12415), .Z(n12285) );
  AOI21_X1 U14700 ( .B1(n12287), .B2(n12286), .A(n12285), .ZN(n12293) );
  AOI21_X1 U14701 ( .B1(n12290), .B2(n12288), .A(n12415), .ZN(n12292) );
  MUX2_X1 U14702 ( .A(n12290), .B(n12289), .S(n12402), .Z(n12291) );
  OAI211_X1 U14703 ( .C1(n12293), .C2(n12292), .A(n7180), .B(n12291), .ZN(
        n12298) );
  MUX2_X1 U14704 ( .A(n12295), .B(n12294), .S(n12402), .Z(n12296) );
  NAND3_X1 U14705 ( .A1(n12298), .A2(n12297), .A3(n12296), .ZN(n12305) );
  INV_X1 U14706 ( .A(n12313), .ZN(n12304) );
  NAND2_X1 U14707 ( .A1(n12442), .A2(n12299), .ZN(n12301) );
  MUX2_X1 U14708 ( .A(n12301), .B(n12300), .S(n12415), .Z(n12302) );
  NAND4_X1 U14709 ( .A1(n12305), .A2(n12304), .A3(n12303), .A4(n12302), .ZN(
        n12317) );
  NAND2_X1 U14710 ( .A1(n12441), .A2(n12415), .ZN(n12309) );
  NAND2_X1 U14711 ( .A1(n12306), .A2(n12402), .ZN(n12308) );
  MUX2_X1 U14712 ( .A(n12309), .B(n12308), .S(n12307), .Z(n12314) );
  INV_X1 U14713 ( .A(n12814), .ZN(n12817) );
  MUX2_X1 U14714 ( .A(n12311), .B(n12310), .S(n12402), .Z(n12312) );
  OAI211_X1 U14715 ( .C1(n12314), .C2(n12313), .A(n12817), .B(n12312), .ZN(
        n12315) );
  INV_X1 U14716 ( .A(n12315), .ZN(n12316) );
  NAND2_X1 U14717 ( .A1(n12317), .A2(n12316), .ZN(n12325) );
  NAND3_X1 U14718 ( .A1(n12325), .A2(n12318), .A3(n12326), .ZN(n12319) );
  NAND2_X1 U14719 ( .A1(n12319), .A2(n12324), .ZN(n12322) );
  INV_X1 U14720 ( .A(n12320), .ZN(n12321) );
  AOI21_X1 U14721 ( .B1(n12322), .B2(n12806), .A(n12321), .ZN(n12331) );
  NAND3_X1 U14722 ( .A1(n12325), .A2(n12324), .A3(n12323), .ZN(n12327) );
  NAND2_X1 U14723 ( .A1(n12327), .A2(n12326), .ZN(n12329) );
  AOI21_X1 U14724 ( .B1(n12329), .B2(n12806), .A(n12328), .ZN(n12330) );
  MUX2_X1 U14725 ( .A(n12331), .B(n12330), .S(n12402), .Z(n12332) );
  NAND2_X1 U14726 ( .A1(n12332), .A2(n12793), .ZN(n12336) );
  MUX2_X1 U14727 ( .A(n12334), .B(n12333), .S(n12402), .Z(n12335) );
  NAND3_X1 U14728 ( .A1(n12336), .A2(n12781), .A3(n12335), .ZN(n12341) );
  OAI21_X1 U14729 ( .B1(n12790), .B2(n12337), .A(n12344), .ZN(n12338) );
  NAND2_X1 U14730 ( .A1(n12338), .A2(n12415), .ZN(n12340) );
  INV_X1 U14731 ( .A(n12343), .ZN(n12339) );
  AOI21_X1 U14732 ( .B1(n12341), .B2(n12340), .A(n12339), .ZN(n12346) );
  AOI21_X1 U14733 ( .B1(n12343), .B2(n12342), .A(n12415), .ZN(n12345) );
  OAI22_X1 U14734 ( .A1(n12346), .A2(n12345), .B1(n12415), .B2(n12344), .ZN(
        n12347) );
  NAND3_X1 U14735 ( .A1(n12347), .A2(n12740), .A3(n12756), .ZN(n12361) );
  INV_X1 U14736 ( .A(n12348), .ZN(n12943) );
  NAND3_X1 U14737 ( .A1(n12355), .A2(n12943), .A3(n12349), .ZN(n12351) );
  NAND2_X1 U14738 ( .A1(n12351), .A2(n12350), .ZN(n12352) );
  OR2_X1 U14739 ( .A1(n12362), .A2(n12352), .ZN(n12358) );
  INV_X1 U14740 ( .A(n12353), .ZN(n12354) );
  NAND2_X1 U14741 ( .A1(n12740), .A2(n12354), .ZN(n12356) );
  NAND3_X1 U14742 ( .A1(n12356), .A2(n12363), .A3(n12355), .ZN(n12357) );
  MUX2_X1 U14743 ( .A(n12358), .B(n12357), .S(n12415), .Z(n12359) );
  INV_X1 U14744 ( .A(n12359), .ZN(n12360) );
  NAND2_X1 U14745 ( .A1(n12361), .A2(n12360), .ZN(n12365) );
  MUX2_X1 U14746 ( .A(n12363), .B(n8697), .S(n12415), .Z(n12364) );
  NAND3_X1 U14747 ( .A1(n12365), .A2(n12711), .A3(n12364), .ZN(n12370) );
  INV_X1 U14748 ( .A(n12703), .ZN(n12369) );
  NAND2_X1 U14749 ( .A1(n12871), .A2(n12727), .ZN(n12367) );
  MUX2_X1 U14750 ( .A(n12367), .B(n12366), .S(n12402), .Z(n12368) );
  NAND3_X1 U14751 ( .A1(n12370), .A2(n12369), .A3(n12368), .ZN(n12375) );
  INV_X1 U14752 ( .A(n12692), .ZN(n12687) );
  NOR2_X1 U14753 ( .A1(n12705), .A2(n12415), .ZN(n12372) );
  NOR2_X1 U14754 ( .A1(n12714), .A2(n12402), .ZN(n12371) );
  OR3_X1 U14755 ( .A1(n12373), .A2(n12372), .A3(n12371), .ZN(n12374) );
  NAND3_X1 U14756 ( .A1(n12375), .A2(n12687), .A3(n12374), .ZN(n12376) );
  NAND3_X1 U14757 ( .A1(n12670), .A2(n12377), .A3(n12376), .ZN(n12381) );
  MUX2_X1 U14758 ( .A(n12379), .B(n12378), .S(n12415), .Z(n12380) );
  AND2_X1 U14759 ( .A1(n12381), .A2(n12380), .ZN(n12385) );
  MUX2_X1 U14760 ( .A(n12383), .B(n12382), .S(n12415), .Z(n12384) );
  OAI211_X1 U14761 ( .C1(n12385), .C2(n12659), .A(n12649), .B(n12384), .ZN(
        n12386) );
  NAND3_X1 U14762 ( .A1(n12639), .A2(n12387), .A3(n12386), .ZN(n12390) );
  OR3_X1 U14763 ( .A1(n12388), .A2(n12402), .A3(n12652), .ZN(n12389) );
  AOI21_X1 U14764 ( .B1(n12390), .B2(n12389), .A(n12628), .ZN(n12392) );
  NOR2_X1 U14765 ( .A1(n12392), .A2(n12391), .ZN(n12401) );
  INV_X1 U14766 ( .A(n12393), .ZN(n12394) );
  AOI21_X1 U14767 ( .B1(n12401), .B2(n12397), .A(n12394), .ZN(n12404) );
  NAND2_X1 U14768 ( .A1(n12396), .A2(n12395), .ZN(n12398) );
  NAND2_X1 U14769 ( .A1(n12398), .A2(n12397), .ZN(n12400) );
  AOI21_X1 U14770 ( .B1(n12401), .B2(n12400), .A(n12399), .ZN(n12403) );
  MUX2_X1 U14771 ( .A(n12404), .B(n12403), .S(n12402), .Z(n12406) );
  NAND2_X1 U14772 ( .A1(n12406), .A2(n12405), .ZN(n12412) );
  INV_X1 U14773 ( .A(n12407), .ZN(n12409) );
  INV_X1 U14774 ( .A(n12410), .ZN(n12408) );
  NAND3_X1 U14775 ( .A1(n12412), .A2(n12411), .A3(n12410), .ZN(n12414) );
  NAND2_X1 U14776 ( .A1(n12414), .A2(n12413), .ZN(n12416) );
  NOR2_X1 U14777 ( .A1(n12421), .A2(n12420), .ZN(n12428) );
  NOR3_X1 U14778 ( .A1(n12423), .A2(n12974), .A3(n12422), .ZN(n12426) );
  OAI21_X1 U14779 ( .B1(n12427), .B2(n12424), .A(P3_B_REG_SCAN_IN), .ZN(n12425) );
  OAI22_X1 U14780 ( .A1(n12428), .A2(n12427), .B1(n12426), .B2(n12425), .ZN(
        P3_U3296) );
  MUX2_X1 U14781 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(n12429), .S(P3_U3897), .Z(
        P3_U3521) );
  MUX2_X1 U14782 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(n12430), .S(P3_U3897), .Z(
        P3_U3520) );
  MUX2_X1 U14783 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12431), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14784 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12432), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14785 ( .A(n12433), .B(P3_DATAO_REG_25__SCAN_IN), .S(n12447), .Z(
        P3_U3516) );
  MUX2_X1 U14786 ( .A(n12434), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12447), .Z(
        P3_U3514) );
  MUX2_X1 U14787 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12435), .S(n12450), .Z(
        P3_U3513) );
  MUX2_X1 U14788 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12714), .S(n12450), .Z(
        P3_U3512) );
  MUX2_X1 U14789 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12436), .S(n12450), .Z(
        P3_U3511) );
  MUX2_X1 U14790 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n12713), .S(n12450), .Z(
        P3_U3510) );
  MUX2_X1 U14791 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12752), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14792 ( .A(n12751), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12447), .Z(
        P3_U3507) );
  MUX2_X1 U14793 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12437), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U14794 ( .A(n12802), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12447), .Z(
        P3_U3505) );
  MUX2_X1 U14795 ( .A(n12438), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12447), .Z(
        P3_U3504) );
  MUX2_X1 U14796 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n12439), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U14797 ( .A(n12440), .B(P3_DATAO_REG_10__SCAN_IN), .S(n12447), .Z(
        P3_U3501) );
  MUX2_X1 U14798 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n12441), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U14799 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12442), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14800 ( .A(n12443), .B(P3_DATAO_REG_7__SCAN_IN), .S(n12447), .Z(
        P3_U3498) );
  MUX2_X1 U14801 ( .A(n12444), .B(P3_DATAO_REG_6__SCAN_IN), .S(n12447), .Z(
        P3_U3497) );
  MUX2_X1 U14802 ( .A(n12445), .B(P3_DATAO_REG_5__SCAN_IN), .S(n12447), .Z(
        P3_U3496) );
  MUX2_X1 U14803 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12446), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14804 ( .A(n12448), .B(P3_DATAO_REG_3__SCAN_IN), .S(n12447), .Z(
        P3_U3494) );
  MUX2_X1 U14805 ( .A(n15068), .B(P3_DATAO_REG_2__SCAN_IN), .S(n12447), .Z(
        P3_U3493) );
  MUX2_X1 U14806 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n12449), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U14807 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n15065), .S(n12450), .Z(
        P3_U3491) );
  INV_X1 U14808 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n12805) );
  AOI21_X1 U14809 ( .B1(n12805), .B2(n12452), .A(n12472), .ZN(n12470) );
  XNOR2_X1 U14810 ( .A(n12483), .B(n12475), .ZN(n12455) );
  NAND2_X1 U14811 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n12455), .ZN(n12477) );
  OAI21_X1 U14812 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n12455), .A(n12477), 
        .ZN(n12468) );
  MUX2_X1 U14813 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12559), .Z(n12482) );
  XNOR2_X1 U14814 ( .A(n12482), .B(n12483), .ZN(n12459) );
  NAND2_X1 U14815 ( .A1(n12457), .A2(n12456), .ZN(n12460) );
  AND2_X1 U14816 ( .A1(n12459), .A2(n12460), .ZN(n12458) );
  NAND2_X1 U14817 ( .A1(n12461), .A2(n12458), .ZN(n12490) );
  INV_X1 U14818 ( .A(n12490), .ZN(n12463) );
  AOI21_X1 U14819 ( .B1(n12461), .B2(n12460), .A(n12459), .ZN(n12462) );
  OAI21_X1 U14820 ( .B1(n12463), .B2(n12462), .A(n14859), .ZN(n12466) );
  AOI21_X1 U14821 ( .B1(n14982), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n12464), 
        .ZN(n12465) );
  OAI211_X1 U14822 ( .C1(n14977), .C2(n12476), .A(n12466), .B(n12465), .ZN(
        n12467) );
  AOI21_X1 U14823 ( .B1(n12468), .B2(n14993), .A(n12467), .ZN(n12469) );
  OAI21_X1 U14824 ( .B1(n12470), .B2(n15005), .A(n12469), .ZN(P3_U3195) );
  NOR2_X1 U14825 ( .A1(n12483), .A2(n12471), .ZN(n12473) );
  NAND2_X1 U14826 ( .A1(n12495), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12507) );
  OAI21_X1 U14827 ( .B1(n12495), .B2(P3_REG2_REG_14__SCAN_IN), .A(n12507), 
        .ZN(n12485) );
  AOI21_X1 U14828 ( .B1(n12474), .B2(n12485), .A(n12501), .ZN(n12500) );
  NAND2_X1 U14829 ( .A1(n12476), .A2(n12475), .ZN(n12478) );
  NAND2_X1 U14830 ( .A1(n12478), .A2(n12477), .ZN(n12481) );
  INV_X1 U14831 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12898) );
  NAND2_X1 U14832 ( .A1(n12479), .A2(n12898), .ZN(n12480) );
  NAND2_X1 U14833 ( .A1(n12495), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12506) );
  AND2_X1 U14834 ( .A1(n12480), .A2(n12506), .ZN(n12487) );
  NAND2_X1 U14835 ( .A1(n12487), .A2(n12481), .ZN(n12504) );
  OAI21_X1 U14836 ( .B1(n12481), .B2(n12487), .A(n12504), .ZN(n12498) );
  INV_X1 U14837 ( .A(n12482), .ZN(n12484) );
  NAND2_X1 U14838 ( .A1(n12484), .A2(n12483), .ZN(n12489) );
  INV_X1 U14839 ( .A(n12485), .ZN(n12486) );
  MUX2_X1 U14840 ( .A(n12487), .B(n12486), .S(n12586), .Z(n12488) );
  NAND3_X1 U14841 ( .A1(n12490), .A2(n12489), .A3(n12488), .ZN(n12509) );
  INV_X1 U14842 ( .A(n12509), .ZN(n12492) );
  AOI21_X1 U14843 ( .B1(n12490), .B2(n12489), .A(n12488), .ZN(n12491) );
  NOR3_X1 U14844 ( .A1(n12492), .A2(n12491), .A3(n14999), .ZN(n12497) );
  AOI21_X1 U14845 ( .B1(n14982), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n12493), 
        .ZN(n12494) );
  OAI21_X1 U14846 ( .B1(n14977), .B2(n12495), .A(n12494), .ZN(n12496) );
  AOI211_X1 U14847 ( .C1(n12498), .C2(n14993), .A(n12497), .B(n12496), .ZN(
        n12499) );
  OAI21_X1 U14848 ( .B1(n12500), .B2(n15005), .A(n12499), .ZN(P3_U3196) );
  INV_X1 U14849 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12503) );
  AOI21_X1 U14850 ( .B1(n12503), .B2(n12502), .A(n12521), .ZN(n12519) );
  NAND2_X1 U14851 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n12505), .ZN(n12526) );
  OAI21_X1 U14852 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n12505), .A(n12526), 
        .ZN(n12517) );
  MUX2_X1 U14853 ( .A(n12507), .B(n12506), .S(n12559), .Z(n12508) );
  XNOR2_X1 U14854 ( .A(n12530), .B(n12525), .ZN(n12511) );
  MUX2_X1 U14855 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12559), .Z(n12510) );
  AOI21_X1 U14856 ( .B1(n12511), .B2(n12510), .A(n12531), .ZN(n12515) );
  INV_X1 U14857 ( .A(n14977), .ZN(n15010) );
  INV_X1 U14858 ( .A(n12525), .ZN(n12532) );
  INV_X1 U14859 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14341) );
  NOR2_X1 U14860 ( .A1(n15014), .A2(n14341), .ZN(n12512) );
  AOI211_X1 U14861 ( .C1(n15010), .C2(n12532), .A(n12513), .B(n12512), .ZN(
        n12514) );
  OAI21_X1 U14862 ( .B1(n12515), .B2(n14999), .A(n12514), .ZN(n12516) );
  AOI21_X1 U14863 ( .B1(n12517), .B2(n14993), .A(n12516), .ZN(n12518) );
  OAI21_X1 U14864 ( .B1(n12519), .B2(n15005), .A(n12518), .ZN(P3_U3197) );
  AND2_X1 U14865 ( .A1(n12525), .A2(n12520), .ZN(n12522) );
  INV_X1 U14866 ( .A(n12550), .ZN(n12547) );
  INV_X1 U14867 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12534) );
  AOI22_X1 U14868 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n12547), .B1(n12550), 
        .B2(n12534), .ZN(n12523) );
  AOI21_X1 U14869 ( .B1(n6464), .B2(n12523), .A(n12552), .ZN(n12545) );
  INV_X1 U14870 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n15253) );
  AOI22_X1 U14871 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12550), .B1(n12547), 
        .B2(n15253), .ZN(n12529) );
  NAND2_X1 U14872 ( .A1(n12525), .A2(n12524), .ZN(n12527) );
  NAND2_X1 U14873 ( .A1(n12527), .A2(n12526), .ZN(n12528) );
  NAND2_X1 U14874 ( .A1(n12529), .A2(n12528), .ZN(n12546) );
  OAI21_X1 U14875 ( .B1(n12529), .B2(n12528), .A(n12546), .ZN(n12543) );
  INV_X1 U14876 ( .A(n12530), .ZN(n12533) );
  MUX2_X1 U14877 ( .A(n12534), .B(n15253), .S(n12559), .Z(n12535) );
  NOR2_X1 U14878 ( .A1(n12547), .A2(n12535), .ZN(n12561) );
  NAND2_X1 U14879 ( .A1(n12547), .A2(n12535), .ZN(n12560) );
  INV_X1 U14880 ( .A(n12560), .ZN(n12536) );
  NOR2_X1 U14881 ( .A1(n12561), .A2(n12536), .ZN(n12537) );
  XNOR2_X1 U14882 ( .A(n12562), .B(n12537), .ZN(n12541) );
  INV_X1 U14883 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n15184) );
  NOR2_X1 U14884 ( .A1(n15014), .A2(n15184), .ZN(n12538) );
  AOI211_X1 U14885 ( .C1(n15010), .C2(n12547), .A(n12539), .B(n12538), .ZN(
        n12540) );
  OAI21_X1 U14886 ( .B1(n12541), .B2(n14999), .A(n12540), .ZN(n12542) );
  AOI21_X1 U14887 ( .B1(n12543), .B2(n14993), .A(n12542), .ZN(n12544) );
  OAI21_X1 U14888 ( .B1(n12545), .B2(n15005), .A(n12544), .ZN(P3_U3198) );
  XNOR2_X1 U14889 ( .A(n12582), .B(P3_REG1_REG_18__SCAN_IN), .ZN(n12578) );
  INV_X1 U14890 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12887) );
  INV_X1 U14891 ( .A(n12548), .ZN(n12549) );
  OAI22_X1 U14892 ( .A1(n14451), .A2(n12887), .B1(n14450), .B2(n12549), .ZN(
        n12579) );
  XOR2_X1 U14893 ( .A(n12578), .B(n12579), .Z(n12573) );
  INV_X1 U14894 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12744) );
  NOR2_X1 U14895 ( .A1(n12582), .A2(n12744), .ZN(n12574) );
  AOI21_X1 U14896 ( .B1(n12582), .B2(n12744), .A(n12574), .ZN(n12555) );
  AND2_X1 U14897 ( .A1(n12550), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n12551) );
  INV_X1 U14898 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14459) );
  OAI21_X1 U14899 ( .B1(n12555), .B2(n12554), .A(n12576), .ZN(n12556) );
  NAND2_X1 U14900 ( .A1(n12556), .A2(n14457), .ZN(n12571) );
  INV_X1 U14901 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n12558) );
  OAI21_X1 U14902 ( .B1(n15014), .B2(n12558), .A(n12557), .ZN(n12569) );
  MUX2_X1 U14903 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12559), .Z(n12566) );
  MUX2_X1 U14904 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12559), .Z(n12564) );
  OAI21_X1 U14905 ( .B1(n12562), .B2(n12561), .A(n12560), .ZN(n14453) );
  XOR2_X1 U14906 ( .A(n12564), .B(n14450), .Z(n14454) );
  NOR2_X1 U14907 ( .A1(n14453), .A2(n14454), .ZN(n14452) );
  AOI21_X1 U14908 ( .B1(n12564), .B2(n12563), .A(n14452), .ZN(n12583) );
  XNOR2_X1 U14909 ( .A(n12583), .B(n12582), .ZN(n12565) );
  NOR2_X1 U14910 ( .A1(n12565), .A2(n12566), .ZN(n12581) );
  AOI21_X1 U14911 ( .B1(n12566), .B2(n12565), .A(n12581), .ZN(n12567) );
  NOR2_X1 U14912 ( .A1(n12567), .A2(n14999), .ZN(n12568) );
  AOI211_X1 U14913 ( .C1(n15010), .C2(n12582), .A(n12569), .B(n12568), .ZN(
        n12570) );
  OAI211_X1 U14914 ( .C1(n12573), .C2(n12572), .A(n12571), .B(n12570), .ZN(
        P3_U3200) );
  INV_X1 U14915 ( .A(n12574), .ZN(n12575) );
  XNOR2_X1 U14916 ( .A(n12594), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12585) );
  AOI22_X1 U14917 ( .A1(n12579), .A2(n12578), .B1(P3_REG1_REG_18__SCAN_IN), 
        .B2(n12577), .ZN(n12580) );
  XNOR2_X1 U14918 ( .A(n12594), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12584) );
  XNOR2_X1 U14919 ( .A(n12580), .B(n12584), .ZN(n12597) );
  AOI21_X1 U14920 ( .B1(n12583), .B2(n12582), .A(n12581), .ZN(n12590) );
  INV_X1 U14921 ( .A(n12584), .ZN(n12588) );
  INV_X1 U14922 ( .A(n12585), .ZN(n12587) );
  MUX2_X1 U14923 ( .A(n12588), .B(n12587), .S(n12586), .Z(n12589) );
  XNOR2_X1 U14924 ( .A(n12590), .B(n12589), .ZN(n12591) );
  NOR2_X1 U14925 ( .A1(n12591), .A2(n14999), .ZN(n12596) );
  NAND2_X1 U14926 ( .A1(n14982), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12592) );
  OAI211_X1 U14927 ( .C1(n14977), .C2(n12594), .A(n12593), .B(n12592), .ZN(
        n12595) );
  OAI21_X1 U14928 ( .B1(n12599), .B2(n15005), .A(n12598), .ZN(P3_U3201) );
  NAND2_X1 U14929 ( .A1(n12603), .A2(n10664), .ZN(n12609) );
  OAI21_X1 U14930 ( .B1(n12901), .B2(n12826), .A(n12609), .ZN(n12605) );
  AOI21_X1 U14931 ( .B1(P3_REG2_REG_31__SCAN_IN), .B2(n12826), .A(n12605), 
        .ZN(n12604) );
  OAI21_X1 U14932 ( .B1(n12903), .B2(n12824), .A(n12604), .ZN(P3_U3202) );
  AOI21_X1 U14933 ( .B1(P3_REG2_REG_30__SCAN_IN), .B2(n12826), .A(n12605), 
        .ZN(n12606) );
  OAI21_X1 U14934 ( .B1(n12906), .B2(n12824), .A(n12606), .ZN(P3_U3203) );
  INV_X1 U14935 ( .A(n12607), .ZN(n12615) );
  NAND2_X1 U14936 ( .A1(n12608), .A2(n15034), .ZN(n12610) );
  OAI211_X1 U14937 ( .C1(n15036), .C2(n12611), .A(n12610), .B(n12609), .ZN(
        n12612) );
  AOI21_X1 U14938 ( .B1(n12613), .B2(n15036), .A(n12612), .ZN(n12614) );
  OAI21_X1 U14939 ( .B1(n12615), .B2(n12829), .A(n12614), .ZN(P3_U3204) );
  INV_X1 U14940 ( .A(n12616), .ZN(n12624) );
  OAI22_X1 U14941 ( .A1(n12618), .A2(n12822), .B1(n15036), .B2(n12617), .ZN(
        n12619) );
  AOI21_X1 U14942 ( .B1(n12620), .B2(n15034), .A(n12619), .ZN(n12623) );
  NAND2_X1 U14943 ( .A1(n12621), .A2(n15036), .ZN(n12622) );
  OAI211_X1 U14944 ( .C1(n12624), .C2(n12829), .A(n12623), .B(n12622), .ZN(
        P3_U3205) );
  AOI21_X1 U14945 ( .B1(n12626), .B2(n12628), .A(n12625), .ZN(n12841) );
  NAND2_X1 U14946 ( .A1(n12842), .A2(n15036), .ZN(n12636) );
  INV_X1 U14947 ( .A(n12630), .ZN(n12632) );
  OAI22_X1 U14948 ( .A1(n12632), .A2(n12822), .B1(n15036), .B2(n12631), .ZN(
        n12633) );
  AOI21_X1 U14949 ( .B1(n12634), .B2(n15034), .A(n12633), .ZN(n12635) );
  OAI211_X1 U14950 ( .C1(n12841), .C2(n12829), .A(n12636), .B(n12635), .ZN(
        P3_U3206) );
  XNOR2_X1 U14951 ( .A(n12637), .B(n12639), .ZN(n12847) );
  INV_X1 U14952 ( .A(n12847), .ZN(n12646) );
  XOR2_X1 U14953 ( .A(n12639), .B(n12638), .Z(n12640) );
  OAI222_X1 U14954 ( .A1(n15044), .A2(n12641), .B1(n15046), .B2(n12662), .C1(
        n12640), .C2(n15072), .ZN(n12846) );
  AOI22_X1 U14955 ( .A1(n12642), .A2(n10664), .B1(n12826), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n12643) );
  OAI21_X1 U14956 ( .B1(n12913), .B2(n12824), .A(n12643), .ZN(n12644) );
  AOI21_X1 U14957 ( .B1(n12846), .B2(n15036), .A(n12644), .ZN(n12645) );
  OAI21_X1 U14958 ( .B1(n12829), .B2(n12646), .A(n12645), .ZN(P3_U3207) );
  XNOR2_X1 U14959 ( .A(n12648), .B(n12647), .ZN(n12851) );
  INV_X1 U14960 ( .A(n12851), .ZN(n12657) );
  XNOR2_X1 U14961 ( .A(n12650), .B(n12649), .ZN(n12651) );
  OAI222_X1 U14962 ( .A1(n15044), .A2(n12652), .B1(n15046), .B2(n12676), .C1(
        n15072), .C2(n12651), .ZN(n12850) );
  AOI22_X1 U14963 ( .A1(n12653), .A2(n10664), .B1(n12826), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n12654) );
  OAI21_X1 U14964 ( .B1(n12917), .B2(n12824), .A(n12654), .ZN(n12655) );
  AOI21_X1 U14965 ( .B1(n12850), .B2(n15036), .A(n12655), .ZN(n12656) );
  OAI21_X1 U14966 ( .B1(n12657), .B2(n12829), .A(n12656), .ZN(P3_U3208) );
  AOI21_X1 U14967 ( .B1(n12659), .B2(n12658), .A(n6480), .ZN(n12854) );
  XNOR2_X1 U14968 ( .A(n12660), .B(n12659), .ZN(n12661) );
  OAI222_X1 U14969 ( .A1(n15044), .A2(n12662), .B1(n15046), .B2(n12691), .C1(
        n12661), .C2(n15072), .ZN(n12855) );
  NAND2_X1 U14970 ( .A1(n12855), .A2(n15036), .ZN(n12669) );
  INV_X1 U14971 ( .A(n12663), .ZN(n12665) );
  OAI22_X1 U14972 ( .A1(n12665), .A2(n12822), .B1(n15036), .B2(n12664), .ZN(
        n12666) );
  AOI21_X1 U14973 ( .B1(n12667), .B2(n15034), .A(n12666), .ZN(n12668) );
  OAI211_X1 U14974 ( .C1(n12854), .C2(n12829), .A(n12669), .B(n12668), .ZN(
        P3_U3209) );
  OR2_X1 U14975 ( .A1(n12671), .A2(n12670), .ZN(n12672) );
  NAND2_X1 U14976 ( .A1(n12673), .A2(n12672), .ZN(n12860) );
  XNOR2_X1 U14977 ( .A(n12674), .B(n7173), .ZN(n12675) );
  NAND2_X1 U14978 ( .A1(n12675), .A2(n15051), .ZN(n12679) );
  OAI22_X1 U14979 ( .A1(n12676), .A2(n15044), .B1(n12702), .B2(n15046), .ZN(
        n12677) );
  INV_X1 U14980 ( .A(n12677), .ZN(n12678) );
  NAND2_X1 U14981 ( .A1(n12679), .A2(n12678), .ZN(n12862) );
  NAND2_X1 U14982 ( .A1(n12862), .A2(n15036), .ZN(n12686) );
  INV_X1 U14983 ( .A(n12680), .ZN(n12682) );
  OAI22_X1 U14984 ( .A1(n12682), .A2(n12822), .B1(n15036), .B2(n12681), .ZN(
        n12683) );
  AOI21_X1 U14985 ( .B1(n12684), .B2(n15034), .A(n12683), .ZN(n12685) );
  OAI211_X1 U14986 ( .C1(n12860), .C2(n12829), .A(n12686), .B(n12685), .ZN(
        P3_U3210) );
  XNOR2_X1 U14987 ( .A(n12688), .B(n12687), .ZN(n12689) );
  OAI222_X1 U14988 ( .A1(n15044), .A2(n12691), .B1(n15046), .B2(n12690), .C1(
        n15072), .C2(n12689), .ZN(n12863) );
  INV_X1 U14989 ( .A(n12863), .ZN(n12699) );
  XNOR2_X1 U14990 ( .A(n12693), .B(n12692), .ZN(n12864) );
  INV_X1 U14991 ( .A(n12694), .ZN(n12926) );
  AOI22_X1 U14992 ( .A1(n12826), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n10664), 
        .B2(n12695), .ZN(n12696) );
  OAI21_X1 U14993 ( .B1(n12926), .B2(n12824), .A(n12696), .ZN(n12697) );
  AOI21_X1 U14994 ( .B1(n12864), .B2(n14476), .A(n12697), .ZN(n12698) );
  OAI21_X1 U14995 ( .B1(n12699), .B2(n12826), .A(n12698), .ZN(P3_U3211) );
  XNOR2_X1 U14996 ( .A(n12700), .B(n12703), .ZN(n12701) );
  OAI222_X1 U14997 ( .A1(n15044), .A2(n12702), .B1(n15046), .B2(n12727), .C1(
        n15072), .C2(n12701), .ZN(n12867) );
  INV_X1 U14998 ( .A(n12867), .ZN(n12710) );
  XNOR2_X1 U14999 ( .A(n12704), .B(n12703), .ZN(n12868) );
  INV_X1 U15000 ( .A(n12705), .ZN(n12930) );
  AOI22_X1 U15001 ( .A1(n12826), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n10664), 
        .B2(n12706), .ZN(n12707) );
  OAI21_X1 U15002 ( .B1(n12930), .B2(n12824), .A(n12707), .ZN(n12708) );
  AOI21_X1 U15003 ( .B1(n12868), .B2(n14476), .A(n12708), .ZN(n12709) );
  OAI21_X1 U15004 ( .B1(n12710), .B2(n12826), .A(n12709), .ZN(P3_U3212) );
  XNOR2_X1 U15005 ( .A(n12712), .B(n12711), .ZN(n12715) );
  AOI222_X1 U15006 ( .A1(n15051), .A2(n12715), .B1(n12714), .B2(n15067), .C1(
        n12713), .C2(n15066), .ZN(n12875) );
  INV_X1 U15007 ( .A(n12716), .ZN(n12717) );
  OAI22_X1 U15008 ( .A1(n15036), .A2(n12718), .B1(n12717), .B2(n12822), .ZN(
        n12719) );
  AOI21_X1 U15009 ( .B1(n12871), .B2(n15034), .A(n12719), .ZN(n12723) );
  NAND2_X1 U15010 ( .A1(n12721), .A2(n12720), .ZN(n12872) );
  NAND3_X1 U15011 ( .A1(n12873), .A2(n12872), .A3(n14476), .ZN(n12722) );
  OAI211_X1 U15012 ( .C1(n12875), .C2(n12826), .A(n12723), .B(n12722), .ZN(
        P3_U3213) );
  XNOR2_X1 U15013 ( .A(n12724), .B(n12729), .ZN(n12725) );
  OAI222_X1 U15014 ( .A1(n15044), .A2(n12727), .B1(n15046), .B2(n12726), .C1(
        n15072), .C2(n12725), .ZN(n12877) );
  INV_X1 U15015 ( .A(n12877), .ZN(n12734) );
  XOR2_X1 U15016 ( .A(n12729), .B(n12728), .Z(n12878) );
  AOI22_X1 U15017 ( .A1(n12826), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n10664), 
        .B2(n12730), .ZN(n12731) );
  OAI21_X1 U15018 ( .B1(n12935), .B2(n12824), .A(n12731), .ZN(n12732) );
  AOI21_X1 U15019 ( .B1(n12878), .B2(n14476), .A(n12732), .ZN(n12733) );
  OAI21_X1 U15020 ( .B1(n12734), .B2(n12826), .A(n12733), .ZN(P3_U3214) );
  NAND2_X1 U15021 ( .A1(n12736), .A2(n12735), .ZN(n12737) );
  INV_X1 U15022 ( .A(n12882), .ZN(n12748) );
  AOI21_X1 U15023 ( .B1(n12740), .B2(n12739), .A(n6533), .ZN(n12741) );
  OAI222_X1 U15024 ( .A1(n15044), .A2(n12742), .B1(n15046), .B2(n12765), .C1(
        n15072), .C2(n12741), .ZN(n12881) );
  NAND2_X1 U15025 ( .A1(n12881), .A2(n15036), .ZN(n12747) );
  OAI22_X1 U15026 ( .A1(n15036), .A2(n12744), .B1(n12743), .B2(n12822), .ZN(
        n12745) );
  AOI21_X1 U15027 ( .B1(n12880), .B2(n15034), .A(n12745), .ZN(n12746) );
  OAI211_X1 U15028 ( .C1(n12748), .C2(n12829), .A(n12747), .B(n12746), .ZN(
        P3_U3215) );
  OAI211_X1 U15029 ( .C1(n12750), .C2(n8872), .A(n12749), .B(n15051), .ZN(
        n12754) );
  AOI22_X1 U15030 ( .A1(n12752), .A2(n15067), .B1(n15066), .B2(n12751), .ZN(
        n12753) );
  NAND2_X1 U15031 ( .A1(n12754), .A2(n12753), .ZN(n12885) );
  INV_X1 U15032 ( .A(n12885), .ZN(n12762) );
  OAI21_X1 U15033 ( .B1(n12757), .B2(n12756), .A(n12755), .ZN(n12886) );
  AOI22_X1 U15034 ( .A1(n12826), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n10664), 
        .B2(n12758), .ZN(n12759) );
  OAI21_X1 U15035 ( .B1(n12943), .B2(n12824), .A(n12759), .ZN(n12760) );
  AOI21_X1 U15036 ( .B1(n12886), .B2(n14476), .A(n12760), .ZN(n12761) );
  OAI21_X1 U15037 ( .B1(n12762), .B2(n12826), .A(n12761), .ZN(P3_U3216) );
  XOR2_X1 U15038 ( .A(n12767), .B(n12763), .Z(n12764) );
  OAI222_X1 U15039 ( .A1(n15044), .A2(n12765), .B1(n15046), .B2(n12790), .C1(
        n12764), .C2(n15072), .ZN(n12889) );
  INV_X1 U15040 ( .A(n12889), .ZN(n12774) );
  OAI21_X1 U15041 ( .B1(n12768), .B2(n12767), .A(n12766), .ZN(n12890) );
  INV_X1 U15042 ( .A(n12769), .ZN(n12947) );
  AOI22_X1 U15043 ( .A1(n12826), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n10664), 
        .B2(n12770), .ZN(n12771) );
  OAI21_X1 U15044 ( .B1(n12947), .B2(n12824), .A(n12771), .ZN(n12772) );
  AOI21_X1 U15045 ( .B1(n12890), .B2(n14476), .A(n12772), .ZN(n12773) );
  OAI21_X1 U15046 ( .B1(n12774), .B2(n12826), .A(n12773), .ZN(P3_U3217) );
  XNOR2_X1 U15047 ( .A(n12775), .B(n12776), .ZN(n12777) );
  OAI222_X1 U15048 ( .A1(n15044), .A2(n12779), .B1(n15046), .B2(n12778), .C1(
        n15072), .C2(n12777), .ZN(n12892) );
  INV_X1 U15049 ( .A(n12892), .ZN(n12786) );
  XNOR2_X1 U15050 ( .A(n12780), .B(n12781), .ZN(n12893) );
  AOI22_X1 U15051 ( .A1(n12826), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n10664), 
        .B2(n12782), .ZN(n12783) );
  OAI21_X1 U15052 ( .B1(n12951), .B2(n12824), .A(n12783), .ZN(n12784) );
  AOI21_X1 U15053 ( .B1(n12893), .B2(n14476), .A(n12784), .ZN(n12785) );
  OAI21_X1 U15054 ( .B1(n12786), .B2(n12826), .A(n12785), .ZN(P3_U3218) );
  XNOR2_X1 U15055 ( .A(n12787), .B(n12788), .ZN(n12789) );
  OAI222_X1 U15056 ( .A1(n15044), .A2(n12790), .B1(n15046), .B2(n14470), .C1(
        n12789), .C2(n15072), .ZN(n12896) );
  INV_X1 U15057 ( .A(n12896), .ZN(n12799) );
  OAI21_X1 U15058 ( .B1(n7529), .B2(n12793), .A(n12792), .ZN(n12897) );
  INV_X1 U15059 ( .A(n12794), .ZN(n12956) );
  AOI22_X1 U15060 ( .A1(n12826), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n10664), 
        .B2(n12795), .ZN(n12796) );
  OAI21_X1 U15061 ( .B1(n12956), .B2(n12824), .A(n12796), .ZN(n12797) );
  AOI21_X1 U15062 ( .B1(n12897), .B2(n14476), .A(n12797), .ZN(n12798) );
  OAI21_X1 U15063 ( .B1(n12799), .B2(n12826), .A(n12798), .ZN(P3_U3219) );
  XNOR2_X1 U15064 ( .A(n12800), .B(n12806), .ZN(n12803) );
  AOI222_X1 U15065 ( .A1(n15051), .A2(n12803), .B1(n12802), .B2(n15067), .C1(
        n12801), .C2(n15066), .ZN(n14481) );
  OAI22_X1 U15066 ( .A1(n15036), .A2(n12805), .B1(n12804), .B2(n12822), .ZN(
        n12809) );
  XOR2_X1 U15067 ( .A(n12807), .B(n12806), .Z(n14480) );
  NOR2_X1 U15068 ( .A1(n14480), .A2(n12829), .ZN(n12808) );
  AOI211_X1 U15069 ( .C1(n15034), .C2(n14484), .A(n12809), .B(n12808), .ZN(
        n12810) );
  OAI21_X1 U15070 ( .B1(n12826), .B2(n14481), .A(n12810), .ZN(P3_U3220) );
  INV_X1 U15071 ( .A(n12811), .ZN(n12812) );
  AOI21_X1 U15072 ( .B1(n12814), .B2(n12813), .A(n12812), .ZN(n14495) );
  INV_X1 U15073 ( .A(n12815), .ZN(n12816) );
  AOI21_X1 U15074 ( .B1(n12817), .B2(n6549), .A(n12816), .ZN(n12818) );
  OAI222_X1 U15075 ( .A1(n15044), .A2(n12820), .B1(n15046), .B2(n12819), .C1(
        n15072), .C2(n12818), .ZN(n14497) );
  NAND2_X1 U15076 ( .A1(n14497), .A2(n15036), .ZN(n12828) );
  INV_X1 U15077 ( .A(n12821), .ZN(n12823) );
  OAI22_X1 U15078 ( .A1(n12824), .A2(n14493), .B1(n12823), .B2(n12822), .ZN(
        n12825) );
  AOI21_X1 U15079 ( .B1(n12826), .B2(P3_REG2_REG_11__SCAN_IN), .A(n12825), 
        .ZN(n12827) );
  OAI211_X1 U15080 ( .C1(n14495), .C2(n12829), .A(n12828), .B(n12827), .ZN(
        P3_U3222) );
  NOR2_X1 U15081 ( .A1(n12901), .A2(n15114), .ZN(n12833) );
  AOI21_X1 U15082 ( .B1(P3_REG1_REG_31__SCAN_IN), .B2(n15114), .A(n12833), 
        .ZN(n12830) );
  OAI21_X1 U15083 ( .B1(n12903), .B2(n12900), .A(n12830), .ZN(P3_U3490) );
  INV_X1 U15084 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n12836) );
  INV_X1 U15085 ( .A(n12900), .ZN(n12831) );
  NAND2_X1 U15086 ( .A1(n12832), .A2(n12831), .ZN(n12835) );
  INV_X1 U15087 ( .A(n12833), .ZN(n12834) );
  OAI211_X1 U15088 ( .C1(n15117), .C2(n12836), .A(n12835), .B(n12834), .ZN(
        P3_U3489) );
  INV_X1 U15089 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n12838) );
  MUX2_X1 U15090 ( .A(n12838), .B(n12837), .S(n15117), .Z(n12839) );
  OAI21_X1 U15091 ( .B1(n12840), .B2(n12900), .A(n12839), .ZN(P3_U3487) );
  INV_X1 U15092 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n12844) );
  INV_X1 U15093 ( .A(n12841), .ZN(n12843) );
  MUX2_X1 U15094 ( .A(n12844), .B(n12907), .S(n15117), .Z(n12845) );
  OAI21_X1 U15095 ( .B1(n12909), .B2(n12900), .A(n12845), .ZN(P3_U3486) );
  INV_X1 U15096 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12848) );
  AOI21_X1 U15097 ( .B1(n12847), .B2(n14490), .A(n12846), .ZN(n12910) );
  MUX2_X1 U15098 ( .A(n12848), .B(n12910), .S(n15117), .Z(n12849) );
  OAI21_X1 U15099 ( .B1(n12913), .B2(n12900), .A(n12849), .ZN(P3_U3485) );
  INV_X1 U15100 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n12852) );
  AOI21_X1 U15101 ( .B1(n14490), .B2(n12851), .A(n12850), .ZN(n12914) );
  MUX2_X1 U15102 ( .A(n12852), .B(n12914), .S(n15117), .Z(n12853) );
  OAI21_X1 U15103 ( .B1(n12917), .B2(n12900), .A(n12853), .ZN(P3_U3484) );
  INV_X1 U15104 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12857) );
  INV_X1 U15105 ( .A(n12854), .ZN(n12856) );
  AOI21_X1 U15106 ( .B1(n14490), .B2(n12856), .A(n12855), .ZN(n12918) );
  MUX2_X1 U15107 ( .A(n12857), .B(n12918), .S(n15117), .Z(n12858) );
  OAI21_X1 U15108 ( .B1(n12921), .B2(n12900), .A(n12858), .ZN(P3_U3483) );
  OAI22_X1 U15109 ( .A1(n12860), .A2(n14494), .B1(n12859), .B2(n15100), .ZN(
        n12861) );
  MUX2_X1 U15110 ( .A(P3_REG1_REG_23__SCAN_IN), .B(n12922), .S(n15117), .Z(
        P3_U3482) );
  INV_X1 U15111 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12865) );
  AOI21_X1 U15112 ( .B1(n14490), .B2(n12864), .A(n12863), .ZN(n12923) );
  MUX2_X1 U15113 ( .A(n12865), .B(n12923), .S(n15117), .Z(n12866) );
  OAI21_X1 U15114 ( .B1(n12926), .B2(n12900), .A(n12866), .ZN(P3_U3481) );
  INV_X1 U15115 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12869) );
  AOI21_X1 U15116 ( .B1(n12868), .B2(n14490), .A(n12867), .ZN(n12927) );
  MUX2_X1 U15117 ( .A(n12869), .B(n12927), .S(n15117), .Z(n12870) );
  OAI21_X1 U15118 ( .B1(n12930), .B2(n12900), .A(n12870), .ZN(P3_U3480) );
  INV_X1 U15119 ( .A(n12871), .ZN(n12876) );
  NAND3_X1 U15120 ( .A1(n12873), .A2(n14490), .A3(n12872), .ZN(n12874) );
  OAI211_X1 U15121 ( .C1(n12876), .C2(n15100), .A(n12875), .B(n12874), .ZN(
        n12931) );
  MUX2_X1 U15122 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n12931), .S(n15117), .Z(
        P3_U3479) );
  INV_X1 U15123 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n15255) );
  AOI21_X1 U15124 ( .B1(n14490), .B2(n12878), .A(n12877), .ZN(n12932) );
  MUX2_X1 U15125 ( .A(n15255), .B(n12932), .S(n15117), .Z(n12879) );
  OAI21_X1 U15126 ( .B1(n12900), .B2(n12935), .A(n12879), .ZN(P3_U3478) );
  INV_X1 U15127 ( .A(n12880), .ZN(n12939) );
  INV_X1 U15128 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12883) );
  AOI21_X1 U15129 ( .B1(n12882), .B2(n14490), .A(n12881), .ZN(n12936) );
  MUX2_X1 U15130 ( .A(n12883), .B(n12936), .S(n15117), .Z(n12884) );
  OAI21_X1 U15131 ( .B1(n12939), .B2(n12900), .A(n12884), .ZN(P3_U3477) );
  AOI21_X1 U15132 ( .B1(n14490), .B2(n12886), .A(n12885), .ZN(n12940) );
  MUX2_X1 U15133 ( .A(n12887), .B(n12940), .S(n15117), .Z(n12888) );
  OAI21_X1 U15134 ( .B1(n12943), .B2(n12900), .A(n12888), .ZN(P3_U3476) );
  AOI21_X1 U15135 ( .B1(n14490), .B2(n12890), .A(n12889), .ZN(n12944) );
  MUX2_X1 U15136 ( .A(n15253), .B(n12944), .S(n15117), .Z(n12891) );
  OAI21_X1 U15137 ( .B1(n12947), .B2(n12900), .A(n12891), .ZN(P3_U3475) );
  INV_X1 U15138 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12894) );
  AOI21_X1 U15139 ( .B1(n14490), .B2(n12893), .A(n12892), .ZN(n12948) );
  MUX2_X1 U15140 ( .A(n12894), .B(n12948), .S(n15117), .Z(n12895) );
  OAI21_X1 U15141 ( .B1(n12951), .B2(n12900), .A(n12895), .ZN(P3_U3474) );
  AOI21_X1 U15142 ( .B1(n14490), .B2(n12897), .A(n12896), .ZN(n12952) );
  MUX2_X1 U15143 ( .A(n12898), .B(n12952), .S(n15117), .Z(n12899) );
  OAI21_X1 U15144 ( .B1(n12956), .B2(n12900), .A(n12899), .ZN(P3_U3473) );
  NOR2_X1 U15145 ( .A1(n12901), .A2(n15110), .ZN(n12904) );
  AOI21_X1 U15146 ( .B1(n15110), .B2(P3_REG0_REG_31__SCAN_IN), .A(n12904), 
        .ZN(n12902) );
  OAI21_X1 U15147 ( .B1(n12903), .B2(n12955), .A(n12902), .ZN(P3_U3458) );
  AOI21_X1 U15148 ( .B1(n15110), .B2(P3_REG0_REG_30__SCAN_IN), .A(n12904), 
        .ZN(n12905) );
  OAI21_X1 U15149 ( .B1(n12906), .B2(n12955), .A(n12905), .ZN(P3_U3457) );
  INV_X1 U15150 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12911) );
  MUX2_X1 U15151 ( .A(n12911), .B(n12910), .S(n15108), .Z(n12912) );
  OAI21_X1 U15152 ( .B1(n12913), .B2(n12955), .A(n12912), .ZN(P3_U3453) );
  INV_X1 U15153 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n12915) );
  MUX2_X1 U15154 ( .A(n12915), .B(n12914), .S(n15108), .Z(n12916) );
  OAI21_X1 U15155 ( .B1(n12917), .B2(n12955), .A(n12916), .ZN(P3_U3452) );
  INV_X1 U15156 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n12919) );
  MUX2_X1 U15157 ( .A(n12919), .B(n12918), .S(n15108), .Z(n12920) );
  OAI21_X1 U15158 ( .B1(n12921), .B2(n12955), .A(n12920), .ZN(P3_U3451) );
  MUX2_X1 U15159 ( .A(n12922), .B(P3_REG0_REG_23__SCAN_IN), .S(n15110), .Z(
        P3_U3450) );
  INV_X1 U15160 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12924) );
  MUX2_X1 U15161 ( .A(n12924), .B(n12923), .S(n15108), .Z(n12925) );
  OAI21_X1 U15162 ( .B1(n12926), .B2(n12955), .A(n12925), .ZN(P3_U3449) );
  INV_X1 U15163 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12928) );
  MUX2_X1 U15164 ( .A(n12928), .B(n12927), .S(n15108), .Z(n12929) );
  OAI21_X1 U15165 ( .B1(n12930), .B2(n12955), .A(n12929), .ZN(P3_U3448) );
  MUX2_X1 U15166 ( .A(P3_REG0_REG_20__SCAN_IN), .B(n12931), .S(n15108), .Z(
        P3_U3447) );
  INV_X1 U15167 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n12933) );
  MUX2_X1 U15168 ( .A(n12933), .B(n12932), .S(n15108), .Z(n12934) );
  OAI21_X1 U15169 ( .B1(n12955), .B2(n12935), .A(n12934), .ZN(P3_U3446) );
  INV_X1 U15170 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n12937) );
  MUX2_X1 U15171 ( .A(n12937), .B(n12936), .S(n15108), .Z(n12938) );
  OAI21_X1 U15172 ( .B1(n12939), .B2(n12955), .A(n12938), .ZN(P3_U3444) );
  INV_X1 U15173 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n12941) );
  MUX2_X1 U15174 ( .A(n12941), .B(n12940), .S(n15108), .Z(n12942) );
  OAI21_X1 U15175 ( .B1(n12943), .B2(n12955), .A(n12942), .ZN(P3_U3441) );
  INV_X1 U15176 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n12945) );
  MUX2_X1 U15177 ( .A(n12945), .B(n12944), .S(n15108), .Z(n12946) );
  OAI21_X1 U15178 ( .B1(n12947), .B2(n12955), .A(n12946), .ZN(P3_U3438) );
  INV_X1 U15179 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n12949) );
  MUX2_X1 U15180 ( .A(n12949), .B(n12948), .S(n15108), .Z(n12950) );
  OAI21_X1 U15181 ( .B1(n12951), .B2(n12955), .A(n12950), .ZN(P3_U3435) );
  INV_X1 U15182 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n12953) );
  MUX2_X1 U15183 ( .A(n12953), .B(n12952), .S(n15108), .Z(n12954) );
  OAI21_X1 U15184 ( .B1(n12956), .B2(n12955), .A(n12954), .ZN(P3_U3432) );
  MUX2_X1 U15185 ( .A(n12958), .B(P3_D_REG_1__SCAN_IN), .S(n12957), .Z(
        P3_U3377) );
  MUX2_X1 U15186 ( .A(P3_D_REG_0__SCAN_IN), .B(n12960), .S(n12959), .Z(
        P3_U3376) );
  NAND2_X1 U15187 ( .A1(n12962), .A2(n12961), .ZN(n12965) );
  OR4_X1 U15188 ( .A1(n6793), .A2(P3_IR_REG_30__SCAN_IN), .A3(P3_U3151), .A4(
        n6991), .ZN(n12964) );
  OAI211_X1 U15189 ( .C1(n12966), .C2(n12973), .A(n12965), .B(n12964), .ZN(
        P3_U3264) );
  INV_X1 U15190 ( .A(n12967), .ZN(n12969) );
  OAI222_X1 U15191 ( .A1(n14410), .A2(n12969), .B1(n12968), .B2(P3_U3151), 
        .C1(n15242), .C2(n12973), .ZN(P3_U3266) );
  INV_X1 U15192 ( .A(n12970), .ZN(n12971) );
  MUX2_X1 U15193 ( .A(n12975), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  AOI211_X1 U15194 ( .C1(n12976), .C2(n12978), .A(n13073), .B(n12977), .ZN(
        n12979) );
  INV_X1 U15195 ( .A(n12979), .ZN(n12983) );
  INV_X1 U15196 ( .A(n13243), .ZN(n13202) );
  AOI22_X1 U15197 ( .A1(n13202), .A2(n14522), .B1(n14524), .B2(n13247), .ZN(
        n13328) );
  OAI22_X1 U15198 ( .A1(n13091), .A2(n13328), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12980), .ZN(n12981) );
  AOI21_X1 U15199 ( .B1(n13331), .B2(n13093), .A(n12981), .ZN(n12982) );
  OAI211_X1 U15200 ( .C1(n7069), .C2(n13096), .A(n12983), .B(n12982), .ZN(
        P2_U3188) );
  OAI21_X1 U15201 ( .B1(n12986), .B2(n12985), .A(n12984), .ZN(n12987) );
  NAND2_X1 U15202 ( .A1(n12987), .A2(n14692), .ZN(n12991) );
  NOR2_X1 U15203 ( .A1(n13231), .A2(n13059), .ZN(n12988) );
  AOI21_X1 U15204 ( .B1(n13237), .B2(n14524), .A(n12988), .ZN(n13383) );
  NAND2_X1 U15205 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13177)
         );
  OAI21_X1 U15206 ( .B1(n13091), .B2(n13383), .A(n13177), .ZN(n12989) );
  AOI21_X1 U15207 ( .B1(n13391), .B2(n13093), .A(n12989), .ZN(n12990) );
  OAI211_X1 U15208 ( .C1(n13575), .C2(n13096), .A(n12991), .B(n12990), .ZN(
        P2_U3191) );
  INV_X1 U15209 ( .A(n12992), .ZN(n12993) );
  NOR2_X1 U15210 ( .A1(n13257), .A2(n13390), .ZN(n12994) );
  XOR2_X1 U15211 ( .A(n12995), .B(n12994), .Z(n12996) );
  XNOR2_X1 U15212 ( .A(n13265), .B(n12996), .ZN(n12997) );
  INV_X1 U15213 ( .A(n12998), .ZN(n13268) );
  OAI22_X1 U15214 ( .A1(n13000), .A2(n13059), .B1(n12999), .B2(n13067), .ZN(
        n13263) );
  AOI22_X1 U15215 ( .A1(n14694), .A2(n13263), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13001) );
  OAI21_X1 U15216 ( .B1(n13268), .B2(n14701), .A(n13001), .ZN(n13002) );
  AOI21_X1 U15217 ( .B1(n7062), .B2(n14697), .A(n13002), .ZN(n13003) );
  OAI211_X1 U15218 ( .C1(n13006), .C2(n13005), .A(n13004), .B(n14692), .ZN(
        n13012) );
  INV_X1 U15219 ( .A(n13360), .ZN(n13010) );
  NOR2_X1 U15220 ( .A1(n13243), .A2(n13067), .ZN(n13007) );
  AOI21_X1 U15221 ( .B1(n13237), .B2(n14522), .A(n13007), .ZN(n13496) );
  OAI22_X1 U15222 ( .A1(n13496), .A2(n13091), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13008), .ZN(n13009) );
  AOI21_X1 U15223 ( .B1(n13010), .B2(n13093), .A(n13009), .ZN(n13011) );
  OAI211_X1 U15224 ( .C1(n13567), .C2(n13096), .A(n13012), .B(n13011), .ZN(
        P2_U3195) );
  INV_X1 U15225 ( .A(n13302), .ZN(n13014) );
  OAI22_X1 U15226 ( .A1(n13206), .A2(n13059), .B1(n13253), .B2(n13067), .ZN(
        n13466) );
  AOI22_X1 U15227 ( .A1(n14694), .A2(n13466), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13013) );
  OAI21_X1 U15228 ( .B1(n13014), .B2(n14701), .A(n13013), .ZN(n13019) );
  AOI211_X1 U15229 ( .C1(n13017), .C2(n13016), .A(n13073), .B(n13015), .ZN(
        n13018) );
  AOI211_X1 U15230 ( .C1(n13308), .C2(n14697), .A(n13019), .B(n13018), .ZN(
        n13020) );
  INV_X1 U15231 ( .A(n13020), .ZN(P2_U3197) );
  INV_X1 U15232 ( .A(n13022), .ZN(n13023) );
  AOI21_X1 U15233 ( .B1(n13024), .B2(n13021), .A(n13023), .ZN(n13029) );
  NOR2_X1 U15234 ( .A1(n14701), .A2(n13426), .ZN(n13027) );
  AND2_X1 U15235 ( .A1(n13100), .A2(n14522), .ZN(n13025) );
  AOI21_X1 U15236 ( .B1(n13228), .B2(n14524), .A(n13025), .ZN(n13533) );
  NAND2_X1 U15237 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n14803)
         );
  OAI21_X1 U15238 ( .B1(n13091), .B2(n13533), .A(n14803), .ZN(n13026) );
  AOI211_X1 U15239 ( .C1(n13422), .C2(n14697), .A(n13027), .B(n13026), .ZN(
        n13028) );
  OAI21_X1 U15240 ( .B1(n13029), .B2(n13073), .A(n13028), .ZN(P2_U3198) );
  OAI21_X1 U15241 ( .B1(n13032), .B2(n13031), .A(n13030), .ZN(n13033) );
  NAND2_X1 U15242 ( .A1(n13033), .A2(n14692), .ZN(n13038) );
  AND2_X1 U15243 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n13142) );
  NOR2_X1 U15244 ( .A1(n14701), .A2(n13034), .ZN(n13035) );
  AOI211_X1 U15245 ( .C1(n14694), .C2(n13036), .A(n13142), .B(n13035), .ZN(
        n13037) );
  OAI211_X1 U15246 ( .C1(n13580), .C2(n13096), .A(n13038), .B(n13037), .ZN(
        P2_U3200) );
  OAI21_X1 U15247 ( .B1(n13041), .B2(n13040), .A(n13039), .ZN(n13047) );
  NAND2_X1 U15248 ( .A1(n13313), .A2(n14697), .ZN(n13044) );
  NAND2_X1 U15249 ( .A1(n13245), .A2(n14522), .ZN(n13042) );
  OAI21_X1 U15250 ( .B1(n13250), .B2(n13067), .A(n13042), .ZN(n13316) );
  AOI22_X1 U15251 ( .A1(n14694), .A2(n13316), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13043) );
  OAI211_X1 U15252 ( .C1(n14701), .C2(n13045), .A(n13044), .B(n13043), .ZN(
        n13046) );
  AOI21_X1 U15253 ( .B1(n13047), .B2(n14692), .A(n13046), .ZN(n13048) );
  INV_X1 U15254 ( .A(n13048), .ZN(P2_U3201) );
  NAND2_X1 U15255 ( .A1(n13050), .A2(n13049), .ZN(n13052) );
  XOR2_X1 U15256 ( .A(n13052), .B(n13051), .Z(n13056) );
  OAI22_X1 U15257 ( .A1(n13239), .A2(n13067), .B1(n13233), .B2(n13059), .ZN(
        n13374) );
  AOI22_X1 U15258 ( .A1(n13374), .A2(n14694), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13053) );
  OAI21_X1 U15259 ( .B1(n13375), .B2(n14701), .A(n13053), .ZN(n13054) );
  AOI21_X1 U15260 ( .B1(n13370), .B2(n14697), .A(n13054), .ZN(n13055) );
  OAI21_X1 U15261 ( .B1(n13056), .B2(n13073), .A(n13055), .ZN(P2_U3205) );
  XOR2_X1 U15262 ( .A(n13058), .B(n13057), .Z(n13064) );
  OAI22_X1 U15263 ( .A1(n13239), .A2(n13059), .B1(n13204), .B2(n13067), .ZN(
        n13342) );
  AOI22_X1 U15264 ( .A1(n13342), .A2(n14694), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13060) );
  OAI21_X1 U15265 ( .B1(n13061), .B2(n14701), .A(n13060), .ZN(n13062) );
  AOI21_X1 U15266 ( .B1(n13491), .B2(n14697), .A(n13062), .ZN(n13063) );
  OAI21_X1 U15267 ( .B1(n13064), .B2(n13073), .A(n13063), .ZN(P2_U3207) );
  XNOR2_X1 U15268 ( .A(n13066), .B(n13065), .ZN(n13074) );
  OR2_X1 U15269 ( .A1(n13233), .A2(n13067), .ZN(n13069) );
  NAND2_X1 U15270 ( .A1(n13228), .A2(n14522), .ZN(n13068) );
  NAND2_X1 U15271 ( .A1(n13069), .A2(n13068), .ZN(n13403) );
  NAND2_X1 U15272 ( .A1(n13403), .A2(n14694), .ZN(n13070) );
  NAND2_X1 U15273 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13158)
         );
  OAI211_X1 U15274 ( .C1(n14701), .C2(n13408), .A(n13070), .B(n13158), .ZN(
        n13071) );
  AOI21_X1 U15275 ( .B1(n13416), .B2(n14697), .A(n13071), .ZN(n13072) );
  OAI21_X1 U15276 ( .B1(n13074), .B2(n13073), .A(n13072), .ZN(P2_U3210) );
  AOI22_X1 U15277 ( .A1(n14694), .A2(n13077), .B1(P2_REG3_REG_6__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13082) );
  NAND2_X1 U15278 ( .A1(n13093), .A2(n13078), .ZN(n13081) );
  NAND2_X1 U15279 ( .A1(n14697), .A2(n13079), .ZN(n13080) );
  NAND4_X1 U15280 ( .A1(n13083), .A2(n13082), .A3(n13081), .A4(n13080), .ZN(
        P2_U3211) );
  OAI21_X1 U15281 ( .B1(n13086), .B2(n13085), .A(n13084), .ZN(n13087) );
  NAND2_X1 U15282 ( .A1(n13087), .A2(n14692), .ZN(n13095) );
  INV_X1 U15283 ( .A(n13250), .ZN(n13208) );
  NAND2_X1 U15284 ( .A1(n13208), .A2(n14522), .ZN(n13089) );
  NAND2_X1 U15285 ( .A1(n13256), .A2(n14524), .ZN(n13088) );
  AND2_X1 U15286 ( .A1(n13089), .A2(n13088), .ZN(n13459) );
  OAI22_X1 U15287 ( .A1(n13091), .A2(n13459), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13090), .ZN(n13092) );
  AOI21_X1 U15288 ( .B1(n13293), .B2(n13093), .A(n13092), .ZN(n13094) );
  OAI211_X1 U15289 ( .C1(n13460), .C2(n13096), .A(n13095), .B(n13094), .ZN(
        P2_U3212) );
  MUX2_X1 U15290 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n13097), .S(n6394), .Z(
        P2_U3562) );
  MUX2_X1 U15291 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13215), .S(n6394), .Z(
        P2_U3561) );
  MUX2_X1 U15292 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13098), .S(n6394), .Z(
        P2_U3560) );
  MUX2_X1 U15293 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13217), .S(n6394), .Z(
        P2_U3559) );
  MUX2_X1 U15294 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13256), .S(n6394), .Z(
        P2_U3558) );
  MUX2_X1 U15295 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13252), .S(n6394), .Z(
        P2_U3557) );
  MUX2_X1 U15296 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13208), .S(n6394), .Z(
        P2_U3556) );
  MUX2_X1 U15297 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13247), .S(P2_U3947), .Z(
        P2_U3555) );
  MUX2_X1 U15298 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13245), .S(P2_U3947), .Z(
        P2_U3554) );
  MUX2_X1 U15299 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13202), .S(n6394), .Z(
        P2_U3553) );
  INV_X1 U15300 ( .A(n13239), .ZN(n13199) );
  MUX2_X1 U15301 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13199), .S(n6394), .Z(
        P2_U3552) );
  MUX2_X1 U15302 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13237), .S(n6394), .Z(
        P2_U3551) );
  MUX2_X1 U15303 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13193), .S(n6394), .Z(
        P2_U3550) );
  MUX2_X1 U15304 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13190), .S(n6394), .Z(
        P2_U3549) );
  MUX2_X1 U15305 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13228), .S(n6394), .Z(
        P2_U3548) );
  MUX2_X1 U15306 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n13099), .S(n6394), .Z(
        P2_U3547) );
  MUX2_X1 U15307 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13100), .S(n6394), .Z(
        P2_U3546) );
  MUX2_X1 U15308 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13101), .S(n6394), .Z(
        P2_U3545) );
  MUX2_X1 U15309 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n14525), .S(n6394), .Z(
        P2_U3544) );
  MUX2_X1 U15310 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13102), .S(n6394), .Z(
        P2_U3543) );
  MUX2_X1 U15311 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n14523), .S(n6394), .Z(
        P2_U3542) );
  MUX2_X1 U15312 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13103), .S(n6394), .Z(
        P2_U3541) );
  MUX2_X1 U15313 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n13104), .S(n6394), .Z(
        P2_U3540) );
  MUX2_X1 U15314 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n13105), .S(n6394), .Z(
        P2_U3539) );
  MUX2_X1 U15315 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n13106), .S(n6394), .Z(
        P2_U3538) );
  MUX2_X1 U15316 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n13107), .S(n6394), .Z(
        P2_U3537) );
  MUX2_X1 U15317 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n13108), .S(n6394), .Z(
        P2_U3536) );
  MUX2_X1 U15318 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n13109), .S(n6394), .Z(
        P2_U3535) );
  MUX2_X1 U15319 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n13110), .S(n6394), .Z(
        P2_U3534) );
  MUX2_X1 U15320 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n13111), .S(n6394), .Z(
        P2_U3533) );
  MUX2_X1 U15321 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n8312), .S(n6394), .Z(
        P2_U3532) );
  MUX2_X1 U15322 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8313), .S(n6394), .Z(
        P2_U3531) );
  OAI211_X1 U15323 ( .C1(n13114), .C2(n13113), .A(n14765), .B(n13112), .ZN(
        n13123) );
  AND2_X1 U15324 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3088), .ZN(n13115) );
  AOI21_X1 U15325 ( .B1(n14719), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n13115), .ZN(
        n13122) );
  NAND2_X1 U15326 ( .A1(n14802), .A2(n13116), .ZN(n13121) );
  OAI211_X1 U15327 ( .C1(n13119), .C2(n13118), .A(n14770), .B(n13117), .ZN(
        n13120) );
  NAND4_X1 U15328 ( .A1(n13123), .A2(n13122), .A3(n13121), .A4(n13120), .ZN(
        P2_U3217) );
  NOR2_X1 U15329 ( .A1(n13125), .A2(n13124), .ZN(n13127) );
  NOR2_X1 U15330 ( .A1(n13128), .A2(n14779), .ZN(n13129) );
  INV_X1 U15331 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n14784) );
  XNOR2_X1 U15332 ( .A(n13128), .B(n14779), .ZN(n14785) );
  NOR2_X1 U15333 ( .A1(n14784), .A2(n14785), .ZN(n14783) );
  XNOR2_X1 U15334 ( .A(n14801), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n14797) );
  NOR2_X1 U15335 ( .A1(n14798), .A2(n14797), .ZN(n14796) );
  AOI21_X1 U15336 ( .B1(n14801), .B2(P2_REG2_REG_16__SCAN_IN), .A(n14796), 
        .ZN(n13133) );
  INV_X1 U15337 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13131) );
  NOR2_X1 U15338 ( .A1(n13148), .A2(n13131), .ZN(n13130) );
  AOI21_X1 U15339 ( .B1(n13148), .B2(n13131), .A(n13130), .ZN(n13132) );
  NOR2_X1 U15340 ( .A1(n13133), .A2(n13132), .ZN(n13146) );
  AOI211_X1 U15341 ( .C1(n13133), .C2(n13132), .A(n13146), .B(n14795), .ZN(
        n13141) );
  NOR2_X1 U15342 ( .A1(n13136), .A2(n14779), .ZN(n13137) );
  INV_X1 U15343 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n14781) );
  XNOR2_X1 U15344 ( .A(n14801), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n14793) );
  XNOR2_X1 U15345 ( .A(n13148), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n13138) );
  AOI211_X1 U15346 ( .C1(n13139), .C2(n13138), .A(n13149), .B(n14791), .ZN(
        n13140) );
  NOR2_X1 U15347 ( .A1(n13141), .A2(n13140), .ZN(n13144) );
  AOI21_X1 U15348 ( .B1(n14719), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n13142), 
        .ZN(n13143) );
  OAI211_X1 U15349 ( .C1(n13145), .C2(n14774), .A(n13144), .B(n13143), .ZN(
        P2_U3231) );
  XNOR2_X1 U15350 ( .A(n13163), .B(n13152), .ZN(n13147) );
  NAND2_X1 U15351 ( .A1(n13147), .A2(n13409), .ZN(n13165) );
  OAI21_X1 U15352 ( .B1(n13409), .B2(n13147), .A(n13165), .ZN(n13157) );
  INV_X1 U15353 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n13155) );
  NAND2_X1 U15354 ( .A1(n13148), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n13151) );
  NAND2_X1 U15355 ( .A1(n13151), .A2(n13150), .ZN(n13153) );
  AOI211_X1 U15356 ( .C1(n13155), .C2(n13154), .A(n13167), .B(n14791), .ZN(
        n13156) );
  AOI21_X1 U15357 ( .B1(n14770), .B2(n13157), .A(n13156), .ZN(n13161) );
  INV_X1 U15358 ( .A(n13158), .ZN(n13159) );
  AOI21_X1 U15359 ( .B1(n14719), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n13159), 
        .ZN(n13160) );
  OAI211_X1 U15360 ( .C1(n13162), .C2(n14774), .A(n13161), .B(n13160), .ZN(
        P2_U3232) );
  NAND2_X1 U15361 ( .A1(n13163), .A2(n13162), .ZN(n13164) );
  NAND2_X1 U15362 ( .A1(n13165), .A2(n13164), .ZN(n13166) );
  XNOR2_X1 U15363 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n13166), .ZN(n13173) );
  INV_X1 U15364 ( .A(n13173), .ZN(n13171) );
  XOR2_X1 U15365 ( .A(n13169), .B(n13168), .Z(n13172) );
  OAI21_X1 U15366 ( .B1(n13172), .B2(n14791), .A(n14774), .ZN(n13170) );
  AOI21_X1 U15367 ( .B1(n13171), .B2(n14770), .A(n13170), .ZN(n13176) );
  AOI22_X1 U15368 ( .A1(n13173), .A2(n14770), .B1(n14765), .B2(n13172), .ZN(
        n13175) );
  OAI211_X1 U15369 ( .C1(n14444), .C2(n14805), .A(n13178), .B(n13177), .ZN(
        P2_U3233) );
  OAI211_X1 U15370 ( .C1(n13221), .C2(n13545), .A(n13390), .B(n13179), .ZN(
        n13442) );
  NOR2_X1 U15371 ( .A1(n13545), .A2(n14812), .ZN(n13180) );
  AOI211_X1 U15372 ( .C1(n6388), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13181), .B(
        n13180), .ZN(n13182) );
  OAI21_X1 U15373 ( .B1(n13413), .B2(n13442), .A(n13182), .ZN(P2_U3235) );
  OR2_X1 U15374 ( .A1(n13229), .A2(n13186), .ZN(n13184) );
  NAND2_X1 U15375 ( .A1(n13229), .A2(n13186), .ZN(n13187) );
  NAND2_X1 U15376 ( .A1(n13188), .A2(n13187), .ZN(n13401) );
  NAND2_X1 U15377 ( .A1(n13520), .A2(n13190), .ZN(n13189) );
  OR2_X1 U15378 ( .A1(n13520), .A2(n13190), .ZN(n13191) );
  NAND2_X1 U15379 ( .A1(n13575), .A2(n13193), .ZN(n13192) );
  OR2_X1 U15380 ( .A1(n13575), .A2(n13193), .ZN(n13194) );
  INV_X1 U15381 ( .A(n13368), .ZN(n13195) );
  NAND2_X1 U15382 ( .A1(n13367), .A2(n13195), .ZN(n13198) );
  NAND2_X1 U15383 ( .A1(n13370), .A2(n13196), .ZN(n13197) );
  NOR2_X1 U15384 ( .A1(n13567), .A2(n13199), .ZN(n13201) );
  NAND2_X1 U15385 ( .A1(n13567), .A2(n13199), .ZN(n13200) );
  INV_X1 U15386 ( .A(n13351), .ZN(n13242) );
  NAND2_X1 U15387 ( .A1(n13348), .A2(n13202), .ZN(n13203) );
  NAND2_X1 U15388 ( .A1(n13336), .A2(n13204), .ZN(n13205) );
  AND2_X1 U15389 ( .A1(n13313), .A2(n13206), .ZN(n13207) );
  OR2_X1 U15390 ( .A1(n13555), .A2(n13208), .ZN(n13209) );
  NAND2_X1 U15391 ( .A1(n13210), .A2(n13209), .ZN(n13290) );
  OR2_X1 U15392 ( .A1(n13550), .A2(n13256), .ZN(n13262) );
  AOI22_X1 U15393 ( .A1(n13217), .A2(n14522), .B1(n13216), .B2(n13215), .ZN(
        n13218) );
  INV_X1 U15394 ( .A(n13218), .ZN(n13219) );
  AOI21_X2 U15395 ( .B1(n13220), .B2(n14520), .A(n13219), .ZN(n13448) );
  INV_X1 U15396 ( .A(n13267), .ZN(n13222) );
  AOI211_X1 U15397 ( .C1(n13446), .C2(n13222), .A(n10035), .B(n13221), .ZN(
        n13445) );
  AOI22_X1 U15398 ( .A1(n14819), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n13223), 
        .B2(n14808), .ZN(n13224) );
  OAI21_X1 U15399 ( .B1(n13225), .B2(n14812), .A(n13224), .ZN(n13259) );
  NAND2_X1 U15400 ( .A1(n13229), .A2(n13228), .ZN(n13230) );
  OR2_X1 U15401 ( .A1(n13575), .A2(n13233), .ZN(n13232) );
  NAND2_X1 U15402 ( .A1(n13575), .A2(n13233), .ZN(n13234) );
  NOR2_X1 U15403 ( .A1(n13370), .A2(n13237), .ZN(n13236) );
  NAND2_X1 U15404 ( .A1(n13370), .A2(n13237), .ZN(n13238) );
  INV_X1 U15405 ( .A(n13355), .ZN(n13357) );
  NAND2_X1 U15406 ( .A1(n13567), .A2(n13239), .ZN(n13240) );
  OR2_X1 U15407 ( .A1(n13348), .A2(n13243), .ZN(n13244) );
  AND2_X1 U15408 ( .A1(n13336), .A2(n13245), .ZN(n13246) );
  NAND2_X1 U15409 ( .A1(n13313), .A2(n13247), .ZN(n13248) );
  NAND2_X1 U15410 ( .A1(n13555), .A2(n13250), .ZN(n13251) );
  NOR2_X1 U15411 ( .A1(n13292), .A2(n13252), .ZN(n13254) );
  XNOR2_X1 U15412 ( .A(n13261), .B(n13260), .ZN(n13454) );
  INV_X1 U15413 ( .A(n13263), .ZN(n13264) );
  NOR2_X1 U15414 ( .A1(n13265), .A2(n13281), .ZN(n13266) );
  OR3_X2 U15415 ( .A1(n13267), .A2(n13266), .A3(n10035), .ZN(n13450) );
  OAI22_X1 U15416 ( .A1(n13450), .A2(n8286), .B1(n13407), .B2(n13268), .ZN(
        n13269) );
  OAI21_X1 U15417 ( .B1(n13451), .B2(n13269), .A(n13438), .ZN(n13271) );
  AOI22_X1 U15418 ( .A1(n7062), .A2(n14531), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n6388), .ZN(n13270) );
  OAI211_X1 U15419 ( .C1(n13434), .C2(n13454), .A(n13271), .B(n13270), .ZN(
        P2_U3237) );
  XNOR2_X1 U15420 ( .A(n13272), .B(n13274), .ZN(n13455) );
  NAND2_X1 U15421 ( .A1(n13274), .A2(n13273), .ZN(n13275) );
  NAND2_X1 U15422 ( .A1(n13276), .A2(n13275), .ZN(n13279) );
  INV_X1 U15423 ( .A(n13277), .ZN(n13278) );
  INV_X1 U15424 ( .A(n13457), .ZN(n13286) );
  NOR2_X1 U15425 ( .A1(n13550), .A2(n13291), .ZN(n13280) );
  NOR2_X1 U15426 ( .A1(n13456), .A2(n13413), .ZN(n13285) );
  AOI22_X1 U15427 ( .A1(n14819), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n13282), 
        .B2(n14808), .ZN(n13283) );
  OAI21_X1 U15428 ( .B1(n13550), .B2(n14812), .A(n13283), .ZN(n13284) );
  AOI211_X1 U15429 ( .C1(n13286), .C2(n13438), .A(n13285), .B(n13284), .ZN(
        n13287) );
  OAI21_X1 U15430 ( .B1(n13455), .B2(n13434), .A(n13287), .ZN(P2_U3238) );
  XNOR2_X1 U15431 ( .A(n13288), .B(n13289), .ZN(n13465) );
  XNOR2_X1 U15432 ( .A(n13290), .B(n13289), .ZN(n13463) );
  AOI211_X1 U15433 ( .C1(n13292), .C2(n13305), .A(n10035), .B(n13291), .ZN(
        n13461) );
  NAND2_X1 U15434 ( .A1(n13461), .A2(n14806), .ZN(n13297) );
  INV_X1 U15435 ( .A(n13293), .ZN(n13294) );
  OAI22_X1 U15436 ( .A1(n14819), .A2(n13459), .B1(n13294), .B2(n13407), .ZN(
        n13295) );
  AOI21_X1 U15437 ( .B1(P2_REG2_REG_26__SCAN_IN), .B2(n6388), .A(n13295), .ZN(
        n13296) );
  OAI211_X1 U15438 ( .C1(n13460), .C2(n14812), .A(n13297), .B(n13296), .ZN(
        n13298) );
  AOI21_X1 U15439 ( .B1(n13463), .B2(n13299), .A(n13298), .ZN(n13300) );
  OAI21_X1 U15440 ( .B1(n13465), .B2(n13434), .A(n13300), .ZN(P2_U3239) );
  XNOR2_X1 U15441 ( .A(n7084), .B(n13301), .ZN(n13469) );
  INV_X1 U15442 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n13304) );
  AOI22_X1 U15443 ( .A1(n13438), .A2(n13466), .B1(n13302), .B2(n14808), .ZN(
        n13303) );
  OAI21_X1 U15444 ( .B1(n13304), .B2(n13438), .A(n13303), .ZN(n13307) );
  OAI211_X1 U15445 ( .C1(n13315), .C2(n13555), .A(n13390), .B(n13305), .ZN(
        n13467) );
  NOR2_X1 U15446 ( .A1(n13467), .A2(n13413), .ZN(n13306) );
  AOI211_X1 U15447 ( .C1(n14531), .C2(n13308), .A(n13307), .B(n13306), .ZN(
        n13311) );
  XNOR2_X1 U15448 ( .A(n13309), .B(n7084), .ZN(n13471) );
  NAND2_X1 U15449 ( .A1(n13471), .A2(n14815), .ZN(n13310) );
  OAI211_X1 U15450 ( .C1(n13469), .C2(n13440), .A(n13311), .B(n13310), .ZN(
        P2_U3240) );
  XNOR2_X1 U15451 ( .A(n13321), .B(n13312), .ZN(n13474) );
  INV_X1 U15452 ( .A(n13474), .ZN(n13325) );
  AND2_X1 U15453 ( .A1(n13313), .A2(n13334), .ZN(n13314) );
  OR3_X1 U15454 ( .A1(n13315), .A2(n13314), .A3(n10035), .ZN(n13476) );
  INV_X1 U15455 ( .A(n13316), .ZN(n13475) );
  OAI21_X1 U15456 ( .B1(n13476), .B2(n8286), .A(n13475), .ZN(n13320) );
  AOI22_X1 U15457 ( .A1(n6388), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n13317), 
        .B2(n14808), .ZN(n13318) );
  OAI21_X1 U15458 ( .B1(n13559), .B2(n14812), .A(n13318), .ZN(n13319) );
  AOI21_X1 U15459 ( .B1(n13320), .B2(n13438), .A(n13319), .ZN(n13324) );
  NAND2_X1 U15460 ( .A1(n13322), .A2(n13321), .ZN(n13477) );
  NAND3_X1 U15461 ( .A1(n13478), .A2(n13477), .A3(n14815), .ZN(n13323) );
  OAI211_X1 U15462 ( .C1(n13325), .C2(n13440), .A(n13324), .B(n13323), .ZN(
        P2_U3241) );
  XNOR2_X1 U15463 ( .A(n13326), .B(n13332), .ZN(n13327) );
  INV_X1 U15464 ( .A(n13486), .ZN(n13330) );
  AOI21_X1 U15465 ( .B1(n13331), .B2(n14808), .A(n13330), .ZN(n13340) );
  XNOR2_X1 U15466 ( .A(n13333), .B(n13332), .ZN(n13484) );
  AOI21_X1 U15467 ( .B1(n13336), .B2(n13344), .A(n10035), .ZN(n13335) );
  NAND2_X1 U15468 ( .A1(n13335), .A2(n13334), .ZN(n13485) );
  AOI22_X1 U15469 ( .A1(n13336), .A2(n14531), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(n14819), .ZN(n13337) );
  OAI21_X1 U15470 ( .B1(n13485), .B2(n13413), .A(n13337), .ZN(n13338) );
  AOI21_X1 U15471 ( .B1(n13484), .B2(n14815), .A(n13338), .ZN(n13339) );
  OAI21_X1 U15472 ( .B1(n13340), .B2(n6388), .A(n13339), .ZN(P2_U3242) );
  XNOR2_X1 U15473 ( .A(n13341), .B(n13351), .ZN(n13343) );
  AOI21_X1 U15474 ( .B1(n13343), .B2(n14520), .A(n13342), .ZN(n13493) );
  AOI21_X1 U15475 ( .B1(n13491), .B2(n13359), .A(n10035), .ZN(n13345) );
  AND2_X1 U15476 ( .A1(n13345), .A2(n13344), .ZN(n13490) );
  AOI22_X1 U15477 ( .A1(n14819), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n13346), 
        .B2(n14808), .ZN(n13347) );
  OAI21_X1 U15478 ( .B1(n13348), .B2(n14812), .A(n13347), .ZN(n13353) );
  OAI21_X1 U15479 ( .B1(n7277), .B2(n13351), .A(n13350), .ZN(n13494) );
  NOR2_X1 U15480 ( .A1(n13494), .A2(n13434), .ZN(n13352) );
  AOI211_X1 U15481 ( .C1(n13490), .C2(n14806), .A(n13353), .B(n13352), .ZN(
        n13354) );
  OAI21_X1 U15482 ( .B1(n6388), .B2(n13493), .A(n13354), .ZN(P2_U3243) );
  XNOR2_X1 U15483 ( .A(n13356), .B(n13355), .ZN(n13500) );
  XNOR2_X1 U15484 ( .A(n13358), .B(n13357), .ZN(n13495) );
  OAI211_X1 U15485 ( .C1(n13371), .C2(n13567), .A(n13390), .B(n13359), .ZN(
        n13497) );
  NOR2_X1 U15486 ( .A1(n13497), .A2(n13413), .ZN(n13365) );
  OAI22_X1 U15487 ( .A1(n13496), .A2(n14819), .B1(n13360), .B2(n13407), .ZN(
        n13361) );
  INV_X1 U15488 ( .A(n13361), .ZN(n13363) );
  NAND2_X1 U15489 ( .A1(n14819), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n13362) );
  OAI211_X1 U15490 ( .C1(n13567), .C2(n14812), .A(n13363), .B(n13362), .ZN(
        n13364) );
  AOI211_X1 U15491 ( .C1(n13495), .C2(n14815), .A(n13365), .B(n13364), .ZN(
        n13366) );
  OAI21_X1 U15492 ( .B1(n13500), .B2(n13440), .A(n13366), .ZN(P2_U3244) );
  XNOR2_X1 U15493 ( .A(n13367), .B(n13368), .ZN(n13505) );
  XNOR2_X1 U15494 ( .A(n13369), .B(n13368), .ZN(n13507) );
  NAND2_X1 U15495 ( .A1(n13507), .A2(n14815), .ZN(n13381) );
  INV_X1 U15496 ( .A(n13389), .ZN(n13373) );
  INV_X1 U15497 ( .A(n13371), .ZN(n13372) );
  OAI211_X1 U15498 ( .C1(n13571), .C2(n13373), .A(n13372), .B(n13390), .ZN(
        n13503) );
  INV_X1 U15499 ( .A(n13503), .ZN(n13379) );
  INV_X1 U15500 ( .A(n13374), .ZN(n13504) );
  OAI22_X1 U15501 ( .A1(n13504), .A2(n14819), .B1(n13375), .B2(n13407), .ZN(
        n13376) );
  AOI21_X1 U15502 ( .B1(P2_REG2_REG_20__SCAN_IN), .B2(n6388), .A(n13376), .ZN(
        n13377) );
  OAI21_X1 U15503 ( .B1(n13571), .B2(n14812), .A(n13377), .ZN(n13378) );
  AOI21_X1 U15504 ( .B1(n13379), .B2(n14806), .A(n13378), .ZN(n13380) );
  OAI211_X1 U15505 ( .C1(n13505), .C2(n13440), .A(n13381), .B(n13380), .ZN(
        P2_U3245) );
  XNOR2_X1 U15506 ( .A(n13382), .B(n13386), .ZN(n13385) );
  INV_X1 U15507 ( .A(n13383), .ZN(n13384) );
  AOI21_X1 U15508 ( .B1(n13385), .B2(n14520), .A(n13384), .ZN(n13512) );
  INV_X1 U15509 ( .A(n13386), .ZN(n13387) );
  XNOR2_X1 U15510 ( .A(n13388), .B(n13387), .ZN(n13510) );
  OAI211_X1 U15511 ( .C1(n13411), .C2(n13575), .A(n13390), .B(n13389), .ZN(
        n13511) );
  NOR2_X1 U15512 ( .A1(n13511), .A2(n13413), .ZN(n13394) );
  AOI22_X1 U15513 ( .A1(n14819), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13391), 
        .B2(n14808), .ZN(n13392) );
  OAI21_X1 U15514 ( .B1(n13575), .B2(n14812), .A(n13392), .ZN(n13393) );
  AOI211_X1 U15515 ( .C1(n13510), .C2(n14815), .A(n13394), .B(n13393), .ZN(
        n13395) );
  OAI21_X1 U15516 ( .B1(n6388), .B2(n13512), .A(n13395), .ZN(P2_U3246) );
  NAND2_X1 U15517 ( .A1(n13396), .A2(n13399), .ZN(n13397) );
  NAND2_X1 U15518 ( .A1(n13398), .A2(n13397), .ZN(n13517) );
  INV_X1 U15519 ( .A(n13517), .ZN(n13420) );
  INV_X1 U15520 ( .A(n13399), .ZN(n13400) );
  XNOR2_X1 U15521 ( .A(n13401), .B(n13400), .ZN(n13406) );
  NAND2_X1 U15522 ( .A1(n13517), .A2(n13402), .ZN(n13405) );
  INV_X1 U15523 ( .A(n13403), .ZN(n13404) );
  OAI211_X1 U15524 ( .C1(n13538), .C2(n13406), .A(n13405), .B(n13404), .ZN(
        n13522) );
  NAND2_X1 U15525 ( .A1(n13522), .A2(n13438), .ZN(n13418) );
  OAI22_X1 U15526 ( .A1(n13438), .A2(n13409), .B1(n13408), .B2(n13407), .ZN(
        n13415) );
  NOR2_X1 U15527 ( .A1(n13410), .A2(n13520), .ZN(n13412) );
  NOR2_X1 U15528 ( .A1(n13518), .A2(n13413), .ZN(n13414) );
  AOI211_X1 U15529 ( .C1(n14531), .C2(n13416), .A(n13415), .B(n13414), .ZN(
        n13417) );
  OAI211_X1 U15530 ( .C1(n13420), .C2(n13419), .A(n13418), .B(n13417), .ZN(
        P2_U3247) );
  XNOR2_X1 U15531 ( .A(n13421), .B(n13430), .ZN(n13537) );
  AOI21_X1 U15532 ( .B1(n13423), .B2(n13422), .A(n10035), .ZN(n13425) );
  NAND2_X1 U15533 ( .A1(n13425), .A2(n13424), .ZN(n13534) );
  INV_X1 U15534 ( .A(n13426), .ZN(n13427) );
  NAND2_X1 U15535 ( .A1(n14808), .A2(n13427), .ZN(n13428) );
  OAI211_X1 U15536 ( .C1(n13534), .C2(n8286), .A(n13533), .B(n13428), .ZN(
        n13437) );
  INV_X1 U15537 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13429) );
  OAI22_X1 U15538 ( .A1(n13585), .A2(n14812), .B1(n13429), .B2(n13438), .ZN(
        n13436) );
  NAND2_X1 U15539 ( .A1(n13431), .A2(n13430), .ZN(n13432) );
  NAND2_X1 U15540 ( .A1(n13433), .A2(n13432), .ZN(n13532) );
  NOR2_X1 U15541 ( .A1(n13532), .A2(n13434), .ZN(n13435) );
  AOI211_X1 U15542 ( .C1(n13438), .C2(n13437), .A(n13436), .B(n13435), .ZN(
        n13439) );
  OAI21_X1 U15543 ( .B1(n13440), .B2(n13537), .A(n13439), .ZN(P2_U3249) );
  INV_X1 U15544 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n13443) );
  AND2_X1 U15545 ( .A1(n13442), .A2(n13441), .ZN(n13542) );
  MUX2_X1 U15546 ( .A(n13443), .B(n13542), .S(n14852), .Z(n13444) );
  OAI21_X1 U15547 ( .B1(n13545), .B2(n13541), .A(n13444), .ZN(P2_U3529) );
  AOI21_X1 U15548 ( .B1(n14830), .B2(n13446), .A(n13445), .ZN(n13447) );
  MUX2_X1 U15549 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13546), .S(n14852), .Z(
        P2_U3528) );
  INV_X1 U15550 ( .A(n13450), .ZN(n13452) );
  MUX2_X1 U15551 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13547), .S(n14852), .Z(
        P2_U3527) );
  OAI21_X1 U15552 ( .B1(n13460), .B2(n14841), .A(n13459), .ZN(n13462) );
  AOI211_X1 U15553 ( .C1(n13463), .C2(n14520), .A(n13462), .B(n13461), .ZN(
        n13464) );
  OAI21_X1 U15554 ( .B1(n13531), .B2(n13465), .A(n13464), .ZN(n13551) );
  MUX2_X1 U15555 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13551), .S(n14852), .Z(
        P2_U3525) );
  INV_X1 U15556 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n13472) );
  INV_X1 U15557 ( .A(n13466), .ZN(n13468) );
  OAI211_X1 U15558 ( .C1(n13469), .C2(n13538), .A(n13468), .B(n13467), .ZN(
        n13470) );
  AOI21_X1 U15559 ( .B1(n14845), .B2(n13471), .A(n13470), .ZN(n13552) );
  MUX2_X1 U15560 ( .A(n13472), .B(n13552), .S(n14852), .Z(n13473) );
  OAI21_X1 U15561 ( .B1(n13555), .B2(n13541), .A(n13473), .ZN(P2_U3524) );
  NAND2_X1 U15562 ( .A1(n13474), .A2(n14520), .ZN(n13481) );
  AND2_X1 U15563 ( .A1(n13476), .A2(n13475), .ZN(n13480) );
  NAND3_X1 U15564 ( .A1(n13478), .A2(n13477), .A3(n14845), .ZN(n13479) );
  NAND3_X1 U15565 ( .A1(n13481), .A2(n13480), .A3(n13479), .ZN(n13556) );
  MUX2_X1 U15566 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13556), .S(n14852), .Z(
        n13482) );
  INV_X1 U15567 ( .A(n13482), .ZN(n13483) );
  OAI21_X1 U15568 ( .B1(n13559), .B2(n13541), .A(n13483), .ZN(P2_U3523) );
  NAND2_X1 U15569 ( .A1(n13484), .A2(n14845), .ZN(n13487) );
  NAND3_X1 U15570 ( .A1(n13487), .A2(n13486), .A3(n13485), .ZN(n13560) );
  MUX2_X1 U15571 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13560), .S(n14852), .Z(
        n13488) );
  INV_X1 U15572 ( .A(n13488), .ZN(n13489) );
  OAI21_X1 U15573 ( .B1(n7069), .B2(n13541), .A(n13489), .ZN(P2_U3522) );
  AOI21_X1 U15574 ( .B1(n14830), .B2(n13491), .A(n13490), .ZN(n13492) );
  OAI211_X1 U15575 ( .C1(n13494), .C2(n13531), .A(n13493), .B(n13492), .ZN(
        n13563) );
  MUX2_X1 U15576 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13563), .S(n14852), .Z(
        P2_U3521) );
  NAND2_X1 U15577 ( .A1(n13495), .A2(n14845), .ZN(n13499) );
  AND2_X1 U15578 ( .A1(n13497), .A2(n13496), .ZN(n13498) );
  OAI211_X1 U15579 ( .C1(n13538), .C2(n13500), .A(n13499), .B(n13498), .ZN(
        n13564) );
  MUX2_X1 U15580 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13564), .S(n14852), .Z(
        n13501) );
  INV_X1 U15581 ( .A(n13501), .ZN(n13502) );
  OAI21_X1 U15582 ( .B1(n13567), .B2(n13541), .A(n13502), .ZN(P2_U3520) );
  OAI211_X1 U15583 ( .C1(n13505), .C2(n13538), .A(n13504), .B(n13503), .ZN(
        n13506) );
  AOI21_X1 U15584 ( .B1(n13507), .B2(n14845), .A(n13506), .ZN(n13568) );
  MUX2_X1 U15585 ( .A(n13508), .B(n13568), .S(n14852), .Z(n13509) );
  OAI21_X1 U15586 ( .B1(n13571), .B2(n13541), .A(n13509), .ZN(P2_U3519) );
  NAND2_X1 U15587 ( .A1(n13510), .A2(n14845), .ZN(n13513) );
  NAND3_X1 U15588 ( .A1(n13513), .A2(n13512), .A3(n13511), .ZN(n13572) );
  MUX2_X1 U15589 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13572), .S(n14852), .Z(
        n13514) );
  INV_X1 U15590 ( .A(n13514), .ZN(n13515) );
  OAI21_X1 U15591 ( .B1(n13575), .B2(n13541), .A(n13515), .ZN(P2_U3518) );
  NAND2_X1 U15592 ( .A1(n13517), .A2(n13516), .ZN(n13519) );
  OAI211_X1 U15593 ( .C1(n13520), .C2(n14841), .A(n13519), .B(n13518), .ZN(
        n13521) );
  OR2_X1 U15594 ( .A1(n13522), .A2(n13521), .ZN(n13576) );
  MUX2_X1 U15595 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13576), .S(n14852), .Z(
        P2_U3517) );
  NAND2_X1 U15596 ( .A1(n13523), .A2(n14845), .ZN(n13527) );
  AND2_X1 U15597 ( .A1(n13525), .A2(n13524), .ZN(n13526) );
  OAI211_X1 U15598 ( .C1(n13538), .C2(n13528), .A(n13527), .B(n13526), .ZN(
        n13577) );
  MUX2_X1 U15599 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13577), .S(n14852), .Z(
        n13529) );
  INV_X1 U15600 ( .A(n13529), .ZN(n13530) );
  OAI21_X1 U15601 ( .B1(n13580), .B2(n13541), .A(n13530), .ZN(P2_U3516) );
  OR2_X1 U15602 ( .A1(n13532), .A2(n13531), .ZN(n13536) );
  AND2_X1 U15603 ( .A1(n13534), .A2(n13533), .ZN(n13535) );
  OAI211_X1 U15604 ( .C1(n13538), .C2(n13537), .A(n13536), .B(n13535), .ZN(
        n13581) );
  MUX2_X1 U15605 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13581), .S(n14852), .Z(
        n13539) );
  INV_X1 U15606 ( .A(n13539), .ZN(n13540) );
  OAI21_X1 U15607 ( .B1(n13585), .B2(n13541), .A(n13540), .ZN(P2_U3515) );
  INV_X1 U15608 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n13543) );
  MUX2_X1 U15609 ( .A(n13543), .B(n13542), .S(n14848), .Z(n13544) );
  OAI21_X1 U15610 ( .B1(n13545), .B2(n13584), .A(n13544), .ZN(P2_U3497) );
  MUX2_X1 U15611 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13547), .S(n14848), .Z(
        P2_U3495) );
  MUX2_X1 U15612 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13551), .S(n14848), .Z(
        P2_U3493) );
  INV_X1 U15613 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n13553) );
  MUX2_X1 U15614 ( .A(n13553), .B(n13552), .S(n14848), .Z(n13554) );
  OAI21_X1 U15615 ( .B1(n13555), .B2(n13584), .A(n13554), .ZN(P2_U3492) );
  MUX2_X1 U15616 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13556), .S(n14848), .Z(
        n13557) );
  INV_X1 U15617 ( .A(n13557), .ZN(n13558) );
  OAI21_X1 U15618 ( .B1(n13559), .B2(n13584), .A(n13558), .ZN(P2_U3491) );
  MUX2_X1 U15619 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13560), .S(n14848), .Z(
        n13561) );
  INV_X1 U15620 ( .A(n13561), .ZN(n13562) );
  OAI21_X1 U15621 ( .B1(n7069), .B2(n13584), .A(n13562), .ZN(P2_U3490) );
  MUX2_X1 U15622 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13563), .S(n14848), .Z(
        P2_U3489) );
  MUX2_X1 U15623 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13564), .S(n14848), .Z(
        n13565) );
  INV_X1 U15624 ( .A(n13565), .ZN(n13566) );
  OAI21_X1 U15625 ( .B1(n13567), .B2(n13584), .A(n13566), .ZN(P2_U3488) );
  INV_X1 U15626 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n13569) );
  MUX2_X1 U15627 ( .A(n13569), .B(n13568), .S(n14848), .Z(n13570) );
  OAI21_X1 U15628 ( .B1(n13571), .B2(n13584), .A(n13570), .ZN(P2_U3487) );
  MUX2_X1 U15629 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13572), .S(n14848), .Z(
        n13573) );
  INV_X1 U15630 ( .A(n13573), .ZN(n13574) );
  OAI21_X1 U15631 ( .B1(n13575), .B2(n13584), .A(n13574), .ZN(P2_U3486) );
  MUX2_X1 U15632 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13576), .S(n14848), .Z(
        P2_U3484) );
  MUX2_X1 U15633 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13577), .S(n14848), .Z(
        n13578) );
  INV_X1 U15634 ( .A(n13578), .ZN(n13579) );
  OAI21_X1 U15635 ( .B1(n13580), .B2(n13584), .A(n13579), .ZN(P2_U3481) );
  MUX2_X1 U15636 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13581), .S(n14848), .Z(
        n13582) );
  INV_X1 U15637 ( .A(n13582), .ZN(n13583) );
  OAI21_X1 U15638 ( .B1(n13585), .B2(n13584), .A(n13583), .ZN(P2_U3478) );
  INV_X1 U15639 ( .A(n13586), .ZN(n13590) );
  INV_X1 U15640 ( .A(n7638), .ZN(n13587) );
  NOR4_X1 U15641 ( .A1(n13587), .A2(P2_IR_REG_30__SCAN_IN), .A3(n7827), .A4(
        P2_U3088), .ZN(n13588) );
  AOI21_X1 U15642 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n13602), .A(n13588), 
        .ZN(n13589) );
  OAI21_X1 U15643 ( .B1(n13590), .B2(n13605), .A(n13589), .ZN(P2_U3296) );
  INV_X1 U15644 ( .A(n13591), .ZN(n14286) );
  OAI222_X1 U15645 ( .A1(n13605), .A2(n14286), .B1(n13593), .B2(P2_U3088), 
        .C1(n13592), .C2(n13614), .ZN(P2_U3298) );
  NAND2_X1 U15646 ( .A1(n13595), .A2(n13594), .ZN(n13597) );
  OAI211_X1 U15647 ( .C1(n13614), .C2(n15244), .A(n13597), .B(n13596), .ZN(
        P2_U3299) );
  INV_X1 U15648 ( .A(n13598), .ZN(n14291) );
  OAI222_X1 U15649 ( .A1(n13605), .A2(n14291), .B1(n13600), .B2(P2_U3088), 
        .C1(n13599), .C2(n13614), .ZN(P2_U3300) );
  INV_X1 U15650 ( .A(n13601), .ZN(n14293) );
  AOI22_X1 U15651 ( .A1(n13603), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n13602), .ZN(n13604) );
  OAI21_X1 U15652 ( .B1(n14293), .B2(n13605), .A(n13604), .ZN(P2_U3301) );
  INV_X1 U15653 ( .A(n13606), .ZN(n14296) );
  OAI222_X1 U15654 ( .A1(n13614), .A2(n13608), .B1(n13605), .B2(n14296), .C1(
        P2_U3088), .C2(n13607), .ZN(P2_U3302) );
  INV_X1 U15655 ( .A(n13609), .ZN(n14299) );
  INV_X1 U15656 ( .A(n13610), .ZN(n13611) );
  OAI222_X1 U15657 ( .A1(n13614), .A2(n13613), .B1(n13605), .B2(n14299), .C1(
        P2_U3088), .C2(n13611), .ZN(P2_U3303) );
  INV_X1 U15658 ( .A(n13615), .ZN(n13616) );
  MUX2_X1 U15659 ( .A(n13616), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  OAI21_X1 U15660 ( .B1(n13619), .B2(n13618), .A(n13617), .ZN(n13620) );
  NAND2_X1 U15661 ( .A1(n13620), .A2(n13757), .ZN(n13624) );
  NOR2_X1 U15662 ( .A1(n13763), .A2(n13965), .ZN(n13622) );
  INV_X1 U15663 ( .A(n13961), .ZN(n13925) );
  OAI22_X1 U15664 ( .A1(n13903), .A2(n13765), .B1(n13766), .B2(n13925), .ZN(
        n13621) );
  AOI211_X1 U15665 ( .C1(P1_REG3_REG_27__SCAN_IN), .C2(P1_U3086), .A(n13622), 
        .B(n13621), .ZN(n13623) );
  OAI211_X1 U15666 ( .C1(n13968), .C2(n13741), .A(n13624), .B(n13623), .ZN(
        P1_U3214) );
  INV_X1 U15667 ( .A(n13625), .ZN(n13626) );
  AOI21_X1 U15668 ( .B1(n13628), .B2(n13627), .A(n13626), .ZN(n13636) );
  NAND2_X1 U15669 ( .A1(n13753), .A2(n13629), .ZN(n13630) );
  OAI211_X1 U15670 ( .C1(n13763), .C2(n13632), .A(n13631), .B(n13630), .ZN(
        n13633) );
  AOI21_X1 U15671 ( .B1(n13634), .B2(n13769), .A(n13633), .ZN(n13635) );
  OAI21_X1 U15672 ( .B1(n13636), .B2(n13771), .A(n13635), .ZN(P1_U3215) );
  OAI21_X1 U15673 ( .B1(n13639), .B2(n13638), .A(n13637), .ZN(n13640) );
  NAND2_X1 U15674 ( .A1(n13640), .A2(n13757), .ZN(n13646) );
  NAND2_X1 U15675 ( .A1(n13775), .A2(n14133), .ZN(n13642) );
  OR2_X1 U15676 ( .A1(n14102), .A2(n13921), .ZN(n13641) );
  NAND2_X1 U15677 ( .A1(n13642), .A2(n13641), .ZN(n14198) );
  INV_X1 U15678 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n13643) );
  OAI22_X1 U15679 ( .A1(n13763), .A2(n14018), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13643), .ZN(n13644) );
  AOI21_X1 U15680 ( .B1(n14198), .B2(n13753), .A(n13644), .ZN(n13645) );
  OAI211_X1 U15681 ( .C1(n14197), .C2(n13741), .A(n13646), .B(n13645), .ZN(
        P1_U3216) );
  INV_X1 U15682 ( .A(n14086), .ZN(n14229) );
  OAI21_X1 U15683 ( .B1(n6433), .B2(n13648), .A(n13647), .ZN(n13649) );
  NAND3_X1 U15684 ( .A1(n6538), .A2(n13757), .A3(n13649), .ZN(n13653) );
  NAND2_X1 U15685 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n15237)
         );
  INV_X1 U15686 ( .A(n15237), .ZN(n13651) );
  OAI22_X1 U15687 ( .A1(n14080), .A2(n13766), .B1(n13765), .B2(n14079), .ZN(
        n13650) );
  AOI211_X1 U15688 ( .C1(n13711), .C2(n14090), .A(n13651), .B(n13650), .ZN(
        n13652) );
  OAI211_X1 U15689 ( .C1(n14229), .C2(n13741), .A(n13653), .B(n13652), .ZN(
        P1_U3219) );
  AOI21_X1 U15690 ( .B1(n13655), .B2(n13654), .A(n6430), .ZN(n13660) );
  OAI22_X1 U15691 ( .A1(n14050), .A2(n13763), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13656), .ZN(n13658) );
  INV_X1 U15692 ( .A(n13775), .ZN(n14043) );
  OAI22_X1 U15693 ( .A1(n14043), .A2(n13766), .B1(n14080), .B2(n13765), .ZN(
        n13657) );
  AOI211_X1 U15694 ( .C1(n14212), .C2(n13769), .A(n13658), .B(n13657), .ZN(
        n13659) );
  OAI21_X1 U15695 ( .B1(n13660), .B2(n13771), .A(n13659), .ZN(P1_U3223) );
  OAI211_X1 U15696 ( .C1(n13664), .C2(n13663), .A(n13662), .B(n13757), .ZN(
        n13672) );
  INV_X1 U15697 ( .A(n13665), .ZN(n13670) );
  OAI22_X1 U15698 ( .A1(n13667), .A2(n13765), .B1(n13766), .B2(n13666), .ZN(
        n13668) );
  AOI211_X1 U15699 ( .C1(n13711), .C2(n13670), .A(n13669), .B(n13668), .ZN(
        n13671) );
  OAI211_X1 U15700 ( .C1(n6823), .C2(n13741), .A(n13672), .B(n13671), .ZN(
        P1_U3224) );
  OAI21_X1 U15701 ( .B1(n13675), .B2(n13674), .A(n13673), .ZN(n13681) );
  NAND2_X1 U15702 ( .A1(n13922), .A2(n13769), .ZN(n13679) );
  OR2_X1 U15703 ( .A1(n14078), .A2(n13921), .ZN(n13677) );
  OR2_X1 U15704 ( .A1(n14102), .A2(n13903), .ZN(n13676) );
  NAND2_X1 U15705 ( .A1(n13677), .A2(n13676), .ZN(n14185) );
  AOI22_X1 U15706 ( .A1(n13753), .A2(n14185), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13678) );
  OAI211_X1 U15707 ( .C1(n13763), .C2(n13989), .A(n13679), .B(n13678), .ZN(
        n13680) );
  AOI21_X1 U15708 ( .B1(n13681), .B2(n13757), .A(n13680), .ZN(n13682) );
  INV_X1 U15709 ( .A(n13682), .ZN(P1_U3225) );
  OAI21_X1 U15710 ( .B1(n13684), .B2(n13683), .A(n13694), .ZN(n13685) );
  NAND2_X1 U15711 ( .A1(n13685), .A2(n13757), .ZN(n13691) );
  INV_X1 U15712 ( .A(n14137), .ZN(n13689) );
  OAI22_X1 U15713 ( .A1(n13686), .A2(n13765), .B1(n13766), .B2(n13892), .ZN(
        n13687) );
  AOI211_X1 U15714 ( .C1(n13711), .C2(n13689), .A(n13688), .B(n13687), .ZN(
        n13690) );
  OAI211_X1 U15715 ( .C1(n7217), .C2(n13741), .A(n13691), .B(n13690), .ZN(
        P1_U3226) );
  AND3_X1 U15716 ( .A1(n13694), .A2(n13693), .A3(n13692), .ZN(n13695) );
  OAI21_X1 U15717 ( .B1(n13696), .B2(n13695), .A(n13757), .ZN(n13702) );
  NAND2_X1 U15718 ( .A1(n13913), .A2(n14135), .ZN(n13698) );
  NAND2_X1 U15719 ( .A1(n13889), .A2(n14133), .ZN(n13697) );
  AND2_X1 U15720 ( .A1(n13698), .A2(n13697), .ZN(n14241) );
  OAI21_X1 U15721 ( .B1(n14241), .B2(n13709), .A(n13699), .ZN(n13700) );
  AOI21_X1 U15722 ( .B1(n14121), .B2(n13711), .A(n13700), .ZN(n13701) );
  OAI211_X1 U15723 ( .C1(n14242), .C2(n13741), .A(n13702), .B(n13701), .ZN(
        P1_U3228) );
  OAI21_X1 U15724 ( .B1(n13705), .B2(n13704), .A(n13703), .ZN(n13706) );
  NAND2_X1 U15725 ( .A1(n13706), .A2(n13757), .ZN(n13713) );
  INV_X1 U15726 ( .A(n13707), .ZN(n14010) );
  AOI22_X1 U15727 ( .A1(n14133), .A2(n14037), .B1(n14135), .B2(n13773), .ZN(
        n14004) );
  INV_X1 U15728 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n13708) );
  OAI22_X1 U15729 ( .A1(n14004), .A2(n13709), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13708), .ZN(n13710) );
  AOI21_X1 U15730 ( .B1(n14010), .B2(n13711), .A(n13710), .ZN(n13712) );
  OAI211_X1 U15731 ( .C1(n14012), .C2(n13741), .A(n13713), .B(n13712), .ZN(
        P1_U3229) );
  XOR2_X1 U15732 ( .A(n13714), .B(n13715), .Z(n13716) );
  NAND2_X1 U15733 ( .A1(n13716), .A2(n13757), .ZN(n13722) );
  INV_X1 U15734 ( .A(n13766), .ZN(n13720) );
  NOR2_X1 U15735 ( .A1(n13765), .A2(n14103), .ZN(n13719) );
  OAI22_X1 U15736 ( .A1(n13763), .A2(n14056), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13717), .ZN(n13718) );
  AOI211_X1 U15737 ( .C1(n13720), .C2(n14062), .A(n13719), .B(n13718), .ZN(
        n13721) );
  OAI211_X1 U15738 ( .C1(n14218), .C2(n13741), .A(n13722), .B(n13721), .ZN(
        P1_U3233) );
  XNOR2_X1 U15739 ( .A(n13724), .B(n13723), .ZN(n13730) );
  NAND2_X1 U15740 ( .A1(n14561), .A2(n13753), .ZN(n13725) );
  OAI211_X1 U15741 ( .C1(n13763), .C2(n13727), .A(n13726), .B(n13725), .ZN(
        n13728) );
  AOI21_X1 U15742 ( .B1(n14562), .B2(n13769), .A(n13728), .ZN(n13729) );
  OAI21_X1 U15743 ( .B1(n13730), .B2(n13771), .A(n13729), .ZN(P1_U3234) );
  INV_X1 U15744 ( .A(n13731), .ZN(n13735) );
  NOR3_X1 U15745 ( .A1(n6430), .A2(n13733), .A3(n13732), .ZN(n13734) );
  OAI21_X1 U15746 ( .B1(n13735), .B2(n13734), .A(n13757), .ZN(n13740) );
  NOR2_X1 U15747 ( .A1(n14030), .A2(n13763), .ZN(n13738) );
  INV_X1 U15748 ( .A(n14062), .ZN(n13736) );
  OAI22_X1 U15749 ( .A1(n13736), .A2(n13765), .B1(n13919), .B2(n13766), .ZN(
        n13737) );
  AOI211_X1 U15750 ( .C1(P1_REG3_REG_22__SCAN_IN), .C2(P1_U3086), .A(n13738), 
        .B(n13737), .ZN(n13739) );
  OAI211_X1 U15751 ( .C1(n13741), .C2(n14033), .A(n13740), .B(n13739), .ZN(
        P1_U3235) );
  AOI21_X1 U15752 ( .B1(n13743), .B2(n13742), .A(n6433), .ZN(n13747) );
  NAND2_X1 U15753 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n13843)
         );
  OAI21_X1 U15754 ( .B1(n13763), .B2(n14107), .A(n13843), .ZN(n13745) );
  OAI22_X1 U15755 ( .A1(n13892), .A2(n13765), .B1(n13766), .B2(n14103), .ZN(
        n13744) );
  AOI211_X1 U15756 ( .C1(n14237), .C2(n13769), .A(n13745), .B(n13744), .ZN(
        n13746) );
  OAI21_X1 U15757 ( .B1(n13747), .B2(n13771), .A(n13746), .ZN(P1_U3238) );
  OAI21_X1 U15758 ( .B1(n13750), .B2(n13749), .A(n13748), .ZN(n13758) );
  NAND2_X1 U15759 ( .A1(n14179), .A2(n13769), .ZN(n13755) );
  OR2_X1 U15760 ( .A1(n14102), .A2(n13924), .ZN(n13752) );
  OR2_X1 U15761 ( .A1(n14078), .A2(n13923), .ZN(n13751) );
  NAND2_X1 U15762 ( .A1(n13752), .A2(n13751), .ZN(n14178) );
  AOI22_X1 U15763 ( .A1(n13753), .A2(n14178), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13754) );
  OAI211_X1 U15764 ( .C1(n13763), .C2(n13978), .A(n13755), .B(n13754), .ZN(
        n13756) );
  AOI21_X1 U15765 ( .B1(n13758), .B2(n13757), .A(n13756), .ZN(n13759) );
  INV_X1 U15766 ( .A(n13759), .ZN(P1_U3240) );
  XNOR2_X1 U15767 ( .A(n13760), .B(n13761), .ZN(n13772) );
  NAND2_X1 U15768 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14605)
         );
  OAI21_X1 U15769 ( .B1(n13763), .B2(n13762), .A(n14605), .ZN(n13768) );
  OAI22_X1 U15770 ( .A1(n13910), .A2(n13766), .B1(n13765), .B2(n13764), .ZN(
        n13767) );
  AOI211_X1 U15771 ( .C1(n13887), .C2(n13769), .A(n13768), .B(n13767), .ZN(
        n13770) );
  OAI21_X1 U15772 ( .B1(n13772), .B2(n13771), .A(n13770), .ZN(P1_U3241) );
  MUX2_X1 U15773 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n13879), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U15774 ( .A(n13933), .B(P1_DATAO_REG_30__SCAN_IN), .S(n13793), .Z(
        P1_U3590) );
  MUX2_X1 U15775 ( .A(n13941), .B(P1_DATAO_REG_29__SCAN_IN), .S(n13793), .Z(
        P1_U3589) );
  MUX2_X1 U15776 ( .A(n13961), .B(P1_DATAO_REG_28__SCAN_IN), .S(n13793), .Z(
        P1_U3588) );
  MUX2_X1 U15777 ( .A(n13942), .B(P1_DATAO_REG_27__SCAN_IN), .S(n13793), .Z(
        P1_U3587) );
  MUX2_X1 U15778 ( .A(n13962), .B(P1_DATAO_REG_26__SCAN_IN), .S(n13793), .Z(
        P1_U3586) );
  MUX2_X1 U15779 ( .A(n13773), .B(P1_DATAO_REG_25__SCAN_IN), .S(n13793), .Z(
        P1_U3585) );
  MUX2_X1 U15780 ( .A(n13774), .B(P1_DATAO_REG_24__SCAN_IN), .S(n13793), .Z(
        P1_U3584) );
  MUX2_X1 U15781 ( .A(n14037), .B(P1_DATAO_REG_23__SCAN_IN), .S(n13793), .Z(
        P1_U3583) );
  MUX2_X1 U15782 ( .A(n13775), .B(P1_DATAO_REG_22__SCAN_IN), .S(n13793), .Z(
        P1_U3582) );
  MUX2_X1 U15783 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14062), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U15784 ( .A(n13916), .B(P1_DATAO_REG_20__SCAN_IN), .S(n13793), .Z(
        P1_U3580) );
  MUX2_X1 U15785 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n13896), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15786 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n13913), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U15787 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14136), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U15788 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n13889), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U15789 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14134), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U15790 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13776), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15791 ( .A(n13777), .B(P1_DATAO_REG_13__SCAN_IN), .S(n13793), .Z(
        P1_U3573) );
  MUX2_X1 U15792 ( .A(n13778), .B(P1_DATAO_REG_12__SCAN_IN), .S(n13793), .Z(
        P1_U3572) );
  MUX2_X1 U15793 ( .A(n13779), .B(P1_DATAO_REG_11__SCAN_IN), .S(n13793), .Z(
        P1_U3571) );
  MUX2_X1 U15794 ( .A(n13780), .B(P1_DATAO_REG_10__SCAN_IN), .S(n13793), .Z(
        P1_U3570) );
  MUX2_X1 U15795 ( .A(n13781), .B(P1_DATAO_REG_9__SCAN_IN), .S(n13793), .Z(
        P1_U3569) );
  MUX2_X1 U15796 ( .A(n13782), .B(P1_DATAO_REG_8__SCAN_IN), .S(n13793), .Z(
        P1_U3568) );
  MUX2_X1 U15797 ( .A(n13783), .B(P1_DATAO_REG_7__SCAN_IN), .S(n13793), .Z(
        P1_U3567) );
  MUX2_X1 U15798 ( .A(n13784), .B(P1_DATAO_REG_6__SCAN_IN), .S(n13793), .Z(
        P1_U3566) );
  MUX2_X1 U15799 ( .A(n13785), .B(P1_DATAO_REG_5__SCAN_IN), .S(n13793), .Z(
        P1_U3565) );
  MUX2_X1 U15800 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13786), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U15801 ( .A(n13787), .B(P1_DATAO_REG_3__SCAN_IN), .S(n13793), .Z(
        P1_U3563) );
  MUX2_X1 U15802 ( .A(n13788), .B(P1_DATAO_REG_2__SCAN_IN), .S(n13793), .Z(
        P1_U3562) );
  MUX2_X1 U15803 ( .A(n13789), .B(P1_DATAO_REG_0__SCAN_IN), .S(n13793), .Z(
        P1_U3560) );
  MUX2_X1 U15804 ( .A(n13792), .B(n13791), .S(n13790), .Z(n13797) );
  AOI21_X1 U15805 ( .B1(n7224), .B2(n13794), .A(n13793), .ZN(n13795) );
  OAI21_X1 U15806 ( .B1(n13797), .B2(n13796), .A(n13795), .ZN(n13842) );
  OAI22_X1 U15807 ( .A1(n14607), .A2(n6804), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13798), .ZN(n13799) );
  AOI21_X1 U15808 ( .B1(n13852), .B2(n13800), .A(n13799), .ZN(n13811) );
  MUX2_X1 U15809 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n9689), .S(n13801), .Z(
        n13804) );
  NAND3_X1 U15810 ( .A1(n13804), .A2(n13803), .A3(n13802), .ZN(n13805) );
  NAND3_X1 U15811 ( .A1(n13873), .A2(n13813), .A3(n13805), .ZN(n13810) );
  OAI211_X1 U15812 ( .C1(n13808), .C2(n13807), .A(n14604), .B(n13806), .ZN(
        n13809) );
  NAND4_X1 U15813 ( .A1(n13842), .A2(n13811), .A3(n13810), .A4(n13809), .ZN(
        P1_U3245) );
  MUX2_X1 U15814 ( .A(n9688), .B(P1_REG2_REG_3__SCAN_IN), .S(n13821), .Z(
        n13814) );
  NAND3_X1 U15815 ( .A1(n13814), .A2(n13813), .A3(n13812), .ZN(n13815) );
  NAND3_X1 U15816 ( .A1(n13873), .A2(n13832), .A3(n13815), .ZN(n13825) );
  AND2_X1 U15817 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n13816) );
  AOI21_X1 U15818 ( .B1(n13817), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n13816), .ZN(
        n13824) );
  OAI211_X1 U15819 ( .C1(n13820), .C2(n13819), .A(n14604), .B(n13818), .ZN(
        n13823) );
  NAND2_X1 U15820 ( .A1(n13852), .A2(n13821), .ZN(n13822) );
  NAND4_X1 U15821 ( .A1(n13825), .A2(n13824), .A3(n13823), .A4(n13822), .ZN(
        P1_U3246) );
  OAI21_X1 U15822 ( .B1(n14607), .B2(n14358), .A(n13826), .ZN(n13827) );
  AOI21_X1 U15823 ( .B1(n13852), .B2(n13828), .A(n13827), .ZN(n13841) );
  INV_X1 U15824 ( .A(n13829), .ZN(n13834) );
  NAND3_X1 U15825 ( .A1(n13832), .A2(n13831), .A3(n13830), .ZN(n13833) );
  NAND3_X1 U15826 ( .A1(n13873), .A2(n13834), .A3(n13833), .ZN(n13840) );
  INV_X1 U15827 ( .A(n13835), .ZN(n13836) );
  OAI211_X1 U15828 ( .C1(n13838), .C2(n13837), .A(n14604), .B(n13836), .ZN(
        n13839) );
  NAND4_X1 U15829 ( .A1(n13842), .A2(n13841), .A3(n13840), .A4(n13839), .ZN(
        P1_U3247) );
  INV_X1 U15830 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n13844) );
  OAI21_X1 U15831 ( .B1(n14607), .B2(n13844), .A(n13843), .ZN(n13851) );
  XNOR2_X1 U15832 ( .A(n13858), .B(n13859), .ZN(n13849) );
  NOR2_X1 U15833 ( .A1(n13848), .A2(n13849), .ZN(n13861) );
  AOI211_X1 U15834 ( .C1(n13849), .C2(n13848), .A(n13861), .B(n13847), .ZN(
        n13850) );
  AOI211_X1 U15835 ( .C1(n13852), .C2(n13865), .A(n13851), .B(n13850), .ZN(
        n13857) );
  OAI21_X1 U15836 ( .B1(n11754), .B2(n13854), .A(n13853), .ZN(n13864) );
  XNOR2_X1 U15837 ( .A(n13858), .B(n13864), .ZN(n13855) );
  NAND2_X1 U15838 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n13855), .ZN(n13867) );
  OAI211_X1 U15839 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n13855), .A(n13873), 
        .B(n13867), .ZN(n13856) );
  NAND2_X1 U15840 ( .A1(n13857), .A2(n13856), .ZN(P1_U3261) );
  NOR2_X1 U15841 ( .A1(n13859), .A2(n13858), .ZN(n13860) );
  NOR2_X1 U15842 ( .A1(n13861), .A2(n13860), .ZN(n13863) );
  XOR2_X1 U15843 ( .A(n13863), .B(n13862), .Z(n13874) );
  INV_X1 U15844 ( .A(n13874), .ZN(n13871) );
  NAND2_X1 U15845 ( .A1(n13865), .A2(n13864), .ZN(n13866) );
  NAND2_X1 U15846 ( .A1(n13867), .A2(n13866), .ZN(n13868) );
  XOR2_X1 U15847 ( .A(n13868), .B(P1_REG2_REG_19__SCAN_IN), .Z(n13872) );
  OAI21_X1 U15848 ( .B1(n13872), .B2(n13869), .A(n14598), .ZN(n13870) );
  AOI21_X1 U15849 ( .B1(n13871), .B2(n14604), .A(n13870), .ZN(n13876) );
  AOI22_X1 U15850 ( .A1(n13874), .A2(n14604), .B1(n13873), .B2(n13872), .ZN(
        n13875) );
  OAI211_X1 U15851 ( .C1(n7648), .C2(n14607), .A(n13877), .B(n15237), .ZN(
        P1_U3262) );
  INV_X1 U15852 ( .A(n14167), .ZN(n13949) );
  NOR2_X1 U15853 ( .A1(n14109), .A2(n14086), .ZN(n14088) );
  NAND2_X1 U15854 ( .A1(n14218), .A2(n14088), .ZN(n14067) );
  NOR2_X1 U15855 ( .A1(n14006), .A2(n13922), .ZN(n13977) );
  NAND2_X1 U15856 ( .A1(n14149), .A2(n14146), .ZN(n13881) );
  NAND2_X1 U15857 ( .A1(n13878), .A2(P1_B_REG_SCAN_IN), .ZN(n13932) );
  NAND3_X1 U15858 ( .A1(n14135), .A2(n13879), .A3(n13932), .ZN(n14154) );
  NOR2_X1 U15859 ( .A1(n14091), .A2(n14154), .ZN(n13884) );
  AOI21_X1 U15860 ( .B1(n14091), .B2(P1_REG2_REG_31__SCAN_IN), .A(n13884), 
        .ZN(n13880) );
  OAI211_X1 U15861 ( .C1(n14151), .C2(n14125), .A(n13881), .B(n13880), .ZN(
        P1_U3263) );
  INV_X1 U15862 ( .A(n13930), .ZN(n13883) );
  NAND2_X1 U15863 ( .A1(n13883), .A2(n13882), .ZN(n14153) );
  NAND3_X1 U15864 ( .A1(n14153), .A2(n14146), .A3(n14152), .ZN(n13886) );
  AOI21_X1 U15865 ( .B1(n14091), .B2(P1_REG2_REG_30__SCAN_IN), .A(n13884), 
        .ZN(n13885) );
  OAI211_X1 U15866 ( .C1(n14156), .C2(n14125), .A(n13886), .B(n13885), .ZN(
        P1_U3264) );
  NAND2_X1 U15867 ( .A1(n14131), .A2(n14143), .ZN(n13891) );
  OR2_X1 U15868 ( .A1(n14132), .A2(n13889), .ZN(n13890) );
  OR2_X1 U15869 ( .A1(n14242), .A2(n13892), .ZN(n13893) );
  NOR2_X1 U15870 ( .A1(n14086), .A2(n13896), .ZN(n13897) );
  AND2_X2 U15871 ( .A1(n14071), .A2(n14070), .ZN(n14222) );
  NAND2_X1 U15872 ( .A1(n14179), .A2(n13962), .ZN(n13904) );
  INV_X1 U15873 ( .A(n13905), .ZN(n13954) );
  NAND2_X1 U15874 ( .A1(n14165), .A2(n13906), .ZN(n13907) );
  NAND2_X1 U15875 ( .A1(n14132), .A2(n13910), .ZN(n13911) );
  INV_X1 U15876 ( .A(n14099), .ZN(n13912) );
  NAND2_X1 U15877 ( .A1(n14110), .A2(n13913), .ZN(n13914) );
  NAND2_X1 U15878 ( .A1(n14002), .A2(n14001), .ZN(n14000) );
  XNOR2_X1 U15879 ( .A(n13927), .B(n13926), .ZN(n13928) );
  NAND2_X1 U15880 ( .A1(n14133), .A2(n13961), .ZN(n14157) );
  NAND2_X1 U15881 ( .A1(n14162), .A2(n14157), .ZN(n13929) );
  NAND2_X1 U15882 ( .A1(n13929), .A2(n14613), .ZN(n13939) );
  AOI21_X1 U15883 ( .B1(n13931), .B2(n13947), .A(n13930), .ZN(n14161) );
  NAND3_X1 U15884 ( .A1(n14135), .A2(n13933), .A3(n13932), .ZN(n14158) );
  OAI22_X1 U15885 ( .A1(n14158), .A2(n14009), .B1(n14638), .B2(n13934), .ZN(
        n13935) );
  AOI21_X1 U15886 ( .B1(P1_REG2_REG_29__SCAN_IN), .B2(n14091), .A(n13935), 
        .ZN(n13936) );
  OAI21_X1 U15887 ( .B1(n14159), .B2(n14125), .A(n13936), .ZN(n13937) );
  AOI21_X1 U15888 ( .B1(n14161), .B2(n14146), .A(n13937), .ZN(n13938) );
  OAI211_X1 U15889 ( .C1(n14164), .C2(n14148), .A(n13939), .B(n13938), .ZN(
        P1_U3356) );
  XNOR2_X1 U15890 ( .A(n13940), .B(n13954), .ZN(n13946) );
  NAND2_X1 U15891 ( .A1(n13941), .A2(n14135), .ZN(n13944) );
  NAND2_X1 U15892 ( .A1(n13942), .A2(n14133), .ZN(n13943) );
  AOI21_X1 U15893 ( .B1(n14167), .B2(n6826), .A(n13948), .ZN(n14168) );
  NOR2_X1 U15894 ( .A1(n13949), .A2(n14125), .ZN(n13953) );
  OAI22_X1 U15895 ( .A1(n14613), .A2(n13951), .B1(n13950), .B2(n14638), .ZN(
        n13952) );
  AOI211_X1 U15896 ( .C1(n14168), .C2(n14146), .A(n13953), .B(n13952), .ZN(
        n13957) );
  NAND3_X1 U15897 ( .A1(n14166), .A2(n14165), .A3(n14621), .ZN(n13956) );
  OAI211_X1 U15898 ( .C1(n14170), .C2(n14091), .A(n13957), .B(n13956), .ZN(
        P1_U3265) );
  AOI22_X1 U15899 ( .A1(n14133), .A2(n13962), .B1(n14135), .B2(n13961), .ZN(
        n13963) );
  AOI21_X1 U15900 ( .B1(n14171), .B2(n13976), .A(n13964), .ZN(n14172) );
  INV_X1 U15901 ( .A(n13965), .ZN(n13966) );
  AOI22_X1 U15902 ( .A1(n14091), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n13966), 
        .B2(n14089), .ZN(n13967) );
  OAI21_X1 U15903 ( .B1(n13968), .B2(n14125), .A(n13967), .ZN(n13970) );
  NOR2_X1 U15904 ( .A1(n14174), .A2(n14117), .ZN(n13969) );
  AOI211_X1 U15905 ( .C1(n14172), .C2(n14146), .A(n13970), .B(n13969), .ZN(
        n13971) );
  OAI21_X1 U15906 ( .B1(n13973), .B2(n13974), .A(n13972), .ZN(n14182) );
  XNOR2_X1 U15907 ( .A(n13974), .B(n13975), .ZN(n14175) );
  NAND2_X1 U15908 ( .A1(n14175), .A2(n14128), .ZN(n13986) );
  OAI21_X1 U15909 ( .B1(n13982), .B2(n13977), .A(n13976), .ZN(n14176) );
  INV_X1 U15910 ( .A(n14176), .ZN(n13984) );
  INV_X1 U15911 ( .A(n14178), .ZN(n13979) );
  OAI22_X1 U15912 ( .A1(n14091), .A2(n13979), .B1(n13978), .B2(n14638), .ZN(
        n13980) );
  AOI21_X1 U15913 ( .B1(P1_REG2_REG_26__SCAN_IN), .B2(n14091), .A(n13980), 
        .ZN(n13981) );
  OAI21_X1 U15914 ( .B1(n13982), .B2(n14125), .A(n13981), .ZN(n13983) );
  AOI21_X1 U15915 ( .B1(n13984), .B2(n14146), .A(n13983), .ZN(n13985) );
  OAI211_X1 U15916 ( .C1(n14182), .C2(n14148), .A(n13986), .B(n13985), .ZN(
        P1_U3267) );
  AOI21_X1 U15917 ( .B1(n13994), .B2(n13988), .A(n13987), .ZN(n14191) );
  XNOR2_X1 U15918 ( .A(n14183), .B(n14006), .ZN(n14186) );
  NAND2_X1 U15919 ( .A1(n14091), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n13992) );
  NOR2_X1 U15920 ( .A1(n14638), .A2(n13989), .ZN(n13990) );
  OAI21_X1 U15921 ( .B1(n13990), .B2(n14185), .A(n14613), .ZN(n13991) );
  OAI211_X1 U15922 ( .C1(n14183), .C2(n14125), .A(n13992), .B(n13991), .ZN(
        n13993) );
  AOI21_X1 U15923 ( .B1(n14186), .B2(n14146), .A(n13993), .ZN(n13997) );
  OR2_X1 U15924 ( .A1(n13995), .A2(n13994), .ZN(n14188) );
  NAND3_X1 U15925 ( .A1(n14188), .A2(n14187), .A3(n14621), .ZN(n13996) );
  OAI211_X1 U15926 ( .C1(n14191), .C2(n14633), .A(n13997), .B(n13996), .ZN(
        P1_U3268) );
  AOI21_X1 U15927 ( .B1(n14001), .B2(n13999), .A(n13998), .ZN(n14196) );
  OAI211_X1 U15928 ( .C1(n14002), .C2(n14001), .A(n14000), .B(n14245), .ZN(
        n14003) );
  OAI211_X1 U15929 ( .C1(n14196), .C2(n14105), .A(n14004), .B(n14003), .ZN(
        n14005) );
  INV_X1 U15930 ( .A(n14005), .ZN(n14195) );
  INV_X1 U15931 ( .A(n14006), .ZN(n14007) );
  AOI211_X1 U15932 ( .C1(n14193), .C2(n6819), .A(n14662), .B(n14007), .ZN(
        n14192) );
  NOR2_X1 U15933 ( .A1(n14009), .A2(n14008), .ZN(n14629) );
  AOI22_X1 U15934 ( .A1(n14091), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n14010), 
        .B2(n14089), .ZN(n14011) );
  OAI21_X1 U15935 ( .B1(n14012), .B2(n14125), .A(n14011), .ZN(n14014) );
  NOR2_X1 U15936 ( .A1(n14196), .A2(n14117), .ZN(n14013) );
  AOI211_X1 U15937 ( .C1(n14192), .C2(n14629), .A(n14014), .B(n14013), .ZN(
        n14015) );
  OAI21_X1 U15938 ( .B1(n14091), .B2(n14195), .A(n14015), .ZN(P1_U3269) );
  XNOR2_X1 U15939 ( .A(n14016), .B(n14023), .ZN(n14205) );
  AOI21_X1 U15940 ( .B1(n14017), .B2(n14028), .A(n7210), .ZN(n14200) );
  NAND2_X1 U15941 ( .A1(n14091), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n14021) );
  NOR2_X1 U15942 ( .A1(n14638), .A2(n14018), .ZN(n14019) );
  OAI21_X1 U15943 ( .B1(n14198), .B2(n14019), .A(n14613), .ZN(n14020) );
  OAI211_X1 U15944 ( .C1(n14197), .C2(n14125), .A(n14021), .B(n14020), .ZN(
        n14022) );
  AOI21_X1 U15945 ( .B1(n14200), .B2(n14146), .A(n14022), .ZN(n14026) );
  OR2_X1 U15946 ( .A1(n14024), .A2(n14023), .ZN(n14202) );
  NAND3_X1 U15947 ( .A1(n14202), .A2(n14201), .A3(n14621), .ZN(n14025) );
  OAI211_X1 U15948 ( .C1(n14205), .C2(n14633), .A(n14026), .B(n14025), .ZN(
        P1_U3270) );
  XNOR2_X1 U15949 ( .A(n14027), .B(n14036), .ZN(n14210) );
  INV_X1 U15950 ( .A(n14028), .ZN(n14029) );
  AOI21_X1 U15951 ( .B1(n14206), .B2(n14049), .A(n14029), .ZN(n14207) );
  INV_X1 U15952 ( .A(n14030), .ZN(n14031) );
  AOI22_X1 U15953 ( .A1(n14031), .A2(n14089), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n14091), .ZN(n14032) );
  OAI21_X1 U15954 ( .B1(n14033), .B2(n14125), .A(n14032), .ZN(n14040) );
  OAI21_X1 U15955 ( .B1(n14036), .B2(n14035), .A(n14034), .ZN(n14038) );
  AOI222_X1 U15956 ( .A1(n14245), .A2(n14038), .B1(n14037), .B2(n14135), .C1(
        n14062), .C2(n14133), .ZN(n14209) );
  NOR2_X1 U15957 ( .A1(n14209), .A2(n14091), .ZN(n14039) );
  AOI211_X1 U15958 ( .C1(n14207), .C2(n14146), .A(n14040), .B(n14039), .ZN(
        n14041) );
  OAI21_X1 U15959 ( .B1(n14210), .B2(n14148), .A(n14041), .ZN(P1_U3271) );
  AOI211_X1 U15960 ( .C1(n14047), .C2(n14042), .A(n14672), .B(n6470), .ZN(
        n14045) );
  OAI22_X1 U15961 ( .A1(n14043), .A2(n14102), .B1(n14080), .B2(n14078), .ZN(
        n14044) );
  NOR2_X1 U15962 ( .A1(n14045), .A2(n14044), .ZN(n14215) );
  OAI21_X1 U15963 ( .B1(n14048), .B2(n14047), .A(n14046), .ZN(n14211) );
  AOI21_X1 U15964 ( .B1(n14212), .B2(n14067), .A(n7211), .ZN(n14213) );
  NAND2_X1 U15965 ( .A1(n14213), .A2(n14146), .ZN(n14053) );
  INV_X1 U15966 ( .A(n14050), .ZN(n14051) );
  AOI22_X1 U15967 ( .A1(n14051), .A2(n14089), .B1(n14091), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n14052) );
  OAI211_X1 U15968 ( .C1(n6818), .C2(n14125), .A(n14053), .B(n14052), .ZN(
        n14054) );
  AOI21_X1 U15969 ( .B1(n14211), .B2(n14621), .A(n14054), .ZN(n14055) );
  OAI21_X1 U15970 ( .B1(n14215), .B2(n14091), .A(n14055), .ZN(P1_U3272) );
  INV_X1 U15971 ( .A(n14056), .ZN(n14065) );
  NAND2_X1 U15972 ( .A1(n14057), .A2(n14070), .ZN(n14058) );
  NAND2_X1 U15973 ( .A1(n14058), .A2(n14245), .ZN(n14059) );
  OR2_X1 U15974 ( .A1(n14060), .A2(n14059), .ZN(n14064) );
  NOR2_X1 U15975 ( .A1(n14103), .A2(n14078), .ZN(n14061) );
  AOI21_X1 U15976 ( .B1(n14062), .B2(n14135), .A(n14061), .ZN(n14063) );
  NAND2_X1 U15977 ( .A1(n14064), .A2(n14063), .ZN(n14224) );
  AOI21_X1 U15978 ( .B1(n14065), .B2(n14089), .A(n14224), .ZN(n14075) );
  OR2_X1 U15979 ( .A1(n14218), .A2(n14088), .ZN(n14066) );
  AND2_X1 U15980 ( .A1(n14067), .A2(n14066), .ZN(n14220) );
  INV_X1 U15981 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n14068) );
  OAI22_X1 U15982 ( .A1(n14218), .A2(n14125), .B1(n14068), .B2(n14613), .ZN(
        n14069) );
  AOI21_X1 U15983 ( .B1(n14220), .B2(n14146), .A(n14069), .ZN(n14074) );
  INV_X1 U15984 ( .A(n14222), .ZN(n14072) );
  OR2_X1 U15985 ( .A1(n14071), .A2(n14070), .ZN(n14217) );
  NAND3_X1 U15986 ( .A1(n14072), .A2(n14621), .A3(n14217), .ZN(n14073) );
  OAI211_X1 U15987 ( .C1(n14075), .C2(n14091), .A(n14074), .B(n14073), .ZN(
        P1_U3273) );
  XNOR2_X1 U15988 ( .A(n14076), .B(n14084), .ZN(n14077) );
  NAND2_X1 U15989 ( .A1(n14077), .A2(n14245), .ZN(n14083) );
  OAI22_X1 U15990 ( .A1(n14080), .A2(n14102), .B1(n14079), .B2(n14078), .ZN(
        n14081) );
  INV_X1 U15991 ( .A(n14081), .ZN(n14082) );
  NAND2_X1 U15992 ( .A1(n14083), .A2(n14082), .ZN(n14233) );
  INV_X1 U15993 ( .A(n14233), .ZN(n14096) );
  XNOR2_X1 U15994 ( .A(n14085), .B(n14084), .ZN(n14228) );
  AND2_X1 U15995 ( .A1(n14109), .A2(n14086), .ZN(n14087) );
  OR2_X1 U15996 ( .A1(n14088), .A2(n14087), .ZN(n14230) );
  NOR2_X1 U15997 ( .A1(n14230), .A2(n14111), .ZN(n14094) );
  AOI22_X1 U15998 ( .A1(n14091), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n14090), 
        .B2(n14089), .ZN(n14092) );
  OAI21_X1 U15999 ( .B1(n14229), .B2(n14125), .A(n14092), .ZN(n14093) );
  AOI211_X1 U16000 ( .C1(n14228), .C2(n14621), .A(n14094), .B(n14093), .ZN(
        n14095) );
  OAI21_X1 U16001 ( .B1(n14096), .B2(n14091), .A(n14095), .ZN(P1_U3274) );
  XNOR2_X1 U16002 ( .A(n14097), .B(n14099), .ZN(n14240) );
  AOI21_X1 U16003 ( .B1(n7351), .B2(n14099), .A(n14672), .ZN(n14101) );
  AOI22_X1 U16004 ( .A1(n14101), .A2(n14100), .B1(n14133), .B2(n14136), .ZN(
        n14239) );
  NOR2_X1 U16005 ( .A1(n14103), .A2(n14102), .ZN(n14236) );
  INV_X1 U16006 ( .A(n14236), .ZN(n14104) );
  OAI211_X1 U16007 ( .C1(n14240), .C2(n14105), .A(n14239), .B(n14104), .ZN(
        n14106) );
  NAND2_X1 U16008 ( .A1(n14106), .A2(n14613), .ZN(n14116) );
  INV_X1 U16009 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14108) );
  OAI22_X1 U16010 ( .A1(n14613), .A2(n14108), .B1(n14107), .B2(n14638), .ZN(
        n14113) );
  OAI21_X1 U16011 ( .B1(n14110), .B2(n14120), .A(n14109), .ZN(n14234) );
  NOR2_X1 U16012 ( .A1(n14234), .A2(n14111), .ZN(n14112) );
  AOI211_X1 U16013 ( .C1(n14114), .C2(n14237), .A(n14113), .B(n14112), .ZN(
        n14115) );
  OAI211_X1 U16014 ( .C1(n14240), .C2(n14117), .A(n14116), .B(n14115), .ZN(
        P1_U3275) );
  XNOR2_X1 U16015 ( .A(n14118), .B(n14127), .ZN(n14249) );
  NOR2_X1 U16016 ( .A1(n6530), .A2(n14242), .ZN(n14119) );
  INV_X1 U16017 ( .A(n14121), .ZN(n14122) );
  OAI22_X1 U16018 ( .A1(n14241), .A2(n14091), .B1(n14122), .B2(n14638), .ZN(
        n14123) );
  AOI21_X1 U16019 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n14091), .A(n14123), 
        .ZN(n14124) );
  OAI21_X1 U16020 ( .B1(n14242), .B2(n14125), .A(n14124), .ZN(n14126) );
  AOI21_X1 U16021 ( .B1(n7610), .B2(n14146), .A(n14126), .ZN(n14130) );
  OR2_X1 U16022 ( .A1(n6544), .A2(n14127), .ZN(n14246) );
  NAND3_X1 U16023 ( .A1(n14246), .A2(n14128), .A3(n14244), .ZN(n14129) );
  OAI211_X1 U16024 ( .C1(n14249), .C2(n14148), .A(n14130), .B(n14129), .ZN(
        P1_U3276) );
  XOR2_X1 U16025 ( .A(n14131), .B(n14143), .Z(n14256) );
  AOI21_X1 U16026 ( .B1(n14132), .B2(n6422), .A(n6530), .ZN(n14254) );
  AOI22_X1 U16027 ( .A1(n14136), .A2(n14135), .B1(n14134), .B2(n14133), .ZN(
        n14250) );
  OAI22_X1 U16028 ( .A1(n14091), .A2(n14250), .B1(n14137), .B2(n14638), .ZN(
        n14138) );
  AOI21_X1 U16029 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n14091), .A(n14138), 
        .ZN(n14139) );
  OAI21_X1 U16030 ( .B1(n7217), .B2(n14125), .A(n14139), .ZN(n14145) );
  INV_X1 U16031 ( .A(n14140), .ZN(n14141) );
  AOI21_X1 U16032 ( .B1(n14143), .B2(n14142), .A(n14141), .ZN(n14251) );
  NOR2_X1 U16033 ( .A1(n14251), .A2(n14633), .ZN(n14144) );
  AOI211_X1 U16034 ( .C1(n14254), .C2(n14146), .A(n14145), .B(n14144), .ZN(
        n14147) );
  OAI21_X1 U16035 ( .B1(n14148), .B2(n14256), .A(n14147), .ZN(P1_U3277) );
  NAND2_X1 U16036 ( .A1(n14149), .A2(n14654), .ZN(n14150) );
  OAI211_X1 U16037 ( .C1(n14151), .C2(n14670), .A(n14150), .B(n14154), .ZN(
        n14259) );
  MUX2_X1 U16038 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14259), .S(n14687), .Z(
        P1_U3559) );
  NAND3_X1 U16039 ( .A1(n14153), .A2(n14654), .A3(n14152), .ZN(n14155) );
  OAI211_X1 U16040 ( .C1(n14156), .C2(n14670), .A(n14155), .B(n14154), .ZN(
        n14260) );
  MUX2_X1 U16041 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14260), .S(n14687), .Z(
        P1_U3558) );
  OAI211_X1 U16042 ( .C1(n14159), .C2(n14670), .A(n14158), .B(n14157), .ZN(
        n14160) );
  AOI21_X1 U16043 ( .B1(n14161), .B2(n14654), .A(n14160), .ZN(n14163) );
  MUX2_X1 U16044 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14261), .S(n14687), .Z(
        P1_U3557) );
  NAND3_X1 U16045 ( .A1(n14166), .A2(n14165), .A3(n14677), .ZN(n14169) );
  AOI22_X1 U16046 ( .A1(n14172), .A2(n14654), .B1(n14653), .B2(n14171), .ZN(
        n14173) );
  MUX2_X1 U16047 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14263), .S(n14687), .Z(
        P1_U3555) );
  NAND2_X1 U16048 ( .A1(n14175), .A2(n14245), .ZN(n14181) );
  NOR2_X1 U16049 ( .A1(n14176), .A2(n14662), .ZN(n14177) );
  AOI211_X1 U16050 ( .C1(n14653), .C2(n14179), .A(n14178), .B(n14177), .ZN(
        n14180) );
  OAI211_X1 U16051 ( .C1(n14257), .C2(n14182), .A(n14181), .B(n14180), .ZN(
        n14264) );
  MUX2_X1 U16052 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14264), .S(n14687), .Z(
        P1_U3554) );
  NOR2_X1 U16053 ( .A1(n14183), .A2(n14670), .ZN(n14184) );
  AOI211_X1 U16054 ( .C1(n14186), .C2(n14654), .A(n14185), .B(n14184), .ZN(
        n14190) );
  NAND3_X1 U16055 ( .A1(n14188), .A2(n14187), .A3(n14677), .ZN(n14189) );
  OAI211_X1 U16056 ( .C1(n14191), .C2(n14672), .A(n14190), .B(n14189), .ZN(
        n14265) );
  MUX2_X1 U16057 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14265), .S(n14687), .Z(
        P1_U3553) );
  AOI21_X1 U16058 ( .B1(n14653), .B2(n14193), .A(n14192), .ZN(n14194) );
  OAI211_X1 U16059 ( .C1(n14196), .C2(n14658), .A(n14195), .B(n14194), .ZN(
        n14266) );
  MUX2_X1 U16060 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14266), .S(n14687), .Z(
        P1_U3552) );
  NOR2_X1 U16061 ( .A1(n14197), .A2(n14670), .ZN(n14199) );
  AOI211_X1 U16062 ( .C1(n14200), .C2(n14654), .A(n14199), .B(n14198), .ZN(
        n14204) );
  NAND3_X1 U16063 ( .A1(n14202), .A2(n14201), .A3(n14677), .ZN(n14203) );
  OAI211_X1 U16064 ( .C1(n14205), .C2(n14672), .A(n14204), .B(n14203), .ZN(
        n14267) );
  MUX2_X1 U16065 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14267), .S(n14687), .Z(
        P1_U3551) );
  AOI22_X1 U16066 ( .A1(n14207), .A2(n14654), .B1(n14206), .B2(n14653), .ZN(
        n14208) );
  OAI211_X1 U16067 ( .C1(n14257), .C2(n14210), .A(n14209), .B(n14208), .ZN(
        n14268) );
  MUX2_X1 U16068 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14268), .S(n14687), .Z(
        P1_U3550) );
  INV_X1 U16069 ( .A(n14211), .ZN(n14216) );
  AOI22_X1 U16070 ( .A1(n14213), .A2(n14654), .B1(n14653), .B2(n14212), .ZN(
        n14214) );
  OAI211_X1 U16071 ( .C1(n14257), .C2(n14216), .A(n14215), .B(n14214), .ZN(
        n14269) );
  MUX2_X1 U16072 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14269), .S(n14687), .Z(
        P1_U3549) );
  INV_X1 U16073 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n14226) );
  NAND2_X1 U16074 ( .A1(n14217), .A2(n14677), .ZN(n14223) );
  NOR2_X1 U16075 ( .A1(n14218), .A2(n14670), .ZN(n14219) );
  AOI21_X1 U16076 ( .B1(n14220), .B2(n14654), .A(n14219), .ZN(n14221) );
  OAI21_X1 U16077 ( .B1(n14223), .B2(n14222), .A(n14221), .ZN(n14225) );
  NOR2_X1 U16078 ( .A1(n14225), .A2(n14224), .ZN(n14270) );
  MUX2_X1 U16079 ( .A(n14226), .B(n14270), .S(n14687), .Z(n14227) );
  INV_X1 U16080 ( .A(n14227), .ZN(P1_U3548) );
  AND2_X1 U16081 ( .A1(n14228), .A2(n14677), .ZN(n14232) );
  OAI22_X1 U16082 ( .A1(n14230), .A2(n14662), .B1(n14229), .B2(n14670), .ZN(
        n14231) );
  MUX2_X1 U16083 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14272), .S(n14687), .Z(
        P1_U3547) );
  NOR2_X1 U16084 ( .A1(n14234), .A2(n14662), .ZN(n14235) );
  AOI211_X1 U16085 ( .C1(n14653), .C2(n14237), .A(n14236), .B(n14235), .ZN(
        n14238) );
  OAI211_X1 U16086 ( .C1(n14257), .C2(n14240), .A(n14239), .B(n14238), .ZN(
        n14273) );
  MUX2_X1 U16087 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14273), .S(n14687), .Z(
        P1_U3546) );
  OAI21_X1 U16088 ( .B1(n14242), .B2(n14670), .A(n14241), .ZN(n14243) );
  AOI21_X1 U16089 ( .B1(n7610), .B2(n14654), .A(n14243), .ZN(n14248) );
  NAND3_X1 U16090 ( .A1(n14246), .A2(n14245), .A3(n14244), .ZN(n14247) );
  OAI211_X1 U16091 ( .C1(n14257), .C2(n14249), .A(n14248), .B(n14247), .ZN(
        n14274) );
  MUX2_X1 U16092 ( .A(n14274), .B(P1_REG1_REG_17__SCAN_IN), .S(n14685), .Z(
        P1_U3545) );
  OAI21_X1 U16093 ( .B1(n7217), .B2(n14670), .A(n14250), .ZN(n14253) );
  NOR2_X1 U16094 ( .A1(n14251), .A2(n14672), .ZN(n14252) );
  AOI211_X1 U16095 ( .C1(n14654), .C2(n14254), .A(n14253), .B(n14252), .ZN(
        n14255) );
  OAI21_X1 U16096 ( .B1(n14257), .B2(n14256), .A(n14255), .ZN(n14275) );
  MUX2_X1 U16097 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14275), .S(n14687), .Z(
        P1_U3544) );
  MUX2_X1 U16098 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n14258), .S(n14687), .Z(
        P1_U3528) );
  MUX2_X1 U16099 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14259), .S(n14679), .Z(
        P1_U3527) );
  MUX2_X1 U16100 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14260), .S(n14679), .Z(
        P1_U3526) );
  MUX2_X1 U16101 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14261), .S(n14679), .Z(
        P1_U3525) );
  MUX2_X1 U16102 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14263), .S(n14679), .Z(
        P1_U3523) );
  MUX2_X1 U16103 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14264), .S(n14679), .Z(
        P1_U3522) );
  MUX2_X1 U16104 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14265), .S(n14679), .Z(
        P1_U3521) );
  MUX2_X1 U16105 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14266), .S(n14679), .Z(
        P1_U3520) );
  MUX2_X1 U16106 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14267), .S(n14679), .Z(
        P1_U3519) );
  MUX2_X1 U16107 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14268), .S(n14679), .Z(
        P1_U3518) );
  MUX2_X1 U16108 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14269), .S(n14679), .Z(
        P1_U3517) );
  MUX2_X1 U16109 ( .A(n15155), .B(n14270), .S(n14679), .Z(n14271) );
  INV_X1 U16110 ( .A(n14271), .ZN(P1_U3516) );
  MUX2_X1 U16111 ( .A(n14272), .B(P1_REG0_REG_19__SCAN_IN), .S(n14678), .Z(
        P1_U3515) );
  MUX2_X1 U16112 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14273), .S(n14679), .Z(
        P1_U3513) );
  MUX2_X1 U16113 ( .A(n14274), .B(P1_REG0_REG_17__SCAN_IN), .S(n14678), .Z(
        P1_U3510) );
  MUX2_X1 U16114 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14275), .S(n14679), .Z(
        P1_U3507) );
  INV_X1 U16115 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n14276) );
  NAND3_X1 U16116 ( .A1(n14276), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n14277) );
  INV_X1 U16117 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n15130) );
  OAI22_X1 U16118 ( .A1(n14278), .A2(n14277), .B1(n15130), .B2(n14298), .ZN(
        n14279) );
  AOI21_X1 U16119 ( .B1(n13586), .B2(n14280), .A(n14279), .ZN(n14281) );
  INV_X1 U16120 ( .A(n14281), .ZN(P1_U3324) );
  OAI222_X1 U16121 ( .A1(P1_U3086), .A2(n14284), .B1(n14300), .B2(n14283), 
        .C1(n14282), .C2(n14298), .ZN(P1_U3325) );
  OAI222_X1 U16122 ( .A1(P1_U3086), .A2(n14287), .B1(n14300), .B2(n14286), 
        .C1(n14285), .C2(n14298), .ZN(P1_U3326) );
  NAND2_X1 U16123 ( .A1(n14288), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n14289) );
  OAI211_X1 U16124 ( .C1(n14291), .C2(n14300), .A(n14290), .B(n14289), .ZN(
        P1_U3328) );
  OAI222_X1 U16125 ( .A1(n14294), .A2(P1_U3086), .B1(n14300), .B2(n14293), 
        .C1(n14292), .C2(n14298), .ZN(P1_U3329) );
  OAI222_X1 U16126 ( .A1(P1_U3086), .A2(n14297), .B1(n14300), .B2(n14296), 
        .C1(n14295), .C2(n14298), .ZN(P1_U3330) );
  OAI222_X1 U16127 ( .A1(P1_U3086), .A2(n14301), .B1(n14300), .B2(n14299), 
        .C1(n7156), .C2(n14298), .ZN(P1_U3331) );
  MUX2_X1 U16128 ( .A(n14304), .B(n14303), .S(P1_U3086), .Z(P1_U3333) );
  INV_X1 U16129 ( .A(n14305), .ZN(n14306) );
  MUX2_X1 U16130 ( .A(n14306), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XNOR2_X1 U16131 ( .A(n12558), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(n14446) );
  INV_X1 U16132 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14345) );
  INV_X1 U16133 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n14339) );
  XNOR2_X1 U16134 ( .A(n14339), .B(P1_ADDR_REG_14__SCAN_IN), .ZN(n14351) );
  INV_X1 U16135 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n15238) );
  INV_X1 U16136 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n14336) );
  INV_X1 U16137 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n15174) );
  INV_X1 U16138 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n15013) );
  XOR2_X1 U16139 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n14311), .Z(n14361) );
  NAND2_X1 U16140 ( .A1(n9595), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14365) );
  INV_X1 U16141 ( .A(n14365), .ZN(n14307) );
  NAND2_X1 U16142 ( .A1(n14307), .A2(n14363), .ZN(n14308) );
  NAND2_X1 U16143 ( .A1(n14361), .A2(n14362), .ZN(n14310) );
  INV_X1 U16144 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14359) );
  NAND2_X1 U16145 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n14312), .ZN(n14313) );
  NAND2_X1 U16146 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n14315), .ZN(n14316) );
  NAND2_X1 U16147 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n14317), .ZN(n14319) );
  INV_X1 U16148 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14373) );
  NOR2_X1 U16149 ( .A1(n14321), .A2(n15232), .ZN(n14323) );
  INV_X1 U16150 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n14324) );
  NOR2_X1 U16151 ( .A1(n14325), .A2(n14324), .ZN(n14327) );
  INV_X1 U16152 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n14329) );
  NOR2_X1 U16153 ( .A1(n14328), .A2(n14329), .ZN(n14331) );
  INV_X1 U16154 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n15202) );
  XOR2_X1 U16155 ( .A(n14329), .B(n14328), .Z(n14356) );
  XNOR2_X1 U16156 ( .A(n15013), .B(P1_ADDR_REG_10__SCAN_IN), .ZN(n14354) );
  XNOR2_X1 U16157 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n14390) );
  NAND2_X1 U16158 ( .A1(n14391), .A2(n14390), .ZN(n14333) );
  OAI21_X1 U16159 ( .B1(n15174), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n14333), 
        .ZN(n14334) );
  INV_X1 U16160 ( .A(n14334), .ZN(n14353) );
  XNOR2_X1 U16161 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(n14336), .ZN(n14352) );
  AND2_X1 U16162 ( .A1(n15238), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n14337) );
  INV_X1 U16163 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15239) );
  XNOR2_X1 U16164 ( .A(n15239), .B(n14341), .ZN(n14348) );
  NAND2_X1 U16165 ( .A1(n14349), .A2(n14348), .ZN(n14340) );
  NAND2_X1 U16166 ( .A1(n11430), .A2(n14346), .ZN(n14343) );
  NOR2_X1 U16167 ( .A1(n11430), .A2(n14346), .ZN(n14342) );
  XNOR2_X1 U16168 ( .A(n14345), .B(P1_ADDR_REG_17__SCAN_IN), .ZN(n14400) );
  NOR2_X1 U16169 ( .A1(n14399), .A2(n14400), .ZN(n14344) );
  AOI21_X1 U16170 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(n14345), .A(n14344), 
        .ZN(n14447) );
  XNOR2_X1 U16171 ( .A(n14446), .B(n14447), .ZN(n14442) );
  XOR2_X1 U16172 ( .A(n15184), .B(P1_ADDR_REG_16__SCAN_IN), .Z(n14347) );
  XOR2_X1 U16173 ( .A(n14347), .B(n14346), .Z(n14591) );
  XOR2_X1 U16174 ( .A(n14349), .B(n14348), .Z(n14587) );
  XNOR2_X1 U16175 ( .A(n14351), .B(n14350), .ZN(n14584) );
  XOR2_X1 U16176 ( .A(n14353), .B(n14352), .Z(n14577) );
  XOR2_X1 U16177 ( .A(n14355), .B(n14354), .Z(n14427) );
  XOR2_X1 U16178 ( .A(n15202), .B(n14356), .Z(n14422) );
  INV_X1 U16179 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n14746) );
  NOR2_X1 U16180 ( .A1(n14370), .A2(n14746), .ZN(n14371) );
  XOR2_X1 U16181 ( .A(n14360), .B(n14359), .Z(n15283) );
  XOR2_X1 U16182 ( .A(n14362), .B(n14361), .Z(n14407) );
  XNOR2_X1 U16183 ( .A(n14365), .B(n14363), .ZN(n14366) );
  INV_X1 U16184 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n14364) );
  NOR2_X1 U16185 ( .A1(n14366), .A2(n14364), .ZN(n14367) );
  OAI21_X1 U16186 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n9595), .A(n14365), .ZN(
        n15277) );
  NAND2_X1 U16187 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15277), .ZN(n15287) );
  XOR2_X1 U16188 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n14366), .Z(n15286) );
  NOR2_X1 U16189 ( .A1(n15287), .A2(n15286), .ZN(n15285) );
  NOR2_X1 U16190 ( .A1(n14367), .A2(n15285), .ZN(n14406) );
  NOR2_X1 U16191 ( .A1(n14407), .A2(n14406), .ZN(n14368) );
  NAND2_X1 U16192 ( .A1(n14407), .A2(n14406), .ZN(n14405) );
  OAI21_X1 U16193 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(n14368), .A(n14405), .ZN(
        n15282) );
  NAND2_X1 U16194 ( .A1(n15283), .A2(n15282), .ZN(n14369) );
  NOR2_X1 U16195 ( .A1(n15283), .A2(n15282), .ZN(n15281) );
  AOI21_X1 U16196 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n14369), .A(n15281), .ZN(
        n15273) );
  NOR2_X1 U16197 ( .A1(n15273), .A2(n15272), .ZN(n15271) );
  NAND2_X1 U16198 ( .A1(n14374), .A2(n14375), .ZN(n14376) );
  INV_X1 U16199 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15275) );
  NOR2_X1 U16200 ( .A1(n14380), .A2(n7160), .ZN(n14381) );
  XOR2_X1 U16201 ( .A(n14377), .B(P3_ADDR_REG_6__SCAN_IN), .Z(n14379) );
  XOR2_X1 U16202 ( .A(n14379), .B(n14378), .Z(n14417) );
  NOR2_X1 U16203 ( .A1(n14417), .A2(n14416), .ZN(n14415) );
  NOR2_X1 U16204 ( .A1(n14384), .A2(n14382), .ZN(n14385) );
  XOR2_X1 U16205 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n14383), .Z(n15280) );
  XOR2_X1 U16206 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n14386), .Z(n14388) );
  NAND2_X1 U16207 ( .A1(n14387), .A2(n14388), .ZN(n14389) );
  INV_X1 U16208 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14419) );
  NAND2_X1 U16209 ( .A1(n14420), .A2(n14419), .ZN(n14418) );
  NAND2_X1 U16210 ( .A1(n14389), .A2(n14418), .ZN(n14423) );
  NAND2_X1 U16211 ( .A1(n14422), .A2(n14423), .ZN(n14421) );
  XNOR2_X1 U16212 ( .A(n14391), .B(n14390), .ZN(n14392) );
  INV_X1 U16213 ( .A(n14572), .ZN(n14573) );
  INV_X1 U16214 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n14575) );
  NAND2_X1 U16215 ( .A1(n14393), .A2(n14392), .ZN(n14574) );
  NAND2_X1 U16216 ( .A1(n14575), .A2(n14574), .ZN(n14571) );
  NAND2_X1 U16217 ( .A1(n14573), .A2(n14571), .ZN(n14578) );
  NAND2_X1 U16218 ( .A1(n14577), .A2(n14578), .ZN(n14576) );
  XNOR2_X1 U16219 ( .A(n15238), .B(P1_ADDR_REG_13__SCAN_IN), .ZN(n14394) );
  XOR2_X1 U16220 ( .A(n14395), .B(n14394), .Z(n14397) );
  NAND2_X1 U16221 ( .A1(n14396), .A2(n14397), .ZN(n14398) );
  INV_X1 U16222 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14778) );
  XOR2_X1 U16223 ( .A(n14400), .B(n14399), .Z(n14402) );
  INV_X1 U16224 ( .A(n14437), .ZN(n14438) );
  INV_X1 U16225 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n14440) );
  INV_X1 U16226 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n15186) );
  AOI21_X1 U16227 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14403) );
  OAI21_X1 U16228 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14403), 
        .ZN(U28) );
  AOI21_X1 U16229 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14404) );
  OAI21_X1 U16230 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14404), 
        .ZN(U29) );
  OAI21_X1 U16231 ( .B1(n14407), .B2(n14406), .A(n14405), .ZN(n14408) );
  XNOR2_X1 U16232 ( .A(n14408), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  OAI22_X1 U16233 ( .A1(n14411), .A2(n14410), .B1(n14409), .B2(n12973), .ZN(
        n14412) );
  INV_X1 U16234 ( .A(n14412), .ZN(n14413) );
  OAI21_X1 U16235 ( .B1(P3_U3151), .B2(n14414), .A(n14413), .ZN(P3_U3285) );
  AOI21_X1 U16236 ( .B1(n14417), .B2(n14416), .A(n14415), .ZN(SUB_1596_U57) );
  OAI21_X1 U16237 ( .B1(n14420), .B2(n14419), .A(n14418), .ZN(SUB_1596_U55) );
  OAI21_X1 U16238 ( .B1(n14423), .B2(n14422), .A(n14421), .ZN(n14424) );
  XNOR2_X1 U16239 ( .A(n14424), .B(P2_ADDR_REG_9__SCAN_IN), .ZN(SUB_1596_U54)
         );
  AOI21_X1 U16240 ( .B1(n14427), .B2(n14426), .A(n14425), .ZN(n14428) );
  XOR2_X1 U16241 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n14428), .Z(SUB_1596_U70)
         );
  OAI22_X1 U16242 ( .A1(n14429), .A2(n14662), .B1(n6823), .B2(n14670), .ZN(
        n14430) );
  AOI21_X1 U16243 ( .B1(n14431), .B2(n14645), .A(n14430), .ZN(n14432) );
  AND2_X1 U16244 ( .A1(n14433), .A2(n14432), .ZN(n14435) );
  INV_X1 U16245 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14434) );
  AOI22_X1 U16246 ( .A1(n14679), .A2(n14435), .B1(n14434), .B2(n14678), .ZN(
        P1_U3495) );
  AOI22_X1 U16247 ( .A1(n14687), .A2(n14435), .B1(n9187), .B2(n14685), .ZN(
        P1_U3540) );
  OAI222_X1 U16248 ( .A1(n14440), .A2(n14439), .B1(n14440), .B2(n14438), .C1(
        n14437), .C2(n14436), .ZN(SUB_1596_U63) );
  XNOR2_X1 U16249 ( .A(n14444), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n14445) );
  NOR2_X1 U16250 ( .A1(n14447), .A2(n14446), .ZN(n14448) );
  AOI21_X1 U16251 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n12558), .A(n14448), 
        .ZN(n14449) );
  AOI22_X1 U16252 ( .A1(n15010), .A2(n14450), .B1(n14982), .B2(
        P3_ADDR_REG_17__SCAN_IN), .ZN(n14464) );
  XOR2_X1 U16253 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n14451), .Z(n14456) );
  AOI211_X1 U16254 ( .C1(n14454), .C2(n14453), .A(n14999), .B(n14452), .ZN(
        n14455) );
  AOI21_X1 U16255 ( .B1(n14456), .B2(n14993), .A(n14455), .ZN(n14463) );
  NAND2_X1 U16256 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(P3_U3151), .ZN(n14462)
         );
  OAI221_X1 U16257 ( .B1(n14460), .B2(n14459), .C1(n14460), .C2(n14458), .A(
        n14457), .ZN(n14461) );
  NAND4_X1 U16258 ( .A1(n14464), .A2(n14463), .A3(n14462), .A4(n14461), .ZN(
        P3_U3199) );
  INV_X1 U16259 ( .A(n14465), .ZN(n14469) );
  AOI21_X1 U16260 ( .B1(n12815), .B2(n14467), .A(n14466), .ZN(n14468) );
  NOR3_X1 U16261 ( .A1(n14469), .A2(n14468), .A3(n15072), .ZN(n14473) );
  OAI22_X1 U16262 ( .A1(n14471), .A2(n15046), .B1(n14470), .B2(n15044), .ZN(
        n14472) );
  NOR2_X1 U16263 ( .A1(n14473), .A2(n14472), .ZN(n14487) );
  XNOR2_X1 U16264 ( .A(n14475), .B(n14474), .ZN(n14491) );
  AOI222_X1 U16265 ( .A1(n14477), .A2(n10664), .B1(n14491), .B2(n14476), .C1(
        n14486), .C2(n15034), .ZN(n14478) );
  OAI221_X1 U16266 ( .B1(n12826), .B2(n14487), .C1(n15036), .C2(n14479), .A(
        n14478), .ZN(P3_U3221) );
  NOR2_X1 U16267 ( .A1(n14480), .A2(n14494), .ZN(n14483) );
  INV_X1 U16268 ( .A(n14481), .ZN(n14482) );
  AOI211_X1 U16269 ( .C1(n15073), .C2(n14484), .A(n14483), .B(n14482), .ZN(
        n14499) );
  INV_X1 U16270 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n14485) );
  AOI22_X1 U16271 ( .A1(n15117), .A2(n14499), .B1(n14485), .B2(n15114), .ZN(
        P3_U3472) );
  INV_X1 U16272 ( .A(n14486), .ZN(n14488) );
  OAI21_X1 U16273 ( .B1(n14488), .B2(n15100), .A(n14487), .ZN(n14489) );
  AOI21_X1 U16274 ( .B1(n14491), .B2(n14490), .A(n14489), .ZN(n14501) );
  AOI22_X1 U16275 ( .A1(n15117), .A2(n14501), .B1(n14492), .B2(n15114), .ZN(
        P3_U3471) );
  OAI22_X1 U16276 ( .A1(n14495), .A2(n14494), .B1(n14493), .B2(n15100), .ZN(
        n14496) );
  NOR2_X1 U16277 ( .A1(n14497), .A2(n14496), .ZN(n14503) );
  INV_X1 U16278 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14498) );
  AOI22_X1 U16279 ( .A1(n15117), .A2(n14503), .B1(n14498), .B2(n15114), .ZN(
        P3_U3470) );
  INV_X1 U16280 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14500) );
  AOI22_X1 U16281 ( .A1(n15110), .A2(n14500), .B1(n14499), .B2(n15108), .ZN(
        P3_U3429) );
  INV_X1 U16282 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14502) );
  AOI22_X1 U16283 ( .A1(n15110), .A2(n14502), .B1(n14501), .B2(n15108), .ZN(
        P3_U3426) );
  INV_X1 U16284 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14504) );
  AOI22_X1 U16285 ( .A1(n15110), .A2(n14504), .B1(n14503), .B2(n15108), .ZN(
        P3_U3423) );
  NAND2_X1 U16286 ( .A1(n14505), .A2(n14506), .ZN(n14507) );
  NAND2_X1 U16287 ( .A1(n14508), .A2(n14507), .ZN(n14509) );
  AOI222_X1 U16288 ( .A1(n14697), .A2(n14511), .B1(n14510), .B2(n14694), .C1(
        n14509), .C2(n14692), .ZN(n14513) );
  OAI211_X1 U16289 ( .C1(n14701), .C2(n14514), .A(n14513), .B(n14512), .ZN(
        P2_U3187) );
  INV_X1 U16290 ( .A(n14515), .ZN(n14516) );
  NAND2_X1 U16291 ( .A1(n14517), .A2(n14516), .ZN(n14518) );
  NAND2_X1 U16292 ( .A1(n14518), .A2(n14532), .ZN(n14521) );
  NAND3_X1 U16293 ( .A1(n14521), .A2(n14520), .A3(n14519), .ZN(n14529) );
  NAND2_X1 U16294 ( .A1(n14523), .A2(n14522), .ZN(n14527) );
  NAND2_X1 U16295 ( .A1(n14525), .A2(n14524), .ZN(n14526) );
  NAND2_X1 U16296 ( .A1(n14527), .A2(n14526), .ZN(n14695) );
  INV_X1 U16297 ( .A(n14695), .ZN(n14528) );
  AND2_X1 U16298 ( .A1(n14529), .A2(n14528), .ZN(n14551) );
  AOI222_X1 U16299 ( .A1(n14696), .A2(n14531), .B1(P2_REG2_REG_12__SCAN_IN), 
        .B2(n6388), .C1(n14808), .C2(n14530), .ZN(n14539) );
  XNOR2_X1 U16300 ( .A(n14533), .B(n14532), .ZN(n14554) );
  AOI21_X1 U16301 ( .B1(n14696), .B2(n14534), .A(n10035), .ZN(n14536) );
  NAND2_X1 U16302 ( .A1(n14536), .A2(n14535), .ZN(n14550) );
  INV_X1 U16303 ( .A(n14550), .ZN(n14537) );
  AOI22_X1 U16304 ( .A1(n14554), .A2(n14815), .B1(n14806), .B2(n14537), .ZN(
        n14538) );
  OAI211_X1 U16305 ( .C1(n6388), .C2(n14551), .A(n14539), .B(n14538), .ZN(
        P2_U3253) );
  OAI22_X1 U16306 ( .A1(n14541), .A2(n10035), .B1(n14540), .B2(n14841), .ZN(
        n14543) );
  AOI211_X1 U16307 ( .C1(n14845), .C2(n14544), .A(n14543), .B(n14542), .ZN(
        n14556) );
  AOI22_X1 U16308 ( .A1(n14852), .A2(n14556), .B1(n14781), .B2(n14850), .ZN(
        P2_U3514) );
  OAI21_X1 U16309 ( .B1(n14546), .B2(n14841), .A(n14545), .ZN(n14548) );
  AOI211_X1 U16310 ( .C1(n14549), .C2(n14845), .A(n14548), .B(n14547), .ZN(
        n14558) );
  AOI22_X1 U16311 ( .A1(n14852), .A2(n14558), .B1(n11187), .B2(n14850), .ZN(
        P2_U3512) );
  INV_X1 U16312 ( .A(n14696), .ZN(n14552) );
  OAI211_X1 U16313 ( .C1(n14552), .C2(n14841), .A(n14551), .B(n14550), .ZN(
        n14553) );
  AOI21_X1 U16314 ( .B1(n14845), .B2(n14554), .A(n14553), .ZN(n14560) );
  AOI22_X1 U16315 ( .A1(n14852), .A2(n14560), .B1(n10288), .B2(n14850), .ZN(
        P2_U3511) );
  INV_X1 U16316 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n14555) );
  AOI22_X1 U16317 ( .A1(n14848), .A2(n14556), .B1(n14555), .B2(n14846), .ZN(
        P2_U3475) );
  INV_X1 U16318 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n14557) );
  AOI22_X1 U16319 ( .A1(n14848), .A2(n14558), .B1(n14557), .B2(n14846), .ZN(
        P2_U3469) );
  INV_X1 U16320 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14559) );
  AOI22_X1 U16321 ( .A1(n14848), .A2(n14560), .B1(n14559), .B2(n14846), .ZN(
        P2_U3466) );
  AOI21_X1 U16322 ( .B1(n14562), .B2(n14653), .A(n14561), .ZN(n14565) );
  NAND2_X1 U16323 ( .A1(n14563), .A2(n14654), .ZN(n14564) );
  OAI211_X1 U16324 ( .C1(n14566), .C2(n14672), .A(n14565), .B(n14564), .ZN(
        n14567) );
  AOI21_X1 U16325 ( .B1(n14568), .B2(n14677), .A(n14567), .ZN(n14570) );
  AOI22_X1 U16326 ( .A1(n14687), .A2(n14570), .B1(n10460), .B2(n14685), .ZN(
        P1_U3541) );
  INV_X1 U16327 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14569) );
  AOI22_X1 U16328 ( .A1(n14679), .A2(n14570), .B1(n14569), .B2(n14678), .ZN(
        P1_U3498) );
  OAI222_X1 U16329 ( .A1(n14575), .A2(n14574), .B1(n14575), .B2(n14573), .C1(
        n14572), .C2(n14571), .ZN(SUB_1596_U69) );
  OAI21_X1 U16330 ( .B1(n14578), .B2(n14577), .A(n14576), .ZN(n14579) );
  XNOR2_X1 U16331 ( .A(n14579), .B(P2_ADDR_REG_12__SCAN_IN), .ZN(SUB_1596_U68)
         );
  OAI21_X1 U16332 ( .B1(n14581), .B2(n14778), .A(n14580), .ZN(SUB_1596_U67) );
  OAI21_X1 U16333 ( .B1(n14584), .B2(n14583), .A(n14582), .ZN(n14585) );
  XNOR2_X1 U16334 ( .A(n14585), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  OAI21_X1 U16335 ( .B1(n14588), .B2(n14587), .A(n14586), .ZN(n14589) );
  XOR2_X1 U16336 ( .A(n14589), .B(n6978), .Z(SUB_1596_U65) );
  INV_X1 U16337 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n15241) );
  AOI21_X1 U16338 ( .B1(n14591), .B2(n14590), .A(n6515), .ZN(n14592) );
  XNOR2_X1 U16339 ( .A(n15241), .B(n14592), .ZN(SUB_1596_U64) );
  OAI21_X1 U16340 ( .B1(n14595), .B2(n14594), .A(n14593), .ZN(n14603) );
  AOI21_X1 U16341 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14597), .A(n14596), 
        .ZN(n14601) );
  OAI22_X1 U16342 ( .A1(n14601), .A2(n14600), .B1(n14599), .B2(n14598), .ZN(
        n14602) );
  AOI21_X1 U16343 ( .B1(n14604), .B2(n14603), .A(n14602), .ZN(n14606) );
  OAI211_X1 U16344 ( .C1(n15239), .C2(n14607), .A(n14606), .B(n14605), .ZN(
        P1_U3258) );
  INV_X1 U16345 ( .A(n14623), .ZN(n14671) );
  INV_X1 U16346 ( .A(n14608), .ZN(n14611) );
  INV_X1 U16347 ( .A(n14609), .ZN(n14610) );
  OAI211_X1 U16348 ( .C1(n14671), .C2(n14611), .A(n14610), .B(n14613), .ZN(
        n14612) );
  OAI21_X1 U16349 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n14613), .A(n14612), 
        .ZN(n14636) );
  NAND2_X1 U16350 ( .A1(n14614), .A2(n14617), .ZN(n14615) );
  NAND2_X1 U16351 ( .A1(n14616), .A2(n14615), .ZN(n14673) );
  OR2_X1 U16352 ( .A1(n14618), .A2(n14617), .ZN(n14619) );
  NAND2_X1 U16353 ( .A1(n14620), .A2(n14619), .ZN(n14676) );
  NAND2_X1 U16354 ( .A1(n14676), .A2(n14621), .ZN(n14632) );
  NAND2_X1 U16355 ( .A1(n14623), .A2(n14622), .ZN(n14624) );
  NAND2_X1 U16356 ( .A1(n14624), .A2(n14654), .ZN(n14625) );
  OR2_X1 U16357 ( .A1(n14626), .A2(n14625), .ZN(n14669) );
  INV_X1 U16358 ( .A(n14627), .ZN(n14628) );
  NAND2_X1 U16359 ( .A1(n14669), .A2(n14628), .ZN(n14630) );
  NAND2_X1 U16360 ( .A1(n14630), .A2(n14629), .ZN(n14631) );
  OAI211_X1 U16361 ( .C1(n14673), .C2(n14633), .A(n14632), .B(n14631), .ZN(
        n14634) );
  INV_X1 U16362 ( .A(n14634), .ZN(n14635) );
  OAI211_X1 U16363 ( .C1(n14638), .C2(n14637), .A(n14636), .B(n14635), .ZN(
        P1_U3283) );
  AND2_X1 U16364 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15229), .ZN(P1_U3294) );
  AND2_X1 U16365 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15229), .ZN(P1_U3295) );
  AND2_X1 U16366 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15229), .ZN(P1_U3296) );
  AND2_X1 U16367 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15229), .ZN(P1_U3297) );
  AND2_X1 U16368 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15229), .ZN(P1_U3298) );
  AND2_X1 U16369 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15229), .ZN(P1_U3299) );
  AND2_X1 U16370 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15229), .ZN(P1_U3300) );
  AND2_X1 U16371 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15229), .ZN(P1_U3301) );
  AND2_X1 U16372 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15229), .ZN(P1_U3302) );
  AND2_X1 U16373 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15229), .ZN(P1_U3303) );
  AND2_X1 U16374 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15229), .ZN(P1_U3304) );
  AND2_X1 U16375 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15229), .ZN(P1_U3305) );
  AND2_X1 U16376 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15229), .ZN(P1_U3306) );
  AND2_X1 U16377 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15229), .ZN(P1_U3307) );
  AND2_X1 U16378 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15229), .ZN(P1_U3308) );
  AND2_X1 U16379 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15229), .ZN(P1_U3309) );
  AND2_X1 U16380 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15229), .ZN(P1_U3310) );
  AND2_X1 U16381 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15229), .ZN(P1_U3311) );
  AND2_X1 U16382 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15229), .ZN(P1_U3313) );
  AND2_X1 U16383 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15229), .ZN(P1_U3314) );
  AND2_X1 U16384 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15229), .ZN(P1_U3315) );
  AND2_X1 U16385 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15229), .ZN(P1_U3316) );
  AND2_X1 U16386 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15229), .ZN(P1_U3317) );
  AND2_X1 U16387 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15229), .ZN(P1_U3318) );
  AND2_X1 U16388 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15229), .ZN(P1_U3319) );
  INV_X1 U16389 ( .A(n15229), .ZN(n14639) );
  INV_X1 U16390 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n15189) );
  NOR2_X1 U16391 ( .A1(n14639), .A2(n15189), .ZN(P1_U3320) );
  AND2_X1 U16392 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15229), .ZN(P1_U3321) );
  AND2_X1 U16393 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15229), .ZN(P1_U3322) );
  AND2_X1 U16394 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15229), .ZN(P1_U3323) );
  OAI22_X1 U16395 ( .A1(n14641), .A2(n14662), .B1(n14640), .B2(n14670), .ZN(
        n14643) );
  AOI211_X1 U16396 ( .C1(n14645), .C2(n14644), .A(n14643), .B(n14642), .ZN(
        n14680) );
  AOI22_X1 U16397 ( .A1(n14679), .A2(n14680), .B1(n9046), .B2(n14678), .ZN(
        P1_U3465) );
  OAI22_X1 U16398 ( .A1(n14647), .A2(n14662), .B1(n14646), .B2(n14670), .ZN(
        n14650) );
  INV_X1 U16399 ( .A(n14648), .ZN(n14649) );
  AOI211_X1 U16400 ( .C1(n14677), .C2(n14651), .A(n14650), .B(n14649), .ZN(
        n14682) );
  AOI22_X1 U16401 ( .A1(n14679), .A2(n14682), .B1(n9073), .B2(n14678), .ZN(
        P1_U3471) );
  AOI22_X1 U16402 ( .A1(n14655), .A2(n14654), .B1(n14653), .B2(n14652), .ZN(
        n14656) );
  OAI211_X1 U16403 ( .C1(n14659), .C2(n14658), .A(n14657), .B(n14656), .ZN(
        n14660) );
  INV_X1 U16404 ( .A(n14660), .ZN(n14683) );
  INV_X1 U16405 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n14661) );
  AOI22_X1 U16406 ( .A1(n14679), .A2(n14683), .B1(n14661), .B2(n14678), .ZN(
        P1_U3477) );
  OAI22_X1 U16407 ( .A1(n14663), .A2(n14662), .B1(n6810), .B2(n14670), .ZN(
        n14665) );
  AOI211_X1 U16408 ( .C1(n14677), .C2(n14666), .A(n14665), .B(n14664), .ZN(
        n14684) );
  INV_X1 U16409 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14667) );
  AOI22_X1 U16410 ( .A1(n14679), .A2(n14684), .B1(n14667), .B2(n14678), .ZN(
        P1_U3483) );
  OAI211_X1 U16411 ( .C1(n14671), .C2(n14670), .A(n14669), .B(n14668), .ZN(
        n14675) );
  NOR2_X1 U16412 ( .A1(n14673), .A2(n14672), .ZN(n14674) );
  AOI211_X1 U16413 ( .C1(n14677), .C2(n14676), .A(n14675), .B(n14674), .ZN(
        n14686) );
  AOI22_X1 U16414 ( .A1(n14679), .A2(n14686), .B1(n9156), .B2(n14678), .ZN(
        P1_U3489) );
  AOI22_X1 U16415 ( .A1(n14687), .A2(n14680), .B1(n9045), .B2(n14685), .ZN(
        P1_U3530) );
  INV_X1 U16416 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n14681) );
  AOI22_X1 U16417 ( .A1(n14687), .A2(n14682), .B1(n14681), .B2(n14685), .ZN(
        P1_U3532) );
  AOI22_X1 U16418 ( .A1(n14687), .A2(n14683), .B1(n9706), .B2(n14685), .ZN(
        P1_U3534) );
  AOI22_X1 U16419 ( .A1(n14687), .A2(n14684), .B1(n9710), .B2(n14685), .ZN(
        P1_U3536) );
  AOI22_X1 U16420 ( .A1(n14687), .A2(n14686), .B1(n9962), .B2(n14685), .ZN(
        P1_U3538) );
  NOR2_X1 U16421 ( .A1(n14719), .A2(P2_U3947), .ZN(P2_U3087) );
  NAND2_X1 U16422 ( .A1(n14689), .A2(n14688), .ZN(n14690) );
  XNOR2_X1 U16423 ( .A(n14691), .B(n14690), .ZN(n14693) );
  AOI222_X1 U16424 ( .A1(n14697), .A2(n14696), .B1(n14695), .B2(n14694), .C1(
        n14693), .C2(n14692), .ZN(n14699) );
  OAI211_X1 U16425 ( .C1(n14701), .C2(n14700), .A(n14699), .B(n14698), .ZN(
        P2_U3196) );
  INV_X1 U16426 ( .A(n14702), .ZN(n14704) );
  OAI21_X1 U16427 ( .B1(n14704), .B2(n14703), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n14705) );
  OAI21_X1 U16428 ( .B1(P2_STATE_REG_SCAN_IN), .B2(P2_REG3_REG_1__SCAN_IN), 
        .A(n14705), .ZN(n14718) );
  OAI211_X1 U16429 ( .C1(n14708), .C2(n14707), .A(n14770), .B(n14706), .ZN(
        n14709) );
  INV_X1 U16430 ( .A(n14709), .ZN(n14716) );
  NAND2_X1 U16431 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n14714) );
  INV_X1 U16432 ( .A(n14710), .ZN(n14713) );
  INV_X1 U16433 ( .A(n14711), .ZN(n14712) );
  AOI211_X1 U16434 ( .C1(n14714), .C2(n14713), .A(n14712), .B(n14791), .ZN(
        n14715) );
  AOI211_X1 U16435 ( .C1(n14719), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n14716), .B(
        n14715), .ZN(n14717) );
  NAND2_X1 U16436 ( .A1(n14718), .A2(n14717), .ZN(P2_U3215) );
  AOI22_X1 U16437 ( .A1(n14719), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n14732) );
  OAI21_X1 U16438 ( .B1(n14722), .B2(n14721), .A(n14720), .ZN(n14729) );
  OAI211_X1 U16439 ( .C1(n14725), .C2(n14724), .A(n14770), .B(n14723), .ZN(
        n14728) );
  NAND2_X1 U16440 ( .A1(n14802), .A2(n14726), .ZN(n14727) );
  OAI211_X1 U16441 ( .C1(n14791), .C2(n14729), .A(n14728), .B(n14727), .ZN(
        n14730) );
  INV_X1 U16442 ( .A(n14730), .ZN(n14731) );
  NAND2_X1 U16443 ( .A1(n14732), .A2(n14731), .ZN(P2_U3216) );
  OAI21_X1 U16444 ( .B1(n14735), .B2(n14734), .A(n14733), .ZN(n14742) );
  OAI211_X1 U16445 ( .C1(n14738), .C2(n14737), .A(n14770), .B(n14736), .ZN(
        n14741) );
  NAND2_X1 U16446 ( .A1(n14802), .A2(n14739), .ZN(n14740) );
  OAI211_X1 U16447 ( .C1(n14791), .C2(n14742), .A(n14741), .B(n14740), .ZN(
        n14743) );
  INV_X1 U16448 ( .A(n14743), .ZN(n14745) );
  NAND2_X1 U16449 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n14744) );
  OAI211_X1 U16450 ( .C1(n14805), .C2(n14746), .A(n14745), .B(n14744), .ZN(
        P2_U3218) );
  INV_X1 U16451 ( .A(n14747), .ZN(n14748) );
  OAI211_X1 U16452 ( .C1(n14750), .C2(n14749), .A(n14770), .B(n14748), .ZN(
        n14757) );
  NOR2_X1 U16453 ( .A1(n14752), .A2(n14751), .ZN(n14753) );
  NOR2_X1 U16454 ( .A1(n14754), .A2(n14753), .ZN(n14755) );
  NAND2_X1 U16455 ( .A1(n14765), .A2(n14755), .ZN(n14756) );
  OAI211_X1 U16456 ( .C1(n14774), .C2(n6617), .A(n14757), .B(n14756), .ZN(
        n14758) );
  INV_X1 U16457 ( .A(n14758), .ZN(n14760) );
  NAND2_X1 U16458 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n14759) );
  OAI211_X1 U16459 ( .C1(n14805), .C2(n15275), .A(n14760), .B(n14759), .ZN(
        P2_U3219) );
  AOI21_X1 U16460 ( .B1(n14763), .B2(n14762), .A(n14761), .ZN(n14764) );
  NAND2_X1 U16461 ( .A1(n14765), .A2(n14764), .ZN(n14772) );
  AOI21_X1 U16462 ( .B1(n14768), .B2(n14767), .A(n14766), .ZN(n14769) );
  NAND2_X1 U16463 ( .A1(n14770), .A2(n14769), .ZN(n14771) );
  OAI211_X1 U16464 ( .C1(n14774), .C2(n14773), .A(n14772), .B(n14771), .ZN(
        n14775) );
  INV_X1 U16465 ( .A(n14775), .ZN(n14777) );
  NAND2_X1 U16466 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n14776)
         );
  OAI211_X1 U16467 ( .C1(n14778), .C2(n14805), .A(n14777), .B(n14776), .ZN(
        P2_U3227) );
  INV_X1 U16468 ( .A(n14779), .ZN(n14788) );
  AOI211_X1 U16469 ( .C1(n14782), .C2(n14781), .A(n14780), .B(n14791), .ZN(
        n14787) );
  AOI211_X1 U16470 ( .C1(n14785), .C2(n14784), .A(n14783), .B(n14795), .ZN(
        n14786) );
  AOI211_X1 U16471 ( .C1(n14802), .C2(n14788), .A(n14787), .B(n14786), .ZN(
        n14790) );
  NAND2_X1 U16472 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3088), .ZN(n14789)
         );
  OAI211_X1 U16473 ( .C1(n6978), .C2(n14805), .A(n14790), .B(n14789), .ZN(
        P2_U3229) );
  AOI211_X1 U16474 ( .C1(n14794), .C2(n14793), .A(n14792), .B(n14791), .ZN(
        n14800) );
  AOI211_X1 U16475 ( .C1(n14798), .C2(n14797), .A(n14796), .B(n14795), .ZN(
        n14799) );
  AOI211_X1 U16476 ( .C1(n14802), .C2(n14801), .A(n14800), .B(n14799), .ZN(
        n14804) );
  OAI211_X1 U16477 ( .C1(n15241), .C2(n14805), .A(n14804), .B(n14803), .ZN(
        P2_U3230) );
  NAND2_X1 U16478 ( .A1(n14807), .A2(n14806), .ZN(n14811) );
  AOI22_X1 U16479 ( .A1(n14819), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n14809), 
        .B2(n14808), .ZN(n14810) );
  OAI211_X1 U16480 ( .C1(n14813), .C2(n14812), .A(n14811), .B(n14810), .ZN(
        n14814) );
  AOI21_X1 U16481 ( .B1(n14816), .B2(n14815), .A(n14814), .ZN(n14817) );
  OAI21_X1 U16482 ( .B1(n6388), .B2(n14818), .A(n14817), .ZN(P2_U3258) );
  INV_X1 U16483 ( .A(n14827), .ZN(n14824) );
  AND2_X1 U16484 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14821), .ZN(P2_U3266) );
  AND2_X1 U16485 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14821), .ZN(P2_U3267) );
  AND2_X1 U16486 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14821), .ZN(P2_U3268) );
  AND2_X1 U16487 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14821), .ZN(P2_U3269) );
  AND2_X1 U16488 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14821), .ZN(P2_U3270) );
  AND2_X1 U16489 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14821), .ZN(P2_U3271) );
  AND2_X1 U16490 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14821), .ZN(P2_U3272) );
  AND2_X1 U16491 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14821), .ZN(P2_U3273) );
  AND2_X1 U16492 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14821), .ZN(P2_U3274) );
  AND2_X1 U16493 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14821), .ZN(P2_U3275) );
  AND2_X1 U16494 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14821), .ZN(P2_U3276) );
  AND2_X1 U16495 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14821), .ZN(P2_U3277) );
  AND2_X1 U16496 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14821), .ZN(P2_U3278) );
  AND2_X1 U16497 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14821), .ZN(P2_U3279) );
  AND2_X1 U16498 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14821), .ZN(P2_U3280) );
  AND2_X1 U16499 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14821), .ZN(P2_U3281) );
  AND2_X1 U16500 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14821), .ZN(P2_U3282) );
  AND2_X1 U16501 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14821), .ZN(P2_U3283) );
  AND2_X1 U16502 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14821), .ZN(P2_U3284) );
  AND2_X1 U16503 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14821), .ZN(P2_U3285) );
  AND2_X1 U16504 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14821), .ZN(P2_U3286) );
  AND2_X1 U16505 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14821), .ZN(P2_U3287) );
  AND2_X1 U16506 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14821), .ZN(P2_U3288) );
  AND2_X1 U16507 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14821), .ZN(P2_U3289) );
  AND2_X1 U16508 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14821), .ZN(P2_U3290) );
  AND2_X1 U16509 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14821), .ZN(P2_U3291) );
  AND2_X1 U16510 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14821), .ZN(P2_U3292) );
  AND2_X1 U16511 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14821), .ZN(P2_U3293) );
  AND2_X1 U16512 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14821), .ZN(P2_U3294) );
  AND2_X1 U16513 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14821), .ZN(P2_U3295) );
  OAI21_X1 U16514 ( .B1(n14827), .B2(n14823), .A(n14822), .ZN(P2_U3416) );
  AOI22_X1 U16515 ( .A1(n14827), .A2(n14826), .B1(n14825), .B2(n14824), .ZN(
        P2_U3417) );
  INV_X1 U16516 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n14828) );
  AOI22_X1 U16517 ( .A1(n14848), .A2(n14829), .B1(n14828), .B2(n14846), .ZN(
        P2_U3430) );
  NAND2_X1 U16518 ( .A1(n14831), .A2(n14830), .ZN(n14832) );
  OAI211_X1 U16519 ( .C1(n14835), .C2(n14834), .A(n14833), .B(n14832), .ZN(
        n14836) );
  NOR2_X1 U16520 ( .A1(n14837), .A2(n14836), .ZN(n14849) );
  INV_X1 U16521 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n14838) );
  AOI22_X1 U16522 ( .A1(n14848), .A2(n14849), .B1(n14838), .B2(n14846), .ZN(
        P2_U3454) );
  OAI211_X1 U16523 ( .C1(n14842), .C2(n14841), .A(n14840), .B(n14839), .ZN(
        n14843) );
  AOI21_X1 U16524 ( .B1(n14845), .B2(n14844), .A(n14843), .ZN(n14851) );
  INV_X1 U16525 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n14847) );
  AOI22_X1 U16526 ( .A1(n14848), .A2(n14851), .B1(n14847), .B2(n14846), .ZN(
        P2_U3463) );
  AOI22_X1 U16527 ( .A1(n14852), .A2(n14849), .B1(n6632), .B2(n14850), .ZN(
        P2_U3507) );
  AOI22_X1 U16528 ( .A1(n14852), .A2(n14851), .B1(n10177), .B2(n14850), .ZN(
        P2_U3510) );
  NOR2_X1 U16529 ( .A1(P3_U3897), .A2(n14982), .ZN(P3_U3150) );
  AOI21_X1 U16530 ( .B1(n11488), .B2(n14854), .A(n14853), .ZN(n14871) );
  INV_X1 U16531 ( .A(n14855), .ZN(n14857) );
  NOR3_X1 U16532 ( .A1(n14858), .A2(n14857), .A3(n14856), .ZN(n14861) );
  INV_X1 U16533 ( .A(n14878), .ZN(n14860) );
  OAI21_X1 U16534 ( .B1(n14861), .B2(n14860), .A(n14859), .ZN(n14862) );
  OAI21_X1 U16535 ( .B1(n14977), .B2(n14863), .A(n14862), .ZN(n14864) );
  AOI211_X1 U16536 ( .C1(P3_ADDR_REG_3__SCAN_IN), .C2(n14982), .A(n14865), .B(
        n14864), .ZN(n14870) );
  OAI21_X1 U16537 ( .B1(P3_REG1_REG_3__SCAN_IN), .B2(n14867), .A(n14866), .ZN(
        n14868) );
  NAND2_X1 U16538 ( .A1(n14993), .A2(n14868), .ZN(n14869) );
  OAI211_X1 U16539 ( .C1(n14871), .C2(n15005), .A(n14870), .B(n14869), .ZN(
        P3_U3185) );
  AOI21_X1 U16540 ( .B1(n14873), .B2(n14872), .A(n6564), .ZN(n14890) );
  INV_X1 U16541 ( .A(n14874), .ZN(n14875) );
  NOR2_X1 U16542 ( .A1(n14876), .A2(n14875), .ZN(n14879) );
  INV_X1 U16543 ( .A(n14898), .ZN(n14877) );
  AOI21_X1 U16544 ( .B1(n14879), .B2(n14878), .A(n14877), .ZN(n14881) );
  OAI22_X1 U16545 ( .A1(n14881), .A2(n14999), .B1(n14880), .B2(n14977), .ZN(
        n14882) );
  AOI211_X1 U16546 ( .C1(P3_ADDR_REG_4__SCAN_IN), .C2(n14982), .A(n14883), .B(
        n14882), .ZN(n14889) );
  OAI21_X1 U16547 ( .B1(n14886), .B2(n14885), .A(n14884), .ZN(n14887) );
  NAND2_X1 U16548 ( .A1(n14993), .A2(n14887), .ZN(n14888) );
  OAI211_X1 U16549 ( .C1(n14890), .C2(n15005), .A(n14889), .B(n14888), .ZN(
        P3_U3186) );
  AOI21_X1 U16550 ( .B1(n14893), .B2(n14892), .A(n14891), .ZN(n14909) );
  INV_X1 U16551 ( .A(n14894), .ZN(n14895) );
  NOR2_X1 U16552 ( .A1(n14896), .A2(n14895), .ZN(n14899) );
  INV_X1 U16553 ( .A(n14917), .ZN(n14897) );
  AOI21_X1 U16554 ( .B1(n14899), .B2(n14898), .A(n14897), .ZN(n14901) );
  OAI22_X1 U16555 ( .A1(n14901), .A2(n14999), .B1(n14900), .B2(n14977), .ZN(
        n14902) );
  AOI211_X1 U16556 ( .C1(P3_ADDR_REG_5__SCAN_IN), .C2(n14982), .A(n14903), .B(
        n14902), .ZN(n14908) );
  OAI21_X1 U16557 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n14905), .A(n14904), .ZN(
        n14906) );
  NAND2_X1 U16558 ( .A1(n14993), .A2(n14906), .ZN(n14907) );
  OAI211_X1 U16559 ( .C1(n14909), .C2(n15005), .A(n14908), .B(n14907), .ZN(
        P3_U3187) );
  AOI21_X1 U16560 ( .B1(n14912), .B2(n14911), .A(n14910), .ZN(n14929) );
  INV_X1 U16561 ( .A(n14913), .ZN(n14914) );
  NOR2_X1 U16562 ( .A1(n14915), .A2(n14914), .ZN(n14918) );
  INV_X1 U16563 ( .A(n14937), .ZN(n14916) );
  AOI21_X1 U16564 ( .B1(n14918), .B2(n14917), .A(n14916), .ZN(n14920) );
  OAI22_X1 U16565 ( .A1(n14920), .A2(n14999), .B1(n14919), .B2(n14977), .ZN(
        n14921) );
  AOI211_X1 U16566 ( .C1(P3_ADDR_REG_6__SCAN_IN), .C2(n14982), .A(n14922), .B(
        n14921), .ZN(n14928) );
  OAI21_X1 U16567 ( .B1(n14925), .B2(n14924), .A(n14923), .ZN(n14926) );
  NAND2_X1 U16568 ( .A1(n14926), .A2(n14993), .ZN(n14927) );
  OAI211_X1 U16569 ( .C1(n14929), .C2(n15005), .A(n14928), .B(n14927), .ZN(
        P3_U3188) );
  AOI21_X1 U16570 ( .B1(n14932), .B2(n14931), .A(n14930), .ZN(n14948) );
  INV_X1 U16571 ( .A(n14933), .ZN(n14934) );
  NOR2_X1 U16572 ( .A1(n14935), .A2(n14934), .ZN(n14938) );
  INV_X1 U16573 ( .A(n14955), .ZN(n14936) );
  AOI21_X1 U16574 ( .B1(n14938), .B2(n14937), .A(n14936), .ZN(n14940) );
  OAI22_X1 U16575 ( .A1(n14940), .A2(n14999), .B1(n14939), .B2(n14977), .ZN(
        n14941) );
  AOI211_X1 U16576 ( .C1(P3_ADDR_REG_7__SCAN_IN), .C2(n14982), .A(n14942), .B(
        n14941), .ZN(n14947) );
  OAI21_X1 U16577 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n14944), .A(n14943), .ZN(
        n14945) );
  NAND2_X1 U16578 ( .A1(n14945), .A2(n14993), .ZN(n14946) );
  OAI211_X1 U16579 ( .C1(n14948), .C2(n15005), .A(n14947), .B(n14946), .ZN(
        P3_U3189) );
  AOI21_X1 U16580 ( .B1(n14950), .B2(n14949), .A(n6558), .ZN(n14967) );
  INV_X1 U16581 ( .A(n14951), .ZN(n14952) );
  NOR2_X1 U16582 ( .A1(n14953), .A2(n14952), .ZN(n14956) );
  INV_X1 U16583 ( .A(n14975), .ZN(n14954) );
  AOI21_X1 U16584 ( .B1(n14956), .B2(n14955), .A(n14954), .ZN(n14958) );
  OAI22_X1 U16585 ( .A1(n14958), .A2(n14999), .B1(n14957), .B2(n14977), .ZN(
        n14959) );
  AOI211_X1 U16586 ( .C1(P3_ADDR_REG_8__SCAN_IN), .C2(n14982), .A(n14960), .B(
        n14959), .ZN(n14966) );
  OAI21_X1 U16587 ( .B1(n14963), .B2(n14962), .A(n14961), .ZN(n14964) );
  NAND2_X1 U16588 ( .A1(n14964), .A2(n14993), .ZN(n14965) );
  OAI211_X1 U16589 ( .C1(n14967), .C2(n15005), .A(n14966), .B(n14965), .ZN(
        P3_U3190) );
  AOI21_X1 U16590 ( .B1(n14970), .B2(n14969), .A(n14968), .ZN(n14988) );
  INV_X1 U16591 ( .A(n14971), .ZN(n14972) );
  NOR2_X1 U16592 ( .A1(n14973), .A2(n14972), .ZN(n14976) );
  INV_X1 U16593 ( .A(n14998), .ZN(n14974) );
  AOI21_X1 U16594 ( .B1(n14976), .B2(n14975), .A(n14974), .ZN(n14979) );
  OAI22_X1 U16595 ( .A1(n14979), .A2(n14999), .B1(n14978), .B2(n14977), .ZN(
        n14980) );
  AOI211_X1 U16596 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n14982), .A(n14981), .B(
        n14980), .ZN(n14987) );
  OAI21_X1 U16597 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n14984), .A(n14983), .ZN(
        n14985) );
  NAND2_X1 U16598 ( .A1(n14985), .A2(n14993), .ZN(n14986) );
  OAI211_X1 U16599 ( .C1(n14988), .C2(n15005), .A(n14987), .B(n14986), .ZN(
        P3_U3191) );
  OAI21_X1 U16600 ( .B1(n14991), .B2(n14990), .A(n14989), .ZN(n14994) );
  AOI21_X1 U16601 ( .B1(n14994), .B2(n14993), .A(n14992), .ZN(n15012) );
  INV_X1 U16602 ( .A(n14995), .ZN(n14996) );
  NAND3_X1 U16603 ( .A1(n14998), .A2(n14997), .A3(n14996), .ZN(n15000) );
  AOI21_X1 U16604 ( .B1(n15001), .B2(n15000), .A(n14999), .ZN(n15008) );
  AOI21_X1 U16605 ( .B1(n15004), .B2(n15003), .A(n15002), .ZN(n15006) );
  NOR2_X1 U16606 ( .A1(n15006), .A2(n15005), .ZN(n15007) );
  AOI211_X1 U16607 ( .C1(n15010), .C2(n15009), .A(n15008), .B(n15007), .ZN(
        n15011) );
  OAI211_X1 U16608 ( .C1(n15014), .C2(n15013), .A(n15012), .B(n15011), .ZN(
        P3_U3192) );
  INV_X1 U16609 ( .A(n15015), .ZN(n15032) );
  OAI21_X1 U16610 ( .B1(n15032), .B2(n15017), .A(n15016), .ZN(n15020) );
  AOI222_X1 U16611 ( .A1(n15036), .A2(n15020), .B1(n15019), .B2(n10664), .C1(
        n15018), .C2(n15034), .ZN(n15021) );
  OAI21_X1 U16612 ( .B1(n15036), .B2(n15022), .A(n15021), .ZN(P3_U3225) );
  OAI21_X1 U16613 ( .B1(n15032), .B2(n15024), .A(n15023), .ZN(n15027) );
  AOI222_X1 U16614 ( .A1(n15036), .A2(n15027), .B1(n15026), .B2(n10664), .C1(
        n15025), .C2(n15034), .ZN(n15028) );
  OAI21_X1 U16615 ( .B1(n15036), .B2(n15029), .A(n15028), .ZN(P3_U3227) );
  OAI21_X1 U16616 ( .B1(n15032), .B2(n15031), .A(n15030), .ZN(n15037) );
  AOI222_X1 U16617 ( .A1(n15037), .A2(n15036), .B1(n15035), .B2(n15034), .C1(
        n15033), .C2(n10664), .ZN(n15038) );
  OAI21_X1 U16618 ( .B1(n15036), .B2(n15039), .A(n15038), .ZN(P3_U3229) );
  OR2_X1 U16619 ( .A1(n15041), .A2(n15040), .ZN(n15042) );
  NAND2_X1 U16620 ( .A1(n15043), .A2(n15042), .ZN(n15086) );
  OAI22_X1 U16621 ( .A1(n15047), .A2(n15046), .B1(n15045), .B2(n15044), .ZN(
        n15048) );
  AOI21_X1 U16622 ( .B1(n15086), .B2(n15106), .A(n15048), .ZN(n15054) );
  XNOR2_X1 U16623 ( .A(n15050), .B(n15049), .ZN(n15052) );
  NAND2_X1 U16624 ( .A1(n15052), .A2(n15051), .ZN(n15053) );
  NAND2_X1 U16625 ( .A1(n15054), .A2(n15053), .ZN(n15090) );
  INV_X1 U16626 ( .A(n15086), .ZN(n15058) );
  INV_X1 U16627 ( .A(n15076), .ZN(n15057) );
  NAND2_X1 U16628 ( .A1(n15055), .A2(n15073), .ZN(n15087) );
  OAI22_X1 U16629 ( .A1(n15058), .A2(n15057), .B1(n15056), .B2(n15087), .ZN(
        n15059) );
  AOI211_X1 U16630 ( .C1(n10664), .C2(P3_REG3_REG_2__SCAN_IN), .A(n15090), .B(
        n15059), .ZN(n15060) );
  AOI22_X1 U16631 ( .A1(n12826), .A2(n15061), .B1(n15060), .B2(n15036), .ZN(
        P3_U3231) );
  XNOR2_X1 U16632 ( .A(n15063), .B(n15062), .ZN(n15071) );
  XNOR2_X1 U16633 ( .A(n15064), .B(n15063), .ZN(n15084) );
  NAND2_X1 U16634 ( .A1(n15084), .A2(n15106), .ZN(n15070) );
  AOI22_X1 U16635 ( .A1(n15068), .A2(n15067), .B1(n15066), .B2(n15065), .ZN(
        n15069) );
  OAI211_X1 U16636 ( .C1(n15072), .C2(n15071), .A(n15070), .B(n15069), .ZN(
        n15082) );
  INV_X1 U16637 ( .A(n15082), .ZN(n15079) );
  AND2_X1 U16638 ( .A1(n15074), .A2(n15073), .ZN(n15083) );
  AOI22_X1 U16639 ( .A1(n10664), .A2(P3_REG3_REG_1__SCAN_IN), .B1(n15083), 
        .B2(n15075), .ZN(n15078) );
  NAND2_X1 U16640 ( .A1(n15084), .A2(n15076), .ZN(n15077) );
  AND3_X1 U16641 ( .A1(n15079), .A2(n15078), .A3(n15077), .ZN(n15080) );
  AOI22_X1 U16642 ( .A1(n12826), .A2(n15081), .B1(n15080), .B2(n15036), .ZN(
        P3_U3232) );
  INV_X1 U16643 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15085) );
  AOI211_X1 U16644 ( .C1(n15099), .C2(n15084), .A(n15083), .B(n15082), .ZN(
        n15111) );
  AOI22_X1 U16645 ( .A1(n15110), .A2(n15085), .B1(n15111), .B2(n15108), .ZN(
        P3_U3393) );
  NAND2_X1 U16646 ( .A1(n15086), .A2(n15099), .ZN(n15088) );
  NAND2_X1 U16647 ( .A1(n15088), .A2(n15087), .ZN(n15089) );
  NOR2_X1 U16648 ( .A1(n15090), .A2(n15089), .ZN(n15112) );
  INV_X1 U16649 ( .A(n15112), .ZN(n15091) );
  OAI22_X1 U16650 ( .A1(n15108), .A2(P3_REG0_REG_2__SCAN_IN), .B1(n15091), 
        .B2(n15110), .ZN(n15092) );
  INV_X1 U16651 ( .A(n15092), .ZN(P3_U3396) );
  INV_X1 U16652 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15098) );
  NAND2_X1 U16653 ( .A1(n15097), .A2(n15099), .ZN(n15093) );
  OAI211_X1 U16654 ( .C1(n15100), .C2(n15095), .A(n15094), .B(n15093), .ZN(
        n15096) );
  AOI21_X1 U16655 ( .B1(n15097), .B2(n15106), .A(n15096), .ZN(n15113) );
  AOI22_X1 U16656 ( .A1(n15110), .A2(n15098), .B1(n15113), .B2(n15108), .ZN(
        P3_U3417) );
  INV_X1 U16657 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15109) );
  INV_X1 U16658 ( .A(n15107), .ZN(n15103) );
  INV_X1 U16659 ( .A(n15099), .ZN(n15102) );
  OAI22_X1 U16660 ( .A1(n15103), .A2(n15102), .B1(n15101), .B2(n15100), .ZN(
        n15104) );
  AOI211_X1 U16661 ( .C1(n15107), .C2(n15106), .A(n15105), .B(n15104), .ZN(
        n15116) );
  AOI22_X1 U16662 ( .A1(n15110), .A2(n15109), .B1(n15116), .B2(n15108), .ZN(
        P3_U3420) );
  AOI22_X1 U16663 ( .A1(n15117), .A2(n15111), .B1(n10717), .B2(n15114), .ZN(
        P3_U3460) );
  AOI22_X1 U16664 ( .A1(n15117), .A2(n15112), .B1(n10713), .B2(n15114), .ZN(
        P3_U3461) );
  AOI22_X1 U16665 ( .A1(n15117), .A2(n15113), .B1(n11519), .B2(n15114), .ZN(
        P3_U3468) );
  AOI22_X1 U16666 ( .A1(n15117), .A2(n15116), .B1(n15115), .B2(n15114), .ZN(
        P3_U3469) );
  AOI22_X1 U16667 ( .A1(n15246), .A2(keyinput59), .B1(keyinput24), .B2(n9034), 
        .ZN(n15118) );
  OAI221_X1 U16668 ( .B1(n15246), .B2(keyinput59), .C1(n9034), .C2(keyinput24), 
        .A(n15118), .ZN(n15127) );
  AOI22_X1 U16669 ( .A1(n15239), .A2(keyinput58), .B1(n9329), .B2(keyinput51), 
        .ZN(n15119) );
  OAI221_X1 U16670 ( .B1(n15239), .B2(keyinput58), .C1(n9329), .C2(keyinput51), 
        .A(n15119), .ZN(n15126) );
  AOI22_X1 U16671 ( .A1(n15275), .A2(keyinput0), .B1(n15121), .B2(keyinput16), 
        .ZN(n15120) );
  OAI221_X1 U16672 ( .B1(n15275), .B2(keyinput0), .C1(n15121), .C2(keyinput16), 
        .A(n15120), .ZN(n15125) );
  AOI22_X1 U16673 ( .A1(n15241), .A2(keyinput48), .B1(n15123), .B2(keyinput41), 
        .ZN(n15122) );
  OAI221_X1 U16674 ( .B1(n15241), .B2(keyinput48), .C1(n15123), .C2(keyinput41), .A(n15122), .ZN(n15124) );
  NOR4_X1 U16675 ( .A1(n15127), .A2(n15126), .A3(n15125), .A4(n15124), .ZN(
        n15167) );
  AOI22_X1 U16676 ( .A1(n15243), .A2(keyinput4), .B1(keyinput3), .B2(n9710), 
        .ZN(n15128) );
  OAI221_X1 U16677 ( .B1(n15243), .B2(keyinput4), .C1(n9710), .C2(keyinput3), 
        .A(n15128), .ZN(n15137) );
  AOI22_X1 U16678 ( .A1(n15254), .A2(keyinput7), .B1(keyinput62), .B2(n15130), 
        .ZN(n15129) );
  OAI221_X1 U16679 ( .B1(n15254), .B2(keyinput7), .C1(n15130), .C2(keyinput62), 
        .A(n15129), .ZN(n15136) );
  XOR2_X1 U16680 ( .A(n10991), .B(keyinput29), .Z(n15134) );
  XNOR2_X1 U16681 ( .A(keyinput26), .B(P1_REG0_REG_1__SCAN_IN), .ZN(n15133) );
  XNOR2_X1 U16682 ( .A(P2_IR_REG_19__SCAN_IN), .B(keyinput27), .ZN(n15132) );
  XNOR2_X1 U16683 ( .A(P3_IR_REG_17__SCAN_IN), .B(keyinput40), .ZN(n15131) );
  NAND4_X1 U16684 ( .A1(n15134), .A2(n15133), .A3(n15132), .A4(n15131), .ZN(
        n15135) );
  NOR3_X1 U16685 ( .A1(n15137), .A2(n15136), .A3(n15135), .ZN(n15166) );
  INV_X1 U16686 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n15140) );
  INV_X1 U16687 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n15139) );
  AOI22_X1 U16688 ( .A1(n15140), .A2(keyinput38), .B1(n15139), .B2(keyinput43), 
        .ZN(n15138) );
  OAI221_X1 U16689 ( .B1(n15140), .B2(keyinput38), .C1(n15139), .C2(keyinput43), .A(n15138), .ZN(n15146) );
  XNOR2_X1 U16690 ( .A(n15141), .B(keyinput32), .ZN(n15145) );
  XNOR2_X1 U16691 ( .A(n15142), .B(keyinput23), .ZN(n15144) );
  XNOR2_X1 U16692 ( .A(n15256), .B(keyinput50), .ZN(n15143) );
  OR4_X1 U16693 ( .A1(n15146), .A2(n15145), .A3(n15144), .A4(n15143), .ZN(
        n15150) );
  AOI22_X1 U16694 ( .A1(n15247), .A2(keyinput18), .B1(keyinput35), .B2(n15238), 
        .ZN(n15147) );
  OAI221_X1 U16695 ( .B1(n15247), .B2(keyinput18), .C1(n15238), .C2(keyinput35), .A(n15147), .ZN(n15149) );
  XNOR2_X1 U16696 ( .A(n6802), .B(keyinput55), .ZN(n15148) );
  NOR3_X1 U16697 ( .A1(n15150), .A2(n15149), .A3(n15148), .ZN(n15165) );
  INV_X1 U16698 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n15153) );
  AOI22_X1 U16699 ( .A1(n15153), .A2(keyinput53), .B1(n15152), .B2(keyinput44), 
        .ZN(n15151) );
  OAI221_X1 U16700 ( .B1(n15153), .B2(keyinput53), .C1(n15152), .C2(keyinput44), .A(n15151), .ZN(n15163) );
  AOI22_X1 U16701 ( .A1(n11758), .A2(keyinput46), .B1(n15155), .B2(keyinput60), 
        .ZN(n15154) );
  OAI221_X1 U16702 ( .B1(n11758), .B2(keyinput46), .C1(n15155), .C2(keyinput60), .A(n15154), .ZN(n15162) );
  INV_X1 U16703 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n15157) );
  AOI22_X1 U16704 ( .A1(n15157), .A2(keyinput28), .B1(n15244), .B2(keyinput56), 
        .ZN(n15156) );
  OAI221_X1 U16705 ( .B1(n15157), .B2(keyinput28), .C1(n15244), .C2(keyinput56), .A(n15156), .ZN(n15161) );
  XNOR2_X1 U16706 ( .A(P3_REG1_REG_16__SCAN_IN), .B(keyinput6), .ZN(n15159) );
  XNOR2_X1 U16707 ( .A(P3_IR_REG_29__SCAN_IN), .B(keyinput22), .ZN(n15158) );
  NAND2_X1 U16708 ( .A1(n15159), .A2(n15158), .ZN(n15160) );
  NOR4_X1 U16709 ( .A1(n15163), .A2(n15162), .A3(n15161), .A4(n15160), .ZN(
        n15164) );
  NAND4_X1 U16710 ( .A1(n15167), .A2(n15166), .A3(n15165), .A4(n15164), .ZN(
        n15228) );
  AOI22_X1 U16711 ( .A1(n15169), .A2(keyinput10), .B1(keyinput39), .B2(n9187), 
        .ZN(n15168) );
  OAI221_X1 U16712 ( .B1(n15169), .B2(keyinput10), .C1(n9187), .C2(keyinput39), 
        .A(n15168), .ZN(n15172) );
  XNOR2_X1 U16713 ( .A(n15170), .B(keyinput57), .ZN(n15171) );
  NOR2_X1 U16714 ( .A1(n15172), .A2(n15171), .ZN(n15182) );
  AOI22_X1 U16715 ( .A1(n15255), .A2(keyinput20), .B1(keyinput36), .B2(n15174), 
        .ZN(n15173) );
  OAI221_X1 U16716 ( .B1(n15255), .B2(keyinput20), .C1(n15174), .C2(keyinput36), .A(n15173), .ZN(n15175) );
  INV_X1 U16717 ( .A(n15175), .ZN(n15181) );
  AOI22_X1 U16718 ( .A1(n15177), .A2(keyinput5), .B1(keyinput63), .B2(n12558), 
        .ZN(n15176) );
  OAI221_X1 U16719 ( .B1(n15177), .B2(keyinput5), .C1(n12558), .C2(keyinput63), 
        .A(n15176), .ZN(n15178) );
  INV_X1 U16720 ( .A(n15178), .ZN(n15180) );
  XNOR2_X1 U16721 ( .A(P3_IR_REG_11__SCAN_IN), .B(keyinput42), .ZN(n15179) );
  AND4_X1 U16722 ( .A1(n15182), .A2(n15181), .A3(n15180), .A4(n15179), .ZN(
        n15226) );
  AOI22_X1 U16723 ( .A1(n15184), .A2(keyinput33), .B1(n15240), .B2(keyinput1), 
        .ZN(n15183) );
  OAI221_X1 U16724 ( .B1(n15184), .B2(keyinput33), .C1(n15240), .C2(keyinput1), 
        .A(n15183), .ZN(n15196) );
  INV_X1 U16725 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n15187) );
  AOI22_X1 U16726 ( .A1(n15187), .A2(keyinput17), .B1(keyinput14), .B2(n15186), 
        .ZN(n15185) );
  OAI221_X1 U16727 ( .B1(n15187), .B2(keyinput17), .C1(n15186), .C2(keyinput14), .A(n15185), .ZN(n15195) );
  AOI22_X1 U16728 ( .A1(n15190), .A2(keyinput15), .B1(n15189), .B2(keyinput2), 
        .ZN(n15188) );
  OAI221_X1 U16729 ( .B1(n15190), .B2(keyinput15), .C1(n15189), .C2(keyinput2), 
        .A(n15188), .ZN(n15194) );
  XOR2_X1 U16730 ( .A(n12664), .B(keyinput30), .Z(n15192) );
  XNOR2_X1 U16731 ( .A(SI_6_), .B(keyinput49), .ZN(n15191) );
  NAND2_X1 U16732 ( .A1(n15192), .A2(n15191), .ZN(n15193) );
  NOR4_X1 U16733 ( .A1(n15196), .A2(n15195), .A3(n15194), .A4(n15193), .ZN(
        n15225) );
  AOI22_X1 U16734 ( .A1(n13409), .A2(keyinput45), .B1(keyinput54), .B2(n9342), 
        .ZN(n15197) );
  OAI221_X1 U16735 ( .B1(n13409), .B2(keyinput45), .C1(n9342), .C2(keyinput54), 
        .A(n15197), .ZN(n15208) );
  AOI22_X1 U16736 ( .A1(n15245), .A2(keyinput21), .B1(keyinput9), .B2(n15199), 
        .ZN(n15198) );
  OAI221_X1 U16737 ( .B1(n15245), .B2(keyinput21), .C1(n15199), .C2(keyinput9), 
        .A(n15198), .ZN(n15207) );
  AOI22_X1 U16738 ( .A1(n15201), .A2(keyinput31), .B1(keyinput19), .B2(n13304), 
        .ZN(n15200) );
  OAI221_X1 U16739 ( .B1(n15201), .B2(keyinput31), .C1(n13304), .C2(keyinput19), .A(n15200), .ZN(n15206) );
  XOR2_X1 U16740 ( .A(n15202), .B(keyinput37), .Z(n15204) );
  XNOR2_X1 U16741 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(keyinput34), .ZN(n15203)
         );
  NAND2_X1 U16742 ( .A1(n15204), .A2(n15203), .ZN(n15205) );
  NOR4_X1 U16743 ( .A1(n15208), .A2(n15207), .A3(n15206), .A4(n15205), .ZN(
        n15224) );
  INV_X1 U16744 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n15210) );
  AOI22_X1 U16745 ( .A1(n15210), .A2(keyinput12), .B1(keyinput13), .B2(n15242), 
        .ZN(n15209) );
  OAI221_X1 U16746 ( .B1(n15210), .B2(keyinput12), .C1(n15242), .C2(keyinput13), .A(n15209), .ZN(n15215) );
  XNOR2_X1 U16747 ( .A(n15211), .B(keyinput11), .ZN(n15214) );
  XNOR2_X1 U16748 ( .A(n15212), .B(keyinput8), .ZN(n15213) );
  OR3_X1 U16749 ( .A1(n15215), .A2(n15214), .A3(n15213), .ZN(n15222) );
  AOI22_X1 U16750 ( .A1(P1_U3086), .A2(keyinput61), .B1(keyinput25), .B2(
        n15217), .ZN(n15216) );
  OAI221_X1 U16751 ( .B1(P1_U3086), .B2(keyinput61), .C1(n15217), .C2(
        keyinput25), .A(n15216), .ZN(n15221) );
  INV_X1 U16752 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n15219) );
  AOI22_X1 U16753 ( .A1(n15232), .A2(keyinput52), .B1(n15219), .B2(keyinput47), 
        .ZN(n15218) );
  OAI221_X1 U16754 ( .B1(n15232), .B2(keyinput52), .C1(n15219), .C2(keyinput47), .A(n15218), .ZN(n15220) );
  NOR3_X1 U16755 ( .A1(n15222), .A2(n15221), .A3(n15220), .ZN(n15223) );
  NAND4_X1 U16756 ( .A1(n15226), .A2(n15225), .A3(n15224), .A4(n15223), .ZN(
        n15227) );
  NOR2_X1 U16757 ( .A1(n15228), .A2(n15227), .ZN(n15231) );
  NAND2_X1 U16758 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15229), .ZN(n15230) );
  XNOR2_X1 U16759 ( .A(n15231), .B(n15230), .ZN(n15270) );
  NOR3_X1 U16760 ( .A1(P3_REG3_REG_25__SCAN_IN), .A2(P3_DATAO_REG_24__SCAN_IN), 
        .A3(n15232), .ZN(n15235) );
  NOR4_X1 U16761 ( .A1(P3_D_REG_22__SCAN_IN), .A2(P3_IR_REG_29__SCAN_IN), .A3(
        P3_DATAO_REG_12__SCAN_IN), .A4(P3_DATAO_REG_17__SCAN_IN), .ZN(n15234)
         );
  NOR4_X1 U16762 ( .A1(P3_IR_REG_11__SCAN_IN), .A2(P2_REG0_REG_28__SCAN_IN), 
        .A3(P2_REG1_REG_24__SCAN_IN), .A4(P2_REG0_REG_29__SCAN_IN), .ZN(n15233) );
  NAND4_X1 U16763 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(n15235), .A3(n15234), .A4(
        n15233), .ZN(n15236) );
  NOR4_X1 U16764 ( .A1(n15237), .A2(n6802), .A3(n15275), .A4(n15236), .ZN(
        n15268) );
  AND4_X1 U16765 ( .A1(n9034), .A2(n15240), .A3(n15239), .A4(n15238), .ZN(
        n15252) );
  AND4_X1 U16766 ( .A1(n15244), .A2(n15243), .A3(n15242), .A4(n15241), .ZN(
        n15251) );
  NOR2_X1 U16767 ( .A1(SI_6_), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n15250) );
  NAND4_X1 U16768 ( .A1(n15247), .A2(n15246), .A3(n15245), .A4(n9035), .ZN(
        n15248) );
  NOR3_X1 U16769 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(P2_REG1_REG_21__SCAN_IN), 
        .A3(n15248), .ZN(n15249) );
  AND4_X1 U16770 ( .A1(n15252), .A2(n15251), .A3(n15250), .A4(n15249), .ZN(
        n15267) );
  NAND4_X1 U16771 ( .A1(n15254), .A2(n10991), .A3(n15253), .A4(n12558), .ZN(
        n15260) );
  NAND4_X1 U16772 ( .A1(P3_D_REG_5__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .A3(
        P2_REG0_REG_19__SCAN_IN), .A4(P1_REG2_REG_23__SCAN_IN), .ZN(n15259) );
  NAND4_X1 U16773 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_REG1_REG_21__SCAN_IN), 
        .A3(P1_REG0_REG_20__SCAN_IN), .A4(P1_REG0_REG_9__SCAN_IN), .ZN(n15258)
         );
  NAND4_X1 U16774 ( .A1(n15256), .A2(n15255), .A3(P3_REG3_REG_23__SCAN_IN), 
        .A4(P3_REG1_REG_4__SCAN_IN), .ZN(n15257) );
  NOR4_X1 U16775 ( .A1(n15260), .A2(n15259), .A3(n15258), .A4(n15257), .ZN(
        n15266) );
  NAND4_X1 U16776 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .A3(P3_ADDR_REG_11__SCAN_IN), .A4(P1_ADDR_REG_9__SCAN_IN), .ZN(n15264)
         );
  NAND4_X1 U16777 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(P1_REG2_REG_24__SCAN_IN), 
        .A3(P1_REG1_REG_12__SCAN_IN), .A4(P3_ADDR_REG_16__SCAN_IN), .ZN(n15263) );
  NAND4_X1 U16778 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_REG3_REG_17__SCAN_IN), 
        .A3(P2_DATAO_REG_31__SCAN_IN), .A4(P2_REG2_REG_25__SCAN_IN), .ZN(
        n15262) );
  NAND4_X1 U16779 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(P3_REG2_REG_24__SCAN_IN), 
        .A3(SI_30_), .A4(P2_ADDR_REG_18__SCAN_IN), .ZN(n15261) );
  NOR4_X1 U16780 ( .A1(n15264), .A2(n15263), .A3(n15262), .A4(n15261), .ZN(
        n15265) );
  NAND4_X1 U16781 ( .A1(n15268), .A2(n15267), .A3(n15266), .A4(n15265), .ZN(
        n15269) );
  XNOR2_X1 U16782 ( .A(n15270), .B(n15269), .ZN(P1_U3312) );
  AOI21_X1 U16783 ( .B1(n15273), .B2(n15272), .A(n15271), .ZN(SUB_1596_U59) );
  OAI21_X1 U16784 ( .B1(n15276), .B2(n15275), .A(n15274), .ZN(SUB_1596_U58) );
  XOR2_X1 U16785 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15277), .Z(SUB_1596_U53) );
  AOI21_X1 U16786 ( .B1(n15280), .B2(n15279), .A(n15278), .ZN(SUB_1596_U56) );
  AOI21_X1 U16787 ( .B1(n15283), .B2(n15282), .A(n15281), .ZN(n15284) );
  XOR2_X1 U16788 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15284), .Z(SUB_1596_U60) );
  AOI21_X1 U16789 ( .B1(n15287), .B2(n15286), .A(n15285), .ZN(SUB_1596_U5) );
  XNOR2_X1 U9673 ( .A(n8971), .B(P1_IR_REG_30__SCAN_IN), .ZN(n8975) );
  INV_X1 U7181 ( .A(n9842), .ZN(n6707) );
  CLKBUF_X2 U7139 ( .A(n9023), .Z(n9459) );
  CLKBUF_X3 U9816 ( .A(n9226), .Z(n9500) );
endmodule

