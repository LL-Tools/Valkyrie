

module b22_C_gen_AntiSAT_k_256_10 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, 
        keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, 
        keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, 
        keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, 
        keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, 
        keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, 
        keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, 
        keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, 
        keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104, 
        keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108, 
        keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112, 
        keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116, 
        keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120, 
        keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124, 
        keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, 
        keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, 
        keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, 
        keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, 
        keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, 
        keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, 
        keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, 
        keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, 
        SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, 
        SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, 
        SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, 
        SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, 
        P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, 
        P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, 
        P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, 
        P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, 
        P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, 
        P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, 
        P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, 
        P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, 
        P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, 
        P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, 
        P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, 
        P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, 
        P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, 
        P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, 
        P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, 
        P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, 
        P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, 
        P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, 
        P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, 
        P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, 
        P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, 
        P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, 
        P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, 
        P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, 
        P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, 
        P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, 
        P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, 
        P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, 
        P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, 
        P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, 
        P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, 
        P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, 
        P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, 
        P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, 
        P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, 
        P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, 
        P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, 
        P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, 
        P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, 
        P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, 
        P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, 
        P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, 
        P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, 
        P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, 
        P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, 
        P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, 
        P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, 
        P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0,
         keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5,
         keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10,
         keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15,
         keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20,
         keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25,
         keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30,
         keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35,
         keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40,
         keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45,
         keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50,
         keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55,
         keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60,
         keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65,
         keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70,
         keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75,
         keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80,
         keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85,
         keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90,
         keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95,
         keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100,
         keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104,
         keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108,
         keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112,
         keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116,
         keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120,
         keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124,
         keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1,
         keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6,
         keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11,
         keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16,
         keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21,
         keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26,
         keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31,
         keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36,
         keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41,
         keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46,
         keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51,
         keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56,
         keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61,
         keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66,
         keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71,
         keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76,
         keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81,
         keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86,
         keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91,
         keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96,
         keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100,
         keyinput_g101, keyinput_g102, keyinput_g103, keyinput_g104,
         keyinput_g105, keyinput_g106, keyinput_g107, keyinput_g108,
         keyinput_g109, keyinput_g110, keyinput_g111, keyinput_g112,
         keyinput_g113, keyinput_g114, keyinput_g115, keyinput_g116,
         keyinput_g117, keyinput_g118, keyinput_g119, keyinput_g120,
         keyinput_g121, keyinput_g122, keyinput_g123, keyinput_g124,
         keyinput_g125, keyinput_g126, keyinput_g127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755;

  INV_X4 U7419 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NAND3_X1 U7420 ( .A1(n6908), .A2(n6907), .A3(n6920), .ZN(n10147) );
  NAND2_X1 U7421 ( .A1(n7218), .A2(n7219), .ZN(n14279) );
  NAND2_X1 U7422 ( .A1(n8539), .A2(n8538), .ZN(n14343) );
  CLKBUF_X1 U7423 ( .A(n13747), .Z(n6684) );
  AOI21_X1 U7424 ( .B1(n13730), .B2(n9265), .A(n9212), .ZN(n13750) );
  NAND2_X2 U7425 ( .A1(n8184), .A2(n12685), .ZN(n14972) );
  INV_X1 U7426 ( .A(n6671), .ZN(n12780) );
  CLKBUF_X2 U7428 ( .A(n10244), .Z(n12882) );
  NAND2_X1 U7431 ( .A1(n6752), .A2(n8811), .ZN(n9273) );
  BUF_X1 U7433 ( .A(n10589), .Z(n13111) );
  INV_X2 U7434 ( .A(n9374), .ZN(n11159) );
  INV_X1 U7435 ( .A(n10243), .ZN(n8299) );
  OAI21_X1 U7436 ( .B1(n9420), .B2(n9421), .A(n6759), .ZN(n7118) );
  OR3_X2 U7437 ( .A1(n12572), .A2(n12123), .A3(n12387), .ZN(n10503) );
  NAND4_X1 U7438 ( .A1(n8318), .A2(n8317), .A3(n8316), .A4(n8315), .ZN(n14166)
         );
  INV_X1 U7439 ( .A(n7763), .ZN(n8115) );
  NAND4_X2 U7440 ( .A1(n8292), .A2(n8291), .A3(n8290), .A4(n8289), .ZN(n14169)
         );
  INV_X1 U7441 ( .A(n8464), .ZN(n8319) );
  INV_X2 U7442 ( .A(n8296), .ZN(n8325) );
  BUF_X2 U7443 ( .A(n7861), .Z(n12766) );
  INV_X1 U7445 ( .A(n7992), .ZN(n10203) );
  AND4_X1 U7446 ( .A1(n8284), .A2(n8283), .A3(n8282), .A4(n8281), .ZN(n10576)
         );
  BUF_X1 U7447 ( .A(n12579), .Z(n6682) );
  OAI21_X1 U7448 ( .B1(n12040), .B2(n8435), .A(n10072), .ZN(n12073) );
  NAND2_X2 U7449 ( .A1(n7328), .A2(n7329), .ZN(n14593) );
  NAND2_X1 U7450 ( .A1(n10503), .A2(n12577), .ZN(n13114) );
  XOR2_X1 U7451 ( .A(n11261), .B(n14660), .Z(n6671) );
  INV_X4 U7452 ( .A(n14397), .ZN(n6677) );
  INV_X2 U7454 ( .A(n12579), .ZN(n12764) );
  INV_X1 U7455 ( .A(n10589), .ZN(n13102) );
  INV_X1 U7456 ( .A(n11160), .ZN(n13173) );
  OR2_X1 U7457 ( .A1(n9031), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9051) );
  INV_X1 U7458 ( .A(n13112), .ZN(n13068) );
  INV_X2 U7459 ( .A(n6706), .ZN(n13115) );
  OR2_X1 U7460 ( .A1(n8623), .A2(n8622), .ZN(n8626) );
  INV_X1 U7461 ( .A(n9189), .ZN(n11521) );
  BUF_X1 U7462 ( .A(n8841), .Z(n9266) );
  INV_X1 U7463 ( .A(n8916), .ZN(n9189) );
  INV_X1 U7464 ( .A(n13178), .ZN(n15687) );
  NAND2_X1 U7465 ( .A1(n9059), .A2(n9058), .ZN(n9062) );
  OAI21_X1 U7466 ( .B1(n6758), .B2(n7449), .A(n7447), .ZN(n10129) );
  OR2_X1 U7467 ( .A1(n8696), .A2(n8637), .ZN(n8638) );
  OAI21_X1 U7468 ( .B1(n8516), .B2(n8515), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8517) );
  NAND2_X2 U7470 ( .A1(n7710), .A2(n7708), .ZN(n7744) );
  OR2_X1 U7471 ( .A1(n14810), .A2(n15004), .ZN(n14811) );
  AND2_X1 U7472 ( .A1(n14853), .A2(n14841), .ZN(n14839) );
  NAND2_X1 U7473 ( .A1(n8626), .A2(n8625), .ZN(n9846) );
  INV_X1 U7474 ( .A(n11252), .ZN(n13356) );
  INV_X1 U7475 ( .A(n8839), .ZN(n6679) );
  MUX2_X1 U7476 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n10187), .S(n15741), .Z(
        n10188) );
  CLKBUF_X1 U7477 ( .A(n10243), .Z(n10812) );
  NAND2_X1 U7478 ( .A1(n8741), .A2(n8713), .ZN(n14434) );
  NAND2_X1 U7479 ( .A1(n8541), .A2(n8540), .ZN(n14338) );
  NAND2_X1 U7480 ( .A1(n14523), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6891) );
  INV_X1 U7481 ( .A(n7779), .ZN(n12758) );
  NAND2_X1 U7482 ( .A1(n7965), .A2(n7964), .ZN(n14991) );
  OAI21_X1 U7483 ( .B1(n8221), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8220) );
  INV_X1 U7484 ( .A(n13724), .ZN(n13526) );
  AOI211_X1 U7485 ( .C1(n14428), .C2(n14366), .A(n14288), .B(n14287), .ZN(
        n14432) );
  NAND3_X1 U7486 ( .A1(n7506), .A2(n7505), .A3(n7175), .ZN(n6672) );
  NAND3_X1 U7487 ( .A1(n7506), .A2(n7505), .A3(n6928), .ZN(n6673) );
  OR2_X1 U7488 ( .A1(n10856), .A2(n10881), .ZN(n6674) );
  INV_X4 U7489 ( .A(n14398), .ZN(n12878) );
  XNOR2_X2 U7490 ( .A(n6891), .B(n6890), .ZN(n7310) );
  INV_X1 U7491 ( .A(n8296), .ZN(n6675) );
  NAND2_X1 U7492 ( .A1(n10535), .A2(n10046), .ZN(n8296) );
  XNOR2_X2 U7493 ( .A(n9385), .B(n9796), .ZN(n9428) );
  NOR2_X2 U7494 ( .A1(n13584), .A2(n13585), .ZN(n13604) );
  OAI21_X2 U7495 ( .B1(n9304), .B2(n7511), .A(n7509), .ZN(n13745) );
  AOI21_X2 U7496 ( .B1(n14685), .B2(n14684), .A(n14683), .ZN(n14682) );
  OR2_X2 U7497 ( .A1(n14434), .A2(n8697), .ZN(n9876) );
  INV_X1 U7498 ( .A(n14664), .ZN(n10603) );
  AND2_X2 U7499 ( .A1(n13379), .A2(n14046), .ZN(n8841) );
  XNOR2_X2 U7500 ( .A(n8786), .B(n8785), .ZN(n13379) );
  XNOR2_X2 U7501 ( .A(n9473), .B(n6851), .ZN(n9475) );
  XNOR2_X2 U7502 ( .A(n8798), .B(n8797), .ZN(n13354) );
  OAI21_X2 U7503 ( .B1(n9337), .B2(n7520), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n7372) );
  AOI21_X2 U7504 ( .B1(n13314), .B2(n13313), .A(n13342), .ZN(n13348) );
  XNOR2_X1 U7505 ( .A(n8659), .B(n11019), .ZN(n10999) );
  XNOR2_X2 U7506 ( .A(n12608), .B(n8165), .ZN(n12781) );
  NOR4_X2 U7507 ( .A1(n13342), .A2(n13341), .A3(n13340), .A4(n13339), .ZN(
        n13343) );
  XNOR2_X1 U7508 ( .A(n7739), .B(P1_IR_REG_2__SCAN_IN), .ZN(n14681) );
  XNOR2_X2 U7509 ( .A(n8151), .B(P1_IR_REG_22__SCAN_IN), .ZN(n15097) );
  OAI222_X1 U7510 ( .A1(n13377), .A2(n12969), .B1(P1_U3086), .B2(n12968), .C1(
        n13140), .C2(n13374), .ZN(P1_U3325) );
  XNOR2_X2 U7511 ( .A(n7700), .B(n12962), .ZN(n12968) );
  OAI21_X2 U7512 ( .B1(n9472), .B2(n15448), .A(n15247), .ZN(n15253) );
  INV_X2 U7513 ( .A(n8806), .ZN(n6676) );
  NAND2_X2 U7514 ( .A1(n7622), .A2(n7621), .ZN(n7624) );
  INV_X4 U7515 ( .A(n8806), .ZN(n10046) );
  NAND2_X2 U7516 ( .A1(n8383), .A2(n8382), .ZN(n11995) );
  AND2_X1 U7517 ( .A1(n7400), .A2(n15741), .ZN(n7371) );
  AOI21_X1 U7518 ( .B1(n14807), .B2(n6966), .A(n14806), .ZN(n15006) );
  NAND2_X1 U7519 ( .A1(n7405), .A2(n7404), .ZN(n13701) );
  NAND2_X1 U7520 ( .A1(n6692), .A2(n6753), .ZN(n7500) );
  OAI21_X1 U7521 ( .B1(n10147), .B2(n13288), .A(n10148), .ZN(n10175) );
  AOI21_X1 U7522 ( .B1(n10147), .B2(n10148), .A(n7363), .ZN(n13698) );
  NAND2_X1 U7523 ( .A1(n14260), .A2(n8595), .ZN(n14243) );
  AND2_X1 U7524 ( .A1(n9316), .A2(n9315), .ZN(n13700) );
  OR2_X1 U7525 ( .A1(n13288), .A2(n13292), .ZN(n13335) );
  MUX2_X1 U7526 ( .A(n14766), .B(n14765), .S(n14764), .Z(n14768) );
  INV_X1 U7527 ( .A(n13783), .ZN(n13784) );
  CLKBUF_X1 U7528 ( .A(n13795), .Z(n13825) );
  NAND2_X1 U7529 ( .A1(n9206), .A2(n9205), .ZN(n13427) );
  OR2_X1 U7530 ( .A1(n15126), .A2(n15127), .ZN(n13654) );
  AOI21_X1 U7531 ( .B1(n14892), .B2(n7528), .A(n7527), .ZN(n7526) );
  OR2_X1 U7532 ( .A1(n9180), .A2(n13760), .ZN(n13741) );
  XNOR2_X1 U7533 ( .A(n13766), .B(n13747), .ZN(n13760) );
  NAND2_X1 U7534 ( .A1(n9175), .A2(n9174), .ZN(n13766) );
  NAND2_X1 U7535 ( .A1(n8074), .A2(n8073), .ZN(n14883) );
  OAI21_X1 U7536 ( .B1(n7479), .B2(n6716), .A(n7480), .ZN(n9919) );
  OR2_X1 U7537 ( .A1(n8085), .A2(n8084), .ZN(n8088) );
  NAND2_X1 U7538 ( .A1(n6948), .A2(n13569), .ZN(n6947) );
  AND2_X1 U7539 ( .A1(n7312), .A2(n7311), .ZN(n12428) );
  XNOR2_X1 U7540 ( .A(n7047), .B(n14707), .ZN(n15259) );
  AND2_X1 U7541 ( .A1(n9412), .A2(n9413), .ZN(n9410) );
  NOR2_X1 U7542 ( .A1(n11759), .A2(n11760), .ZN(n14694) );
  AND2_X2 U7543 ( .A1(n12391), .A2(n13220), .ZN(n12392) );
  NAND2_X1 U7544 ( .A1(n7943), .A2(n7942), .ZN(n7959) );
  NAND2_X1 U7545 ( .A1(n7940), .A2(n7939), .ZN(n7943) );
  NAND2_X1 U7546 ( .A1(n7423), .A2(n6733), .ZN(n7940) );
  NAND2_X1 U7547 ( .A1(n7317), .A2(n7316), .ZN(n11350) );
  NAND2_X1 U7548 ( .A1(n6973), .A2(n8167), .ZN(n11478) );
  AND2_X1 U7549 ( .A1(n7011), .A2(n11641), .ZN(n7010) );
  NAND2_X1 U7550 ( .A1(n7833), .A2(n7832), .ZN(n12632) );
  INV_X1 U7551 ( .A(n12789), .ZN(n11625) );
  NOR2_X1 U7552 ( .A1(n9234), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9250) );
  OAI21_X1 U7553 ( .B1(n7860), .B2(n7859), .A(n7663), .ZN(n7875) );
  NAND2_X1 U7554 ( .A1(n7849), .A2(n7848), .ZN(n12641) );
  OR2_X1 U7555 ( .A1(n9221), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9234) );
  AOI21_X1 U7556 ( .B1(n12144), .B2(n11719), .A(n11718), .ZN(n11723) );
  XNOR2_X1 U7557 ( .A(n9022), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n9021) );
  NAND2_X2 U7558 ( .A1(n11366), .A2(n13914), .ZN(n15703) );
  NOR2_X1 U7559 ( .A1(n10602), .A2(n10601), .ZN(n10693) );
  OAI21_X1 U7560 ( .B1(n9437), .B2(n15109), .A(n15106), .ZN(n9438) );
  AND2_X1 U7561 ( .A1(n6960), .A2(n6959), .ZN(n11261) );
  INV_X1 U7562 ( .A(n10905), .ZN(n11464) );
  NAND2_X2 U7563 ( .A1(n14784), .A2(n14982), .ZN(n14913) );
  INV_X1 U7564 ( .A(n13535), .ZN(n15691) );
  NAND2_X1 U7565 ( .A1(n13535), .A2(n11173), .ZN(n13176) );
  NAND2_X1 U7566 ( .A1(n7376), .A2(n7374), .ZN(n8995) );
  INV_X2 U7567 ( .A(n13532), .ZN(n6678) );
  INV_X1 U7568 ( .A(n11578), .ZN(n11818) );
  NAND2_X1 U7569 ( .A1(n8822), .A2(n8821), .ZN(n15697) );
  NAND4_X1 U7570 ( .A1(n8805), .A2(n8804), .A3(n8803), .A4(n8802), .ZN(n13536)
         );
  NAND4_X1 U7571 ( .A1(n8304), .A2(n8303), .A3(n8302), .A4(n8301), .ZN(n14167)
         );
  OR2_X1 U7572 ( .A1(n15379), .A2(n15378), .ZN(n7096) );
  INV_X1 U7573 ( .A(n10590), .ZN(n15295) );
  OR2_X1 U7574 ( .A1(n6878), .A2(n6877), .ZN(n10590) );
  BUF_X2 U7575 ( .A(n8823), .Z(n8860) );
  AND2_X1 U7576 ( .A1(n7098), .A2(n7097), .ZN(n15379) );
  INV_X1 U7577 ( .A(n13114), .ZN(n10821) );
  BUF_X4 U7578 ( .A(n8312), .Z(n8582) );
  NAND2_X1 U7579 ( .A1(n7634), .A2(n7633), .ZN(n7752) );
  BUF_X2 U7580 ( .A(n8843), .Z(n9134) );
  BUF_X2 U7581 ( .A(n8310), .Z(n8405) );
  INV_X1 U7582 ( .A(n7723), .ZN(n7861) );
  CLKBUF_X3 U7583 ( .A(n13114), .Z(n6681) );
  AND2_X2 U7584 ( .A1(n10336), .A2(n11708), .ZN(n14398) );
  AND2_X1 U7585 ( .A1(n8270), .A2(n8269), .ZN(n8312) );
  INV_X1 U7586 ( .A(n10589), .ZN(n6680) );
  NAND2_X1 U7587 ( .A1(n7710), .A2(n13376), .ZN(n7784) );
  BUF_X2 U7588 ( .A(n8650), .Z(n11007) );
  AOI21_X1 U7589 ( .B1(n7642), .B2(n7419), .A(n6756), .ZN(n7418) );
  INV_X2 U7590 ( .A(n10357), .ZN(n7986) );
  CLKBUF_X1 U7591 ( .A(n8464), .Z(n10056) );
  XNOR2_X1 U7592 ( .A(n8644), .B(n8643), .ZN(n8713) );
  CLKBUF_X1 U7593 ( .A(n8206), .Z(n12993) );
  OR2_X2 U7594 ( .A1(n12770), .A2(n8198), .ZN(n14958) );
  XNOR2_X1 U7595 ( .A(n8268), .B(P2_IR_REG_29__SCAN_IN), .ZN(n8269) );
  INV_X1 U7596 ( .A(n12968), .ZN(n7710) );
  NAND2_X1 U7597 ( .A1(n8267), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8268) );
  INV_X1 U7598 ( .A(n15275), .ZN(n14764) );
  NAND2_X1 U7599 ( .A1(n8649), .A2(n8648), .ZN(n8697) );
  AOI21_X1 U7600 ( .B1(n7390), .B2(n7069), .A(n7068), .ZN(n7067) );
  XNOR2_X1 U7601 ( .A(n7703), .B(n7702), .ZN(n13376) );
  INV_X2 U7602 ( .A(n14037), .ZN(n12850) );
  XNOR2_X1 U7603 ( .A(n7625), .B(SI_1_), .ZN(n7722) );
  NAND2_X1 U7604 ( .A1(n12961), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7700) );
  AND2_X2 U7605 ( .A1(n7985), .A2(n8145), .ZN(n15275) );
  NAND2_X1 U7606 ( .A1(n7287), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7000) );
  NAND2_X1 U7607 ( .A1(n8727), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8277) );
  OAI21_X1 U7608 ( .B1(n8145), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8144) );
  AND2_X1 U7609 ( .A1(n7693), .A2(n7683), .ZN(n7692) );
  NAND2_X1 U7610 ( .A1(n8150), .A2(n7023), .ZN(n8145) );
  INV_X1 U7611 ( .A(n8717), .ZN(n8264) );
  NOR2_X1 U7612 ( .A1(n7601), .A2(P3_IR_REG_24__SCAN_IN), .ZN(n7177) );
  AND4_X1 U7613 ( .A1(n7689), .A2(n7893), .A3(n9594), .A4(n9733), .ZN(n7690)
         );
  AND3_X1 U7614 ( .A1(n7685), .A2(n7684), .A3(n7682), .ZN(n7570) );
  AND2_X1 U7615 ( .A1(n8294), .A2(n7458), .ZN(n7457) );
  AND4_X1 U7616 ( .A1(n8964), .A2(n9026), .A3(n9009), .A4(n8761), .ZN(n7593)
         );
  INV_X1 U7617 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n14769) );
  INV_X1 U7618 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n7893) );
  NOR2_X1 U7619 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n7685) );
  NOR2_X1 U7620 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n7684) );
  NOR2_X1 U7621 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n7686) );
  INV_X4 U7622 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X2 U7623 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9733) );
  XOR2_X1 U7624 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), .Z(
        n9420) );
  NOR2_X1 U7625 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n8781) );
  NOR2_X2 U7626 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n7960) );
  INV_X4 U7627 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7524) );
  XNOR2_X1 U7628 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8816) );
  INV_X1 U7629 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n9026) );
  INV_X1 U7630 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n9009) );
  INV_X1 U7631 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n8219) );
  INV_X1 U7632 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n8222) );
  INV_X1 U7633 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8231) );
  NOR2_X1 U7634 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n7678) );
  INV_X1 U7635 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8780) );
  INV_X1 U7636 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8779) );
  AOI21_X1 U7637 ( .B1(n14215), .B2(n15520), .A(n9868), .ZN(n10164) );
  XNOR2_X1 U7638 ( .A(n9851), .B(n10094), .ZN(n14215) );
  NAND2_X2 U7640 ( .A1(n14632), .A2(n14631), .ZN(n14630) );
  NOR2_X2 U7641 ( .A1(n9118), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9132) );
  NAND4_X4 U7642 ( .A1(n7719), .A2(n7718), .A3(n7717), .A4(n7716), .ZN(n14663)
         );
  AND2_X1 U7643 ( .A1(n12968), .A2(n13376), .ZN(n7779) );
  XNOR2_X2 U7644 ( .A(n7742), .B(n12589), .ZN(n12587) );
  INV_X2 U7645 ( .A(n14662), .ZN(n7742) );
  XNOR2_X1 U7646 ( .A(n8220), .B(n8219), .ZN(n12572) );
  NOR2_X2 U7647 ( .A1(n9051), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9067) );
  XNOR2_X2 U7648 ( .A(n7720), .B(n7055), .ZN(n14672) );
  NOR2_X1 U7649 ( .A1(n9306), .A2(n13724), .ZN(n13288) );
  AND2_X2 U7650 ( .A1(n9227), .A2(n9226), .ZN(n13724) );
  MUX2_X1 U7651 ( .A(n8198), .B(n8213), .S(n12759), .Z(n12579) );
  XNOR2_X2 U7652 ( .A(n11199), .B(n11196), .ZN(n11337) );
  NAND2_X1 U7653 ( .A1(n6913), .A2(n6915), .ZN(n6911) );
  OR2_X1 U7654 ( .A1(n13960), .A2(n13449), .ZN(n13256) );
  OR2_X1 U7655 ( .A1(n14032), .A2(n13896), .ZN(n9289) );
  NAND2_X1 U7656 ( .A1(n9126), .A2(n9125), .ZN(n9127) );
  INV_X1 U7657 ( .A(n7076), .ZN(n7075) );
  OAI21_X1 U7658 ( .B1(n9061), .B2(n7077), .A(n9089), .ZN(n7076) );
  NAND2_X1 U7659 ( .A1(n10439), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8889) );
  OAI21_X1 U7660 ( .B1(n12312), .B2(n8675), .A(n8674), .ZN(n12375) );
  OR2_X1 U7661 ( .A1(n14991), .A2(n14648), .ZN(n8184) );
  NAND2_X1 U7662 ( .A1(n7427), .A2(n6704), .ZN(n7429) );
  INV_X1 U7663 ( .A(n7146), .ZN(n11952) );
  OAI21_X1 U7664 ( .B1(n11653), .B2(n11652), .A(n6757), .ZN(n7146) );
  INV_X1 U7665 ( .A(n9134), .ZN(n9265) );
  NAND2_X1 U7666 ( .A1(n8790), .A2(n14046), .ZN(n8823) );
  XNOR2_X1 U7667 ( .A(n8770), .B(P3_IR_REG_19__SCAN_IN), .ZN(n13666) );
  AOI21_X1 U7668 ( .B1(n9094), .B2(n7388), .A(n7387), .ZN(n7386) );
  INV_X1 U7669 ( .A(n9108), .ZN(n7387) );
  INV_X1 U7670 ( .A(n9091), .ZN(n7388) );
  INV_X1 U7671 ( .A(n9094), .ZN(n7389) );
  INV_X1 U7672 ( .A(n7694), .ZN(n7770) );
  NAND2_X1 U7673 ( .A1(n7190), .A2(n10590), .ZN(n7188) );
  OR2_X1 U7674 ( .A1(n7193), .A2(n12667), .ZN(n7192) );
  INV_X1 U7675 ( .A(n9992), .ZN(n7488) );
  OR2_X1 U7676 ( .A1(n15275), .A2(n15097), .ZN(n7185) );
  NOR2_X1 U7677 ( .A1(n9386), .A2(n9387), .ZN(n9388) );
  NAND2_X1 U7678 ( .A1(n8790), .A2(n8794), .ZN(n8843) );
  NAND2_X1 U7679 ( .A1(n13336), .A2(n7364), .ZN(n7363) );
  NAND2_X1 U7680 ( .A1(n13288), .A2(n10148), .ZN(n7364) );
  NOR2_X1 U7681 ( .A1(n7511), .A2(n6838), .ZN(n6837) );
  INV_X1 U7682 ( .A(n9312), .ZN(n6838) );
  NOR2_X1 U7683 ( .A1(n13786), .A2(n7495), .ZN(n7494) );
  INV_X1 U7684 ( .A(n7497), .ZN(n7495) );
  INV_X1 U7685 ( .A(n9283), .ZN(n7508) );
  NAND2_X1 U7686 ( .A1(n7062), .A2(n9006), .ZN(n9022) );
  NAND2_X1 U7687 ( .A1(n9004), .A2(n9003), .ZN(n7062) );
  AOI21_X1 U7688 ( .B1(n7067), .B2(n7391), .A(n7378), .ZN(n7064) );
  NAND2_X1 U7689 ( .A1(n10585), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8981) );
  NAND2_X1 U7690 ( .A1(n10455), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8923) );
  NOR2_X1 U7691 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n10943) );
  AOI21_X1 U7692 ( .B1(n10021), .B2(n7463), .A(n7461), .ZN(n7460) );
  AOI22_X1 U7693 ( .A1(n7450), .A2(n7455), .B1(n7451), .B2(n7453), .ZN(n7448)
         );
  NAND2_X1 U7694 ( .A1(n10067), .A2(n7454), .ZN(n7453) );
  INV_X1 U7695 ( .A(n7455), .ZN(n7454) );
  AND2_X1 U7696 ( .A1(n10032), .A2(n7456), .ZN(n7455) );
  INV_X1 U7697 ( .A(n7310), .ZN(n8270) );
  INV_X1 U7698 ( .A(n7309), .ZN(n6887) );
  NOR2_X1 U7699 ( .A1(n12409), .A2(n14475), .ZN(n6986) );
  OAI21_X1 U7700 ( .B1(n12103), .B2(n8423), .A(n7265), .ZN(n12040) );
  OR2_X1 U7701 ( .A1(n12257), .A2(n14159), .ZN(n7265) );
  INV_X1 U7702 ( .A(n11317), .ZN(n8349) );
  NOR2_X1 U7703 ( .A1(n14307), .A2(n14430), .ZN(n14289) );
  NAND2_X1 U7704 ( .A1(n6889), .A2(n7277), .ZN(n14392) );
  AOI21_X1 U7705 ( .B1(n7279), .B2(n7281), .A(n6736), .ZN(n7277) );
  NAND2_X1 U7706 ( .A1(n8678), .A2(n7279), .ZN(n6889) );
  NAND3_X1 U7707 ( .A1(n6701), .A2(n8264), .A3(n7288), .ZN(n7287) );
  INV_X1 U7708 ( .A(n8062), .ZN(n7568) );
  INV_X1 U7709 ( .A(n8183), .ZN(n6983) );
  OR2_X1 U7710 ( .A1(n15225), .A2(n12999), .ZN(n12669) );
  OR2_X1 U7711 ( .A1(n14664), .A2(n15274), .ZN(n12777) );
  INV_X1 U7712 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n7689) );
  NAND2_X1 U7713 ( .A1(n7427), .A2(n8106), .ZN(n8124) );
  XNOR2_X1 U7714 ( .A(n8086), .B(SI_24_), .ZN(n8085) );
  INV_X1 U7715 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n7962) );
  AOI21_X1 U7716 ( .B1(n7412), .B2(n7032), .A(n7031), .ZN(n7030) );
  INV_X1 U7717 ( .A(n7650), .ZN(n7032) );
  NAND2_X1 U7718 ( .A1(n7034), .A2(n7650), .ZN(n7817) );
  NAND2_X1 U7719 ( .A1(n7803), .A2(n7648), .ZN(n7034) );
  XNOR2_X1 U7720 ( .A(n7643), .B(SI_5_), .ZN(n7420) );
  AND2_X1 U7721 ( .A1(n12352), .A2(n12355), .ZN(n12353) );
  OR2_X1 U7722 ( .A1(n12983), .A2(n12982), .ZN(n12984) );
  AOI21_X1 U7723 ( .B1(n11954), .B2(n6689), .A(n7181), .ZN(n7179) );
  INV_X1 U7724 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8756) );
  NAND2_X1 U7725 ( .A1(n6921), .A2(n9213), .ZN(n6920) );
  NAND2_X1 U7726 ( .A1(n6910), .A2(n6912), .ZN(n6908) );
  AND4_X1 U7727 ( .A1(n9138), .A2(n9137), .A3(n9136), .A4(n9135), .ZN(n13789)
         );
  NAND2_X1 U7728 ( .A1(n13963), .A2(n13256), .ZN(n13816) );
  NOR2_X1 U7729 ( .A1(n13521), .A2(n13878), .ZN(n6839) );
  OR2_X1 U7730 ( .A1(n9327), .A2(n13267), .ZN(n15690) );
  AND2_X1 U7731 ( .A1(n7397), .A2(n7402), .ZN(n7399) );
  OR2_X1 U7732 ( .A1(n13689), .A2(n15726), .ZN(n7397) );
  CLKBUF_X1 U7733 ( .A(n8980), .Z(n13150) );
  INV_X1 U7734 ( .A(n13150), .ZN(n9115) );
  INV_X1 U7735 ( .A(n9145), .ZN(n13149) );
  NAND2_X1 U7736 ( .A1(n11252), .A2(n11160), .ZN(n15719) );
  AND2_X1 U7737 ( .A1(n14035), .A2(n11103), .ZN(n11118) );
  NAND2_X1 U7738 ( .A1(n9246), .A2(n9245), .ZN(n9257) );
  OR2_X1 U7739 ( .A1(n9244), .A2(n9243), .ZN(n9246) );
  XNOR2_X1 U7740 ( .A(n9335), .B(P3_IR_REG_26__SCAN_IN), .ZN(n9346) );
  NAND2_X1 U7741 ( .A1(n6708), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9335) );
  CLKBUF_X1 U7742 ( .A(n9337), .Z(n9338) );
  NAND2_X1 U7743 ( .A1(n9127), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9139) );
  AOI21_X1 U7744 ( .B1(n7386), .B2(n7389), .A(n7385), .ZN(n7384) );
  INV_X1 U7745 ( .A(n9111), .ZN(n7385) );
  AND2_X1 U7746 ( .A1(n7593), .A2(n7368), .ZN(n7367) );
  INV_X1 U7747 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n7368) );
  NAND2_X1 U7748 ( .A1(n7394), .A2(n6804), .ZN(n9059) );
  INV_X1 U7749 ( .A(n9044), .ZN(n7396) );
  NAND2_X1 U7750 ( .A1(n8903), .A2(n6714), .ZN(n8924) );
  NAND2_X1 U7751 ( .A1(n8890), .A2(n8889), .ZN(n8901) );
  AND2_X1 U7752 ( .A1(n14051), .A2(n6797), .ZN(n7257) );
  NAND2_X1 U7753 ( .A1(n10234), .A2(n7213), .ZN(n10244) );
  NAND2_X1 U7754 ( .A1(n14084), .A2(n14083), .ZN(n14082) );
  XNOR2_X1 U7755 ( .A(n10244), .B(n10753), .ZN(n10238) );
  NAND2_X1 U7756 ( .A1(n7310), .A2(n8269), .ZN(n8367) );
  INV_X1 U7757 ( .A(n8405), .ZN(n8572) );
  OR2_X1 U7758 ( .A1(n15366), .A2(n15365), .ZN(n7098) );
  NAND2_X1 U7759 ( .A1(n14281), .A2(n7266), .ZN(n14260) );
  AND2_X1 U7760 ( .A1(n14264), .A2(n8588), .ZN(n7266) );
  AOI21_X1 U7761 ( .B1(n7226), .B2(n14342), .A(n6723), .ZN(n7225) );
  OR2_X1 U7762 ( .A1(n14338), .A2(n14355), .ZN(n7229) );
  AND2_X1 U7763 ( .A1(n7229), .A2(n7228), .ZN(n7226) );
  NOR2_X1 U7764 ( .A1(n12317), .A2(n12321), .ZN(n12318) );
  OAI21_X1 U7765 ( .B1(n12042), .B2(n7301), .A(n7297), .ZN(n12312) );
  AOI21_X1 U7766 ( .B1(n7300), .B2(n7299), .A(n7298), .ZN(n7297) );
  INV_X1 U7767 ( .A(n8671), .ZN(n7299) );
  INV_X1 U7768 ( .A(n10071), .ZN(n7298) );
  NAND2_X1 U7769 ( .A1(n10535), .A2(n8806), .ZN(n8464) );
  INV_X1 U7770 ( .A(n7287), .ZN(n8275) );
  NAND2_X1 U7771 ( .A1(n7326), .A2(n7327), .ZN(n7325) );
  OAI21_X1 U7772 ( .B1(n13119), .B2(n7345), .A(n7344), .ZN(n7343) );
  NAND2_X1 U7773 ( .A1(n13119), .A2(n7348), .ZN(n7344) );
  NOR2_X1 U7774 ( .A1(n7346), .A2(n14533), .ZN(n7345) );
  NAND2_X1 U7775 ( .A1(n10357), .A2(n8806), .ZN(n7723) );
  NAND2_X1 U7776 ( .A1(n15213), .A2(n12444), .ZN(n12449) );
  OR2_X1 U7777 ( .A1(n7912), .A2(n7911), .ZN(n7933) );
  INV_X1 U7778 ( .A(n12538), .ZN(n7327) );
  NAND2_X1 U7779 ( .A1(n10357), .A2(n10046), .ZN(n7694) );
  NOR2_X1 U7780 ( .A1(n15194), .A2(n15193), .ZN(n13018) );
  NAND2_X1 U7781 ( .A1(n7059), .A2(n7058), .ZN(n7057) );
  NAND2_X1 U7782 ( .A1(n14681), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7058) );
  INV_X1 U7783 ( .A(n6870), .ZN(n6869) );
  OAI21_X1 U7784 ( .B1(n6871), .B2(n6687), .A(n8102), .ZN(n6870) );
  NAND2_X1 U7785 ( .A1(n6862), .A2(n6861), .ZN(n14908) );
  AOI21_X1 U7786 ( .B1(n6691), .B2(n6864), .A(n6747), .ZN(n6861) );
  AND2_X1 U7787 ( .A1(n15048), .A2(n14647), .ZN(n8015) );
  NAND2_X1 U7788 ( .A1(n12460), .A2(n6984), .ZN(n12551) );
  OR2_X1 U7789 ( .A1(n12234), .A2(n12999), .ZN(n7591) );
  NAND2_X1 U7790 ( .A1(n12768), .A2(n12767), .ZN(n14774) );
  XNOR2_X1 U7791 ( .A(n8623), .B(n8127), .ZN(n12474) );
  OR2_X1 U7792 ( .A1(n7877), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n7892) );
  NAND2_X1 U7793 ( .A1(n7113), .A2(n7112), .ZN(n9455) );
  NAND2_X1 U7794 ( .A1(n7114), .A2(n15436), .ZN(n7113) );
  NAND2_X1 U7795 ( .A1(n15113), .A2(n15114), .ZN(n7114) );
  OAI21_X1 U7796 ( .B1(n13676), .B2(n15583), .A(n6827), .ZN(n6826) );
  INV_X1 U7797 ( .A(n13680), .ZN(n6827) );
  NAND2_X1 U7798 ( .A1(n7498), .A2(n13874), .ZN(n7501) );
  INV_X1 U7799 ( .A(n13335), .ZN(n7504) );
  NAND2_X1 U7800 ( .A1(n7313), .A2(n7314), .ZN(n10601) );
  NAND3_X1 U7801 ( .A1(n10507), .A2(n10506), .A3(n6706), .ZN(n7314) );
  NAND2_X1 U7802 ( .A1(n10599), .A2(n10600), .ZN(n7313) );
  INV_X1 U7803 ( .A(n12808), .ZN(n10208) );
  NAND2_X1 U7804 ( .A1(n9936), .A2(n9938), .ZN(n7478) );
  NAND2_X1 U7805 ( .A1(n9947), .A2(n9949), .ZN(n7474) );
  NAND2_X1 U7806 ( .A1(n12690), .A2(n12689), .ZN(n6821) );
  NAND2_X1 U7807 ( .A1(n12703), .A2(n12705), .ZN(n7202) );
  NAND2_X1 U7808 ( .A1(n7471), .A2(n10010), .ZN(n7469) );
  NOR2_X1 U7809 ( .A1(n7471), .A2(n10010), .ZN(n7470) );
  NAND2_X1 U7810 ( .A1(n12727), .A2(n12725), .ZN(n7211) );
  OR2_X1 U7811 ( .A1(n14264), .A2(n6847), .ZN(n6846) );
  OR4_X1 U7812 ( .A1(n10088), .A2(n14391), .A3(n14365), .A4(n10087), .ZN(
        n10089) );
  AND2_X1 U7813 ( .A1(n10084), .A2(n6843), .ZN(n10085) );
  NAND2_X1 U7814 ( .A1(n13838), .A2(n13251), .ZN(n6906) );
  NAND2_X1 U7815 ( .A1(n7462), .A2(n10027), .ZN(n7461) );
  NAND2_X1 U7816 ( .A1(n7464), .A2(n7463), .ZN(n7462) );
  INV_X1 U7817 ( .A(n7282), .ZN(n7281) );
  NOR2_X1 U7818 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n8260) );
  AND3_X1 U7819 ( .A1(n6823), .A2(n8259), .A3(n8258), .ZN(n7276) );
  NOR2_X1 U7820 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n6823) );
  NOR2_X1 U7821 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n8258) );
  NAND2_X1 U7822 ( .A1(n12736), .A2(n12738), .ZN(n7209) );
  INV_X1 U7823 ( .A(n7786), .ZN(n7565) );
  NAND2_X1 U7824 ( .A1(n8088), .A2(n6734), .ZN(n7427) );
  INV_X1 U7825 ( .A(n8104), .ZN(n7428) );
  AND2_X1 U7826 ( .A1(n7439), .A2(n8006), .ZN(n7438) );
  NAND2_X1 U7827 ( .A1(n7440), .A2(n6713), .ZN(n7439) );
  NOR2_X1 U7828 ( .A1(n7420), .A2(n7757), .ZN(n7416) );
  INV_X1 U7829 ( .A(n7420), .ZN(n7642) );
  AOI21_X1 U7830 ( .B1(n7628), .B2(n7629), .A(n7627), .ZN(n7631) );
  INV_X1 U7831 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n9809) );
  INV_X1 U7832 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n9806) );
  OR2_X1 U7833 ( .A1(n12918), .A2(n13469), .ZN(n12921) );
  NOR2_X1 U7834 ( .A1(n6796), .A2(n7158), .ZN(n7157) );
  INV_X1 U7835 ( .A(n12912), .ZN(n7158) );
  AND2_X1 U7836 ( .A1(n13466), .A2(n12921), .ZN(n12919) );
  NAND2_X1 U7837 ( .A1(n7168), .A2(n7170), .ZN(n7167) );
  INV_X1 U7838 ( .A(n12353), .ZN(n7168) );
  NAND2_X1 U7839 ( .A1(n11160), .A2(n11159), .ZN(n11161) );
  NOR2_X1 U7840 ( .A1(n15579), .A2(n6824), .ZN(n11904) );
  NOR2_X1 U7841 ( .A1(n15578), .A2(n11856), .ZN(n6824) );
  OR2_X1 U7842 ( .A1(n13707), .A2(n10177), .ZN(n9316) );
  INV_X1 U7843 ( .A(n6913), .ZN(n6912) );
  OR2_X1 U7844 ( .A1(n13427), .A2(n13750), .ZN(n13290) );
  INV_X1 U7845 ( .A(n13269), .ZN(n6917) );
  OR2_X1 U7846 ( .A1(n13414), .A2(n13801), .ZN(n13737) );
  OR2_X1 U7847 ( .A1(n9295), .A2(n9294), .ZN(n9296) );
  INV_X1 U7848 ( .A(n6926), .ZN(n6925) );
  OR2_X1 U7849 ( .A1(n13911), .A2(n6925), .ZN(n6924) );
  AND2_X1 U7850 ( .A1(n9038), .A2(n13230), .ZN(n7365) );
  OAI21_X1 U7851 ( .B1(n7351), .B2(n6902), .A(n13217), .ZN(n6901) );
  INV_X1 U7852 ( .A(n13212), .ZN(n6902) );
  INV_X1 U7853 ( .A(n13216), .ZN(n6899) );
  INV_X1 U7854 ( .A(n7517), .ZN(n7516) );
  NAND2_X1 U7855 ( .A1(n7518), .A2(n13323), .ZN(n7517) );
  INV_X1 U7856 ( .A(n7519), .ZN(n7518) );
  AOI21_X1 U7857 ( .B1(n7352), .B2(n12023), .A(n7515), .ZN(n7351) );
  INV_X1 U7858 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8784) );
  OR2_X1 U7859 ( .A1(n9160), .A2(n12122), .ZN(n9202) );
  NOR2_X1 U7860 ( .A1(n8769), .A2(P3_IR_REG_19__SCAN_IN), .ZN(n8766) );
  OR2_X1 U7861 ( .A1(n8783), .A2(P3_IR_REG_18__SCAN_IN), .ZN(n8769) );
  INV_X1 U7862 ( .A(n9073), .ZN(n7077) );
  INV_X1 U7863 ( .A(n8944), .ZN(n7068) );
  INV_X1 U7864 ( .A(n7070), .ZN(n7069) );
  INV_X1 U7865 ( .A(n8923), .ZN(n7392) );
  INV_X1 U7866 ( .A(n8905), .ZN(n7393) );
  NAND2_X1 U7867 ( .A1(n7239), .A2(n7238), .ZN(n7043) );
  AND2_X1 U7868 ( .A1(n7242), .A2(n14090), .ZN(n7238) );
  AND2_X1 U7869 ( .A1(n10318), .A2(n14125), .ZN(n6828) );
  INV_X1 U7870 ( .A(n14105), .ZN(n7217) );
  INV_X1 U7871 ( .A(n14058), .ZN(n7216) );
  AND2_X1 U7872 ( .A1(n7241), .A2(n7240), .ZN(n7239) );
  INV_X1 U7873 ( .A(n12498), .ZN(n7240) );
  OR2_X1 U7874 ( .A1(n7243), .A2(n7242), .ZN(n7241) );
  AOI211_X1 U7875 ( .C1(n10111), .C2(n11007), .A(n10110), .B(n10109), .ZN(
        n10132) );
  AND2_X1 U7876 ( .A1(n15471), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7104) );
  INV_X1 U7877 ( .A(n6888), .ZN(n6886) );
  AND2_X1 U7878 ( .A1(n6727), .A2(n8690), .ZN(n7309) );
  AND2_X1 U7879 ( .A1(n10090), .A2(n8688), .ZN(n6888) );
  INV_X1 U7880 ( .A(n14365), .ZN(n7295) );
  NOR2_X1 U7881 ( .A1(n11782), .A2(n15533), .ZN(n11783) );
  NAND2_X1 U7882 ( .A1(n14347), .A2(n6731), .ZN(n14307) );
  AND2_X1 U7883 ( .A1(n8263), .A2(n7286), .ZN(n7285) );
  AND2_X1 U7884 ( .A1(n8266), .A2(n8265), .ZN(n7286) );
  INV_X1 U7885 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8266) );
  AND3_X1 U7886 ( .A1(n6993), .A2(n6992), .A3(n6991), .ZN(n8263) );
  INV_X1 U7887 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6993) );
  INV_X1 U7888 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8642) );
  NOR2_X1 U7889 ( .A1(n7048), .A2(n14694), .ZN(n7047) );
  NOR2_X1 U7890 ( .A1(n14695), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7048) );
  NAND2_X1 U7891 ( .A1(n7144), .A2(n14817), .ZN(n7143) );
  NAND2_X1 U7892 ( .A1(n6970), .A2(n6972), .ZN(n6969) );
  INV_X1 U7893 ( .A(n6971), .ZN(n6970) );
  OAI21_X1 U7894 ( .B1(n6972), .B2(n8190), .A(n7525), .ZN(n6971) );
  AOI21_X1 U7895 ( .B1(n7526), .B2(n12801), .A(n14866), .ZN(n7525) );
  NOR2_X1 U7896 ( .A1(n14941), .A2(n7579), .ZN(n7578) );
  INV_X1 U7897 ( .A(n8185), .ZN(n7540) );
  AND2_X1 U7898 ( .A1(n6766), .A2(n6981), .ZN(n6980) );
  NAND2_X1 U7899 ( .A1(n6982), .A2(n8183), .ZN(n6981) );
  INV_X1 U7900 ( .A(n6984), .ZN(n6982) );
  NOR2_X1 U7901 ( .A1(n12553), .A2(n6985), .ZN(n6984) );
  INV_X1 U7902 ( .A(n8181), .ZN(n6985) );
  NOR2_X1 U7903 ( .A1(n11625), .A2(n7559), .ZN(n7558) );
  NAND2_X1 U7904 ( .A1(n12789), .A2(n7562), .ZN(n7561) );
  INV_X1 U7905 ( .A(n7842), .ZN(n7562) );
  NOR2_X1 U7906 ( .A1(n12632), .A2(n12641), .ZN(n7140) );
  OAI21_X1 U7907 ( .B1(n11480), .B2(n12785), .A(n6859), .ZN(n11433) );
  AOI21_X1 U7908 ( .B1(n11599), .B2(n6860), .A(n6754), .ZN(n6859) );
  INV_X1 U7909 ( .A(n7815), .ZN(n6860) );
  INV_X1 U7910 ( .A(n8166), .ZN(n6975) );
  INV_X1 U7911 ( .A(n10771), .ZN(n12778) );
  NAND2_X1 U7912 ( .A1(n10928), .A2(n8164), .ZN(n6976) );
  NOR2_X1 U7913 ( .A1(n12770), .A2(n14764), .ZN(n10222) );
  AND2_X1 U7914 ( .A1(n7984), .A2(n7680), .ZN(n6978) );
  INV_X1 U7915 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n7680) );
  NAND2_X1 U7916 ( .A1(n8150), .A2(n6690), .ZN(n7982) );
  XNOR2_X1 U7917 ( .A(n8000), .B(SI_18_), .ZN(n7974) );
  NAND2_X1 U7918 ( .A1(n7037), .A2(n7035), .ZN(n7921) );
  AOI21_X1 U7919 ( .B1(n7039), .B2(n7041), .A(n7036), .ZN(n7035) );
  INV_X1 U7920 ( .A(n7040), .ZN(n7039) );
  AND2_X1 U7921 ( .A1(n7685), .A2(n7684), .ZN(n7571) );
  NAND2_X1 U7922 ( .A1(n7659), .A2(n7658), .ZN(n7860) );
  NAND2_X1 U7923 ( .A1(n7647), .A2(n7646), .ZN(n7803) );
  NAND2_X1 U7924 ( .A1(n7638), .A2(n7637), .ZN(n7758) );
  NOR2_X1 U7925 ( .A1(n9390), .A2(n9391), .ZN(n9392) );
  XNOR2_X1 U7926 ( .A(n9392), .B(n9393), .ZN(n9432) );
  OAI22_X2 U7927 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n9716), .B1(n9435), .B2(
        n9396), .ZN(n9397) );
  AOI22_X1 U7928 ( .A1(n15272), .A2(P3_ADDR_REG_15__SCAN_IN), .B1(n9468), .B2(
        n9470), .ZN(n9473) );
  INV_X1 U7929 ( .A(n12977), .ZN(n7151) );
  OR2_X1 U7930 ( .A1(n13393), .A2(n6684), .ZN(n13392) );
  AND2_X1 U7931 ( .A1(n12928), .A2(n13405), .ZN(n12929) );
  NOR2_X1 U7932 ( .A1(n13511), .A2(n13878), .ZN(n12905) );
  INV_X1 U7933 ( .A(n13842), .ZN(n13449) );
  AND2_X1 U7934 ( .A1(n12939), .A2(n12938), .ZN(n13455) );
  OR2_X1 U7935 ( .A1(n12937), .A2(n12936), .ZN(n12938) );
  NAND2_X1 U7936 ( .A1(n9151), .A2(n9150), .ZN(n9186) );
  NOR2_X1 U7937 ( .A1(n12507), .A2(n7171), .ZN(n7170) );
  INV_X1 U7938 ( .A(n7173), .ZN(n7172) );
  OR2_X1 U7939 ( .A1(n11950), .A2(n11949), .ZN(n11951) );
  NOR2_X1 U7940 ( .A1(n11953), .A2(n11954), .ZN(n12025) );
  NAND2_X1 U7941 ( .A1(n12949), .A2(n13430), .ZN(n13432) );
  INV_X1 U7942 ( .A(n13878), .ZN(n13510) );
  OR2_X1 U7943 ( .A1(n9370), .A2(n13702), .ZN(n13310) );
  NAND2_X1 U7944 ( .A1(n7357), .A2(n7355), .ZN(n13133) );
  NAND2_X1 U7945 ( .A1(n7360), .A2(n7356), .ZN(n7355) );
  NAND2_X1 U7946 ( .A1(n7361), .A2(n9213), .ZN(n7356) );
  NAND2_X1 U7947 ( .A1(n13161), .A2(n13160), .ZN(n13162) );
  OAI21_X1 U7948 ( .B1(n10881), .B2(n11222), .A(n10862), .ZN(n10863) );
  INV_X1 U7949 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8757) );
  INV_X1 U7950 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n7523) );
  NAND2_X1 U7951 ( .A1(n15568), .A2(n6709), .ZN(n6953) );
  NAND2_X1 U7952 ( .A1(n6952), .A2(n6709), .ZN(n6951) );
  OR2_X1 U7953 ( .A1(n15609), .A2(n15608), .ZN(n6949) );
  AOI21_X1 U7954 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n15649), .A(n15642), .ZN(
        n11845) );
  NOR2_X1 U7955 ( .A1(n12260), .A2(n7269), .ZN(n12327) );
  AND2_X1 U7956 ( .A1(n12262), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7269) );
  AOI21_X1 U7957 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n13540), .A(n13537), .ZN(
        n13555) );
  INV_X1 U7958 ( .A(n7272), .ZN(n13603) );
  NAND2_X1 U7959 ( .A1(n9312), .A2(n7406), .ZN(n7405) );
  NAND2_X1 U7960 ( .A1(n13761), .A2(n6837), .ZN(n7404) );
  NAND2_X1 U7961 ( .A1(n10169), .A2(n9314), .ZN(n7406) );
  NAND2_X1 U7962 ( .A1(n9318), .A2(n9317), .ZN(n13705) );
  INV_X1 U7963 ( .A(n13701), .ZN(n9318) );
  OR2_X1 U7964 ( .A1(n12931), .A2(n13788), .ZN(n13757) );
  NAND2_X1 U7965 ( .A1(n13774), .A2(n9302), .ZN(n9304) );
  NAND2_X1 U7966 ( .A1(n12931), .A2(n9301), .ZN(n9302) );
  NAND2_X1 U7967 ( .A1(n9304), .A2(n6799), .ZN(n13761) );
  AOI21_X1 U7968 ( .B1(n7586), .B2(n9299), .A(n6807), .ZN(n7497) );
  NAND2_X1 U7969 ( .A1(n13272), .A2(n13273), .ZN(n13798) );
  AND4_X1 U7970 ( .A1(n9123), .A2(n9122), .A3(n9121), .A4(n9120), .ZN(n13827)
         );
  NAND2_X1 U7971 ( .A1(n13858), .A2(n13857), .ZN(n13856) );
  AND4_X1 U7972 ( .A1(n9072), .A2(n9071), .A3(n9070), .A4(n9069), .ZN(n13864)
         );
  NOR2_X1 U7973 ( .A1(n13236), .A2(n6927), .ZN(n6926) );
  INV_X1 U7974 ( .A(n13231), .ZN(n6927) );
  NAND2_X1 U7975 ( .A1(n13912), .A2(n13911), .ZN(n13910) );
  AND4_X1 U7976 ( .A1(n8993), .A2(n8992), .A3(n8991), .A4(n8990), .ZN(n13897)
         );
  NAND2_X1 U7977 ( .A1(n11824), .A2(n7588), .ZN(n12153) );
  AOI21_X1 U7978 ( .B1(n13317), .B2(n7354), .A(n7353), .ZN(n7352) );
  INV_X1 U7979 ( .A(n13202), .ZN(n7354) );
  INV_X1 U7980 ( .A(n13206), .ZN(n7353) );
  NAND2_X1 U7981 ( .A1(n7350), .A2(n7351), .ZN(n12156) );
  AND2_X1 U7982 ( .A1(n11691), .A2(n9284), .ZN(n12006) );
  CLKBUF_X1 U7983 ( .A(n11691), .Z(n11692) );
  NAND2_X1 U7984 ( .A1(n9327), .A2(n13305), .ZN(n15689) );
  AND2_X1 U7985 ( .A1(n11493), .A2(n9278), .ZN(n9277) );
  AND2_X1 U7986 ( .A1(n8820), .A2(n7610), .ZN(n8822) );
  INV_X1 U7987 ( .A(n15690), .ZN(n13880) );
  NAND2_X1 U7988 ( .A1(n9220), .A2(n9219), .ZN(n9306) );
  NAND2_X1 U7989 ( .A1(n9107), .A2(n9106), .ZN(n13963) );
  OR2_X1 U7990 ( .A1(n8980), .A2(n10392), .ZN(n8930) );
  NOR2_X1 U7991 ( .A1(n9378), .A2(n9377), .ZN(n11115) );
  INV_X1 U7992 ( .A(n15689), .ZN(n13877) );
  NAND2_X1 U7993 ( .A1(n13138), .A2(n13137), .ZN(n13148) );
  OR2_X1 U7994 ( .A1(n13136), .A2(n13135), .ZN(n13138) );
  NAND4_X1 U7995 ( .A1(n7506), .A2(n7505), .A3(n7177), .A4(n6929), .ZN(n8787)
         );
  AND2_X1 U7996 ( .A1(n6930), .A2(n8797), .ZN(n6929) );
  OAI21_X1 U7997 ( .B1(n9229), .B2(n9228), .A(n9230), .ZN(n9244) );
  NOR2_X1 U7998 ( .A1(n7601), .A2(P3_IR_REG_17__SCAN_IN), .ZN(n7175) );
  XNOR2_X1 U7999 ( .A(n9334), .B(n9333), .ZN(n10855) );
  OAI21_X1 U8000 ( .B1(n9332), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9334) );
  NAND2_X1 U8001 ( .A1(n8771), .A2(n8780), .ZN(n9332) );
  NAND2_X1 U8002 ( .A1(n7380), .A2(n7381), .ZN(n9157) );
  AOI21_X1 U8003 ( .B1(n9139), .B2(P2_DATAO_REG_20__SCAN_IN), .A(n7382), .ZN(
        n7381) );
  INV_X1 U8004 ( .A(n9142), .ZN(n7382) );
  OAI21_X1 U8005 ( .B1(n9127), .B2(P1_DATAO_REG_20__SCAN_IN), .A(n9139), .ZN(
        n9128) );
  OR2_X1 U8006 ( .A1(n9128), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9140) );
  OAI21_X1 U8007 ( .B1(n9062), .B2(n7077), .A(n7075), .ZN(n9092) );
  AND2_X1 U8008 ( .A1(n9108), .A2(n9093), .ZN(n9094) );
  AND2_X1 U8009 ( .A1(n9073), .A2(n9060), .ZN(n9061) );
  NAND2_X1 U8010 ( .A1(n9062), .A2(n9061), .ZN(n9074) );
  NAND2_X1 U8011 ( .A1(n7607), .A2(n7593), .ZN(n8762) );
  NAND2_X1 U8012 ( .A1(n7395), .A2(n6698), .ZN(n7394) );
  NAND2_X1 U8013 ( .A1(n9022), .A2(n10817), .ZN(n9023) );
  NAND2_X1 U8014 ( .A1(n9021), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7395) );
  NAND2_X1 U8015 ( .A1(n8997), .A2(n8996), .ZN(n9004) );
  NAND2_X1 U8016 ( .A1(n8995), .A2(n8994), .ZN(n8997) );
  INV_X1 U8017 ( .A(n8958), .ZN(n7379) );
  AND2_X1 U8018 ( .A1(n8981), .A2(n8960), .ZN(n8961) );
  AND2_X1 U8019 ( .A1(n8958), .A2(n8946), .ZN(n8947) );
  NAND2_X1 U8020 ( .A1(n8948), .A2(n8947), .ZN(n8959) );
  NAND2_X1 U8021 ( .A1(n7063), .A2(n7067), .ZN(n8948) );
  OR2_X1 U8022 ( .A1(n8901), .A2(n7391), .ZN(n7063) );
  NOR2_X1 U8023 ( .A1(n7392), .A2(n7071), .ZN(n7070) );
  INV_X1 U8024 ( .A(n8900), .ZN(n7071) );
  AND2_X1 U8025 ( .A1(n8944), .A2(n8925), .ZN(n8926) );
  NAND2_X1 U8026 ( .A1(n8924), .A2(n8923), .ZN(n8927) );
  NAND2_X1 U8027 ( .A1(n8901), .A2(n8900), .ZN(n8903) );
  AND2_X1 U8028 ( .A1(n8889), .A2(n8872), .ZN(n8887) );
  AOI21_X1 U8029 ( .B1(n12063), .B2(n10301), .A(n7587), .ZN(n12203) );
  NOR2_X1 U8030 ( .A1(n12861), .A2(n12860), .ZN(n12862) );
  XNOR2_X1 U8031 ( .A(n10905), .B(n10244), .ZN(n10246) );
  AND2_X1 U8032 ( .A1(n14167), .A2(n12878), .ZN(n10245) );
  NAND2_X1 U8033 ( .A1(n11748), .A2(n11747), .ZN(n7253) );
  XNOR2_X1 U8034 ( .A(n11019), .B(n12882), .ZN(n10256) );
  NAND2_X1 U8035 ( .A1(n10898), .A2(n10254), .ZN(n10899) );
  NAND2_X1 U8036 ( .A1(n10884), .A2(n7261), .ZN(n11232) );
  AND2_X1 U8037 ( .A1(n10267), .A2(n10263), .ZN(n7261) );
  NAND2_X1 U8038 ( .A1(n14082), .A2(n12873), .ZN(n14136) );
  AND2_X1 U8039 ( .A1(n10098), .A2(n10142), .ZN(n10534) );
  NAND2_X1 U8040 ( .A1(n10132), .A2(n10130), .ZN(n7431) );
  NAND2_X1 U8041 ( .A1(n6842), .A2(n10141), .ZN(n6841) );
  INV_X1 U8042 ( .A(n10100), .ZN(n6842) );
  NOR2_X1 U8043 ( .A1(n7450), .A2(n7451), .ZN(n7449) );
  AND2_X1 U8044 ( .A1(n10066), .A2(n7448), .ZN(n7447) );
  NAND2_X1 U8045 ( .A1(n15369), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7097) );
  OR2_X1 U8046 ( .A1(n11536), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7093) );
  AOI21_X1 U8047 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n12217), .A(n12210), .ZN(
        n12211) );
  NOR2_X1 U8048 ( .A1(n14190), .A2(n14191), .ZN(n14192) );
  INV_X1 U8049 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7024) );
  AND2_X1 U8050 ( .A1(n14270), .A2(n6994), .ZN(n14210) );
  NOR2_X1 U8051 ( .A1(n10063), .A2(n6995), .ZN(n6994) );
  INV_X1 U8052 ( .A(n6996), .ZN(n6995) );
  OAI21_X1 U8053 ( .B1(n8695), .B2(n7306), .A(n7304), .ZN(n7308) );
  AOI21_X1 U8054 ( .B1(n7307), .B2(n7305), .A(n6743), .ZN(n7304) );
  NAND2_X1 U8055 ( .A1(n14243), .A2(n8607), .ZN(n8609) );
  NAND2_X1 U8056 ( .A1(n8694), .A2(n14242), .ZN(n14253) );
  AOI21_X1 U8057 ( .B1(n7222), .B2(n7220), .A(n6699), .ZN(n7219) );
  NAND2_X1 U8058 ( .A1(n14333), .A2(n6888), .ZN(n14328) );
  AND2_X1 U8059 ( .A1(n8677), .A2(n6718), .ZN(n7284) );
  NAND2_X1 U8060 ( .A1(n7283), .A2(n6718), .ZN(n7282) );
  INV_X1 U8061 ( .A(n14153), .ZN(n14129) );
  OR2_X1 U8062 ( .A1(n12375), .A2(n8676), .ZN(n8678) );
  NAND2_X1 U8063 ( .A1(n12318), .A2(n6986), .ZN(n12564) );
  INV_X1 U8064 ( .A(n12370), .ZN(n7236) );
  NAND2_X1 U8065 ( .A1(n8454), .A2(n8453), .ZN(n12321) );
  NAND2_X1 U8066 ( .A1(n12078), .A2(n12246), .ZN(n12317) );
  NAND2_X1 U8067 ( .A1(n12104), .A2(n8670), .ZN(n12042) );
  NAND2_X1 U8068 ( .A1(n8412), .A2(n8411), .ZN(n12103) );
  NAND2_X1 U8069 ( .A1(n12106), .A2(n12105), .ZN(n12104) );
  NAND2_X1 U8070 ( .A1(n11775), .A2(n8669), .ZN(n12106) );
  INV_X1 U8071 ( .A(n14368), .ZN(n14323) );
  INV_X1 U8072 ( .A(n14369), .ZN(n14325) );
  NOR2_X1 U8073 ( .A1(n11380), .A2(n15523), .ZN(n11739) );
  AND2_X1 U8074 ( .A1(n10075), .A2(n10074), .ZN(n11269) );
  INV_X1 U8075 ( .A(n11318), .ZN(n7251) );
  NAND2_X1 U8076 ( .A1(n8654), .A2(n8653), .ZN(n10850) );
  INV_X1 U8077 ( .A(n10743), .ZN(n8286) );
  AND2_X1 U8078 ( .A1(n8697), .A2(n8713), .ZN(n10336) );
  XNOR2_X1 U8079 ( .A(n7213), .B(n10142), .ZN(n7212) );
  NAND2_X1 U8080 ( .A1(n10058), .A2(n10057), .ZN(n14202) );
  NAND2_X1 U8081 ( .A1(n8520), .A2(n8519), .ZN(n14375) );
  NAND2_X1 U8082 ( .A1(n8329), .A2(n8328), .ZN(n11074) );
  NAND2_X1 U8083 ( .A1(n8264), .A2(n6701), .ZN(n8727) );
  INV_X1 U8084 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8643) );
  NAND2_X1 U8085 ( .A1(n7262), .A2(n6710), .ZN(n8646) );
  AND2_X1 U8086 ( .A1(n8326), .A2(n7263), .ZN(n7262) );
  NOR2_X1 U8087 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n7263) );
  OAI21_X1 U8088 ( .B1(n14533), .B2(n7021), .A(n7020), .ZN(n7019) );
  NOR2_X1 U8089 ( .A1(n14621), .A2(n7349), .ZN(n7021) );
  NAND2_X1 U8090 ( .A1(n14533), .A2(n13099), .ZN(n7020) );
  NOR2_X1 U8091 ( .A1(n12428), .A2(n12427), .ZN(n15181) );
  NOR2_X1 U8092 ( .A1(n14558), .A2(n7006), .ZN(n7005) );
  INV_X1 U8093 ( .A(n13053), .ZN(n7006) );
  INV_X1 U8094 ( .A(n7336), .ZN(n7335) );
  OAI21_X1 U8095 ( .B1(n14604), .B2(n7337), .A(n14540), .ZN(n7336) );
  INV_X1 U8096 ( .A(n13064), .ZN(n7337) );
  AND2_X1 U8097 ( .A1(n12541), .A2(n6776), .ZN(n7326) );
  NOR2_X1 U8098 ( .A1(n7851), .A2(n10918), .ZN(n7867) );
  NAND2_X1 U8099 ( .A1(n15181), .A2(n15180), .ZN(n15210) );
  NOR2_X1 U8100 ( .A1(n11344), .A2(n7319), .ZN(n7318) );
  INV_X1 U8101 ( .A(n11338), .ZN(n7319) );
  NOR2_X1 U8102 ( .A1(n11344), .A2(n11196), .ZN(n7321) );
  INV_X1 U8103 ( .A(n11189), .ZN(n11191) );
  NAND2_X1 U8104 ( .A1(n15172), .A2(n13008), .ZN(n13015) );
  AND2_X1 U8105 ( .A1(n7536), .A2(n7534), .ZN(n8165) );
  NOR2_X1 U8106 ( .A1(n7535), .A2(n6732), .ZN(n7534) );
  INV_X1 U8107 ( .A(n7537), .ZN(n7536) );
  NOR2_X1 U8108 ( .A1(n10210), .A2(n10476), .ZN(n7535) );
  INV_X1 U8109 ( .A(n7691), .ZN(n7927) );
  NAND2_X1 U8110 ( .A1(n7054), .A2(n7053), .ZN(n7052) );
  NAND2_X1 U8111 ( .A1(n14733), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n7053) );
  INV_X1 U8112 ( .A(n14732), .ZN(n7054) );
  NAND2_X1 U8113 ( .A1(n7052), .A2(n14751), .ZN(n7051) );
  NAND2_X1 U8114 ( .A1(n8109), .A2(n8108), .ZN(n14622) );
  INV_X1 U8115 ( .A(n8082), .ZN(n7566) );
  NOR2_X1 U8116 ( .A1(n6744), .A2(n6872), .ZN(n6871) );
  NAND2_X1 U8117 ( .A1(n7996), .A2(n14597), .ZN(n7997) );
  OAI21_X1 U8118 ( .B1(n14970), .B2(n7973), .A(n8184), .ZN(n14957) );
  NAND2_X1 U8119 ( .A1(n14957), .A2(n14956), .ZN(n14955) );
  NOR2_X1 U8120 ( .A1(n12413), .A2(n7554), .ZN(n7553) );
  INV_X1 U8121 ( .A(n7591), .ZN(n7554) );
  OR2_X1 U8122 ( .A1(n13009), .A2(n14650), .ZN(n7556) );
  NOR2_X1 U8123 ( .A1(n7543), .A2(n12798), .ZN(n7542) );
  OR2_X1 U8124 ( .A1(n12175), .A2(n6873), .ZN(n12226) );
  INV_X1 U8125 ( .A(n6876), .ZN(n6873) );
  AND2_X1 U8126 ( .A1(n12177), .A2(n12178), .ZN(n12175) );
  INV_X1 U8127 ( .A(n8170), .ZN(n7529) );
  NAND2_X1 U8128 ( .A1(n8169), .A2(n7559), .ZN(n11429) );
  NAND2_X1 U8129 ( .A1(n11606), .A2(n7140), .ZN(n11804) );
  OR2_X1 U8130 ( .A1(n12632), .A2(n14655), .ZN(n7842) );
  NAND2_X1 U8131 ( .A1(n11433), .A2(n12788), .ZN(n11432) );
  OR2_X1 U8132 ( .A1(n12599), .A2(n14660), .ZN(n7768) );
  OR2_X1 U8133 ( .A1(n12593), .A2(n14661), .ZN(n7756) );
  INV_X1 U8134 ( .A(n14871), .ZN(n14975) );
  AND2_X1 U8135 ( .A1(n8156), .A2(n8155), .ZN(n11583) );
  AND3_X1 U8136 ( .A1(n14810), .A2(n8214), .A3(n15049), .ZN(n14821) );
  OAI21_X1 U8137 ( .B1(n9846), .B2(n7444), .A(n7442), .ZN(n10055) );
  AOI21_X1 U8138 ( .B1(n7445), .B2(n7443), .A(n6812), .ZN(n7442) );
  INV_X1 U8139 ( .A(n7445), .ZN(n7444) );
  AND2_X1 U8140 ( .A1(n7691), .A2(n7692), .ZN(n7699) );
  NOR2_X1 U8141 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n7548) );
  NAND2_X1 U8142 ( .A1(n8088), .A2(n8087), .ZN(n8105) );
  AND2_X1 U8143 ( .A1(n6690), .A2(n7984), .ZN(n7023) );
  INV_X1 U8144 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8146) );
  XNOR2_X1 U8145 ( .A(n7974), .B(n8001), .ZN(n11388) );
  XNOR2_X1 U8146 ( .A(n7758), .B(n7757), .ZN(n10423) );
  XOR2_X1 U8147 ( .A(P3_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n9419) );
  NAND2_X1 U8148 ( .A1(n9430), .A2(n9431), .ZN(n9434) );
  XNOR2_X1 U8149 ( .A(n9432), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n9433) );
  XNOR2_X1 U8150 ( .A(n9401), .B(P1_ADDR_REG_10__SCAN_IN), .ZN(n9414) );
  NAND2_X1 U8151 ( .A1(n15234), .A2(n7121), .ZN(n7123) );
  OAI21_X1 U8152 ( .B1(n15234), .B2(n7121), .A(n7125), .ZN(n7122) );
  NOR2_X1 U8153 ( .A1(n15248), .A2(n15249), .ZN(n9472) );
  INV_X1 U8154 ( .A(n7131), .ZN(n7130) );
  AND3_X1 U8155 ( .A1(n8912), .A2(n8911), .A3(n8910), .ZN(n12030) );
  NAND2_X1 U8156 ( .A1(n12354), .A2(n12353), .ZN(n12506) );
  AND3_X1 U8157 ( .A1(n8968), .A2(n8967), .A3(n8966), .ZN(n15730) );
  OR2_X1 U8158 ( .A1(n13150), .A2(SI_10_), .ZN(n8967) );
  AND3_X1 U8159 ( .A1(n8838), .A2(n8837), .A3(n8836), .ZN(n11287) );
  NAND2_X1 U8160 ( .A1(n11281), .A2(n7615), .ZN(n11572) );
  NAND2_X1 U8161 ( .A1(n9117), .A2(n9116), .ZN(n13817) );
  NAND2_X1 U8162 ( .A1(n9147), .A2(n9146), .ZN(n13414) );
  OR2_X1 U8163 ( .A1(n13150), .A2(n11099), .ZN(n9146) );
  OR2_X1 U8164 ( .A1(n11100), .A2(n9145), .ZN(n9147) );
  AND4_X1 U8165 ( .A1(n8883), .A2(n8882), .A3(n8881), .A4(n8880), .ZN(n12028)
         );
  INV_X1 U8166 ( .A(n8859), .ZN(n11696) );
  AND3_X1 U8167 ( .A1(n8858), .A2(n8857), .A3(n8856), .ZN(n11578) );
  INV_X1 U8168 ( .A(n13523), .ZN(n13492) );
  NAND2_X1 U8169 ( .A1(n9050), .A2(n9049), .ZN(n13521) );
  XNOR2_X1 U8170 ( .A(n11839), .B(n15599), .ZN(n15588) );
  XNOR2_X1 U8171 ( .A(n12327), .B(n12328), .ZN(n12261) );
  NAND2_X1 U8172 ( .A1(n6957), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n7268) );
  INV_X1 U8173 ( .A(n12261), .ZN(n6957) );
  OAI22_X1 U8174 ( .A1(n12261), .A2(n6958), .B1(n6719), .B2(n12330), .ZN(
        n13537) );
  OR2_X1 U8175 ( .A1(n12330), .A2(n12528), .ZN(n6958) );
  NAND2_X1 U8176 ( .A1(n13655), .A2(n6938), .ZN(n6937) );
  INV_X1 U8177 ( .A(n6943), .ZN(n6938) );
  OAI21_X1 U8178 ( .B1(n13654), .B2(n6943), .A(n6941), .ZN(n6940) );
  NAND2_X1 U8179 ( .A1(n6942), .A2(n13668), .ZN(n6941) );
  INV_X1 U8180 ( .A(n6944), .ZN(n6942) );
  INV_X1 U8181 ( .A(n9330), .ZN(n7402) );
  NAND2_X1 U8182 ( .A1(n9099), .A2(n9098), .ZN(n13960) );
  NAND2_X1 U8183 ( .A1(n11681), .A2(n11680), .ZN(n13919) );
  AND2_X1 U8184 ( .A1(n11118), .A2(n11117), .ZN(n15702) );
  OR2_X1 U8185 ( .A1(n11366), .A2(n11365), .ZN(n13913) );
  NOR2_X1 U8186 ( .A1(n7500), .A2(n15739), .ZN(n7499) );
  NAND2_X1 U8187 ( .A1(n7501), .A2(n15734), .ZN(n6932) );
  INV_X1 U8188 ( .A(n9306), .ZN(n13715) );
  NAND2_X1 U8189 ( .A1(n9029), .A2(n9028), .ZN(n14032) );
  NAND2_X1 U8190 ( .A1(n15734), .A2(n15731), .ZN(n14033) );
  AND2_X1 U8191 ( .A1(n7149), .A2(n9347), .ZN(n14036) );
  NAND2_X1 U8192 ( .A1(n7148), .A2(n7147), .ZN(n7149) );
  AND2_X1 U8193 ( .A1(n9346), .A2(n9345), .ZN(n7147) );
  NAND2_X1 U8194 ( .A1(n6673), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8798) );
  INV_X1 U8195 ( .A(n13545), .ZN(n13540) );
  NAND2_X1 U8196 ( .A1(n8611), .A2(n8610), .ZN(n14415) );
  NAND2_X1 U8197 ( .A1(n7258), .A2(n7257), .ZN(n14050) );
  AND2_X1 U8198 ( .A1(n7258), .A2(n6797), .ZN(n14052) );
  XNOR2_X1 U8199 ( .A(n12862), .B(n12863), .ZN(n14059) );
  NAND2_X1 U8200 ( .A1(n14059), .A2(n14058), .ZN(n14057) );
  NAND2_X1 U8201 ( .A1(n8628), .A2(n8627), .ZN(n12892) );
  NAND2_X1 U8202 ( .A1(n8427), .A2(n8426), .ZN(n12051) );
  NAND2_X1 U8203 ( .A1(n8479), .A2(n8478), .ZN(n14475) );
  NAND2_X1 U8204 ( .A1(n10242), .A2(n10241), .ZN(n10659) );
  NAND2_X1 U8205 ( .A1(n8340), .A2(n8339), .ZN(n11685) );
  OR2_X1 U8206 ( .A1(n8487), .A2(n8486), .ZN(n14154) );
  NAND2_X1 U8207 ( .A1(n8311), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8274) );
  NAND2_X1 U8208 ( .A1(n8310), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8271) );
  AND2_X1 U8209 ( .A1(n12212), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n14190) );
  NOR2_X1 U8210 ( .A1(n15454), .A2(n15453), .ZN(n15452) );
  NAND2_X1 U8211 ( .A1(n14200), .A2(n15484), .ZN(n7085) );
  OAI21_X1 U8212 ( .B1(n14199), .B2(n15461), .A(n7091), .ZN(n7090) );
  AOI21_X1 U8213 ( .B1(n14198), .B2(n15484), .A(n7092), .ZN(n7091) );
  NAND2_X1 U8214 ( .A1(n6883), .A2(n6882), .ZN(n8710) );
  AND2_X1 U8215 ( .A1(n14227), .A2(n7307), .ZN(n9852) );
  NOR2_X1 U8216 ( .A1(n12890), .A2(n14387), .ZN(n6894) );
  NAND2_X1 U8217 ( .A1(n7224), .A2(n7225), .ZN(n14298) );
  NAND2_X1 U8218 ( .A1(n14343), .A2(n7226), .ZN(n7224) );
  INV_X1 U8219 ( .A(n12892), .ZN(n12853) );
  NAND2_X1 U8220 ( .A1(n10052), .A2(n10051), .ZN(n14484) );
  NAND2_X1 U8221 ( .A1(n8275), .A2(n6730), .ZN(n14523) );
  INV_X1 U8222 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7482) );
  INV_X1 U8223 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10384) );
  NAND2_X1 U8224 ( .A1(n7007), .A2(n7010), .ZN(n11926) );
  OR2_X1 U8225 ( .A1(n11350), .A2(n7013), .ZN(n7007) );
  NOR2_X1 U8226 ( .A1(n7341), .A2(n15212), .ZN(n7339) );
  AND2_X1 U8227 ( .A1(n7343), .A2(n6724), .ZN(n7341) );
  NAND2_X1 U8228 ( .A1(n7343), .A2(n7347), .ZN(n7342) );
  NAND2_X1 U8229 ( .A1(n13119), .A2(n14533), .ZN(n7347) );
  AOI21_X1 U8230 ( .B1(n7010), .B2(n7013), .A(n6760), .ZN(n7008) );
  NOR2_X1 U8231 ( .A1(n7694), .A2(n6849), .ZN(n6877) );
  NAND2_X1 U8232 ( .A1(n14593), .A2(n13053), .ZN(n14557) );
  NAND2_X1 U8233 ( .A1(n14630), .A2(n13018), .ZN(n15196) );
  AND4_X1 U8234 ( .A1(n7938), .A2(n7937), .A3(n7936), .A4(n7935), .ZN(n15192)
         );
  INV_X1 U8235 ( .A(n11261), .ZN(n12599) );
  INV_X1 U8236 ( .A(n15098), .ZN(n7315) );
  NAND2_X1 U8237 ( .A1(n8008), .A2(n8007), .ZN(n15048) );
  AND2_X1 U8238 ( .A1(n14627), .A2(n15224), .ZN(n15218) );
  OR2_X1 U8239 ( .A1(n12771), .A2(n12993), .ZN(n14869) );
  AND4_X1 U8240 ( .A1(n7918), .A2(n7917), .A3(n7916), .A4(n7915), .ZN(n12999)
         );
  INV_X1 U8241 ( .A(n8165), .ZN(n14659) );
  INV_X1 U8242 ( .A(n10360), .ZN(n7056) );
  NOR2_X1 U8243 ( .A1(n7050), .A2(n7049), .ZN(n14746) );
  INV_X1 U8244 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n7049) );
  OAI21_X1 U8245 ( .B1(n7052), .B2(n14751), .A(n7051), .ZN(n7050) );
  OR2_X1 U8246 ( .A1(n14770), .A2(n14958), .ZN(n14994) );
  NOR2_X1 U8247 ( .A1(n8143), .A2(n8142), .ZN(n8210) );
  NAND2_X1 U8248 ( .A1(n7880), .A2(n7879), .ZN(n12653) );
  INV_X1 U8249 ( .A(n15277), .ZN(n14982) );
  NOR2_X1 U8250 ( .A1(n15330), .A2(n6966), .ZN(n6962) );
  AND2_X1 U8251 ( .A1(n7544), .A2(n15332), .ZN(n6964) );
  INV_X1 U8252 ( .A(n14774), .ZN(n15075) );
  NAND2_X1 U8253 ( .A1(n14994), .A2(n14999), .ZN(n15073) );
  OR2_X1 U8254 ( .A1(n15113), .A2(n15114), .ZN(n7112) );
  AND2_X1 U8255 ( .A1(n9455), .A2(n9456), .ZN(n15234) );
  AND2_X1 U8256 ( .A1(n9464), .A2(n9463), .ZN(n15241) );
  XNOR2_X1 U8257 ( .A(n9475), .B(P3_ADDR_REG_16__SCAN_IN), .ZN(n15252) );
  NAND2_X1 U8258 ( .A1(n6858), .A2(n6712), .ZN(n7110) );
  AND2_X1 U8259 ( .A1(n7110), .A2(n15494), .ZN(n7109) );
  NAND2_X1 U8260 ( .A1(n12610), .A2(n7196), .ZN(n7195) );
  OR2_X1 U8261 ( .A1(n9892), .A2(n7485), .ZN(n7484) );
  INV_X1 U8262 ( .A(n9891), .ZN(n7485) );
  NAND2_X1 U8263 ( .A1(n12621), .A2(n7207), .ZN(n7206) );
  OR2_X1 U8264 ( .A1(n9916), .A2(n7481), .ZN(n7480) );
  NAND2_X1 U8265 ( .A1(n12642), .A2(n12644), .ZN(n7200) );
  NAND2_X1 U8266 ( .A1(n9925), .A2(n9927), .ZN(n7476) );
  MUX2_X1 U8267 ( .A(n13267), .B(n13175), .S(n13174), .Z(n13182) );
  AND2_X1 U8268 ( .A1(n12668), .A2(n6773), .ZN(n7193) );
  AND2_X1 U8269 ( .A1(n14972), .A2(n12674), .ZN(n12679) );
  AND2_X1 U8270 ( .A1(n13893), .A2(n13233), .ZN(n6830) );
  NAND2_X1 U8271 ( .A1(n7488), .A2(n9991), .ZN(n7487) );
  NAND2_X1 U8272 ( .A1(n12714), .A2(n12716), .ZN(n7204) );
  NAND2_X1 U8273 ( .A1(n13786), .A2(n13274), .ZN(n6832) );
  NOR2_X1 U8274 ( .A1(n12075), .A2(n6844), .ZN(n6843) );
  NAND2_X1 U8275 ( .A1(n12041), .A2(n12105), .ZN(n6844) );
  OR2_X1 U8276 ( .A1(n13746), .A2(n7082), .ZN(n7081) );
  INV_X1 U8277 ( .A(n13740), .ZN(n7082) );
  OR2_X1 U8278 ( .A1(n9290), .A2(n13332), .ZN(n9292) );
  AOI21_X1 U8279 ( .B1(n7470), .B2(n7469), .A(n7467), .ZN(n7466) );
  OR2_X1 U8280 ( .A1(n12976), .A2(n12975), .ZN(n12979) );
  OR2_X1 U8281 ( .A1(n13298), .A2(n13297), .ZN(n13308) );
  MUX2_X1 U8282 ( .A(n13296), .B(n13295), .S(n13305), .Z(n13298) );
  AND2_X1 U8283 ( .A1(n10091), .A2(n6845), .ZN(n10093) );
  NOR2_X1 U8284 ( .A1(n14251), .A2(n6846), .ZN(n6845) );
  AND2_X1 U8285 ( .A1(n10022), .A2(n7465), .ZN(n7464) );
  NAND2_X1 U8286 ( .A1(n10020), .A2(n10023), .ZN(n7463) );
  INV_X1 U8287 ( .A(n7280), .ZN(n7279) );
  OAI21_X1 U8288 ( .B1(n7284), .B2(n7281), .A(n8679), .ZN(n7280) );
  INV_X1 U8289 ( .A(n8192), .ZN(n7528) );
  INV_X1 U8290 ( .A(n14865), .ZN(n7527) );
  NAND2_X1 U8291 ( .A1(n8072), .A2(n8071), .ZN(n8086) );
  NAND2_X1 U8292 ( .A1(n8066), .A2(n8065), .ZN(n8072) );
  INV_X1 U8293 ( .A(n8028), .ZN(n8031) );
  AND2_X1 U8294 ( .A1(n7673), .A2(n7425), .ZN(n7424) );
  NAND2_X1 U8295 ( .A1(n7426), .A2(n7670), .ZN(n7425) );
  INV_X1 U8296 ( .A(n7668), .ZN(n7426) );
  NAND2_X1 U8297 ( .A1(n7424), .A2(n7036), .ZN(n7422) );
  INV_X1 U8298 ( .A(n7667), .ZN(n7041) );
  OAI21_X1 U8299 ( .B1(n7604), .B2(n7041), .A(n7668), .ZN(n7040) );
  NAND2_X1 U8300 ( .A1(n7664), .A2(n10436), .ZN(n7667) );
  NAND2_X1 U8301 ( .A1(n7660), .A2(n10422), .ZN(n7663) );
  NOR2_X1 U8302 ( .A1(n7033), .A2(n7802), .ZN(n7029) );
  INV_X1 U8303 ( .A(n7412), .ZN(n7033) );
  INV_X1 U8304 ( .A(n7413), .ZN(n7031) );
  AOI21_X1 U8305 ( .B1(n7654), .B2(n7414), .A(n6755), .ZN(n7413) );
  INV_X1 U8306 ( .A(n7653), .ZN(n7414) );
  NOR2_X1 U8307 ( .A1(n7826), .A2(n7816), .ZN(n7412) );
  INV_X1 U8308 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7616) );
  AND2_X1 U8309 ( .A1(n12297), .A2(n13533), .ZN(n12298) );
  NOR2_X1 U8310 ( .A1(n7362), .A2(n13292), .ZN(n7361) );
  INV_X1 U8311 ( .A(n13304), .ZN(n7362) );
  NOR2_X1 U8312 ( .A1(n7359), .A2(n13721), .ZN(n7358) );
  AND2_X1 U8313 ( .A1(n13989), .A2(n13158), .ZN(n13340) );
  INV_X1 U8314 ( .A(n11838), .ZN(n6952) );
  NAND2_X1 U8315 ( .A1(n15618), .A2(n11905), .ZN(n11906) );
  NAND2_X1 U8316 ( .A1(n15652), .A2(n11908), .ZN(n11909) );
  NAND2_X1 U8317 ( .A1(n12263), .A2(n12264), .ZN(n12332) );
  OAI21_X1 U8318 ( .B1(n13545), .B2(n8989), .A(n13544), .ZN(n13559) );
  NAND2_X1 U8319 ( .A1(n13586), .A2(n13592), .ZN(n13615) );
  NAND2_X1 U8320 ( .A1(n13638), .A2(n6816), .ZN(n13641) );
  OR2_X1 U8321 ( .A1(n9311), .A2(n10170), .ZN(n9312) );
  XNOR2_X1 U8322 ( .A(n12971), .B(n13299), .ZN(n13336) );
  NOR2_X1 U8323 ( .A1(n13336), .A2(n7411), .ZN(n7410) );
  INV_X1 U8324 ( .A(n10166), .ZN(n7411) );
  NAND2_X1 U8325 ( .A1(n7410), .A2(n7409), .ZN(n9313) );
  INV_X1 U8326 ( .A(n10165), .ZN(n7409) );
  NAND2_X1 U8327 ( .A1(n6922), .A2(n9214), .ZN(n6921) );
  AOI21_X1 U8328 ( .B1(n13782), .B2(n9201), .A(n7614), .ZN(n13719) );
  AOI21_X1 U8329 ( .B1(n6916), .B2(n9124), .A(n6914), .ZN(n6913) );
  INV_X1 U8330 ( .A(n13272), .ZN(n6914) );
  OR2_X1 U8331 ( .A1(n13804), .A2(n13789), .ZN(n13272) );
  AND2_X1 U8332 ( .A1(n13268), .A2(n13269), .ZN(n13315) );
  NAND2_X1 U8333 ( .A1(n15691), .A2(n11672), .ZN(n13174) );
  NAND2_X1 U8334 ( .A1(n13174), .A2(n13176), .ZN(n11169) );
  XNOR2_X1 U8335 ( .A(n9273), .B(n15697), .ZN(n13178) );
  AOI21_X1 U8336 ( .B1(n6905), .B2(n13247), .A(n13260), .ZN(n6904) );
  AND2_X1 U8337 ( .A1(n13847), .A2(n6906), .ZN(n6905) );
  NOR2_X1 U8338 ( .A1(n7521), .A2(P3_IR_REG_17__SCAN_IN), .ZN(n6930) );
  NAND2_X1 U8339 ( .A1(n7177), .A2(n7522), .ZN(n7176) );
  AOI21_X1 U8340 ( .B1(n7075), .B2(n7077), .A(n7074), .ZN(n7073) );
  INV_X1 U8341 ( .A(n7386), .ZN(n7074) );
  INV_X1 U8342 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8758) );
  NOR2_X1 U8343 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_6__SCAN_IN), .ZN(
        n8760) );
  NOR2_X1 U8344 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n8759) );
  INV_X1 U8345 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n9007) );
  NOR2_X1 U8346 ( .A1(n8998), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n9008) );
  INV_X1 U8347 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9005) );
  OR2_X1 U8348 ( .A1(n8921), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n8938) );
  CLKBUF_X1 U8349 ( .A(n8884), .Z(n8885) );
  NOR2_X1 U8350 ( .A1(n8429), .A2(n8428), .ZN(n8440) );
  AOI21_X1 U8351 ( .B1(n10067), .B2(n6805), .A(n7452), .ZN(n7451) );
  INV_X1 U8352 ( .A(n10035), .ZN(n7452) );
  NOR2_X1 U8353 ( .A1(n6805), .A2(n10067), .ZN(n7450) );
  INV_X1 U8354 ( .A(n7307), .ZN(n7306) );
  OR2_X1 U8355 ( .A1(n14238), .A2(n6693), .ZN(n6884) );
  NOR2_X1 U8356 ( .A1(n12892), .A2(n6997), .ZN(n6996) );
  INV_X1 U8357 ( .A(n6998), .ZN(n6997) );
  NOR2_X1 U8358 ( .A1(n14415), .A2(n14420), .ZN(n6998) );
  INV_X1 U8359 ( .A(n7222), .ZN(n7221) );
  NOR2_X1 U8360 ( .A1(n7223), .A2(n14297), .ZN(n7222) );
  INV_X1 U8361 ( .A(n7225), .ZN(n7223) );
  INV_X1 U8362 ( .A(n7226), .ZN(n7220) );
  NOR2_X1 U8363 ( .A1(n6988), .A2(n14443), .ZN(n6987) );
  INV_X1 U8364 ( .A(n6989), .ZN(n6988) );
  NOR2_X1 U8365 ( .A1(n14338), .A2(n14454), .ZN(n6989) );
  NAND2_X1 U8366 ( .A1(n8682), .A2(n8681), .ZN(n7296) );
  AND2_X1 U8367 ( .A1(n8482), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8493) );
  INV_X1 U8368 ( .A(n8672), .ZN(n7302) );
  NAND2_X1 U8369 ( .A1(n11783), .A2(n12116), .ZN(n12048) );
  NOR2_X1 U8370 ( .A1(n8385), .A2(n8384), .ZN(n8401) );
  NAND2_X1 U8371 ( .A1(n11776), .A2(n11777), .ZN(n11775) );
  INV_X1 U8372 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8384) );
  OAI21_X1 U8373 ( .B1(n8349), .B2(n7250), .A(n8360), .ZN(n7249) );
  NAND2_X1 U8374 ( .A1(n11324), .A2(n11329), .ZN(n11271) );
  NOR2_X1 U8375 ( .A1(n10807), .A2(n10812), .ZN(n10848) );
  NOR2_X2 U8376 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n8514) );
  INV_X1 U8377 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n8379) );
  OR2_X1 U8378 ( .A1(n8363), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n8378) );
  AOI21_X1 U8379 ( .B1(n14533), .B2(n7349), .A(n6763), .ZN(n7348) );
  AND2_X1 U8380 ( .A1(n12823), .A2(n12822), .ZN(n12834) );
  OAI21_X1 U8381 ( .B1(n10203), .B2(n11213), .A(n7785), .ZN(n7537) );
  INV_X1 U8382 ( .A(n14803), .ZN(n13101) );
  INV_X1 U8383 ( .A(n14643), .ZN(n13091) );
  AND2_X1 U8384 ( .A1(n14898), .A2(n14645), .ZN(n8062) );
  NAND2_X1 U8385 ( .A1(n14915), .A2(n8044), .ZN(n8045) );
  NAND2_X1 U8386 ( .A1(n7567), .A2(n12801), .ZN(n7569) );
  INV_X1 U8387 ( .A(n14891), .ZN(n7567) );
  NOR2_X1 U8388 ( .A1(n12802), .A2(n8015), .ZN(n7576) );
  NAND2_X1 U8389 ( .A1(n14953), .A2(n7578), .ZN(n6863) );
  INV_X1 U8390 ( .A(n7578), .ZN(n6864) );
  OR2_X1 U8391 ( .A1(n14915), .A2(n14888), .ZN(n8192) );
  NAND2_X1 U8392 ( .A1(n13017), .A2(n14579), .ZN(n7555) );
  NOR2_X1 U8393 ( .A1(n13009), .A2(n15200), .ZN(n7138) );
  NOR2_X1 U8394 ( .A1(n12668), .A2(n7905), .ZN(n6876) );
  AOI21_X1 U8395 ( .B1(n11552), .B2(n7565), .A(n6745), .ZN(n7563) );
  NAND2_X1 U8396 ( .A1(n11587), .A2(n7743), .ZN(n10770) );
  NAND2_X1 U8397 ( .A1(n10590), .A2(n6865), .ZN(n8154) );
  INV_X1 U8398 ( .A(n15274), .ZN(n12578) );
  AOI21_X1 U8399 ( .B1(n9845), .B2(n9848), .A(n7446), .ZN(n7445) );
  INV_X1 U8400 ( .A(n10041), .ZN(n7446) );
  INV_X1 U8401 ( .A(n9848), .ZN(n7443) );
  NOR2_X1 U8402 ( .A1(n7999), .A2(n7441), .ZN(n7440) );
  INV_X1 U8403 ( .A(n7958), .ZN(n7441) );
  NAND2_X1 U8404 ( .A1(n7437), .A2(n7438), .ZN(n8034) );
  NAND2_X1 U8405 ( .A1(n7959), .A2(n7440), .ZN(n7437) );
  XNOR2_X1 U8406 ( .A(n7941), .B(SI_16_), .ZN(n7939) );
  INV_X1 U8407 ( .A(n7641), .ZN(n7419) );
  INV_X1 U8408 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n7688) );
  NAND2_X1 U8409 ( .A1(n7624), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6848) );
  AND2_X1 U8410 ( .A1(n7116), .A2(n7115), .ZN(n9385) );
  NAND2_X1 U8411 ( .A1(n9384), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n7115) );
  INV_X1 U8412 ( .A(n9419), .ZN(n7117) );
  XNOR2_X1 U8413 ( .A(n9388), .B(n9389), .ZN(n9416) );
  OAI21_X1 U8414 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n9806), .A(n9400), .ZN(
        n9401) );
  NAND2_X1 U8415 ( .A1(n15237), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n7124) );
  NAND2_X1 U8416 ( .A1(n12127), .A2(n7184), .ZN(n7182) );
  NAND2_X1 U8417 ( .A1(n11083), .A2(n13176), .ZN(n11166) );
  OR2_X1 U8418 ( .A1(n12927), .A2(n12926), .ZN(n13405) );
  NAND2_X1 U8419 ( .A1(n7156), .A2(n6741), .ZN(n13406) );
  OR2_X1 U8420 ( .A1(n13503), .A2(n6796), .ZN(n7160) );
  AOI21_X1 U8421 ( .B1(n7592), .B2(n13909), .A(n7170), .ZN(n7169) );
  INV_X1 U8422 ( .A(n7166), .ZN(n7165) );
  OAI21_X1 U8423 ( .B1(n7172), .B2(n13529), .A(n7167), .ZN(n7166) );
  INV_X1 U8424 ( .A(n12905), .ZN(n7161) );
  AND2_X1 U8425 ( .A1(n13429), .A2(n12944), .ZN(n13456) );
  NOR2_X1 U8426 ( .A1(n9177), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9208) );
  AND2_X1 U8427 ( .A1(n6896), .A2(n9274), .ZN(n11083) );
  INV_X1 U8428 ( .A(n13536), .ZN(n6896) );
  AND2_X1 U8429 ( .A1(n9132), .A2(n13471), .ZN(n9151) );
  OR2_X1 U8430 ( .A1(n9186), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9188) );
  XNOR2_X1 U8431 ( .A(n13364), .B(n11672), .ZN(n7155) );
  OR2_X1 U8432 ( .A1(n8843), .A2(n11177), .ZN(n8792) );
  NOR2_X1 U8433 ( .A1(n10858), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11218) );
  OR2_X1 U8434 ( .A1(n10872), .A2(n10871), .ZN(n10938) );
  OAI21_X1 U8435 ( .B1(P3_IR_REG_1__SCAN_IN), .B2(n10939), .A(n10938), .ZN(
        n10940) );
  XNOR2_X1 U8436 ( .A(n11901), .B(n15561), .ZN(n15562) );
  AOI21_X1 U8437 ( .B1(n15562), .B2(P3_REG1_REG_3__SCAN_IN), .A(n6852), .ZN(
        n15581) );
  AND2_X1 U8438 ( .A1(n11901), .A2(n11902), .ZN(n6852) );
  NOR2_X1 U8439 ( .A1(n15581), .A2(n15580), .ZN(n15579) );
  AOI21_X1 U8440 ( .B1(n15573), .B2(n15572), .A(n15571), .ZN(n15594) );
  XOR2_X1 U8441 ( .A(n11906), .B(n15633), .Z(n15637) );
  AND2_X1 U8442 ( .A1(n6949), .A2(n11841), .ZN(n11842) );
  INV_X1 U8443 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n12129) );
  NOR2_X1 U8444 ( .A1(n11842), .A2(n11875), .ZN(n11843) );
  AOI21_X1 U8445 ( .B1(n15646), .B2(n15645), .A(n15644), .ZN(n15665) );
  OR2_X1 U8446 ( .A1(n15659), .A2(n11846), .ZN(n6946) );
  XNOR2_X1 U8447 ( .A(n12328), .B(n12332), .ZN(n12265) );
  NOR2_X1 U8448 ( .A1(n12272), .A2(n12271), .ZN(n12342) );
  XNOR2_X1 U8449 ( .A(n13559), .B(n13566), .ZN(n13546) );
  NAND2_X1 U8450 ( .A1(n13546), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n13561) );
  OR2_X1 U8451 ( .A1(n13556), .A2(n13557), .ZN(n6948) );
  NAND2_X1 U8452 ( .A1(n13564), .A2(n13570), .ZN(n13586) );
  NAND2_X1 U8453 ( .A1(n6947), .A2(n13591), .ZN(n7272) );
  NOR2_X1 U8454 ( .A1(n13595), .A2(n13596), .ZN(n13609) );
  OAI21_X1 U8455 ( .B1(n6955), .B2(n13604), .A(n6954), .ZN(n13650) );
  NAND2_X1 U8456 ( .A1(n13606), .A2(n6956), .ZN(n6954) );
  XNOR2_X1 U8457 ( .A(n13641), .B(n15130), .ZN(n15129) );
  AOI21_X1 U8458 ( .B1(n15128), .B2(n13643), .A(n13642), .ZN(n13671) );
  NOR2_X1 U8459 ( .A1(n13671), .A2(n6825), .ZN(n13675) );
  NOR2_X1 U8460 ( .A1(n13664), .A2(n13965), .ZN(n6825) );
  AOI21_X1 U8461 ( .B1(n13633), .B2(n13649), .A(n15134), .ZN(n13665) );
  NAND2_X1 U8462 ( .A1(n13652), .A2(n13660), .ZN(n6944) );
  NAND2_X1 U8463 ( .A1(n13662), .A2(n6944), .ZN(n6943) );
  AND2_X1 U8464 ( .A1(n13310), .A2(n13306), .ZN(n13338) );
  OR2_X1 U8465 ( .A1(n13690), .A2(n9251), .ZN(n13708) );
  INV_X1 U8466 ( .A(n13336), .ZN(n13297) );
  NAND2_X1 U8467 ( .A1(n9313), .A2(n7408), .ZN(n10170) );
  NAND2_X1 U8468 ( .A1(n7410), .A2(n10150), .ZN(n7408) );
  INV_X1 U8469 ( .A(n7510), .ZN(n7509) );
  OAI21_X1 U8470 ( .B1(n6799), .B2(n7511), .A(n13746), .ZN(n7510) );
  AND2_X1 U8471 ( .A1(n13757), .A2(n13739), .ZN(n13773) );
  NAND2_X1 U8472 ( .A1(n6909), .A2(n6913), .ZN(n13782) );
  NAND2_X1 U8473 ( .A1(n13816), .A2(n6916), .ZN(n6909) );
  INV_X1 U8474 ( .A(n13315), .ZN(n13815) );
  OR2_X1 U8475 ( .A1(n9100), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9118) );
  INV_X1 U8476 ( .A(n13831), .ZN(n9106) );
  NOR2_X1 U8477 ( .A1(n13825), .A2(n9106), .ZN(n13824) );
  NAND2_X1 U8478 ( .A1(n9081), .A2(n9635), .ZN(n9100) );
  AND2_X1 U8479 ( .A1(n9067), .A2(n13441), .ZN(n9081) );
  AND2_X1 U8480 ( .A1(n13240), .A2(n13250), .ZN(n13865) );
  AND2_X1 U8481 ( .A1(n7365), .A2(n6924), .ZN(n6923) );
  AND2_X1 U8482 ( .A1(n7490), .A2(n7489), .ZN(n13876) );
  OAI21_X1 U8483 ( .B1(n13894), .B2(n7491), .A(n15142), .ZN(n7490) );
  NOR2_X1 U8484 ( .A1(n8987), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9014) );
  AND4_X1 U8485 ( .A1(n9036), .A2(n9035), .A3(n9034), .A4(n9033), .ZN(n13896)
         );
  AOI21_X1 U8486 ( .B1(n13907), .B2(n13906), .A(n7492), .ZN(n13894) );
  AND2_X1 U8487 ( .A1(n13483), .A2(n12897), .ZN(n7492) );
  OAI22_X1 U8488 ( .A1(n12524), .A2(n13909), .B1(n9288), .B2(n15150), .ZN(
        n13907) );
  AND2_X1 U8489 ( .A1(n12524), .A2(n13909), .ZN(n9288) );
  OR2_X1 U8490 ( .A1(n8970), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8987) );
  AND2_X1 U8491 ( .A1(n13227), .A2(n13226), .ZN(n13327) );
  AOI21_X1 U8492 ( .B1(n6900), .B2(n6902), .A(n6899), .ZN(n6898) );
  INV_X1 U8493 ( .A(n6901), .ZN(n6900) );
  INV_X1 U8494 ( .A(n7514), .ZN(n7513) );
  OAI21_X1 U8495 ( .B1(n7517), .B2(n7515), .A(n9287), .ZN(n7514) );
  NAND2_X1 U8496 ( .A1(n8932), .A2(n8931), .ZN(n8952) );
  AND2_X1 U8497 ( .A1(n8913), .A2(n12129), .ZN(n8932) );
  OR2_X1 U8498 ( .A1(n12152), .A2(n7517), .ZN(n12280) );
  NOR2_X1 U8499 ( .A1(n12153), .A2(n13326), .ZN(n12152) );
  OR2_X1 U8500 ( .A1(n8878), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8894) );
  NOR2_X1 U8501 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8861) );
  AND2_X1 U8502 ( .A1(n8778), .A2(n9366), .ZN(n13728) );
  INV_X1 U8503 ( .A(n11083), .ZN(n13172) );
  AND2_X1 U8504 ( .A1(n11159), .A2(n13666), .ZN(n11501) );
  AND4_X1 U8505 ( .A1(n11118), .A2(n9372), .A3(n9376), .A4(n9378), .ZN(n11364)
         );
  NAND2_X1 U8506 ( .A1(n13146), .A2(n13145), .ZN(n13159) );
  OR2_X1 U8507 ( .A1(n13126), .A2(n10182), .ZN(n10183) );
  AND2_X1 U8508 ( .A1(n13728), .A2(n10182), .ZN(n15726) );
  NAND2_X1 U8509 ( .A1(n9262), .A2(n9261), .ZN(n13136) );
  INV_X1 U8510 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8797) );
  NAND2_X1 U8511 ( .A1(n8784), .A2(n7522), .ZN(n7520) );
  NAND2_X1 U8512 ( .A1(n7407), .A2(n9217), .ZN(n9229) );
  NAND2_X1 U8513 ( .A1(n9216), .A2(n9215), .ZN(n7407) );
  AND2_X1 U8514 ( .A1(n8766), .A2(n8764), .ZN(n8771) );
  OR2_X1 U8515 ( .A1(n9025), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n9047) );
  AOI21_X1 U8516 ( .B1(n7377), .B2(n7379), .A(n7375), .ZN(n7374) );
  NAND2_X1 U8517 ( .A1(n7065), .A2(n7064), .ZN(n7376) );
  INV_X1 U8518 ( .A(n8981), .ZN(n7375) );
  OR2_X1 U8519 ( .A1(n8977), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n8998) );
  INV_X1 U8520 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8964) );
  NOR2_X1 U8521 ( .A1(n8938), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n8942) );
  AND2_X1 U8522 ( .A1(n8870), .A2(n8853), .ZN(n8868) );
  AND2_X1 U8523 ( .A1(n8830), .A2(n8819), .ZN(n8828) );
  OR2_X1 U8524 ( .A1(n14040), .A2(n10943), .ZN(n7270) );
  NAND2_X1 U8525 ( .A1(n7373), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8814) );
  INV_X1 U8526 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n7373) );
  OR2_X1 U8527 ( .A1(n8456), .A2(n8455), .ZN(n8470) );
  AND3_X1 U8528 ( .A1(n14128), .A2(n7043), .A3(n6828), .ZN(n6855) );
  NAND2_X1 U8529 ( .A1(n10308), .A2(n6740), .ZN(n7042) );
  OR2_X1 U8530 ( .A1(n8354), .A2(n11094), .ZN(n8369) );
  INV_X1 U8531 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8368) );
  NOR2_X1 U8532 ( .A1(n7217), .A2(n7216), .ZN(n7215) );
  OR2_X1 U8533 ( .A1(n10309), .A2(n12401), .ZN(n7243) );
  AND2_X1 U8534 ( .A1(n10309), .A2(n12401), .ZN(n7242) );
  AND2_X1 U8535 ( .A1(n10282), .A2(n11242), .ZN(n7259) );
  NAND2_X1 U8536 ( .A1(n11244), .A2(n11243), .ZN(n7260) );
  AND2_X1 U8537 ( .A1(n10295), .A2(n10289), .ZN(n7252) );
  NOR2_X1 U8538 ( .A1(n8544), .A2(n8542), .ZN(n8557) );
  OR2_X1 U8539 ( .A1(n8417), .A2(n11303), .ZN(n8429) );
  XNOR2_X1 U8540 ( .A(n12409), .B(n12877), .ZN(n10309) );
  NAND2_X1 U8541 ( .A1(n15344), .A2(n10977), .ZN(n7105) );
  AOI21_X1 U8542 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(n15344), .A(n15339), .ZN(
        n14173) );
  AND2_X1 U8543 ( .A1(n7096), .A2(n7095), .ZN(n15391) );
  NAND2_X1 U8544 ( .A1(n15382), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7095) );
  OR2_X1 U8545 ( .A1(n8639), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n8363) );
  AND2_X1 U8546 ( .A1(n10984), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7099) );
  OR2_X1 U8547 ( .A1(n11979), .A2(n11980), .ZN(n12219) );
  AND2_X1 U8548 ( .A1(n12221), .A2(n12222), .ZN(n14183) );
  INV_X1 U8549 ( .A(n15488), .ZN(n7103) );
  INV_X1 U8550 ( .A(n10092), .ZN(n8696) );
  NOR2_X1 U8551 ( .A1(n8696), .A2(n6693), .ZN(n7307) );
  NAND2_X1 U8552 ( .A1(n8695), .A2(n6685), .ZN(n6883) );
  AOI21_X1 U8553 ( .B1(n6685), .B2(n6693), .A(n14395), .ZN(n6882) );
  NAND2_X1 U8554 ( .A1(n14270), .A2(n6998), .ZN(n14231) );
  AND2_X1 U8555 ( .A1(n14289), .A2(n14495), .ZN(n14270) );
  NAND2_X1 U8556 ( .A1(n14270), .A2(n14249), .ZN(n14244) );
  OAI21_X1 U8557 ( .B1(n14333), .B2(n6887), .A(n6885), .ZN(n8692) );
  AOI21_X1 U8558 ( .B1(n7309), .B2(n6886), .A(n6762), .ZN(n6885) );
  NAND2_X1 U8559 ( .A1(n14328), .A2(n7309), .ZN(n14262) );
  NAND2_X1 U8560 ( .A1(n14328), .A2(n8690), .ZN(n14300) );
  NAND2_X1 U8561 ( .A1(n14347), .A2(n6987), .ZN(n14316) );
  AOI21_X1 U8562 ( .B1(n7293), .B2(n8680), .A(n7292), .ZN(n7291) );
  INV_X1 U8563 ( .A(n8685), .ZN(n7292) );
  NAND2_X1 U8564 ( .A1(n14347), .A2(n8712), .ZN(n14348) );
  NAND2_X1 U8565 ( .A1(n7296), .A2(n8683), .ZN(n14364) );
  AOI21_X1 U8566 ( .B1(n7234), .B2(n7233), .A(n6695), .ZN(n7232) );
  NOR2_X1 U8567 ( .A1(n12048), .A2(n12051), .ZN(n12078) );
  AND2_X1 U8568 ( .A1(n10534), .A2(n8705), .ZN(n14369) );
  AND2_X1 U8569 ( .A1(n10534), .A2(n8706), .ZN(n14368) );
  OR2_X1 U8570 ( .A1(n11271), .A2(n11088), .ZN(n11380) );
  NOR2_X1 U8571 ( .A1(n11073), .A2(n11074), .ZN(n11324) );
  INV_X1 U8572 ( .A(n10235), .ZN(n10748) );
  OR2_X1 U8573 ( .A1(n10576), .A2(n10746), .ZN(n10550) );
  NAND2_X1 U8574 ( .A1(n10576), .A2(n10746), .ZN(n10235) );
  INV_X1 U8575 ( .A(n15520), .ZN(n14478) );
  INV_X1 U8576 ( .A(n15525), .ZN(n15532) );
  NOR2_X1 U8577 ( .A1(n8639), .A2(n7290), .ZN(n7289) );
  XNOR2_X1 U8578 ( .A(n8640), .B(P2_IR_REG_20__SCAN_IN), .ZN(n10077) );
  NAND2_X1 U8579 ( .A1(n7264), .A2(n6710), .ZN(n8641) );
  INV_X1 U8580 ( .A(n8639), .ZN(n7264) );
  INV_X1 U8581 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n7458) );
  INV_X1 U8582 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7459) );
  INV_X1 U8583 ( .A(n8054), .ZN(n8055) );
  NAND2_X1 U8584 ( .A1(n8055), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8076) );
  INV_X1 U8585 ( .A(n7348), .ZN(n7346) );
  INV_X1 U8586 ( .A(n6705), .ZN(n7013) );
  NAND2_X1 U8587 ( .A1(n7012), .A2(n6705), .ZN(n7011) );
  INV_X1 U8588 ( .A(n11349), .ZN(n7012) );
  XNOR2_X1 U8589 ( .A(n10593), .B(n6706), .ZN(n10594) );
  INV_X1 U8590 ( .A(n8095), .ZN(n8096) );
  INV_X1 U8591 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7780) );
  NOR2_X1 U8592 ( .A1(n7781), .A2(n7780), .ZN(n7796) );
  NOR2_X1 U8593 ( .A1(n8010), .A2(n8009), .ZN(n8023) );
  INV_X1 U8594 ( .A(n12449), .ZN(n12452) );
  NAND2_X1 U8595 ( .A1(n8037), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8054) );
  NAND2_X1 U8596 ( .A1(n14603), .A2(n14604), .ZN(n14602) );
  NAND2_X1 U8597 ( .A1(n12748), .A2(n12750), .ZN(n7198) );
  INV_X1 U8598 ( .A(n12754), .ZN(n10210) );
  INV_X1 U8599 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10918) );
  NOR2_X1 U8600 ( .A1(n11053), .A2(n7046), .ZN(n11055) );
  AND2_X1 U8601 ( .A1(n11054), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7046) );
  NAND2_X1 U8602 ( .A1(n11055), .A2(n11056), .ZN(n11419) );
  NOR2_X1 U8603 ( .A1(n7045), .A2(n7044), .ZN(n11422) );
  NOR2_X1 U8604 ( .A1(n11420), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7044) );
  INV_X1 U8605 ( .A(n11419), .ZN(n7045) );
  OR2_X1 U8606 ( .A1(n11423), .A2(n11422), .ZN(n11715) );
  INV_X1 U8607 ( .A(n7047), .ZN(n14696) );
  XNOR2_X1 U8608 ( .A(n14755), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n14756) );
  NOR2_X1 U8609 ( .A1(n7142), .A2(n7143), .ZN(n7141) );
  NAND2_X1 U8610 ( .A1(n15079), .A2(n14826), .ZN(n7142) );
  NOR2_X1 U8611 ( .A1(n14810), .A2(n7143), .ZN(n14778) );
  NAND2_X1 U8612 ( .A1(n10197), .A2(n10196), .ZN(n14809) );
  NAND2_X1 U8613 ( .A1(n8122), .A2(n6696), .ZN(n10220) );
  NAND2_X1 U8614 ( .A1(n10220), .A2(n7573), .ZN(n14808) );
  NOR2_X1 U8615 ( .A1(n14799), .A2(n7574), .ZN(n7573) );
  INV_X1 U8616 ( .A(n10219), .ZN(n7574) );
  NAND2_X1 U8617 ( .A1(n8122), .A2(n8121), .ZN(n8141) );
  INV_X1 U8618 ( .A(n12806), .ZN(n14831) );
  NAND2_X1 U8619 ( .A1(n6869), .A2(n6687), .ZN(n6867) );
  NAND2_X1 U8620 ( .A1(n6969), .A2(n8193), .ZN(n6968) );
  INV_X1 U8621 ( .A(n14883), .ZN(n14880) );
  INV_X1 U8622 ( .A(n8076), .ZN(n8077) );
  OAI21_X1 U8623 ( .B1(n8191), .B2(n6972), .A(n6970), .ZN(n14868) );
  NAND2_X1 U8624 ( .A1(n7569), .A2(n6711), .ZN(n14863) );
  NAND2_X1 U8625 ( .A1(n14893), .A2(n8212), .ZN(n14894) );
  INV_X1 U8626 ( .A(n7569), .ZN(n14890) );
  NAND2_X1 U8627 ( .A1(n14903), .A2(n8192), .ZN(n14886) );
  NAND2_X1 U8628 ( .A1(n14886), .A2(n14892), .ZN(n14885) );
  NOR2_X1 U8629 ( .A1(n14924), .A2(n15035), .ZN(n14893) );
  NAND2_X1 U8630 ( .A1(n8191), .A2(n8190), .ZN(n14903) );
  NOR2_X1 U8631 ( .A1(n14959), .A2(n15048), .ZN(n14943) );
  NAND2_X1 U8632 ( .A1(n7539), .A2(n7538), .ZN(n14933) );
  NAND2_X1 U8633 ( .A1(n6764), .A2(n12692), .ZN(n7538) );
  OR2_X1 U8634 ( .A1(n14986), .A2(n14965), .ZN(n14959) );
  NAND3_X1 U8635 ( .A1(n12228), .A2(n6688), .A3(n7137), .ZN(n14986) );
  NAND2_X1 U8636 ( .A1(n12228), .A2(n6688), .ZN(n14985) );
  NAND2_X1 U8637 ( .A1(n7966), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n7990) );
  NOR2_X1 U8638 ( .A1(n7933), .A2(n7706), .ZN(n7950) );
  AND2_X1 U8639 ( .A1(n7950), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n7966) );
  INV_X1 U8640 ( .A(n6874), .ZN(n12554) );
  OAI22_X1 U8641 ( .A1(n12175), .A2(n6875), .B1(n7549), .B2(n7551), .ZN(n6874)
         );
  NAND2_X1 U8642 ( .A1(n7550), .A2(n6876), .ZN(n6875) );
  AND2_X1 U8643 ( .A1(n12798), .A2(n7553), .ZN(n7549) );
  NAND2_X1 U8644 ( .A1(n12228), .A2(n8211), .ZN(n12465) );
  AND2_X1 U8645 ( .A1(n7881), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7899) );
  AND2_X1 U8646 ( .A1(n6694), .A2(n11606), .ZN(n12135) );
  INV_X1 U8647 ( .A(n7533), .ZN(n7532) );
  AND2_X1 U8648 ( .A1(n7530), .A2(n6794), .ZN(n7531) );
  NAND2_X1 U8649 ( .A1(n7557), .A2(n7560), .ZN(n11803) );
  AND2_X1 U8650 ( .A1(n7561), .A2(n7858), .ZN(n7560) );
  OR2_X1 U8651 ( .A1(n7836), .A2(n7704), .ZN(n7851) );
  NOR2_X1 U8652 ( .A1(n6751), .A2(n6975), .ZN(n6974) );
  AND2_X1 U8653 ( .A1(n10926), .A2(n11148), .ZN(n11549) );
  NOR2_X1 U8654 ( .A1(n10836), .A2(n12599), .ZN(n10926) );
  INV_X1 U8655 ( .A(n14869), .ZN(n14974) );
  NOR2_X1 U8656 ( .A1(n10590), .A2(n12578), .ZN(n11590) );
  NAND2_X1 U8657 ( .A1(n11563), .A2(n7729), .ZN(n11588) );
  NAND2_X1 U8658 ( .A1(n8155), .A2(n8154), .ZN(n12775) );
  NAND2_X1 U8659 ( .A1(n12775), .A2(n11564), .ZN(n11563) );
  INV_X1 U8660 ( .A(n14795), .ZN(n10218) );
  AND2_X1 U8661 ( .A1(n14812), .A2(n14811), .ZN(n15003) );
  OR2_X1 U8662 ( .A1(n14839), .A2(n14838), .ZN(n15011) );
  NAND2_X1 U8663 ( .A1(n6976), .A2(n8166), .ZN(n11553) );
  XNOR2_X1 U8664 ( .A(n10055), .B(n10054), .ZN(n12960) );
  XNOR2_X1 U8665 ( .A(n9846), .B(n9845), .ZN(n12494) );
  NOR2_X1 U8666 ( .A1(n8148), .A2(n7679), .ZN(n8224) );
  XNOR2_X1 U8667 ( .A(n8124), .B(n8107), .ZN(n12384) );
  OAI21_X2 U8668 ( .B1(n7959), .B2(n7436), .A(n7432), .ZN(n8066) );
  AOI21_X1 U8669 ( .B1(n7435), .B2(n7434), .A(n7433), .ZN(n7432) );
  INV_X1 U8670 ( .A(n8033), .ZN(n7433) );
  INV_X1 U8671 ( .A(n7440), .ZN(n7434) );
  MUX2_X1 U8672 ( .A(n7983), .B(P1_IR_REG_31__SCAN_IN), .S(n7984), .Z(n7985)
         );
  NAND2_X1 U8673 ( .A1(n7982), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7983) );
  XNOR2_X1 U8674 ( .A(n7926), .B(n7925), .ZN(n11078) );
  NAND2_X1 U8675 ( .A1(n7415), .A2(n7653), .ZN(n7827) );
  NAND2_X1 U8676 ( .A1(n7817), .A2(n7651), .ZN(n7415) );
  OR2_X1 U8677 ( .A1(n7771), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n7773) );
  NAND2_X1 U8678 ( .A1(n7421), .A2(n7641), .ZN(n7769) );
  NAND2_X1 U8679 ( .A1(n7758), .A2(n7639), .ZN(n7421) );
  AND2_X1 U8680 ( .A1(n6850), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n9422) );
  INV_X1 U8681 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n11219) );
  XNOR2_X1 U8682 ( .A(n9416), .B(n7119), .ZN(n9417) );
  INV_X1 U8683 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n7119) );
  NOR2_X1 U8684 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n9432), .ZN(n9394) );
  INV_X1 U8685 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n9716) );
  XOR2_X1 U8686 ( .A(n9592), .B(n9397), .Z(n9439) );
  NOR2_X1 U8687 ( .A1(n9445), .A2(n9446), .ZN(n9449) );
  AND2_X1 U8688 ( .A1(n6857), .A2(n6856), .ZN(n9412) );
  NAND2_X1 U8689 ( .A1(n9460), .A2(P3_ADDR_REG_13__SCAN_IN), .ZN(n6856) );
  INV_X1 U8690 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n6851) );
  NOR2_X1 U8691 ( .A1(n12025), .A2(n7183), .ZN(n12128) );
  INV_X1 U8692 ( .A(n12981), .ZN(n7152) );
  OAI21_X1 U8693 ( .B1(n13481), .B2(n13477), .A(n13478), .ZN(n13385) );
  NAND2_X1 U8694 ( .A1(n13385), .A2(n13384), .ZN(n13383) );
  OAI21_X1 U8695 ( .B1(n12941), .B2(n12940), .A(n13455), .ZN(n13393) );
  INV_X1 U8696 ( .A(n7159), .ZN(n13399) );
  AOI21_X1 U8697 ( .B1(n13502), .B2(n13503), .A(n6796), .ZN(n7159) );
  NAND2_X1 U8698 ( .A1(n9249), .A2(n9248), .ZN(n13707) );
  INV_X1 U8699 ( .A(n7180), .ZN(n12300) );
  OAI21_X1 U8700 ( .B1(n12025), .B2(n7182), .A(n6715), .ZN(n7180) );
  NAND2_X1 U8701 ( .A1(n7164), .A2(n7162), .ZN(n13440) );
  INV_X1 U8702 ( .A(n7163), .ZN(n7162) );
  NAND2_X1 U8703 ( .A1(n13385), .A2(n6726), .ZN(n7164) );
  OAI21_X1 U8704 ( .B1(n12905), .B2(n12903), .A(n12904), .ZN(n7163) );
  AND3_X1 U8705 ( .A1(n8877), .A2(n8876), .A3(n8875), .ZN(n11660) );
  NAND2_X1 U8706 ( .A1(n11572), .A2(n11571), .ZN(n11653) );
  AND4_X1 U8707 ( .A1(n8957), .A2(n8956), .A3(n8955), .A4(n8954), .ZN(n12526)
         );
  NAND2_X1 U8708 ( .A1(n9131), .A2(n9130), .ZN(n13804) );
  OR2_X1 U8709 ( .A1(n13150), .A2(n11026), .ZN(n9130) );
  OR2_X1 U8710 ( .A1(n11027), .A2(n9145), .ZN(n9131) );
  NAND2_X1 U8711 ( .A1(n12506), .A2(n7170), .ZN(n12896) );
  INV_X1 U8712 ( .A(n13495), .ZN(n13516) );
  AND4_X1 U8713 ( .A1(n8867), .A2(n8866), .A3(n8865), .A4(n8864), .ZN(n12007)
         );
  AND4_X1 U8714 ( .A1(n8899), .A2(n8898), .A3(n8897), .A4(n8896), .ZN(n12155)
         );
  OR2_X1 U8715 ( .A1(n11172), .A2(n15690), .ZN(n13495) );
  OR2_X1 U8716 ( .A1(n11172), .A2(n15689), .ZN(n13514) );
  NAND2_X1 U8717 ( .A1(n11114), .A2(n11118), .ZN(n13523) );
  NAND2_X1 U8718 ( .A1(n13914), .A2(n11121), .ZN(n13520) );
  AOI21_X1 U8719 ( .B1(n13164), .B2(n13163), .A(n13162), .ZN(n13165) );
  NAND2_X1 U8720 ( .A1(n13133), .A2(n13310), .ZN(n13164) );
  OAI211_X1 U8721 ( .C1(n11521), .C2(n13942), .A(n9179), .B(n9178), .ZN(n13747) );
  AND3_X1 U8722 ( .A1(n9155), .A2(n9154), .A3(n9153), .ZN(n13801) );
  INV_X1 U8723 ( .A(n13789), .ZN(n13812) );
  NAND4_X1 U8724 ( .A1(n9105), .A2(n9104), .A3(n9103), .A4(n9102), .ZN(n13842)
         );
  INV_X1 U8725 ( .A(n13828), .ZN(n13852) );
  NAND4_X1 U8726 ( .A1(n9056), .A2(n9055), .A3(n9054), .A4(n9053), .ZN(n13878)
         );
  INV_X1 U8727 ( .A(n13896), .ZN(n13528) );
  INV_X1 U8728 ( .A(n13897), .ZN(n13483) );
  INV_X1 U8729 ( .A(n12526), .ZN(n13530) );
  NAND2_X1 U8730 ( .A1(n14035), .A2(n10233), .ZN(n13532) );
  NOR2_X1 U8731 ( .A1(n10859), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11222) );
  AOI21_X1 U8732 ( .B1(n10957), .B2(n10956), .A(n10955), .ZN(n15557) );
  NOR2_X1 U8733 ( .A1(n15551), .A2(n11838), .ZN(n15567) );
  AND2_X1 U8734 ( .A1(n11840), .A2(n11864), .ZN(n6950) );
  INV_X1 U8735 ( .A(n6949), .ZN(n15607) );
  XNOR2_X1 U8736 ( .A(n11842), .B(n11875), .ZN(n15626) );
  NOR2_X1 U8737 ( .A1(n15626), .A2(n11874), .ZN(n15625) );
  OAI21_X1 U8738 ( .B1(n15626), .B2(n7274), .A(n7273), .ZN(n15642) );
  NAND2_X1 U8739 ( .A1(n7275), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7274) );
  NAND2_X1 U8740 ( .A1(n11843), .A2(n7275), .ZN(n7273) );
  INV_X1 U8741 ( .A(n15643), .ZN(n7275) );
  XNOR2_X1 U8742 ( .A(n11845), .B(n11910), .ZN(n15660) );
  NOR2_X1 U8743 ( .A1(n15660), .A2(n15661), .ZN(n15659) );
  AND2_X1 U8744 ( .A1(n6946), .A2(n6945), .ZN(n12260) );
  INV_X1 U8745 ( .A(n11848), .ZN(n6945) );
  INV_X1 U8746 ( .A(n6946), .ZN(n11849) );
  INV_X1 U8747 ( .A(n7268), .ZN(n12329) );
  NOR2_X1 U8748 ( .A1(n13538), .A2(n13899), .ZN(n13556) );
  INV_X1 U8749 ( .A(n6947), .ZN(n13582) );
  INV_X1 U8750 ( .A(n6948), .ZN(n13558) );
  XNOR2_X1 U8751 ( .A(n7272), .B(n13616), .ZN(n13584) );
  NOR2_X1 U8752 ( .A1(n13604), .A2(n13605), .ZN(n13607) );
  XNOR2_X1 U8753 ( .A(n13650), .B(n15130), .ZN(n15126) );
  INV_X1 U8754 ( .A(n13654), .ZN(n15125) );
  XNOR2_X1 U8755 ( .A(n13699), .B(n13700), .ZN(n13929) );
  AOI21_X1 U8756 ( .B1(n13706), .B2(n13705), .A(n13704), .ZN(n13928) );
  XNOR2_X1 U8757 ( .A(n10147), .B(n13335), .ZN(n13717) );
  AND2_X1 U8758 ( .A1(n13742), .A2(n13741), .ZN(n13744) );
  AND2_X1 U8759 ( .A1(n9304), .A2(n9303), .ZN(n13762) );
  NAND2_X1 U8760 ( .A1(n7496), .A2(n7497), .ZN(n13785) );
  NAND2_X1 U8761 ( .A1(n6918), .A2(n13269), .ZN(n13803) );
  NAND2_X1 U8762 ( .A1(n6919), .A2(n13268), .ZN(n6918) );
  INV_X1 U8763 ( .A(n13816), .ZN(n6919) );
  NAND2_X1 U8764 ( .A1(n13856), .A2(n13251), .ZN(n13848) );
  NAND2_X1 U8765 ( .A1(n9066), .A2(n9065), .ZN(n13971) );
  NAND2_X1 U8766 ( .A1(n7366), .A2(n13230), .ZN(n13884) );
  NAND2_X1 U8767 ( .A1(n13910), .A2(n6926), .ZN(n7366) );
  NAND2_X1 U8768 ( .A1(n13910), .A2(n13231), .ZN(n13892) );
  NAND2_X1 U8769 ( .A1(n12156), .A2(n13212), .ZN(n12279) );
  OAI21_X1 U8770 ( .B1(n12001), .B2(n12023), .A(n7352), .ZN(n12157) );
  NAND2_X1 U8771 ( .A1(n11829), .A2(n13317), .ZN(n11828) );
  NAND2_X1 U8772 ( .A1(n12001), .A2(n13202), .ZN(n11829) );
  NAND2_X1 U8773 ( .A1(n11396), .A2(n9283), .ZN(n11694) );
  NAND2_X1 U8774 ( .A1(n13152), .A2(n13151), .ZN(n13924) );
  INV_X1 U8775 ( .A(n13159), .ZN(n13986) );
  INV_X1 U8776 ( .A(n13924), .ZN(n13989) );
  NAND2_X1 U8777 ( .A1(n15732), .A2(n7080), .ZN(n7079) );
  INV_X1 U8778 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n7080) );
  INV_X1 U8779 ( .A(n13427), .ZN(n13997) );
  OR2_X1 U8780 ( .A1(n13150), .A2(n9183), .ZN(n9184) );
  OAI211_X1 U8781 ( .C1(n11910), .C2(n10856), .A(n8951), .B(n8950), .ZN(n12295) );
  OR2_X1 U8782 ( .A1(n8980), .A2(SI_9_), .ZN(n8951) );
  INV_X1 U8783 ( .A(n12030), .ZN(n11945) );
  INV_X1 U8784 ( .A(n11660), .ZN(n11795) );
  AND2_X1 U8785 ( .A1(n9351), .A2(n9350), .ZN(n14034) );
  AND2_X1 U8786 ( .A1(n10855), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14035) );
  OR2_X1 U8787 ( .A1(n14039), .A2(n14040), .ZN(n8786) );
  XNOR2_X1 U8788 ( .A(n8789), .B(n8788), .ZN(n14046) );
  INV_X1 U8789 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8788) );
  INV_X1 U8790 ( .A(n9343), .ZN(n12037) );
  NAND2_X1 U8791 ( .A1(n9339), .A2(n9338), .ZN(n11939) );
  NAND2_X1 U8792 ( .A1(n9140), .A2(n9139), .ZN(n9143) );
  INV_X1 U8793 ( .A(SI_20_), .ZN(n11026) );
  INV_X1 U8794 ( .A(n13666), .ZN(n13679) );
  OAI21_X1 U8795 ( .B1(n9092), .B2(n7389), .A(n7386), .ZN(n9112) );
  NAND2_X1 U8796 ( .A1(n9095), .A2(n9094), .ZN(n9109) );
  NAND2_X1 U8797 ( .A1(n9092), .A2(n9091), .ZN(n9095) );
  NAND2_X1 U8798 ( .A1(n9074), .A2(n9073), .ZN(n9090) );
  INV_X1 U8799 ( .A(SI_16_), .ZN(n10572) );
  INV_X1 U8800 ( .A(SI_15_), .ZN(n10497) );
  NAND2_X1 U8801 ( .A1(n7394), .A2(n9041), .ZN(n9045) );
  INV_X1 U8802 ( .A(SI_14_), .ZN(n10457) );
  NAND2_X1 U8803 ( .A1(n7395), .A2(n9023), .ZN(n9042) );
  INV_X1 U8804 ( .A(SI_12_), .ZN(n10436) );
  INV_X1 U8805 ( .A(SI_11_), .ZN(n10422) );
  INV_X1 U8806 ( .A(SI_10_), .ZN(n10415) );
  OAI21_X1 U8807 ( .B1(n8948), .B2(n7379), .A(n7377), .ZN(n8982) );
  NAND2_X1 U8808 ( .A1(n8959), .A2(n8958), .ZN(n8962) );
  NAND2_X1 U8809 ( .A1(n7066), .A2(n7390), .ZN(n8945) );
  NAND2_X1 U8810 ( .A1(n8901), .A2(n7070), .ZN(n7066) );
  INV_X1 U8811 ( .A(n11896), .ZN(n15649) );
  NAND2_X1 U8812 ( .A1(n8903), .A2(n8902), .ZN(n8906) );
  INV_X1 U8813 ( .A(n11897), .ZN(n15615) );
  NAND2_X1 U8814 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n6933) );
  AND2_X1 U8815 ( .A1(n8630), .A2(n8615), .ZN(n14233) );
  NAND2_X1 U8816 ( .A1(n11446), .A2(n10283), .ZN(n11616) );
  NAND2_X1 U8817 ( .A1(n8400), .A2(n8399), .ZN(n15533) );
  NAND2_X1 U8818 ( .A1(n10248), .A2(n10247), .ZN(n10249) );
  INV_X1 U8819 ( .A(n10245), .ZN(n10248) );
  INV_X1 U8820 ( .A(n10246), .ZN(n10247) );
  NAND2_X1 U8821 ( .A1(n7256), .A2(n7255), .ZN(n12886) );
  AOI21_X1 U8822 ( .B1(n7257), .B2(n14137), .A(n12881), .ZN(n7255) );
  NAND2_X1 U8823 ( .A1(n8366), .A2(n8365), .ZN(n15523) );
  NAND2_X1 U8824 ( .A1(n8590), .A2(n8589), .ZN(n14085) );
  AOI21_X1 U8825 ( .B1(n10308), .B2(n7243), .A(n7242), .ZN(n12497) );
  NAND2_X1 U8826 ( .A1(n8577), .A2(n8576), .ZN(n14430) );
  NAND2_X1 U8827 ( .A1(n14106), .A2(n14105), .ZN(n14104) );
  NAND2_X1 U8828 ( .A1(n12865), .A2(n14057), .ZN(n14106) );
  AND2_X1 U8829 ( .A1(n10899), .A2(n10255), .ZN(n10794) );
  NAND2_X1 U8830 ( .A1(n7260), .A2(n11242), .ZN(n11448) );
  AND2_X1 U8831 ( .A1(n10348), .A2(n10347), .ZN(n14131) );
  NAND2_X1 U8832 ( .A1(n8439), .A2(n8438), .ZN(n12080) );
  OR2_X1 U8833 ( .A1(n10264), .A2(n10265), .ZN(n10266) );
  NAND2_X1 U8834 ( .A1(n10884), .A2(n10263), .ZN(n11234) );
  NAND2_X1 U8835 ( .A1(n7027), .A2(n7026), .ZN(n7258) );
  INV_X1 U8836 ( .A(n14137), .ZN(n7026) );
  NAND2_X1 U8837 ( .A1(n14136), .A2(n14137), .ZN(n7025) );
  XNOR2_X1 U8838 ( .A(n10308), .B(n10309), .ZN(n12402) );
  NAND2_X1 U8839 ( .A1(n10339), .A2(n14387), .ZN(n14146) );
  AOI21_X1 U8840 ( .B1(n10135), .B2(n10134), .A(n10133), .ZN(n7430) );
  OAI21_X1 U8841 ( .B1(n14318), .B2(n8564), .A(n8563), .ZN(n14335) );
  INV_X1 U8842 ( .A(n7098), .ZN(n15364) );
  INV_X1 U8843 ( .A(n7096), .ZN(n15377) );
  NOR2_X1 U8844 ( .A1(n7102), .A2(n7101), .ZN(n7100) );
  INV_X1 U8845 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7101) );
  OAI21_X1 U8846 ( .B1(n11295), .B2(P2_REG2_REG_9__SCAN_IN), .A(n11290), .ZN(
        n15429) );
  NOR2_X1 U8847 ( .A1(n15429), .A2(n15430), .ZN(n15428) );
  NOR2_X1 U8848 ( .A1(n15428), .A2(n7094), .ZN(n11294) );
  AND2_X1 U8849 ( .A1(n15433), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7094) );
  OR2_X1 U8850 ( .A1(n11975), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6836) );
  AND2_X1 U8851 ( .A1(n12211), .A2(n12214), .ZN(n7108) );
  NOR2_X1 U8852 ( .A1(n14193), .A2(n15438), .ZN(n15454) );
  NOR2_X1 U8853 ( .A1(n15452), .A2(n6822), .ZN(n15464) );
  AND2_X1 U8854 ( .A1(n15457), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6822) );
  OR2_X1 U8855 ( .A1(n14203), .A2(n12878), .ZN(n14405) );
  NAND2_X1 U8856 ( .A1(n9864), .A2(n9863), .ZN(n14222) );
  NOR2_X1 U8857 ( .A1(n14238), .A2(n7246), .ZN(n7245) );
  INV_X1 U8858 ( .A(n8608), .ZN(n7246) );
  NAND2_X1 U8859 ( .A1(n8609), .A2(n8608), .ZN(n14239) );
  AND2_X1 U8860 ( .A1(n14281), .A2(n14280), .ZN(n14428) );
  NAND2_X1 U8861 ( .A1(n14333), .A2(n8688), .ZN(n14322) );
  NAND2_X1 U8862 ( .A1(n7230), .A2(n7226), .ZN(n14315) );
  OR2_X1 U8863 ( .A1(n14343), .A2(n14342), .ZN(n7230) );
  NAND2_X1 U8864 ( .A1(n7254), .A2(n8529), .ZN(n14346) );
  NAND2_X1 U8865 ( .A1(n7278), .A2(n7282), .ZN(n12562) );
  NAND2_X1 U8866 ( .A1(n8678), .A2(n7284), .ZN(n7278) );
  NAND2_X1 U8867 ( .A1(n8678), .A2(n8677), .ZN(n12483) );
  NAND2_X1 U8868 ( .A1(n12318), .A2(n8711), .ZN(n12487) );
  NAND2_X1 U8869 ( .A1(n7235), .A2(n7234), .ZN(n12480) );
  AND2_X1 U8870 ( .A1(n7235), .A2(n7237), .ZN(n12481) );
  NAND2_X1 U8871 ( .A1(n7236), .A2(n12374), .ZN(n7235) );
  NAND2_X1 U8872 ( .A1(n7303), .A2(n8672), .ZN(n12074) );
  NAND2_X1 U8873 ( .A1(n12042), .A2(n8671), .ZN(n7303) );
  NAND2_X1 U8874 ( .A1(n11320), .A2(n8350), .ZN(n11270) );
  NAND2_X2 U8875 ( .A1(n8323), .A2(n8322), .ZN(n11019) );
  OR2_X1 U8876 ( .A1(n8464), .A2(n10384), .ZN(n8279) );
  INV_X1 U8877 ( .A(n14202), .ZN(n14489) );
  AND2_X1 U8878 ( .A1(n14439), .A2(n14438), .ZN(n14497) );
  NAND2_X1 U8879 ( .A1(n8416), .A2(n8415), .ZN(n12257) );
  AND2_X1 U8880 ( .A1(n10343), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15512) );
  OAI21_X1 U8881 ( .B1(n8751), .B2(n8750), .A(n8749), .ZN(n15511) );
  INV_X1 U8882 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n6890) );
  INV_X1 U8883 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n12000) );
  NAND2_X1 U8884 ( .A1(n8648), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8644) );
  INV_X1 U8885 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11814) );
  MUX2_X1 U8886 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8647), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n8649) );
  INV_X1 U8887 ( .A(n10077), .ZN(n11708) );
  INV_X1 U8888 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n11023) );
  INV_X1 U8889 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11079) );
  INV_X1 U8890 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n11046) );
  INV_X1 U8891 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10682) );
  INV_X1 U8892 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10583) );
  INV_X1 U8893 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10518) );
  INV_X1 U8894 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10461) );
  INV_X1 U8895 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10453) );
  INV_X1 U8896 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10445) );
  INV_X1 U8897 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10439) );
  INV_X1 U8898 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10427) );
  INV_X1 U8899 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10407) );
  NAND2_X1 U8900 ( .A1(n8293), .A2(n8294), .ZN(n8305) );
  INV_X1 U8901 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10409) );
  XNOR2_X1 U8902 ( .A(n8295), .B(n8294), .ZN(n10978) );
  NAND2_X1 U8903 ( .A1(n11638), .A2(n6705), .ZN(n11642) );
  NAND2_X1 U8904 ( .A1(n7018), .A2(n15179), .ZN(n7017) );
  NAND2_X1 U8905 ( .A1(n7019), .A2(n7022), .ZN(n7018) );
  OR2_X1 U8906 ( .A1(n14533), .A2(n7349), .ZN(n7022) );
  NOR2_X1 U8907 ( .A1(n6686), .A2(n15212), .ZN(n7016) );
  NAND2_X1 U8908 ( .A1(n8129), .A2(n8128), .ZN(n14537) );
  INV_X1 U8909 ( .A(n7326), .ZN(n7004) );
  NAND2_X1 U8910 ( .A1(n7910), .A2(n7909), .ZN(n15225) );
  NAND2_X1 U8911 ( .A1(n14602), .A2(n13064), .ZN(n14539) );
  NOR2_X1 U8912 ( .A1(n10819), .A2(n10818), .ZN(n7003) );
  XNOR2_X1 U8913 ( .A(n11189), .B(n7002), .ZN(n10823) );
  NAND2_X1 U8914 ( .A1(n7332), .A2(n13042), .ZN(n14548) );
  INV_X1 U8915 ( .A(n14546), .ZN(n7332) );
  NAND2_X1 U8916 ( .A1(n8022), .A2(n8021), .ZN(n14928) );
  NAND2_X1 U8917 ( .A1(n12452), .A2(n12451), .ZN(n12539) );
  NAND2_X1 U8918 ( .A1(n8093), .A2(n8092), .ZN(n15017) );
  AOI22_X1 U8919 ( .A1(n11337), .A2(n11338), .B1(n11199), .B2(n11200), .ZN(
        n11345) );
  NAND2_X1 U8920 ( .A1(n14575), .A2(n14576), .ZN(n14574) );
  NAND2_X1 U8921 ( .A1(n15196), .A2(n13021), .ZN(n14575) );
  AOI21_X1 U8922 ( .B1(n7335), .B2(n7337), .A(n6806), .ZN(n7334) );
  INV_X1 U8923 ( .A(n12094), .ZN(n7311) );
  INV_X1 U8924 ( .A(n7312), .ZN(n12095) );
  INV_X1 U8925 ( .A(n7330), .ZN(n7329) );
  OAI21_X1 U8926 ( .B1(n13042), .B2(n7331), .A(n14594), .ZN(n7330) );
  NAND2_X1 U8927 ( .A1(n14548), .A2(n13046), .ZN(n14595) );
  NAND2_X1 U8928 ( .A1(n12539), .A2(n12538), .ZN(n12540) );
  AND2_X1 U8929 ( .A1(n15096), .A2(n10357), .ZN(n15035) );
  NAND2_X1 U8930 ( .A1(n7322), .A2(n7323), .ZN(n14613) );
  AOI21_X1 U8931 ( .B1(n14576), .B2(n7324), .A(n6761), .ZN(n7323) );
  INV_X1 U8932 ( .A(n13021), .ZN(n7324) );
  AOI21_X1 U8933 ( .B1(n11199), .B2(n7321), .A(n7320), .ZN(n7317) );
  INV_X1 U8934 ( .A(n11343), .ZN(n7320) );
  NAND2_X1 U8935 ( .A1(n11350), .A2(n11349), .ZN(n11638) );
  NAND2_X1 U8936 ( .A1(n10828), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15222) );
  OR2_X1 U8937 ( .A1(n10825), .A2(P1_U3086), .ZN(n12843) );
  OR2_X1 U8938 ( .A1(n12758), .A2(n7745), .ZN(n7746) );
  OR2_X1 U8939 ( .A1(n7784), .A2(n10462), .ZN(n7725) );
  INV_X1 U8940 ( .A(n7057), .ZN(n10361) );
  NOR2_X1 U8941 ( .A1(n10474), .A2(n6720), .ZN(n10676) );
  NOR2_X1 U8942 ( .A1(n10566), .A2(n10565), .ZN(n10564) );
  NOR2_X1 U8943 ( .A1(n10522), .A2(n10521), .ZN(n10641) );
  NOR2_X1 U8944 ( .A1(n10519), .A2(n7061), .ZN(n10522) );
  AND2_X1 U8945 ( .A1(n10523), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7061) );
  NOR2_X1 U8946 ( .A1(n10641), .A2(n7060), .ZN(n10645) );
  AND2_X1 U8947 ( .A1(n10642), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7060) );
  NAND2_X1 U8948 ( .A1(n10645), .A2(n10644), .ZN(n10726) );
  AOI21_X1 U8949 ( .B1(n10723), .B2(n10722), .A(n10721), .ZN(n10916) );
  OR2_X1 U8950 ( .A1(n11758), .A2(n11757), .ZN(n11759) );
  AOI211_X1 U8951 ( .C1(n11722), .C2(n11756), .A(n11768), .B(n11724), .ZN(
        n11770) );
  INV_X1 U8952 ( .A(n7051), .ZN(n14745) );
  INV_X1 U8953 ( .A(n14756), .ZN(n14761) );
  AOI211_X1 U8954 ( .C1(n12747), .C2(n14811), .A(n14958), .B(n14778), .ZN(
        n14795) );
  NAND2_X1 U8955 ( .A1(n14801), .A2(n7600), .ZN(n14807) );
  INV_X1 U8956 ( .A(n14622), .ZN(n14841) );
  OAI21_X1 U8957 ( .B1(n14906), .B2(n6687), .A(n6869), .ZN(n14847) );
  INV_X1 U8958 ( .A(n6868), .ZN(n14848) );
  AOI21_X1 U8959 ( .B1(n14906), .B2(n6871), .A(n6687), .ZN(n6868) );
  AND2_X1 U8960 ( .A1(n7577), .A2(n7575), .ZN(n14919) );
  INV_X1 U8961 ( .A(n8015), .ZN(n7575) );
  INV_X1 U8962 ( .A(n7577), .ZN(n14939) );
  NAND2_X1 U8963 ( .A1(n7541), .A2(n8185), .ZN(n14954) );
  NAND2_X1 U8964 ( .A1(n14971), .A2(n14972), .ZN(n7541) );
  NAND2_X1 U8965 ( .A1(n11388), .A2(n12766), .ZN(n7965) );
  NAND2_X1 U8966 ( .A1(n12460), .A2(n8181), .ZN(n12548) );
  NAND2_X1 U8967 ( .A1(n12464), .A2(n12798), .ZN(n12463) );
  NAND2_X1 U8968 ( .A1(n7552), .A2(n7556), .ZN(n12464) );
  NAND2_X1 U8969 ( .A1(n12226), .A2(n7553), .ZN(n7552) );
  NAND2_X1 U8970 ( .A1(n8179), .A2(n12670), .ZN(n12462) );
  NAND2_X1 U8971 ( .A1(n12226), .A2(n7591), .ZN(n12414) );
  NAND2_X1 U8972 ( .A1(n11429), .A2(n7533), .ZN(n11624) );
  NAND2_X1 U8973 ( .A1(n11606), .A2(n12093), .ZN(n11626) );
  NAND2_X1 U8974 ( .A1(n11623), .A2(n12789), .ZN(n11622) );
  NAND2_X1 U8975 ( .A1(n11432), .A2(n7842), .ZN(n11623) );
  NAND2_X1 U8976 ( .A1(n11546), .A2(n11552), .ZN(n11545) );
  NAND2_X1 U8977 ( .A1(n10924), .A2(n7786), .ZN(n11546) );
  AND2_X1 U8978 ( .A1(n11143), .A2(n11142), .ZN(n15277) );
  NAND2_X1 U8979 ( .A1(n7897), .A2(n7896), .ZN(n12662) );
  NAND2_X1 U8980 ( .A1(n7544), .A2(n6879), .ZN(n10228) );
  INV_X1 U8981 ( .A(n6880), .ZN(n6879) );
  OAI21_X1 U8982 ( .B1(n14798), .B2(n15286), .A(n15324), .ZN(n6880) );
  INV_X1 U8983 ( .A(n14537), .ZN(n14826) );
  NAND2_X1 U8984 ( .A1(n8216), .A2(n8215), .ZN(n8255) );
  AOI21_X1 U8985 ( .B1(n12751), .B2(P2_DATAO_REG_4__SCAN_IN), .A(n6721), .ZN(
        n6959) );
  NAND2_X1 U8986 ( .A1(n10423), .A2(n12766), .ZN(n6960) );
  XNOR2_X1 U8987 ( .A(n10049), .B(n10048), .ZN(n14521) );
  OAI22_X1 U8988 ( .A1(n10055), .A2(n10053), .B1(n10045), .B2(n13381), .ZN(
        n10049) );
  INV_X1 U8989 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n12962) );
  NOR2_X1 U8990 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n7545) );
  NAND2_X1 U8991 ( .A1(n8227), .A2(n6748), .ZN(n7546) );
  NOR2_X1 U8992 ( .A1(n7699), .A2(n7548), .ZN(n7547) );
  INV_X1 U8993 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11816) );
  NAND2_X1 U8994 ( .A1(n8145), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8147) );
  INV_X1 U8995 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n11064) );
  INV_X1 U8996 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n11025) );
  INV_X1 U8997 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n11081) );
  INV_X1 U8998 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n11048) );
  AND2_X1 U8999 ( .A1(n7878), .A2(n7892), .ZN(n11712) );
  INV_X1 U9000 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10684) );
  INV_X1 U9001 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10585) );
  INV_X1 U9002 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10516) );
  INV_X1 U9003 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10459) );
  INV_X1 U9004 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10455) );
  INV_X1 U9005 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10447) );
  INV_X1 U9006 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10441) );
  INV_X1 U9007 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10424) );
  INV_X1 U9008 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10404) );
  INV_X1 U9009 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10402) );
  NAND2_X1 U9010 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n7055) );
  INV_X1 U9011 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7617) );
  INV_X1 U9012 ( .A(n7118), .ZN(n9418) );
  XNOR2_X1 U9013 ( .A(n9417), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n15743) );
  INV_X1 U9014 ( .A(n7111), .ZN(n15107) );
  OAI21_X1 U9015 ( .B1(n15744), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6750), .ZN(
        n7111) );
  XNOR2_X1 U9016 ( .A(n9449), .B(n6834), .ZN(n15111) );
  INV_X1 U9017 ( .A(n9450), .ZN(n6834) );
  NOR2_X1 U9018 ( .A1(n15241), .A2(n9465), .ZN(n15245) );
  OAI21_X1 U9019 ( .B1(n7128), .B2(n9472), .A(n7127), .ZN(n15122) );
  NAND2_X1 U9020 ( .A1(n7130), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n7128) );
  NAND2_X1 U9021 ( .A1(n15253), .A2(n7134), .ZN(n7129) );
  AND2_X1 U9022 ( .A1(n7268), .A2(n6719), .ZN(n12331) );
  NAND2_X1 U9023 ( .A1(n6940), .A2(n13655), .ZN(n6939) );
  AND2_X1 U9024 ( .A1(n7400), .A2(n7402), .ZN(n13696) );
  AND2_X1 U9025 ( .A1(n10180), .A2(n10181), .ZN(n13132) );
  NAND2_X1 U9026 ( .A1(n15739), .A2(n9269), .ZN(n7369) );
  NAND2_X1 U9027 ( .A1(n7503), .A2(n7502), .ZN(n10157) );
  NAND2_X1 U9028 ( .A1(n15739), .A2(n10156), .ZN(n7502) );
  NAND2_X1 U9029 ( .A1(n7398), .A2(n7401), .ZN(n9382) );
  OR2_X1 U9030 ( .A1(n15734), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n7401) );
  OAI21_X1 U9031 ( .B1(n7500), .B2(n6932), .A(n6931), .ZN(n10159) );
  NAND2_X1 U9032 ( .A1(n15732), .A2(n10158), .ZN(n6931) );
  NOR2_X1 U9033 ( .A1(n7088), .A2(n6819), .ZN(n7087) );
  NAND2_X1 U9034 ( .A1(n7090), .A2(n11007), .ZN(n7089) );
  AOI21_X1 U9035 ( .B1(n12856), .B2(n15498), .A(n12855), .ZN(n6892) );
  OAI21_X1 U9036 ( .B1(n12854), .B2(n6894), .A(n14397), .ZN(n6893) );
  OR2_X1 U9037 ( .A1(n12857), .A2(n14362), .ZN(n6895) );
  OAI21_X1 U9038 ( .B1(n12853), .B2(n14472), .A(n9839), .ZN(n9840) );
  AOI21_X1 U9039 ( .B1(n10063), .B2(n10162), .A(n10161), .ZN(n10163) );
  NAND2_X1 U9040 ( .A1(n7599), .A2(n8753), .ZN(n8754) );
  OAI21_X1 U9041 ( .B1(n12957), .B2(n10385), .A(n7106), .ZN(P2_U3326) );
  NOR2_X1 U9042 ( .A1(n12959), .A2(n10384), .ZN(n7107) );
  NAND2_X1 U9043 ( .A1(n7342), .A2(n15179), .ZN(n7340) );
  INV_X1 U9044 ( .A(n7050), .ZN(n14734) );
  NAND2_X1 U9045 ( .A1(n6965), .A2(n7597), .ZN(P1_U3557) );
  AOI21_X1 U9046 ( .B1(n7544), .B2(n6962), .A(n6810), .ZN(n6961) );
  OAI21_X1 U9047 ( .B1(n15073), .B2(n10226), .A(n7136), .ZN(n15074) );
  NAND2_X1 U9048 ( .A1(n10226), .A2(n12757), .ZN(n7136) );
  INV_X1 U9049 ( .A(n7112), .ZN(n15112) );
  NOR2_X1 U9050 ( .A1(n15238), .A2(n15237), .ZN(n15236) );
  NOR2_X1 U9051 ( .A1(n9457), .A2(n15234), .ZN(n15238) );
  NOR2_X1 U9052 ( .A1(n15099), .A2(n15100), .ZN(n6835) );
  NOR2_X1 U9053 ( .A1(n7109), .A2(n15100), .ZN(n9834) );
  AND2_X1 U9054 ( .A1(n8696), .A2(n6884), .ZN(n6685) );
  INV_X1 U9055 ( .A(n7592), .ZN(n7171) );
  AND2_X1 U9056 ( .A1(n7019), .A2(n6749), .ZN(n6686) );
  NOR2_X2 U9057 ( .A1(n12577), .A2(n8152), .ZN(n6706) );
  NOR2_X1 U9058 ( .A1(n6711), .A2(n7566), .ZN(n6687) );
  INV_X1 U9059 ( .A(n13326), .ZN(n7515) );
  INV_X1 U9060 ( .A(n14238), .ZN(n7305) );
  INV_X1 U9061 ( .A(n8367), .ZN(n8314) );
  INV_X1 U9062 ( .A(n12803), .ZN(n14866) );
  AND2_X1 U9063 ( .A1(n7138), .A2(n13022), .ZN(n6688) );
  INV_X1 U9064 ( .A(n11190), .ZN(n7002) );
  INV_X1 U9065 ( .A(n7391), .ZN(n7390) );
  OAI21_X1 U9066 ( .B1(n6714), .B2(n7392), .A(n8926), .ZN(n7391) );
  NOR2_X1 U9067 ( .A1(n7182), .A2(n12298), .ZN(n6689) );
  AND2_X1 U9068 ( .A1(n7960), .A2(n7962), .ZN(n6690) );
  AND2_X1 U9069 ( .A1(n7576), .A2(n6863), .ZN(n6691) );
  AND2_X1 U9070 ( .A1(n10154), .A2(n10155), .ZN(n6692) );
  INV_X1 U9071 ( .A(n13099), .ZN(n7349) );
  AND2_X1 U9072 ( .A1(n14415), .A2(n14141), .ZN(n6693) );
  NAND2_X1 U9073 ( .A1(n10195), .A2(n10194), .ZN(n15004) );
  INV_X1 U9074 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10417) );
  AND2_X1 U9075 ( .A1(n7140), .A2(n7139), .ZN(n6694) );
  AND2_X1 U9076 ( .A1(n14475), .A2(n14154), .ZN(n6695) );
  AND2_X1 U9077 ( .A1(n12807), .A2(n8121), .ZN(n6696) );
  AND2_X1 U9078 ( .A1(n13653), .A2(n13660), .ZN(n6697) );
  AND2_X1 U9079 ( .A1(n9023), .A2(n6803), .ZN(n6698) );
  AND2_X1 U9080 ( .A1(n7227), .A2(n14326), .ZN(n6699) );
  INV_X1 U9081 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n7698) );
  INV_X1 U9082 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8265) );
  INV_X1 U9083 ( .A(n13017), .ZN(n15200) );
  AND2_X1 U9084 ( .A1(n7697), .A2(n7696), .ZN(n13017) );
  AND2_X1 U9085 ( .A1(n6986), .A2(n14518), .ZN(n6700) );
  AND2_X1 U9086 ( .A1(n7285), .A2(n8326), .ZN(n6701) );
  NAND2_X1 U9087 ( .A1(n8796), .A2(n8795), .ZN(n13535) );
  NOR2_X1 U9088 ( .A1(n12980), .A2(n12973), .ZN(n6702) );
  INV_X1 U9089 ( .A(n12609), .ZN(n7196) );
  NOR2_X1 U9090 ( .A1(n12667), .A2(n6771), .ZN(n6703) );
  NAND2_X1 U9091 ( .A1(n8566), .A2(n8565), .ZN(n14306) );
  INV_X1 U9092 ( .A(n14306), .ZN(n7227) );
  INV_X1 U9093 ( .A(n10090), .ZN(n7228) );
  INV_X1 U9094 ( .A(n10020), .ZN(n7465) );
  INV_X1 U9095 ( .A(n12482), .ZN(n7283) );
  OR2_X1 U9096 ( .A1(n13817), .A2(n13827), .ZN(n13268) );
  AND2_X1 U9097 ( .A1(n7148), .A2(n9346), .ZN(n9348) );
  AND2_X1 U9098 ( .A1(n8106), .A2(SI_26_), .ZN(n6704) );
  OR2_X1 U9099 ( .A1(n11637), .A2(n11636), .ZN(n6705) );
  INV_X1 U9100 ( .A(n12788), .ZN(n7559) );
  INV_X1 U9101 ( .A(n15237), .ZN(n7121) );
  NAND2_X1 U9102 ( .A1(n14955), .A2(n7578), .ZN(n7577) );
  INV_X1 U9103 ( .A(n7213), .ZN(n10710) );
  OR2_X1 U9104 ( .A1(n8697), .A2(n10077), .ZN(n7213) );
  NOR2_X1 U9105 ( .A1(n9081), .A2(n9068), .ZN(n6707) );
  NAND2_X2 U9106 ( .A1(n7754), .A2(n7753), .ZN(n12593) );
  OR2_X1 U9107 ( .A1(n8783), .A2(n7176), .ZN(n6708) );
  OR2_X1 U9108 ( .A1(n15578), .A2(n11857), .ZN(n6709) );
  INV_X1 U9109 ( .A(n9876), .ZN(n10061) );
  XNOR2_X1 U9110 ( .A(n8147), .B(n8146), .ZN(n8213) );
  NAND2_X1 U9111 ( .A1(n13761), .A2(n10149), .ZN(n10168) );
  AND2_X1 U9112 ( .A1(n7472), .A2(n7276), .ZN(n6710) );
  AND2_X1 U9113 ( .A1(n14866), .A2(n7568), .ZN(n6711) );
  NOR2_X1 U9114 ( .A1(n15123), .A2(n9486), .ZN(n6712) );
  NOR2_X1 U9115 ( .A1(n7957), .A2(SI_17_), .ZN(n6713) );
  AND2_X1 U9116 ( .A1(n7393), .A2(n8902), .ZN(n6714) );
  NAND2_X1 U9117 ( .A1(n12126), .A2(n12155), .ZN(n6715) );
  AND2_X1 U9118 ( .A1(n9909), .A2(n9908), .ZN(n6716) );
  INV_X1 U9119 ( .A(n7436), .ZN(n7435) );
  NAND2_X1 U9120 ( .A1(n7438), .A2(n6802), .ZN(n7436) );
  NAND2_X1 U9121 ( .A1(n9957), .A2(n9972), .ZN(n6717) );
  CLKBUF_X3 U9122 ( .A(n10821), .Z(n13103) );
  OR2_X1 U9123 ( .A1(n14475), .A2(n12405), .ZN(n6718) );
  OR2_X1 U9124 ( .A1(n12328), .A2(n12327), .ZN(n6719) );
  AND2_X1 U9125 ( .A1(n10475), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6720) );
  NAND2_X1 U9126 ( .A1(n8492), .A2(n8491), .ZN(n12565) );
  INV_X1 U9127 ( .A(n12565), .ZN(n14518) );
  NAND2_X1 U9128 ( .A1(n7931), .A2(n7930), .ZN(n13009) );
  INV_X1 U9129 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n9796) );
  INV_X1 U9130 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7288) );
  NAND2_X1 U9131 ( .A1(n13379), .A2(n8794), .ZN(n8916) );
  AND2_X1 U9132 ( .A1(n7986), .A2(n10483), .ZN(n6721) );
  NAND2_X1 U9133 ( .A1(n12769), .A2(n10503), .ZN(n10589) );
  XNOR2_X1 U9134 ( .A(n8768), .B(P3_IR_REG_20__SCAN_IN), .ZN(n9374) );
  INV_X1 U9135 ( .A(n7670), .ZN(n7036) );
  NOR3_X1 U9136 ( .A1(n12682), .A2(n12681), .A3(n12680), .ZN(n6722) );
  INV_X1 U9137 ( .A(n12802), .ZN(n14920) );
  XNOR2_X1 U9138 ( .A(n14415), .B(n14255), .ZN(n14238) );
  INV_X1 U9139 ( .A(n13531), .ZN(n12357) );
  INV_X1 U9140 ( .A(n12622), .ZN(n7207) );
  AND2_X1 U9141 ( .A1(n14443), .A2(n14335), .ZN(n6723) );
  OR2_X1 U9142 ( .A1(n13119), .A2(n7346), .ZN(n6724) );
  AND2_X1 U9143 ( .A1(n10218), .A2(n10217), .ZN(n6725) );
  AND2_X1 U9144 ( .A1(n7161), .A2(n13384), .ZN(n6726) );
  NOR2_X1 U9145 ( .A1(n14299), .A2(n14283), .ZN(n6727) );
  INV_X1 U9146 ( .A(n12801), .ZN(n14892) );
  AND2_X1 U9147 ( .A1(n13191), .A2(n13200), .ZN(n13316) );
  NOR2_X1 U9148 ( .A1(n10046), .A2(n10379), .ZN(n6728) );
  NOR2_X1 U9149 ( .A1(n6676), .A2(n10394), .ZN(n6729) );
  OR2_X1 U9150 ( .A1(n13009), .A2(n15192), .ZN(n12670) );
  INV_X1 U9151 ( .A(n12670), .ZN(n7543) );
  AND2_X1 U9152 ( .A1(n8276), .A2(n7482), .ZN(n6730) );
  AND2_X1 U9153 ( .A1(n6987), .A2(n7227), .ZN(n6731) );
  NAND2_X1 U9154 ( .A1(n8531), .A2(n8530), .ZN(n14454) );
  NAND2_X1 U9155 ( .A1(n8597), .A2(n8596), .ZN(n14420) );
  AND2_X1 U9156 ( .A1(n10200), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6732) );
  XNOR2_X1 U9157 ( .A(n7655), .B(SI_9_), .ZN(n7826) );
  AND2_X1 U9158 ( .A1(n7422), .A2(n7677), .ZN(n6733) );
  AND2_X1 U9159 ( .A1(n8087), .A2(n7428), .ZN(n6734) );
  AND2_X1 U9160 ( .A1(n7501), .A2(n6692), .ZN(n6735) );
  AND2_X1 U9161 ( .A1(n12565), .A2(n14129), .ZN(n6736) );
  NAND2_X1 U9162 ( .A1(n8556), .A2(n8555), .ZN(n14443) );
  AND2_X1 U9163 ( .A1(n10220), .A2(n10219), .ZN(n6737) );
  NAND2_X1 U9164 ( .A1(n14270), .A2(n6996), .ZN(n6999) );
  INV_X1 U9165 ( .A(n7757), .ZN(n7639) );
  XNOR2_X1 U9166 ( .A(n7640), .B(SI_4_), .ZN(n7757) );
  NOR2_X1 U9167 ( .A1(n13607), .A2(n13606), .ZN(n6738) );
  AOI21_X1 U9168 ( .B1(n6715), .B2(n12299), .A(n12298), .ZN(n7181) );
  AND2_X1 U9169 ( .A1(n7230), .A2(n7229), .ZN(n6739) );
  AND2_X1 U9170 ( .A1(n7239), .A2(n14090), .ZN(n6740) );
  NAND2_X1 U9171 ( .A1(n13290), .A2(n9213), .ZN(n13721) );
  NAND2_X1 U9172 ( .A1(n7949), .A2(n7948), .ZN(n14573) );
  INV_X1 U9173 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7522) );
  INV_X1 U9174 ( .A(n7184), .ZN(n7183) );
  AND2_X1 U9175 ( .A1(n12919), .A2(n7160), .ZN(n6741) );
  INV_X1 U9176 ( .A(n12668), .ZN(n12795) );
  AND2_X1 U9177 ( .A1(n12669), .A2(n12666), .ZN(n12668) );
  AND2_X1 U9178 ( .A1(n13737), .A2(n13736), .ZN(n13786) );
  AND2_X1 U9179 ( .A1(n13004), .A2(n7325), .ZN(n6742) );
  INV_X1 U9180 ( .A(n7154), .ZN(n11179) );
  NAND2_X1 U9181 ( .A1(n7155), .A2(n15691), .ZN(n7154) );
  AND2_X1 U9182 ( .A1(n12853), .A2(n14228), .ZN(n6743) );
  NAND2_X1 U9183 ( .A1(n12801), .A2(n8082), .ZN(n6744) );
  NOR2_X1 U9184 ( .A1(n12611), .A2(n14658), .ZN(n6745) );
  AND2_X1 U9185 ( .A1(n7296), .A2(n7293), .ZN(n6746) );
  NOR2_X1 U9186 ( .A1(n14928), .A2(n14646), .ZN(n6747) );
  AND2_X1 U9187 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n6748) );
  AND4_X1 U9188 ( .A1(n8848), .A2(n8847), .A3(n8846), .A4(n8845), .ZN(n9282)
         );
  NAND2_X1 U9189 ( .A1(n14533), .A2(n14621), .ZN(n6749) );
  INV_X1 U9190 ( .A(n7551), .ZN(n7550) );
  OAI21_X1 U9191 ( .B1(n7556), .B2(n8180), .A(n7555), .ZN(n7551) );
  OR2_X1 U9192 ( .A1(n9434), .A2(n9433), .ZN(n6750) );
  AND2_X1 U9193 ( .A1(n12611), .A2(n11346), .ZN(n6751) );
  AND3_X1 U9194 ( .A1(n8812), .A2(n8813), .A3(n7493), .ZN(n6752) );
  NAND2_X1 U9195 ( .A1(n13717), .A2(n15716), .ZN(n6753) );
  NOR2_X1 U9196 ( .A1(n12623), .A2(n14656), .ZN(n6754) );
  AND2_X1 U9197 ( .A1(n7655), .A2(SI_9_), .ZN(n6755) );
  AND2_X1 U9198 ( .A1(n7643), .A2(SI_5_), .ZN(n6756) );
  OR2_X1 U9199 ( .A1(n11655), .A2(n11654), .ZN(n6757) );
  INV_X1 U9200 ( .A(n7378), .ZN(n7377) );
  OAI21_X1 U9201 ( .B1(n8947), .B2(n7379), .A(n8961), .ZN(n7378) );
  AND2_X1 U9202 ( .A1(n10031), .A2(n10030), .ZN(n6758) );
  INV_X1 U9203 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7702) );
  NAND2_X1 U9204 ( .A1(n9383), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n6759) );
  AND2_X1 U9205 ( .A1(n11925), .A2(n11924), .ZN(n6760) );
  AND2_X1 U9206 ( .A1(n13029), .A2(n13028), .ZN(n6761) );
  NAND2_X1 U9207 ( .A1(n14261), .A2(n14263), .ZN(n6762) );
  AND2_X1 U9208 ( .A1(n13110), .A2(n13109), .ZN(n6763) );
  INV_X1 U9209 ( .A(n7614), .ZN(n6922) );
  NOR2_X1 U9210 ( .A1(n9200), .A2(n9199), .ZN(n7614) );
  INV_X1 U9211 ( .A(n7301), .ZN(n7300) );
  OR2_X1 U9212 ( .A1(n8673), .A2(n7302), .ZN(n7301) );
  INV_X1 U9213 ( .A(n7360), .ZN(n7359) );
  AOI21_X1 U9214 ( .B1(n13304), .B2(n7363), .A(n13303), .ZN(n7360) );
  INV_X1 U9215 ( .A(n14953), .ZN(n14956) );
  AND2_X1 U9216 ( .A1(n12691), .A2(n12692), .ZN(n14953) );
  AND2_X1 U9217 ( .A1(n12753), .A2(n12752), .ZN(n15079) );
  INV_X1 U9218 ( .A(n15079), .ZN(n7145) );
  OR2_X1 U9219 ( .A1(n14956), .A2(n7540), .ZN(n6764) );
  NAND2_X1 U9220 ( .A1(n12551), .A2(n8183), .ZN(n14971) );
  AND2_X1 U9221 ( .A1(n10319), .A2(n10320), .ZN(n6765) );
  AND2_X1 U9222 ( .A1(n14972), .A2(n12692), .ZN(n6766) );
  AND2_X1 U9223 ( .A1(n14663), .A2(n14664), .ZN(n6767) );
  AND2_X1 U9224 ( .A1(n9414), .A2(n9415), .ZN(n6768) );
  NOR2_X1 U9225 ( .A1(n7611), .A2(n12482), .ZN(n7234) );
  AND2_X1 U9226 ( .A1(n10181), .A2(n15734), .ZN(n6769) );
  AND2_X1 U9227 ( .A1(n9201), .A2(n9213), .ZN(n6770) );
  AND2_X1 U9228 ( .A1(n12664), .A2(n12665), .ZN(n6771) );
  AND2_X1 U9229 ( .A1(n8529), .A2(n7609), .ZN(n6772) );
  OR2_X1 U9230 ( .A1(n12664), .A2(n12665), .ZN(n6773) );
  AND2_X1 U9231 ( .A1(n13802), .A2(n13270), .ZN(n6774) );
  INV_X1 U9232 ( .A(n13046), .ZN(n7331) );
  AND2_X1 U9233 ( .A1(n7258), .A2(n7025), .ZN(n6775) );
  OR2_X1 U9234 ( .A1(n12451), .A2(n7327), .ZN(n6776) );
  AND2_X1 U9235 ( .A1(n14281), .A2(n8588), .ZN(n6777) );
  OR2_X1 U9236 ( .A1(n7488), .A2(n9991), .ZN(n6778) );
  OR2_X1 U9237 ( .A1(n9893), .A2(n9891), .ZN(n6779) );
  INV_X1 U9238 ( .A(n7276), .ZN(n8424) );
  OR2_X1 U9239 ( .A1(n12727), .A2(n12725), .ZN(n6780) );
  OR2_X1 U9240 ( .A1(n9949), .A2(n9947), .ZN(n6781) );
  OR2_X1 U9241 ( .A1(n9927), .A2(n9925), .ZN(n6782) );
  OR2_X1 U9242 ( .A1(n12750), .A2(n12748), .ZN(n6783) );
  OR2_X1 U9243 ( .A1(n12716), .A2(n12714), .ZN(n6784) );
  OR2_X1 U9244 ( .A1(n12705), .A2(n12703), .ZN(n6785) );
  AND2_X1 U9245 ( .A1(n6867), .A2(n8103), .ZN(n6786) );
  INV_X1 U9246 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n7984) );
  OR2_X1 U9247 ( .A1(n12738), .A2(n12736), .ZN(n6787) );
  AND2_X1 U9248 ( .A1(n6702), .A2(n7150), .ZN(n6788) );
  OR2_X1 U9249 ( .A1(n7196), .A2(n12610), .ZN(n6789) );
  OR2_X1 U9250 ( .A1(n9936), .A2(n9938), .ZN(n6790) );
  OR2_X1 U9251 ( .A1(n12642), .A2(n12644), .ZN(n6791) );
  OR2_X1 U9252 ( .A1(n12621), .A2(n7207), .ZN(n6792) );
  NAND2_X1 U9253 ( .A1(n7481), .A2(n9916), .ZN(n6793) );
  OR2_X1 U9254 ( .A1(n12641), .A2(n15207), .ZN(n6794) );
  INV_X1 U9255 ( .A(n7133), .ZN(n7132) );
  NAND2_X1 U9256 ( .A1(n15252), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n7133) );
  INV_X1 U9257 ( .A(n7294), .ZN(n7293) );
  NAND2_X1 U9258 ( .A1(n7295), .A2(n8683), .ZN(n7294) );
  NAND2_X1 U9259 ( .A1(n12087), .A2(n12088), .ZN(n6795) );
  INV_X1 U9260 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8799) );
  INV_X1 U9261 ( .A(n7784), .ZN(n7763) );
  INV_X1 U9262 ( .A(n12374), .ZN(n7233) );
  INV_X1 U9263 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6849) );
  INV_X1 U9264 ( .A(n13529), .ZN(n13909) );
  AND2_X1 U9265 ( .A1(n12915), .A2(n13842), .ZN(n6796) );
  NAND2_X1 U9266 ( .A1(n12876), .A2(n12875), .ZN(n6797) );
  OAI21_X1 U9267 ( .B1(n12452), .B2(n7327), .A(n7326), .ZN(n13005) );
  NAND4_X1 U9268 ( .A1(n9020), .A2(n9019), .A3(n9018), .A4(n9017), .ZN(n13879)
         );
  INV_X1 U9269 ( .A(n13879), .ZN(n7491) );
  INV_X1 U9270 ( .A(n12882), .ZN(n12877) );
  INV_X1 U9271 ( .A(n14991), .ZN(n7137) );
  AND2_X1 U9272 ( .A1(n12228), .A2(n7138), .ZN(n6798) );
  INV_X1 U9273 ( .A(n12971), .ZN(n13300) );
  NAND2_X1 U9274 ( .A1(n9233), .A2(n9232), .ZN(n12971) );
  AND2_X1 U9275 ( .A1(n9305), .A2(n9303), .ZN(n6799) );
  INV_X1 U9276 ( .A(n15670), .ZN(n11910) );
  AND3_X1 U9277 ( .A1(n7760), .A2(n7571), .A3(n7572), .ZN(n7862) );
  AND2_X1 U9278 ( .A1(n12318), .A2(n6700), .ZN(n6800) );
  INV_X1 U9279 ( .A(n10149), .ZN(n7511) );
  NAND2_X1 U9280 ( .A1(n12913), .A2(n12912), .ZN(n13502) );
  NAND2_X1 U9281 ( .A1(n13383), .A2(n12903), .ZN(n13509) );
  NAND2_X1 U9282 ( .A1(n10199), .A2(n10198), .ZN(n12747) );
  INV_X1 U9283 ( .A(n12747), .ZN(n7144) );
  NOR2_X1 U9284 ( .A1(n14400), .A2(n14375), .ZN(n14347) );
  INV_X1 U9285 ( .A(n10011), .ZN(n7471) );
  NAND2_X1 U9286 ( .A1(n7505), .A2(n7506), .ZN(n9076) );
  NOR2_X1 U9287 ( .A1(n12175), .A2(n7905), .ZN(n6801) );
  INV_X1 U9288 ( .A(n6916), .ZN(n6915) );
  NOR2_X1 U9289 ( .A1(n13798), .A2(n6917), .ZN(n6916) );
  INV_X1 U9290 ( .A(n10016), .ZN(n7467) );
  NAND2_X1 U9291 ( .A1(n14347), .A2(n6989), .ZN(n6990) );
  AND2_X1 U9292 ( .A1(n7606), .A2(n7613), .ZN(n6802) );
  NAND2_X1 U9293 ( .A1(n11048), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n6803) );
  AND2_X1 U9294 ( .A1(n7396), .A2(n9041), .ZN(n6804) );
  AND2_X1 U9295 ( .A1(n10034), .A2(n10033), .ZN(n6805) );
  AND2_X1 U9296 ( .A1(n13071), .A2(n13070), .ZN(n6806) );
  AND2_X1 U9297 ( .A1(n13804), .A2(n13812), .ZN(n6807) );
  OAI21_X1 U9298 ( .B1(n10308), .B2(n7242), .A(n7239), .ZN(n7244) );
  OR2_X1 U9299 ( .A1(n8885), .A2(n8762), .ZN(n6808) );
  NAND2_X1 U9300 ( .A1(n8150), .A2(n7960), .ZN(n6809) );
  INV_X1 U9301 ( .A(n10063), .ZN(n14220) );
  AND2_X1 U9302 ( .A1(n9185), .A2(n9184), .ZN(n14006) );
  INV_X1 U9303 ( .A(n14006), .ZN(n12931) );
  INV_X1 U9304 ( .A(n13838), .ZN(n13857) );
  INV_X1 U9305 ( .A(n15734), .ZN(n15732) );
  INV_X1 U9306 ( .A(n15741), .ZN(n15739) );
  NOR2_X1 U9307 ( .A1(n12789), .A2(n7529), .ZN(n7533) );
  AND2_X1 U9308 ( .A1(n15330), .A2(n10225), .ZN(n6810) );
  INV_X1 U9309 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6991) );
  NAND2_X1 U9310 ( .A1(n7253), .A2(n10289), .ZN(n12014) );
  NAND2_X1 U9311 ( .A1(n7289), .A2(n8264), .ZN(n6811) );
  INV_X1 U9312 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6992) );
  AND2_X1 U9313 ( .A1(n8700), .A2(n8631), .ZN(n12887) );
  OAI21_X1 U9314 ( .B1(n12354), .B2(n7171), .A(n7172), .ZN(n7174) );
  AND2_X1 U9315 ( .A1(n10043), .A2(n14048), .ZN(n6812) );
  NOR2_X1 U9316 ( .A1(n12152), .A2(n7519), .ZN(n6813) );
  AND2_X1 U9317 ( .A1(n11429), .A2(n8170), .ZN(n6814) );
  AND2_X1 U9318 ( .A1(n13655), .A2(n13668), .ZN(n6815) );
  INV_X1 U9319 ( .A(n7611), .ZN(n7237) );
  NAND2_X1 U9320 ( .A1(n15512), .A2(n10338), .ZN(n14387) );
  NAND2_X1 U9321 ( .A1(n7866), .A2(n7865), .ZN(n15217) );
  INV_X1 U9322 ( .A(n15217), .ZN(n7139) );
  INV_X1 U9323 ( .A(n15489), .ZN(n7092) );
  OR2_X1 U9324 ( .A1(n13640), .A2(n13639), .ZN(n6816) );
  NOR2_X1 U9325 ( .A1(n15625), .A2(n11843), .ZN(n6817) );
  AND2_X1 U9326 ( .A1(n14201), .A2(n11708), .ZN(n10347) );
  INV_X1 U9327 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7125) );
  INV_X1 U9328 ( .A(n15286), .ZN(n6966) );
  NOR2_X1 U9329 ( .A1(n11179), .A2(n11165), .ZN(n6818) );
  INV_X1 U9330 ( .A(n7271), .ZN(n6956) );
  NOR2_X1 U9331 ( .A1(n13640), .A2(n13854), .ZN(n7271) );
  INV_X1 U9332 ( .A(n15407), .ZN(n7102) );
  AND2_X1 U9333 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6819) );
  NOR2_X1 U9334 ( .A1(n15567), .A2(n15568), .ZN(n6820) );
  NAND2_X1 U9335 ( .A1(n14688), .A2(n14689), .ZN(n7059) );
  INV_X1 U9336 ( .A(n7267), .ZN(n11217) );
  NAND2_X1 U9337 ( .A1(n11223), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n7267) );
  NOR2_X1 U9338 ( .A1(n8787), .A2(P3_IR_REG_29__SCAN_IN), .ZN(n14039) );
  INV_X1 U9339 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6850) );
  AND2_X1 U9340 ( .A1(n10503), .A2(n10431), .ZN(n11142) );
  INV_X1 U9341 ( .A(n14136), .ZN(n7027) );
  NAND2_X1 U9342 ( .A1(n12864), .A2(n12863), .ZN(n12865) );
  OAI21_X1 U9343 ( .B1(n14118), .B2(n14114), .A(n14115), .ZN(n14077) );
  OAI211_X1 U9344 ( .C1(n14052), .C2(n14051), .A(n14050), .B(n14103), .ZN(
        n14056) );
  NAND2_X1 U9345 ( .A1(n14067), .A2(n14066), .ZN(n14065) );
  NAND2_X1 U9346 ( .A1(n6853), .A2(n7214), .ZN(n14084) );
  AOI21_X1 U9347 ( .B1(n13681), .B2(n15666), .A(n6826), .ZN(n13682) );
  OAI21_X1 U9348 ( .B1(n6722), .B2(n6821), .A(n14953), .ZN(n12694) );
  NAND2_X1 U9349 ( .A1(n7038), .A2(n7667), .ZN(n7890) );
  NOR2_X1 U9350 ( .A1(n15391), .A2(n15390), .ZN(n15389) );
  NAND2_X1 U9351 ( .A1(n10988), .A2(n10987), .ZN(n11290) );
  NOR2_X1 U9352 ( .A1(n15404), .A2(n15403), .ZN(n15402) );
  NOR2_X1 U9353 ( .A1(n15353), .A2(n15352), .ZN(n15351) );
  NAND2_X1 U9354 ( .A1(n11535), .A2(n7093), .ZN(n11537) );
  NAND2_X1 U9355 ( .A1(n7086), .A2(n7085), .ZN(n7084) );
  NAND2_X1 U9356 ( .A1(n11971), .A2(n6836), .ZN(n11972) );
  NOR2_X1 U9357 ( .A1(n15464), .A2(n15463), .ZN(n15462) );
  NOR2_X1 U9358 ( .A1(n15411), .A2(n7099), .ZN(n10988) );
  NAND2_X1 U9359 ( .A1(n11537), .A2(n11538), .ZN(n11971) );
  NAND3_X1 U9360 ( .A1(n7083), .A2(n7089), .A3(n7087), .ZN(P2_U3233) );
  NOR2_X1 U9361 ( .A1(n15462), .A2(n7104), .ZN(n14195) );
  NOR2_X1 U9362 ( .A1(n14173), .A2(n14172), .ZN(n14171) );
  NAND2_X1 U9363 ( .A1(n11294), .A2(n11293), .ZN(n11535) );
  NAND2_X1 U9364 ( .A1(n14199), .A2(n15478), .ZN(n7086) );
  NOR2_X1 U9365 ( .A1(n15413), .A2(n15412), .ZN(n15411) );
  NAND2_X1 U9366 ( .A1(n10995), .A2(n8324), .ZN(n11068) );
  NAND2_X1 U9367 ( .A1(n10846), .A2(n8309), .ZN(n10996) );
  NAND2_X1 U9368 ( .A1(n10745), .A2(n8288), .ZN(n10806) );
  NAND2_X1 U9369 ( .A1(n8337), .A2(n8336), .ZN(n11318) );
  NAND2_X1 U9370 ( .A1(n10847), .A2(n10851), .ZN(n10846) );
  NAND3_X1 U9371 ( .A1(n7472), .A2(n7276), .A3(n7595), .ZN(n8717) );
  NAND2_X1 U9373 ( .A1(n14363), .A2(n8528), .ZN(n7254) );
  NAND2_X1 U9374 ( .A1(n14237), .A2(n8620), .ZN(n8637) );
  XNOR2_X1 U9375 ( .A(n8223), .B(n8222), .ZN(n12123) );
  NAND2_X1 U9376 ( .A1(n7009), .A2(n7008), .ZN(n11927) );
  NOR2_X1 U9377 ( .A1(n10693), .A2(n10692), .ZN(n10699) );
  INV_X1 U9378 ( .A(n12086), .ZN(n7001) );
  NAND2_X1 U9379 ( .A1(n7001), .A2(n6795), .ZN(n7312) );
  NOR2_X1 U9380 ( .A1(n10820), .A2(n7003), .ZN(n10824) );
  NAND2_X1 U9381 ( .A1(n10824), .A2(n10823), .ZN(n11193) );
  NAND2_X1 U9382 ( .A1(n13617), .A2(n13618), .ZN(n13619) );
  NAND2_X1 U9383 ( .A1(n15654), .A2(n15653), .ZN(n15652) );
  NAND2_X1 U9384 ( .A1(n11912), .A2(n11913), .ZN(n12263) );
  NAND2_X1 U9385 ( .A1(n11232), .A2(n10268), .ZN(n11091) );
  OAI22_X1 U9386 ( .A1(n11616), .A2(n11615), .B1(n10285), .B2(n10284), .ZN(
        n11748) );
  INV_X1 U9387 ( .A(n6854), .ZN(n6853) );
  NAND2_X1 U9388 ( .A1(n7875), .A2(n7604), .ZN(n7038) );
  NAND2_X1 U9389 ( .A1(n7028), .A2(n7030), .ZN(n7845) );
  NAND2_X1 U9390 ( .A1(n7417), .A2(n7418), .ZN(n7788) );
  AOI21_X1 U9391 ( .B1(n7042), .B2(n6855), .A(n6765), .ZN(n14067) );
  OAI21_X1 U9392 ( .B1(n12865), .B2(n7217), .A(n12869), .ZN(n6854) );
  OR3_X1 U9393 ( .A1(n13286), .A2(n13285), .A3(n13721), .ZN(n13294) );
  OAI21_X1 U9394 ( .B1(n13242), .B2(n13241), .A(n13267), .ZN(n13249) );
  INV_X1 U9395 ( .A(n13346), .ZN(n13350) );
  NAND2_X1 U9396 ( .A1(n6829), .A2(n13238), .ZN(n13245) );
  OAI22_X1 U9397 ( .A1(n13187), .A2(n13186), .B1(n13185), .B2(n13267), .ZN(
        n13188) );
  AOI211_X1 U9398 ( .C1(n13305), .C2(n13304), .A(n13303), .B(n13302), .ZN(
        n13312) );
  AND2_X2 U9399 ( .A1(n7367), .A2(n7607), .ZN(n7506) );
  OAI21_X1 U9400 ( .B1(n13235), .B2(n13234), .A(n6830), .ZN(n6829) );
  INV_X1 U9401 ( .A(n6831), .ZN(n13276) );
  AOI21_X1 U9402 ( .B1(n13271), .B2(n6774), .A(n6832), .ZN(n6831) );
  NAND2_X1 U9403 ( .A1(n13350), .A2(n13349), .ZN(n13351) );
  NAND2_X1 U9404 ( .A1(n6833), .A2(n9440), .ZN(n9444) );
  NAND2_X1 U9405 ( .A1(n15749), .A2(n15748), .ZN(n6833) );
  NOR2_X1 U9406 ( .A1(n9455), .A2(n9456), .ZN(n15233) );
  XNOR2_X1 U9407 ( .A(n9434), .B(n9433), .ZN(n15744) );
  XNOR2_X1 U9408 ( .A(n6835), .B(n15494), .ZN(SUB_1596_U62) );
  NAND2_X1 U9409 ( .A1(n7129), .A2(n7133), .ZN(n9479) );
  NOR2_X1 U9410 ( .A1(n9464), .A2(n9463), .ZN(n15240) );
  NAND3_X1 U9411 ( .A1(n7120), .A2(n7122), .A3(n7123), .ZN(n9464) );
  NAND2_X1 U9412 ( .A1(n14943), .A2(n15090), .ZN(n14924) );
  OAI22_X1 U9413 ( .A1(n7723), .A2(n10385), .B1(n14672), .B2(n10357), .ZN(
        n6878) );
  NOR2_X1 U9414 ( .A1(n7699), .A2(n7863), .ZN(n7135) );
  NAND2_X1 U9415 ( .A1(n6963), .A2(n6961), .ZN(n6965) );
  NOR2_X2 U9416 ( .A1(n14894), .A2(n14883), .ZN(n14852) );
  NOR2_X4 U9417 ( .A1(n11605), .A2(n12623), .ZN(n11606) );
  NOR2_X4 U9418 ( .A1(n12227), .A2(n15225), .ZN(n12228) );
  XNOR2_X1 U9419 ( .A(n14192), .B(n15437), .ZN(n15439) );
  NAND2_X1 U9420 ( .A1(n7084), .A2(n14201), .ZN(n7083) );
  XNOR2_X1 U9421 ( .A(n14195), .B(n7103), .ZN(n15477) );
  NOR2_X1 U9422 ( .A1(n14191), .A2(n7108), .ZN(n12212) );
  NOR2_X1 U9423 ( .A1(n15402), .A2(n7100), .ZN(n15413) );
  AOI21_X1 U9424 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n15394), .A(n15389), .ZN(
        n15404) );
  NAND2_X1 U9425 ( .A1(n12006), .A2(n12005), .ZN(n12004) );
  NAND2_X1 U9426 ( .A1(n11394), .A2(n9281), .ZN(n11396) );
  INV_X1 U9427 ( .A(n13862), .ZN(n6840) );
  AOI21_X1 U9428 ( .B1(n15730), .B2(n13530), .A(n12392), .ZN(n12524) );
  NAND2_X1 U9429 ( .A1(n7496), .A2(n7494), .ZN(n13783) );
  NAND2_X1 U9430 ( .A1(n7399), .A2(n7371), .ZN(n7370) );
  NAND2_X1 U9431 ( .A1(n7370), .A2(n7369), .ZN(n9371) );
  AND2_X2 U9432 ( .A1(n13189), .A2(n13184), .ZN(n13319) );
  NAND2_X1 U9433 ( .A1(n13894), .A2(n7491), .ZN(n7489) );
  OAI22_X2 U9434 ( .A1(n6840), .A2(n6839), .B1(n13510), .B2(n14028), .ZN(
        n13851) );
  AOI21_X1 U9435 ( .B1(n10109), .B2(n10101), .A(n6841), .ZN(n10135) );
  NAND3_X1 U9436 ( .A1(n14342), .A2(n10090), .A3(n14297), .ZN(n6847) );
  NAND2_X1 U9437 ( .A1(n7431), .A2(n7430), .ZN(n10136) );
  OAI21_X2 U9438 ( .B1(n7624), .B2(n6849), .A(n6848), .ZN(n7625) );
  NAND2_X2 U9439 ( .A1(n12202), .A2(n10307), .ZN(n10308) );
  OAI21_X1 U9440 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n9809), .A(n9399), .ZN(
        n9447) );
  NAND2_X1 U9441 ( .A1(n9461), .A2(n9409), .ZN(n6857) );
  INV_X1 U9442 ( .A(n9480), .ZN(n6858) );
  NAND2_X1 U9443 ( .A1(n15620), .A2(n15619), .ZN(n15618) );
  XNOR2_X2 U9444 ( .A(n6933), .B(n7524), .ZN(n10881) );
  NAND2_X1 U9445 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(n7618), .ZN(n7622) );
  NAND2_X1 U9446 ( .A1(n7118), .A2(n7117), .ZN(n7116) );
  OAI21_X1 U9447 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n9405), .A(n9404), .ZN(
        n9458) );
  NOR2_X1 U9448 ( .A1(n9403), .A2(n6768), .ZN(n9454) );
  NOR2_X1 U9449 ( .A1(n9428), .A2(P1_ADDR_REG_3__SCAN_IN), .ZN(n9386) );
  NOR2_X1 U9450 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n9416), .ZN(n9390) );
  OAI21_X1 U9451 ( .B1(n7134), .B2(n7132), .A(n9478), .ZN(n7131) );
  OAI21_X2 U9452 ( .B1(n9439), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n9398), .ZN(
        n9442) );
  NAND2_X1 U9453 ( .A1(n11480), .A2(n7815), .ZN(n11598) );
  NAND2_X1 U9454 ( .A1(n7558), .A2(n11433), .ZN(n7557) );
  NAND2_X1 U9455 ( .A1(n14957), .A2(n6691), .ZN(n6862) );
  NOR2_X2 U9456 ( .A1(n6977), .A2(n7679), .ZN(n7693) );
  AND2_X2 U9457 ( .A1(n7862), .A2(n7690), .ZN(n7691) );
  INV_X1 U9458 ( .A(n14663), .ZN(n6865) );
  NAND2_X1 U9459 ( .A1(n14906), .A2(n6869), .ZN(n6866) );
  NAND2_X1 U9460 ( .A1(n6786), .A2(n6866), .ZN(n14830) );
  NAND2_X1 U9461 ( .A1(n14906), .A2(n8045), .ZN(n14891) );
  INV_X1 U9462 ( .A(n8045), .ZN(n6872) );
  NAND2_X2 U9463 ( .A1(n8206), .A2(n10214), .ZN(n10357) );
  AND2_X2 U9464 ( .A1(n10224), .A2(n6725), .ZN(n7544) );
  NAND2_X1 U9465 ( .A1(n8658), .A2(n11000), .ZN(n8661) );
  NAND2_X1 U9466 ( .A1(n6881), .A2(n8657), .ZN(n11000) );
  NAND2_X1 U9467 ( .A1(n10850), .A2(n8655), .ZN(n6881) );
  NAND2_X1 U9468 ( .A1(n8695), .A2(n14238), .ZN(n14227) );
  NAND3_X1 U9469 ( .A1(n6895), .A2(n6893), .A3(n6892), .ZN(P2_U3237) );
  INV_X1 U9470 ( .A(n11173), .ZN(n11672) );
  AND3_X2 U9471 ( .A1(n8800), .A2(n8801), .A3(n6674), .ZN(n11173) );
  NAND2_X1 U9472 ( .A1(n7350), .A2(n6900), .ZN(n6897) );
  NAND2_X1 U9473 ( .A1(n6897), .A2(n6898), .ZN(n12390) );
  NAND2_X1 U9474 ( .A1(n13858), .A2(n6905), .ZN(n6903) );
  NAND2_X1 U9475 ( .A1(n6903), .A2(n6904), .ZN(n13832) );
  NAND2_X1 U9476 ( .A1(n13816), .A2(n6910), .ZN(n6907) );
  AND2_X2 U9477 ( .A1(n6770), .A2(n6911), .ZN(n6910) );
  OAI21_X1 U9478 ( .B1(n13912), .B2(n6925), .A(n6923), .ZN(n9040) );
  AND2_X1 U9479 ( .A1(n7177), .A2(n6930), .ZN(n6928) );
  NAND4_X1 U9480 ( .A1(n7506), .A2(n7505), .A3(n7177), .A4(n8763), .ZN(n9337)
         );
  AOI21_X1 U9481 ( .B1(n13654), .B2(n13653), .A(n13652), .ZN(n13661) );
  NAND3_X1 U9482 ( .A1(n13682), .A2(n6939), .A3(n6934), .ZN(P3_U3201) );
  INV_X1 U9483 ( .A(n6935), .ZN(n6934) );
  OAI21_X1 U9484 ( .B1(n6937), .B2(n6697), .A(n6936), .ZN(n6935) );
  NAND3_X1 U9485 ( .A1(n6697), .A2(n13654), .A3(n6815), .ZN(n6936) );
  NOR2_X1 U9486 ( .A1(n15587), .A2(n6950), .ZN(n15609) );
  OAI21_X1 U9487 ( .B1(n15551), .B2(n6951), .A(n6953), .ZN(n11839) );
  OR2_X1 U9488 ( .A1(n13605), .A2(n7271), .ZN(n6955) );
  NAND2_X1 U9489 ( .A1(n14798), .A2(n6964), .ZN(n6963) );
  INV_X1 U9490 ( .A(n6967), .ZN(n14851) );
  AOI21_X2 U9491 ( .B1(n8191), .B2(n6970), .A(n6968), .ZN(n6967) );
  INV_X1 U9492 ( .A(n7526), .ZN(n6972) );
  NAND2_X1 U9493 ( .A1(n6976), .A2(n6974), .ZN(n6973) );
  OAI22_X1 U9494 ( .A1(n11478), .A2(n11481), .B1(n14657), .B2(n11476), .ZN(
        n11600) );
  NAND4_X1 U9495 ( .A1(n6978), .A2(n7960), .A3(n7678), .A4(n8146), .ZN(n6977)
         );
  NAND4_X1 U9496 ( .A1(n7960), .A2(n7678), .A3(n8146), .A4(n7984), .ZN(n8148)
         );
  NAND2_X1 U9497 ( .A1(n6979), .A2(n6980), .ZN(n7539) );
  OR2_X2 U9498 ( .A1(n12460), .A2(n6983), .ZN(n6979) );
  XNOR2_X2 U9499 ( .A(n7135), .B(P1_IR_REG_28__SCAN_IN), .ZN(n8206) );
  NAND3_X1 U9500 ( .A1(n14513), .A2(n6700), .A3(n12318), .ZN(n14400) );
  INV_X1 U9501 ( .A(n6990), .ZN(n14337) );
  INV_X1 U9502 ( .A(n6999), .ZN(n9865) );
  XNOR2_X2 U9503 ( .A(n7000), .B(n8276), .ZN(n8705) );
  NAND2_X2 U9504 ( .A1(n11193), .A2(n11192), .ZN(n11199) );
  OAI21_X2 U9505 ( .B1(n12449), .B2(n7004), .A(n6742), .ZN(n15172) );
  NAND2_X1 U9506 ( .A1(n14593), .A2(n7005), .ZN(n14555) );
  NAND2_X2 U9507 ( .A1(n14555), .A2(n13059), .ZN(n14603) );
  NAND2_X1 U9508 ( .A1(n11350), .A2(n7010), .ZN(n7009) );
  OR2_X1 U9509 ( .A1(n14620), .A2(n7017), .ZN(n7015) );
  NAND3_X1 U9510 ( .A1(n7015), .A2(n7014), .A3(n14538), .ZN(P1_U3214) );
  NAND2_X1 U9511 ( .A1(n14620), .A2(n7016), .ZN(n7014) );
  NAND2_X1 U9512 ( .A1(n14620), .A2(n14621), .ZN(n13100) );
  NAND3_X1 U9513 ( .A1(n7024), .A2(n7619), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n7620) );
  NOR2_X1 U9514 ( .A1(n15493), .A2(n7024), .ZN(n7088) );
  NAND2_X1 U9515 ( .A1(n7803), .A2(n7029), .ZN(n7028) );
  NAND2_X1 U9516 ( .A1(n7875), .A2(n7039), .ZN(n7037) );
  NAND2_X2 U9517 ( .A1(n8469), .A2(n8468), .ZN(n12409) );
  MUX2_X1 U9518 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n8806), .Z(n7640) );
  AND2_X1 U9519 ( .A1(n7057), .A2(n7056), .ZN(n10474) );
  NAND2_X1 U9520 ( .A1(n8901), .A2(n7067), .ZN(n7065) );
  NAND2_X1 U9521 ( .A1(n9062), .A2(n7075), .ZN(n7072) );
  NAND2_X1 U9522 ( .A1(n7072), .A2(n7073), .ZN(n7383) );
  NAND3_X1 U9523 ( .A1(n10180), .A2(n6769), .A3(n10183), .ZN(n7078) );
  NAND3_X1 U9524 ( .A1(n10180), .A2(n10181), .A3(n10183), .ZN(n10187) );
  NAND2_X1 U9525 ( .A1(n7078), .A2(n7079), .ZN(n10186) );
  NAND3_X1 U9526 ( .A1(n9193), .A2(n7081), .A3(n13281), .ZN(n9198) );
  OR2_X2 U9527 ( .A1(n13746), .A2(n13741), .ZN(n9193) );
  OAI21_X1 U9528 ( .B1(n15344), .B2(n10977), .A(n7105), .ZN(n15338) );
  XNOR2_X2 U9529 ( .A(n8278), .B(P2_IR_REG_1__SCAN_IN), .ZN(n15344) );
  MUX2_X1 U9530 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n10962), .S(n15344), .Z(
        n15336) );
  NAND2_X1 U9531 ( .A1(n8518), .A2(n15344), .ZN(n7605) );
  AOI21_X1 U9532 ( .B1(n15344), .B2(P2_STATE_REG_SCAN_IN), .A(n7107), .ZN(
        n7106) );
  INV_X1 U9533 ( .A(n7110), .ZN(n15099) );
  OR2_X2 U9534 ( .A1(n9480), .A2(n15123), .ZN(n9485) );
  NAND2_X1 U9535 ( .A1(n9457), .A2(n7124), .ZN(n7120) );
  NAND2_X1 U9536 ( .A1(n15247), .A2(n7133), .ZN(n7126) );
  NAND2_X1 U9537 ( .A1(n7126), .A2(n7130), .ZN(n7127) );
  NAND2_X1 U9538 ( .A1(n15253), .A2(n15252), .ZN(n15251) );
  OR2_X1 U9539 ( .A1(n15252), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n7134) );
  NAND3_X1 U9540 ( .A1(n6694), .A2(n15117), .A3(n11606), .ZN(n12179) );
  NAND2_X1 U9541 ( .A1(n14839), .A2(n7141), .ZN(n14777) );
  NAND2_X1 U9542 ( .A1(n14839), .A2(n14826), .ZN(n14810) );
  NAND2_X1 U9543 ( .A1(n12037), .A2(n9344), .ZN(n7148) );
  OAI21_X1 U9544 ( .B1(n13432), .B2(n7152), .A(n6788), .ZN(n12986) );
  NAND2_X1 U9545 ( .A1(n12981), .A2(n7151), .ZN(n7150) );
  NAND2_X1 U9546 ( .A1(n12950), .A2(n12981), .ZN(n12974) );
  NAND2_X1 U9547 ( .A1(n13432), .A2(n12977), .ZN(n12950) );
  NAND3_X1 U9548 ( .A1(n7153), .A2(n11168), .A3(n7154), .ZN(n11180) );
  INV_X1 U9549 ( .A(n11165), .ZN(n7153) );
  NAND2_X1 U9550 ( .A1(n12913), .A2(n7157), .ZN(n7156) );
  OAI21_X1 U9551 ( .B1(n12354), .B2(n7169), .A(n7165), .ZN(n13418) );
  OAI21_X1 U9552 ( .B1(n12353), .B2(n7171), .A(n12507), .ZN(n7173) );
  NAND3_X1 U9553 ( .A1(n7506), .A2(n7505), .A3(n8763), .ZN(n8783) );
  NAND2_X1 U9554 ( .A1(n11953), .A2(n6689), .ZN(n7178) );
  NAND2_X1 U9555 ( .A1(n7178), .A2(n7179), .ZN(n12301) );
  NAND2_X1 U9556 ( .A1(n12026), .A2(n13534), .ZN(n7184) );
  NAND2_X1 U9557 ( .A1(n12576), .A2(n7185), .ZN(n12759) );
  OAI211_X1 U9558 ( .C1(n12581), .C2(n12584), .A(n12580), .B(n7186), .ZN(n7187) );
  NAND3_X1 U9559 ( .A1(n6683), .A2(n6767), .A3(n12582), .ZN(n7186) );
  INV_X1 U9560 ( .A(n7187), .ZN(n7189) );
  NAND3_X1 U9561 ( .A1(n7189), .A2(n7608), .A3(n7188), .ZN(n12588) );
  OAI22_X1 U9562 ( .A1(n12581), .A2(n14664), .B1(n6683), .B2(n14663), .ZN(
        n7190) );
  NAND3_X1 U9563 ( .A1(n12661), .A2(n12660), .A3(n6703), .ZN(n7191) );
  NAND2_X1 U9564 ( .A1(n7191), .A2(n7192), .ZN(n12672) );
  NAND2_X1 U9565 ( .A1(n7194), .A2(n6789), .ZN(n12614) );
  NAND3_X1 U9566 ( .A1(n12607), .A2(n12606), .A3(n7195), .ZN(n7194) );
  NAND3_X1 U9567 ( .A1(n12746), .A2(n6783), .A3(n12745), .ZN(n7197) );
  NAND2_X1 U9568 ( .A1(n7197), .A2(n7198), .ZN(n12841) );
  NAND2_X1 U9569 ( .A1(n7199), .A2(n7200), .ZN(n12647) );
  NAND3_X1 U9570 ( .A1(n12640), .A2(n6791), .A3(n12639), .ZN(n7199) );
  NAND2_X1 U9571 ( .A1(n7201), .A2(n7202), .ZN(n12709) );
  NAND3_X1 U9572 ( .A1(n12702), .A2(n6785), .A3(n12701), .ZN(n7201) );
  NAND2_X1 U9573 ( .A1(n7203), .A2(n7204), .ZN(n12719) );
  NAND3_X1 U9574 ( .A1(n12712), .A2(n6784), .A3(n12713), .ZN(n7203) );
  NAND2_X1 U9575 ( .A1(n7205), .A2(n7206), .ZN(n12626) );
  NAND3_X1 U9576 ( .A1(n12619), .A2(n6792), .A3(n12618), .ZN(n7205) );
  NAND2_X1 U9577 ( .A1(n7208), .A2(n7209), .ZN(n12741) );
  NAND3_X1 U9578 ( .A1(n12735), .A2(n6787), .A3(n12734), .ZN(n7208) );
  NAND2_X1 U9579 ( .A1(n7210), .A2(n7211), .ZN(n12730) );
  NAND3_X1 U9580 ( .A1(n12724), .A2(n6780), .A3(n12723), .ZN(n7210) );
  NAND2_X1 U9581 ( .A1(n12605), .A2(n12604), .ZN(n12606) );
  AND4_X4 U9582 ( .A1(n7690), .A2(n7570), .A3(n7760), .A4(n7572), .ZN(n8150)
         );
  NAND2_X1 U9583 ( .A1(n12707), .A2(n12706), .ZN(n12713) );
  NAND2_X2 U9584 ( .A1(n7212), .A2(n14201), .ZN(n10234) );
  NAND2_X1 U9585 ( .A1(n14059), .A2(n7215), .ZN(n7214) );
  NAND2_X1 U9586 ( .A1(n12370), .A2(n7234), .ZN(n7231) );
  NAND2_X1 U9587 ( .A1(n7231), .A2(n7232), .ZN(n12560) );
  INV_X1 U9588 ( .A(n7244), .ZN(n14091) );
  NAND2_X1 U9589 ( .A1(n8609), .A2(n7245), .ZN(n14237) );
  NAND2_X1 U9590 ( .A1(n7247), .A2(n7248), .ZN(n8362) );
  NAND2_X1 U9591 ( .A1(n11318), .A2(n8350), .ZN(n7247) );
  INV_X1 U9592 ( .A(n7249), .ZN(n7248) );
  INV_X1 U9593 ( .A(n8350), .ZN(n7250) );
  NAND2_X1 U9594 ( .A1(n7251), .A2(n8349), .ZN(n11320) );
  NAND2_X1 U9595 ( .A1(n7253), .A2(n7252), .ZN(n12063) );
  NAND2_X1 U9596 ( .A1(n7254), .A2(n6772), .ZN(n8539) );
  NAND2_X1 U9597 ( .A1(n14136), .A2(n7257), .ZN(n7256) );
  NAND3_X1 U9598 ( .A1(n10793), .A2(n10899), .A3(n10255), .ZN(n10792) );
  NAND2_X1 U9599 ( .A1(n10792), .A2(n10259), .ZN(n10885) );
  NAND2_X1 U9600 ( .A1(n7260), .A2(n7259), .ZN(n11446) );
  INV_X1 U9601 ( .A(n8646), .ZN(n8645) );
  NAND2_X1 U9602 ( .A1(n8326), .A2(n8265), .ZN(n8639) );
  INV_X2 U9603 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8294) );
  MUX2_X1 U9604 ( .A(n11224), .B(n15671), .S(P3_IR_REG_0__SCAN_IN), .Z(n11225)
         );
  XNOR2_X2 U9605 ( .A(n7270), .B(P3_IR_REG_2__SCAN_IN), .ZN(n11900) );
  INV_X1 U9606 ( .A(n8263), .ZN(n7290) );
  OAI21_X1 U9607 ( .B1(n8682), .B2(n7294), .A(n7291), .ZN(n14353) );
  INV_X1 U9608 ( .A(n7308), .ZN(n9853) );
  NAND2_X1 U9609 ( .A1(n10507), .A2(n10506), .ZN(n10599) );
  MUX2_X1 U9610 ( .A(n10666), .B(n7315), .S(n10357), .Z(n15274) );
  NAND2_X1 U9611 ( .A1(n11337), .A2(n7318), .ZN(n7316) );
  NAND3_X1 U9612 ( .A1(n14630), .A2(n13018), .A3(n14576), .ZN(n7322) );
  NAND2_X1 U9613 ( .A1(n14546), .A2(n13046), .ZN(n7328) );
  NAND2_X1 U9614 ( .A1(n14603), .A2(n7335), .ZN(n7333) );
  NAND2_X1 U9615 ( .A1(n7333), .A2(n7334), .ZN(n14585) );
  NAND2_X1 U9616 ( .A1(n13100), .A2(n7339), .ZN(n7338) );
  OAI211_X1 U9617 ( .C1(n13100), .C2(n7340), .A(n7338), .B(n13123), .ZN(
        P1_U3220) );
  NAND2_X1 U9618 ( .A1(n12001), .A2(n7352), .ZN(n7350) );
  NAND2_X1 U9619 ( .A1(n13719), .A2(n7358), .ZN(n7357) );
  INV_X2 U9620 ( .A(n9274), .ZN(n11368) );
  NAND2_X2 U9621 ( .A1(n13354), .A2(n13667), .ZN(n8835) );
  XNOR2_X2 U9622 ( .A(n7372), .B(n8799), .ZN(n13667) );
  INV_X1 U9623 ( .A(n8814), .ZN(n8815) );
  NAND2_X1 U9624 ( .A1(n9128), .A2(n9139), .ZN(n7380) );
  NAND2_X1 U9625 ( .A1(n9157), .A2(n9156), .ZN(n9182) );
  NAND2_X1 U9626 ( .A1(n7383), .A2(n7384), .ZN(n9126) );
  NAND2_X1 U9627 ( .A1(n9331), .A2(n13874), .ZN(n7400) );
  NAND3_X1 U9628 ( .A1(n7399), .A2(n7400), .A3(n15734), .ZN(n7398) );
  NAND2_X1 U9629 ( .A1(n9161), .A2(n9202), .ZN(n9203) );
  NAND2_X1 U9630 ( .A1(n7403), .A2(n9159), .ZN(n9160) );
  NAND2_X1 U9631 ( .A1(n9173), .A2(n9172), .ZN(n7403) );
  NAND2_X1 U9632 ( .A1(n7758), .A2(n7416), .ZN(n7417) );
  NAND2_X1 U9633 ( .A1(n7890), .A2(n7424), .ZN(n7423) );
  NAND2_X1 U9634 ( .A1(n7429), .A2(n8123), .ZN(n8126) );
  OAI21_X2 U9635 ( .B1(n7959), .B2(n6713), .A(n7958), .ZN(n8000) );
  OAI21_X1 U9636 ( .B1(n9846), .B2(n9845), .A(n9848), .ZN(n10042) );
  INV_X1 U9637 ( .A(n10034), .ZN(n7456) );
  NAND3_X1 U9638 ( .A1(n7459), .A2(n8293), .A3(n8294), .ZN(n8320) );
  AND3_X2 U9639 ( .A1(n7459), .A2(n8293), .A3(n7457), .ZN(n8326) );
  OAI21_X1 U9640 ( .B1(n10021), .B2(n7464), .A(n7463), .ZN(n10026) );
  INV_X1 U9641 ( .A(n7460), .ZN(n10025) );
  OAI21_X1 U9642 ( .B1(n10012), .B2(n7470), .A(n7469), .ZN(n10015) );
  NAND2_X1 U9643 ( .A1(n7468), .A2(n7466), .ZN(n10014) );
  NAND2_X1 U9644 ( .A1(n10012), .A2(n7469), .ZN(n7468) );
  AND4_X2 U9645 ( .A1(n8514), .A2(n8513), .A3(n8261), .A4(n8260), .ZN(n7472)
         );
  NAND2_X1 U9646 ( .A1(n7473), .A2(n7474), .ZN(n9959) );
  NAND3_X1 U9647 ( .A1(n9946), .A2(n6781), .A3(n9945), .ZN(n7473) );
  NAND2_X1 U9648 ( .A1(n7475), .A2(n7476), .ZN(n9930) );
  NAND3_X1 U9649 ( .A1(n9924), .A2(n6782), .A3(n9923), .ZN(n7475) );
  NAND2_X1 U9650 ( .A1(n7477), .A2(n7478), .ZN(n9941) );
  NAND3_X1 U9651 ( .A1(n9935), .A2(n6790), .A3(n9934), .ZN(n7477) );
  NAND2_X1 U9652 ( .A1(n9914), .A2(n6793), .ZN(n7479) );
  INV_X1 U9653 ( .A(n9915), .ZN(n7481) );
  NAND2_X1 U9654 ( .A1(n8275), .A2(n8276), .ZN(n8267) );
  NAND3_X1 U9655 ( .A1(n9889), .A2(n9890), .A3(n6779), .ZN(n7483) );
  NAND2_X1 U9656 ( .A1(n7483), .A2(n7484), .ZN(n9897) );
  NAND3_X1 U9657 ( .A1(n9990), .A2(n9989), .A3(n6778), .ZN(n7486) );
  NAND2_X1 U9658 ( .A1(n7486), .A2(n7487), .ZN(n9996) );
  INV_X2 U9659 ( .A(n8823), .ZN(n9321) );
  OR2_X1 U9660 ( .A1(n8823), .A2(n10951), .ZN(n7493) );
  NAND2_X1 U9661 ( .A1(n13795), .A2(n7586), .ZN(n7496) );
  XNOR2_X1 U9662 ( .A(n10152), .B(n7504), .ZN(n7498) );
  NAND2_X1 U9663 ( .A1(n7499), .A2(n7501), .ZN(n7503) );
  INV_X2 U9664 ( .A(n8884), .ZN(n7505) );
  NAND2_X1 U9665 ( .A1(n11396), .A2(n7507), .ZN(n11691) );
  NOR2_X1 U9666 ( .A1(n13316), .A2(n7508), .ZN(n7507) );
  NAND2_X1 U9667 ( .A1(n12153), .A2(n7516), .ZN(n7512) );
  NAND2_X1 U9668 ( .A1(n7512), .A2(n7513), .ZN(n12391) );
  AND2_X1 U9669 ( .A1(n12304), .A2(n13210), .ZN(n7519) );
  NAND3_X1 U9670 ( .A1(n8784), .A2(n7522), .A3(n8799), .ZN(n7521) );
  NAND3_X1 U9671 ( .A1(n10417), .A2(n7524), .A3(n8756), .ZN(n8833) );
  NAND4_X1 U9672 ( .A1(n8756), .A2(n7524), .A3(n7523), .A4(n8757), .ZN(n8854)
         );
  NAND3_X1 U9673 ( .A1(n11625), .A2(n8170), .A3(n12788), .ZN(n7530) );
  OAI21_X2 U9674 ( .B1(n8169), .B2(n7532), .A(n7531), .ZN(n11800) );
  NAND2_X2 U9675 ( .A1(n8179), .A2(n7542), .ZN(n12460) );
  AND2_X4 U9676 ( .A1(n12968), .A2(n7708), .ZN(n12754) );
  NAND3_X1 U9677 ( .A1(n7708), .A2(n12968), .A3(P1_REG1_REG_2__SCAN_IN), .ZN(
        n7732) );
  NAND2_X1 U9678 ( .A1(n12754), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7717) );
  NAND2_X1 U9679 ( .A1(n12754), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7726) );
  XNOR2_X2 U9680 ( .A(n10209), .B(n10208), .ZN(n14798) );
  NAND3_X1 U9681 ( .A1(n7692), .A2(n7691), .A3(n7698), .ZN(n7701) );
  NAND3_X1 U9682 ( .A1(n7692), .A2(n7691), .A3(n7545), .ZN(n12961) );
  NAND2_X2 U9683 ( .A1(n7547), .A2(n7546), .ZN(n10214) );
  NAND2_X1 U9684 ( .A1(n7564), .A2(n7563), .ZN(n11479) );
  NAND3_X1 U9685 ( .A1(n10925), .A2(n11552), .A3(n12781), .ZN(n7564) );
  NAND2_X1 U9686 ( .A1(n10925), .A2(n12781), .ZN(n10924) );
  NOR2_X1 U9687 ( .A1(n14890), .A2(n8062), .ZN(n14864) );
  AND2_X1 U9688 ( .A1(n7687), .A2(n7686), .ZN(n7572) );
  AND2_X2 U9689 ( .A1(n7738), .A2(n7688), .ZN(n7760) );
  NAND2_X1 U9690 ( .A1(n14955), .A2(n7997), .ZN(n14940) );
  INV_X1 U9691 ( .A(n7997), .ZN(n7579) );
  NAND2_X1 U9692 ( .A1(n10659), .A2(n10658), .ZN(n10898) );
  INV_X1 U9693 ( .A(n8269), .ZN(n14529) );
  OR2_X1 U9694 ( .A1(n9888), .A2(n9887), .ZN(n9889) );
  NAND2_X1 U9695 ( .A1(n12841), .A2(n12837), .ZN(n12838) );
  NAND2_X1 U9696 ( .A1(n14036), .A2(n11160), .ZN(n11158) );
  NAND2_X1 U9697 ( .A1(n11162), .A2(n11161), .ZN(n11164) );
  NAND2_X1 U9698 ( .A1(n11158), .A2(n9374), .ZN(n11162) );
  NAND2_X1 U9699 ( .A1(n8637), .A2(n8696), .ZN(n9844) );
  AND2_X1 U9700 ( .A1(n12937), .A2(n13788), .ZN(n12934) );
  INV_X1 U9701 ( .A(n14958), .ZN(n10508) );
  INV_X1 U9702 ( .A(n10595), .ZN(n10596) );
  NAND2_X1 U9703 ( .A1(n8221), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8223) );
  AOI21_X2 U9704 ( .B1(n12560), .B2(n12561), .A(n8499), .ZN(n14384) );
  XNOR2_X1 U9705 ( .A(n8144), .B(P1_IR_REG_21__SCAN_IN), .ZN(n8198) );
  OAI211_X2 U9706 ( .C1(n10417), .C2(n10856), .A(n8810), .B(n8809), .ZN(n9274)
         );
  NAND4_X4 U9707 ( .A1(n8274), .A2(n8273), .A3(n8272), .A4(n8271), .ZN(n14170)
         );
  OR2_X1 U9708 ( .A1(n8823), .A2(n11678), .ZN(n8791) );
  AND2_X2 U9709 ( .A1(n8198), .A2(n8213), .ZN(n12577) );
  NAND2_X1 U9710 ( .A1(n8150), .A2(n7693), .ZN(n8227) );
  AND2_X1 U9711 ( .A1(n8141), .A2(n8197), .ZN(n8142) );
  OR2_X2 U9712 ( .A1(n10589), .A2(n10508), .ZN(n10697) );
  AND2_X1 U9713 ( .A1(n7596), .A2(n9870), .ZN(n7580) );
  AND2_X2 U9714 ( .A1(n9836), .A2(n9835), .ZN(n15550) );
  NAND2_X2 U9715 ( .A1(n8835), .A2(n10046), .ZN(n8980) );
  NAND2_X1 U9716 ( .A1(n11181), .A2(n11182), .ZN(n11281) );
  AND2_X1 U9717 ( .A1(n8841), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n7581) );
  INV_X1 U9718 ( .A(n8841), .ZN(n9030) );
  INV_X1 U9719 ( .A(n15703), .ZN(n13921) );
  INV_X1 U9720 ( .A(n13983), .ZN(n10189) );
  OR2_X1 U9721 ( .A1(n13692), .A2(n13983), .ZN(n7582) );
  OR2_X1 U9722 ( .A1(n13715), .A2(n13983), .ZN(n7583) );
  OR2_X1 U9723 ( .A1(n13715), .A2(n14033), .ZN(n7584) );
  OR2_X1 U9724 ( .A1(n13692), .A2(n14033), .ZN(n7585) );
  AND2_X1 U9725 ( .A1(n13798), .A2(n9298), .ZN(n7586) );
  INV_X1 U9726 ( .A(n14965), .ZN(n7996) );
  AND2_X1 U9727 ( .A1(n8699), .A2(n8698), .ZN(n14395) );
  INV_X1 U9728 ( .A(n14395), .ZN(n14358) );
  AND3_X1 U9729 ( .A1(n7995), .A2(n7994), .A3(n7993), .ZN(n14597) );
  AND2_X1 U9730 ( .A1(n10300), .A2(n10299), .ZN(n7587) );
  OR2_X1 U9731 ( .A1(n12155), .A2(n11945), .ZN(n7588) );
  OR2_X1 U9732 ( .A1(n14826), .A2(n15046), .ZN(n7589) );
  OR2_X1 U9733 ( .A1(n14826), .A2(n15089), .ZN(n7590) );
  OR2_X1 U9734 ( .A1(n12505), .A2(n12526), .ZN(n7592) );
  OR2_X1 U9735 ( .A1(n9861), .A2(n14204), .ZN(n7594) );
  AND3_X1 U9736 ( .A1(n8642), .A2(n8262), .A3(n8643), .ZN(n7595) );
  OR2_X1 U9737 ( .A1(n14220), .A2(n14472), .ZN(n7596) );
  OR2_X1 U9738 ( .A1(n7144), .A2(n15046), .ZN(n7597) );
  OR2_X1 U9739 ( .A1(n7144), .A2(n15089), .ZN(n7598) );
  OR2_X1 U9740 ( .A1(n12853), .A2(n14517), .ZN(n7599) );
  OR2_X1 U9741 ( .A1(n14800), .A2(n14799), .ZN(n7600) );
  NAND4_X1 U9742 ( .A1(n8782), .A2(n8781), .A3(n8780), .A4(n8779), .ZN(n7601)
         );
  INV_X1 U9743 ( .A(n14893), .ZN(n14909) );
  INV_X1 U9744 ( .A(n15035), .ZN(n14915) );
  AND2_X1 U9745 ( .A1(n12814), .A2(n12815), .ZN(n7602) );
  INV_X1 U9746 ( .A(n14850), .ZN(n8102) );
  INV_X1 U9747 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9383) );
  INV_X1 U9748 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n8217) );
  INV_X1 U9749 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9384) );
  NOR2_X1 U9750 ( .A1(n14271), .A2(n14270), .ZN(n7603) );
  AND2_X1 U9751 ( .A1(n7667), .A2(n7666), .ZN(n7604) );
  INV_X1 U9752 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n8931) );
  OR2_X1 U9753 ( .A1(n6677), .A2(n11007), .ZN(n14214) );
  NAND2_X1 U9754 ( .A1(n15543), .A2(n15532), .ZN(n14517) );
  OR2_X1 U9755 ( .A1(n8029), .A2(SI_20_), .ZN(n7606) );
  INV_X1 U9756 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n9389) );
  AND4_X1 U9757 ( .A1(n8760), .A2(n8759), .A3(n9007), .A4(n8978), .ZN(n7607)
         );
  OR2_X1 U9758 ( .A1(n12586), .A2(n12585), .ZN(n7608) );
  INV_X1 U9759 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8862) );
  OR2_X1 U9760 ( .A1(n14454), .A2(n14370), .ZN(n7609) );
  INV_X1 U9761 ( .A(n14454), .ZN(n8712) );
  OR2_X1 U9762 ( .A1(n8835), .A2(n11900), .ZN(n7610) );
  NOR2_X1 U9763 ( .A1(n12409), .A2(n14155), .ZN(n7611) );
  INV_X1 U9764 ( .A(n12409), .ZN(n8711) );
  AND2_X1 U9765 ( .A1(n9961), .A2(n9960), .ZN(n7612) );
  OR2_X1 U9766 ( .A1(n8031), .A2(SI_21_), .ZN(n7613) );
  AND3_X1 U9767 ( .A1(n9192), .A2(n9191), .A3(n9190), .ZN(n13788) );
  INV_X1 U9768 ( .A(n13788), .ZN(n9301) );
  AND2_X1 U9769 ( .A1(n11280), .A2(n11282), .ZN(n7615) );
  AND2_X2 U9770 ( .A1(n8254), .A2(n8253), .ZN(n15324) );
  INV_X1 U9771 ( .A(n15324), .ZN(n10226) );
  AND3_X2 U9772 ( .A1(n11140), .A2(n8253), .A3(n11137), .ZN(n15332) );
  INV_X1 U9773 ( .A(n9880), .ZN(n9881) );
  OR2_X1 U9774 ( .A1(n9897), .A2(n9896), .ZN(n9898) );
  AND2_X1 U9775 ( .A1(n12688), .A2(n12687), .ZN(n12689) );
  NOR2_X1 U9776 ( .A1(n7612), .A2(n6717), .ZN(n9958) );
  NAND2_X1 U9777 ( .A1(n12722), .A2(n12721), .ZN(n12723) );
  INV_X1 U9778 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8761) );
  INV_X1 U9779 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8262) );
  OR2_X1 U9780 ( .A1(n9273), .A2(n11178), .ZN(n9276) );
  INV_X1 U9781 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7681) );
  INV_X1 U9782 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7619) );
  INV_X1 U9783 ( .A(n12295), .ZN(n9286) );
  NAND2_X1 U9784 ( .A1(n9189), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8824) );
  INV_X1 U9785 ( .A(n10809), .ZN(n10076) );
  INV_X1 U9786 ( .A(n12593), .ZN(n7755) );
  OR2_X1 U9787 ( .A1(n15217), .A2(n14653), .ZN(n7874) );
  AND2_X1 U9788 ( .A1(n7682), .A2(n7681), .ZN(n7683) );
  INV_X1 U9789 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n13441) );
  OR2_X1 U9790 ( .A1(n9309), .A2(n9308), .ZN(n10166) );
  INV_X1 U9791 ( .A(n13760), .ZN(n9305) );
  INV_X1 U9792 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n9635) );
  INV_X1 U9793 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8763) );
  NOR2_X1 U9794 ( .A1(n8470), .A2(n12403), .ZN(n8482) );
  INV_X1 U9795 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8428) );
  NAND2_X1 U9796 ( .A1(n11374), .A2(n11375), .ZN(n11373) );
  INV_X1 U9797 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8276) );
  NAND2_X1 U9798 ( .A1(n11191), .A2(n7002), .ZN(n11192) );
  NOR2_X1 U9799 ( .A1(n10503), .A2(n10504), .ZN(n10505) );
  INV_X1 U9800 ( .A(n12807), .ZN(n8197) );
  NAND2_X1 U9801 ( .A1(n11583), .A2(n8157), .ZN(n8159) );
  INV_X1 U9802 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9594) );
  INV_X1 U9803 ( .A(n7826), .ZN(n7654) );
  NAND2_X1 U9804 ( .A1(n7620), .A2(n14769), .ZN(n7621) );
  INV_X1 U9805 ( .A(n14046), .ZN(n8794) );
  AND2_X1 U9806 ( .A1(n9250), .A2(n13367), .ZN(n13690) );
  AND2_X1 U9807 ( .A1(n10167), .A2(n10166), .ZN(n10173) );
  NAND2_X1 U9808 ( .A1(n13745), .A2(n10150), .ZN(n13722) );
  INV_X1 U9809 ( .A(n14034), .ZN(n11359) );
  OR2_X1 U9810 ( .A1(n8980), .A2(SI_11_), .ZN(n8985) );
  INV_X1 U9811 ( .A(n11235), .ZN(n10267) );
  OR2_X1 U9812 ( .A1(n8369), .A2(n8368), .ZN(n8385) );
  NAND2_X1 U9813 ( .A1(n10246), .A2(n10245), .ZN(n10255) );
  INV_X1 U9814 ( .A(n12016), .ZN(n10295) );
  OR2_X1 U9815 ( .A1(n8630), .A2(n8629), .ZN(n8700) );
  NAND2_X1 U9816 ( .A1(n8493), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8507) );
  OR2_X1 U9817 ( .A1(n8507), .A2(n8506), .ZN(n8522) );
  INV_X1 U9818 ( .A(n14166), .ZN(n8659) );
  NAND2_X1 U9819 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n8096), .ZN(n8113) );
  INV_X1 U9820 ( .A(n8036), .ZN(n8037) );
  INV_X1 U9821 ( .A(n13376), .ZN(n7708) );
  INV_X1 U9822 ( .A(n14642), .ZN(n13113) );
  NAND2_X1 U9823 ( .A1(n8077), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8095) );
  INV_X1 U9824 ( .A(n13009), .ZN(n8211) );
  OR2_X1 U9825 ( .A1(n7809), .A2(n7808), .ZN(n7836) );
  INV_X1 U9826 ( .A(n14809), .ZN(n14799) );
  OR2_X1 U9827 ( .A1(n12653), .A2(n14652), .ZN(n7887) );
  OR2_X1 U9828 ( .A1(n12641), .A2(n14654), .ZN(n7858) );
  OR2_X1 U9829 ( .A1(n12608), .A2(n14659), .ZN(n7786) );
  NAND2_X1 U9830 ( .A1(n14663), .A2(n15295), .ZN(n8155) );
  NAND2_X1 U9831 ( .A1(n8126), .A2(n8125), .ZN(n8623) );
  INV_X1 U9832 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9605) );
  OAI21_X1 U9833 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n9407), .A(n9406), .ZN(
        n9461) );
  OR2_X1 U9834 ( .A1(n13150), .A2(n12310), .ZN(n9232) );
  AND2_X1 U9835 ( .A1(n12977), .A2(n12948), .ZN(n13430) );
  NAND2_X1 U9836 ( .A1(n11570), .A2(n6679), .ZN(n11571) );
  OR2_X1 U9837 ( .A1(n13150), .A2(n12150), .ZN(n9219) );
  AND2_X1 U9838 ( .A1(n11525), .A2(n9271), .ZN(n13702) );
  AOI21_X1 U9839 ( .B1(P3_REG2_REG_2__SCAN_IN), .B2(n11835), .A(n11834), .ZN(
        n11836) );
  AND2_X1 U9840 ( .A1(n11837), .A2(n11902), .ZN(n11838) );
  INV_X1 U9841 ( .A(n15674), .ZN(n15591) );
  AND2_X1 U9842 ( .A1(n10857), .A2(n10856), .ZN(n10866) );
  OR2_X1 U9843 ( .A1(n13150), .A2(n11937), .ZN(n9162) );
  INV_X1 U9844 ( .A(n13332), .ZN(n13847) );
  AND4_X1 U9845 ( .A1(n9087), .A2(n9086), .A3(n9085), .A4(n9084), .ZN(n13828)
         );
  AND2_X1 U9846 ( .A1(n9289), .A2(n9037), .ZN(n13883) );
  AND2_X1 U9847 ( .A1(n11362), .A2(n11361), .ZN(n11363) );
  INV_X1 U9848 ( .A(n11501), .ZN(n15698) );
  OR2_X1 U9849 ( .A1(n13684), .A2(n13683), .ZN(n13984) );
  OR2_X1 U9850 ( .A1(n13150), .A2(n12038), .ZN(n9205) );
  OR2_X1 U9851 ( .A1(n13150), .A2(n11408), .ZN(n9174) );
  INV_X1 U9852 ( .A(n10856), .ZN(n9114) );
  INV_X1 U9853 ( .A(n13874), .ZN(n15696) );
  AND2_X1 U9854 ( .A1(n11084), .A2(n11110), .ZN(n9380) );
  INV_X1 U9855 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n8785) );
  AND2_X1 U9856 ( .A1(n9125), .A2(n9110), .ZN(n9111) );
  AND2_X1 U9857 ( .A1(n8851), .A2(n8832), .ZN(n8849) );
  INV_X1 U9858 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n11094) );
  NAND2_X1 U9859 ( .A1(n10255), .A2(n10249), .ZN(n10901) );
  INV_X1 U9860 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10891) );
  INV_X1 U9861 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n11303) );
  INV_X1 U9862 ( .A(n8713), .ZN(n10142) );
  AND2_X1 U9863 ( .A1(n8557), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8567) );
  OR2_X1 U9864 ( .A1(n8522), .A2(n8521), .ZN(n8544) );
  OR2_X1 U9865 ( .A1(n11531), .A2(n11532), .ZN(n11977) );
  NAND2_X1 U9866 ( .A1(n9854), .A2(n14358), .ZN(n9864) );
  INV_X1 U9867 ( .A(n14347), .ZN(n14374) );
  NAND2_X1 U9868 ( .A1(n14397), .A2(n11008), .ZN(n15503) );
  OR2_X1 U9869 ( .A1(n15543), .A2(n8752), .ZN(n8753) );
  INV_X1 U9870 ( .A(n14155), .ZN(n12485) );
  INV_X1 U9871 ( .A(n11783), .ZN(n12113) );
  OR2_X1 U9872 ( .A1(n8516), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n8476) );
  NOR2_X2 U9873 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n8293) );
  NAND2_X1 U9874 ( .A1(n7899), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7912) );
  OR2_X1 U9875 ( .A1(n7990), .A2(n7989), .ZN(n8010) );
  INV_X1 U9876 ( .A(n14615), .ZN(n15205) );
  NAND2_X1 U9877 ( .A1(n12774), .A2(n7602), .ZN(n12840) );
  INV_X1 U9878 ( .A(n7744), .ZN(n7992) );
  NOR2_X1 U9879 ( .A1(n11716), .A2(n11717), .ZN(n11758) );
  NAND2_X1 U9880 ( .A1(n14803), .A2(n14974), .ZN(n14804) );
  NAND2_X1 U9881 ( .A1(n14908), .A2(n14907), .ZN(n14906) );
  INV_X1 U9882 ( .A(n12794), .ZN(n12553) );
  NAND2_X1 U9883 ( .A1(n14913), .A2(n11147), .ZN(n14949) );
  OR2_X1 U9884 ( .A1(n10500), .A2(P1_D_REG_0__SCAN_IN), .ZN(n8249) );
  AND2_X1 U9885 ( .A1(n8213), .A2(n14764), .ZN(n8251) );
  INV_X1 U9886 ( .A(n12632), .ZN(n12093) );
  INV_X1 U9887 ( .A(n12785), .ZN(n11599) );
  OR2_X1 U9888 ( .A1(n12771), .A2(n10465), .ZN(n14871) );
  XNOR2_X1 U9889 ( .A(n8066), .B(SI_22_), .ZN(n8554) );
  AND2_X1 U9890 ( .A1(n11108), .A2(n11107), .ZN(n11278) );
  AOI21_X1 U9891 ( .B1(n13708), .B2(n9265), .A(n9255), .ZN(n10177) );
  INV_X1 U9892 ( .A(n13827), .ZN(n12923) );
  INV_X1 U9893 ( .A(n15583), .ZN(n15677) );
  NAND2_X1 U9894 ( .A1(n9080), .A2(n9079), .ZN(n13967) );
  NAND2_X1 U9895 ( .A1(n9375), .A2(n13166), .ZN(n13874) );
  INV_X1 U9896 ( .A(n13913), .ZN(n13901) );
  INV_X1 U9897 ( .A(n15702), .ZN(n13914) );
  AND2_X1 U9898 ( .A1(n9368), .A2(n9367), .ZN(n9369) );
  INV_X1 U9899 ( .A(n15719), .ZN(n15731) );
  INV_X1 U9900 ( .A(n15726), .ZN(n15724) );
  INV_X1 U9901 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8978) );
  OR2_X1 U9902 ( .A1(n10538), .A2(n10537), .ZN(n10543) );
  AND2_X1 U9903 ( .A1(n8546), .A2(n8545), .ZN(n14339) );
  INV_X1 U9904 ( .A(n14148), .ZN(n14103) );
  NAND2_X1 U9905 ( .A1(n10553), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14140) );
  NOR2_X1 U9906 ( .A1(n10341), .A2(n15514), .ZN(n10348) );
  AND2_X1 U9907 ( .A1(n8575), .A2(n8574), .ZN(n14326) );
  INV_X1 U9908 ( .A(n8582), .ZN(n8564) );
  NAND2_X1 U9909 ( .A1(n10539), .A2(n10540), .ZN(n15461) );
  INV_X1 U9910 ( .A(n15461), .ZN(n15478) );
  INV_X1 U9911 ( .A(n10088), .ZN(n14354) );
  INV_X1 U9912 ( .A(n14214), .ZN(n15498) );
  NAND2_X1 U9913 ( .A1(n10709), .A2(n14387), .ZN(n14397) );
  INV_X1 U9914 ( .A(n14517), .ZN(n10162) );
  AND2_X1 U9915 ( .A1(n8748), .A2(n15513), .ZN(n9836) );
  AND2_X1 U9916 ( .A1(n8729), .A2(n8750), .ZN(n15508) );
  AND2_X1 U9917 ( .A1(n15183), .A2(n14974), .ZN(n14587) );
  AND2_X1 U9918 ( .A1(n7867), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7881) );
  AND2_X1 U9919 ( .A1(n10827), .A2(n11142), .ZN(n14627) );
  INV_X1 U9920 ( .A(n15212), .ZN(n15179) );
  OR2_X1 U9921 ( .A1(n10203), .A2(n14837), .ZN(n8117) );
  AND4_X1 U9922 ( .A1(n7715), .A2(n7714), .A3(n7713), .A4(n7712), .ZN(n14579)
         );
  AND2_X1 U9923 ( .A1(n10470), .A2(n10362), .ZN(n14762) );
  NAND2_X1 U9924 ( .A1(n14805), .A2(n14804), .ZN(n14806) );
  INV_X1 U9925 ( .A(n12797), .ZN(n12413) );
  INV_X1 U9926 ( .A(n14958), .ZN(n15049) );
  INV_X1 U9927 ( .A(n14949), .ZN(n14992) );
  AND2_X1 U9928 ( .A1(n8249), .A2(n10430), .ZN(n11137) );
  AND2_X1 U9929 ( .A1(n12763), .A2(n12576), .ZN(n15286) );
  NAND2_X1 U9930 ( .A1(n11145), .A2(n10223), .ZN(n15321) );
  NAND2_X1 U9931 ( .A1(n8236), .A2(n8235), .ZN(n10500) );
  AND2_X1 U9932 ( .A1(n7846), .A2(n7831), .ZN(n10909) );
  AND2_X1 U9933 ( .A1(n10868), .A2(n10867), .ZN(n15674) );
  AND2_X1 U9934 ( .A1(n11278), .A2(n13359), .ZN(n13518) );
  AOI21_X1 U9935 ( .B1(n13353), .B2(n13352), .A(n13351), .ZN(n13360) );
  INV_X1 U9936 ( .A(n13723), .ZN(n13763) );
  INV_X1 U9937 ( .A(n13864), .ZN(n13843) );
  INV_X1 U9938 ( .A(n15666), .ZN(n15595) );
  OR2_X1 U9939 ( .A1(n10869), .A2(n10864), .ZN(n15681) );
  INV_X1 U9940 ( .A(n13919), .ZN(n13905) );
  NAND2_X1 U9941 ( .A1(n12971), .A2(n10189), .ZN(n10190) );
  NAND2_X1 U9942 ( .A1(n15741), .A2(n15731), .ZN(n13983) );
  AND2_X2 U9943 ( .A1(n11364), .A2(n9369), .ZN(n15741) );
  NAND2_X1 U9944 ( .A1(n12971), .A2(n10184), .ZN(n10185) );
  INV_X1 U9945 ( .A(n13521), .ZN(n14028) );
  AND2_X2 U9946 ( .A1(n9381), .A2(n11118), .ZN(n15734) );
  CLKBUF_X1 U9947 ( .A(n10610), .Z(n10628) );
  INV_X1 U9948 ( .A(SI_18_), .ZN(n10739) );
  INV_X1 U9949 ( .A(SI_13_), .ZN(n10449) );
  CLKBUF_X1 U9950 ( .A(n14049), .Z(n13382) );
  INV_X1 U9951 ( .A(n14146), .ZN(n14102) );
  NAND2_X1 U9952 ( .A1(n10348), .A2(n10333), .ZN(n14148) );
  INV_X1 U9953 ( .A(n14326), .ZN(n14152) );
  INV_X1 U9954 ( .A(n15484), .ZN(n15465) );
  INV_X1 U9955 ( .A(n15333), .ZN(n15493) );
  INV_X1 U9956 ( .A(n9840), .ZN(n9841) );
  INV_X1 U9957 ( .A(n15550), .ZN(n15548) );
  INV_X1 U9958 ( .A(n14085), .ZN(n14495) );
  INV_X1 U9959 ( .A(n14390), .ZN(n14513) );
  AND2_X2 U9960 ( .A1(n9836), .A2(n15511), .ZN(n15543) );
  INV_X1 U9961 ( .A(n15543), .ZN(n15541) );
  OR2_X1 U9962 ( .A1(n15514), .A2(n15508), .ZN(n15509) );
  INV_X1 U9963 ( .A(n15512), .ZN(n15514) );
  INV_X1 U9964 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n12167) );
  INV_X1 U9965 ( .A(n8650), .ZN(n14201) );
  INV_X1 U9966 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10764) );
  INV_X1 U9967 ( .A(n15271), .ZN(n14737) );
  INV_X1 U9968 ( .A(n12662), .ZN(n12663) );
  NAND2_X1 U9969 ( .A1(n10511), .A2(n10510), .ZN(n15212) );
  OR2_X1 U9970 ( .A1(n7972), .A2(n7971), .ZN(n14648) );
  OR2_X1 U9971 ( .A1(n10503), .A2(n10232), .ZN(n14640) );
  INV_X1 U9972 ( .A(n14762), .ZN(n15266) );
  INV_X1 U9973 ( .A(n14944), .ZN(n14988) );
  INV_X1 U9974 ( .A(n15332), .ZN(n15330) );
  INV_X1 U9975 ( .A(n14928), .ZN(n15090) );
  AND2_X1 U9976 ( .A1(n10354), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10431) );
  INV_X1 U9977 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11389) );
  INV_X1 U9978 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10817) );
  XNOR2_X1 U9979 ( .A(n9832), .B(n9831), .ZN(n9833) );
  INV_X1 U9980 ( .A(n13532), .ZN(P3_U3897) );
  AND2_X1 U9981 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10537), .ZN(P2_U3947) );
  INV_X1 U9982 ( .A(n8755), .ZN(P2_U3495) );
  NAND2_X1 U9983 ( .A1(n8252), .A2(n7589), .ZN(P1_U3555) );
  NAND2_X1 U9984 ( .A1(n8257), .A2(n7590), .ZN(P1_U3523) );
  XNOR2_X1 U9985 ( .A(n9834), .B(n9833), .ZN(SUB_1596_U4) );
  NAND3_X1 U9986 ( .A1(n7617), .A2(n7616), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n7618) );
  INV_X2 U9987 ( .A(n7624), .ZN(n8806) );
  MUX2_X1 U9988 ( .A(n10402), .B(n10409), .S(n10046), .Z(n7736) );
  INV_X1 U9989 ( .A(n7736), .ZN(n7630) );
  MUX2_X1 U9990 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(P1_DATAO_REG_0__SCAN_IN), 
        .S(n7624), .Z(n7623) );
  NAND2_X1 U9991 ( .A1(n7623), .A2(SI_0_), .ZN(n7721) );
  INV_X1 U9992 ( .A(n7721), .ZN(n7629) );
  INV_X1 U9993 ( .A(n7722), .ZN(n7628) );
  INV_X1 U9994 ( .A(n7625), .ZN(n7626) );
  INV_X1 U9995 ( .A(SI_1_), .ZN(n10378) );
  NOR2_X1 U9996 ( .A1(n7626), .A2(n10378), .ZN(n7627) );
  XNOR2_X1 U9997 ( .A(n7631), .B(SI_2_), .ZN(n7737) );
  NAND2_X1 U9998 ( .A1(n7630), .A2(n7737), .ZN(n7634) );
  INV_X1 U9999 ( .A(n7631), .ZN(n7632) );
  NAND2_X1 U10000 ( .A1(n7632), .A2(SI_2_), .ZN(n7633) );
  MUX2_X1 U10001 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n6676), .Z(n7636) );
  XNOR2_X1 U10002 ( .A(n7636), .B(SI_3_), .ZN(n7751) );
  INV_X1 U10003 ( .A(n7751), .ZN(n7635) );
  NAND2_X1 U10004 ( .A1(n7752), .A2(n7635), .ZN(n7638) );
  NAND2_X1 U10005 ( .A1(n7636), .A2(SI_3_), .ZN(n7637) );
  NAND2_X1 U10006 ( .A1(n7640), .A2(SI_4_), .ZN(n7641) );
  MUX2_X1 U10007 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n10046), .Z(n7643) );
  MUX2_X1 U10008 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n10046), .Z(n7645) );
  XNOR2_X1 U10009 ( .A(n7645), .B(SI_6_), .ZN(n7787) );
  INV_X1 U10010 ( .A(n7787), .ZN(n7644) );
  NAND2_X1 U10011 ( .A1(n7788), .A2(n7644), .ZN(n7647) );
  NAND2_X1 U10012 ( .A1(n7645), .A2(SI_6_), .ZN(n7646) );
  MUX2_X1 U10013 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n6676), .Z(n7649) );
  XNOR2_X1 U10014 ( .A(n7649), .B(SI_7_), .ZN(n7802) );
  INV_X1 U10015 ( .A(n7802), .ZN(n7648) );
  NAND2_X1 U10016 ( .A1(n7649), .A2(SI_7_), .ZN(n7650) );
  MUX2_X1 U10017 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n10046), .Z(n7652) );
  XNOR2_X1 U10018 ( .A(n7652), .B(SI_8_), .ZN(n7816) );
  INV_X1 U10019 ( .A(n7816), .ZN(n7651) );
  NAND2_X1 U10020 ( .A1(n7652), .A2(SI_8_), .ZN(n7653) );
  MUX2_X1 U10021 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n10046), .Z(n7655) );
  MUX2_X1 U10022 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n6676), .Z(n7843) );
  INV_X1 U10023 ( .A(n7843), .ZN(n7656) );
  NAND2_X1 U10024 ( .A1(n7656), .A2(n10415), .ZN(n7657) );
  NAND2_X1 U10025 ( .A1(n7845), .A2(n7657), .ZN(n7659) );
  NAND2_X1 U10026 ( .A1(n7843), .A2(SI_10_), .ZN(n7658) );
  MUX2_X1 U10027 ( .A(n10684), .B(n10682), .S(n10046), .Z(n7660) );
  INV_X1 U10028 ( .A(n7660), .ZN(n7661) );
  NAND2_X1 U10029 ( .A1(n7661), .A2(SI_11_), .ZN(n7662) );
  NAND2_X1 U10030 ( .A1(n7663), .A2(n7662), .ZN(n7859) );
  MUX2_X1 U10031 ( .A(n9005), .B(n10764), .S(n10046), .Z(n7664) );
  INV_X1 U10032 ( .A(n7664), .ZN(n7665) );
  NAND2_X1 U10033 ( .A1(n7665), .A2(SI_12_), .ZN(n7666) );
  MUX2_X1 U10034 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n10046), .Z(n7888) );
  NAND2_X1 U10035 ( .A1(n7888), .A2(SI_13_), .ZN(n7668) );
  INV_X1 U10036 ( .A(n7888), .ZN(n7669) );
  NAND2_X1 U10037 ( .A1(n7669), .A2(n10449), .ZN(n7670) );
  MUX2_X1 U10038 ( .A(n11048), .B(n11046), .S(n10046), .Z(n7919) );
  MUX2_X1 U10039 ( .A(n11081), .B(n11079), .S(n10046), .Z(n7924) );
  INV_X1 U10040 ( .A(n7924), .ZN(n7671) );
  NAND2_X1 U10041 ( .A1(n7671), .A2(SI_15_), .ZN(n7675) );
  OAI21_X1 U10042 ( .B1(n7919), .B2(n10457), .A(n7675), .ZN(n7672) );
  INV_X1 U10043 ( .A(n7672), .ZN(n7673) );
  INV_X1 U10044 ( .A(n7919), .ZN(n7674) );
  NOR2_X1 U10045 ( .A1(n7674), .A2(SI_14_), .ZN(n7676) );
  AOI22_X1 U10046 ( .A1(n7676), .A2(n7675), .B1(n10497), .B2(n7924), .ZN(n7677) );
  MUX2_X1 U10047 ( .A(n11025), .B(n11023), .S(n10046), .Z(n7941) );
  XNOR2_X1 U10048 ( .A(n7940), .B(n7939), .ZN(n11021) );
  NAND4_X1 U10049 ( .A1(n8217), .A2(n8231), .A3(n8222), .A4(n8219), .ZN(n7679)
         );
  INV_X1 U10050 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n7682) );
  NOR2_X1 U10051 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n7687) );
  NOR2_X2 U10052 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n7738) );
  NAND2_X1 U10053 ( .A1(n11021), .A2(n12766), .ZN(n7697) );
  INV_X1 U10054 ( .A(n8150), .ZN(n7946) );
  NAND2_X1 U10055 ( .A1(n7946), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7695) );
  XNOR2_X1 U10056 ( .A(n7695), .B(P1_IR_REG_16__SCAN_IN), .ZN(n14716) );
  AOI22_X1 U10057 ( .A1(n12751), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7986), 
        .B2(n14716), .ZN(n7696) );
  NAND2_X1 U10058 ( .A1(n7701), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7703) );
  NAND2_X1 U10059 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n7781) );
  NAND2_X1 U10060 ( .A1(n7796), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7809) );
  INV_X1 U10061 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7808) );
  NAND2_X1 U10062 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .ZN(n7704) );
  INV_X1 U10063 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7911) );
  INV_X1 U10064 ( .A(n7933), .ZN(n7705) );
  AOI21_X1 U10065 ( .B1(n7705), .B2(P1_REG3_REG_15__SCAN_IN), .A(
        P1_REG3_REG_16__SCAN_IN), .ZN(n7707) );
  NAND2_X1 U10066 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_REG3_REG_16__SCAN_IN), 
        .ZN(n7706) );
  OR2_X1 U10067 ( .A1(n7707), .A2(n7950), .ZN(n15203) );
  INV_X1 U10068 ( .A(n15203), .ZN(n12466) );
  NAND2_X1 U10069 ( .A1(n7992), .A2(n12466), .ZN(n7715) );
  INV_X1 U10070 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7709) );
  OR2_X1 U10071 ( .A1(n10210), .A2(n7709), .ZN(n7714) );
  INV_X1 U10072 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n14720) );
  OR2_X1 U10073 ( .A1(n8115), .A2(n14720), .ZN(n7713) );
  INV_X1 U10074 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n7711) );
  OR2_X1 U10075 ( .A1(n12758), .A2(n7711), .ZN(n7712) );
  INV_X1 U10076 ( .A(n14579), .ZN(n14649) );
  INV_X1 U10077 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n14665) );
  OR2_X1 U10078 ( .A1(n7744), .A2(n14665), .ZN(n7719) );
  INV_X1 U10079 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n14673) );
  OR2_X1 U10080 ( .A1(n7784), .A2(n14673), .ZN(n7718) );
  INV_X1 U10081 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10353) );
  NAND2_X1 U10082 ( .A1(n7779), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n7716) );
  INV_X1 U10083 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n7720) );
  XNOR2_X1 U10084 ( .A(n7722), .B(n7721), .ZN(n10385) );
  INV_X1 U10085 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10467) );
  OR2_X1 U10086 ( .A1(n7744), .A2(n10467), .ZN(n7727) );
  INV_X1 U10087 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10504) );
  INV_X1 U10088 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10462) );
  NAND2_X1 U10089 ( .A1(n7779), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n7724) );
  NAND4_X2 U10090 ( .A1(n7727), .A2(n7726), .A3(n7725), .A4(n7724), .ZN(n14664) );
  NOR2_X1 U10091 ( .A1(n6676), .A2(n9810), .ZN(n7728) );
  INV_X1 U10092 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8807) );
  XNOR2_X1 U10093 ( .A(n7728), .B(n8807), .ZN(n15098) );
  NAND2_X1 U10094 ( .A1(n14664), .A2(n12578), .ZN(n11564) );
  OR2_X1 U10095 ( .A1(n14663), .A2(n10590), .ZN(n7729) );
  NAND2_X1 U10096 ( .A1(n7779), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n7735) );
  INV_X1 U10097 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n14679) );
  OR2_X1 U10098 ( .A1(n7744), .A2(n14679), .ZN(n7734) );
  INV_X1 U10099 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7730) );
  OR2_X1 U10100 ( .A1(n7784), .A2(n7730), .ZN(n7733) );
  INV_X1 U10101 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n7731) );
  NAND4_X2 U10102 ( .A1(n7735), .A2(n7734), .A3(n7733), .A4(n7732), .ZN(n14662) );
  XNOR2_X1 U10103 ( .A(n7737), .B(n7736), .ZN(n10400) );
  NAND2_X1 U10104 ( .A1(n7861), .A2(n10400), .ZN(n7741) );
  INV_X1 U10105 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n7863) );
  OR2_X1 U10106 ( .A1(n7738), .A2(n7863), .ZN(n7739) );
  NAND2_X1 U10107 ( .A1(n7986), .A2(n14681), .ZN(n7740) );
  OAI211_X1 U10108 ( .C1(n7694), .C2(n10402), .A(n7741), .B(n7740), .ZN(n12589) );
  NAND2_X1 U10109 ( .A1(n11588), .A2(n12587), .ZN(n11587) );
  OR2_X1 U10110 ( .A1(n14662), .A2(n12589), .ZN(n7743) );
  NAND2_X1 U10111 ( .A1(n12754), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7749) );
  OR2_X1 U10112 ( .A1(n7744), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n7748) );
  INV_X1 U10113 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10480) );
  OR2_X1 U10114 ( .A1(n7784), .A2(n10480), .ZN(n7747) );
  INV_X1 U10115 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7745) );
  NAND4_X1 U10116 ( .A1(n7749), .A2(n7748), .A3(n7747), .A4(n7746), .ZN(n14661) );
  OR2_X1 U10117 ( .A1(n7760), .A2(n7863), .ZN(n7750) );
  XNOR2_X1 U10118 ( .A(n7750), .B(P1_IR_REG_3__SCAN_IN), .ZN(n10475) );
  AOI22_X1 U10119 ( .A1(n7770), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n7986), .B2(
        n10475), .ZN(n7754) );
  XNOR2_X1 U10120 ( .A(n7752), .B(n7751), .ZN(n10403) );
  NAND2_X1 U10121 ( .A1(n10403), .A2(n7861), .ZN(n7753) );
  XNOR2_X2 U10122 ( .A(n14661), .B(n7755), .ZN(n10771) );
  NAND2_X1 U10123 ( .A1(n10770), .A2(n10771), .ZN(n10769) );
  NAND2_X1 U10124 ( .A1(n10769), .A2(n7756), .ZN(n10835) );
  INV_X1 U10125 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n7759) );
  NAND2_X1 U10126 ( .A1(n7760), .A2(n7759), .ZN(n7771) );
  NAND2_X1 U10127 ( .A1(n7771), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7761) );
  XNOR2_X1 U10128 ( .A(n7761), .B(P1_IR_REG_4__SCAN_IN), .ZN(n10483) );
  NAND2_X1 U10129 ( .A1(n12754), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7767) );
  INV_X1 U10130 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7762) );
  OR2_X1 U10131 ( .A1(n12758), .A2(n7762), .ZN(n7766) );
  OAI21_X1 U10132 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n7781), .ZN(n11336) );
  OR2_X1 U10133 ( .A1(n10203), .A2(n11336), .ZN(n7765) );
  INV_X1 U10134 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10482) );
  OR2_X1 U10135 ( .A1(n7784), .A2(n10482), .ZN(n7764) );
  NAND2_X1 U10136 ( .A1(n10835), .A2(n12780), .ZN(n10834) );
  NAND2_X1 U10137 ( .A1(n10834), .A2(n7768), .ZN(n10925) );
  XNOR2_X1 U10138 ( .A(n7769), .B(n7420), .ZN(n10437) );
  NAND2_X1 U10139 ( .A1(n10437), .A2(n12766), .ZN(n7778) );
  NAND2_X1 U10140 ( .A1(n7773), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7772) );
  MUX2_X1 U10141 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7772), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n7776) );
  INV_X1 U10142 ( .A(n7773), .ZN(n7775) );
  INV_X1 U10143 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n7774) );
  NAND2_X1 U10144 ( .A1(n7775), .A2(n7774), .ZN(n7790) );
  NAND2_X1 U10145 ( .A1(n7776), .A2(n7790), .ZN(n10484) );
  INV_X1 U10146 ( .A(n10484), .ZN(n10561) );
  AOI22_X1 U10147 ( .A1(n12751), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n7986), 
        .B2(n10561), .ZN(n7777) );
  NAND2_X1 U10148 ( .A1(n7778), .A2(n7777), .ZN(n12608) );
  INV_X1 U10149 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10476) );
  AND2_X1 U10150 ( .A1(n7781), .A2(n7780), .ZN(n7782) );
  OR2_X1 U10151 ( .A1(n7782), .A2(n7796), .ZN(n11213) );
  INV_X1 U10152 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7783) );
  OR2_X1 U10153 ( .A1(n7784), .A2(n7783), .ZN(n7785) );
  XNOR2_X1 U10154 ( .A(n7788), .B(n7787), .ZN(n10443) );
  NAND2_X1 U10155 ( .A1(n10443), .A2(n12766), .ZN(n7794) );
  NAND2_X1 U10156 ( .A1(n7790), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7789) );
  MUX2_X1 U10157 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7789), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n7792) );
  INV_X1 U10158 ( .A(n7790), .ZN(n7791) );
  NAND2_X1 U10159 ( .A1(n7791), .A2(n9605), .ZN(n7804) );
  AND2_X1 U10160 ( .A1(n7792), .A2(n7804), .ZN(n10523) );
  AOI22_X1 U10161 ( .A1(n12751), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n7986), 
        .B2(n10523), .ZN(n7793) );
  NAND2_X1 U10162 ( .A1(n7794), .A2(n7793), .ZN(n12611) );
  NAND2_X1 U10163 ( .A1(n12754), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7801) );
  INV_X1 U10164 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7795) );
  OR2_X1 U10165 ( .A1(n12758), .A2(n7795), .ZN(n7800) );
  OR2_X1 U10166 ( .A1(n7796), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7797) );
  NAND2_X1 U10167 ( .A1(n7809), .A2(n7797), .ZN(n11351) );
  OR2_X1 U10168 ( .A1(n10203), .A2(n11351), .ZN(n7799) );
  INV_X1 U10169 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10485) );
  OR2_X1 U10170 ( .A1(n8115), .A2(n10485), .ZN(n7798) );
  NAND4_X1 U10171 ( .A1(n7801), .A2(n7800), .A3(n7799), .A4(n7798), .ZN(n14658) );
  XNOR2_X1 U10172 ( .A(n12611), .B(n14658), .ZN(n12783) );
  INV_X1 U10173 ( .A(n12783), .ZN(n11552) );
  XNOR2_X1 U10174 ( .A(n7803), .B(n7802), .ZN(n10452) );
  NAND2_X1 U10175 ( .A1(n10452), .A2(n12766), .ZN(n7806) );
  NAND2_X1 U10176 ( .A1(n7804), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7818) );
  XNOR2_X1 U10177 ( .A(n7818), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10642) );
  AOI22_X1 U10178 ( .A1(n12751), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7986), 
        .B2(n10642), .ZN(n7805) );
  NAND2_X1 U10179 ( .A1(n7806), .A2(n7805), .ZN(n12620) );
  NAND2_X1 U10180 ( .A1(n12754), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7814) );
  INV_X1 U10181 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7807) );
  OR2_X1 U10182 ( .A1(n12758), .A2(n7807), .ZN(n7813) );
  NAND2_X1 U10183 ( .A1(n7809), .A2(n7808), .ZN(n7810) );
  NAND2_X1 U10184 ( .A1(n7836), .A2(n7810), .ZN(n11643) );
  OR2_X1 U10185 ( .A1(n10203), .A2(n11643), .ZN(n7812) );
  INV_X1 U10186 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n11487) );
  OR2_X1 U10187 ( .A1(n8115), .A2(n11487), .ZN(n7811) );
  NAND4_X1 U10188 ( .A1(n7814), .A2(n7813), .A3(n7812), .A4(n7811), .ZN(n14657) );
  XNOR2_X1 U10189 ( .A(n12620), .B(n14657), .ZN(n12784) );
  INV_X1 U10190 ( .A(n12784), .ZN(n11481) );
  NAND2_X1 U10191 ( .A1(n11479), .A2(n11481), .ZN(n11480) );
  OR2_X1 U10192 ( .A1(n12620), .A2(n14657), .ZN(n7815) );
  XNOR2_X1 U10193 ( .A(n7817), .B(n7816), .ZN(n10458) );
  NAND2_X1 U10194 ( .A1(n10458), .A2(n12766), .ZN(n7821) );
  INV_X1 U10195 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n9763) );
  NAND2_X1 U10196 ( .A1(n7818), .A2(n9763), .ZN(n7819) );
  NAND2_X1 U10197 ( .A1(n7819), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7828) );
  XNOR2_X1 U10198 ( .A(n7828), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10727) );
  AOI22_X1 U10199 ( .A1(n12751), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7986), 
        .B2(n10727), .ZN(n7820) );
  NAND2_X2 U10200 ( .A1(n7821), .A2(n7820), .ZN(n12623) );
  NAND2_X1 U10201 ( .A1(n10200), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n7825) );
  INV_X1 U10202 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10643) );
  OR2_X1 U10203 ( .A1(n10210), .A2(n10643), .ZN(n7824) );
  INV_X1 U10204 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7835) );
  XNOR2_X1 U10205 ( .A(n7836), .B(n7835), .ZN(n11932) );
  OR2_X1 U10206 ( .A1(n10203), .A2(n11932), .ZN(n7823) );
  INV_X1 U10207 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n11609) );
  OR2_X1 U10208 ( .A1(n8115), .A2(n11609), .ZN(n7822) );
  NAND4_X1 U10209 ( .A1(n7825), .A2(n7824), .A3(n7823), .A4(n7822), .ZN(n14656) );
  XNOR2_X1 U10210 ( .A(n12623), .B(n14656), .ZN(n12785) );
  XNOR2_X1 U10211 ( .A(n7827), .B(n7826), .ZN(n10515) );
  NAND2_X1 U10212 ( .A1(n10515), .A2(n7861), .ZN(n7833) );
  INV_X1 U10213 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9744) );
  NAND2_X1 U10214 ( .A1(n7828), .A2(n9744), .ZN(n7829) );
  NAND2_X1 U10215 ( .A1(n7829), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7830) );
  INV_X1 U10216 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9732) );
  NAND2_X1 U10217 ( .A1(n7830), .A2(n9732), .ZN(n7846) );
  OR2_X1 U10218 ( .A1(n7830), .A2(n9732), .ZN(n7831) );
  AOI22_X1 U10219 ( .A1(n12751), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7986), 
        .B2(n10909), .ZN(n7832) );
  NAND2_X1 U10220 ( .A1(n10200), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n7841) );
  INV_X1 U10221 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10725) );
  OR2_X1 U10222 ( .A1(n10210), .A2(n10725), .ZN(n7840) );
  INV_X1 U10223 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7834) );
  OAI21_X1 U10224 ( .B1(n7836), .B2(n7835), .A(n7834), .ZN(n7837) );
  NAND2_X1 U10225 ( .A1(n7837), .A2(n7851), .ZN(n12099) );
  OR2_X1 U10226 ( .A1(n10203), .A2(n12099), .ZN(n7839) );
  INV_X1 U10227 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n11439) );
  OR2_X1 U10228 ( .A1(n8115), .A2(n11439), .ZN(n7838) );
  NAND4_X1 U10229 ( .A1(n7841), .A2(n7840), .A3(n7839), .A4(n7838), .ZN(n14655) );
  INV_X1 U10230 ( .A(n14655), .ZN(n12092) );
  XNOR2_X1 U10231 ( .A(n12632), .B(n12092), .ZN(n12788) );
  XNOR2_X1 U10232 ( .A(n7843), .B(SI_10_), .ZN(n7844) );
  XNOR2_X1 U10233 ( .A(n7845), .B(n7844), .ZN(n10581) );
  NAND2_X1 U10234 ( .A1(n10581), .A2(n7861), .ZN(n7849) );
  NAND2_X1 U10235 ( .A1(n7846), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7847) );
  XNOR2_X1 U10236 ( .A(n7847), .B(P1_IR_REG_10__SCAN_IN), .ZN(n11054) );
  AOI22_X1 U10237 ( .A1(n12751), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n11054), 
        .B2(n7986), .ZN(n7848) );
  NAND2_X1 U10238 ( .A1(n12754), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7857) );
  INV_X1 U10239 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7850) );
  OR2_X1 U10240 ( .A1(n12758), .A2(n7850), .ZN(n7856) );
  INV_X1 U10241 ( .A(n7867), .ZN(n7853) );
  NAND2_X1 U10242 ( .A1(n7851), .A2(n10918), .ZN(n7852) );
  NAND2_X1 U10243 ( .A1(n7853), .A2(n7852), .ZN(n15190) );
  OR2_X1 U10244 ( .A1(n10203), .A2(n15190), .ZN(n7855) );
  INV_X1 U10245 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10913) );
  OR2_X1 U10246 ( .A1(n8115), .A2(n10913), .ZN(n7854) );
  NAND4_X1 U10247 ( .A1(n7857), .A2(n7856), .A3(n7855), .A4(n7854), .ZN(n14654) );
  INV_X1 U10248 ( .A(n14654), .ZN(n15207) );
  XNOR2_X1 U10249 ( .A(n12641), .B(n15207), .ZN(n12789) );
  XNOR2_X1 U10250 ( .A(n7860), .B(n7859), .ZN(n10681) );
  NAND2_X1 U10251 ( .A1(n10681), .A2(n12766), .ZN(n7866) );
  OR2_X1 U10252 ( .A1(n7862), .A2(n7863), .ZN(n7864) );
  XNOR2_X1 U10253 ( .A(n7864), .B(P1_IR_REG_11__SCAN_IN), .ZN(n11420) );
  AOI22_X1 U10254 ( .A1(n12751), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7986), 
        .B2(n11420), .ZN(n7865) );
  NAND2_X1 U10255 ( .A1(n10200), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7873) );
  NOR2_X1 U10256 ( .A1(n7867), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7868) );
  OR2_X1 U10257 ( .A1(n7881), .A2(n7868), .ZN(n15221) );
  OR2_X1 U10258 ( .A1(n10203), .A2(n15221), .ZN(n7872) );
  INV_X1 U10259 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7869) );
  OR2_X1 U10260 ( .A1(n8115), .A2(n7869), .ZN(n7871) );
  INV_X1 U10261 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n11052) );
  OR2_X1 U10262 ( .A1(n10210), .A2(n11052), .ZN(n7870) );
  NAND4_X1 U10263 ( .A1(n7873), .A2(n7872), .A3(n7871), .A4(n7870), .ZN(n14653) );
  INV_X1 U10264 ( .A(n14653), .ZN(n8171) );
  XNOR2_X1 U10265 ( .A(n15217), .B(n8171), .ZN(n12790) );
  NAND2_X1 U10266 ( .A1(n11803), .A2(n12790), .ZN(n11802) );
  NAND2_X1 U10267 ( .A1(n11802), .A2(n7874), .ZN(n12139) );
  XNOR2_X1 U10268 ( .A(n7875), .B(n7604), .ZN(n10736) );
  NAND2_X1 U10269 ( .A1(n10736), .A2(n12766), .ZN(n7880) );
  NAND2_X1 U10270 ( .A1(n7862), .A2(n9733), .ZN(n7877) );
  NAND2_X1 U10271 ( .A1(n7877), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7876) );
  MUX2_X1 U10272 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7876), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n7878) );
  AOI22_X1 U10273 ( .A1(n12751), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n7986), 
        .B2(n11712), .ZN(n7879) );
  NAND2_X1 U10274 ( .A1(n10200), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7886) );
  INV_X1 U10275 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n11713) );
  OR2_X1 U10276 ( .A1(n10210), .A2(n11713), .ZN(n7885) );
  NOR2_X1 U10277 ( .A1(n7881), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7882) );
  OR2_X1 U10278 ( .A1(n7899), .A2(n7882), .ZN(n12454) );
  OR2_X1 U10279 ( .A1(n7744), .A2(n12454), .ZN(n7884) );
  INV_X1 U10280 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n12144) );
  OR2_X1 U10281 ( .A1(n8115), .A2(n12144), .ZN(n7883) );
  NAND4_X1 U10282 ( .A1(n7886), .A2(n7885), .A3(n7884), .A4(n7883), .ZN(n14652) );
  XNOR2_X1 U10283 ( .A(n12653), .B(n14652), .ZN(n12791) );
  INV_X1 U10284 ( .A(n12791), .ZN(n12138) );
  NAND2_X1 U10285 ( .A1(n12139), .A2(n12138), .ZN(n12137) );
  NAND2_X1 U10286 ( .A1(n12137), .A2(n7887), .ZN(n12177) );
  XNOR2_X1 U10287 ( .A(n7888), .B(n10449), .ZN(n7889) );
  XNOR2_X1 U10288 ( .A(n7890), .B(n7889), .ZN(n10814) );
  NAND2_X1 U10289 ( .A1(n10814), .A2(n12766), .ZN(n7897) );
  NAND2_X1 U10290 ( .A1(n7892), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7891) );
  MUX2_X1 U10291 ( .A(n7891), .B(P1_IR_REG_31__SCAN_IN), .S(n7893), .Z(n7895)
         );
  INV_X1 U10292 ( .A(n7892), .ZN(n7894) );
  NAND2_X1 U10293 ( .A1(n7894), .A2(n7893), .ZN(n7906) );
  NAND2_X1 U10294 ( .A1(n7895), .A2(n7906), .ZN(n11756) );
  INV_X1 U10295 ( .A(n11756), .ZN(n11721) );
  AOI22_X1 U10296 ( .A1(n12751), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n7986), 
        .B2(n11721), .ZN(n7896) );
  NAND2_X1 U10297 ( .A1(n12754), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7904) );
  INV_X1 U10298 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n7898) );
  OR2_X1 U10299 ( .A1(n12758), .A2(n7898), .ZN(n7903) );
  OR2_X1 U10300 ( .A1(n7899), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7900) );
  NAND2_X1 U10301 ( .A1(n7912), .A2(n7900), .ZN(n12168) );
  OR2_X1 U10302 ( .A1(n7744), .A2(n12168), .ZN(n7902) );
  INV_X1 U10303 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11722) );
  OR2_X1 U10304 ( .A1(n8115), .A2(n11722), .ZN(n7901) );
  NAND4_X1 U10305 ( .A1(n7904), .A2(n7903), .A3(n7902), .A4(n7901), .ZN(n14651) );
  XNOR2_X1 U10306 ( .A(n12662), .B(n14651), .ZN(n12792) );
  INV_X1 U10307 ( .A(n12792), .ZN(n12178) );
  INV_X1 U10308 ( .A(n14651), .ZN(n15168) );
  NOR2_X1 U10309 ( .A1(n12662), .A2(n14651), .ZN(n7905) );
  XNOR2_X1 U10310 ( .A(n7921), .B(SI_14_), .ZN(n7920) );
  XNOR2_X1 U10311 ( .A(n7920), .B(n7919), .ZN(n11045) );
  NAND2_X1 U10312 ( .A1(n11045), .A2(n12766), .ZN(n7910) );
  NAND2_X1 U10313 ( .A1(n7906), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7907) );
  MUX2_X1 U10314 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7907), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n7908) );
  AND2_X1 U10315 ( .A1(n7908), .A2(n7927), .ZN(n14695) );
  AOI22_X1 U10316 ( .A1(n12751), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n7986), 
        .B2(n14695), .ZN(n7909) );
  NAND2_X1 U10317 ( .A1(n10200), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n7918) );
  NAND2_X1 U10318 ( .A1(n7912), .A2(n7911), .ZN(n7913) );
  NAND2_X1 U10319 ( .A1(n7933), .A2(n7913), .ZN(n15178) );
  OR2_X1 U10320 ( .A1(n7744), .A2(n15178), .ZN(n7917) );
  INV_X1 U10321 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11763) );
  OR2_X1 U10322 ( .A1(n8115), .A2(n11763), .ZN(n7916) );
  INV_X1 U10323 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7914) );
  OR2_X1 U10324 ( .A1(n10210), .A2(n7914), .ZN(n7915) );
  NAND2_X1 U10325 ( .A1(n15225), .A2(n12999), .ZN(n12666) );
  INV_X1 U10326 ( .A(n15225), .ZN(n12234) );
  NAND2_X1 U10327 ( .A1(n7920), .A2(n7919), .ZN(n7923) );
  NAND2_X1 U10328 ( .A1(n7921), .A2(n10457), .ZN(n7922) );
  NAND2_X1 U10329 ( .A1(n7923), .A2(n7922), .ZN(n7926) );
  XNOR2_X1 U10330 ( .A(n7924), .B(SI_15_), .ZN(n7925) );
  NAND2_X1 U10331 ( .A1(n11078), .A2(n12766), .ZN(n7931) );
  NAND2_X1 U10332 ( .A1(n7927), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7928) );
  MUX2_X1 U10333 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7928), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n7929) );
  AND2_X1 U10334 ( .A1(n7929), .A2(n7946), .ZN(n15262) );
  AOI22_X1 U10335 ( .A1(n12751), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n7986), 
        .B2(n15262), .ZN(n7930) );
  NAND2_X1 U10336 ( .A1(n10200), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n7938) );
  INV_X1 U10337 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n15258) );
  OR2_X1 U10338 ( .A1(n10210), .A2(n15258), .ZN(n7937) );
  INV_X1 U10339 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7932) );
  XNOR2_X1 U10340 ( .A(n7933), .B(n7932), .ZN(n12417) );
  OR2_X1 U10341 ( .A1(n7744), .A2(n12417), .ZN(n7936) );
  INV_X1 U10342 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7934) );
  OR2_X1 U10343 ( .A1(n8115), .A2(n7934), .ZN(n7935) );
  NAND2_X1 U10344 ( .A1(n13009), .A2(n15192), .ZN(n12675) );
  NAND2_X1 U10345 ( .A1(n12670), .A2(n12675), .ZN(n12797) );
  INV_X1 U10346 ( .A(n15192), .ZN(n14650) );
  XNOR2_X1 U10347 ( .A(n15200), .B(n14579), .ZN(n12798) );
  NAND2_X1 U10348 ( .A1(n7941), .A2(n10572), .ZN(n7942) );
  MUX2_X1 U10349 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(P1_DATAO_REG_17__SCAN_IN), 
        .S(n10046), .Z(n7957) );
  INV_X1 U10350 ( .A(n7957), .ZN(n7944) );
  XNOR2_X1 U10351 ( .A(n7944), .B(SI_17_), .ZN(n7945) );
  XNOR2_X1 U10352 ( .A(n7959), .B(n7945), .ZN(n11063) );
  NAND2_X1 U10353 ( .A1(n11063), .A2(n12766), .ZN(n7949) );
  OAI21_X1 U10354 ( .B1(n7946), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7947) );
  XNOR2_X1 U10355 ( .A(n7947), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14733) );
  AOI22_X1 U10356 ( .A1(n12751), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n7986), 
        .B2(n14733), .ZN(n7948) );
  NOR2_X1 U10357 ( .A1(n7950), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n7951) );
  OR2_X1 U10358 ( .A1(n7966), .A2(n7951), .ZN(n12555) );
  INV_X1 U10359 ( .A(n12555), .ZN(n14581) );
  NAND2_X1 U10360 ( .A1(n14581), .A2(n7992), .ZN(n7956) );
  NAND2_X1 U10361 ( .A1(n12754), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n7955) );
  INV_X1 U10362 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n7952) );
  OR2_X1 U10363 ( .A1(n12758), .A2(n7952), .ZN(n7954) );
  INV_X1 U10364 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14722) );
  OR2_X1 U10365 ( .A1(n8115), .A2(n14722), .ZN(n7953) );
  NAND4_X1 U10366 ( .A1(n7956), .A2(n7955), .A3(n7954), .A4(n7953), .ZN(n14973) );
  NAND2_X1 U10367 ( .A1(n14573), .A2(n14973), .ZN(n12683) );
  NOR2_X1 U10368 ( .A1(n14573), .A2(n14973), .ZN(n12673) );
  AOI21_X1 U10369 ( .B1(n12554), .B2(n12683), .A(n12673), .ZN(n14970) );
  NAND2_X1 U10370 ( .A1(n7957), .A2(SI_17_), .ZN(n7958) );
  MUX2_X1 U10371 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n10046), .Z(n8001) );
  NAND2_X1 U10372 ( .A1(n6809), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7961) );
  MUX2_X1 U10373 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7961), .S(
        P1_IR_REG_18__SCAN_IN), .Z(n7963) );
  AND2_X1 U10374 ( .A1(n7963), .A2(n7982), .ZN(n14751) );
  AOI22_X1 U10375 ( .A1(n12751), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n7986), 
        .B2(n14751), .ZN(n7964) );
  OR2_X1 U10376 ( .A1(n7966), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n7967) );
  NAND2_X1 U10377 ( .A1(n7990), .A2(n7967), .ZN(n14983) );
  NAND2_X1 U10378 ( .A1(n7763), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7968) );
  OAI21_X1 U10379 ( .B1(n14983), .B2(n10203), .A(n7968), .ZN(n7972) );
  INV_X1 U10380 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n7970) );
  NAND2_X1 U10381 ( .A1(n12754), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n7969) );
  OAI21_X1 U10382 ( .B1(n12758), .B2(n7970), .A(n7969), .ZN(n7971) );
  NAND2_X1 U10383 ( .A1(n14991), .A2(n14648), .ZN(n12685) );
  INV_X1 U10384 ( .A(n12685), .ZN(n7973) );
  INV_X1 U10385 ( .A(n7974), .ZN(n7975) );
  NAND2_X1 U10386 ( .A1(n7975), .A2(n8001), .ZN(n7977) );
  NAND2_X1 U10387 ( .A1(n8000), .A2(SI_18_), .ZN(n7976) );
  NAND2_X1 U10388 ( .A1(n7977), .A2(n7976), .ZN(n7981) );
  MUX2_X1 U10389 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n6676), .Z(n7978) );
  NAND2_X1 U10390 ( .A1(n7978), .A2(SI_19_), .ZN(n8004) );
  INV_X1 U10391 ( .A(n7978), .ZN(n7979) );
  INV_X1 U10392 ( .A(SI_19_), .ZN(n10784) );
  NAND2_X1 U10393 ( .A1(n7979), .A2(n10784), .ZN(n8002) );
  NAND2_X1 U10394 ( .A1(n8004), .A2(n8002), .ZN(n7980) );
  XNOR2_X2 U10395 ( .A(n7981), .B(n7980), .ZN(n11596) );
  NAND2_X1 U10396 ( .A1(n11596), .A2(n12766), .ZN(n7988) );
  AOI22_X1 U10397 ( .A1(n12751), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n15275), 
        .B2(n7986), .ZN(n7987) );
  NAND2_X2 U10398 ( .A1(n7988), .A2(n7987), .ZN(n14965) );
  INV_X1 U10399 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n7989) );
  NAND2_X1 U10400 ( .A1(n7990), .A2(n7989), .ZN(n7991) );
  AND2_X1 U10401 ( .A1(n8010), .A2(n7991), .ZN(n14961) );
  NAND2_X1 U10402 ( .A1(n14961), .A2(n7992), .ZN(n7995) );
  AOI22_X1 U10403 ( .A1(n10200), .A2(P1_REG0_REG_19__SCAN_IN), .B1(n12754), 
        .B2(P1_REG1_REG_19__SCAN_IN), .ZN(n7994) );
  NAND2_X1 U10404 ( .A1(n7763), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n7993) );
  OR2_X1 U10405 ( .A1(n14965), .A2(n14597), .ZN(n12691) );
  NAND2_X1 U10406 ( .A1(n14965), .A2(n14597), .ZN(n12692) );
  INV_X1 U10407 ( .A(n14597), .ZN(n14976) );
  INV_X1 U10408 ( .A(n8001), .ZN(n7998) );
  OAI21_X1 U10409 ( .B1(n10739), .B2(n7998), .A(n8004), .ZN(n7999) );
  NOR2_X1 U10410 ( .A1(n8001), .A2(SI_18_), .ZN(n8005) );
  INV_X1 U10411 ( .A(n8002), .ZN(n8003) );
  AOI21_X1 U10412 ( .B1(n8005), .B2(n8004), .A(n8003), .ZN(n8006) );
  XNOR2_X1 U10413 ( .A(n8034), .B(n11026), .ZN(n8016) );
  MUX2_X1 U10414 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n6676), .Z(n8029) );
  XNOR2_X1 U10415 ( .A(n8016), .B(n8029), .ZN(n11707) );
  NAND2_X1 U10416 ( .A1(n11707), .A2(n12766), .ZN(n8008) );
  NAND2_X1 U10417 ( .A1(n12751), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8007) );
  INV_X1 U10418 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8009) );
  NAND2_X1 U10419 ( .A1(n8010), .A2(n8009), .ZN(n8012) );
  INV_X1 U10420 ( .A(n8023), .ZN(n8011) );
  NAND2_X1 U10421 ( .A1(n8012), .A2(n8011), .ZN(n14945) );
  AOI22_X1 U10422 ( .A1(n10200), .A2(P1_REG0_REG_20__SCAN_IN), .B1(n12754), 
        .B2(P1_REG1_REG_20__SCAN_IN), .ZN(n8014) );
  NAND2_X1 U10423 ( .A1(n7763), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8013) );
  OAI211_X1 U10424 ( .C1(n14945), .C2(n10203), .A(n8014), .B(n8013), .ZN(
        n14647) );
  INV_X1 U10425 ( .A(n14647), .ZN(n8186) );
  XNOR2_X1 U10426 ( .A(n15048), .B(n8186), .ZN(n14934) );
  INV_X1 U10427 ( .A(n14934), .ZN(n14941) );
  INV_X1 U10428 ( .A(n8016), .ZN(n8018) );
  NOR2_X1 U10429 ( .A1(n8034), .A2(n11026), .ZN(n8017) );
  AOI21_X1 U10430 ( .B1(n8018), .B2(n8029), .A(n8017), .ZN(n8020) );
  MUX2_X1 U10431 ( .A(n11816), .B(n11814), .S(n6676), .Z(n8028) );
  XNOR2_X1 U10432 ( .A(n8028), .B(SI_21_), .ZN(n8019) );
  XNOR2_X1 U10433 ( .A(n8020), .B(n8019), .ZN(n11813) );
  NAND2_X1 U10434 ( .A1(n11813), .A2(n12766), .ZN(n8022) );
  NAND2_X1 U10435 ( .A1(n12751), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8021) );
  NAND2_X1 U10436 ( .A1(n12754), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n8027) );
  INV_X1 U10437 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n15087) );
  OR2_X1 U10438 ( .A1(n12758), .A2(n15087), .ZN(n8026) );
  NAND2_X1 U10439 ( .A1(n8023), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8036) );
  OAI21_X1 U10440 ( .B1(P1_REG3_REG_21__SCAN_IN), .B2(n8023), .A(n8036), .ZN(
        n14925) );
  OR2_X1 U10441 ( .A1(n7744), .A2(n14925), .ZN(n8025) );
  INV_X1 U10442 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n14926) );
  OR2_X1 U10443 ( .A1(n8115), .A2(n14926), .ZN(n8024) );
  NAND4_X1 U10444 ( .A1(n8027), .A2(n8026), .A3(n8025), .A4(n8024), .ZN(n14646) );
  XNOR2_X1 U10445 ( .A(n14928), .B(n14646), .ZN(n12802) );
  INV_X1 U10446 ( .A(n8029), .ZN(n8030) );
  NOR2_X1 U10447 ( .A1(n8030), .A2(n11026), .ZN(n8032) );
  AOI22_X1 U10448 ( .A1(n8032), .A2(n7613), .B1(n8031), .B2(SI_21_), .ZN(n8033) );
  OR2_X1 U10449 ( .A1(n8554), .A2(n10046), .ZN(n8035) );
  XNOR2_X1 U10450 ( .A(n8035), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15096) );
  NAND2_X1 U10451 ( .A1(n10200), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8042) );
  INV_X1 U10452 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n14911) );
  OR2_X1 U10453 ( .A1(n8115), .A2(n14911), .ZN(n8041) );
  OAI21_X1 U10454 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n8037), .A(n8054), .ZN(
        n14910) );
  OR2_X1 U10455 ( .A1(n7744), .A2(n14910), .ZN(n8040) );
  INV_X1 U10456 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n8038) );
  OR2_X1 U10457 ( .A1(n10210), .A2(n8038), .ZN(n8039) );
  NAND4_X1 U10458 ( .A1(n8042), .A2(n8041), .A3(n8040), .A4(n8039), .ZN(n14888) );
  NAND2_X1 U10459 ( .A1(n14915), .A2(n14888), .ZN(n8043) );
  NAND2_X1 U10460 ( .A1(n8192), .A2(n8043), .ZN(n14907) );
  INV_X1 U10461 ( .A(n14888), .ZN(n8044) );
  INV_X1 U10462 ( .A(n8554), .ZN(n8046) );
  MUX2_X1 U10463 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n6676), .Z(n8553) );
  NAND2_X1 U10464 ( .A1(n8046), .A2(n8553), .ZN(n8048) );
  NAND2_X1 U10465 ( .A1(n8066), .A2(SI_22_), .ZN(n8047) );
  NAND2_X1 U10466 ( .A1(n8048), .A2(n8047), .ZN(n8050) );
  MUX2_X1 U10467 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n10046), .Z(n8068) );
  XNOR2_X1 U10468 ( .A(n8068), .B(SI_23_), .ZN(n8049) );
  XNOR2_X2 U10469 ( .A(n8050), .B(n8049), .ZN(n12058) );
  NAND2_X1 U10470 ( .A1(n12058), .A2(n12766), .ZN(n8052) );
  NAND2_X1 U10471 ( .A1(n12751), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8051) );
  NAND2_X2 U10472 ( .A1(n8052), .A2(n8051), .ZN(n14898) );
  NAND2_X1 U10473 ( .A1(n12754), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n8060) );
  INV_X1 U10474 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n8053) );
  OR2_X1 U10475 ( .A1(n12758), .A2(n8053), .ZN(n8059) );
  OAI21_X1 U10476 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n8055), .A(n8076), .ZN(
        n14896) );
  OR2_X1 U10477 ( .A1(n7744), .A2(n14896), .ZN(n8058) );
  INV_X1 U10478 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n8056) );
  OR2_X1 U10479 ( .A1(n8115), .A2(n8056), .ZN(n8057) );
  NAND4_X1 U10480 ( .A1(n8060), .A2(n8059), .A3(n8058), .A4(n8057), .ZN(n14645) );
  INV_X1 U10481 ( .A(n14645), .ZN(n14870) );
  NAND2_X1 U10482 ( .A1(n14898), .A2(n14870), .ZN(n14865) );
  OR2_X1 U10483 ( .A1(n14898), .A2(n14870), .ZN(n8061) );
  NAND2_X1 U10484 ( .A1(n14865), .A2(n8061), .ZN(n12801) );
  INV_X1 U10485 ( .A(n8068), .ZN(n8063) );
  INV_X1 U10486 ( .A(SI_23_), .ZN(n11408) );
  NAND2_X1 U10487 ( .A1(n8063), .A2(n11408), .ZN(n8069) );
  OAI21_X1 U10488 ( .B1(n8553), .B2(SI_22_), .A(n8069), .ZN(n8064) );
  INV_X1 U10489 ( .A(n8064), .ZN(n8065) );
  INV_X1 U10490 ( .A(n8553), .ZN(n8067) );
  INV_X1 U10491 ( .A(SI_22_), .ZN(n9183) );
  NOR2_X1 U10492 ( .A1(n8067), .A2(n9183), .ZN(n8070) );
  AOI22_X1 U10493 ( .A1(n8070), .A2(n8069), .B1(n8068), .B2(SI_23_), .ZN(n8071) );
  MUX2_X1 U10494 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n10046), .Z(n8083) );
  XNOR2_X1 U10495 ( .A(n8085), .B(n8083), .ZN(n12120) );
  NAND2_X1 U10496 ( .A1(n12120), .A2(n12766), .ZN(n8074) );
  NAND2_X1 U10497 ( .A1(n12751), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8073) );
  NAND2_X1 U10498 ( .A1(n12754), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8081) );
  INV_X1 U10499 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n8075) );
  OR2_X1 U10500 ( .A1(n12758), .A2(n8075), .ZN(n8080) );
  OAI21_X1 U10501 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n8077), .A(n8095), .ZN(
        n14876) );
  OR2_X1 U10502 ( .A1(n7744), .A2(n14876), .ZN(n8079) );
  INV_X1 U10503 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n14877) );
  OR2_X1 U10504 ( .A1(n8115), .A2(n14877), .ZN(n8078) );
  NAND4_X1 U10505 ( .A1(n8081), .A2(n8080), .A3(n8079), .A4(n8078), .ZN(n14887) );
  XNOR2_X1 U10506 ( .A(n14883), .B(n14887), .ZN(n12803) );
  INV_X1 U10507 ( .A(n14887), .ZN(n13072) );
  NAND2_X1 U10508 ( .A1(n14880), .A2(n13072), .ZN(n8082) );
  INV_X1 U10509 ( .A(n8083), .ZN(n8084) );
  NAND2_X1 U10510 ( .A1(n8086), .A2(SI_24_), .ZN(n8087) );
  INV_X1 U10511 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n12574) );
  MUX2_X1 U10512 ( .A(n12574), .B(n12167), .S(n10046), .Z(n8089) );
  INV_X1 U10513 ( .A(SI_25_), .ZN(n12038) );
  NAND2_X1 U10514 ( .A1(n8089), .A2(n12038), .ZN(n8106) );
  INV_X1 U10515 ( .A(n8089), .ZN(n8090) );
  NAND2_X1 U10516 ( .A1(n8090), .A2(SI_25_), .ZN(n8091) );
  NAND2_X1 U10517 ( .A1(n8106), .A2(n8091), .ZN(n8104) );
  XNOR2_X1 U10518 ( .A(n8105), .B(n8104), .ZN(n12165) );
  NAND2_X1 U10519 ( .A1(n12165), .A2(n12766), .ZN(n8093) );
  NAND2_X1 U10520 ( .A1(n12751), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8092) );
  NAND2_X1 U10521 ( .A1(n12754), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8100) );
  INV_X1 U10522 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n8094) );
  OR2_X1 U10523 ( .A1(n12758), .A2(n8094), .ZN(n8099) );
  OAI21_X1 U10524 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n8096), .A(n8113), .ZN(
        n14854) );
  OR2_X1 U10525 ( .A1(n7744), .A2(n14854), .ZN(n8098) );
  INV_X1 U10526 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n14855) );
  OR2_X1 U10527 ( .A1(n8115), .A2(n14855), .ZN(n8097) );
  NAND4_X1 U10528 ( .A1(n8100), .A2(n8099), .A3(n8098), .A4(n8097), .ZN(n14644) );
  NAND2_X1 U10529 ( .A1(n15017), .A2(n14644), .ZN(n8103) );
  OR2_X1 U10530 ( .A1(n15017), .A2(n14644), .ZN(n8101) );
  NAND2_X1 U10531 ( .A1(n8103), .A2(n8101), .ZN(n14850) );
  INV_X1 U10532 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n12389) );
  INV_X1 U10533 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n12385) );
  MUX2_X1 U10534 ( .A(n12389), .B(n12385), .S(n10046), .Z(n8123) );
  XNOR2_X1 U10535 ( .A(n8123), .B(SI_26_), .ZN(n8107) );
  NAND2_X1 U10536 ( .A1(n12384), .A2(n12766), .ZN(n8109) );
  NAND2_X1 U10537 ( .A1(n12751), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8108) );
  NAND2_X1 U10538 ( .A1(n10200), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8119) );
  INV_X1 U10539 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n8110) );
  OR2_X1 U10540 ( .A1(n10210), .A2(n8110), .ZN(n8118) );
  INV_X1 U10541 ( .A(n8113), .ZN(n8111) );
  NAND2_X1 U10542 ( .A1(n8111), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8133) );
  INV_X1 U10543 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8112) );
  NAND2_X1 U10544 ( .A1(n8113), .A2(n8112), .ZN(n8114) );
  NAND2_X1 U10545 ( .A1(n8133), .A2(n8114), .ZN(n14837) );
  INV_X1 U10546 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n14840) );
  OR2_X1 U10547 ( .A1(n8115), .A2(n14840), .ZN(n8116) );
  NAND4_X1 U10548 ( .A1(n8119), .A2(n8118), .A3(n8117), .A4(n8116), .ZN(n14643) );
  NAND2_X1 U10549 ( .A1(n14622), .A2(n13091), .ZN(n8195) );
  OR2_X1 U10550 ( .A1(n14622), .A2(n13091), .ZN(n8120) );
  NAND2_X1 U10551 ( .A1(n8195), .A2(n8120), .ZN(n12806) );
  NAND2_X1 U10552 ( .A1(n14830), .A2(n12806), .ZN(n8122) );
  NAND2_X1 U10553 ( .A1(n14622), .A2(n14643), .ZN(n8121) );
  INV_X1 U10554 ( .A(SI_26_), .ZN(n12150) );
  NAND2_X1 U10555 ( .A1(n8124), .A2(n12150), .ZN(n8125) );
  INV_X1 U10556 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n12475) );
  INV_X1 U10557 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n12479) );
  MUX2_X1 U10558 ( .A(n12475), .B(n12479), .S(n10046), .Z(n8621) );
  XNOR2_X1 U10559 ( .A(n8621), .B(SI_27_), .ZN(n8127) );
  NAND2_X1 U10560 ( .A1(n12474), .A2(n12766), .ZN(n8129) );
  NAND2_X1 U10561 ( .A1(n12751), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8128) );
  NAND2_X1 U10562 ( .A1(n10200), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8139) );
  INV_X1 U10563 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n8130) );
  OR2_X1 U10564 ( .A1(n10210), .A2(n8130), .ZN(n8138) );
  INV_X1 U10565 ( .A(n8133), .ZN(n8131) );
  NAND2_X1 U10566 ( .A1(n8131), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n10201) );
  INV_X1 U10567 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8132) );
  NAND2_X1 U10568 ( .A1(n8133), .A2(n8132), .ZN(n8134) );
  NAND2_X1 U10569 ( .A1(n10201), .A2(n8134), .ZN(n14822) );
  OR2_X1 U10570 ( .A1(n7744), .A2(n14822), .ZN(n8137) );
  INV_X1 U10571 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n8135) );
  OR2_X1 U10572 ( .A1(n8115), .A2(n8135), .ZN(n8136) );
  NAND4_X1 U10573 ( .A1(n8139), .A2(n8138), .A3(n8137), .A4(n8136), .ZN(n14803) );
  NAND2_X1 U10574 ( .A1(n14537), .A2(n13101), .ZN(n10192) );
  OR2_X1 U10575 ( .A1(n14537), .A2(n13101), .ZN(n8140) );
  NAND2_X1 U10576 ( .A1(n10192), .A2(n8140), .ZN(n12807) );
  INV_X1 U10577 ( .A(n10220), .ZN(n8143) );
  INV_X1 U10578 ( .A(n8148), .ZN(n8149) );
  NAND2_X1 U10579 ( .A1(n8150), .A2(n8149), .ZN(n8218) );
  NAND2_X1 U10580 ( .A1(n8218), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8151) );
  AND2_X1 U10581 ( .A1(n14764), .A2(n15097), .ZN(n8152) );
  NAND2_X1 U10582 ( .A1(n12577), .A2(n15097), .ZN(n8153) );
  NAND2_X1 U10583 ( .A1(n13115), .A2(n8153), .ZN(n11145) );
  NAND2_X1 U10584 ( .A1(n8154), .A2(n12777), .ZN(n8156) );
  INV_X1 U10585 ( .A(n12587), .ZN(n8157) );
  INV_X1 U10586 ( .A(n12589), .ZN(n15301) );
  OR2_X1 U10587 ( .A1(n14662), .A2(n15301), .ZN(n8158) );
  NAND2_X1 U10588 ( .A1(n8159), .A2(n8158), .ZN(n10768) );
  NAND2_X1 U10589 ( .A1(n10768), .A2(n12778), .ZN(n8161) );
  OR2_X1 U10590 ( .A1(n14661), .A2(n7755), .ZN(n8160) );
  NAND2_X1 U10591 ( .A1(n8161), .A2(n8160), .ZN(n10833) );
  NAND2_X1 U10592 ( .A1(n10833), .A2(n6671), .ZN(n8163) );
  INV_X1 U10593 ( .A(n14660), .ZN(n11197) );
  NAND2_X1 U10594 ( .A1(n11197), .A2(n12599), .ZN(n8162) );
  NAND2_X1 U10595 ( .A1(n8163), .A2(n8162), .ZN(n10928) );
  INV_X1 U10596 ( .A(n12781), .ZN(n8164) );
  NAND2_X1 U10597 ( .A1(n12608), .A2(n8165), .ZN(n8166) );
  INV_X1 U10598 ( .A(n14658), .ZN(n11346) );
  OR2_X1 U10599 ( .A1(n12611), .A2(n11346), .ZN(n8167) );
  INV_X1 U10600 ( .A(n12620), .ZN(n11476) );
  OR2_X2 U10601 ( .A1(n11600), .A2(n11599), .ZN(n11602) );
  INV_X1 U10602 ( .A(n14656), .ZN(n11645) );
  OR2_X1 U10603 ( .A1(n12623), .A2(n11645), .ZN(n8168) );
  NAND2_X1 U10604 ( .A1(n11602), .A2(n8168), .ZN(n11431) );
  INV_X1 U10605 ( .A(n11431), .ZN(n8169) );
  NAND2_X1 U10606 ( .A1(n12632), .A2(n12092), .ZN(n8170) );
  INV_X1 U10607 ( .A(n12790), .ZN(n11799) );
  NAND2_X1 U10608 ( .A1(n11800), .A2(n11799), .ZN(n8173) );
  OR2_X1 U10609 ( .A1(n15217), .A2(n8171), .ZN(n8172) );
  NAND2_X1 U10610 ( .A1(n8173), .A2(n8172), .ZN(n12136) );
  NAND2_X1 U10611 ( .A1(n12136), .A2(n12791), .ZN(n8175) );
  INV_X1 U10612 ( .A(n14652), .ZN(n15204) );
  OR2_X1 U10613 ( .A1(n12653), .A2(n15204), .ZN(n8174) );
  NAND2_X1 U10614 ( .A1(n8175), .A2(n8174), .ZN(n12171) );
  NAND2_X1 U10615 ( .A1(n12171), .A2(n12792), .ZN(n8177) );
  OR2_X1 U10616 ( .A1(n12662), .A2(n15168), .ZN(n8176) );
  NAND2_X1 U10617 ( .A1(n8177), .A2(n8176), .ZN(n12237) );
  NAND2_X1 U10618 ( .A1(n12237), .A2(n12668), .ZN(n8178) );
  NAND2_X1 U10619 ( .A1(n8178), .A2(n12669), .ZN(n12412) );
  NAND2_X1 U10620 ( .A1(n12412), .A2(n12413), .ZN(n8179) );
  INV_X1 U10621 ( .A(n12798), .ZN(n8180) );
  OR2_X1 U10622 ( .A1(n13017), .A2(n14649), .ZN(n8181) );
  INV_X1 U10623 ( .A(n12673), .ZN(n8182) );
  NAND2_X1 U10624 ( .A1(n8182), .A2(n12683), .ZN(n12794) );
  INV_X1 U10625 ( .A(n14973), .ZN(n15191) );
  OR2_X1 U10626 ( .A1(n14573), .A2(n15191), .ZN(n8183) );
  INV_X1 U10627 ( .A(n14648), .ZN(n12549) );
  OR2_X1 U10628 ( .A1(n14991), .A2(n12549), .ZN(n8185) );
  NAND2_X1 U10629 ( .A1(n14933), .A2(n14941), .ZN(n14937) );
  OR2_X1 U10630 ( .A1(n15048), .A2(n8186), .ZN(n8187) );
  NAND2_X1 U10631 ( .A1(n14937), .A2(n8187), .ZN(n14921) );
  NAND2_X1 U10632 ( .A1(n14921), .A2(n12802), .ZN(n8189) );
  INV_X1 U10633 ( .A(n14646), .ZN(n14596) );
  OR2_X1 U10634 ( .A1(n14596), .A2(n14928), .ZN(n8188) );
  NAND2_X1 U10635 ( .A1(n8189), .A2(n8188), .ZN(n14905) );
  INV_X1 U10636 ( .A(n14905), .ZN(n8191) );
  INV_X1 U10637 ( .A(n14907), .ZN(n8190) );
  NAND2_X1 U10638 ( .A1(n14883), .A2(n13072), .ZN(n8193) );
  NAND2_X1 U10639 ( .A1(n14851), .A2(n14850), .ZN(n14849) );
  INV_X1 U10640 ( .A(n14644), .ZN(n14872) );
  NAND2_X1 U10641 ( .A1(n15017), .A2(n14872), .ZN(n8194) );
  NAND2_X1 U10642 ( .A1(n14849), .A2(n8194), .ZN(n14832) );
  NAND2_X1 U10643 ( .A1(n14832), .A2(n14831), .ZN(n14834) );
  NAND2_X1 U10644 ( .A1(n14834), .A2(n8195), .ZN(n8196) );
  NAND2_X1 U10645 ( .A1(n8196), .A2(n8197), .ZN(n10193) );
  OAI21_X1 U10646 ( .B1(n8197), .B2(n8196), .A(n10193), .ZN(n8208) );
  INV_X1 U10647 ( .A(n8213), .ZN(n12812) );
  NAND2_X1 U10648 ( .A1(n8198), .A2(n12812), .ZN(n12763) );
  NAND2_X1 U10649 ( .A1(n15275), .A2(n15097), .ZN(n12576) );
  NAND2_X1 U10650 ( .A1(n10200), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8205) );
  INV_X1 U10651 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n8199) );
  OR2_X1 U10652 ( .A1(n10210), .A2(n8199), .ZN(n8204) );
  INV_X1 U10653 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8200) );
  XNOR2_X1 U10654 ( .A(n10201), .B(n8200), .ZN(n14813) );
  OR2_X1 U10655 ( .A1(n7744), .A2(n14813), .ZN(n8203) );
  INV_X1 U10656 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n8201) );
  OR2_X1 U10657 ( .A1(n8115), .A2(n8201), .ZN(n8202) );
  NAND4_X1 U10658 ( .A1(n8205), .A2(n8204), .A3(n8203), .A4(n8202), .ZN(n14642) );
  NAND2_X1 U10659 ( .A1(n8198), .A2(n15097), .ZN(n12771) );
  INV_X1 U10660 ( .A(n12993), .ZN(n10465) );
  OAI22_X1 U10661 ( .A1(n13113), .A2(n14871), .B1(n13091), .B2(n14869), .ZN(
        n8207) );
  AOI21_X1 U10662 ( .B1(n8208), .B2(n6966), .A(n8207), .ZN(n8209) );
  OAI21_X1 U10663 ( .B1(n8210), .B2(n11145), .A(n8209), .ZN(n14828) );
  INV_X1 U10664 ( .A(n14828), .ZN(n8216) );
  INV_X1 U10665 ( .A(n12653), .ZN(n15117) );
  NAND2_X1 U10666 ( .A1(n11590), .A2(n15301), .ZN(n11589) );
  OR2_X1 U10667 ( .A1(n11589), .A2(n12593), .ZN(n10836) );
  INV_X1 U10668 ( .A(n12608), .ZN(n11148) );
  INV_X1 U10669 ( .A(n12611), .ZN(n11548) );
  NAND2_X1 U10670 ( .A1(n11549), .A2(n11548), .ZN(n11547) );
  OR2_X1 U10671 ( .A1(n11547), .A2(n12620), .ZN(n11605) );
  OR2_X1 U10672 ( .A1(n12179), .A2(n12662), .ZN(n12227) );
  INV_X1 U10673 ( .A(n14573), .ZN(n13022) );
  INV_X1 U10674 ( .A(n14898), .ZN(n8212) );
  INV_X1 U10675 ( .A(n15017), .ZN(n14859) );
  AND2_X2 U10676 ( .A1(n14852), .A2(n14859), .ZN(n14853) );
  OR2_X1 U10677 ( .A1(n14839), .A2(n14826), .ZN(n8214) );
  INV_X1 U10678 ( .A(n15097), .ZN(n12575) );
  NAND2_X1 U10679 ( .A1(n8213), .A2(n12575), .ZN(n12770) );
  INV_X1 U10680 ( .A(n14821), .ZN(n8215) );
  NOR2_X2 U10681 ( .A1(n8218), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n8229) );
  NAND2_X1 U10682 ( .A1(n8229), .A2(n8231), .ZN(n8221) );
  NAND2_X1 U10683 ( .A1(n8150), .A2(n8224), .ZN(n8225) );
  NAND2_X1 U10684 ( .A1(n8225), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8226) );
  MUX2_X1 U10685 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8226), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n8228) );
  NAND2_X1 U10686 ( .A1(n8228), .A2(n8227), .ZN(n12387) );
  INV_X1 U10687 ( .A(n8229), .ZN(n8230) );
  NAND2_X1 U10688 ( .A1(n8230), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8232) );
  XNOR2_X1 U10689 ( .A(n8232), .B(n8231), .ZN(n10354) );
  OAI211_X1 U10690 ( .C1(n12771), .C2(n8251), .A(n10503), .B(n10354), .ZN(
        n10825) );
  INV_X1 U10691 ( .A(n12843), .ZN(n11140) );
  OR2_X1 U10692 ( .A1(n12123), .A2(P1_B_REG_SCAN_IN), .ZN(n8234) );
  INV_X1 U10693 ( .A(n12387), .ZN(n8233) );
  AND2_X1 U10694 ( .A1(n8234), .A2(n8233), .ZN(n8236) );
  NAND3_X1 U10695 ( .A1(n12572), .A2(P1_B_REG_SCAN_IN), .A3(n12123), .ZN(n8235) );
  NAND2_X1 U10696 ( .A1(n12572), .A2(n12387), .ZN(n10501) );
  OAI21_X1 U10697 ( .B1(n10500), .B2(P1_D_REG_1__SCAN_IN), .A(n10501), .ZN(
        n8248) );
  INV_X1 U10698 ( .A(n8198), .ZN(n12813) );
  NAND2_X1 U10699 ( .A1(n10222), .A2(n12813), .ZN(n11141) );
  NOR4_X1 U10700 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n8240) );
  NOR4_X1 U10701 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n8239) );
  NOR4_X1 U10702 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n8238) );
  NOR4_X1 U10703 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n8237) );
  NAND4_X1 U10704 ( .A1(n8240), .A2(n8239), .A3(n8238), .A4(n8237), .ZN(n8246)
         );
  NOR2_X1 U10705 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n8244) );
  NOR4_X1 U10706 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n8243) );
  NOR4_X1 U10707 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n8242) );
  NOR4_X1 U10708 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n8241) );
  NAND4_X1 U10709 ( .A1(n8244), .A2(n8243), .A3(n8242), .A4(n8241), .ZN(n8245)
         );
  NOR2_X1 U10710 ( .A1(n8246), .A2(n8245), .ZN(n10498) );
  OR2_X1 U10711 ( .A1(n10500), .A2(n10498), .ZN(n8247) );
  AND3_X1 U10712 ( .A1(n8248), .A2(n11141), .A3(n8247), .ZN(n8253) );
  NAND2_X1 U10713 ( .A1(n12123), .A2(n12387), .ZN(n10430) );
  MUX2_X1 U10714 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n8255), .S(n15332), .Z(
        n8250) );
  INV_X1 U10715 ( .A(n8250), .ZN(n8252) );
  OR2_X1 U10716 ( .A1(n8198), .A2(n15097), .ZN(n15273) );
  NOR2_X2 U10717 ( .A1(n15273), .A2(n8251), .ZN(n15224) );
  NAND2_X1 U10718 ( .A1(n15332), .A2(n15224), .ZN(n15046) );
  NOR2_X1 U10719 ( .A1(n12843), .A2(n11137), .ZN(n8254) );
  MUX2_X1 U10720 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n8255), .S(n15324), .Z(
        n8256) );
  INV_X1 U10721 ( .A(n8256), .ZN(n8257) );
  NAND2_X1 U10722 ( .A1(n15324), .A2(n15224), .ZN(n15089) );
  NOR2_X1 U10723 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n8259) );
  NOR2_X2 U10724 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), 
        .ZN(n8513) );
  NOR2_X1 U10725 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), 
        .ZN(n8261) );
  AND2_X2 U10726 ( .A1(n7310), .A2(n14529), .ZN(n8311) );
  NAND2_X1 U10727 ( .A1(n8314), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8273) );
  NAND2_X1 U10728 ( .A1(n8312), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n8272) );
  AND2_X2 U10729 ( .A1(n8270), .A2(n14529), .ZN(n8310) );
  XNOR2_X2 U10730 ( .A(n8277), .B(n7288), .ZN(n12477) );
  NAND2_X4 U10731 ( .A1(n8705), .A2(n12477), .ZN(n10535) );
  OR2_X1 U10732 ( .A1(n8296), .A2(n10385), .ZN(n8280) );
  NAND2_X1 U10733 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8278) );
  NAND3_X2 U10734 ( .A1(n8280), .A2(n8279), .A3(n7605), .ZN(n10753) );
  XNOR2_X2 U10735 ( .A(n14170), .B(n10753), .ZN(n10749) );
  INV_X1 U10736 ( .A(n10749), .ZN(n8287) );
  NAND2_X1 U10737 ( .A1(n8312), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8284) );
  NAND2_X1 U10738 ( .A1(n8314), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8283) );
  NAND2_X1 U10739 ( .A1(n8310), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8282) );
  NAND2_X1 U10740 ( .A1(n8311), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8281) );
  NAND2_X1 U10741 ( .A1(n10046), .A2(SI_0_), .ZN(n8285) );
  XNOR2_X1 U10742 ( .A(n8285), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n14532) );
  MUX2_X1 U10743 ( .A(P2_IR_REG_0__SCAN_IN), .B(n14532), .S(n10535), .Z(n10746) );
  INV_X1 U10744 ( .A(n10746), .ZN(n10236) );
  NOR2_X1 U10745 ( .A1(n10576), .A2(n10236), .ZN(n10743) );
  NAND2_X1 U10746 ( .A1(n8287), .A2(n8286), .ZN(n10745) );
  INV_X1 U10747 ( .A(n14170), .ZN(n10554) );
  INV_X1 U10748 ( .A(n10753), .ZN(n15502) );
  NAND2_X1 U10749 ( .A1(n10554), .A2(n15502), .ZN(n8288) );
  NAND2_X1 U10750 ( .A1(n8311), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8292) );
  NAND2_X1 U10751 ( .A1(n8582), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n8291) );
  NAND2_X1 U10752 ( .A1(n8314), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8290) );
  NAND2_X1 U10753 ( .A1(n8310), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8289) );
  INV_X1 U10754 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n14522) );
  OR2_X1 U10755 ( .A1(n8293), .A2(n14522), .ZN(n8295) );
  NAND2_X1 U10756 ( .A1(n6675), .A2(n10400), .ZN(n8298) );
  OR2_X1 U10757 ( .A1(n8464), .A2(n10409), .ZN(n8297) );
  OAI211_X1 U10758 ( .C1(n10535), .C2(n10978), .A(n8298), .B(n8297), .ZN(
        n10243) );
  XNOR2_X2 U10759 ( .A(n14169), .B(n8299), .ZN(n10809) );
  NAND2_X1 U10760 ( .A1(n10806), .A2(n10809), .ZN(n10805) );
  INV_X1 U10761 ( .A(n14169), .ZN(n10577) );
  NAND2_X1 U10762 ( .A1(n10577), .A2(n8299), .ZN(n8300) );
  NAND2_X1 U10763 ( .A1(n10805), .A2(n8300), .ZN(n10847) );
  NAND2_X1 U10764 ( .A1(n8311), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8304) );
  INV_X1 U10765 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n11030) );
  NAND2_X1 U10766 ( .A1(n8312), .A2(n11030), .ZN(n8303) );
  NAND2_X1 U10767 ( .A1(n8314), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8302) );
  NAND2_X1 U10768 ( .A1(n8310), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n8301) );
  NAND2_X1 U10769 ( .A1(n10403), .A2(n8325), .ZN(n8308) );
  INV_X4 U10770 ( .A(n10535), .ZN(n8518) );
  NAND2_X1 U10771 ( .A1(n8305), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8306) );
  XNOR2_X1 U10772 ( .A(n8306), .B(P2_IR_REG_3__SCAN_IN), .ZN(n15356) );
  AOI22_X1 U10773 ( .A1(n8319), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n8518), .B2(
        n15356), .ZN(n8307) );
  NAND2_X2 U10774 ( .A1(n8308), .A2(n8307), .ZN(n10905) );
  XNOR2_X2 U10775 ( .A(n14167), .B(n11464), .ZN(n10851) );
  INV_X1 U10776 ( .A(n14167), .ZN(n8656) );
  NAND2_X1 U10777 ( .A1(n8656), .A2(n11464), .ZN(n8309) );
  NAND2_X1 U10778 ( .A1(n8405), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n8318) );
  NAND2_X1 U10779 ( .A1(n8311), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8317) );
  NAND2_X1 U10780 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8330) );
  OAI21_X1 U10781 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n8330), .ZN(n11009) );
  INV_X1 U10782 ( .A(n11009), .ZN(n8313) );
  NAND2_X1 U10783 ( .A1(n8582), .A2(n8313), .ZN(n8316) );
  INV_X2 U10784 ( .A(n8367), .ZN(n9855) );
  NAND2_X1 U10785 ( .A1(n9855), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8315) );
  NAND2_X1 U10786 ( .A1(n10423), .A2(n8325), .ZN(n8323) );
  NAND2_X1 U10787 ( .A1(n8320), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8321) );
  XNOR2_X1 U10788 ( .A(n8321), .B(P2_IR_REG_4__SCAN_IN), .ZN(n15369) );
  AOI22_X1 U10789 ( .A1(n8319), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n8518), .B2(
        n15369), .ZN(n8322) );
  NAND2_X1 U10790 ( .A1(n10996), .A2(n10999), .ZN(n10995) );
  OR2_X1 U10791 ( .A1(n14166), .A2(n11019), .ZN(n8324) );
  NAND2_X1 U10792 ( .A1(n10437), .A2(n8325), .ZN(n8329) );
  OR2_X1 U10793 ( .A1(n8326), .A2(n14522), .ZN(n8327) );
  XNOR2_X1 U10794 ( .A(n8327), .B(P2_IR_REG_5__SCAN_IN), .ZN(n15382) );
  AOI22_X1 U10795 ( .A1(n8319), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8518), .B2(
        n15382), .ZN(n8328) );
  INV_X1 U10796 ( .A(n11074), .ZN(n11127) );
  NAND2_X1 U10797 ( .A1(n8405), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8335) );
  NAND2_X1 U10798 ( .A1(n9856), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8334) );
  NOR2_X1 U10799 ( .A1(n8330), .A2(n10891), .ZN(n8341) );
  INV_X1 U10800 ( .A(n8341), .ZN(n8343) );
  NAND2_X1 U10801 ( .A1(n8330), .A2(n10891), .ZN(n8331) );
  AND2_X1 U10802 ( .A1(n8343), .A2(n8331), .ZN(n11125) );
  NAND2_X1 U10803 ( .A1(n8582), .A2(n11125), .ZN(n8333) );
  NAND2_X1 U10804 ( .A1(n9855), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8332) );
  NAND4_X1 U10805 ( .A1(n8335), .A2(n8334), .A3(n8333), .A4(n8332), .ZN(n14165) );
  INV_X1 U10806 ( .A(n14165), .ZN(n11228) );
  OAI21_X1 U10807 ( .B1(n11068), .B2(n11127), .A(n11228), .ZN(n8337) );
  NAND2_X1 U10808 ( .A1(n11068), .A2(n11127), .ZN(n8336) );
  NAND2_X1 U10809 ( .A1(n10443), .A2(n8325), .ZN(n8340) );
  NAND2_X1 U10810 ( .A1(n8639), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8338) );
  XNOR2_X1 U10811 ( .A(n8338), .B(P2_IR_REG_6__SCAN_IN), .ZN(n15394) );
  AOI22_X1 U10812 ( .A1(n8319), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8518), .B2(
        n15394), .ZN(n8339) );
  NAND2_X1 U10813 ( .A1(n9856), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8348) );
  NAND2_X1 U10814 ( .A1(n8405), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8347) );
  NAND2_X1 U10815 ( .A1(n8341), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8354) );
  INV_X1 U10816 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8342) );
  NAND2_X1 U10817 ( .A1(n8343), .A2(n8342), .ZN(n8344) );
  AND2_X1 U10818 ( .A1(n8354), .A2(n8344), .ZN(n11327) );
  NAND2_X1 U10819 ( .A1(n8582), .A2(n11327), .ZN(n8346) );
  NAND2_X1 U10820 ( .A1(n9855), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8345) );
  NAND4_X1 U10821 ( .A1(n8348), .A2(n8347), .A3(n8346), .A4(n8345), .ZN(n14164) );
  XNOR2_X1 U10822 ( .A(n11685), .B(n14164), .ZN(n11317) );
  NAND2_X1 U10823 ( .A1(n11685), .A2(n14164), .ZN(n8350) );
  NAND2_X1 U10824 ( .A1(n10452), .A2(n8325), .ZN(n8353) );
  NAND2_X1 U10825 ( .A1(n8363), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8351) );
  XNOR2_X1 U10826 ( .A(n8351), .B(P2_IR_REG_7__SCAN_IN), .ZN(n15407) );
  AOI22_X1 U10827 ( .A1(n8319), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8518), .B2(
        n15407), .ZN(n8352) );
  NAND2_X1 U10828 ( .A1(n8353), .A2(n8352), .ZN(n11088) );
  NAND2_X1 U10829 ( .A1(n8405), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8359) );
  NAND2_X1 U10830 ( .A1(n9856), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8358) );
  NAND2_X1 U10831 ( .A1(n8354), .A2(n11094), .ZN(n8355) );
  AND2_X1 U10832 ( .A1(n8369), .A2(n8355), .ZN(n11272) );
  NAND2_X1 U10833 ( .A1(n8582), .A2(n11272), .ZN(n8357) );
  NAND2_X1 U10834 ( .A1(n9855), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8356) );
  NAND4_X1 U10835 ( .A1(n8359), .A2(n8358), .A3(n8357), .A4(n8356), .ZN(n14163) );
  OR2_X1 U10836 ( .A1(n11088), .A2(n14163), .ZN(n8360) );
  NAND2_X1 U10837 ( .A1(n11088), .A2(n14163), .ZN(n8361) );
  NAND2_X1 U10838 ( .A1(n8362), .A2(n8361), .ZN(n11372) );
  NAND2_X1 U10839 ( .A1(n10458), .A2(n8325), .ZN(n8366) );
  NAND2_X1 U10840 ( .A1(n8378), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8364) );
  XNOR2_X1 U10841 ( .A(n8364), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10984) );
  AOI22_X1 U10842 ( .A1(n8319), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8518), .B2(
        n10984), .ZN(n8365) );
  NAND2_X1 U10843 ( .A1(n8311), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8374) );
  NAND2_X1 U10844 ( .A1(n9855), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8373) );
  NAND2_X1 U10845 ( .A1(n8369), .A2(n8368), .ZN(n8370) );
  NAND2_X1 U10846 ( .A1(n8385), .A2(n8370), .ZN(n11247) );
  INV_X1 U10847 ( .A(n11247), .ZN(n11383) );
  NAND2_X1 U10848 ( .A1(n8582), .A2(n11383), .ZN(n8372) );
  NAND2_X1 U10849 ( .A1(n8405), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8371) );
  NAND4_X1 U10850 ( .A1(n8374), .A2(n8373), .A3(n8372), .A4(n8371), .ZN(n14162) );
  INV_X1 U10851 ( .A(n14162), .ZN(n11093) );
  NAND2_X1 U10852 ( .A1(n15523), .A2(n11093), .ZN(n8667) );
  OR2_X1 U10853 ( .A1(n15523), .A2(n11093), .ZN(n8375) );
  NAND2_X1 U10854 ( .A1(n8667), .A2(n8375), .ZN(n10081) );
  NAND2_X1 U10855 ( .A1(n11372), .A2(n10081), .ZN(n8377) );
  NAND2_X1 U10856 ( .A1(n15523), .A2(n14162), .ZN(n8376) );
  NAND2_X1 U10857 ( .A1(n8377), .A2(n8376), .ZN(n11732) );
  NAND2_X1 U10858 ( .A1(n10515), .A2(n8325), .ZN(n8383) );
  INV_X1 U10859 ( .A(n8378), .ZN(n8380) );
  NAND2_X1 U10860 ( .A1(n8380), .A2(n8379), .ZN(n8395) );
  NAND2_X1 U10861 ( .A1(n8395), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8381) );
  XNOR2_X1 U10862 ( .A(n8381), .B(P2_IR_REG_9__SCAN_IN), .ZN(n11295) );
  AOI22_X1 U10863 ( .A1(n8319), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8518), .B2(
        n11295), .ZN(n8382) );
  NAND2_X1 U10864 ( .A1(n8405), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8390) );
  BUF_X2 U10865 ( .A(n8311), .Z(n9856) );
  NAND2_X1 U10866 ( .A1(n9856), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8389) );
  INV_X1 U10867 ( .A(n8401), .ZN(n8403) );
  NAND2_X1 U10868 ( .A1(n8385), .A2(n8384), .ZN(n8386) );
  AND2_X1 U10869 ( .A1(n8403), .A2(n8386), .ZN(n11742) );
  NAND2_X1 U10870 ( .A1(n8582), .A2(n11742), .ZN(n8388) );
  NAND2_X1 U10871 ( .A1(n9855), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8387) );
  NAND4_X1 U10872 ( .A1(n8390), .A2(n8389), .A3(n8388), .A4(n8387), .ZN(n14161) );
  INV_X1 U10873 ( .A(n14161), .ZN(n8391) );
  NAND2_X1 U10874 ( .A1(n11995), .A2(n8391), .ZN(n8668) );
  OR2_X1 U10875 ( .A1(n11995), .A2(n8391), .ZN(n8392) );
  NAND2_X1 U10876 ( .A1(n8668), .A2(n8392), .ZN(n11731) );
  NAND2_X1 U10877 ( .A1(n11732), .A2(n11731), .ZN(n8394) );
  NAND2_X1 U10878 ( .A1(n11995), .A2(n14161), .ZN(n8393) );
  NAND2_X1 U10879 ( .A1(n8394), .A2(n8393), .ZN(n11774) );
  NAND2_X1 U10880 ( .A1(n10581), .A2(n8325), .ZN(n8400) );
  INV_X1 U10881 ( .A(n8395), .ZN(n8397) );
  INV_X1 U10882 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8396) );
  NAND2_X1 U10883 ( .A1(n8397), .A2(n8396), .ZN(n8413) );
  NAND2_X1 U10884 ( .A1(n8413), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8398) );
  XNOR2_X1 U10885 ( .A(n8398), .B(P2_IR_REG_10__SCAN_IN), .ZN(n15433) );
  AOI22_X1 U10886 ( .A1(n8319), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n8518), 
        .B2(n15433), .ZN(n8399) );
  NAND2_X1 U10887 ( .A1(n9856), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8409) );
  NAND2_X1 U10888 ( .A1(n9855), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8408) );
  NAND2_X1 U10889 ( .A1(n8401), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8417) );
  INV_X1 U10890 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8402) );
  NAND2_X1 U10891 ( .A1(n8403), .A2(n8402), .ZN(n8404) );
  AND2_X1 U10892 ( .A1(n8417), .A2(n8404), .ZN(n11785) );
  NAND2_X1 U10893 ( .A1(n8582), .A2(n11785), .ZN(n8407) );
  NAND2_X1 U10894 ( .A1(n8405), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n8406) );
  NAND4_X1 U10895 ( .A1(n8409), .A2(n8408), .A3(n8407), .A4(n8406), .ZN(n14160) );
  INV_X1 U10896 ( .A(n14160), .ZN(n12108) );
  NAND2_X1 U10897 ( .A1(n15533), .A2(n12108), .ZN(n8669) );
  OR2_X1 U10898 ( .A1(n15533), .A2(n12108), .ZN(n8410) );
  NAND2_X1 U10899 ( .A1(n8669), .A2(n8410), .ZN(n10083) );
  NAND2_X1 U10900 ( .A1(n11774), .A2(n10083), .ZN(n8412) );
  NAND2_X1 U10901 ( .A1(n15533), .A2(n14160), .ZN(n8411) );
  NAND2_X1 U10902 ( .A1(n10681), .A2(n8325), .ZN(n8416) );
  OAI21_X1 U10903 ( .B1(n8413), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8414) );
  XNOR2_X1 U10904 ( .A(n8414), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11536) );
  AOI22_X1 U10905 ( .A1(n8319), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n11536), 
        .B2(n8518), .ZN(n8415) );
  NAND2_X1 U10906 ( .A1(n9856), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n8422) );
  NAND2_X1 U10907 ( .A1(n8417), .A2(n11303), .ZN(n8418) );
  AND2_X1 U10908 ( .A1(n8429), .A2(n8418), .ZN(n12114) );
  NAND2_X1 U10909 ( .A1(n8582), .A2(n12114), .ZN(n8421) );
  NAND2_X1 U10910 ( .A1(n9855), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8420) );
  NAND2_X1 U10911 ( .A1(n8405), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8419) );
  NAND4_X1 U10912 ( .A1(n8422), .A2(n8421), .A3(n8420), .A4(n8419), .ZN(n14159) );
  AND2_X1 U10913 ( .A1(n12257), .A2(n14159), .ZN(n8423) );
  NAND2_X1 U10914 ( .A1(n10736), .A2(n8325), .ZN(n8427) );
  OR2_X2 U10915 ( .A1(n8639), .A2(n8424), .ZN(n8436) );
  NAND2_X1 U10916 ( .A1(n8436), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8425) );
  XNOR2_X1 U10917 ( .A(n8425), .B(P2_IR_REG_12__SCAN_IN), .ZN(n11975) );
  AOI22_X1 U10918 ( .A1(n8319), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8518), 
        .B2(n11975), .ZN(n8426) );
  NAND2_X1 U10919 ( .A1(n8405), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n8434) );
  NAND2_X1 U10920 ( .A1(n9856), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8433) );
  INV_X1 U10921 ( .A(n8440), .ZN(n8442) );
  NAND2_X1 U10922 ( .A1(n8429), .A2(n8428), .ZN(n8430) );
  AND2_X1 U10923 ( .A1(n8442), .A2(n8430), .ZN(n12050) );
  NAND2_X1 U10924 ( .A1(n8582), .A2(n12050), .ZN(n8432) );
  NAND2_X1 U10925 ( .A1(n9855), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8431) );
  NAND4_X1 U10926 ( .A1(n8434), .A2(n8433), .A3(n8432), .A4(n8431), .ZN(n14158) );
  OR2_X1 U10927 ( .A1(n12051), .A2(n14158), .ZN(n10073) );
  INV_X1 U10928 ( .A(n10073), .ZN(n8435) );
  NAND2_X1 U10929 ( .A1(n12051), .A2(n14158), .ZN(n10072) );
  NAND2_X1 U10930 ( .A1(n10814), .A2(n8325), .ZN(n8439) );
  NOR2_X2 U10931 ( .A1(n8436), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n8451) );
  OR2_X1 U10932 ( .A1(n8451), .A2(n14522), .ZN(n8437) );
  XNOR2_X1 U10933 ( .A(n8437), .B(P2_IR_REG_13__SCAN_IN), .ZN(n12217) );
  AOI22_X1 U10934 ( .A1(n8319), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8518), 
        .B2(n12217), .ZN(n8438) );
  NAND2_X1 U10935 ( .A1(n8405), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8447) );
  NAND2_X1 U10936 ( .A1(n8311), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n8446) );
  NAND2_X1 U10937 ( .A1(n8440), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8456) );
  INV_X1 U10938 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8441) );
  NAND2_X1 U10939 ( .A1(n8442), .A2(n8441), .ZN(n8443) );
  AND2_X1 U10940 ( .A1(n8456), .A2(n8443), .ZN(n12079) );
  NAND2_X1 U10941 ( .A1(n8582), .A2(n12079), .ZN(n8445) );
  NAND2_X1 U10942 ( .A1(n9855), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8444) );
  NAND4_X1 U10943 ( .A1(n8447), .A2(n8446), .A3(n8445), .A4(n8444), .ZN(n14157) );
  AND2_X1 U10944 ( .A1(n12080), .A2(n14157), .ZN(n8449) );
  OR2_X1 U10945 ( .A1(n12080), .A2(n14157), .ZN(n8448) );
  OAI21_X1 U10946 ( .B1(n12073), .B2(n8449), .A(n8448), .ZN(n12316) );
  INV_X1 U10947 ( .A(n12316), .ZN(n8462) );
  NAND2_X1 U10948 ( .A1(n11045), .A2(n8325), .ZN(n8454) );
  INV_X1 U10949 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n8450) );
  NAND2_X1 U10950 ( .A1(n8451), .A2(n8450), .ZN(n8516) );
  NAND2_X1 U10951 ( .A1(n8516), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8452) );
  XNOR2_X1 U10952 ( .A(n8452), .B(P2_IR_REG_14__SCAN_IN), .ZN(n14184) );
  AOI22_X1 U10953 ( .A1(n8319), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8518), 
        .B2(n14184), .ZN(n8453) );
  NAND2_X1 U10954 ( .A1(n8405), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8461) );
  NAND2_X1 U10955 ( .A1(n9856), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n8460) );
  INV_X1 U10956 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8455) );
  NAND2_X1 U10957 ( .A1(n8456), .A2(n8455), .ZN(n8457) );
  AND2_X1 U10958 ( .A1(n8470), .A2(n8457), .ZN(n12320) );
  NAND2_X1 U10959 ( .A1(n8582), .A2(n12320), .ZN(n8459) );
  NAND2_X1 U10960 ( .A1(n9855), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8458) );
  NAND4_X1 U10961 ( .A1(n8461), .A2(n8460), .A3(n8459), .A4(n8458), .ZN(n14156) );
  OR2_X1 U10962 ( .A1(n12321), .A2(n14156), .ZN(n10069) );
  NAND2_X1 U10963 ( .A1(n8462), .A2(n10069), .ZN(n8463) );
  NAND2_X1 U10964 ( .A1(n12321), .A2(n14156), .ZN(n10068) );
  NAND2_X1 U10965 ( .A1(n8463), .A2(n10068), .ZN(n12370) );
  NAND2_X1 U10966 ( .A1(n11078), .A2(n8325), .ZN(n8469) );
  NAND2_X1 U10967 ( .A1(n8476), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8466) );
  INV_X1 U10968 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8465) );
  XNOR2_X1 U10969 ( .A(n8466), .B(n8465), .ZN(n15437) );
  OAI22_X1 U10970 ( .A1(n10056), .A2(n11079), .B1(n15437), .B2(n10535), .ZN(
        n8467) );
  INV_X1 U10971 ( .A(n8467), .ZN(n8468) );
  NAND2_X1 U10972 ( .A1(n8405), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8475) );
  NAND2_X1 U10973 ( .A1(n9856), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n8474) );
  INV_X1 U10974 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n12403) );
  INV_X1 U10975 ( .A(n8482), .ZN(n8484) );
  NAND2_X1 U10976 ( .A1(n8470), .A2(n12403), .ZN(n8471) );
  AND2_X1 U10977 ( .A1(n8484), .A2(n8471), .ZN(n12371) );
  NAND2_X1 U10978 ( .A1(n8582), .A2(n12371), .ZN(n8473) );
  NAND2_X1 U10979 ( .A1(n9855), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8472) );
  NAND4_X1 U10980 ( .A1(n8475), .A2(n8474), .A3(n8473), .A4(n8472), .ZN(n14155) );
  XNOR2_X1 U10981 ( .A(n12409), .B(n12485), .ZN(n12374) );
  NAND2_X1 U10982 ( .A1(n11021), .A2(n8325), .ZN(n8479) );
  NOR2_X1 U10983 ( .A1(n8476), .A2(P2_IR_REG_15__SCAN_IN), .ZN(n8489) );
  OR2_X1 U10984 ( .A1(n8489), .A2(n14522), .ZN(n8477) );
  XNOR2_X1 U10985 ( .A(n8477), .B(P2_IR_REG_16__SCAN_IN), .ZN(n15457) );
  AOI22_X1 U10986 ( .A1(n15457), .A2(n8518), .B1(n8319), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n8478) );
  NAND2_X1 U10987 ( .A1(n9856), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n8481) );
  NAND2_X1 U10988 ( .A1(n9855), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8480) );
  NAND2_X1 U10989 ( .A1(n8481), .A2(n8480), .ZN(n8487) );
  INV_X1 U10990 ( .A(n8493), .ZN(n8495) );
  INV_X1 U10991 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8483) );
  NAND2_X1 U10992 ( .A1(n8484), .A2(n8483), .ZN(n8485) );
  NAND2_X1 U10993 ( .A1(n8495), .A2(n8485), .ZN(n12500) );
  INV_X1 U10994 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n12489) );
  OAI22_X1 U10995 ( .A1(n12500), .A2(n8564), .B1(n8572), .B2(n12489), .ZN(
        n8486) );
  XNOR2_X1 U10996 ( .A(n14475), .B(n14154), .ZN(n12482) );
  NAND2_X1 U10997 ( .A1(n11063), .A2(n8325), .ZN(n8492) );
  INV_X1 U10998 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8488) );
  NAND2_X1 U10999 ( .A1(n8489), .A2(n8488), .ZN(n8500) );
  NAND2_X1 U11000 ( .A1(n8500), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8490) );
  XNOR2_X1 U11001 ( .A(n8490), .B(P2_IR_REG_17__SCAN_IN), .ZN(n15471) );
  AOI22_X1 U11002 ( .A1(n15471), .A2(n8518), .B1(n8319), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n8491) );
  INV_X1 U11003 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n14470) );
  INV_X1 U11004 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8494) );
  NAND2_X1 U11005 ( .A1(n8495), .A2(n8494), .ZN(n8496) );
  NAND2_X1 U11006 ( .A1(n8507), .A2(n8496), .ZN(n12566) );
  OR2_X1 U11007 ( .A1(n12566), .A2(n8564), .ZN(n8498) );
  AOI22_X1 U11008 ( .A1(n8405), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n9856), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n8497) );
  OAI211_X1 U11009 ( .C1(n8367), .C2(n14470), .A(n8498), .B(n8497), .ZN(n14153) );
  XNOR2_X1 U11010 ( .A(n12565), .B(n14129), .ZN(n12561) );
  AND2_X1 U11011 ( .A1(n12565), .A2(n14153), .ZN(n8499) );
  NAND2_X1 U11012 ( .A1(n11388), .A2(n8325), .ZN(n8505) );
  OAI21_X1 U11013 ( .B1(n8500), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8502) );
  INV_X1 U11014 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8501) );
  XNOR2_X1 U11015 ( .A(n8502), .B(n8501), .ZN(n15488) );
  INV_X1 U11016 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11391) );
  OAI22_X1 U11017 ( .A1(n15488), .A2(n10535), .B1(n10056), .B2(n11391), .ZN(
        n8503) );
  INV_X1 U11018 ( .A(n8503), .ZN(n8504) );
  NAND2_X2 U11019 ( .A1(n8505), .A2(n8504), .ZN(n14390) );
  INV_X1 U11020 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n15480) );
  INV_X1 U11021 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8506) );
  NAND2_X1 U11022 ( .A1(n8507), .A2(n8506), .ZN(n8508) );
  NAND2_X1 U11023 ( .A1(n8522), .A2(n8508), .ZN(n14386) );
  OR2_X1 U11024 ( .A1(n14386), .A2(n8564), .ZN(n8510) );
  AOI22_X1 U11025 ( .A1(n8405), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9856), .B2(
        P2_REG0_REG_18__SCAN_IN), .ZN(n8509) );
  OAI211_X1 U11026 ( .C1(n8367), .C2(n15480), .A(n8510), .B(n8509), .ZN(n14367) );
  INV_X1 U11027 ( .A(n14367), .ZN(n14071) );
  XNOR2_X1 U11028 ( .A(n14390), .B(n14071), .ZN(n14391) );
  NAND2_X1 U11029 ( .A1(n14384), .A2(n14391), .ZN(n14383) );
  OR2_X1 U11030 ( .A1(n14390), .A2(n14367), .ZN(n8511) );
  NAND2_X1 U11031 ( .A1(n14383), .A2(n8511), .ZN(n14363) );
  NAND2_X1 U11032 ( .A1(n11596), .A2(n8325), .ZN(n8520) );
  INV_X1 U11033 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8512) );
  NAND3_X1 U11034 ( .A1(n8514), .A2(n8513), .A3(n8512), .ZN(n8515) );
  XNOR2_X1 U11035 ( .A(n8517), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8650) );
  AOI22_X1 U11036 ( .A1(n8319), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n11007), 
        .B2(n8518), .ZN(n8519) );
  INV_X1 U11037 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8521) );
  NAND2_X1 U11038 ( .A1(n8522), .A2(n8521), .ZN(n8523) );
  NAND2_X1 U11039 ( .A1(n8544), .A2(n8523), .ZN(n14069) );
  INV_X1 U11040 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n14461) );
  NAND2_X1 U11041 ( .A1(n8311), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8525) );
  NAND2_X1 U11042 ( .A1(n8405), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8524) );
  OAI211_X1 U11043 ( .C1(n14461), .C2(n8367), .A(n8525), .B(n8524), .ZN(n8526)
         );
  INV_X1 U11044 ( .A(n8526), .ZN(n8527) );
  OAI21_X1 U11045 ( .B1(n14069), .B2(n8564), .A(n8527), .ZN(n14356) );
  NAND2_X1 U11046 ( .A1(n14375), .A2(n14356), .ZN(n8528) );
  OR2_X1 U11047 ( .A1(n14375), .A2(n14356), .ZN(n8529) );
  NAND2_X1 U11048 ( .A1(n11707), .A2(n8325), .ZN(n8531) );
  INV_X1 U11049 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11709) );
  OR2_X1 U11050 ( .A1(n10056), .A2(n11709), .ZN(n8530) );
  XNOR2_X1 U11051 ( .A(n8544), .B(P2_REG3_REG_20__SCAN_IN), .ZN(n14350) );
  NAND2_X1 U11052 ( .A1(n14350), .A2(n8582), .ZN(n8537) );
  INV_X1 U11053 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8534) );
  NAND2_X1 U11054 ( .A1(n9855), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8533) );
  NAND2_X1 U11055 ( .A1(n9856), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8532) );
  OAI211_X1 U11056 ( .C1(n8572), .C2(n8534), .A(n8533), .B(n8532), .ZN(n8535)
         );
  INV_X1 U11057 ( .A(n8535), .ZN(n8536) );
  NAND2_X1 U11058 ( .A1(n8537), .A2(n8536), .ZN(n14370) );
  NAND2_X1 U11059 ( .A1(n14454), .A2(n14370), .ZN(n8538) );
  NAND2_X1 U11060 ( .A1(n11813), .A2(n8325), .ZN(n8541) );
  OR2_X1 U11061 ( .A1(n10056), .A2(n11814), .ZN(n8540) );
  NAND2_X1 U11062 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(P2_REG3_REG_21__SCAN_IN), 
        .ZN(n8542) );
  INV_X1 U11063 ( .A(n8557), .ZN(n8546) );
  INV_X1 U11064 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n14119) );
  INV_X1 U11065 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8543) );
  OAI21_X1 U11066 ( .B1(n8544), .B2(n14119), .A(n8543), .ZN(n8545) );
  NAND2_X1 U11067 ( .A1(n14339), .A2(n8582), .ZN(n8552) );
  INV_X1 U11068 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8549) );
  NAND2_X1 U11069 ( .A1(n9856), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8548) );
  NAND2_X1 U11070 ( .A1(n9855), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8547) );
  OAI211_X1 U11071 ( .C1(n8572), .C2(n8549), .A(n8548), .B(n8547), .ZN(n8550)
         );
  INV_X1 U11072 ( .A(n8550), .ZN(n8551) );
  NAND2_X1 U11073 ( .A1(n8552), .A2(n8551), .ZN(n14355) );
  XNOR2_X1 U11074 ( .A(n14338), .B(n14355), .ZN(n14342) );
  XNOR2_X1 U11075 ( .A(n8554), .B(n8553), .ZN(n11998) );
  NAND2_X1 U11076 ( .A1(n11998), .A2(n8325), .ZN(n8556) );
  OR2_X1 U11077 ( .A1(n10056), .A2(n12000), .ZN(n8555) );
  NOR2_X1 U11078 ( .A1(n8557), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8558) );
  OR2_X1 U11079 ( .A1(n8567), .A2(n8558), .ZN(n14318) );
  INV_X1 U11080 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8561) );
  NAND2_X1 U11081 ( .A1(n9856), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8560) );
  NAND2_X1 U11082 ( .A1(n9855), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8559) );
  OAI211_X1 U11083 ( .C1(n8561), .C2(n8572), .A(n8560), .B(n8559), .ZN(n8562)
         );
  INV_X1 U11084 ( .A(n8562), .ZN(n8563) );
  XNOR2_X1 U11085 ( .A(n14443), .B(n14335), .ZN(n10090) );
  NAND2_X1 U11086 ( .A1(n12058), .A2(n8325), .ZN(n8566) );
  INV_X1 U11087 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n12061) );
  OR2_X1 U11088 ( .A1(n10056), .A2(n12061), .ZN(n8565) );
  OR2_X1 U11089 ( .A1(n8567), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8568) );
  NAND2_X1 U11090 ( .A1(n8567), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8579) );
  AND2_X1 U11091 ( .A1(n8568), .A2(n8579), .ZN(n14309) );
  NAND2_X1 U11092 ( .A1(n14309), .A2(n8582), .ZN(n8575) );
  INV_X1 U11093 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8571) );
  NAND2_X1 U11094 ( .A1(n9855), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8570) );
  NAND2_X1 U11095 ( .A1(n9856), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8569) );
  OAI211_X1 U11096 ( .C1(n8572), .C2(n8571), .A(n8570), .B(n8569), .ZN(n8573)
         );
  INV_X1 U11097 ( .A(n8573), .ZN(n8574) );
  XNOR2_X1 U11098 ( .A(n14306), .B(n14152), .ZN(n14297) );
  NAND2_X1 U11099 ( .A1(n12120), .A2(n8325), .ZN(n8577) );
  INV_X1 U11100 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n12122) );
  OR2_X1 U11101 ( .A1(n10056), .A2(n12122), .ZN(n8576) );
  NAND2_X1 U11102 ( .A1(n8405), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8586) );
  NAND2_X1 U11103 ( .A1(n9856), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8585) );
  INV_X1 U11104 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8578) );
  NAND2_X1 U11105 ( .A1(n8578), .A2(n8579), .ZN(n8581) );
  INV_X1 U11106 ( .A(n8579), .ZN(n8580) );
  NAND2_X1 U11107 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(n8580), .ZN(n8601) );
  AND2_X1 U11108 ( .A1(n8581), .A2(n8601), .ZN(n14290) );
  NAND2_X1 U11109 ( .A1(n8582), .A2(n14290), .ZN(n8584) );
  NAND2_X1 U11110 ( .A1(n9855), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8583) );
  NAND4_X1 U11111 ( .A1(n8586), .A2(n8585), .A3(n8584), .A4(n8583), .ZN(n14151) );
  INV_X1 U11112 ( .A(n14151), .ZN(n14268) );
  NAND2_X1 U11113 ( .A1(n14430), .A2(n14268), .ZN(n14263) );
  OR2_X1 U11114 ( .A1(n14430), .A2(n14268), .ZN(n8587) );
  NAND2_X1 U11115 ( .A1(n14263), .A2(n8587), .ZN(n14283) );
  INV_X1 U11116 ( .A(n14283), .ZN(n14278) );
  OR2_X2 U11117 ( .A1(n14279), .A2(n14278), .ZN(n14281) );
  NAND2_X1 U11118 ( .A1(n14430), .A2(n14151), .ZN(n8588) );
  NAND2_X1 U11119 ( .A1(n12165), .A2(n8325), .ZN(n8590) );
  OR2_X1 U11120 ( .A1(n10056), .A2(n12167), .ZN(n8589) );
  NAND2_X1 U11121 ( .A1(n8405), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8594) );
  NAND2_X1 U11122 ( .A1(n8311), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8593) );
  XNOR2_X1 U11123 ( .A(n8601), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n14272) );
  NAND2_X1 U11124 ( .A1(n8582), .A2(n14272), .ZN(n8592) );
  NAND2_X1 U11125 ( .A1(n9855), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8591) );
  NAND4_X1 U11126 ( .A1(n8594), .A2(n8593), .A3(n8592), .A4(n8591), .ZN(n14254) );
  INV_X1 U11127 ( .A(n14254), .ZN(n14286) );
  XNOR2_X1 U11128 ( .A(n14085), .B(n14286), .ZN(n14264) );
  INV_X1 U11129 ( .A(n14264), .ZN(n8691) );
  OR2_X1 U11130 ( .A1(n14085), .A2(n14254), .ZN(n8595) );
  NAND2_X1 U11131 ( .A1(n12384), .A2(n8325), .ZN(n8597) );
  OR2_X1 U11132 ( .A1(n10056), .A2(n12385), .ZN(n8596) );
  NAND2_X1 U11133 ( .A1(n8310), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8606) );
  NAND2_X1 U11134 ( .A1(n9856), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8605) );
  INV_X1 U11135 ( .A(n8601), .ZN(n8599) );
  AND2_X1 U11136 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(P2_REG3_REG_25__SCAN_IN), 
        .ZN(n8598) );
  NAND2_X1 U11137 ( .A1(n8599), .A2(n8598), .ZN(n8614) );
  INV_X1 U11138 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8600) );
  INV_X1 U11139 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n14138) );
  OAI21_X1 U11140 ( .B1(n8601), .B2(n8600), .A(n14138), .ZN(n8602) );
  AND2_X1 U11141 ( .A1(n8614), .A2(n8602), .ZN(n14247) );
  NAND2_X1 U11142 ( .A1(n8582), .A2(n14247), .ZN(n8604) );
  NAND2_X1 U11143 ( .A1(n9855), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8603) );
  NAND4_X1 U11144 ( .A1(n8606), .A2(n8605), .A3(n8604), .A4(n8603), .ZN(n14229) );
  NAND2_X1 U11145 ( .A1(n14420), .A2(n14229), .ZN(n8607) );
  OR2_X1 U11146 ( .A1(n14420), .A2(n14229), .ZN(n8608) );
  NAND2_X1 U11147 ( .A1(n12474), .A2(n8325), .ZN(n8611) );
  OR2_X1 U11148 ( .A1(n10056), .A2(n12479), .ZN(n8610) );
  NAND2_X1 U11149 ( .A1(n8405), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8619) );
  NAND2_X1 U11150 ( .A1(n9856), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8618) );
  INV_X1 U11151 ( .A(n8614), .ZN(n8612) );
  NAND2_X1 U11152 ( .A1(n8612), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8630) );
  INV_X1 U11153 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8613) );
  NAND2_X1 U11154 ( .A1(n8614), .A2(n8613), .ZN(n8615) );
  NAND2_X1 U11155 ( .A1(n8582), .A2(n14233), .ZN(n8617) );
  NAND2_X1 U11156 ( .A1(n9855), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8616) );
  NAND4_X1 U11157 ( .A1(n8619), .A2(n8618), .A3(n8617), .A4(n8616), .ZN(n14255) );
  NAND2_X1 U11158 ( .A1(n14415), .A2(n14255), .ZN(n8620) );
  INV_X1 U11159 ( .A(n8621), .ZN(n8624) );
  NOR2_X1 U11160 ( .A1(n8624), .A2(SI_27_), .ZN(n8622) );
  NAND2_X1 U11161 ( .A1(n8624), .A2(SI_27_), .ZN(n8625) );
  MUX2_X1 U11162 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n6676), .Z(n9847) );
  XNOR2_X1 U11163 ( .A(n9847), .B(SI_28_), .ZN(n9845) );
  NAND2_X1 U11164 ( .A1(n12494), .A2(n8325), .ZN(n8628) );
  INV_X1 U11165 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9260) );
  OR2_X1 U11166 ( .A1(n10056), .A2(n9260), .ZN(n8627) );
  NAND2_X1 U11167 ( .A1(n9856), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8635) );
  NAND2_X1 U11168 ( .A1(n9855), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8634) );
  INV_X1 U11169 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8629) );
  NAND2_X1 U11170 ( .A1(n8630), .A2(n8629), .ZN(n8631) );
  NAND2_X1 U11171 ( .A1(n8582), .A2(n12887), .ZN(n8633) );
  NAND2_X1 U11172 ( .A1(n8310), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8632) );
  NAND4_X1 U11173 ( .A1(n8635), .A2(n8634), .A3(n8633), .A4(n8632), .ZN(n14228) );
  NAND2_X1 U11174 ( .A1(n12892), .A2(n14228), .ZN(n9843) );
  OR2_X1 U11175 ( .A1(n12892), .A2(n14228), .ZN(n8636) );
  NAND2_X1 U11176 ( .A1(n9843), .A2(n8636), .ZN(n10092) );
  NAND2_X1 U11177 ( .A1(n9844), .A2(n8638), .ZN(n12857) );
  NAND2_X1 U11178 ( .A1(n8641), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8640) );
  AND2_X2 U11179 ( .A1(n11007), .A2(n11708), .ZN(n8741) );
  NAND2_X1 U11180 ( .A1(n8645), .A2(n8642), .ZN(n8648) );
  NAND2_X1 U11181 ( .A1(n8646), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8647) );
  NAND2_X1 U11182 ( .A1(n14434), .A2(n10234), .ZN(n15520) );
  INV_X1 U11183 ( .A(n10851), .ZN(n8655) );
  NAND2_X1 U11184 ( .A1(n10748), .A2(n10749), .ZN(n8652) );
  NAND2_X1 U11185 ( .A1(n10554), .A2(n10753), .ZN(n8651) );
  NAND2_X1 U11186 ( .A1(n8652), .A2(n8651), .ZN(n10808) );
  NAND2_X1 U11187 ( .A1(n10808), .A2(n10076), .ZN(n8654) );
  NAND2_X1 U11188 ( .A1(n10577), .A2(n10812), .ZN(n8653) );
  NAND2_X1 U11189 ( .A1(n8656), .A2(n10905), .ZN(n8657) );
  INV_X1 U11190 ( .A(n10999), .ZN(n8658) );
  NAND2_X1 U11191 ( .A1(n8659), .A2(n11019), .ZN(n8660) );
  NAND2_X1 U11192 ( .A1(n8661), .A2(n8660), .ZN(n11069) );
  XNOR2_X1 U11193 ( .A(n11074), .B(n14165), .ZN(n11070) );
  NAND2_X1 U11194 ( .A1(n11069), .A2(n11070), .ZN(n8663) );
  NAND2_X1 U11195 ( .A1(n11074), .A2(n11228), .ZN(n8662) );
  NAND2_X1 U11196 ( .A1(n8663), .A2(n8662), .ZN(n11316) );
  NAND2_X1 U11197 ( .A1(n11316), .A2(n11317), .ZN(n8665) );
  INV_X1 U11198 ( .A(n14164), .ZN(n11092) );
  NAND2_X1 U11199 ( .A1(n11685), .A2(n11092), .ZN(n8664) );
  NAND2_X1 U11200 ( .A1(n8665), .A2(n8664), .ZN(n11266) );
  INV_X1 U11201 ( .A(n14163), .ZN(n11229) );
  OR2_X1 U11202 ( .A1(n11088), .A2(n11229), .ZN(n10075) );
  NAND2_X1 U11203 ( .A1(n11266), .A2(n10075), .ZN(n8666) );
  NAND2_X1 U11204 ( .A1(n11088), .A2(n11229), .ZN(n10074) );
  NAND2_X1 U11205 ( .A1(n8666), .A2(n10074), .ZN(n11374) );
  INV_X1 U11206 ( .A(n10081), .ZN(n11375) );
  NAND2_X1 U11207 ( .A1(n11373), .A2(n8667), .ZN(n11734) );
  INV_X1 U11208 ( .A(n11731), .ZN(n11735) );
  NAND2_X1 U11209 ( .A1(n11734), .A2(n11735), .ZN(n11733) );
  NAND2_X1 U11210 ( .A1(n11733), .A2(n8668), .ZN(n11776) );
  INV_X1 U11211 ( .A(n10083), .ZN(n11777) );
  XNOR2_X1 U11212 ( .A(n12257), .B(n14159), .ZN(n12105) );
  INV_X1 U11213 ( .A(n14159), .ZN(n12043) );
  NAND2_X1 U11214 ( .A1(n12257), .A2(n12043), .ZN(n8670) );
  INV_X1 U11215 ( .A(n14158), .ZN(n12107) );
  OR2_X1 U11216 ( .A1(n12051), .A2(n12107), .ZN(n8671) );
  NAND2_X1 U11217 ( .A1(n12051), .A2(n12107), .ZN(n8672) );
  INV_X1 U11218 ( .A(n14157), .ZN(n12314) );
  NAND2_X1 U11219 ( .A1(n12080), .A2(n12314), .ZN(n10070) );
  INV_X1 U11220 ( .A(n10070), .ZN(n8673) );
  OR2_X1 U11221 ( .A1(n12080), .A2(n12314), .ZN(n10071) );
  INV_X1 U11222 ( .A(n14156), .ZN(n12406) );
  NOR2_X1 U11223 ( .A1(n12321), .A2(n12406), .ZN(n8675) );
  NAND2_X1 U11224 ( .A1(n12321), .A2(n12406), .ZN(n8674) );
  AND2_X1 U11225 ( .A1(n12409), .A2(n12485), .ZN(n8676) );
  OR2_X1 U11226 ( .A1(n12409), .A2(n12485), .ZN(n8677) );
  INV_X1 U11227 ( .A(n14154), .ZN(n12405) );
  OR2_X1 U11228 ( .A1(n12565), .A2(n14129), .ZN(n8679) );
  INV_X1 U11229 ( .A(n14392), .ZN(n8682) );
  AND2_X1 U11230 ( .A1(n14390), .A2(n14071), .ZN(n8680) );
  INV_X1 U11231 ( .A(n8680), .ZN(n8681) );
  OR2_X1 U11232 ( .A1(n14390), .A2(n14071), .ZN(n8683) );
  INV_X1 U11233 ( .A(n14356), .ZN(n14130) );
  NAND2_X1 U11234 ( .A1(n14375), .A2(n14130), .ZN(n8685) );
  OR2_X1 U11235 ( .A1(n14375), .A2(n14130), .ZN(n8684) );
  NAND2_X1 U11236 ( .A1(n8685), .A2(n8684), .ZN(n14365) );
  INV_X1 U11237 ( .A(n14370), .ZN(n14070) );
  NAND2_X1 U11238 ( .A1(n14454), .A2(n14070), .ZN(n8687) );
  OR2_X1 U11239 ( .A1(n14454), .A2(n14070), .ZN(n8686) );
  NAND2_X1 U11240 ( .A1(n8687), .A2(n8686), .ZN(n10088) );
  NAND2_X1 U11241 ( .A1(n14353), .A2(n14354), .ZN(n14352) );
  NAND2_X1 U11242 ( .A1(n14352), .A2(n8687), .ZN(n14334) );
  NAND2_X1 U11243 ( .A1(n14334), .A2(n14342), .ZN(n14333) );
  INV_X1 U11244 ( .A(n14355), .ZN(n14324) );
  NAND2_X1 U11245 ( .A1(n14338), .A2(n14324), .ZN(n8688) );
  INV_X1 U11246 ( .A(n14335), .ZN(n8689) );
  OR2_X1 U11247 ( .A1(n14443), .A2(n8689), .ZN(n8690) );
  INV_X1 U11248 ( .A(n14297), .ZN(n14299) );
  NAND2_X1 U11249 ( .A1(n14306), .A2(n14326), .ZN(n14282) );
  OR2_X1 U11250 ( .A1(n14283), .A2(n14282), .ZN(n14261) );
  NAND2_X1 U11251 ( .A1(n8692), .A2(n8691), .ZN(n14266) );
  NAND2_X1 U11252 ( .A1(n14085), .A2(n14286), .ZN(n14250) );
  NAND2_X1 U11253 ( .A1(n14266), .A2(n14250), .ZN(n8694) );
  INV_X1 U11254 ( .A(n14229), .ZN(n14269) );
  NAND2_X1 U11255 ( .A1(n14420), .A2(n14269), .ZN(n14225) );
  OR2_X1 U11256 ( .A1(n14420), .A2(n14269), .ZN(n8693) );
  NAND2_X1 U11257 ( .A1(n14225), .A2(n8693), .ZN(n14251) );
  INV_X1 U11258 ( .A(n14251), .ZN(n14242) );
  NAND2_X1 U11259 ( .A1(n14253), .A2(n14225), .ZN(n8695) );
  INV_X1 U11260 ( .A(n14255), .ZN(n14141) );
  OR2_X1 U11261 ( .A1(n14201), .A2(n8713), .ZN(n8699) );
  NOR2_X1 U11262 ( .A1(n8697), .A2(n11708), .ZN(n10111) );
  INV_X1 U11263 ( .A(n10111), .ZN(n8698) );
  NAND2_X1 U11264 ( .A1(n9856), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8704) );
  NAND2_X1 U11265 ( .A1(n9855), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8703) );
  INV_X1 U11266 ( .A(n8700), .ZN(n14217) );
  NAND2_X1 U11267 ( .A1(n8582), .A2(n14217), .ZN(n8702) );
  NAND2_X1 U11268 ( .A1(n8310), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8701) );
  NAND4_X1 U11269 ( .A1(n8704), .A2(n8703), .A3(n8702), .A4(n8701), .ZN(n14150) );
  INV_X1 U11270 ( .A(n8697), .ZN(n10098) );
  NAND2_X1 U11271 ( .A1(n14150), .A2(n14369), .ZN(n8708) );
  INV_X1 U11272 ( .A(n8705), .ZN(n8706) );
  NAND2_X1 U11273 ( .A1(n14255), .A2(n14368), .ZN(n8707) );
  NAND2_X1 U11274 ( .A1(n8708), .A2(n8707), .ZN(n12888) );
  INV_X1 U11275 ( .A(n12888), .ZN(n8709) );
  OAI21_X1 U11276 ( .B1(n9852), .B2(n8710), .A(n8709), .ZN(n12854) );
  INV_X1 U11277 ( .A(n12080), .ZN(n12246) );
  INV_X1 U11278 ( .A(n11995), .ZN(n11992) );
  OR2_X1 U11279 ( .A1(n10753), .A2(n10746), .ZN(n10807) );
  AND2_X1 U11280 ( .A1(n10848), .A2(n11464), .ZN(n11004) );
  INV_X1 U11281 ( .A(n11019), .ZN(n11459) );
  NAND2_X1 U11282 ( .A1(n11004), .A2(n11459), .ZN(n11073) );
  INV_X1 U11283 ( .A(n11685), .ZN(n11329) );
  NAND2_X1 U11284 ( .A1(n11992), .A2(n11739), .ZN(n11782) );
  INV_X1 U11285 ( .A(n14443), .ZN(n14321) );
  INV_X1 U11286 ( .A(n14420), .ZN(n14249) );
  NAND2_X1 U11287 ( .A1(n14231), .A2(n12892), .ZN(n8714) );
  NAND2_X1 U11288 ( .A1(n8714), .A2(n14398), .ZN(n8715) );
  NOR2_X1 U11289 ( .A1(n9865), .A2(n8715), .ZN(n12856) );
  NOR2_X1 U11290 ( .A1(n12854), .A2(n12856), .ZN(n8716) );
  OAI21_X1 U11291 ( .B1(n12857), .B2(n14478), .A(n8716), .ZN(n9837) );
  NOR2_X1 U11292 ( .A1(n8639), .A2(n8717), .ZN(n8744) );
  NAND2_X1 U11293 ( .A1(n8744), .A2(n6991), .ZN(n8719) );
  NAND2_X1 U11294 ( .A1(n8719), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8718) );
  MUX2_X1 U11295 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8718), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n8721) );
  INV_X1 U11296 ( .A(n8719), .ZN(n8720) );
  NAND2_X1 U11297 ( .A1(n8720), .A2(n6992), .ZN(n8722) );
  NAND2_X1 U11298 ( .A1(n8721), .A2(n8722), .ZN(n12121) );
  XNOR2_X1 U11299 ( .A(n12121), .B(P2_B_REG_SCAN_IN), .ZN(n8725) );
  NAND2_X1 U11300 ( .A1(n8722), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8723) );
  MUX2_X1 U11301 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8723), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8724) );
  NAND2_X1 U11302 ( .A1(n8724), .A2(n6811), .ZN(n12166) );
  NAND2_X1 U11303 ( .A1(n8725), .A2(n12166), .ZN(n8729) );
  NAND2_X1 U11304 ( .A1(n6811), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8726) );
  MUX2_X1 U11305 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8726), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8728) );
  NAND2_X1 U11306 ( .A1(n8728), .A2(n8727), .ZN(n12386) );
  INV_X1 U11307 ( .A(n12386), .ZN(n8750) );
  NOR4_X1 U11308 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n8738) );
  OR4_X1 U11309 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n8735) );
  NOR4_X1 U11310 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n8733) );
  NOR4_X1 U11311 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n8732) );
  NOR4_X1 U11312 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8731) );
  NOR4_X1 U11313 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n8730) );
  NAND4_X1 U11314 ( .A1(n8733), .A2(n8732), .A3(n8731), .A4(n8730), .ZN(n8734)
         );
  NOR4_X1 U11315 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n8735), .A4(n8734), .ZN(n8737) );
  NOR4_X1 U11316 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n8736) );
  NAND3_X1 U11317 ( .A1(n8738), .A2(n8737), .A3(n8736), .ZN(n8739) );
  AND2_X1 U11318 ( .A1(n15508), .A2(n8739), .ZN(n10331) );
  INV_X1 U11319 ( .A(n10347), .ZN(n10141) );
  NAND2_X1 U11320 ( .A1(n10141), .A2(n10534), .ZN(n10342) );
  INV_X1 U11321 ( .A(n10342), .ZN(n8740) );
  OR2_X1 U11322 ( .A1(n10331), .A2(n8740), .ZN(n10705) );
  NAND2_X1 U11323 ( .A1(n8741), .A2(n10336), .ZN(n10340) );
  INV_X1 U11324 ( .A(n10340), .ZN(n10338) );
  NOR2_X1 U11325 ( .A1(n10705), .A2(n10338), .ZN(n8748) );
  INV_X1 U11326 ( .A(n12166), .ZN(n8743) );
  NOR2_X1 U11327 ( .A1(n12121), .A2(n12386), .ZN(n8742) );
  NAND2_X1 U11328 ( .A1(n8743), .A2(n8742), .ZN(n10231) );
  OR2_X1 U11329 ( .A1(n8744), .A2(n14522), .ZN(n8745) );
  XNOR2_X1 U11330 ( .A(n8745), .B(n6991), .ZN(n10533) );
  AND2_X1 U11331 ( .A1(n10231), .A2(n10533), .ZN(n10343) );
  INV_X1 U11332 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15515) );
  NAND2_X1 U11333 ( .A1(n15508), .A2(n15515), .ZN(n8747) );
  NAND2_X1 U11334 ( .A1(n12166), .A2(n12386), .ZN(n8746) );
  NAND2_X1 U11335 ( .A1(n8747), .A2(n8746), .ZN(n10706) );
  AND2_X1 U11336 ( .A1(n15512), .A2(n10706), .ZN(n15513) );
  INV_X1 U11337 ( .A(n12121), .ZN(n8751) );
  INV_X1 U11338 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15510) );
  NAND2_X1 U11339 ( .A1(n15508), .A2(n15510), .ZN(n8749) );
  NAND2_X1 U11340 ( .A1(n10141), .A2(n10336), .ZN(n15525) );
  INV_X1 U11341 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8752) );
  AOI21_X1 U11342 ( .B1(n9837), .B2(n15543), .A(n8754), .ZN(n8755) );
  NOR2_X2 U11343 ( .A1(n8854), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n8873) );
  NAND2_X1 U11344 ( .A1(n8873), .A2(n8758), .ZN(n8884) );
  INV_X1 U11345 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8764) );
  NAND2_X1 U11346 ( .A1(n9332), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8765) );
  XNOR2_X2 U11347 ( .A(n8765), .B(n8779), .ZN(n11252) );
  INV_X1 U11348 ( .A(n8766), .ZN(n8767) );
  NAND2_X1 U11349 ( .A1(n8767), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8768) );
  NAND2_X1 U11350 ( .A1(n8769), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8770) );
  OAI21_X1 U11351 ( .B1(n11252), .B2(n9374), .A(n13666), .ZN(n8774) );
  INV_X1 U11352 ( .A(n8771), .ZN(n8772) );
  NAND2_X1 U11353 ( .A1(n8772), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8773) );
  XNOR2_X2 U11354 ( .A(n8773), .B(n8780), .ZN(n11160) );
  NAND2_X1 U11355 ( .A1(n8774), .A2(n11160), .ZN(n8776) );
  OAI21_X1 U11356 ( .B1(n9374), .B2(n13173), .A(n11252), .ZN(n8775) );
  NAND2_X1 U11357 ( .A1(n8776), .A2(n8775), .ZN(n11109) );
  INV_X1 U11358 ( .A(n11163), .ZN(n13347) );
  AND2_X1 U11359 ( .A1(n15719), .A2(n13347), .ZN(n8777) );
  NAND2_X1 U11360 ( .A1(n11109), .A2(n8777), .ZN(n8778) );
  OR3_X1 U11361 ( .A1(n11252), .A2(n13666), .A3(n11159), .ZN(n9366) );
  NAND2_X1 U11362 ( .A1(n11252), .A2(n11501), .ZN(n10182) );
  NOR2_X1 U11363 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), 
        .ZN(n8782) );
  NAND2_X1 U11364 ( .A1(n8787), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8789) );
  INV_X1 U11365 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n11177) );
  INV_X1 U11366 ( .A(n13379), .ZN(n8790) );
  INV_X1 U11367 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n11678) );
  NAND2_X1 U11368 ( .A1(n8792), .A2(n8791), .ZN(n8793) );
  NOR2_X1 U11369 ( .A1(n8793), .A2(n7581), .ZN(n8796) );
  INV_X1 U11370 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10871) );
  OR2_X1 U11371 ( .A1(n8916), .A2(n10871), .ZN(n8795) );
  BUF_X2 U11372 ( .A(n8835), .Z(n10856) );
  OR2_X1 U11373 ( .A1(n8980), .A2(n10378), .ZN(n8801) );
  XNOR2_X1 U11374 ( .A(n8816), .B(n8814), .ZN(n10379) );
  NAND2_X1 U11375 ( .A1(n10856), .A2(n6728), .ZN(n8800) );
  NAND2_X1 U11376 ( .A1(n9321), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8805) );
  NAND2_X1 U11377 ( .A1(n8841), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8804) );
  INV_X1 U11378 ( .A(n8843), .ZN(n8915) );
  NAND2_X1 U11379 ( .A1(n8915), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8803) );
  NAND2_X1 U11380 ( .A1(n9189), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8802) );
  OR2_X1 U11381 ( .A1(n8980), .A2(n9810), .ZN(n8810) );
  NAND2_X4 U11382 ( .A1(n8835), .A2(n8806), .ZN(n9145) );
  NAND2_X1 U11383 ( .A1(n8807), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8808) );
  AND2_X1 U11384 ( .A1(n8814), .A2(n8808), .ZN(n10416) );
  OR2_X1 U11385 ( .A1(n9145), .A2(n10416), .ZN(n8809) );
  NAND2_X1 U11386 ( .A1(n11166), .A2(n13174), .ZN(n15688) );
  NAND2_X1 U11387 ( .A1(n8915), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8813) );
  NAND2_X1 U11388 ( .A1(n8841), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8812) );
  NAND2_X1 U11389 ( .A1(n9189), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8811) );
  NAND2_X1 U11390 ( .A1(n8816), .A2(n8815), .ZN(n8818) );
  NAND2_X1 U11391 ( .A1(n10384), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8817) );
  NAND2_X1 U11392 ( .A1(n8818), .A2(n8817), .ZN(n8829) );
  NAND2_X1 U11393 ( .A1(n10409), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8830) );
  NAND2_X1 U11394 ( .A1(n10402), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8819) );
  XNOR2_X1 U11395 ( .A(n8829), .B(n8828), .ZN(n10394) );
  NAND2_X1 U11396 ( .A1(n10856), .A2(n6729), .ZN(n8820) );
  OR2_X1 U11397 ( .A1(n8980), .A2(SI_2_), .ZN(n8821) );
  NAND2_X1 U11398 ( .A1(n15688), .A2(n15687), .ZN(n15686) );
  OR2_X1 U11399 ( .A1(n9273), .A2(n15697), .ZN(n13179) );
  NAND2_X1 U11400 ( .A1(n15686), .A2(n13179), .ZN(n11491) );
  NAND2_X1 U11401 ( .A1(n8841), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8827) );
  INV_X1 U11402 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n11852) );
  OR2_X1 U11403 ( .A1(n8860), .A2(n11852), .ZN(n8826) );
  OR2_X1 U11404 ( .A1(n8843), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n8825) );
  AND4_X2 U11405 ( .A1(n8827), .A2(n8826), .A3(n8825), .A4(n8824), .ZN(n8839)
         );
  OR2_X1 U11406 ( .A1(n8980), .A2(SI_3_), .ZN(n8838) );
  NAND2_X1 U11407 ( .A1(n8829), .A2(n8828), .ZN(n8831) );
  NAND2_X1 U11408 ( .A1(n8831), .A2(n8830), .ZN(n8850) );
  NAND2_X1 U11409 ( .A1(n10407), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8851) );
  NAND2_X1 U11410 ( .A1(n10404), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8832) );
  XNOR2_X1 U11411 ( .A(n8850), .B(n8849), .ZN(n10410) );
  OR2_X1 U11412 ( .A1(n9145), .A2(n10410), .ZN(n8837) );
  NAND2_X1 U11413 ( .A1(n8833), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8834) );
  XNOR2_X1 U11414 ( .A(n8834), .B(P3_IR_REG_3__SCAN_IN), .ZN(n15561) );
  OR2_X1 U11415 ( .A1(n8835), .A2(n15561), .ZN(n8836) );
  NAND2_X1 U11416 ( .A1(n8839), .A2(n11287), .ZN(n13189) );
  INV_X1 U11417 ( .A(n11287), .ZN(n15713) );
  NAND2_X1 U11418 ( .A1(n6679), .A2(n15713), .ZN(n13184) );
  NAND2_X1 U11419 ( .A1(n11491), .A2(n13319), .ZN(n8840) );
  NAND2_X1 U11420 ( .A1(n8840), .A2(n13189), .ZN(n11393) );
  NAND2_X1 U11421 ( .A1(n9321), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8848) );
  INV_X1 U11422 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n8842) );
  OR2_X1 U11423 ( .A1(n9030), .A2(n8842), .ZN(n8847) );
  AND2_X1 U11424 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8844) );
  NOR2_X1 U11425 ( .A1(n8861), .A2(n8844), .ZN(n11817) );
  OR2_X1 U11426 ( .A1(n9134), .A2(n11817), .ZN(n8846) );
  INV_X1 U11427 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n11856) );
  OR2_X1 U11428 ( .A1(n8916), .A2(n11856), .ZN(n8845) );
  OR2_X1 U11429 ( .A1(n8980), .A2(SI_4_), .ZN(n8858) );
  NAND2_X1 U11430 ( .A1(n8850), .A2(n8849), .ZN(n8852) );
  NAND2_X1 U11431 ( .A1(n8852), .A2(n8851), .ZN(n8869) );
  NAND2_X1 U11432 ( .A1(n10427), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8870) );
  NAND2_X1 U11433 ( .A1(n10424), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8853) );
  XNOR2_X1 U11434 ( .A(n8869), .B(n8868), .ZN(n10380) );
  OR2_X1 U11435 ( .A1(n9145), .A2(n10380), .ZN(n8857) );
  NAND2_X1 U11436 ( .A1(n8854), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8855) );
  XNOR2_X1 U11437 ( .A(n8855), .B(P3_IR_REG_4__SCAN_IN), .ZN(n15578) );
  OR2_X1 U11438 ( .A1(n10856), .A2(n15578), .ZN(n8856) );
  NAND2_X1 U11439 ( .A1(n9282), .A2(n11578), .ZN(n13192) );
  INV_X1 U11440 ( .A(n9282), .ZN(n8859) );
  NAND2_X1 U11441 ( .A1(n8859), .A2(n11818), .ZN(n13193) );
  NAND2_X1 U11442 ( .A1(n13192), .A2(n13193), .ZN(n11397) );
  NAND2_X1 U11443 ( .A1(n11393), .A2(n9280), .ZN(n11392) );
  NAND2_X1 U11444 ( .A1(n11392), .A2(n13192), .ZN(n11698) );
  NAND2_X1 U11445 ( .A1(n8841), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8867) );
  INV_X1 U11446 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n11862) );
  OR2_X1 U11447 ( .A1(n8860), .A2(n11862), .ZN(n8866) );
  NAND2_X1 U11448 ( .A1(n8861), .A2(n8862), .ZN(n8878) );
  OR2_X1 U11449 ( .A1(n8862), .A2(n8861), .ZN(n8863) );
  AND2_X1 U11450 ( .A1(n8878), .A2(n8863), .ZN(n11699) );
  OR2_X1 U11451 ( .A1(n9134), .A2(n11699), .ZN(n8865) );
  INV_X1 U11452 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15601) );
  OR2_X1 U11453 ( .A1(n8916), .A2(n15601), .ZN(n8864) );
  OR2_X1 U11454 ( .A1(n8980), .A2(SI_5_), .ZN(n8877) );
  NAND2_X1 U11455 ( .A1(n8869), .A2(n8868), .ZN(n8871) );
  NAND2_X1 U11456 ( .A1(n8871), .A2(n8870), .ZN(n8888) );
  NAND2_X1 U11457 ( .A1(n10441), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8872) );
  XNOR2_X1 U11458 ( .A(n8888), .B(n8887), .ZN(n10386) );
  OR2_X1 U11459 ( .A1(n9145), .A2(n10386), .ZN(n8876) );
  OR2_X1 U11460 ( .A1(n8873), .A2(n14040), .ZN(n8874) );
  XNOR2_X1 U11461 ( .A(n8874), .B(P3_IR_REG_5__SCAN_IN), .ZN(n15599) );
  OR2_X1 U11462 ( .A1(n10856), .A2(n15599), .ZN(n8875) );
  NAND2_X1 U11463 ( .A1(n12007), .A2(n11660), .ZN(n13191) );
  INV_X1 U11464 ( .A(n12007), .ZN(n11949) );
  NAND2_X1 U11465 ( .A1(n11949), .A2(n11795), .ZN(n13200) );
  NAND2_X1 U11466 ( .A1(n11698), .A2(n13316), .ZN(n11697) );
  NAND2_X1 U11467 ( .A1(n11697), .A2(n13191), .ZN(n12002) );
  NAND2_X1 U11468 ( .A1(n8841), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8883) );
  INV_X1 U11469 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11868) );
  OR2_X1 U11470 ( .A1(n8860), .A2(n11868), .ZN(n8882) );
  NAND2_X1 U11471 ( .A1(n8878), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8879) );
  AND2_X1 U11472 ( .A1(n8894), .A2(n8879), .ZN(n12003) );
  OR2_X1 U11473 ( .A1(n9134), .A2(n12003), .ZN(n8881) );
  INV_X1 U11474 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n11867) );
  OR2_X1 U11475 ( .A1(n8916), .A2(n11867), .ZN(n8880) );
  NAND2_X1 U11476 ( .A1(n8885), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8886) );
  XNOR2_X1 U11477 ( .A(n8886), .B(P3_IR_REG_6__SCAN_IN), .ZN(n11897) );
  INV_X1 U11478 ( .A(SI_6_), .ZN(n10418) );
  OR2_X1 U11479 ( .A1(n8980), .A2(n10418), .ZN(n8893) );
  NAND2_X1 U11480 ( .A1(n8888), .A2(n8887), .ZN(n8890) );
  XNOR2_X1 U11481 ( .A(n10445), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n8891) );
  XNOR2_X1 U11482 ( .A(n8901), .B(n8891), .ZN(n10419) );
  OR2_X1 U11483 ( .A1(n9145), .A2(n10419), .ZN(n8892) );
  OAI211_X1 U11484 ( .C1(n10856), .C2(n15615), .A(n8893), .B(n8892), .ZN(
        n11958) );
  NAND2_X1 U11485 ( .A1(n12028), .A2(n11958), .ZN(n13202) );
  INV_X1 U11486 ( .A(n12028), .ZN(n13534) );
  INV_X1 U11487 ( .A(n11958), .ZN(n15720) );
  NAND2_X1 U11488 ( .A1(n13534), .A2(n15720), .ZN(n13201) );
  NAND2_X1 U11489 ( .A1(n13202), .A2(n13201), .ZN(n12005) );
  INV_X1 U11490 ( .A(n12005), .ZN(n13322) );
  NAND2_X1 U11491 ( .A1(n12002), .A2(n13322), .ZN(n12001) );
  NAND2_X1 U11492 ( .A1(n9266), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8899) );
  INV_X1 U11493 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11874) );
  OR2_X1 U11494 ( .A1(n8860), .A2(n11874), .ZN(n8898) );
  NOR2_X2 U11495 ( .A1(n8894), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8913) );
  AND2_X1 U11496 ( .A1(n8894), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8895) );
  NOR2_X1 U11497 ( .A1(n8913), .A2(n8895), .ZN(n12033) );
  OR2_X1 U11498 ( .A1(n9134), .A2(n12033), .ZN(n8897) );
  INV_X1 U11499 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n11873) );
  OR2_X1 U11500 ( .A1(n11521), .A2(n11873), .ZN(n8896) );
  OR2_X1 U11501 ( .A1(n8980), .A2(SI_7_), .ZN(n8912) );
  NAND2_X1 U11502 ( .A1(n10447), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8900) );
  NAND2_X1 U11503 ( .A1(n10445), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8902) );
  NAND2_X1 U11504 ( .A1(n10453), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8904) );
  NAND2_X1 U11505 ( .A1(n8923), .A2(n8904), .ZN(n8905) );
  NAND2_X1 U11506 ( .A1(n8906), .A2(n8905), .ZN(n8907) );
  AND2_X1 U11507 ( .A1(n8924), .A2(n8907), .ZN(n10389) );
  OR2_X1 U11508 ( .A1(n9145), .A2(n10389), .ZN(n8911) );
  OR2_X1 U11509 ( .A1(n8885), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n8921) );
  NAND2_X1 U11510 ( .A1(n8921), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8909) );
  INV_X1 U11511 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8908) );
  XNOR2_X1 U11512 ( .A(n8909), .B(n8908), .ZN(n15633) );
  INV_X1 U11513 ( .A(n15633), .ZN(n11875) );
  OR2_X1 U11514 ( .A1(n10856), .A2(n11875), .ZN(n8910) );
  NAND2_X1 U11515 ( .A1(n12155), .A2(n12030), .ZN(n13206) );
  INV_X1 U11516 ( .A(n12155), .ZN(n10765) );
  NAND2_X1 U11517 ( .A1(n10765), .A2(n11945), .ZN(n13207) );
  NAND2_X1 U11518 ( .A1(n13206), .A2(n13207), .ZN(n12023) );
  INV_X1 U11519 ( .A(n12023), .ZN(n13317) );
  INV_X1 U11520 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n12161) );
  OR2_X1 U11521 ( .A1(n8860), .A2(n12161), .ZN(n8920) );
  NAND2_X1 U11522 ( .A1(n9266), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8919) );
  NOR2_X1 U11523 ( .A1(n8913), .A2(n12129), .ZN(n8914) );
  OR2_X1 U11524 ( .A1(n8932), .A2(n8914), .ZN(n12158) );
  NAND2_X1 U11525 ( .A1(n8915), .A2(n12158), .ZN(n8918) );
  INV_X1 U11526 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n11879) );
  OR2_X1 U11527 ( .A1(n8916), .A2(n11879), .ZN(n8917) );
  NAND4_X1 U11528 ( .A1(n8920), .A2(n8919), .A3(n8918), .A4(n8917), .ZN(n13533) );
  NAND2_X1 U11529 ( .A1(n8938), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8922) );
  XNOR2_X1 U11530 ( .A(n8922), .B(P3_IR_REG_8__SCAN_IN), .ZN(n11896) );
  INV_X1 U11531 ( .A(SI_8_), .ZN(n10392) );
  NAND2_X1 U11532 ( .A1(n10459), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8944) );
  NAND2_X1 U11533 ( .A1(n10461), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8925) );
  OR2_X1 U11534 ( .A1(n8927), .A2(n8926), .ZN(n8928) );
  NAND2_X1 U11535 ( .A1(n8945), .A2(n8928), .ZN(n10393) );
  OR2_X1 U11536 ( .A1(n9145), .A2(n10393), .ZN(n8929) );
  OAI211_X1 U11537 ( .C1(n10856), .C2(n15649), .A(n8930), .B(n8929), .ZN(
        n12159) );
  XNOR2_X1 U11538 ( .A(n13533), .B(n12159), .ZN(n13326) );
  INV_X1 U11539 ( .A(n13533), .ZN(n12304) );
  NAND2_X1 U11540 ( .A1(n12304), .A2(n12159), .ZN(n13212) );
  NAND2_X1 U11541 ( .A1(n9266), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8937) );
  NAND2_X1 U11542 ( .A1(n9321), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8936) );
  OR2_X1 U11543 ( .A1(n8932), .A2(n8931), .ZN(n8933) );
  AND2_X1 U11544 ( .A1(n8952), .A2(n8933), .ZN(n12308) );
  OR2_X1 U11545 ( .A1(n9134), .A2(n12308), .ZN(n8935) );
  INV_X1 U11546 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11884) );
  OR2_X1 U11547 ( .A1(n11521), .A2(n11884), .ZN(n8934) );
  NAND4_X1 U11548 ( .A1(n8937), .A2(n8936), .A3(n8935), .A4(n8934), .ZN(n13531) );
  INV_X1 U11549 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n14040) );
  NOR2_X1 U11550 ( .A1(n8942), .A2(n14040), .ZN(n8939) );
  MUX2_X1 U11551 ( .A(n14040), .B(n8939), .S(P3_IR_REG_9__SCAN_IN), .Z(n8940)
         );
  INV_X1 U11552 ( .A(n8940), .ZN(n8943) );
  INV_X1 U11553 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8941) );
  NAND2_X1 U11554 ( .A1(n8942), .A2(n8941), .ZN(n8977) );
  NAND2_X1 U11555 ( .A1(n8943), .A2(n8977), .ZN(n15670) );
  NAND2_X1 U11556 ( .A1(n10516), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8958) );
  NAND2_X1 U11557 ( .A1(n10518), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8946) );
  OR2_X1 U11558 ( .A1(n8948), .A2(n8947), .ZN(n8949) );
  AND2_X1 U11559 ( .A1(n8959), .A2(n8949), .ZN(n10397) );
  OR2_X1 U11560 ( .A1(n9145), .A2(n10397), .ZN(n8950) );
  NAND2_X1 U11561 ( .A1(n13531), .A2(n12295), .ZN(n13217) );
  NAND2_X1 U11562 ( .A1(n12357), .A2(n9286), .ZN(n13216) );
  NAND2_X1 U11563 ( .A1(n9266), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8957) );
  INV_X1 U11564 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n12395) );
  OR2_X1 U11565 ( .A1(n8860), .A2(n12395), .ZN(n8956) );
  OR2_X2 U11566 ( .A1(n8952), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8970) );
  NAND2_X1 U11567 ( .A1(n8952), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8953) );
  AND2_X1 U11568 ( .A1(n8970), .A2(n8953), .ZN(n12396) );
  OR2_X1 U11569 ( .A1(n9134), .A2(n12396), .ZN(n8955) );
  INV_X1 U11570 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11888) );
  OR2_X1 U11571 ( .A1(n11521), .A2(n11888), .ZN(n8954) );
  NAND2_X1 U11572 ( .A1(n10583), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8960) );
  OR2_X1 U11573 ( .A1(n8962), .A2(n8961), .ZN(n8963) );
  AND2_X1 U11574 ( .A1(n8982), .A2(n8963), .ZN(n10413) );
  OR2_X1 U11575 ( .A1(n9145), .A2(n10413), .ZN(n8968) );
  NAND2_X1 U11576 ( .A1(n8977), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8965) );
  XNOR2_X1 U11577 ( .A(n8965), .B(n8964), .ZN(n12262) );
  INV_X1 U11578 ( .A(n12262), .ZN(n11895) );
  OR2_X1 U11579 ( .A1(n10856), .A2(n11895), .ZN(n8966) );
  INV_X1 U11580 ( .A(n15730), .ZN(n12397) );
  NAND2_X1 U11581 ( .A1(n13530), .A2(n12397), .ZN(n13222) );
  NAND2_X1 U11582 ( .A1(n12390), .A2(n13222), .ZN(n8969) );
  NAND2_X1 U11583 ( .A1(n12526), .A2(n15730), .ZN(n13221) );
  NAND2_X1 U11584 ( .A1(n8969), .A2(n13221), .ZN(n12523) );
  NAND2_X1 U11585 ( .A1(n9266), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8976) );
  INV_X1 U11586 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n12528) );
  OR2_X1 U11587 ( .A1(n8860), .A2(n12528), .ZN(n8975) );
  NAND2_X1 U11588 ( .A1(n8970), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8971) );
  AND2_X1 U11589 ( .A1(n8987), .A2(n8971), .ZN(n12527) );
  OR2_X1 U11590 ( .A1(n9134), .A2(n12527), .ZN(n8974) );
  INV_X1 U11591 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n8972) );
  OR2_X1 U11592 ( .A1(n11521), .A2(n8972), .ZN(n8973) );
  NAND4_X1 U11593 ( .A1(n8976), .A2(n8975), .A3(n8974), .A4(n8973), .ZN(n13529) );
  NAND2_X1 U11594 ( .A1(n8998), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8979) );
  XNOR2_X1 U11595 ( .A(n8979), .B(n8978), .ZN(n12339) );
  INV_X1 U11596 ( .A(n12339), .ZN(n12328) );
  XNOR2_X1 U11597 ( .A(n10682), .B(P2_DATAO_REG_11__SCAN_IN), .ZN(n8983) );
  XNOR2_X1 U11598 ( .A(n8995), .B(n8983), .ZN(n10420) );
  OR2_X1 U11599 ( .A1(n9145), .A2(n10420), .ZN(n8984) );
  OAI211_X1 U11600 ( .C1(n12328), .C2(n10856), .A(n8985), .B(n8984), .ZN(
        n15150) );
  INV_X1 U11601 ( .A(n15150), .ZN(n12530) );
  NAND2_X1 U11602 ( .A1(n13909), .A2(n12530), .ZN(n13227) );
  NAND2_X1 U11603 ( .A1(n13529), .A2(n15150), .ZN(n13226) );
  NAND2_X1 U11604 ( .A1(n12523), .A2(n13327), .ZN(n8986) );
  NAND2_X1 U11605 ( .A1(n8986), .A2(n13227), .ZN(n13912) );
  NAND2_X1 U11606 ( .A1(n9266), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8993) );
  INV_X1 U11607 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n13916) );
  OR2_X1 U11608 ( .A1(n8860), .A2(n13916), .ZN(n8992) );
  AND2_X1 U11609 ( .A1(n8987), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8988) );
  NOR2_X1 U11610 ( .A1(n9014), .A2(n8988), .ZN(n13915) );
  OR2_X1 U11611 ( .A1(n9134), .A2(n13915), .ZN(n8991) );
  INV_X1 U11612 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n8989) );
  OR2_X1 U11613 ( .A1(n11521), .A2(n8989), .ZN(n8990) );
  NAND2_X1 U11614 ( .A1(n10682), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8994) );
  NAND2_X1 U11615 ( .A1(n10684), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8996) );
  XNOR2_X1 U11616 ( .A(n9005), .B(P1_DATAO_REG_12__SCAN_IN), .ZN(n9002) );
  XNOR2_X1 U11617 ( .A(n9004), .B(n9002), .ZN(n10434) );
  NAND2_X1 U11618 ( .A1(n10434), .A2(n13149), .ZN(n9001) );
  OR2_X1 U11619 ( .A1(n9008), .A2(n14040), .ZN(n8999) );
  XNOR2_X1 U11620 ( .A(n8999), .B(P3_IR_REG_12__SCAN_IN), .ZN(n13545) );
  OR2_X1 U11621 ( .A1(n10856), .A2(n13540), .ZN(n9000) );
  OAI211_X1 U11622 ( .C1(n13150), .C2(n10436), .A(n9001), .B(n9000), .ZN(
        n12897) );
  NAND2_X1 U11623 ( .A1(n13897), .A2(n12897), .ZN(n13231) );
  INV_X1 U11624 ( .A(n12897), .ZN(n15146) );
  NAND2_X1 U11625 ( .A1(n13483), .A2(n15146), .ZN(n13232) );
  NAND2_X1 U11626 ( .A1(n13231), .A2(n13232), .ZN(n13906) );
  INV_X1 U11627 ( .A(n13906), .ZN(n13911) );
  INV_X1 U11628 ( .A(n9002), .ZN(n9003) );
  NAND2_X1 U11629 ( .A1(n9005), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n9006) );
  XNOR2_X1 U11630 ( .A(n9021), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n10448) );
  NAND2_X1 U11631 ( .A1(n10448), .A2(n13149), .ZN(n9012) );
  NAND2_X1 U11632 ( .A1(n9008), .A2(n9007), .ZN(n9025) );
  NAND2_X1 U11633 ( .A1(n9025), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9010) );
  XNOR2_X1 U11634 ( .A(n9009), .B(n9010), .ZN(n13560) );
  AOI22_X1 U11635 ( .A1(n9115), .A2(n10449), .B1(n9114), .B2(n13560), .ZN(
        n9011) );
  NAND2_X1 U11636 ( .A1(n9012), .A2(n9011), .ZN(n15142) );
  NAND2_X1 U11637 ( .A1(n9321), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n9020) );
  NAND2_X1 U11638 ( .A1(n9266), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n9019) );
  INV_X1 U11639 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n9013) );
  OR2_X1 U11640 ( .A1(n9014), .A2(n9013), .ZN(n9015) );
  NAND2_X1 U11641 ( .A1(n9014), .A2(n9013), .ZN(n9031) );
  AND2_X1 U11642 ( .A1(n9015), .A2(n9031), .ZN(n13898) );
  OR2_X1 U11643 ( .A1(n9134), .A2(n13898), .ZN(n9018) );
  INV_X1 U11644 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n9016) );
  OR2_X1 U11645 ( .A1(n11521), .A2(n9016), .ZN(n9017) );
  NOR2_X1 U11646 ( .A1(n15142), .A2(n13879), .ZN(n13236) );
  NAND2_X1 U11647 ( .A1(n15142), .A2(n13879), .ZN(n13230) );
  XNOR2_X1 U11648 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n9024) );
  XNOR2_X1 U11649 ( .A(n9042), .B(n9024), .ZN(n10456) );
  NAND2_X1 U11650 ( .A1(n10456), .A2(n13149), .ZN(n9029) );
  NAND2_X1 U11651 ( .A1(n9047), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9027) );
  XNOR2_X1 U11652 ( .A(n9027), .B(n9026), .ZN(n13583) );
  AOI22_X1 U11653 ( .A1(n9115), .A2(n10457), .B1(n9114), .B2(n13583), .ZN(
        n9028) );
  NAND2_X1 U11654 ( .A1(n9321), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n9036) );
  INV_X1 U11655 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n14030) );
  OR2_X1 U11656 ( .A1(n9030), .A2(n14030), .ZN(n9035) );
  NAND2_X1 U11657 ( .A1(n9031), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9032) );
  AND2_X1 U11658 ( .A1(n9051), .A2(n9032), .ZN(n13885) );
  OR2_X1 U11659 ( .A1(n9134), .A2(n13885), .ZN(n9034) );
  INV_X1 U11660 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n13981) );
  OR2_X1 U11661 ( .A1(n11521), .A2(n13981), .ZN(n9033) );
  NAND2_X1 U11662 ( .A1(n14032), .A2(n13896), .ZN(n9037) );
  INV_X1 U11663 ( .A(n13883), .ZN(n9038) );
  OR2_X1 U11664 ( .A1(n14032), .A2(n13528), .ZN(n9039) );
  NAND2_X1 U11665 ( .A1(n9040), .A2(n9039), .ZN(n13866) );
  NAND2_X1 U11666 ( .A1(n11046), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n9041) );
  NAND2_X1 U11667 ( .A1(n11081), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n9058) );
  NAND2_X1 U11668 ( .A1(n11079), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n9043) );
  NAND2_X1 U11669 ( .A1(n9058), .A2(n9043), .ZN(n9044) );
  NAND2_X1 U11670 ( .A1(n9045), .A2(n9044), .ZN(n9046) );
  NAND2_X1 U11671 ( .A1(n9059), .A2(n9046), .ZN(n10496) );
  OR2_X1 U11672 ( .A1(n10496), .A2(n9145), .ZN(n9050) );
  OAI21_X1 U11673 ( .B1(n9047), .B2(P3_IR_REG_14__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9048) );
  XNOR2_X1 U11674 ( .A(n9048), .B(P3_IR_REG_15__SCAN_IN), .ZN(n13610) );
  AOI22_X1 U11675 ( .A1(n9115), .A2(SI_15_), .B1(n9114), .B2(n13610), .ZN(
        n9049) );
  NAND2_X1 U11676 ( .A1(n9266), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n9056) );
  INV_X1 U11677 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13977) );
  OR2_X1 U11678 ( .A1(n11521), .A2(n13977), .ZN(n9055) );
  AND2_X1 U11679 ( .A1(n9051), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9052) );
  NOR2_X1 U11680 ( .A1(n9067), .A2(n9052), .ZN(n13867) );
  OR2_X1 U11681 ( .A1(n9134), .A2(n13867), .ZN(n9054) );
  INV_X1 U11682 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n13585) );
  OR2_X1 U11683 ( .A1(n8860), .A2(n13585), .ZN(n9053) );
  OR2_X1 U11684 ( .A1(n13521), .A2(n13510), .ZN(n13240) );
  NAND2_X1 U11685 ( .A1(n13521), .A2(n13510), .ZN(n13250) );
  NAND2_X1 U11686 ( .A1(n13866), .A2(n13865), .ZN(n9057) );
  NAND2_X1 U11687 ( .A1(n9057), .A2(n13250), .ZN(n13858) );
  NAND2_X1 U11688 ( .A1(n11025), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n9073) );
  NAND2_X1 U11689 ( .A1(n11023), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n9060) );
  OR2_X1 U11690 ( .A1(n9062), .A2(n9061), .ZN(n9063) );
  NAND2_X1 U11691 ( .A1(n9074), .A2(n9063), .ZN(n10571) );
  OR2_X1 U11692 ( .A1(n10571), .A2(n9145), .ZN(n9066) );
  NAND2_X1 U11693 ( .A1(n6808), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9064) );
  XNOR2_X1 U11694 ( .A(n9064), .B(P3_IR_REG_16__SCAN_IN), .ZN(n13640) );
  AOI22_X1 U11695 ( .A1(n9115), .A2(SI_16_), .B1(n9114), .B2(n13640), .ZN(
        n9065) );
  NAND2_X1 U11696 ( .A1(n9266), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n9072) );
  INV_X1 U11697 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13854) );
  OR2_X1 U11698 ( .A1(n8860), .A2(n13854), .ZN(n9071) );
  NOR2_X1 U11699 ( .A1(n9067), .A2(n13441), .ZN(n9068) );
  OR2_X1 U11700 ( .A1(n9134), .A2(n6707), .ZN(n9070) );
  INV_X1 U11701 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13639) );
  OR2_X1 U11702 ( .A1(n11521), .A2(n13639), .ZN(n9069) );
  OR2_X1 U11703 ( .A1(n13971), .A2(n13864), .ZN(n13252) );
  NAND2_X1 U11704 ( .A1(n13971), .A2(n13864), .ZN(n13251) );
  NAND2_X1 U11705 ( .A1(n13252), .A2(n13251), .ZN(n13838) );
  NAND2_X1 U11706 ( .A1(n11064), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n9091) );
  INV_X1 U11707 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11067) );
  NAND2_X1 U11708 ( .A1(n11067), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n9075) );
  NAND2_X1 U11709 ( .A1(n9091), .A2(n9075), .ZN(n9088) );
  XNOR2_X1 U11710 ( .A(n9090), .B(n9088), .ZN(n10688) );
  NAND2_X1 U11711 ( .A1(n10688), .A2(n13149), .ZN(n9080) );
  NAND2_X1 U11712 ( .A1(n9076), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9077) );
  MUX2_X1 U11713 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9077), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n9078) );
  NAND2_X1 U11714 ( .A1(n9078), .A2(n8783), .ZN(n13649) );
  INV_X1 U11715 ( .A(n13649), .ZN(n15130) );
  AOI22_X1 U11716 ( .A1(n9115), .A2(SI_17_), .B1(n9114), .B2(n15130), .ZN(
        n9079) );
  NAND2_X1 U11717 ( .A1(n9266), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n9087) );
  INV_X1 U11718 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n15127) );
  OR2_X1 U11719 ( .A1(n8860), .A2(n15127), .ZN(n9086) );
  OR2_X1 U11720 ( .A1(n9081), .A2(n9635), .ZN(n9082) );
  AND2_X1 U11721 ( .A1(n9100), .A2(n9082), .ZN(n13845) );
  OR2_X1 U11722 ( .A1(n9134), .A2(n13845), .ZN(n9085) );
  INV_X1 U11723 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n9083) );
  OR2_X1 U11724 ( .A1(n11521), .A2(n9083), .ZN(n9084) );
  OR2_X1 U11725 ( .A1(n13967), .A2(n13828), .ZN(n13258) );
  NAND2_X1 U11726 ( .A1(n13967), .A2(n13828), .ZN(n13255) );
  NAND2_X1 U11727 ( .A1(n13258), .A2(n13255), .ZN(n13332) );
  INV_X1 U11728 ( .A(n13832), .ZN(n9107) );
  INV_X1 U11729 ( .A(n9088), .ZN(n9089) );
  NAND2_X1 U11730 ( .A1(n11389), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n9108) );
  NAND2_X1 U11731 ( .A1(n11391), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n9093) );
  OR2_X1 U11732 ( .A1(n9095), .A2(n9094), .ZN(n9096) );
  NAND2_X1 U11733 ( .A1(n9109), .A2(n9096), .ZN(n10738) );
  OR2_X1 U11734 ( .A1(n10738), .A2(n9145), .ZN(n9099) );
  NAND2_X1 U11735 ( .A1(n8783), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9097) );
  XNOR2_X1 U11736 ( .A(n9097), .B(P3_IR_REG_18__SCAN_IN), .ZN(n13664) );
  AOI22_X1 U11737 ( .A1(n9115), .A2(SI_18_), .B1(n9114), .B2(n13664), .ZN(
        n9098) );
  NAND2_X1 U11738 ( .A1(n9321), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n9105) );
  NAND2_X1 U11739 ( .A1(n9266), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n9104) );
  NAND2_X1 U11740 ( .A1(n9189), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n9103) );
  NAND2_X1 U11741 ( .A1(n9100), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9101) );
  AND2_X1 U11742 ( .A1(n9118), .A2(n9101), .ZN(n13829) );
  OR2_X1 U11743 ( .A1(n9134), .A2(n13829), .ZN(n9102) );
  NAND2_X1 U11744 ( .A1(n13960), .A2(n13449), .ZN(n13262) );
  NAND2_X1 U11745 ( .A1(n13256), .A2(n13262), .ZN(n13831) );
  INV_X1 U11746 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11597) );
  NAND2_X1 U11747 ( .A1(n11597), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n9125) );
  INV_X1 U11748 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n12958) );
  NAND2_X1 U11749 ( .A1(n12958), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n9110) );
  OR2_X1 U11750 ( .A1(n9112), .A2(n9111), .ZN(n9113) );
  NAND2_X1 U11751 ( .A1(n9126), .A2(n9113), .ZN(n10785) );
  OR2_X1 U11752 ( .A1(n10785), .A2(n9145), .ZN(n9117) );
  AOI22_X1 U11753 ( .A1(n9115), .A2(SI_19_), .B1(n9114), .B2(n13666), .ZN(
        n9116) );
  NAND2_X1 U11754 ( .A1(n9266), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n9123) );
  AND2_X1 U11755 ( .A1(n9118), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9119) );
  NOR2_X1 U11756 ( .A1(n9132), .A2(n9119), .ZN(n13818) );
  OR2_X1 U11757 ( .A1(n13818), .A2(n9134), .ZN(n9122) );
  INV_X1 U11758 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13958) );
  OR2_X1 U11759 ( .A1(n11521), .A2(n13958), .ZN(n9121) );
  INV_X1 U11760 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13819) );
  OR2_X1 U11761 ( .A1(n8860), .A2(n13819), .ZN(n9120) );
  INV_X1 U11762 ( .A(n13268), .ZN(n9124) );
  NAND2_X1 U11763 ( .A1(n13817), .A2(n13827), .ZN(n13269) );
  NAND2_X1 U11764 ( .A1(n9128), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9129) );
  NAND2_X1 U11765 ( .A1(n9140), .A2(n9129), .ZN(n11027) );
  INV_X1 U11766 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n13471) );
  NOR2_X1 U11767 ( .A1(n9132), .A2(n13471), .ZN(n9133) );
  OR2_X1 U11768 ( .A1(n9151), .A2(n9133), .ZN(n13805) );
  NAND2_X1 U11769 ( .A1(n13805), .A2(n9265), .ZN(n9138) );
  NAND2_X1 U11770 ( .A1(n9321), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n9137) );
  NAND2_X1 U11771 ( .A1(n9266), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n9136) );
  INV_X1 U11772 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13954) );
  OR2_X1 U11773 ( .A1(n11521), .A2(n13954), .ZN(n9135) );
  NAND2_X1 U11774 ( .A1(n13804), .A2(n13789), .ZN(n13273) );
  NAND2_X1 U11775 ( .A1(n11816), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9156) );
  NAND2_X1 U11776 ( .A1(n11814), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9141) );
  AND2_X1 U11777 ( .A1(n9156), .A2(n9141), .ZN(n9142) );
  OR2_X1 U11778 ( .A1(n9143), .A2(n9142), .ZN(n9144) );
  NAND2_X1 U11779 ( .A1(n9157), .A2(n9144), .ZN(n11100) );
  INV_X1 U11780 ( .A(SI_21_), .ZN(n11099) );
  NAND2_X1 U11781 ( .A1(n9266), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n9149) );
  NAND2_X1 U11782 ( .A1(n9321), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n9148) );
  AND2_X1 U11783 ( .A1(n9149), .A2(n9148), .ZN(n9155) );
  INV_X1 U11784 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n9150) );
  OR2_X1 U11785 ( .A1(n9151), .A2(n9150), .ZN(n9152) );
  NAND2_X1 U11786 ( .A1(n9186), .A2(n9152), .ZN(n13790) );
  NAND2_X1 U11787 ( .A1(n13790), .A2(n9265), .ZN(n9154) );
  NAND2_X1 U11788 ( .A1(n9189), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n9153) );
  NAND2_X1 U11789 ( .A1(n13414), .A2(n13801), .ZN(n13736) );
  XNOR2_X1 U11790 ( .A(n12000), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n9181) );
  NAND2_X1 U11791 ( .A1(n12000), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n9158) );
  OAI21_X2 U11792 ( .B1(n9182), .B2(n9181), .A(n9158), .ZN(n9173) );
  XNOR2_X1 U11793 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n9172) );
  NAND2_X1 U11794 ( .A1(n12061), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9159) );
  NAND2_X1 U11795 ( .A1(n9160), .A2(n12122), .ZN(n9161) );
  INV_X1 U11796 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n12125) );
  XNOR2_X1 U11797 ( .A(n9203), .B(n12125), .ZN(n11936) );
  NAND2_X1 U11798 ( .A1(n11936), .A2(n13149), .ZN(n9163) );
  INV_X1 U11799 ( .A(SI_24_), .ZN(n11937) );
  NAND2_X2 U11800 ( .A1(n9163), .A2(n9162), .ZN(n13937) );
  OR2_X2 U11801 ( .A1(n9188), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9177) );
  INV_X1 U11802 ( .A(n9208), .ZN(n9165) );
  NAND2_X1 U11803 ( .A1(n9177), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9164) );
  NAND2_X1 U11804 ( .A1(n9165), .A2(n9164), .ZN(n13751) );
  NAND2_X1 U11805 ( .A1(n13751), .A2(n9265), .ZN(n9171) );
  INV_X1 U11806 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n9168) );
  NAND2_X1 U11807 ( .A1(n9266), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n9167) );
  NAND2_X1 U11808 ( .A1(n9321), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n9166) );
  OAI211_X1 U11809 ( .C1(n11521), .C2(n9168), .A(n9167), .B(n9166), .ZN(n9169)
         );
  INV_X1 U11810 ( .A(n9169), .ZN(n9170) );
  AND2_X2 U11811 ( .A1(n9171), .A2(n9170), .ZN(n13723) );
  NAND2_X1 U11812 ( .A1(n13937), .A2(n13723), .ZN(n13281) );
  XNOR2_X2 U11813 ( .A(n13937), .B(n13723), .ZN(n13746) );
  XNOR2_X1 U11814 ( .A(n9173), .B(n9172), .ZN(n11406) );
  NAND2_X1 U11815 ( .A1(n11406), .A2(n13149), .ZN(n9175) );
  INV_X1 U11816 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13942) );
  NAND2_X1 U11817 ( .A1(n9188), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9176) );
  NAND2_X1 U11818 ( .A1(n9177), .A2(n9176), .ZN(n13767) );
  NAND2_X1 U11819 ( .A1(n13767), .A2(n9265), .ZN(n9179) );
  AOI22_X1 U11820 ( .A1(n9266), .A2(P3_REG0_REG_23__SCAN_IN), .B1(n9321), .B2(
        P3_REG2_REG_23__SCAN_IN), .ZN(n9178) );
  INV_X1 U11821 ( .A(n13747), .ZN(n13776) );
  OR2_X1 U11822 ( .A1(n13766), .A2(n13776), .ZN(n13283) );
  INV_X1 U11823 ( .A(n13283), .ZN(n9180) );
  XNOR2_X1 U11824 ( .A(n9182), .B(n9181), .ZN(n11254) );
  NAND2_X1 U11825 ( .A1(n11254), .A2(n13149), .ZN(n9185) );
  NAND2_X1 U11826 ( .A1(n9186), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9187) );
  NAND2_X1 U11827 ( .A1(n9188), .A2(n9187), .ZN(n13777) );
  NAND2_X1 U11828 ( .A1(n13777), .A2(n9265), .ZN(n9192) );
  AOI22_X1 U11829 ( .A1(n9266), .A2(P3_REG0_REG_22__SCAN_IN), .B1(n9321), .B2(
        P3_REG2_REG_22__SCAN_IN), .ZN(n9191) );
  NAND2_X1 U11830 ( .A1(n9189), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n9190) );
  AND2_X1 U11831 ( .A1(n13757), .A2(n13283), .ZN(n13740) );
  INV_X1 U11832 ( .A(n9198), .ZN(n9196) );
  NAND2_X1 U11833 ( .A1(n12931), .A2(n13788), .ZN(n13739) );
  AND2_X1 U11834 ( .A1(n13739), .A2(n9193), .ZN(n9194) );
  AND2_X1 U11835 ( .A1(n9194), .A2(n13281), .ZN(n9195) );
  OR2_X2 U11836 ( .A1(n9196), .A2(n9195), .ZN(n9197) );
  AND2_X1 U11837 ( .A1(n13736), .A2(n9197), .ZN(n9201) );
  INV_X1 U11838 ( .A(n9197), .ZN(n9200) );
  AND2_X1 U11839 ( .A1(n13737), .A2(n9198), .ZN(n9199) );
  OAI21_X1 U11840 ( .B1(n9203), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n9202), .ZN(
        n9216) );
  XNOR2_X1 U11841 ( .A(n12167), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n9204) );
  XNOR2_X1 U11842 ( .A(n9216), .B(n9204), .ZN(n12036) );
  NAND2_X1 U11843 ( .A1(n12036), .A2(n13149), .ZN(n9206) );
  INV_X1 U11844 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n9207) );
  NAND2_X1 U11845 ( .A1(n9208), .A2(n9207), .ZN(n9221) );
  OR2_X1 U11846 ( .A1(n9208), .A2(n9207), .ZN(n9209) );
  NAND2_X1 U11847 ( .A1(n9221), .A2(n9209), .ZN(n13730) );
  INV_X1 U11848 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13934) );
  NAND2_X1 U11849 ( .A1(n9321), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n9211) );
  NAND2_X1 U11850 ( .A1(n9266), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n9210) );
  OAI211_X1 U11851 ( .C1(n13934), .C2(n11521), .A(n9211), .B(n9210), .ZN(n9212) );
  NAND2_X1 U11852 ( .A1(n13427), .A2(n13750), .ZN(n9213) );
  INV_X1 U11853 ( .A(n13721), .ZN(n9214) );
  INV_X1 U11854 ( .A(n9213), .ZN(n13287) );
  NAND2_X1 U11855 ( .A1(n12167), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9215) );
  NAND2_X1 U11856 ( .A1(n12574), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9217) );
  XNOR2_X1 U11857 ( .A(n12385), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n9218) );
  XNOR2_X1 U11858 ( .A(n9229), .B(n9218), .ZN(n12148) );
  NAND2_X1 U11859 ( .A1(n12148), .A2(n13149), .ZN(n9220) );
  NAND2_X1 U11860 ( .A1(n9221), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9222) );
  NAND2_X1 U11861 ( .A1(n9234), .A2(n9222), .ZN(n13713) );
  NAND2_X1 U11862 ( .A1(n13713), .A2(n9265), .ZN(n9227) );
  INV_X1 U11863 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n10156) );
  NAND2_X1 U11864 ( .A1(n9266), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n9224) );
  NAND2_X1 U11865 ( .A1(n9321), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n9223) );
  OAI211_X1 U11866 ( .C1(n11521), .C2(n10156), .A(n9224), .B(n9223), .ZN(n9225) );
  INV_X1 U11867 ( .A(n9225), .ZN(n9226) );
  NAND2_X1 U11868 ( .A1(n9306), .A2(n13724), .ZN(n10148) );
  AND2_X1 U11869 ( .A1(n12389), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9228) );
  NAND2_X1 U11870 ( .A1(n12385), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9230) );
  XNOR2_X1 U11871 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n9231) );
  XNOR2_X1 U11872 ( .A(n9244), .B(n9231), .ZN(n12309) );
  NAND2_X1 U11873 ( .A1(n12309), .A2(n13149), .ZN(n9233) );
  INV_X1 U11874 ( .A(SI_27_), .ZN(n12310) );
  INV_X1 U11875 ( .A(n9250), .ZN(n9236) );
  NAND2_X1 U11876 ( .A1(n9234), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9235) );
  NAND2_X1 U11877 ( .A1(n9236), .A2(n9235), .ZN(n13127) );
  NAND2_X1 U11878 ( .A1(n13127), .A2(n9265), .ZN(n9242) );
  INV_X1 U11879 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n9239) );
  NAND2_X1 U11880 ( .A1(n9266), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n9238) );
  NAND2_X1 U11881 ( .A1(n9321), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n9237) );
  OAI211_X1 U11882 ( .C1(n9239), .C2(n11521), .A(n9238), .B(n9237), .ZN(n9240)
         );
  INV_X1 U11883 ( .A(n9240), .ZN(n9241) );
  NAND2_X2 U11884 ( .A1(n9242), .A2(n9241), .ZN(n13299) );
  AND2_X1 U11885 ( .A1(n12479), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9243) );
  NAND2_X1 U11886 ( .A1(n12475), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9245) );
  XNOR2_X1 U11887 ( .A(n9260), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n9247) );
  XNOR2_X1 U11888 ( .A(n9257), .B(n9247), .ZN(n12848) );
  NAND2_X1 U11889 ( .A1(n12848), .A2(n13149), .ZN(n9249) );
  INV_X1 U11890 ( .A(SI_28_), .ZN(n12851) );
  OR2_X1 U11891 ( .A1(n13150), .A2(n12851), .ZN(n9248) );
  INV_X1 U11892 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n13367) );
  NOR2_X1 U11893 ( .A1(n9250), .A2(n13367), .ZN(n9251) );
  INV_X1 U11894 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n9254) );
  NAND2_X1 U11895 ( .A1(n9266), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n9253) );
  NAND2_X1 U11896 ( .A1(n9321), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n9252) );
  OAI211_X1 U11897 ( .C1(n9254), .C2(n11521), .A(n9253), .B(n9252), .ZN(n9255)
         );
  NAND2_X1 U11898 ( .A1(n13707), .A2(n10177), .ZN(n9315) );
  INV_X1 U11899 ( .A(n9315), .ZN(n9256) );
  NOR2_X1 U11900 ( .A1(n13300), .A2(n13299), .ZN(n13697) );
  NOR2_X1 U11901 ( .A1(n9256), .A2(n13697), .ZN(n13304) );
  INV_X1 U11902 ( .A(n9316), .ZN(n13303) );
  INV_X1 U11903 ( .A(n9257), .ZN(n9259) );
  INV_X1 U11904 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12995) );
  NAND2_X1 U11905 ( .A1(n12995), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9258) );
  NAND2_X1 U11906 ( .A1(n9259), .A2(n9258), .ZN(n9262) );
  NAND2_X1 U11907 ( .A1(n9260), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9261) );
  XNOR2_X1 U11908 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n13134) );
  XNOR2_X1 U11909 ( .A(n13136), .B(n13134), .ZN(n14045) );
  NAND2_X1 U11910 ( .A1(n14045), .A2(n13149), .ZN(n9264) );
  INV_X1 U11911 ( .A(SI_29_), .ZN(n14048) );
  OR2_X1 U11912 ( .A1(n13150), .A2(n14048), .ZN(n9263) );
  NAND2_X1 U11913 ( .A1(n9264), .A2(n9263), .ZN(n9370) );
  NAND2_X1 U11914 ( .A1(n13690), .A2(n9265), .ZN(n11525) );
  INV_X1 U11915 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9269) );
  NAND2_X1 U11916 ( .A1(n9266), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9268) );
  NAND2_X1 U11917 ( .A1(n9321), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n9267) );
  OAI211_X1 U11918 ( .C1(n11521), .C2(n9269), .A(n9268), .B(n9267), .ZN(n9270)
         );
  INV_X1 U11919 ( .A(n9270), .ZN(n9271) );
  NAND2_X1 U11920 ( .A1(n9370), .A2(n13702), .ZN(n13306) );
  INV_X1 U11921 ( .A(n13338), .ZN(n9272) );
  XNOR2_X1 U11922 ( .A(n13133), .B(n9272), .ZN(n13689) );
  INV_X1 U11923 ( .A(n12159), .ZN(n13210) );
  NAND2_X1 U11924 ( .A1(n15691), .A2(n11173), .ZN(n15684) );
  INV_X1 U11925 ( .A(n15697), .ZN(n11178) );
  AND2_X1 U11926 ( .A1(n15684), .A2(n9276), .ZN(n9275) );
  NAND2_X1 U11927 ( .A1(n13536), .A2(n9274), .ZN(n11673) );
  NAND2_X1 U11928 ( .A1(n11169), .A2(n11673), .ZN(n15683) );
  NAND2_X1 U11929 ( .A1(n9275), .A2(n15683), .ZN(n11492) );
  NAND2_X1 U11930 ( .A1(n15687), .A2(n9276), .ZN(n11493) );
  NAND2_X1 U11931 ( .A1(n6679), .A2(n11287), .ZN(n9278) );
  NAND2_X1 U11932 ( .A1(n11492), .A2(n9277), .ZN(n11394) );
  INV_X1 U11933 ( .A(n11397), .ZN(n9280) );
  NAND2_X1 U11934 ( .A1(n9278), .A2(n13319), .ZN(n11395) );
  INV_X1 U11935 ( .A(n11395), .ZN(n9279) );
  NOR2_X1 U11936 ( .A1(n9280), .A2(n9279), .ZN(n9281) );
  NAND2_X1 U11937 ( .A1(n8859), .A2(n11578), .ZN(n9283) );
  NAND2_X1 U11938 ( .A1(n12007), .A2(n11795), .ZN(n9284) );
  NAND2_X1 U11939 ( .A1(n11958), .A2(n13534), .ZN(n9285) );
  NAND2_X1 U11940 ( .A1(n12004), .A2(n9285), .ZN(n11825) );
  NAND2_X1 U11941 ( .A1(n11825), .A2(n12023), .ZN(n11824) );
  XNOR2_X1 U11942 ( .A(n13531), .B(n12295), .ZN(n13323) );
  NAND2_X1 U11943 ( .A1(n13531), .A2(n9286), .ZN(n9287) );
  NAND2_X1 U11944 ( .A1(n13221), .A2(n13222), .ZN(n13220) );
  NAND2_X1 U11945 ( .A1(n13876), .A2(n13883), .ZN(n13875) );
  NAND2_X1 U11946 ( .A1(n13875), .A2(n9289), .ZN(n13862) );
  NAND2_X1 U11947 ( .A1(n13967), .A2(n13852), .ZN(n9293) );
  INV_X1 U11948 ( .A(n9293), .ZN(n9290) );
  AND2_X1 U11949 ( .A1(n13838), .A2(n9292), .ZN(n9291) );
  NAND2_X1 U11950 ( .A1(n13851), .A2(n9291), .ZN(n9297) );
  INV_X1 U11951 ( .A(n9292), .ZN(n9295) );
  NAND2_X1 U11952 ( .A1(n13971), .A2(n13843), .ZN(n13839) );
  AND2_X1 U11953 ( .A1(n13839), .A2(n9293), .ZN(n9294) );
  NAND2_X1 U11954 ( .A1(n9297), .A2(n9296), .ZN(n13795) );
  NAND2_X1 U11955 ( .A1(n13817), .A2(n12923), .ZN(n13797) );
  NAND2_X1 U11956 ( .A1(n13797), .A2(n13831), .ZN(n9299) );
  NOR2_X1 U11957 ( .A1(n13960), .A2(n13842), .ZN(n13796) );
  OAI21_X1 U11958 ( .B1(n13315), .B2(n13796), .A(n13797), .ZN(n9298) );
  INV_X1 U11959 ( .A(n13414), .ZN(n14010) );
  NAND2_X1 U11960 ( .A1(n14010), .A2(n13801), .ZN(n9300) );
  NAND2_X1 U11961 ( .A1(n13783), .A2(n9300), .ZN(n13774) );
  NAND2_X1 U11962 ( .A1(n14006), .A2(n13788), .ZN(n9303) );
  NAND2_X1 U11963 ( .A1(n13766), .A2(n6684), .ZN(n10149) );
  INV_X1 U11964 ( .A(n13299), .ZN(n13703) );
  NAND2_X1 U11965 ( .A1(n13300), .A2(n13703), .ZN(n9314) );
  INV_X1 U11966 ( .A(n9314), .ZN(n9311) );
  NAND2_X1 U11967 ( .A1(n13715), .A2(n13724), .ZN(n9310) );
  INV_X1 U11968 ( .A(n9310), .ZN(n9309) );
  INV_X1 U11969 ( .A(n13750), .ZN(n13527) );
  NAND2_X1 U11970 ( .A1(n13427), .A2(n13527), .ZN(n10151) );
  NAND2_X1 U11971 ( .A1(n9306), .A2(n13526), .ZN(n9307) );
  AND2_X1 U11972 ( .A1(n10151), .A2(n9307), .ZN(n9308) );
  AND2_X1 U11973 ( .A1(n13721), .A2(n9310), .ZN(n10165) );
  NAND2_X1 U11974 ( .A1(n13937), .A2(n13763), .ZN(n10150) );
  AND2_X1 U11975 ( .A1(n9313), .A2(n13746), .ZN(n10169) );
  INV_X1 U11976 ( .A(n13700), .ZN(n9317) );
  INV_X1 U11977 ( .A(n10177), .ZN(n13525) );
  NAND2_X1 U11978 ( .A1(n13707), .A2(n13525), .ZN(n9319) );
  NAND2_X1 U11979 ( .A1(n13705), .A2(n9319), .ZN(n9320) );
  XNOR2_X1 U11980 ( .A(n9320), .B(n13338), .ZN(n9331) );
  NAND2_X1 U11981 ( .A1(n13356), .A2(n13666), .ZN(n9375) );
  NAND2_X1 U11982 ( .A1(n13173), .A2(n9374), .ZN(n13166) );
  INV_X1 U11983 ( .A(n13354), .ZN(n9328) );
  INV_X1 U11984 ( .A(n13667), .ZN(n13590) );
  NAND2_X1 U11985 ( .A1(n9328), .A2(n13590), .ZN(n10864) );
  NAND2_X1 U11986 ( .A1(n10856), .A2(n10864), .ZN(n9327) );
  NAND2_X4 U11987 ( .A1(n13356), .A2(n13173), .ZN(n13267) );
  INV_X1 U11988 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n9324) );
  NAND2_X1 U11989 ( .A1(n9321), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n9323) );
  NAND2_X1 U11990 ( .A1(n9266), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9322) );
  OAI211_X1 U11991 ( .C1(n9324), .C2(n11521), .A(n9323), .B(n9322), .ZN(n9325)
         );
  INV_X1 U11992 ( .A(n9325), .ZN(n9326) );
  AND2_X1 U11993 ( .A1(n11525), .A2(n9326), .ZN(n13153) );
  INV_X4 U11994 ( .A(n13267), .ZN(n13305) );
  AND2_X1 U11995 ( .A1(n9328), .A2(P3_B_REG_SCAN_IN), .ZN(n9329) );
  OR2_X1 U11996 ( .A1(n15689), .A2(n9329), .ZN(n13683) );
  OAI22_X1 U11997 ( .A1(n10177), .A2(n15690), .B1(n13153), .B2(n13683), .ZN(
        n9330) );
  INV_X1 U11998 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9333) );
  NAND2_X1 U11999 ( .A1(n6672), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9336) );
  MUX2_X1 U12000 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9336), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n9339) );
  INV_X1 U12001 ( .A(n11939), .ZN(n9342) );
  NAND2_X1 U12002 ( .A1(n9338), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9340) );
  MUX2_X1 U12003 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9340), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n9341) );
  AND2_X1 U12004 ( .A1(n9341), .A2(n6708), .ZN(n9343) );
  NAND3_X1 U12005 ( .A1(n9346), .A2(n9342), .A3(n9343), .ZN(n11103) );
  XNOR2_X1 U12006 ( .A(n11939), .B(P3_B_REG_SCAN_IN), .ZN(n9344) );
  INV_X1 U12007 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n9345) );
  INV_X1 U12008 ( .A(n9346), .ZN(n12149) );
  NAND2_X1 U12009 ( .A1(n12149), .A2(n11939), .ZN(n9347) );
  INV_X1 U12010 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n9349) );
  NAND2_X1 U12011 ( .A1(n9348), .A2(n9349), .ZN(n9351) );
  NAND2_X1 U12012 ( .A1(n12149), .A2(n12037), .ZN(n9350) );
  NAND2_X1 U12013 ( .A1(n14036), .A2(n14034), .ZN(n9372) );
  NOR2_X1 U12014 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .ZN(
        n9355) );
  NOR4_X1 U12015 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n9354) );
  NOR4_X1 U12016 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n9353) );
  NOR4_X1 U12017 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n9352) );
  NAND4_X1 U12018 ( .A1(n9355), .A2(n9354), .A3(n9353), .A4(n9352), .ZN(n9361)
         );
  NOR4_X1 U12019 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n9359) );
  NOR4_X1 U12020 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n9358) );
  NOR4_X1 U12021 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n9357) );
  NOR4_X1 U12022 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n9356) );
  NAND4_X1 U12023 ( .A1(n9359), .A2(n9358), .A3(n9357), .A4(n9356), .ZN(n9360)
         );
  OAI21_X1 U12024 ( .B1(n9361), .B2(n9360), .A(n9348), .ZN(n9376) );
  INV_X1 U12025 ( .A(n14036), .ZN(n9362) );
  NAND2_X1 U12026 ( .A1(n9362), .A2(n11359), .ZN(n9378) );
  OAI22_X1 U12027 ( .A1(n15719), .A2(n9374), .B1(n13666), .B2(n11252), .ZN(
        n9363) );
  NAND2_X1 U12028 ( .A1(n9363), .A2(n11163), .ZN(n9364) );
  NAND2_X1 U12029 ( .A1(n9364), .A2(n13267), .ZN(n9365) );
  NAND2_X1 U12030 ( .A1(n9365), .A2(n11359), .ZN(n9368) );
  OR2_X1 U12031 ( .A1(n13267), .A2(n13347), .ZN(n11101) );
  NAND2_X1 U12032 ( .A1(n13267), .A2(n9366), .ZN(n11360) );
  NAND2_X1 U12033 ( .A1(n11101), .A2(n11360), .ZN(n11358) );
  NAND2_X1 U12034 ( .A1(n11358), .A2(n14034), .ZN(n9367) );
  INV_X1 U12035 ( .A(n9370), .ZN(n13692) );
  NAND2_X1 U12036 ( .A1(n9371), .A2(n7582), .ZN(P3_U3488) );
  INV_X1 U12037 ( .A(n9372), .ZN(n9373) );
  NAND2_X1 U12038 ( .A1(n9373), .A2(n9376), .ZN(n11120) );
  OR2_X1 U12039 ( .A1(n13267), .A2(n11163), .ZN(n11084) );
  NAND2_X1 U12040 ( .A1(n11160), .A2(n9374), .ZN(n13345) );
  OR2_X1 U12041 ( .A1(n9375), .A2(n13345), .ZN(n11110) );
  INV_X1 U12042 ( .A(n9376), .ZN(n9377) );
  NAND2_X1 U12043 ( .A1(n11115), .A2(n11109), .ZN(n9379) );
  OAI21_X1 U12044 ( .B1(n11120), .B2(n9380), .A(n9379), .ZN(n9381) );
  NAND2_X1 U12045 ( .A1(n9382), .A2(n7585), .ZN(P3_U3456) );
  INV_X1 U12046 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n9474) );
  INV_X1 U12047 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15272) );
  INV_X1 U12048 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n9469) );
  NAND2_X1 U12049 ( .A1(n9469), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n9468) );
  INV_X1 U12050 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n9411) );
  XOR2_X1 U12051 ( .A(n9411), .B(P1_ADDR_REG_14__SCAN_IN), .Z(n9413) );
  INV_X1 U12052 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9460) );
  INV_X1 U12053 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n9407) );
  XOR2_X1 U12054 ( .A(P1_ADDR_REG_12__SCAN_IN), .B(n9407), .Z(n9459) );
  INV_X1 U12055 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n9405) );
  XOR2_X1 U12056 ( .A(n9806), .B(P1_ADDR_REG_9__SCAN_IN), .Z(n9448) );
  XOR2_X1 U12057 ( .A(n9809), .B(P1_ADDR_REG_8__SCAN_IN), .Z(n9441) );
  INV_X1 U12058 ( .A(n9422), .ZN(n9421) );
  NOR2_X1 U12059 ( .A1(n9385), .A2(n9796), .ZN(n9387) );
  NOR2_X1 U12060 ( .A1(n9388), .A2(n9389), .ZN(n9391) );
  INV_X1 U12061 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n9393) );
  NOR2_X1 U12062 ( .A1(n9392), .A2(n9393), .ZN(n9395) );
  NOR2_X2 U12063 ( .A1(n9395), .A2(n9394), .ZN(n9435) );
  AND2_X1 U12064 ( .A1(n9716), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9396) );
  NAND2_X1 U12065 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n9397), .ZN(n9398) );
  INV_X1 U12066 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n9592) );
  NAND2_X1 U12067 ( .A1(n9441), .A2(n9442), .ZN(n9399) );
  NAND2_X1 U12068 ( .A1(n9448), .A2(n9447), .ZN(n9400) );
  INV_X1 U12069 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9402) );
  NOR2_X1 U12070 ( .A1(n9401), .A2(n9402), .ZN(n9403) );
  INV_X1 U12071 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n9415) );
  XOR2_X1 U12072 ( .A(P1_ADDR_REG_11__SCAN_IN), .B(n9405), .Z(n9453) );
  NAND2_X1 U12073 ( .A1(n9454), .A2(n9453), .ZN(n9404) );
  NAND2_X1 U12074 ( .A1(n9459), .A2(n9458), .ZN(n9406) );
  INV_X1 U12075 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n9408) );
  NAND2_X1 U12076 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n9408), .ZN(n9409) );
  AOI21_X2 U12077 ( .B1(n9411), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n9410), .ZN(
        n9470) );
  INV_X1 U12078 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n9467) );
  XOR2_X1 U12079 ( .A(n9413), .B(n9412), .Z(n15244) );
  INV_X1 U12080 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n15436) );
  XOR2_X1 U12081 ( .A(n9415), .B(n9414), .Z(n15114) );
  INV_X1 U12082 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n15372) );
  OR2_X1 U12083 ( .A1(n15372), .A2(n9417), .ZN(n9431) );
  INV_X1 U12084 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15359) );
  INV_X1 U12085 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n9427) );
  XNOR2_X1 U12086 ( .A(n9419), .B(n9418), .ZN(n15103) );
  XNOR2_X1 U12087 ( .A(n9421), .B(n9420), .ZN(n9423) );
  NAND2_X1 U12088 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n9423), .ZN(n9425) );
  AOI21_X1 U12089 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n11219), .A(n9422), .ZN(
        n15747) );
  INV_X1 U12090 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15746) );
  NOR2_X1 U12091 ( .A1(n15747), .A2(n15746), .ZN(n15755) );
  XOR2_X1 U12092 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n9423), .Z(n15754) );
  NAND2_X1 U12093 ( .A1(n15755), .A2(n15754), .ZN(n9424) );
  NAND2_X1 U12094 ( .A1(n9425), .A2(n9424), .ZN(n15104) );
  NAND2_X1 U12095 ( .A1(n15103), .A2(n15104), .ZN(n9426) );
  NOR2_X1 U12096 ( .A1(n15103), .A2(n15104), .ZN(n15102) );
  AOI21_X1 U12097 ( .B1(n9427), .B2(n9426), .A(n15102), .ZN(n15752) );
  XNOR2_X1 U12098 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n9428), .ZN(n15751) );
  NAND2_X1 U12099 ( .A1(n15752), .A2(n15751), .ZN(n9429) );
  NOR2_X1 U12100 ( .A1(n15752), .A2(n15751), .ZN(n15750) );
  AOI21_X1 U12101 ( .B1(n15359), .B2(n9429), .A(n15750), .ZN(n15742) );
  NAND2_X1 U12102 ( .A1(n15743), .A2(n15742), .ZN(n9430) );
  NOR2_X1 U12103 ( .A1(n15107), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9437) );
  XOR2_X1 U12104 ( .A(n9716), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n9436) );
  XNOR2_X1 U12105 ( .A(n9436), .B(n9435), .ZN(n15109) );
  NAND2_X1 U12106 ( .A1(n15107), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n15106) );
  NAND2_X1 U12107 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n9438), .ZN(n9440) );
  INV_X1 U12108 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n15410) );
  XNOR2_X1 U12109 ( .A(n15410), .B(n9438), .ZN(n15749) );
  XNOR2_X1 U12110 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9439), .ZN(n15748) );
  XNOR2_X1 U12111 ( .A(n9442), .B(n9441), .ZN(n9443) );
  NOR2_X1 U12112 ( .A1(n9444), .A2(n9443), .ZN(n9446) );
  XNOR2_X1 U12113 ( .A(n9444), .B(n9443), .ZN(n15110) );
  NOR2_X1 U12114 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n15110), .ZN(n9445) );
  XNOR2_X1 U12115 ( .A(n9448), .B(n9447), .ZN(n9450) );
  NAND2_X1 U12116 ( .A1(n9449), .A2(n9450), .ZN(n9452) );
  NAND2_X1 U12117 ( .A1(n15111), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n9451) );
  NAND2_X1 U12118 ( .A1(n9452), .A2(n9451), .ZN(n15113) );
  XOR2_X1 U12119 ( .A(n9454), .B(n9453), .Z(n9456) );
  NOR2_X1 U12120 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n15233), .ZN(n9457) );
  XNOR2_X1 U12121 ( .A(n9459), .B(n9458), .ZN(n15237) );
  XOR2_X1 U12122 ( .A(n9460), .B(P3_ADDR_REG_13__SCAN_IN), .Z(n9462) );
  XOR2_X1 U12123 ( .A(n9462), .B(n9461), .Z(n9463) );
  NOR2_X1 U12124 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(n15240), .ZN(n9465) );
  NAND2_X1 U12125 ( .A1(n15244), .A2(n15245), .ZN(n9466) );
  NOR2_X1 U12126 ( .A1(n15244), .A2(n15245), .ZN(n15243) );
  AOI21_X2 U12127 ( .B1(n9467), .B2(n9466), .A(n15243), .ZN(n15248) );
  OAI21_X1 U12128 ( .B1(n9469), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n9468), .ZN(
        n9471) );
  XOR2_X1 U12129 ( .A(n9471), .B(n9470), .Z(n15249) );
  INV_X1 U12130 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n15448) );
  NAND2_X1 U12131 ( .A1(n15248), .A2(n15249), .ZN(n15247) );
  INV_X1 U12132 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n15460) );
  INV_X1 U12133 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n15133) );
  NAND2_X1 U12134 ( .A1(n9473), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9477) );
  NAND2_X1 U12135 ( .A1(n9475), .A2(n9474), .ZN(n9476) );
  NAND2_X1 U12136 ( .A1(n9477), .A2(n9476), .ZN(n9481) );
  XNOR2_X1 U12137 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n9481), .ZN(n9482) );
  XNOR2_X1 U12138 ( .A(n15133), .B(n9482), .ZN(n9478) );
  NOR2_X1 U12139 ( .A1(n9479), .A2(n9478), .ZN(n15123) );
  NOR2_X1 U12140 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n15122), .ZN(n9480) );
  NOR2_X1 U12141 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n9481), .ZN(n9484) );
  NOR2_X1 U12142 ( .A1(n15133), .A2(n9482), .ZN(n9483) );
  NOR2_X1 U12143 ( .A1(n9484), .A2(n9483), .ZN(n9488) );
  INV_X1 U12144 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9490) );
  XNOR2_X1 U12145 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(n9490), .ZN(n9487) );
  XOR2_X1 U12146 ( .A(n9488), .B(n9487), .Z(n9486) );
  AND2_X2 U12147 ( .A1(n9485), .A2(n9486), .ZN(n15100) );
  NOR2_X1 U12148 ( .A1(n9488), .A2(n9487), .ZN(n9489) );
  AOI21_X1 U12149 ( .B1(P3_ADDR_REG_18__SCAN_IN), .B2(n9490), .A(n9489), .ZN(
        n9493) );
  XNOR2_X1 U12150 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n9491) );
  XNOR2_X1 U12151 ( .A(n14769), .B(n9491), .ZN(n9492) );
  XNOR2_X1 U12152 ( .A(n9493), .B(n9492), .ZN(n9832) );
  AOI22_X1 U12153 ( .A1(keyinput_f82), .A2(P3_DATAO_REG_14__SCAN_IN), .B1(
        keyinput_f68), .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n9494) );
  OAI221_X1 U12154 ( .B1(keyinput_f82), .B2(P3_DATAO_REG_14__SCAN_IN), .C1(
        keyinput_f68), .C2(P3_DATAO_REG_28__SCAN_IN), .A(n9494), .ZN(n9501) );
  AOI22_X1 U12155 ( .A1(keyinput_f70), .A2(P3_DATAO_REG_26__SCAN_IN), .B1(
        P1_IR_REG_2__SCAN_IN), .B2(keyinput_f109), .ZN(n9495) );
  OAI221_X1 U12156 ( .B1(keyinput_f70), .B2(P3_DATAO_REG_26__SCAN_IN), .C1(
        P1_IR_REG_2__SCAN_IN), .C2(keyinput_f109), .A(n9495), .ZN(n9500) );
  AOI22_X1 U12157 ( .A1(keyinput_f95), .A2(P3_DATAO_REG_1__SCAN_IN), .B1(
        P1_IR_REG_13__SCAN_IN), .B2(keyinput_f120), .ZN(n9496) );
  OAI221_X1 U12158 ( .B1(keyinput_f95), .B2(P3_DATAO_REG_1__SCAN_IN), .C1(
        P1_IR_REG_13__SCAN_IN), .C2(keyinput_f120), .A(n9496), .ZN(n9499) );
  AOI22_X1 U12159 ( .A1(P3_ADDR_REG_0__SCAN_IN), .A2(keyinput_f97), .B1(
        keyinput_f78), .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n9497) );
  OAI221_X1 U12160 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(keyinput_f97), .C1(
        keyinput_f78), .C2(P3_DATAO_REG_18__SCAN_IN), .A(n9497), .ZN(n9498) );
  NOR4_X1 U12161 ( .A1(n9501), .A2(n9500), .A3(n9499), .A4(n9498), .ZN(n9654)
         );
  AOI22_X1 U12162 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(keyinput_f101), .B1(
        P3_REG3_REG_19__SCAN_IN), .B2(keyinput_f41), .ZN(n9502) );
  OAI221_X1 U12163 ( .B1(P3_ADDR_REG_4__SCAN_IN), .B2(keyinput_f101), .C1(
        P3_REG3_REG_19__SCAN_IN), .C2(keyinput_f41), .A(n9502), .ZN(n9527) );
  OAI22_X1 U12164 ( .A1(SI_16_), .A2(keyinput_f16), .B1(SI_6_), .B2(
        keyinput_f26), .ZN(n9503) );
  AOI221_X1 U12165 ( .B1(SI_16_), .B2(keyinput_f16), .C1(keyinput_f26), .C2(
        SI_6_), .A(n9503), .ZN(n9507) );
  AOI22_X1 U12166 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(keyinput_f51), .B1(
        P3_B_REG_SCAN_IN), .B2(keyinput_f64), .ZN(n9504) );
  OAI221_X1 U12167 ( .B1(P3_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .C1(
        P3_B_REG_SCAN_IN), .C2(keyinput_f64), .A(n9504), .ZN(n9505) );
  AOI21_X1 U12168 ( .B1(keyinput_f4), .B2(n12851), .A(n9505), .ZN(n9506) );
  OAI211_X1 U12169 ( .C1(keyinput_f4), .C2(n12851), .A(n9507), .B(n9506), .ZN(
        n9526) );
  OAI22_X1 U12170 ( .A1(SI_29_), .A2(keyinput_f3), .B1(keyinput_f15), .B2(
        SI_17_), .ZN(n9508) );
  AOI221_X1 U12171 ( .B1(SI_29_), .B2(keyinput_f3), .C1(SI_17_), .C2(
        keyinput_f15), .A(n9508), .ZN(n9515) );
  OAI22_X1 U12172 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(keyinput_f60), .B1(
        keyinput_f6), .B2(SI_26_), .ZN(n9509) );
  AOI221_X1 U12173 ( .B1(P3_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .C1(
        SI_26_), .C2(keyinput_f6), .A(n9509), .ZN(n9514) );
  OAI22_X1 U12174 ( .A1(SI_0_), .A2(keyinput_f32), .B1(
        P3_DATAO_REG_24__SCAN_IN), .B2(keyinput_f72), .ZN(n9510) );
  AOI221_X1 U12175 ( .B1(SI_0_), .B2(keyinput_f32), .C1(keyinput_f72), .C2(
        P3_DATAO_REG_24__SCAN_IN), .A(n9510), .ZN(n9513) );
  OAI22_X1 U12176 ( .A1(P3_REG3_REG_28__SCAN_IN), .A2(keyinput_f42), .B1(
        keyinput_f85), .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n9511) );
  AOI221_X1 U12177 ( .B1(P3_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .C1(
        P3_DATAO_REG_11__SCAN_IN), .C2(keyinput_f85), .A(n9511), .ZN(n9512) );
  NAND4_X1 U12178 ( .A1(n9515), .A2(n9514), .A3(n9513), .A4(n9512), .ZN(n9525)
         );
  OAI22_X1 U12179 ( .A1(keyinput_f71), .A2(P3_DATAO_REG_25__SCAN_IN), .B1(
        P3_RD_REG_SCAN_IN), .B2(keyinput_f33), .ZN(n9516) );
  AOI221_X1 U12180 ( .B1(keyinput_f71), .B2(P3_DATAO_REG_25__SCAN_IN), .C1(
        keyinput_f33), .C2(P3_RD_REG_SCAN_IN), .A(n9516), .ZN(n9523) );
  OAI22_X1 U12181 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(keyinput_f43), .B1(SI_2_), 
        .B2(keyinput_f30), .ZN(n9517) );
  AOI221_X1 U12182 ( .B1(P3_REG3_REG_8__SCAN_IN), .B2(keyinput_f43), .C1(
        keyinput_f30), .C2(SI_2_), .A(n9517), .ZN(n9522) );
  OAI22_X1 U12183 ( .A1(P3_REG3_REG_25__SCAN_IN), .A2(keyinput_f47), .B1(
        keyinput_f96), .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n9518) );
  AOI221_X1 U12184 ( .B1(P3_REG3_REG_25__SCAN_IN), .B2(keyinput_f47), .C1(
        P3_DATAO_REG_0__SCAN_IN), .C2(keyinput_f96), .A(n9518), .ZN(n9521) );
  OAI22_X1 U12185 ( .A1(SI_31_), .A2(keyinput_f1), .B1(
        P3_DATAO_REG_29__SCAN_IN), .B2(keyinput_f67), .ZN(n9519) );
  AOI221_X1 U12186 ( .B1(SI_31_), .B2(keyinput_f1), .C1(keyinput_f67), .C2(
        P3_DATAO_REG_29__SCAN_IN), .A(n9519), .ZN(n9520) );
  NAND4_X1 U12187 ( .A1(n9523), .A2(n9522), .A3(n9521), .A4(n9520), .ZN(n9524)
         );
  NOR4_X1 U12188 ( .A1(n9527), .A2(n9526), .A3(n9525), .A4(n9524), .ZN(n9653)
         );
  OAI22_X1 U12189 ( .A1(SI_9_), .A2(keyinput_f23), .B1(
        P3_DATAO_REG_19__SCAN_IN), .B2(keyinput_f77), .ZN(n9528) );
  AOI221_X1 U12190 ( .B1(SI_9_), .B2(keyinput_f23), .C1(keyinput_f77), .C2(
        P3_DATAO_REG_19__SCAN_IN), .A(n9528), .ZN(n9535) );
  OAI22_X1 U12191 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(keyinput_f112), .B1(
        P3_DATAO_REG_16__SCAN_IN), .B2(keyinput_f80), .ZN(n9529) );
  AOI221_X1 U12192 ( .B1(P1_IR_REG_5__SCAN_IN), .B2(keyinput_f112), .C1(
        keyinput_f80), .C2(P3_DATAO_REG_16__SCAN_IN), .A(n9529), .ZN(n9534) );
  OAI22_X1 U12193 ( .A1(P3_DATAO_REG_5__SCAN_IN), .A2(keyinput_f91), .B1(
        P3_ADDR_REG_6__SCAN_IN), .B2(keyinput_f103), .ZN(n9530) );
  AOI221_X1 U12194 ( .B1(P3_DATAO_REG_5__SCAN_IN), .B2(keyinput_f91), .C1(
        keyinput_f103), .C2(P3_ADDR_REG_6__SCAN_IN), .A(n9530), .ZN(n9533) );
  OAI22_X1 U12195 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(keyinput_f61), .B1(
        P1_IR_REG_15__SCAN_IN), .B2(keyinput_f122), .ZN(n9531) );
  AOI221_X1 U12196 ( .B1(P3_REG3_REG_6__SCAN_IN), .B2(keyinput_f61), .C1(
        keyinput_f122), .C2(P1_IR_REG_15__SCAN_IN), .A(n9531), .ZN(n9532) );
  NAND4_X1 U12197 ( .A1(n9535), .A2(n9534), .A3(n9533), .A4(n9532), .ZN(n9563)
         );
  OAI22_X1 U12198 ( .A1(P3_REG3_REG_7__SCAN_IN), .A2(keyinput_f35), .B1(
        keyinput_f121), .B2(P1_IR_REG_14__SCAN_IN), .ZN(n9536) );
  AOI221_X1 U12199 ( .B1(P3_REG3_REG_7__SCAN_IN), .B2(keyinput_f35), .C1(
        P1_IR_REG_14__SCAN_IN), .C2(keyinput_f121), .A(n9536), .ZN(n9543) );
  OAI22_X1 U12200 ( .A1(P3_STATE_REG_SCAN_IN), .A2(keyinput_f34), .B1(
        keyinput_f98), .B2(P3_ADDR_REG_1__SCAN_IN), .ZN(n9537) );
  AOI221_X1 U12201 ( .B1(P3_STATE_REG_SCAN_IN), .B2(keyinput_f34), .C1(
        P3_ADDR_REG_1__SCAN_IN), .C2(keyinput_f98), .A(n9537), .ZN(n9542) );
  OAI22_X1 U12202 ( .A1(P3_REG3_REG_5__SCAN_IN), .A2(keyinput_f49), .B1(
        P1_IR_REG_16__SCAN_IN), .B2(keyinput_f123), .ZN(n9538) );
  AOI221_X1 U12203 ( .B1(P3_REG3_REG_5__SCAN_IN), .B2(keyinput_f49), .C1(
        keyinput_f123), .C2(P1_IR_REG_16__SCAN_IN), .A(n9538), .ZN(n9541) );
  OAI22_X1 U12204 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(keyinput_f48), .B1(
        keyinput_f46), .B2(P3_REG3_REG_12__SCAN_IN), .ZN(n9539) );
  AOI221_X1 U12205 ( .B1(P3_REG3_REG_16__SCAN_IN), .B2(keyinput_f48), .C1(
        P3_REG3_REG_12__SCAN_IN), .C2(keyinput_f46), .A(n9539), .ZN(n9540) );
  NAND4_X1 U12206 ( .A1(n9543), .A2(n9542), .A3(n9541), .A4(n9540), .ZN(n9562)
         );
  OAI22_X1 U12207 ( .A1(SI_13_), .A2(keyinput_f19), .B1(keyinput_f73), .B2(
        P3_DATAO_REG_23__SCAN_IN), .ZN(n9544) );
  AOI221_X1 U12208 ( .B1(SI_13_), .B2(keyinput_f19), .C1(
        P3_DATAO_REG_23__SCAN_IN), .C2(keyinput_f73), .A(n9544), .ZN(n9551) );
  OAI22_X1 U12209 ( .A1(keyinput_f105), .A2(P3_ADDR_REG_8__SCAN_IN), .B1(
        keyinput_f87), .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n9545) );
  AOI221_X1 U12210 ( .B1(keyinput_f105), .B2(P3_ADDR_REG_8__SCAN_IN), .C1(
        P3_DATAO_REG_9__SCAN_IN), .C2(keyinput_f87), .A(n9545), .ZN(n9550) );
  OAI22_X1 U12211 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(keyinput_f108), .B1(
        P3_ADDR_REG_5__SCAN_IN), .B2(keyinput_f102), .ZN(n9546) );
  AOI221_X1 U12212 ( .B1(P1_IR_REG_1__SCAN_IN), .B2(keyinput_f108), .C1(
        keyinput_f102), .C2(P3_ADDR_REG_5__SCAN_IN), .A(n9546), .ZN(n9549) );
  OAI22_X1 U12213 ( .A1(P3_REG3_REG_2__SCAN_IN), .A2(keyinput_f59), .B1(
        keyinput_f12), .B2(SI_20_), .ZN(n9547) );
  AOI221_X1 U12214 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(keyinput_f59), .C1(
        SI_20_), .C2(keyinput_f12), .A(n9547), .ZN(n9548) );
  NAND4_X1 U12215 ( .A1(n9551), .A2(n9550), .A3(n9549), .A4(n9548), .ZN(n9561)
         );
  OAI22_X1 U12216 ( .A1(P3_REG3_REG_26__SCAN_IN), .A2(keyinput_f62), .B1(
        SI_27_), .B2(keyinput_f5), .ZN(n9552) );
  AOI221_X1 U12217 ( .B1(P3_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .C1(
        keyinput_f5), .C2(SI_27_), .A(n9552), .ZN(n9559) );
  OAI22_X1 U12218 ( .A1(P3_REG3_REG_1__SCAN_IN), .A2(keyinput_f44), .B1(
        keyinput_f115), .B2(P1_IR_REG_8__SCAN_IN), .ZN(n9553) );
  AOI221_X1 U12219 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(keyinput_f44), .C1(
        P1_IR_REG_8__SCAN_IN), .C2(keyinput_f115), .A(n9553), .ZN(n9558) );
  OAI22_X1 U12220 ( .A1(P3_REG3_REG_21__SCAN_IN), .A2(keyinput_f45), .B1(
        keyinput_f116), .B2(P1_IR_REG_9__SCAN_IN), .ZN(n9554) );
  AOI221_X1 U12221 ( .B1(P3_REG3_REG_21__SCAN_IN), .B2(keyinput_f45), .C1(
        P1_IR_REG_9__SCAN_IN), .C2(keyinput_f116), .A(n9554), .ZN(n9557) );
  OAI22_X1 U12222 ( .A1(SI_12_), .A2(keyinput_f20), .B1(P1_IR_REG_20__SCAN_IN), 
        .B2(keyinput_f127), .ZN(n9555) );
  AOI221_X1 U12223 ( .B1(SI_12_), .B2(keyinput_f20), .C1(keyinput_f127), .C2(
        P1_IR_REG_20__SCAN_IN), .A(n9555), .ZN(n9556) );
  NAND4_X1 U12224 ( .A1(n9559), .A2(n9558), .A3(n9557), .A4(n9556), .ZN(n9560)
         );
  NOR4_X1 U12225 ( .A1(n9563), .A2(n9562), .A3(n9561), .A4(n9560), .ZN(n9652)
         );
  OAI22_X1 U12226 ( .A1(P3_REG3_REG_23__SCAN_IN), .A2(keyinput_f38), .B1(
        P3_DATAO_REG_8__SCAN_IN), .B2(keyinput_f88), .ZN(n9564) );
  AOI221_X1 U12227 ( .B1(P3_REG3_REG_23__SCAN_IN), .B2(keyinput_f38), .C1(
        keyinput_f88), .C2(P3_DATAO_REG_8__SCAN_IN), .A(n9564), .ZN(n9571) );
  OAI22_X1 U12228 ( .A1(SI_25_), .A2(keyinput_f7), .B1(SI_19_), .B2(
        keyinput_f13), .ZN(n9565) );
  AOI221_X1 U12229 ( .B1(SI_25_), .B2(keyinput_f7), .C1(keyinput_f13), .C2(
        SI_19_), .A(n9565), .ZN(n9570) );
  OAI22_X1 U12230 ( .A1(P3_REG3_REG_11__SCAN_IN), .A2(keyinput_f58), .B1(
        keyinput_f75), .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n9566) );
  AOI221_X1 U12231 ( .B1(P3_REG3_REG_11__SCAN_IN), .B2(keyinput_f58), .C1(
        P3_DATAO_REG_21__SCAN_IN), .C2(keyinput_f75), .A(n9566), .ZN(n9569) );
  OAI22_X1 U12232 ( .A1(SI_23_), .A2(keyinput_f9), .B1(keyinput_f29), .B2(
        SI_3_), .ZN(n9567) );
  AOI221_X1 U12233 ( .B1(SI_23_), .B2(keyinput_f9), .C1(SI_3_), .C2(
        keyinput_f29), .A(n9567), .ZN(n9568) );
  NAND4_X1 U12234 ( .A1(n9571), .A2(n9570), .A3(n9569), .A4(n9568), .ZN(n9650)
         );
  INV_X1 U12235 ( .A(P3_WR_REG_SCAN_IN), .ZN(n9808) );
  XNOR2_X1 U12236 ( .A(keyinput_f0), .B(n9808), .ZN(n9578) );
  INV_X1 U12237 ( .A(P3_DATAO_REG_2__SCAN_IN), .ZN(n10718) );
  XNOR2_X1 U12238 ( .A(n10718), .B(keyinput_f94), .ZN(n9577) );
  XNOR2_X1 U12239 ( .A(SI_5_), .B(keyinput_f27), .ZN(n9575) );
  XNOR2_X1 U12240 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_f110), .ZN(n9574) );
  XNOR2_X1 U12241 ( .A(P3_REG3_REG_27__SCAN_IN), .B(keyinput_f36), .ZN(n9573)
         );
  XNOR2_X1 U12242 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_f126), .ZN(n9572)
         );
  NAND4_X1 U12243 ( .A1(n9575), .A2(n9574), .A3(n9573), .A4(n9572), .ZN(n9576)
         );
  OR3_X1 U12244 ( .A1(n9578), .A2(n9577), .A3(n9576), .ZN(n9583) );
  AOI22_X1 U12245 ( .A1(n10415), .A2(keyinput_f22), .B1(n11937), .B2(
        keyinput_f8), .ZN(n9579) );
  OAI221_X1 U12246 ( .B1(n10415), .B2(keyinput_f22), .C1(n11937), .C2(
        keyinput_f8), .A(n9579), .ZN(n9582) );
  INV_X1 U12247 ( .A(P3_DATAO_REG_27__SCAN_IN), .ZN(n11445) );
  INV_X1 U12248 ( .A(P3_DATAO_REG_3__SCAN_IN), .ZN(n10720) );
  AOI22_X1 U12249 ( .A1(n11445), .A2(keyinput_f69), .B1(keyinput_f93), .B2(
        n10720), .ZN(n9580) );
  OAI221_X1 U12250 ( .B1(n11445), .B2(keyinput_f69), .C1(n10720), .C2(
        keyinput_f93), .A(n9580), .ZN(n9581) );
  NOR3_X1 U12251 ( .A1(n9583), .A2(n9582), .A3(n9581), .ZN(n9602) );
  AOI22_X1 U12252 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(keyinput_f111), .B1(SI_1_), 
        .B2(keyinput_f31), .ZN(n9584) );
  OAI221_X1 U12253 ( .B1(P1_IR_REG_4__SCAN_IN), .B2(keyinput_f111), .C1(SI_1_), 
        .C2(keyinput_f31), .A(n9584), .ZN(n9591) );
  INV_X1 U12254 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n11576) );
  AOI22_X1 U12255 ( .A1(n11576), .A2(keyinput_f52), .B1(keyinput_f14), .B2(
        n10739), .ZN(n9585) );
  OAI221_X1 U12256 ( .B1(n11576), .B2(keyinput_f52), .C1(n10739), .C2(
        keyinput_f14), .A(n9585), .ZN(n9590) );
  INV_X1 U12257 ( .A(P3_DATAO_REG_20__SCAN_IN), .ZN(n10804) );
  AOI22_X1 U12258 ( .A1(n10804), .A2(keyinput_f76), .B1(n10457), .B2(
        keyinput_f18), .ZN(n9586) );
  OAI221_X1 U12259 ( .B1(n10804), .B2(keyinput_f76), .C1(n10457), .C2(
        keyinput_f18), .A(n9586), .ZN(n9589) );
  INV_X1 U12260 ( .A(SI_30_), .ZN(n13381) );
  INV_X1 U12261 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n13494) );
  AOI22_X1 U12262 ( .A1(n13381), .A2(keyinput_f2), .B1(n13494), .B2(
        keyinput_f57), .ZN(n9587) );
  OAI221_X1 U12263 ( .B1(n13381), .B2(keyinput_f2), .C1(n13494), .C2(
        keyinput_f57), .A(n9587), .ZN(n9588) );
  NOR4_X1 U12264 ( .A1(n9591), .A2(n9590), .A3(n9589), .A4(n9588), .ZN(n9601)
         );
  XOR2_X1 U12265 ( .A(keyinput_f104), .B(n9592), .Z(n9600) );
  INV_X1 U12266 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n11914) );
  AOI22_X1 U12267 ( .A1(n10422), .A2(keyinput_f21), .B1(n11914), .B2(
        keyinput_f39), .ZN(n9593) );
  OAI221_X1 U12268 ( .B1(n10422), .B2(keyinput_f21), .C1(n11914), .C2(
        keyinput_f39), .A(n9593), .ZN(n9598) );
  XOR2_X1 U12269 ( .A(SI_22_), .B(keyinput_f10), .Z(n9597) );
  XNOR2_X1 U12270 ( .A(n9594), .B(keyinput_f119), .ZN(n9596) );
  XNOR2_X1 U12271 ( .A(n10497), .B(keyinput_f17), .ZN(n9595) );
  NOR4_X1 U12272 ( .A1(n9598), .A2(n9597), .A3(n9596), .A4(n9595), .ZN(n9599)
         );
  NAND4_X1 U12273 ( .A1(n9602), .A2(n9601), .A3(n9600), .A4(n9599), .ZN(n9649)
         );
  INV_X1 U12274 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n13386) );
  OAI22_X1 U12275 ( .A1(n13386), .A2(keyinput_f37), .B1(n9013), .B2(
        keyinput_f56), .ZN(n9603) );
  AOI221_X1 U12276 ( .B1(n13386), .B2(keyinput_f37), .C1(keyinput_f56), .C2(
        n9013), .A(n9603), .ZN(n9612) );
  INV_X1 U12277 ( .A(P3_DATAO_REG_22__SCAN_IN), .ZN(n10883) );
  INV_X1 U12278 ( .A(P3_DATAO_REG_7__SCAN_IN), .ZN(n10767) );
  OAI22_X1 U12279 ( .A1(n10883), .A2(keyinput_f74), .B1(n10767), .B2(
        keyinput_f89), .ZN(n9604) );
  AOI221_X1 U12280 ( .B1(n10883), .B2(keyinput_f74), .C1(keyinput_f89), .C2(
        n10767), .A(n9604), .ZN(n9611) );
  INV_X1 U12281 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n10791) );
  XNOR2_X1 U12282 ( .A(n10791), .B(keyinput_f79), .ZN(n9609) );
  XOR2_X1 U12283 ( .A(SI_21_), .B(keyinput_f11), .Z(n9608) );
  INV_X1 U12284 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10666) );
  XNOR2_X1 U12285 ( .A(n10666), .B(keyinput_f107), .ZN(n9607) );
  XNOR2_X1 U12286 ( .A(n9605), .B(keyinput_f113), .ZN(n9606) );
  NOR4_X1 U12287 ( .A1(n9609), .A2(n9608), .A3(n9607), .A4(n9606), .ZN(n9610)
         );
  NAND3_X1 U12288 ( .A1(n9612), .A2(n9611), .A3(n9610), .ZN(n9648) );
  INV_X1 U12289 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n11284) );
  INV_X1 U12290 ( .A(P3_DATAO_REG_12__SCAN_IN), .ZN(n10789) );
  AOI22_X1 U12291 ( .A1(n11284), .A2(keyinput_f40), .B1(keyinput_f84), .B2(
        n10789), .ZN(n9613) );
  OAI221_X1 U12292 ( .B1(n11284), .B2(keyinput_f40), .C1(n10789), .C2(
        keyinput_f84), .A(n9613), .ZN(n9621) );
  INV_X1 U12293 ( .A(P3_DATAO_REG_13__SCAN_IN), .ZN(n10760) );
  INV_X1 U12294 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n11527) );
  AOI22_X1 U12295 ( .A1(n10760), .A2(keyinput_f83), .B1(keyinput_f65), .B2(
        n11527), .ZN(n9614) );
  OAI221_X1 U12296 ( .B1(n10760), .B2(keyinput_f83), .C1(n11527), .C2(
        keyinput_f65), .A(n9614), .ZN(n9620) );
  INV_X1 U12297 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n9616) );
  AOI22_X1 U12298 ( .A1(n9616), .A2(keyinput_f99), .B1(n8931), .B2(
        keyinput_f53), .ZN(n9615) );
  OAI221_X1 U12299 ( .B1(n9616), .B2(keyinput_f99), .C1(n8931), .C2(
        keyinput_f53), .A(n9615), .ZN(n9619) );
  INV_X1 U12300 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9753) );
  AOI22_X1 U12301 ( .A1(n9733), .A2(keyinput_f118), .B1(n9753), .B2(
        keyinput_f124), .ZN(n9617) );
  OAI221_X1 U12302 ( .B1(n9733), .B2(keyinput_f118), .C1(n9753), .C2(
        keyinput_f124), .A(n9617), .ZN(n9618) );
  NOR4_X1 U12303 ( .A1(n9621), .A2(n9620), .A3(n9619), .A4(n9618), .ZN(n9646)
         );
  INV_X1 U12304 ( .A(P3_DATAO_REG_15__SCAN_IN), .ZN(n10756) );
  OAI22_X1 U12305 ( .A1(keyinput_f106), .A2(n9806), .B1(n10756), .B2(
        keyinput_f81), .ZN(n9622) );
  AOI221_X1 U12306 ( .B1(n9806), .B2(keyinput_f106), .C1(n10756), .C2(
        keyinput_f81), .A(n9622), .ZN(n9645) );
  INV_X1 U12307 ( .A(P3_DATAO_REG_10__SCAN_IN), .ZN(n9624) );
  AOI22_X1 U12308 ( .A1(n9624), .A2(keyinput_f86), .B1(keyinput_f100), .B2(
        n9796), .ZN(n9623) );
  OAI221_X1 U12309 ( .B1(n9624), .B2(keyinput_f86), .C1(n9796), .C2(
        keyinput_f100), .A(n9623), .ZN(n9630) );
  XNOR2_X1 U12310 ( .A(SI_8_), .B(keyinput_f24), .ZN(n9628) );
  XNOR2_X1 U12311 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_f114), .ZN(n9627) );
  XNOR2_X1 U12312 ( .A(P3_REG3_REG_20__SCAN_IN), .B(keyinput_f55), .ZN(n9626)
         );
  XNOR2_X1 U12313 ( .A(SI_7_), .B(keyinput_f25), .ZN(n9625) );
  NAND4_X1 U12314 ( .A1(n9628), .A2(n9627), .A3(n9626), .A4(n9625), .ZN(n9629)
         );
  NOR2_X1 U12315 ( .A1(n9630), .A2(n9629), .ZN(n9644) );
  INV_X1 U12316 ( .A(P3_DATAO_REG_4__SCAN_IN), .ZN(n10758) );
  AOI22_X1 U12317 ( .A1(n11367), .A2(keyinput_f54), .B1(keyinput_f92), .B2(
        n10758), .ZN(n9631) );
  OAI221_X1 U12318 ( .B1(n11367), .B2(keyinput_f54), .C1(n10758), .C2(
        keyinput_f92), .A(n9631), .ZN(n9642) );
  INV_X1 U12319 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n11510) );
  INV_X1 U12320 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n13513) );
  AOI22_X1 U12321 ( .A1(n11510), .A2(keyinput_f66), .B1(n13513), .B2(
        keyinput_f63), .ZN(n9632) );
  OAI221_X1 U12322 ( .B1(n11510), .B2(keyinput_f66), .C1(n13513), .C2(
        keyinput_f63), .A(n9632), .ZN(n9641) );
  INV_X1 U12323 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n9634) );
  AOI22_X1 U12324 ( .A1(n9635), .A2(keyinput_f50), .B1(keyinput_f117), .B2(
        n9634), .ZN(n9633) );
  OAI221_X1 U12325 ( .B1(n9635), .B2(keyinput_f50), .C1(n9634), .C2(
        keyinput_f117), .A(n9633), .ZN(n9640) );
  INV_X1 U12326 ( .A(P3_DATAO_REG_6__SCAN_IN), .ZN(n9636) );
  XOR2_X1 U12327 ( .A(n9636), .B(keyinput_f90), .Z(n9638) );
  XNOR2_X1 U12328 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_f125), .ZN(n9637)
         );
  NAND2_X1 U12329 ( .A1(n9638), .A2(n9637), .ZN(n9639) );
  NOR4_X1 U12330 ( .A1(n9642), .A2(n9641), .A3(n9640), .A4(n9639), .ZN(n9643)
         );
  NAND4_X1 U12331 ( .A1(n9646), .A2(n9645), .A3(n9644), .A4(n9643), .ZN(n9647)
         );
  NOR4_X1 U12332 ( .A1(n9650), .A2(n9649), .A3(n9648), .A4(n9647), .ZN(n9651)
         );
  NAND4_X1 U12333 ( .A1(n9654), .A2(n9653), .A3(n9652), .A4(n9651), .ZN(n9829)
         );
  INV_X1 U12334 ( .A(keyinput_f28), .ZN(n9655) );
  MUX2_X1 U12335 ( .A(keyinput_f28), .B(n9655), .S(SI_4_), .Z(n9828) );
  XOR2_X1 U12336 ( .A(SI_4_), .B(keyinput_g28), .Z(n9827) );
  XNOR2_X1 U12337 ( .A(n11527), .B(keyinput_g65), .ZN(n9662) );
  AOI22_X1 U12338 ( .A1(P3_DATAO_REG_15__SCAN_IN), .A2(keyinput_g81), .B1(
        P1_IR_REG_19__SCAN_IN), .B2(keyinput_g126), .ZN(n9656) );
  OAI221_X1 U12339 ( .B1(P3_DATAO_REG_15__SCAN_IN), .B2(keyinput_g81), .C1(
        P1_IR_REG_19__SCAN_IN), .C2(keyinput_g126), .A(n9656), .ZN(n9661) );
  AOI22_X1 U12340 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(keyinput_g99), .B1(SI_16_), .B2(keyinput_g16), .ZN(n9657) );
  OAI221_X1 U12341 ( .B1(P3_ADDR_REG_2__SCAN_IN), .B2(keyinput_g99), .C1(
        SI_16_), .C2(keyinput_g16), .A(n9657), .ZN(n9660) );
  AOI22_X1 U12342 ( .A1(P3_DATAO_REG_26__SCAN_IN), .A2(keyinput_g70), .B1(
        P3_REG3_REG_26__SCAN_IN), .B2(keyinput_g62), .ZN(n9658) );
  OAI221_X1 U12343 ( .B1(P3_DATAO_REG_26__SCAN_IN), .B2(keyinput_g70), .C1(
        P3_REG3_REG_26__SCAN_IN), .C2(keyinput_g62), .A(n9658), .ZN(n9659) );
  NOR4_X1 U12344 ( .A1(n9662), .A2(n9661), .A3(n9660), .A4(n9659), .ZN(n9690)
         );
  AOI22_X1 U12345 ( .A1(P3_DATAO_REG_30__SCAN_IN), .A2(keyinput_g66), .B1(
        P3_ADDR_REG_7__SCAN_IN), .B2(keyinput_g104), .ZN(n9663) );
  OAI221_X1 U12346 ( .B1(P3_DATAO_REG_30__SCAN_IN), .B2(keyinput_g66), .C1(
        P3_ADDR_REG_7__SCAN_IN), .C2(keyinput_g104), .A(n9663), .ZN(n9670) );
  AOI22_X1 U12347 ( .A1(P3_DATAO_REG_28__SCAN_IN), .A2(keyinput_g68), .B1(
        P1_IR_REG_0__SCAN_IN), .B2(keyinput_g107), .ZN(n9664) );
  OAI221_X1 U12348 ( .B1(P3_DATAO_REG_28__SCAN_IN), .B2(keyinput_g68), .C1(
        P1_IR_REG_0__SCAN_IN), .C2(keyinput_g107), .A(n9664), .ZN(n9669) );
  AOI22_X1 U12349 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(keyinput_g117), .B1(
        P3_REG3_REG_10__SCAN_IN), .B2(keyinput_g39), .ZN(n9665) );
  OAI221_X1 U12350 ( .B1(P1_IR_REG_10__SCAN_IN), .B2(keyinput_g117), .C1(
        P3_REG3_REG_10__SCAN_IN), .C2(keyinput_g39), .A(n9665), .ZN(n9668) );
  AOI22_X1 U12351 ( .A1(P3_DATAO_REG_11__SCAN_IN), .A2(keyinput_g85), .B1(
        SI_23_), .B2(keyinput_g9), .ZN(n9666) );
  OAI221_X1 U12352 ( .B1(P3_DATAO_REG_11__SCAN_IN), .B2(keyinput_g85), .C1(
        SI_23_), .C2(keyinput_g9), .A(n9666), .ZN(n9667) );
  NOR4_X1 U12353 ( .A1(n9670), .A2(n9669), .A3(n9668), .A4(n9667), .ZN(n9689)
         );
  AOI22_X1 U12354 ( .A1(P3_DATAO_REG_16__SCAN_IN), .A2(keyinput_g80), .B1(
        SI_30_), .B2(keyinput_g2), .ZN(n9671) );
  OAI221_X1 U12355 ( .B1(P3_DATAO_REG_16__SCAN_IN), .B2(keyinput_g80), .C1(
        SI_30_), .C2(keyinput_g2), .A(n9671), .ZN(n9678) );
  AOI22_X1 U12356 ( .A1(P3_DATAO_REG_22__SCAN_IN), .A2(keyinput_g74), .B1(
        SI_17_), .B2(keyinput_g15), .ZN(n9672) );
  OAI221_X1 U12357 ( .B1(P3_DATAO_REG_22__SCAN_IN), .B2(keyinput_g74), .C1(
        SI_17_), .C2(keyinput_g15), .A(n9672), .ZN(n9677) );
  AOI22_X1 U12358 ( .A1(SI_12_), .A2(keyinput_g20), .B1(
        P3_REG3_REG_12__SCAN_IN), .B2(keyinput_g46), .ZN(n9673) );
  OAI221_X1 U12359 ( .B1(SI_12_), .B2(keyinput_g20), .C1(
        P3_REG3_REG_12__SCAN_IN), .C2(keyinput_g46), .A(n9673), .ZN(n9676) );
  AOI22_X1 U12360 ( .A1(P3_DATAO_REG_27__SCAN_IN), .A2(keyinput_g69), .B1(
        P3_DATAO_REG_24__SCAN_IN), .B2(keyinput_g72), .ZN(n9674) );
  OAI221_X1 U12361 ( .B1(P3_DATAO_REG_27__SCAN_IN), .B2(keyinput_g69), .C1(
        P3_DATAO_REG_24__SCAN_IN), .C2(keyinput_g72), .A(n9674), .ZN(n9675) );
  NOR4_X1 U12362 ( .A1(n9678), .A2(n9677), .A3(n9676), .A4(n9675), .ZN(n9688)
         );
  AOI22_X1 U12363 ( .A1(P3_DATAO_REG_6__SCAN_IN), .A2(keyinput_g90), .B1(
        P3_REG3_REG_7__SCAN_IN), .B2(keyinput_g35), .ZN(n9679) );
  OAI221_X1 U12364 ( .B1(P3_DATAO_REG_6__SCAN_IN), .B2(keyinput_g90), .C1(
        P3_REG3_REG_7__SCAN_IN), .C2(keyinput_g35), .A(n9679), .ZN(n9686) );
  AOI22_X1 U12365 ( .A1(P3_DATAO_REG_14__SCAN_IN), .A2(keyinput_g82), .B1(
        SI_11_), .B2(keyinput_g21), .ZN(n9680) );
  OAI221_X1 U12366 ( .B1(P3_DATAO_REG_14__SCAN_IN), .B2(keyinput_g82), .C1(
        SI_11_), .C2(keyinput_g21), .A(n9680), .ZN(n9685) );
  AOI22_X1 U12367 ( .A1(P3_DATAO_REG_12__SCAN_IN), .A2(keyinput_g84), .B1(
        P3_ADDR_REG_4__SCAN_IN), .B2(keyinput_g101), .ZN(n9681) );
  OAI221_X1 U12368 ( .B1(P3_DATAO_REG_12__SCAN_IN), .B2(keyinput_g84), .C1(
        P3_ADDR_REG_4__SCAN_IN), .C2(keyinput_g101), .A(n9681), .ZN(n9684) );
  AOI22_X1 U12369 ( .A1(P3_DATAO_REG_9__SCAN_IN), .A2(keyinput_g87), .B1(
        P3_DATAO_REG_29__SCAN_IN), .B2(keyinput_g67), .ZN(n9682) );
  OAI221_X1 U12370 ( .B1(P3_DATAO_REG_9__SCAN_IN), .B2(keyinput_g87), .C1(
        P3_DATAO_REG_29__SCAN_IN), .C2(keyinput_g67), .A(n9682), .ZN(n9683) );
  NOR4_X1 U12371 ( .A1(n9686), .A2(n9685), .A3(n9684), .A4(n9683), .ZN(n9687)
         );
  NAND4_X1 U12372 ( .A1(n9690), .A2(n9689), .A3(n9688), .A4(n9687), .ZN(n9825)
         );
  AOI22_X1 U12373 ( .A1(P3_DATAO_REG_21__SCAN_IN), .A2(keyinput_g75), .B1(
        P3_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .ZN(n9691) );
  OAI221_X1 U12374 ( .B1(P3_DATAO_REG_21__SCAN_IN), .B2(keyinput_g75), .C1(
        P3_REG3_REG_15__SCAN_IN), .C2(keyinput_g63), .A(n9691), .ZN(n9698) );
  AOI22_X1 U12375 ( .A1(P3_DATAO_REG_0__SCAN_IN), .A2(keyinput_g96), .B1(
        SI_21_), .B2(keyinput_g11), .ZN(n9692) );
  OAI221_X1 U12376 ( .B1(P3_DATAO_REG_0__SCAN_IN), .B2(keyinput_g96), .C1(
        SI_21_), .C2(keyinput_g11), .A(n9692), .ZN(n9697) );
  AOI22_X1 U12377 ( .A1(SI_25_), .A2(keyinput_g7), .B1(P3_STATE_REG_SCAN_IN), 
        .B2(keyinput_g34), .ZN(n9693) );
  OAI221_X1 U12378 ( .B1(SI_25_), .B2(keyinput_g7), .C1(P3_STATE_REG_SCAN_IN), 
        .C2(keyinput_g34), .A(n9693), .ZN(n9696) );
  AOI22_X1 U12379 ( .A1(P3_DATAO_REG_17__SCAN_IN), .A2(keyinput_g79), .B1(
        P3_DATAO_REG_3__SCAN_IN), .B2(keyinput_g93), .ZN(n9694) );
  OAI221_X1 U12380 ( .B1(P3_DATAO_REG_17__SCAN_IN), .B2(keyinput_g79), .C1(
        P3_DATAO_REG_3__SCAN_IN), .C2(keyinput_g93), .A(n9694), .ZN(n9695) );
  NOR4_X1 U12381 ( .A1(n9698), .A2(n9697), .A3(n9696), .A4(n9695), .ZN(n9728)
         );
  AOI22_X1 U12382 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(keyinput_g98), .B1(
        P3_DATAO_REG_1__SCAN_IN), .B2(keyinput_g95), .ZN(n9699) );
  OAI221_X1 U12383 ( .B1(P3_ADDR_REG_1__SCAN_IN), .B2(keyinput_g98), .C1(
        P3_DATAO_REG_1__SCAN_IN), .C2(keyinput_g95), .A(n9699), .ZN(n9706) );
  AOI22_X1 U12384 ( .A1(P3_DATAO_REG_10__SCAN_IN), .A2(keyinput_g86), .B1(
        P3_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .ZN(n9700) );
  OAI221_X1 U12385 ( .B1(P3_DATAO_REG_10__SCAN_IN), .B2(keyinput_g86), .C1(
        P3_REG3_REG_22__SCAN_IN), .C2(keyinput_g57), .A(n9700), .ZN(n9705) );
  AOI22_X1 U12386 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(keyinput_g119), .B1(
        P3_REG3_REG_23__SCAN_IN), .B2(keyinput_g38), .ZN(n9701) );
  OAI221_X1 U12387 ( .B1(P1_IR_REG_12__SCAN_IN), .B2(keyinput_g119), .C1(
        P3_REG3_REG_23__SCAN_IN), .C2(keyinput_g38), .A(n9701), .ZN(n9704) );
  AOI22_X1 U12388 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(keyinput_g125), .B1(
        P3_REG3_REG_6__SCAN_IN), .B2(keyinput_g61), .ZN(n9702) );
  OAI221_X1 U12389 ( .B1(P1_IR_REG_18__SCAN_IN), .B2(keyinput_g125), .C1(
        P3_REG3_REG_6__SCAN_IN), .C2(keyinput_g61), .A(n9702), .ZN(n9703) );
  NOR4_X1 U12390 ( .A1(n9706), .A2(n9705), .A3(n9704), .A4(n9703), .ZN(n9727)
         );
  AOI22_X1 U12391 ( .A1(P3_DATAO_REG_8__SCAN_IN), .A2(keyinput_g88), .B1(
        P3_DATAO_REG_25__SCAN_IN), .B2(keyinput_g71), .ZN(n9707) );
  OAI221_X1 U12392 ( .B1(P3_DATAO_REG_8__SCAN_IN), .B2(keyinput_g88), .C1(
        P3_DATAO_REG_25__SCAN_IN), .C2(keyinput_g71), .A(n9707), .ZN(n9714) );
  AOI22_X1 U12393 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(keyinput_g102), .B1(
        SI_29_), .B2(keyinput_g3), .ZN(n9708) );
  OAI221_X1 U12394 ( .B1(P3_ADDR_REG_5__SCAN_IN), .B2(keyinput_g102), .C1(
        SI_29_), .C2(keyinput_g3), .A(n9708), .ZN(n9713) );
  AOI22_X1 U12395 ( .A1(P3_REG3_REG_2__SCAN_IN), .A2(keyinput_g59), .B1(
        P3_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .ZN(n9709) );
  OAI221_X1 U12396 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .C1(
        P3_REG3_REG_19__SCAN_IN), .C2(keyinput_g41), .A(n9709), .ZN(n9712) );
  AOI22_X1 U12397 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(keyinput_g127), .B1(SI_10_), .B2(keyinput_g22), .ZN(n9710) );
  OAI221_X1 U12398 ( .B1(P1_IR_REG_20__SCAN_IN), .B2(keyinput_g127), .C1(
        SI_10_), .C2(keyinput_g22), .A(n9710), .ZN(n9711) );
  NOR4_X1 U12399 ( .A1(n9714), .A2(n9713), .A3(n9712), .A4(n9711), .ZN(n9726)
         );
  AOI22_X1 U12400 ( .A1(n11576), .A2(keyinput_g52), .B1(keyinput_g103), .B2(
        n9716), .ZN(n9715) );
  OAI221_X1 U12401 ( .B1(n11576), .B2(keyinput_g52), .C1(n9716), .C2(
        keyinput_g103), .A(n9715), .ZN(n9724) );
  AOI22_X1 U12402 ( .A1(n13441), .A2(keyinput_g48), .B1(keyinput_g92), .B2(
        n10758), .ZN(n9717) );
  OAI221_X1 U12403 ( .B1(n13441), .B2(keyinput_g48), .C1(n10758), .C2(
        keyinput_g92), .A(n9717), .ZN(n9723) );
  INV_X1 U12404 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n12266) );
  XOR2_X1 U12405 ( .A(n12266), .B(keyinput_g58), .Z(n9721) );
  XNOR2_X1 U12406 ( .A(SI_6_), .B(keyinput_g26), .ZN(n9720) );
  XNOR2_X1 U12407 ( .A(SI_2_), .B(keyinput_g30), .ZN(n9719) );
  XNOR2_X1 U12408 ( .A(P3_REG3_REG_14__SCAN_IN), .B(keyinput_g37), .ZN(n9718)
         );
  NAND4_X1 U12409 ( .A1(n9721), .A2(n9720), .A3(n9719), .A4(n9718), .ZN(n9722)
         );
  NOR3_X1 U12410 ( .A1(n9724), .A2(n9723), .A3(n9722), .ZN(n9725) );
  NAND4_X1 U12411 ( .A1(n9728), .A2(n9727), .A3(n9726), .A4(n9725), .ZN(n9824)
         );
  INV_X1 U12412 ( .A(SI_31_), .ZN(n14044) );
  AOI22_X1 U12413 ( .A1(n14044), .A2(keyinput_g1), .B1(keyinput_g94), .B2(
        n10718), .ZN(n9729) );
  OAI221_X1 U12414 ( .B1(n14044), .B2(keyinput_g1), .C1(n10718), .C2(
        keyinput_g94), .A(n9729), .ZN(n9739) );
  AOI22_X1 U12415 ( .A1(n9207), .A2(keyinput_g47), .B1(keyinput_g40), .B2(
        n11284), .ZN(n9730) );
  OAI221_X1 U12416 ( .B1(n9207), .B2(keyinput_g47), .C1(n11284), .C2(
        keyinput_g40), .A(n9730), .ZN(n9738) );
  AOI22_X1 U12417 ( .A1(n9733), .A2(keyinput_g118), .B1(keyinput_g116), .B2(
        n9732), .ZN(n9731) );
  OAI221_X1 U12418 ( .B1(n9733), .B2(keyinput_g118), .C1(n9732), .C2(
        keyinput_g116), .A(n9731), .ZN(n9737) );
  XNOR2_X1 U12419 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_g113), .ZN(n9735) );
  XNOR2_X1 U12420 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_g108), .ZN(n9734) );
  NAND2_X1 U12421 ( .A1(n9735), .A2(n9734), .ZN(n9736) );
  NOR4_X1 U12422 ( .A1(n9739), .A2(n9738), .A3(n9737), .A4(n9736), .ZN(n9775)
         );
  INV_X1 U12423 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n9741) );
  AOI22_X1 U12424 ( .A1(n9741), .A2(keyinput_g60), .B1(keyinput_g54), .B2(
        n11367), .ZN(n9740) );
  OAI221_X1 U12425 ( .B1(n9741), .B2(keyinput_g60), .C1(n11367), .C2(
        keyinput_g54), .A(n9740), .ZN(n9750) );
  INV_X1 U12426 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n11015) );
  AOI22_X1 U12427 ( .A1(n11219), .A2(keyinput_g97), .B1(keyinput_g73), .B2(
        n11015), .ZN(n9742) );
  OAI221_X1 U12428 ( .B1(n11219), .B2(keyinput_g97), .C1(n11015), .C2(
        keyinput_g73), .A(n9742), .ZN(n9749) );
  AOI22_X1 U12429 ( .A1(n8862), .A2(keyinput_g49), .B1(keyinput_g115), .B2(
        n9744), .ZN(n9743) );
  OAI221_X1 U12430 ( .B1(n8862), .B2(keyinput_g49), .C1(n9744), .C2(
        keyinput_g115), .A(n9743), .ZN(n9748) );
  XNOR2_X1 U12431 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_g120), .ZN(n9746)
         );
  XNOR2_X1 U12432 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_g110), .ZN(n9745) );
  NAND2_X1 U12433 ( .A1(n9746), .A2(n9745), .ZN(n9747) );
  NOR4_X1 U12434 ( .A1(n9750), .A2(n9749), .A3(n9748), .A4(n9747), .ZN(n9774)
         );
  INV_X1 U12435 ( .A(P3_DATAO_REG_18__SCAN_IN), .ZN(n10762) );
  AOI22_X1 U12436 ( .A1(n10762), .A2(keyinput_g78), .B1(keyinput_g89), .B2(
        n10767), .ZN(n9751) );
  OAI221_X1 U12437 ( .B1(n10762), .B2(keyinput_g78), .C1(n10767), .C2(
        keyinput_g89), .A(n9751), .ZN(n9760) );
  AOI22_X1 U12438 ( .A1(n8931), .A2(keyinput_g53), .B1(keyinput_g124), .B2(
        n9753), .ZN(n9752) );
  OAI221_X1 U12439 ( .B1(n8931), .B2(keyinput_g53), .C1(n9753), .C2(
        keyinput_g124), .A(n9752), .ZN(n9759) );
  AOI22_X1 U12440 ( .A1(n13367), .A2(keyinput_g42), .B1(keyinput_g43), .B2(
        n12129), .ZN(n9754) );
  OAI221_X1 U12441 ( .B1(n13367), .B2(keyinput_g42), .C1(n12129), .C2(
        keyinput_g43), .A(n9754), .ZN(n9758) );
  XNOR2_X1 U12442 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_g121), .ZN(n9756)
         );
  XNOR2_X1 U12443 ( .A(P3_REG3_REG_17__SCAN_IN), .B(keyinput_g50), .ZN(n9755)
         );
  NAND2_X1 U12444 ( .A1(n9756), .A2(n9755), .ZN(n9757) );
  NOR4_X1 U12445 ( .A1(n9760), .A2(n9759), .A3(n9758), .A4(n9757), .ZN(n9773)
         );
  INV_X1 U12446 ( .A(P3_B_REG_SCAN_IN), .ZN(n9762) );
  AOI22_X1 U12447 ( .A1(n9762), .A2(keyinput_g64), .B1(keyinput_g8), .B2(
        n11937), .ZN(n9761) );
  OAI221_X1 U12448 ( .B1(n9762), .B2(keyinput_g64), .C1(n11937), .C2(
        keyinput_g8), .A(n9761), .ZN(n9771) );
  XOR2_X1 U12449 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_g122), .Z(n9770) );
  XNOR2_X1 U12450 ( .A(n9763), .B(keyinput_g114), .ZN(n9769) );
  XNOR2_X1 U12451 ( .A(SI_9_), .B(keyinput_g23), .ZN(n9767) );
  XNOR2_X1 U12452 ( .A(SI_19_), .B(keyinput_g13), .ZN(n9766) );
  XNOR2_X1 U12453 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_g109), .ZN(n9765) );
  XNOR2_X1 U12454 ( .A(SI_22_), .B(keyinput_g10), .ZN(n9764) );
  NAND4_X1 U12455 ( .A1(n9767), .A2(n9766), .A3(n9765), .A4(n9764), .ZN(n9768)
         );
  NOR4_X1 U12456 ( .A1(n9771), .A2(n9770), .A3(n9769), .A4(n9768), .ZN(n9772)
         );
  NAND4_X1 U12457 ( .A1(n9775), .A2(n9774), .A3(n9773), .A4(n9772), .ZN(n9823)
         );
  AOI22_X1 U12458 ( .A1(n12150), .A2(keyinput_g6), .B1(n11177), .B2(
        keyinput_g44), .ZN(n9776) );
  OAI221_X1 U12459 ( .B1(n12150), .B2(keyinput_g6), .C1(n11177), .C2(
        keyinput_g44), .A(n9776), .ZN(n9784) );
  INV_X1 U12460 ( .A(P3_DATAO_REG_19__SCAN_IN), .ZN(n10787) );
  AOI22_X1 U12461 ( .A1(n12851), .A2(keyinput_g4), .B1(keyinput_g77), .B2(
        n10787), .ZN(n9777) );
  OAI221_X1 U12462 ( .B1(n12851), .B2(keyinput_g4), .C1(n10787), .C2(
        keyinput_g77), .A(n9777), .ZN(n9783) );
  INV_X1 U12463 ( .A(P3_DATAO_REG_5__SCAN_IN), .ZN(n10742) );
  AOI22_X1 U12464 ( .A1(n10742), .A2(keyinput_g91), .B1(n10739), .B2(
        keyinput_g14), .ZN(n9778) );
  OAI221_X1 U12465 ( .B1(n10742), .B2(keyinput_g91), .C1(n10739), .C2(
        keyinput_g14), .A(n9778), .ZN(n9782) );
  XNOR2_X1 U12466 ( .A(SI_3_), .B(keyinput_g29), .ZN(n9780) );
  XNOR2_X1 U12467 ( .A(SI_20_), .B(keyinput_g12), .ZN(n9779) );
  NAND2_X1 U12468 ( .A1(n9780), .A2(n9779), .ZN(n9781) );
  NOR4_X1 U12469 ( .A1(n9784), .A2(n9783), .A3(n9782), .A4(n9781), .ZN(n9821)
         );
  INV_X1 U12470 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n9786) );
  INV_X1 U12471 ( .A(P3_RD_REG_SCAN_IN), .ZN(n10376) );
  AOI22_X1 U12472 ( .A1(n9786), .A2(keyinput_g51), .B1(keyinput_g33), .B2(
        n10376), .ZN(n9785) );
  OAI221_X1 U12473 ( .B1(n9786), .B2(keyinput_g51), .C1(n10376), .C2(
        keyinput_g33), .A(n9785), .ZN(n9794) );
  AOI22_X1 U12474 ( .A1(n10804), .A2(keyinput_g76), .B1(n9150), .B2(
        keyinput_g45), .ZN(n9787) );
  OAI221_X1 U12475 ( .B1(n10804), .B2(keyinput_g76), .C1(n9150), .C2(
        keyinput_g45), .A(n9787), .ZN(n9793) );
  XNOR2_X1 U12476 ( .A(SI_13_), .B(keyinput_g19), .ZN(n9791) );
  XNOR2_X1 U12477 ( .A(SI_5_), .B(keyinput_g27), .ZN(n9790) );
  XNOR2_X1 U12478 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_g111), .ZN(n9789) );
  XNOR2_X1 U12479 ( .A(SI_7_), .B(keyinput_g25), .ZN(n9788) );
  NAND4_X1 U12480 ( .A1(n9791), .A2(n9790), .A3(n9789), .A4(n9788), .ZN(n9792)
         );
  NOR3_X1 U12481 ( .A1(n9794), .A2(n9793), .A3(n9792), .ZN(n9820) );
  AOI22_X1 U12482 ( .A1(n10760), .A2(keyinput_g83), .B1(keyinput_g100), .B2(
        n9796), .ZN(n9795) );
  OAI221_X1 U12483 ( .B1(n10760), .B2(keyinput_g83), .C1(n9796), .C2(
        keyinput_g100), .A(n9795), .ZN(n9804) );
  AOI22_X1 U12484 ( .A1(n10497), .A2(keyinput_g17), .B1(n13471), .B2(
        keyinput_g55), .ZN(n9797) );
  OAI221_X1 U12485 ( .B1(n10497), .B2(keyinput_g17), .C1(n13471), .C2(
        keyinput_g55), .A(n9797), .ZN(n9803) );
  XOR2_X1 U12486 ( .A(n9013), .B(keyinput_g56), .Z(n9801) );
  XNOR2_X1 U12487 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_g123), .ZN(n9800)
         );
  XNOR2_X1 U12488 ( .A(SI_27_), .B(keyinput_g5), .ZN(n9799) );
  XNOR2_X1 U12489 ( .A(SI_8_), .B(keyinput_g24), .ZN(n9798) );
  NAND4_X1 U12490 ( .A1(n9801), .A2(n9800), .A3(n9799), .A4(n9798), .ZN(n9802)
         );
  NOR3_X1 U12491 ( .A1(n9804), .A2(n9803), .A3(n9802), .ZN(n9819) );
  AOI22_X1 U12492 ( .A1(n10457), .A2(keyinput_g18), .B1(keyinput_g106), .B2(
        n9806), .ZN(n9805) );
  OAI221_X1 U12493 ( .B1(n10457), .B2(keyinput_g18), .C1(n9806), .C2(
        keyinput_g106), .A(n9805), .ZN(n9817) );
  AOI22_X1 U12494 ( .A1(n9809), .A2(keyinput_g105), .B1(keyinput_g0), .B2(
        n9808), .ZN(n9807) );
  OAI221_X1 U12495 ( .B1(n9809), .B2(keyinput_g105), .C1(n9808), .C2(
        keyinput_g0), .A(n9807), .ZN(n9816) );
  INV_X1 U12496 ( .A(SI_0_), .ZN(n9810) );
  XOR2_X1 U12497 ( .A(n9810), .B(keyinput_g32), .Z(n9814) );
  XNOR2_X1 U12498 ( .A(SI_1_), .B(keyinput_g31), .ZN(n9813) );
  XNOR2_X1 U12499 ( .A(P3_REG3_REG_27__SCAN_IN), .B(keyinput_g36), .ZN(n9812)
         );
  XNOR2_X1 U12500 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_g112), .ZN(n9811) );
  NAND4_X1 U12501 ( .A1(n9814), .A2(n9813), .A3(n9812), .A4(n9811), .ZN(n9815)
         );
  NOR3_X1 U12502 ( .A1(n9817), .A2(n9816), .A3(n9815), .ZN(n9818) );
  NAND4_X1 U12503 ( .A1(n9821), .A2(n9820), .A3(n9819), .A4(n9818), .ZN(n9822)
         );
  NOR4_X1 U12504 ( .A1(n9825), .A2(n9824), .A3(n9823), .A4(n9822), .ZN(n9826)
         );
  AOI211_X1 U12505 ( .C1(n9829), .C2(n9828), .A(n9827), .B(n9826), .ZN(n9830)
         );
  INV_X1 U12506 ( .A(n9830), .ZN(n9831) );
  INV_X1 U12507 ( .A(n15511), .ZN(n9835) );
  NAND2_X1 U12508 ( .A1(n9837), .A2(n15550), .ZN(n9842) );
  NAND2_X1 U12509 ( .A1(n15550), .A2(n15532), .ZN(n14472) );
  INV_X1 U12510 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9838) );
  OR2_X1 U12511 ( .A1(n15550), .A2(n9838), .ZN(n9839) );
  NAND2_X1 U12512 ( .A1(n9842), .A2(n9841), .ZN(P2_U3527) );
  NAND2_X1 U12513 ( .A1(n9844), .A2(n9843), .ZN(n9851) );
  OR2_X1 U12514 ( .A1(n9847), .A2(SI_28_), .ZN(n9848) );
  INV_X1 U12515 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n13375) );
  INV_X1 U12516 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14528) );
  MUX2_X1 U12517 ( .A(n13375), .B(n14528), .S(n6676), .Z(n10043) );
  XNOR2_X1 U12518 ( .A(n10043), .B(SI_29_), .ZN(n10041) );
  XNOR2_X2 U12519 ( .A(n10042), .B(n10041), .ZN(n13373) );
  NAND2_X1 U12520 ( .A1(n13373), .A2(n8325), .ZN(n9850) );
  OR2_X1 U12521 ( .A1(n10056), .A2(n14528), .ZN(n9849) );
  NAND2_X2 U12522 ( .A1(n9850), .A2(n9849), .ZN(n10063) );
  XNOR2_X1 U12523 ( .A(n10063), .B(n14150), .ZN(n10094) );
  XNOR2_X1 U12524 ( .A(n9853), .B(n10094), .ZN(n9854) );
  INV_X1 U12525 ( .A(n14228), .ZN(n10037) );
  OR2_X1 U12526 ( .A1(n10037), .A2(n14323), .ZN(n9862) );
  NAND2_X1 U12527 ( .A1(n9855), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n9859) );
  NAND2_X1 U12528 ( .A1(n8310), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9858) );
  NAND2_X1 U12529 ( .A1(n9856), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9857) );
  NAND3_X1 U12530 ( .A1(n9859), .A2(n9858), .A3(n9857), .ZN(n14149) );
  INV_X1 U12531 ( .A(n14149), .ZN(n9861) );
  INV_X1 U12532 ( .A(n12477), .ZN(n10540) );
  NAND2_X1 U12533 ( .A1(n10540), .A2(P2_B_REG_SCAN_IN), .ZN(n9860) );
  NAND2_X1 U12534 ( .A1(n14369), .A2(n9860), .ZN(n14204) );
  AND2_X1 U12535 ( .A1(n9862), .A2(n7594), .ZN(n9863) );
  INV_X1 U12536 ( .A(n14222), .ZN(n9867) );
  AOI211_X1 U12537 ( .C1(n10063), .C2(n6999), .A(n12878), .B(n14210), .ZN(
        n14216) );
  INV_X1 U12538 ( .A(n14216), .ZN(n9866) );
  NAND2_X1 U12539 ( .A1(n9867), .A2(n9866), .ZN(n9868) );
  INV_X1 U12540 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9869) );
  OR2_X1 U12541 ( .A1(n15550), .A2(n9869), .ZN(n9870) );
  OAI21_X1 U12542 ( .B1(n10164), .B2(n15548), .A(n7580), .ZN(P2_U3528) );
  INV_X1 U12543 ( .A(n14415), .ZN(n14235) );
  BUF_X4 U12544 ( .A(n9876), .Z(n10102) );
  MUX2_X1 U12545 ( .A(n14141), .B(n14235), .S(n10102), .Z(n10036) );
  INV_X1 U12546 ( .A(n10036), .ZN(n10067) );
  NAND2_X1 U12547 ( .A1(n10576), .A2(n9876), .ZN(n9871) );
  NAND2_X1 U12548 ( .A1(n9871), .A2(n10550), .ZN(n9873) );
  NAND2_X1 U12549 ( .A1(n10236), .A2(n9876), .ZN(n9872) );
  NAND2_X1 U12550 ( .A1(n9873), .A2(n9872), .ZN(n9875) );
  NAND3_X1 U12551 ( .A1(n10550), .A2(n10710), .A3(n14434), .ZN(n9874) );
  NAND2_X1 U12552 ( .A1(n9875), .A2(n9874), .ZN(n9879) );
  MUX2_X1 U12553 ( .A(n14170), .B(n10753), .S(n9876), .Z(n9880) );
  NAND2_X1 U12554 ( .A1(n9879), .A2(n9880), .ZN(n9878) );
  MUX2_X1 U12555 ( .A(n14170), .B(n10753), .S(n10061), .Z(n9877) );
  NAND2_X1 U12556 ( .A1(n9878), .A2(n9877), .ZN(n9884) );
  INV_X1 U12557 ( .A(n9879), .ZN(n9882) );
  NAND2_X1 U12558 ( .A1(n9882), .A2(n9881), .ZN(n9883) );
  NAND2_X1 U12559 ( .A1(n9884), .A2(n9883), .ZN(n9888) );
  MUX2_X1 U12560 ( .A(n14169), .B(n10812), .S(n10061), .Z(n9887) );
  NAND2_X1 U12561 ( .A1(n9888), .A2(n9887), .ZN(n9886) );
  MUX2_X1 U12562 ( .A(n14169), .B(n10812), .S(n10102), .Z(n9885) );
  NAND2_X1 U12563 ( .A1(n9886), .A2(n9885), .ZN(n9890) );
  MUX2_X1 U12564 ( .A(n14167), .B(n10905), .S(n10102), .Z(n9892) );
  MUX2_X1 U12565 ( .A(n14167), .B(n10905), .S(n10061), .Z(n9891) );
  INV_X1 U12566 ( .A(n9892), .ZN(n9893) );
  MUX2_X1 U12567 ( .A(n14166), .B(n11019), .S(n10104), .Z(n9896) );
  NAND2_X1 U12568 ( .A1(n9897), .A2(n9896), .ZN(n9895) );
  MUX2_X1 U12569 ( .A(n14166), .B(n11019), .S(n10102), .Z(n9894) );
  NAND2_X1 U12570 ( .A1(n9895), .A2(n9894), .ZN(n9899) );
  NAND2_X1 U12571 ( .A1(n9899), .A2(n9898), .ZN(n9902) );
  MUX2_X1 U12572 ( .A(n14165), .B(n11074), .S(n10102), .Z(n9903) );
  NAND2_X1 U12573 ( .A1(n9902), .A2(n9903), .ZN(n9901) );
  MUX2_X1 U12574 ( .A(n14165), .B(n11074), .S(n9993), .Z(n9900) );
  NAND2_X1 U12575 ( .A1(n9901), .A2(n9900), .ZN(n9907) );
  INV_X1 U12576 ( .A(n9902), .ZN(n9905) );
  INV_X1 U12577 ( .A(n9903), .ZN(n9904) );
  NAND2_X1 U12578 ( .A1(n9905), .A2(n9904), .ZN(n9906) );
  NAND2_X1 U12579 ( .A1(n9907), .A2(n9906), .ZN(n9910) );
  INV_X1 U12580 ( .A(n10102), .ZN(n9993) );
  MUX2_X1 U12581 ( .A(n14164), .B(n11685), .S(n9993), .Z(n9911) );
  NAND2_X1 U12582 ( .A1(n9910), .A2(n9911), .ZN(n9909) );
  MUX2_X1 U12583 ( .A(n14164), .B(n11685), .S(n10102), .Z(n9908) );
  INV_X1 U12584 ( .A(n9910), .ZN(n9913) );
  INV_X1 U12585 ( .A(n9911), .ZN(n9912) );
  NAND2_X1 U12586 ( .A1(n9913), .A2(n9912), .ZN(n9914) );
  MUX2_X1 U12587 ( .A(n14163), .B(n11088), .S(n10102), .Z(n9916) );
  INV_X1 U12588 ( .A(n10102), .ZN(n10104) );
  MUX2_X1 U12589 ( .A(n14163), .B(n11088), .S(n9993), .Z(n9915) );
  MUX2_X1 U12590 ( .A(n14162), .B(n15523), .S(n9993), .Z(n9920) );
  NAND2_X1 U12591 ( .A1(n9919), .A2(n9920), .ZN(n9918) );
  MUX2_X1 U12592 ( .A(n14162), .B(n15523), .S(n10102), .Z(n9917) );
  NAND2_X1 U12593 ( .A1(n9918), .A2(n9917), .ZN(n9924) );
  INV_X1 U12594 ( .A(n9919), .ZN(n9922) );
  INV_X1 U12595 ( .A(n9920), .ZN(n9921) );
  NAND2_X1 U12596 ( .A1(n9922), .A2(n9921), .ZN(n9923) );
  MUX2_X1 U12597 ( .A(n14161), .B(n11995), .S(n10102), .Z(n9926) );
  MUX2_X1 U12598 ( .A(n14161), .B(n11995), .S(n9993), .Z(n9925) );
  INV_X1 U12599 ( .A(n9926), .ZN(n9927) );
  MUX2_X1 U12600 ( .A(n14160), .B(n15533), .S(n9993), .Z(n9931) );
  NAND2_X1 U12601 ( .A1(n9930), .A2(n9931), .ZN(n9929) );
  MUX2_X1 U12602 ( .A(n14160), .B(n15533), .S(n10102), .Z(n9928) );
  NAND2_X1 U12603 ( .A1(n9929), .A2(n9928), .ZN(n9935) );
  INV_X1 U12604 ( .A(n9930), .ZN(n9933) );
  INV_X1 U12605 ( .A(n9931), .ZN(n9932) );
  NAND2_X1 U12606 ( .A1(n9933), .A2(n9932), .ZN(n9934) );
  MUX2_X1 U12607 ( .A(n14159), .B(n12257), .S(n10102), .Z(n9937) );
  MUX2_X1 U12608 ( .A(n14159), .B(n12257), .S(n9993), .Z(n9936) );
  INV_X1 U12609 ( .A(n9937), .ZN(n9938) );
  MUX2_X1 U12610 ( .A(n14158), .B(n12051), .S(n9993), .Z(n9942) );
  NAND2_X1 U12611 ( .A1(n9941), .A2(n9942), .ZN(n9940) );
  MUX2_X1 U12612 ( .A(n14158), .B(n12051), .S(n10102), .Z(n9939) );
  NAND2_X1 U12613 ( .A1(n9940), .A2(n9939), .ZN(n9946) );
  INV_X1 U12614 ( .A(n9941), .ZN(n9944) );
  INV_X1 U12615 ( .A(n9942), .ZN(n9943) );
  NAND2_X1 U12616 ( .A1(n9944), .A2(n9943), .ZN(n9945) );
  MUX2_X1 U12617 ( .A(n14157), .B(n12080), .S(n10102), .Z(n9948) );
  MUX2_X1 U12618 ( .A(n14157), .B(n12080), .S(n9993), .Z(n9947) );
  INV_X1 U12619 ( .A(n9948), .ZN(n9949) );
  INV_X1 U12620 ( .A(n12321), .ZN(n12363) );
  MUX2_X1 U12621 ( .A(n12406), .B(n12363), .S(n9993), .Z(n9961) );
  MUX2_X1 U12622 ( .A(n14156), .B(n12321), .S(n10102), .Z(n9960) );
  MUX2_X1 U12623 ( .A(n12485), .B(n8711), .S(n9993), .Z(n9969) );
  MUX2_X1 U12624 ( .A(n14155), .B(n12409), .S(n10102), .Z(n9968) );
  NAND2_X1 U12625 ( .A1(n9969), .A2(n9968), .ZN(n9957) );
  MUX2_X1 U12626 ( .A(n14154), .B(n14475), .S(n9993), .Z(n9974) );
  NAND2_X1 U12627 ( .A1(n9974), .A2(n14153), .ZN(n9950) );
  NAND2_X1 U12628 ( .A1(n12405), .A2(n9993), .ZN(n9952) );
  AOI21_X1 U12629 ( .B1(n9950), .B2(n9952), .A(n14518), .ZN(n9956) );
  NAND2_X1 U12630 ( .A1(n9974), .A2(n14129), .ZN(n9951) );
  OR2_X1 U12631 ( .A1(n14475), .A2(n9993), .ZN(n9962) );
  AOI21_X1 U12632 ( .B1(n9951), .B2(n9962), .A(n12565), .ZN(n9955) );
  NAND2_X1 U12633 ( .A1(n14153), .A2(n10102), .ZN(n9964) );
  OR2_X1 U12634 ( .A1(n14475), .A2(n9964), .ZN(n9954) );
  INV_X1 U12635 ( .A(n9952), .ZN(n9973) );
  NAND2_X1 U12636 ( .A1(n9973), .A2(n14129), .ZN(n9953) );
  NAND2_X1 U12637 ( .A1(n9954), .A2(n9953), .ZN(n9966) );
  OR3_X1 U12638 ( .A1(n9956), .A2(n9955), .A3(n9966), .ZN(n9972) );
  NAND2_X1 U12639 ( .A1(n9959), .A2(n9958), .ZN(n9982) );
  OR3_X1 U12640 ( .A1(n6717), .A2(n9961), .A3(n9960), .ZN(n9980) );
  INV_X1 U12641 ( .A(n9962), .ZN(n9963) );
  NAND2_X1 U12642 ( .A1(n9974), .A2(n9963), .ZN(n9965) );
  NAND2_X1 U12643 ( .A1(n9965), .A2(n9964), .ZN(n9967) );
  AOI22_X1 U12644 ( .A1(n9967), .A2(n14518), .B1(n9974), .B2(n9966), .ZN(n9979) );
  INV_X1 U12645 ( .A(n9968), .ZN(n9971) );
  INV_X1 U12646 ( .A(n9969), .ZN(n9970) );
  NAND3_X1 U12647 ( .A1(n9972), .A2(n9971), .A3(n9970), .ZN(n9978) );
  NAND2_X1 U12648 ( .A1(n9974), .A2(n9973), .ZN(n9975) );
  OAI21_X1 U12649 ( .B1(n10102), .B2(n14153), .A(n9975), .ZN(n9976) );
  NAND2_X1 U12650 ( .A1(n9976), .A2(n12565), .ZN(n9977) );
  AND4_X1 U12651 ( .A1(n9980), .A2(n9979), .A3(n9978), .A4(n9977), .ZN(n9981)
         );
  NAND2_X1 U12652 ( .A1(n9982), .A2(n9981), .ZN(n9985) );
  MUX2_X1 U12653 ( .A(n14367), .B(n14390), .S(n9993), .Z(n9986) );
  NAND2_X1 U12654 ( .A1(n9985), .A2(n9986), .ZN(n9984) );
  MUX2_X1 U12655 ( .A(n14367), .B(n14390), .S(n10102), .Z(n9983) );
  NAND2_X1 U12656 ( .A1(n9984), .A2(n9983), .ZN(n9990) );
  INV_X1 U12657 ( .A(n9985), .ZN(n9988) );
  INV_X1 U12658 ( .A(n9986), .ZN(n9987) );
  NAND2_X1 U12659 ( .A1(n9988), .A2(n9987), .ZN(n9989) );
  MUX2_X1 U12660 ( .A(n14356), .B(n14375), .S(n10102), .Z(n9992) );
  MUX2_X1 U12661 ( .A(n14356), .B(n14375), .S(n9993), .Z(n9991) );
  MUX2_X1 U12662 ( .A(n14370), .B(n14454), .S(n10104), .Z(n9997) );
  NAND2_X1 U12663 ( .A1(n9996), .A2(n9997), .ZN(n9995) );
  MUX2_X1 U12664 ( .A(n14370), .B(n14454), .S(n10102), .Z(n9994) );
  NAND2_X1 U12665 ( .A1(n9995), .A2(n9994), .ZN(n10001) );
  INV_X1 U12666 ( .A(n9996), .ZN(n9999) );
  INV_X1 U12667 ( .A(n9997), .ZN(n9998) );
  NAND2_X1 U12668 ( .A1(n9999), .A2(n9998), .ZN(n10000) );
  NAND2_X1 U12669 ( .A1(n10001), .A2(n10000), .ZN(n10004) );
  MUX2_X1 U12670 ( .A(n14355), .B(n14338), .S(n10102), .Z(n10005) );
  NAND2_X1 U12671 ( .A1(n10004), .A2(n10005), .ZN(n10003) );
  MUX2_X1 U12672 ( .A(n14355), .B(n14338), .S(n10104), .Z(n10002) );
  NAND2_X1 U12673 ( .A1(n10003), .A2(n10002), .ZN(n10009) );
  INV_X1 U12674 ( .A(n10004), .ZN(n10007) );
  INV_X1 U12675 ( .A(n10005), .ZN(n10006) );
  NAND2_X1 U12676 ( .A1(n10007), .A2(n10006), .ZN(n10008) );
  NAND2_X1 U12677 ( .A1(n10009), .A2(n10008), .ZN(n10012) );
  MUX2_X1 U12678 ( .A(n14335), .B(n14443), .S(n9993), .Z(n10011) );
  MUX2_X1 U12679 ( .A(n14335), .B(n14443), .S(n10102), .Z(n10010) );
  MUX2_X1 U12680 ( .A(n14152), .B(n14306), .S(n10102), .Z(n10016) );
  MUX2_X1 U12681 ( .A(n14152), .B(n14306), .S(n9993), .Z(n10013) );
  NAND2_X1 U12682 ( .A1(n10014), .A2(n10013), .ZN(n10019) );
  INV_X1 U12683 ( .A(n10015), .ZN(n10017) );
  NAND2_X1 U12684 ( .A1(n10017), .A2(n7467), .ZN(n10018) );
  NAND2_X1 U12685 ( .A1(n10019), .A2(n10018), .ZN(n10021) );
  MUX2_X1 U12686 ( .A(n14151), .B(n14430), .S(n10104), .Z(n10022) );
  MUX2_X1 U12687 ( .A(n14151), .B(n14430), .S(n10102), .Z(n10020) );
  INV_X1 U12688 ( .A(n10022), .ZN(n10023) );
  MUX2_X1 U12689 ( .A(n14254), .B(n14085), .S(n10102), .Z(n10027) );
  MUX2_X1 U12690 ( .A(n14254), .B(n14085), .S(n9993), .Z(n10024) );
  NAND2_X1 U12691 ( .A1(n10025), .A2(n10024), .ZN(n10031) );
  INV_X1 U12692 ( .A(n10026), .ZN(n10029) );
  INV_X1 U12693 ( .A(n10027), .ZN(n10028) );
  NAND2_X1 U12694 ( .A1(n10029), .A2(n10028), .ZN(n10030) );
  MUX2_X1 U12695 ( .A(n14229), .B(n14420), .S(n9993), .Z(n10032) );
  MUX2_X1 U12696 ( .A(n14229), .B(n14420), .S(n10102), .Z(n10034) );
  INV_X1 U12697 ( .A(n10032), .ZN(n10033) );
  MUX2_X1 U12698 ( .A(n14255), .B(n14415), .S(n9993), .Z(n10035) );
  MUX2_X1 U12699 ( .A(n10037), .B(n12853), .S(n10102), .Z(n10115) );
  MUX2_X1 U12700 ( .A(n14228), .B(n12892), .S(n10104), .Z(n10114) );
  NAND2_X1 U12701 ( .A1(n8314), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n10040) );
  NAND2_X1 U12702 ( .A1(n8310), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n10039) );
  NAND2_X1 U12703 ( .A1(n9856), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n10038) );
  NAND3_X1 U12704 ( .A1(n10040), .A2(n10039), .A3(n10038), .ZN(n14206) );
  NAND2_X1 U12705 ( .A1(n14206), .A2(n10102), .ZN(n10059) );
  MUX2_X1 U12706 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n10046), .Z(n10044) );
  XNOR2_X1 U12707 ( .A(n10044), .B(SI_30_), .ZN(n10053) );
  INV_X1 U12708 ( .A(n10044), .ZN(n10045) );
  MUX2_X1 U12709 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n6676), .Z(n10047) );
  XNOR2_X1 U12710 ( .A(n10047), .B(SI_31_), .ZN(n10048) );
  NAND2_X1 U12711 ( .A1(n14521), .A2(n8325), .ZN(n10052) );
  INV_X1 U12712 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n10050) );
  OR2_X1 U12713 ( .A1(n10056), .A2(n10050), .ZN(n10051) );
  MUX2_X1 U12714 ( .A(n10059), .B(n14206), .S(n14484), .Z(n10065) );
  INV_X1 U12715 ( .A(n10053), .ZN(n10054) );
  NAND2_X1 U12716 ( .A1(n12960), .A2(n8325), .ZN(n10058) );
  INV_X1 U12717 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13139) );
  OR2_X1 U12718 ( .A1(n10056), .A2(n13139), .ZN(n10057) );
  NAND2_X1 U12719 ( .A1(n8741), .A2(n10142), .ZN(n10108) );
  NAND4_X1 U12720 ( .A1(n10059), .A2(n10098), .A3(n10141), .A4(n10108), .ZN(
        n10060) );
  AOI22_X1 U12721 ( .A1(n14202), .A2(n10104), .B1(n14149), .B2(n10060), .ZN(
        n10125) );
  MUX2_X1 U12722 ( .A(n14149), .B(n14202), .S(n10102), .Z(n10124) );
  INV_X1 U12723 ( .A(n14150), .ZN(n10062) );
  MUX2_X1 U12724 ( .A(n10062), .B(n14220), .S(n10104), .Z(n10119) );
  MUX2_X1 U12725 ( .A(n14150), .B(n10063), .S(n10102), .Z(n10118) );
  OAI22_X1 U12726 ( .A1(n10125), .A2(n10124), .B1(n10119), .B2(n10118), .ZN(
        n10064) );
  AND2_X1 U12727 ( .A1(n10065), .A2(n10064), .ZN(n10112) );
  AOI21_X1 U12728 ( .B1(n10115), .B2(n10114), .A(n10112), .ZN(n10066) );
  INV_X1 U12729 ( .A(n14206), .ZN(n10103) );
  XNOR2_X1 U12730 ( .A(n14484), .B(n10103), .ZN(n10113) );
  XOR2_X1 U12731 ( .A(n14149), .B(n14202), .Z(n10096) );
  NAND2_X1 U12732 ( .A1(n10069), .A2(n10068), .ZN(n12315) );
  NAND2_X1 U12733 ( .A1(n10071), .A2(n10070), .ZN(n12075) );
  NAND2_X1 U12734 ( .A1(n10073), .A2(n10072), .ZN(n12041) );
  AND2_X1 U12735 ( .A1(n10550), .A2(n10235), .ZN(n10716) );
  NAND4_X1 U12736 ( .A1(n10749), .A2(n10077), .A3(n10716), .A4(n10076), .ZN(
        n10078) );
  NOR3_X1 U12737 ( .A1(n10078), .A2(n10999), .A3(n10851), .ZN(n10079) );
  NAND4_X1 U12738 ( .A1(n11269), .A2(n10079), .A3(n11317), .A4(n11070), .ZN(
        n10080) );
  OR3_X1 U12739 ( .A1(n11731), .A2(n10081), .A3(n10080), .ZN(n10082) );
  NOR2_X1 U12740 ( .A1(n10083), .A2(n10082), .ZN(n10084) );
  NAND3_X1 U12741 ( .A1(n12315), .A2(n10085), .A3(n12482), .ZN(n10086) );
  OR3_X1 U12742 ( .A1(n12374), .A2(n12561), .A3(n10086), .ZN(n10087) );
  NOR2_X1 U12743 ( .A1(n14283), .A2(n10089), .ZN(n10091) );
  NAND4_X1 U12744 ( .A1(n10094), .A2(n10093), .A3(n10092), .A4(n14238), .ZN(
        n10095) );
  NOR3_X1 U12745 ( .A1(n10113), .A2(n10096), .A3(n10095), .ZN(n10097) );
  XNOR2_X1 U12746 ( .A(n10097), .B(n11007), .ZN(n10099) );
  NOR2_X1 U12747 ( .A1(n10099), .A2(n10098), .ZN(n10109) );
  INV_X1 U12748 ( .A(n8741), .ZN(n10101) );
  OAI22_X1 U12749 ( .A1(n11007), .A2(n8697), .B1(n7213), .B2(n10142), .ZN(
        n10100) );
  OR3_X1 U12750 ( .A1(n14484), .A2(n10103), .A3(n10102), .ZN(n10107) );
  NOR2_X1 U12751 ( .A1(n14206), .A2(n10104), .ZN(n10105) );
  NAND2_X1 U12752 ( .A1(n14484), .A2(n10105), .ZN(n10106) );
  NAND2_X1 U12753 ( .A1(n10107), .A2(n10106), .ZN(n10130) );
  NOR3_X1 U12754 ( .A1(n10129), .A2(n10135), .A3(n10130), .ZN(n10140) );
  INV_X1 U12755 ( .A(n10108), .ZN(n10110) );
  INV_X1 U12756 ( .A(n10112), .ZN(n10123) );
  INV_X1 U12757 ( .A(n10113), .ZN(n10121) );
  INV_X1 U12758 ( .A(n10114), .ZN(n10117) );
  INV_X1 U12759 ( .A(n10115), .ZN(n10116) );
  AOI22_X1 U12760 ( .A1(n10119), .A2(n10118), .B1(n10117), .B2(n10116), .ZN(
        n10120) );
  NAND2_X1 U12761 ( .A1(n10121), .A2(n10120), .ZN(n10122) );
  NAND2_X1 U12762 ( .A1(n10123), .A2(n10122), .ZN(n10127) );
  NAND2_X1 U12763 ( .A1(n10125), .A2(n10124), .ZN(n10126) );
  NAND2_X1 U12764 ( .A1(n10127), .A2(n10126), .ZN(n10131) );
  NOR2_X1 U12765 ( .A1(n10132), .A2(n10131), .ZN(n10128) );
  NAND2_X1 U12766 ( .A1(n10129), .A2(n10128), .ZN(n10137) );
  INV_X1 U12767 ( .A(n10130), .ZN(n10134) );
  INV_X1 U12768 ( .A(n10131), .ZN(n10133) );
  NAND2_X1 U12769 ( .A1(n10137), .A2(n10136), .ZN(n10139) );
  OR2_X1 U12770 ( .A1(n10533), .A2(P2_U3088), .ZN(n12059) );
  INV_X1 U12771 ( .A(n12059), .ZN(n10138) );
  OAI21_X1 U12772 ( .B1(n10140), .B2(n10139), .A(n10138), .ZN(n10146) );
  NOR4_X1 U12773 ( .A1(n15514), .A2(n12477), .A3(n14323), .A4(n10141), .ZN(
        n10144) );
  OAI21_X1 U12774 ( .B1(n10142), .B2(n12059), .A(P2_B_REG_SCAN_IN), .ZN(n10143) );
  OR2_X1 U12775 ( .A1(n10144), .A2(n10143), .ZN(n10145) );
  NAND2_X1 U12776 ( .A1(n10146), .A2(n10145), .ZN(P2_U3328) );
  INV_X1 U12777 ( .A(n10182), .ZN(n15716) );
  INV_X1 U12778 ( .A(n10148), .ZN(n13292) );
  NAND2_X1 U12779 ( .A1(n13722), .A2(n13721), .ZN(n13720) );
  NAND2_X1 U12780 ( .A1(n13720), .A2(n10151), .ZN(n10152) );
  NOR2_X1 U12781 ( .A1(n13750), .A2(n15690), .ZN(n10153) );
  AOI21_X1 U12782 ( .B1(n13299), .B2(n13877), .A(n10153), .ZN(n10155) );
  INV_X1 U12783 ( .A(n13728), .ZN(n15693) );
  NAND2_X1 U12784 ( .A1(n13717), .A2(n15693), .ZN(n10154) );
  NAND2_X1 U12785 ( .A1(n10157), .A2(n7583), .ZN(P3_U3485) );
  INV_X1 U12786 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n10158) );
  NAND2_X1 U12787 ( .A1(n10159), .A2(n7584), .ZN(P3_U3453) );
  INV_X1 U12788 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n10160) );
  NOR2_X1 U12789 ( .A1(n15543), .A2(n10160), .ZN(n10161) );
  OAI21_X1 U12790 ( .B1(n10164), .B2(n15541), .A(n10163), .ZN(P2_U3496) );
  NAND2_X1 U12791 ( .A1(n13722), .A2(n10165), .ZN(n10167) );
  NAND2_X1 U12792 ( .A1(n10168), .A2(n10169), .ZN(n10171) );
  NAND2_X1 U12793 ( .A1(n10171), .A2(n10170), .ZN(n10172) );
  OAI21_X1 U12794 ( .B1(n10173), .B2(n13297), .A(n10172), .ZN(n10174) );
  NAND2_X1 U12795 ( .A1(n10174), .A2(n13874), .ZN(n10181) );
  INV_X1 U12796 ( .A(n10175), .ZN(n10176) );
  AOI21_X2 U12797 ( .B1(n13297), .B2(n10176), .A(n13698), .ZN(n13126) );
  NOR2_X1 U12798 ( .A1(n13126), .A2(n13728), .ZN(n10179) );
  OAI22_X1 U12799 ( .A1(n10177), .A2(n15689), .B1(n13724), .B2(n15690), .ZN(
        n10178) );
  NOR2_X2 U12800 ( .A1(n10179), .A2(n10178), .ZN(n10180) );
  INV_X1 U12801 ( .A(n14033), .ZN(n10184) );
  NAND2_X1 U12802 ( .A1(n10186), .A2(n10185), .ZN(P3_U3454) );
  INV_X1 U12803 ( .A(n10188), .ZN(n10191) );
  NAND2_X1 U12804 ( .A1(n10191), .A2(n10190), .ZN(P3_U3486) );
  NAND2_X1 U12805 ( .A1(n10193), .A2(n10192), .ZN(n14800) );
  NAND2_X1 U12806 ( .A1(n12494), .A2(n12766), .ZN(n10195) );
  NAND2_X1 U12807 ( .A1(n12751), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n10194) );
  NAND2_X1 U12808 ( .A1(n15004), .A2(n13113), .ZN(n10197) );
  OR2_X1 U12809 ( .A1(n15004), .A2(n13113), .ZN(n10196) );
  NAND2_X1 U12810 ( .A1(n14800), .A2(n14799), .ZN(n14801) );
  NAND2_X1 U12811 ( .A1(n14801), .A2(n10197), .ZN(n10209) );
  NAND2_X1 U12812 ( .A1(n13373), .A2(n7861), .ZN(n10199) );
  NAND2_X1 U12813 ( .A1(n12751), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n10198) );
  NAND2_X1 U12814 ( .A1(n12754), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n10207) );
  NAND2_X1 U12815 ( .A1(n10200), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n10206) );
  INV_X1 U12816 ( .A(n10201), .ZN(n10202) );
  NAND2_X1 U12817 ( .A1(n10202), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n14785) );
  OR2_X1 U12818 ( .A1(n10203), .A2(n14785), .ZN(n10205) );
  INV_X1 U12819 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n14789) );
  OR2_X1 U12820 ( .A1(n8115), .A2(n14789), .ZN(n10204) );
  NAND4_X1 U12821 ( .A1(n10207), .A2(n10206), .A3(n10205), .A4(n10204), .ZN(
        n14802) );
  XNOR2_X1 U12822 ( .A(n12747), .B(n14802), .ZN(n12808) );
  NOR2_X1 U12823 ( .A1(n13113), .A2(n14869), .ZN(n14791) );
  INV_X1 U12824 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n15001) );
  OR2_X1 U12825 ( .A1(n10210), .A2(n15001), .ZN(n10213) );
  INV_X1 U12826 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n14779) );
  OR2_X1 U12827 ( .A1(n8115), .A2(n14779), .ZN(n10212) );
  INV_X1 U12828 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n15077) );
  OR2_X1 U12829 ( .A1(n12758), .A2(n15077), .ZN(n10211) );
  AND3_X1 U12830 ( .A1(n10213), .A2(n10212), .A3(n10211), .ZN(n12762) );
  INV_X1 U12831 ( .A(P1_B_REG_SCAN_IN), .ZN(n10215) );
  NOR2_X1 U12832 ( .A1(n10214), .A2(n10215), .ZN(n10216) );
  OR2_X1 U12833 ( .A1(n14871), .A2(n10216), .ZN(n14771) );
  NOR2_X1 U12834 ( .A1(n12762), .A2(n14771), .ZN(n14788) );
  NOR2_X1 U12835 ( .A1(n14791), .A2(n14788), .ZN(n10217) );
  INV_X1 U12836 ( .A(n15004), .ZN(n14817) );
  NAND2_X1 U12837 ( .A1(n14826), .A2(n13101), .ZN(n10219) );
  OAI21_X1 U12838 ( .B1(n14817), .B2(n13113), .A(n14808), .ZN(n10221) );
  XNOR2_X1 U12839 ( .A(n10221), .B(n12808), .ZN(n14783) );
  INV_X1 U12840 ( .A(n10222), .ZN(n10223) );
  NAND2_X1 U12841 ( .A1(n14783), .A2(n15321), .ZN(n10224) );
  INV_X1 U12842 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n10225) );
  OR2_X1 U12843 ( .A1(n15324), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n10227) );
  NAND2_X1 U12844 ( .A1(n10228), .A2(n10227), .ZN(n10229) );
  NAND2_X1 U12845 ( .A1(n10229), .A2(n7598), .ZN(P1_U3525) );
  INV_X1 U12846 ( .A(n10533), .ZN(n10230) );
  NOR2_X1 U12847 ( .A1(n10231), .A2(n10230), .ZN(n10537) );
  INV_X2 U12848 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U12849 ( .A(n10431), .ZN(n10232) );
  INV_X2 U12850 ( .A(n14640), .ZN(P1_U4016) );
  INV_X1 U12851 ( .A(n11103), .ZN(n10233) );
  NAND2_X1 U12852 ( .A1(n14367), .A2(n12878), .ZN(n10312) );
  INV_X1 U12853 ( .A(n10312), .ZN(n10320) );
  XNOR2_X1 U12854 ( .A(n14390), .B(n12882), .ZN(n10319) );
  NAND2_X1 U12855 ( .A1(n10746), .A2(n10336), .ZN(n10712) );
  NAND2_X1 U12856 ( .A1(n10235), .A2(n10712), .ZN(n10551) );
  AND2_X1 U12857 ( .A1(n10244), .A2(n10236), .ZN(n10237) );
  OR2_X1 U12858 ( .A1(n10551), .A2(n10237), .ZN(n10574) );
  NAND2_X1 U12859 ( .A1(n14170), .A2(n12878), .ZN(n10240) );
  XNOR2_X1 U12860 ( .A(n10240), .B(n10238), .ZN(n10573) );
  NAND2_X1 U12861 ( .A1(n10574), .A2(n10573), .ZN(n10242) );
  INV_X1 U12862 ( .A(n10238), .ZN(n10239) );
  NAND2_X1 U12863 ( .A1(n10240), .A2(n10239), .ZN(n10241) );
  NAND2_X1 U12864 ( .A1(n14169), .A2(n12878), .ZN(n10252) );
  XNOR2_X1 U12865 ( .A(n10243), .B(n10244), .ZN(n10250) );
  XNOR2_X1 U12866 ( .A(n10252), .B(n10250), .ZN(n10658) );
  INV_X1 U12867 ( .A(n10250), .ZN(n10251) );
  NAND2_X1 U12868 ( .A1(n10252), .A2(n10251), .ZN(n10897) );
  INV_X1 U12869 ( .A(n10897), .ZN(n10253) );
  NOR2_X1 U12870 ( .A1(n10901), .A2(n10253), .ZN(n10254) );
  NAND2_X1 U12871 ( .A1(n14166), .A2(n12878), .ZN(n10257) );
  XNOR2_X1 U12872 ( .A(n10256), .B(n10257), .ZN(n10793) );
  INV_X1 U12873 ( .A(n10256), .ZN(n10258) );
  NAND2_X1 U12874 ( .A1(n10258), .A2(n10257), .ZN(n10259) );
  XNOR2_X1 U12875 ( .A(n11074), .B(n12882), .ZN(n10260) );
  NAND2_X1 U12876 ( .A1(n14165), .A2(n12878), .ZN(n10261) );
  XNOR2_X1 U12877 ( .A(n10260), .B(n10261), .ZN(n10886) );
  NAND2_X1 U12878 ( .A1(n10885), .A2(n10886), .ZN(n10884) );
  INV_X1 U12879 ( .A(n10260), .ZN(n10262) );
  NAND2_X1 U12880 ( .A1(n10262), .A2(n10261), .ZN(n10263) );
  XNOR2_X1 U12881 ( .A(n11685), .B(n12882), .ZN(n10264) );
  AND2_X1 U12882 ( .A1(n14164), .A2(n12878), .ZN(n10265) );
  NAND2_X1 U12883 ( .A1(n10264), .A2(n10265), .ZN(n10268) );
  NAND2_X1 U12884 ( .A1(n10268), .A2(n10266), .ZN(n11235) );
  XNOR2_X1 U12885 ( .A(n11088), .B(n12882), .ZN(n10271) );
  NAND2_X1 U12886 ( .A1(n14163), .A2(n12878), .ZN(n10269) );
  XNOR2_X1 U12887 ( .A(n10271), .B(n10269), .ZN(n11090) );
  NAND2_X1 U12888 ( .A1(n11091), .A2(n11090), .ZN(n11089) );
  INV_X1 U12889 ( .A(n10269), .ZN(n10270) );
  NAND2_X1 U12890 ( .A1(n10271), .A2(n10270), .ZN(n10272) );
  NAND2_X1 U12891 ( .A1(n11089), .A2(n10272), .ZN(n11244) );
  XNOR2_X1 U12892 ( .A(n15523), .B(n12877), .ZN(n10273) );
  NAND2_X1 U12893 ( .A1(n14162), .A2(n12878), .ZN(n10274) );
  NAND2_X1 U12894 ( .A1(n10273), .A2(n10274), .ZN(n11243) );
  INV_X1 U12895 ( .A(n10273), .ZN(n10276) );
  INV_X1 U12896 ( .A(n10274), .ZN(n10275) );
  NAND2_X1 U12897 ( .A1(n10276), .A2(n10275), .ZN(n11242) );
  XNOR2_X1 U12898 ( .A(n11995), .B(n12877), .ZN(n10277) );
  NAND2_X1 U12899 ( .A1(n14161), .A2(n12878), .ZN(n10278) );
  NAND2_X1 U12900 ( .A1(n10277), .A2(n10278), .ZN(n10283) );
  INV_X1 U12901 ( .A(n10277), .ZN(n10280) );
  INV_X1 U12902 ( .A(n10278), .ZN(n10279) );
  NAND2_X1 U12903 ( .A1(n10280), .A2(n10279), .ZN(n10281) );
  NAND2_X1 U12904 ( .A1(n10283), .A2(n10281), .ZN(n11449) );
  INV_X1 U12905 ( .A(n11449), .ZN(n10282) );
  XNOR2_X1 U12906 ( .A(n15533), .B(n12877), .ZN(n10285) );
  NAND2_X1 U12907 ( .A1(n14160), .A2(n12878), .ZN(n10284) );
  XNOR2_X1 U12908 ( .A(n10285), .B(n10284), .ZN(n11615) );
  XNOR2_X1 U12909 ( .A(n12257), .B(n12882), .ZN(n10288) );
  NAND2_X1 U12910 ( .A1(n14159), .A2(n12878), .ZN(n10286) );
  XNOR2_X1 U12911 ( .A(n10288), .B(n10286), .ZN(n11747) );
  INV_X1 U12912 ( .A(n10286), .ZN(n10287) );
  NAND2_X1 U12913 ( .A1(n10288), .A2(n10287), .ZN(n10289) );
  XNOR2_X1 U12914 ( .A(n12051), .B(n12877), .ZN(n10290) );
  NAND2_X1 U12915 ( .A1(n14158), .A2(n12878), .ZN(n10291) );
  NAND2_X1 U12916 ( .A1(n10290), .A2(n10291), .ZN(n12062) );
  INV_X1 U12917 ( .A(n10290), .ZN(n10293) );
  INV_X1 U12918 ( .A(n10291), .ZN(n10292) );
  NAND2_X1 U12919 ( .A1(n10293), .A2(n10292), .ZN(n10294) );
  NAND2_X1 U12920 ( .A1(n12062), .A2(n10294), .ZN(n12016) );
  XNOR2_X1 U12921 ( .A(n12080), .B(n12877), .ZN(n10297) );
  NAND2_X1 U12922 ( .A1(n14157), .A2(n12878), .ZN(n10298) );
  XNOR2_X1 U12923 ( .A(n10297), .B(n10298), .ZN(n12064) );
  INV_X1 U12924 ( .A(n12064), .ZN(n10296) );
  AND2_X1 U12925 ( .A1(n10296), .A2(n12062), .ZN(n10301) );
  INV_X1 U12926 ( .A(n10297), .ZN(n10300) );
  INV_X1 U12927 ( .A(n10298), .ZN(n10299) );
  XNOR2_X1 U12928 ( .A(n12321), .B(n12877), .ZN(n10302) );
  NAND2_X1 U12929 ( .A1(n14156), .A2(n12878), .ZN(n10303) );
  NAND2_X1 U12930 ( .A1(n10302), .A2(n10303), .ZN(n10307) );
  INV_X1 U12931 ( .A(n10302), .ZN(n10305) );
  INV_X1 U12932 ( .A(n10303), .ZN(n10304) );
  NAND2_X1 U12933 ( .A1(n10305), .A2(n10304), .ZN(n10306) );
  AND2_X1 U12934 ( .A1(n10307), .A2(n10306), .ZN(n12204) );
  NAND2_X1 U12935 ( .A1(n12203), .A2(n12204), .ZN(n12202) );
  NAND2_X1 U12936 ( .A1(n14155), .A2(n12878), .ZN(n12401) );
  XNOR2_X1 U12937 ( .A(n14475), .B(n12877), .ZN(n10311) );
  NAND2_X1 U12938 ( .A1(n14154), .A2(n12878), .ZN(n10310) );
  NAND2_X1 U12939 ( .A1(n10311), .A2(n10310), .ZN(n14092) );
  OAI21_X1 U12940 ( .B1(n10311), .B2(n10310), .A(n14092), .ZN(n12498) );
  XNOR2_X1 U12941 ( .A(n12565), .B(n12882), .ZN(n10313) );
  AND2_X1 U12942 ( .A1(n14153), .A2(n12878), .ZN(n10314) );
  NAND2_X1 U12943 ( .A1(n10313), .A2(n10314), .ZN(n14090) );
  XNOR2_X1 U12944 ( .A(n10319), .B(n10312), .ZN(n14128) );
  INV_X1 U12945 ( .A(n10313), .ZN(n10316) );
  INV_X1 U12946 ( .A(n10314), .ZN(n10315) );
  NAND2_X1 U12947 ( .A1(n10316), .A2(n10315), .ZN(n14125) );
  INV_X1 U12948 ( .A(n14092), .ZN(n10317) );
  NAND2_X1 U12949 ( .A1(n14090), .A2(n10317), .ZN(n10318) );
  AND2_X1 U12950 ( .A1(n14356), .A2(n12878), .ZN(n10322) );
  XNOR2_X1 U12951 ( .A(n14375), .B(n12882), .ZN(n10321) );
  NOR2_X1 U12952 ( .A1(n10321), .A2(n10322), .ZN(n10323) );
  AOI21_X1 U12953 ( .B1(n10322), .B2(n10321), .A(n10323), .ZN(n14066) );
  INV_X1 U12954 ( .A(n10323), .ZN(n10324) );
  NAND2_X1 U12955 ( .A1(n14065), .A2(n10324), .ZN(n14118) );
  XNOR2_X1 U12956 ( .A(n14454), .B(n12882), .ZN(n10326) );
  AND2_X1 U12957 ( .A1(n14370), .A2(n12878), .ZN(n10325) );
  NOR2_X1 U12958 ( .A1(n10326), .A2(n10325), .ZN(n14114) );
  NAND2_X1 U12959 ( .A1(n10326), .A2(n10325), .ZN(n14115) );
  XNOR2_X1 U12960 ( .A(n14338), .B(n12882), .ZN(n10327) );
  NAND2_X1 U12961 ( .A1(n14355), .A2(n12878), .ZN(n10328) );
  XNOR2_X1 U12962 ( .A(n10327), .B(n10328), .ZN(n14076) );
  NAND2_X1 U12963 ( .A1(n14077), .A2(n14076), .ZN(n14075) );
  INV_X1 U12964 ( .A(n10328), .ZN(n10329) );
  NAND2_X1 U12965 ( .A1(n10327), .A2(n10329), .ZN(n10330) );
  NAND2_X1 U12966 ( .A1(n14075), .A2(n10330), .ZN(n12859) );
  XNOR2_X1 U12967 ( .A(n14443), .B(n12882), .ZN(n12858) );
  XNOR2_X1 U12968 ( .A(n12859), .B(n12858), .ZN(n10335) );
  NAND2_X1 U12969 ( .A1(n14335), .A2(n12878), .ZN(n10334) );
  OR3_X1 U12970 ( .A1(n10331), .A2(n15511), .A3(n10706), .ZN(n10341) );
  INV_X1 U12971 ( .A(n10534), .ZN(n10332) );
  AND2_X1 U12972 ( .A1(n15525), .A2(n10332), .ZN(n10333) );
  NOR2_X1 U12973 ( .A1(n10335), .A2(n10334), .ZN(n12861) );
  AOI211_X1 U12974 ( .C1(n10335), .C2(n10334), .A(n14148), .B(n12861), .ZN(
        n10352) );
  INV_X1 U12975 ( .A(n10336), .ZN(n10337) );
  NOR2_X1 U12976 ( .A1(n10337), .A2(n11708), .ZN(n11008) );
  NAND2_X1 U12977 ( .A1(n10348), .A2(n11008), .ZN(n10339) );
  NOR2_X1 U12978 ( .A1(n14321), .A2(n14102), .ZN(n10351) );
  NAND2_X1 U12979 ( .A1(n10341), .A2(n10340), .ZN(n10345) );
  AND2_X1 U12980 ( .A1(n10343), .A2(n10342), .ZN(n10344) );
  NAND2_X1 U12981 ( .A1(n10345), .A2(n10344), .ZN(n10553) );
  INV_X1 U12982 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10346) );
  OAI22_X1 U12983 ( .A1(n14318), .A2(n14140), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10346), .ZN(n10350) );
  AND2_X1 U12984 ( .A1(n14131), .A2(n14369), .ZN(n14108) );
  INV_X1 U12985 ( .A(n14108), .ZN(n14142) );
  AND2_X1 U12986 ( .A1(n14131), .A2(n14368), .ZN(n14109) );
  INV_X1 U12987 ( .A(n14109), .ZN(n14143) );
  OAI22_X1 U12988 ( .A1(n14326), .A2(n14142), .B1(n14324), .B2(n14143), .ZN(
        n10349) );
  OR4_X1 U12989 ( .A1(n10352), .A2(n10351), .A3(n10350), .A4(n10349), .ZN(
        P2_U3207) );
  MUX2_X1 U12990 ( .A(n10353), .B(P1_REG1_REG_1__SCAN_IN), .S(n14672), .Z(
        n14670) );
  NAND3_X1 U12991 ( .A1(n14670), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_REG1_REG_0__SCAN_IN), .ZN(n14668) );
  OAI21_X1 U12992 ( .B1(n14672), .B2(n10353), .A(n14668), .ZN(n14688) );
  MUX2_X1 U12993 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n7731), .S(n14681), .Z(
        n14689) );
  XNOR2_X1 U12994 ( .A(n10475), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n10360) );
  INV_X1 U12995 ( .A(n11142), .ZN(n10355) );
  INV_X1 U12996 ( .A(n10354), .ZN(n10356) );
  NAND2_X1 U12997 ( .A1(n10356), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12846) );
  NAND2_X1 U12998 ( .A1(n10355), .A2(n12846), .ZN(n10370) );
  OR2_X1 U12999 ( .A1(n12771), .A2(n10356), .ZN(n10358) );
  NAND2_X1 U13000 ( .A1(n10358), .A2(n10357), .ZN(n10369) );
  INV_X1 U13001 ( .A(n10369), .ZN(n10359) );
  AND2_X1 U13002 ( .A1(n10370), .A2(n10359), .ZN(n10470) );
  INV_X1 U13003 ( .A(n10470), .ZN(n10368) );
  INV_X1 U13004 ( .A(n10214), .ZN(n10463) );
  OR2_X1 U13005 ( .A1(n10368), .A2(n10463), .ZN(n14759) );
  AOI211_X1 U13006 ( .C1(n10361), .C2(n10360), .A(n10474), .B(n14759), .ZN(
        n10375) );
  NOR2_X1 U13007 ( .A1(n12993), .A2(n10214), .ZN(n10362) );
  MUX2_X1 U13008 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n14673), .S(n14672), .Z(
        n10363) );
  OR3_X1 U13009 ( .A1(n10363), .A2(n10462), .A3(n10666), .ZN(n14685) );
  INV_X1 U13010 ( .A(n14672), .ZN(n14667) );
  NAND2_X1 U13011 ( .A1(n14667), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n14684) );
  MUX2_X1 U13012 ( .A(n7730), .B(P1_REG2_REG_2__SCAN_IN), .S(n14681), .Z(
        n14683) );
  INV_X1 U13013 ( .A(n14681), .ZN(n10401) );
  NOR2_X1 U13014 ( .A1(n10401), .A2(n7730), .ZN(n10365) );
  MUX2_X1 U13015 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10480), .S(n10475), .Z(
        n10364) );
  OAI21_X1 U13016 ( .B1(n14682), .B2(n10365), .A(n10364), .ZN(n10479) );
  INV_X1 U13017 ( .A(n10479), .ZN(n10367) );
  NOR3_X1 U13018 ( .A1(n14682), .A2(n10365), .A3(n10364), .ZN(n10366) );
  NOR3_X1 U13019 ( .A1(n15266), .A2(n10367), .A3(n10366), .ZN(n10374) );
  OR2_X1 U13020 ( .A1(n10368), .A2(n10465), .ZN(n14757) );
  INV_X1 U13021 ( .A(n10475), .ZN(n10481) );
  NOR2_X1 U13022 ( .A1(n14757), .A2(n10481), .ZN(n10373) );
  NAND2_X1 U13023 ( .A1(n10370), .A2(n10369), .ZN(n15271) );
  INV_X1 U13024 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10371) );
  INV_X1 U13025 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n11312) );
  OAI22_X1 U13026 ( .A1(n15271), .A2(n10371), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11312), .ZN(n10372) );
  OR4_X1 U13027 ( .A1(n10375), .A2(n10374), .A3(n10373), .A4(n10372), .ZN(
        P1_U3246) );
  MUX2_X1 U13028 ( .A(P2_RD_REG_SCAN_IN), .B(n7617), .S(P1_RD_REG_SCAN_IN), 
        .Z(n10377) );
  NAND2_X1 U13029 ( .A1(n10377), .A2(n10376), .ZN(U29) );
  NOR2_X1 U13030 ( .A1(n6676), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14037) );
  NAND2_X1 U13031 ( .A1(n10046), .A2(P3_U3151), .ZN(n14049) );
  OAI222_X1 U13032 ( .A1(n12850), .A2(n10379), .B1(n14049), .B2(n10378), .C1(
        P3_U3151), .C2(n10881), .ZN(P3_U3294) );
  INV_X1 U13033 ( .A(n15578), .ZN(n11903) );
  INV_X1 U13034 ( .A(SI_4_), .ZN(n10382) );
  INV_X1 U13035 ( .A(n10380), .ZN(n10381) );
  OAI222_X1 U13036 ( .A1(P3_U3151), .A2(n11903), .B1(n14049), .B2(n10382), 
        .C1(n12850), .C2(n10381), .ZN(P3_U3291) );
  NOR2_X1 U13037 ( .A1(n6676), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14525) );
  INV_X2 U13038 ( .A(n14525), .ZN(n12959) );
  NAND2_X1 U13039 ( .A1(n10046), .A2(P2_U3088), .ZN(n14531) );
  INV_X1 U13040 ( .A(n14531), .ZN(n12057) );
  INV_X1 U13041 ( .A(n12057), .ZN(n12957) );
  NAND2_X1 U13042 ( .A1(n10046), .A2(P1_U3086), .ZN(n13374) );
  INV_X1 U13043 ( .A(n13374), .ZN(n12964) );
  INV_X1 U13044 ( .A(n12964), .ZN(n12476) );
  NOR2_X1 U13045 ( .A1(n6676), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12963) );
  INV_X2 U13046 ( .A(n12963), .ZN(n13377) );
  OAI222_X1 U13047 ( .A1(n12476), .A2(n6849), .B1(n13377), .B2(n10385), .C1(
        n14672), .C2(P1_U3086), .ZN(P1_U3354) );
  INV_X1 U13048 ( .A(n15599), .ZN(n11864) );
  INV_X1 U13049 ( .A(SI_5_), .ZN(n10388) );
  INV_X1 U13050 ( .A(n10386), .ZN(n10387) );
  OAI222_X1 U13051 ( .A1(P3_U3151), .A2(n11864), .B1(n13382), .B2(n10388), 
        .C1(n12850), .C2(n10387), .ZN(P3_U3290) );
  INV_X1 U13052 ( .A(SI_7_), .ZN(n10391) );
  INV_X1 U13053 ( .A(n10389), .ZN(n10390) );
  OAI222_X1 U13054 ( .A1(P3_U3151), .A2(n15633), .B1(n13382), .B2(n10391), 
        .C1(n12850), .C2(n10390), .ZN(P3_U3288) );
  OAI222_X1 U13055 ( .A1(n12850), .A2(n10393), .B1(n13382), .B2(n10392), .C1(
        P3_U3151), .C2(n15649), .ZN(P3_U3287) );
  INV_X1 U13056 ( .A(n11900), .ZN(n11835) );
  INV_X1 U13057 ( .A(SI_2_), .ZN(n10396) );
  INV_X1 U13058 ( .A(n10394), .ZN(n10395) );
  OAI222_X1 U13059 ( .A1(P3_U3151), .A2(n11835), .B1(n13382), .B2(n10396), 
        .C1(n12850), .C2(n10395), .ZN(P3_U3293) );
  INV_X1 U13060 ( .A(SI_9_), .ZN(n10399) );
  INV_X1 U13061 ( .A(n10397), .ZN(n10398) );
  OAI222_X1 U13062 ( .A1(P3_U3151), .A2(n15670), .B1(n13382), .B2(n10399), 
        .C1(n12850), .C2(n10398), .ZN(P3_U3286) );
  INV_X1 U13063 ( .A(n10400), .ZN(n10408) );
  OAI222_X1 U13064 ( .A1(n12476), .A2(n10402), .B1(n13377), .B2(n10408), .C1(
        P1_U3086), .C2(n10401), .ZN(P1_U3353) );
  INV_X1 U13065 ( .A(n10403), .ZN(n10406) );
  OAI222_X1 U13066 ( .A1(n12476), .A2(n10404), .B1(n13377), .B2(n10406), .C1(
        P1_U3086), .C2(n10481), .ZN(P1_U3352) );
  INV_X1 U13067 ( .A(n15356), .ZN(n10405) );
  OAI222_X1 U13068 ( .A1(n12959), .A2(n10407), .B1(n14531), .B2(n10406), .C1(
        P2_U3088), .C2(n10405), .ZN(P2_U3324) );
  OAI222_X1 U13069 ( .A1(n12959), .A2(n10409), .B1(n14531), .B2(n10408), .C1(
        P2_U3088), .C2(n10978), .ZN(P2_U3325) );
  INV_X1 U13070 ( .A(n15561), .ZN(n11902) );
  INV_X1 U13071 ( .A(SI_3_), .ZN(n10412) );
  INV_X1 U13072 ( .A(n10410), .ZN(n10411) );
  OAI222_X1 U13073 ( .A1(P3_U3151), .A2(n11902), .B1(n13382), .B2(n10412), 
        .C1(n12850), .C2(n10411), .ZN(P3_U3292) );
  INV_X1 U13074 ( .A(n10413), .ZN(n10414) );
  OAI222_X1 U13075 ( .A1(P3_U3151), .A2(n12262), .B1(n13382), .B2(n10415), 
        .C1(n12850), .C2(n10414), .ZN(P3_U3285) );
  OAI222_X1 U13076 ( .A1(P3_U3151), .A2(n10417), .B1(n12850), .B2(n10416), 
        .C1(n9810), .C2(n14049), .ZN(P3_U3295) );
  OAI222_X1 U13077 ( .A1(P3_U3151), .A2(n15615), .B1(n12850), .B2(n10419), 
        .C1(n10418), .C2(n14049), .ZN(P3_U3289) );
  INV_X1 U13078 ( .A(n10420), .ZN(n10421) );
  OAI222_X1 U13079 ( .A1(P3_U3151), .A2(n12339), .B1(n13382), .B2(n10422), 
        .C1(n12850), .C2(n10421), .ZN(P3_U3284) );
  INV_X1 U13080 ( .A(n10423), .ZN(n10426) );
  INV_X1 U13081 ( .A(n10483), .ZN(n10673) );
  OAI222_X1 U13082 ( .A1(n12476), .A2(n10424), .B1(n13377), .B2(n10426), .C1(
        P1_U3086), .C2(n10673), .ZN(P1_U3351) );
  INV_X1 U13083 ( .A(n15369), .ZN(n10425) );
  OAI222_X1 U13084 ( .A1(n12959), .A2(n10427), .B1(n14531), .B2(n10426), .C1(
        P2_U3088), .C2(n10425), .ZN(P2_U3323) );
  NAND2_X1 U13085 ( .A1(n11142), .A2(n10500), .ZN(n15284) );
  INV_X1 U13086 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10429) );
  INV_X1 U13087 ( .A(n10501), .ZN(n10428) );
  AOI22_X1 U13088 ( .A1(n15284), .A2(n10429), .B1(n10428), .B2(n10431), .ZN(
        P1_U3446) );
  INV_X1 U13089 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10433) );
  INV_X1 U13090 ( .A(n10430), .ZN(n10432) );
  AOI22_X1 U13091 ( .A1(n15284), .A2(n10433), .B1(n10432), .B2(n10431), .ZN(
        P1_U3445) );
  INV_X1 U13092 ( .A(n10434), .ZN(n10435) );
  OAI222_X1 U13093 ( .A1(P3_U3151), .A2(n13540), .B1(n13382), .B2(n10436), 
        .C1(n12850), .C2(n10435), .ZN(P3_U3283) );
  INV_X1 U13094 ( .A(n10437), .ZN(n10440) );
  INV_X1 U13095 ( .A(n15382), .ZN(n10438) );
  OAI222_X1 U13096 ( .A1(n12959), .A2(n10439), .B1(n14531), .B2(n10440), .C1(
        P2_U3088), .C2(n10438), .ZN(P2_U3322) );
  OAI222_X1 U13097 ( .A1(n12476), .A2(n10441), .B1(n13377), .B2(n10440), .C1(
        P1_U3086), .C2(n10484), .ZN(P1_U3350) );
  NAND2_X1 U13098 ( .A1(n14640), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n10442) );
  OAI21_X1 U13099 ( .B1(n12999), .B2(n14640), .A(n10442), .ZN(P1_U3574) );
  INV_X1 U13100 ( .A(n10443), .ZN(n10446) );
  INV_X1 U13101 ( .A(n15394), .ZN(n10444) );
  OAI222_X1 U13102 ( .A1(n12959), .A2(n10445), .B1(n14531), .B2(n10446), .C1(
        P2_U3088), .C2(n10444), .ZN(P2_U3321) );
  INV_X1 U13103 ( .A(n10523), .ZN(n10492) );
  OAI222_X1 U13104 ( .A1(n12476), .A2(n10447), .B1(n13377), .B2(n10446), .C1(
        P1_U3086), .C2(n10492), .ZN(P1_U3349) );
  NOR2_X1 U13105 ( .A1(n14737), .A2(P1_U4016), .ZN(P1_U3085) );
  OAI222_X1 U13106 ( .A1(P3_U3151), .A2(n13560), .B1(n13382), .B2(n10449), 
        .C1(n12850), .C2(n10448), .ZN(P3_U3282) );
  INV_X1 U13107 ( .A(n10576), .ZN(n10450) );
  NAND2_X1 U13108 ( .A1(n10450), .A2(P2_U3947), .ZN(n10451) );
  OAI21_X1 U13109 ( .B1(n8807), .B2(P2_U3947), .A(n10451), .ZN(P2_U3531) );
  INV_X1 U13110 ( .A(n10452), .ZN(n10454) );
  OAI222_X1 U13111 ( .A1(n12959), .A2(n10453), .B1(n14531), .B2(n10454), .C1(
        P2_U3088), .C2(n7102), .ZN(P2_U3320) );
  INV_X1 U13112 ( .A(n10642), .ZN(n10646) );
  OAI222_X1 U13113 ( .A1(n12476), .A2(n10455), .B1(n13377), .B2(n10454), .C1(
        P1_U3086), .C2(n10646), .ZN(P1_U3348) );
  OAI222_X1 U13114 ( .A1(P3_U3151), .A2(n13583), .B1(n13382), .B2(n10457), 
        .C1(n12850), .C2(n10456), .ZN(P3_U3281) );
  INV_X1 U13115 ( .A(n10458), .ZN(n10460) );
  INV_X1 U13116 ( .A(n10727), .ZN(n10653) );
  OAI222_X1 U13117 ( .A1(n12476), .A2(n10459), .B1(n13377), .B2(n10460), .C1(
        P1_U3086), .C2(n10653), .ZN(P1_U3347) );
  INV_X1 U13118 ( .A(n10984), .ZN(n15418) );
  OAI222_X1 U13119 ( .A1(n12959), .A2(n10461), .B1(n14531), .B2(n10460), .C1(
        P2_U3088), .C2(n15418), .ZN(P2_U3319) );
  NAND2_X1 U13120 ( .A1(n10463), .A2(n10462), .ZN(n10464) );
  NAND2_X1 U13121 ( .A1(n10465), .A2(n10464), .ZN(n10667) );
  AOI21_X1 U13122 ( .B1(n10504), .B2(n10214), .A(n10667), .ZN(n10466) );
  MUX2_X1 U13123 ( .A(n10667), .B(n10466), .S(n10666), .Z(n10469) );
  OAI22_X1 U13124 ( .A1(n15271), .A2(n6850), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10467), .ZN(n10468) );
  AOI21_X1 U13125 ( .B1(n10470), .B2(n10469), .A(n10468), .ZN(n10472) );
  INV_X1 U13126 ( .A(n14759), .ZN(n15260) );
  NAND3_X1 U13127 ( .A1(n15260), .A2(P1_IR_REG_0__SCAN_IN), .A3(n10504), .ZN(
        n10471) );
  NAND2_X1 U13128 ( .A1(n10472), .A2(n10471), .ZN(P1_U3243) );
  INV_X1 U13129 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10473) );
  MUX2_X1 U13130 ( .A(n10473), .B(P1_REG1_REG_6__SCAN_IN), .S(n10523), .Z(
        n10478) );
  XNOR2_X1 U13131 ( .A(n10483), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n10675) );
  NOR2_X1 U13132 ( .A1(n10676), .A2(n10675), .ZN(n10674) );
  AOI21_X1 U13133 ( .B1(n10483), .B2(P1_REG1_REG_4__SCAN_IN), .A(n10674), .ZN(
        n10560) );
  MUX2_X1 U13134 ( .A(n10476), .B(P1_REG1_REG_5__SCAN_IN), .S(n10484), .Z(
        n10559) );
  NAND2_X1 U13135 ( .A1(n10560), .A2(n10559), .ZN(n10558) );
  OAI21_X1 U13136 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n10561), .A(n10558), .ZN(
        n10477) );
  NOR2_X1 U13137 ( .A1(n10477), .A2(n10478), .ZN(n10519) );
  AOI211_X1 U13138 ( .C1(n10478), .C2(n10477), .A(n14759), .B(n10519), .ZN(
        n10495) );
  OAI21_X1 U13139 ( .B1(n10481), .B2(n10480), .A(n10479), .ZN(n10670) );
  MUX2_X1 U13140 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10482), .S(n10483), .Z(
        n10671) );
  AOI22_X1 U13141 ( .A1(n10670), .A2(n10671), .B1(P1_REG2_REG_4__SCAN_IN), 
        .B2(n10483), .ZN(n10566) );
  MUX2_X1 U13142 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n7783), .S(n10484), .Z(
        n10565) );
  NOR2_X1 U13143 ( .A1(n10484), .A2(n7783), .ZN(n10487) );
  MUX2_X1 U13144 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10485), .S(n10523), .Z(
        n10486) );
  OAI21_X1 U13145 ( .B1(n10564), .B2(n10487), .A(n10486), .ZN(n10526) );
  INV_X1 U13146 ( .A(n10526), .ZN(n10489) );
  NOR3_X1 U13147 ( .A1(n10564), .A2(n10487), .A3(n10486), .ZN(n10488) );
  NOR3_X1 U13148 ( .A1(n15266), .A2(n10489), .A3(n10488), .ZN(n10494) );
  AND2_X1 U13149 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10490) );
  AOI21_X1 U13150 ( .B1(n14737), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n10490), .ZN(
        n10491) );
  OAI21_X1 U13151 ( .B1(n10492), .B2(n14757), .A(n10491), .ZN(n10493) );
  OR3_X1 U13152 ( .A1(n10495), .A2(n10494), .A3(n10493), .ZN(P1_U3249) );
  INV_X1 U13153 ( .A(n13610), .ZN(n13616) );
  OAI222_X1 U13154 ( .A1(P3_U3151), .A2(n13616), .B1(n13382), .B2(n10497), 
        .C1(n12850), .C2(n10496), .ZN(P3_U3280) );
  AND2_X1 U13155 ( .A1(n10498), .A2(P1_D_REG_1__SCAN_IN), .ZN(n10499) );
  OR2_X1 U13156 ( .A1(n10500), .A2(n10499), .ZN(n10502) );
  AND2_X1 U13157 ( .A1(n10502), .A2(n10501), .ZN(n11139) );
  NAND2_X1 U13158 ( .A1(n11137), .A2(n11139), .ZN(n10512) );
  NAND2_X1 U13159 ( .A1(n10512), .A2(n11141), .ZN(n10827) );
  INV_X1 U13160 ( .A(n15218), .ZN(n15186) );
  INV_X1 U13161 ( .A(n12577), .ZN(n12769) );
  OR2_X1 U13162 ( .A1(n13111), .A2(n15274), .ZN(n10507) );
  AOI21_X1 U13163 ( .B1(n14664), .B2(n10821), .A(n10505), .ZN(n10506) );
  OAI222_X1 U13164 ( .A1(n15274), .A2(n6681), .B1(n10697), .B2(n10603), .C1(
        n10503), .C2(n10666), .ZN(n10600) );
  XOR2_X1 U13165 ( .A(n10599), .B(n10600), .Z(n10665) );
  INV_X1 U13166 ( .A(n10512), .ZN(n10511) );
  NAND2_X1 U13167 ( .A1(n11142), .A2(n12771), .ZN(n10509) );
  NOR2_X1 U13168 ( .A1(n10509), .A2(n15224), .ZN(n10510) );
  NAND2_X1 U13169 ( .A1(n10665), .A2(n15179), .ZN(n10514) );
  NOR2_X1 U13170 ( .A1(n6865), .A2(n14871), .ZN(n15289) );
  NOR2_X2 U13171 ( .A1(n10512), .A2(n12843), .ZN(n15183) );
  NAND2_X1 U13172 ( .A1(n10827), .A2(n11140), .ZN(n10701) );
  AOI22_X1 U13173 ( .A1(n15289), .A2(n15183), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n10701), .ZN(n10513) );
  OAI211_X1 U13174 ( .C1(n15186), .C2(n15274), .A(n10514), .B(n10513), .ZN(
        P1_U3232) );
  INV_X1 U13175 ( .A(n10515), .ZN(n10517) );
  INV_X1 U13176 ( .A(n10909), .ZN(n10912) );
  OAI222_X1 U13177 ( .A1(n12476), .A2(n10516), .B1(n13377), .B2(n10517), .C1(
        P1_U3086), .C2(n10912), .ZN(P1_U3346) );
  INV_X1 U13178 ( .A(n11295), .ZN(n10990) );
  OAI222_X1 U13179 ( .A1(n12959), .A2(n10518), .B1(n14531), .B2(n10517), .C1(
        P2_U3088), .C2(n10990), .ZN(P2_U3318) );
  INV_X1 U13180 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10520) );
  MUX2_X1 U13181 ( .A(n10520), .B(P1_REG1_REG_7__SCAN_IN), .S(n10642), .Z(
        n10521) );
  AOI211_X1 U13182 ( .C1(n10522), .C2(n10521), .A(n14759), .B(n10641), .ZN(
        n10532) );
  NAND2_X1 U13183 ( .A1(n10523), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10525) );
  MUX2_X1 U13184 ( .A(n11487), .B(P1_REG2_REG_7__SCAN_IN), .S(n10642), .Z(
        n10524) );
  AOI21_X1 U13185 ( .B1(n10526), .B2(n10525), .A(n10524), .ZN(n10649) );
  AND3_X1 U13186 ( .A1(n10526), .A2(n10525), .A3(n10524), .ZN(n10527) );
  NOR3_X1 U13187 ( .A1(n15266), .A2(n10649), .A3(n10527), .ZN(n10531) );
  INV_X1 U13188 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10529) );
  INV_X1 U13189 ( .A(n14757), .ZN(n15263) );
  NAND2_X1 U13190 ( .A1(n15263), .A2(n10642), .ZN(n10528) );
  NAND2_X1 U13191 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n11644) );
  OAI211_X1 U13192 ( .C1(n15271), .C2(n10529), .A(n10528), .B(n11644), .ZN(
        n10530) );
  OR3_X1 U13193 ( .A1(n10532), .A2(n10531), .A3(n10530), .ZN(P1_U3250) );
  NAND2_X1 U13194 ( .A1(n10534), .A2(n10533), .ZN(n10536) );
  AND2_X1 U13195 ( .A1(n10536), .A2(n10535), .ZN(n10538) );
  NOR2_X1 U13196 ( .A1(n10543), .A2(P2_U3088), .ZN(n15333) );
  NOR2_X1 U13197 ( .A1(n8705), .A2(P2_U3088), .ZN(n12495) );
  NAND2_X1 U13198 ( .A1(n10543), .A2(n12495), .ZN(n10541) );
  INV_X1 U13199 ( .A(n10541), .ZN(n10539) );
  NOR2_X2 U13200 ( .A1(n10541), .A2(n10540), .ZN(n15484) );
  AOI22_X1 U13201 ( .A1(n15478), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n15484), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n10547) );
  INV_X1 U13202 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10545) );
  AND2_X1 U13203 ( .A1(n8705), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10542) );
  NAND2_X1 U13204 ( .A1(n10543), .A2(n10542), .ZN(n15489) );
  OAI21_X1 U13205 ( .B1(n15461), .B2(P2_REG2_REG_0__SCAN_IN), .A(n15489), .ZN(
        n10544) );
  AOI21_X1 U13206 ( .B1(n15484), .B2(n10545), .A(n10544), .ZN(n10546) );
  MUX2_X1 U13207 ( .A(n10547), .B(n10546), .S(P2_IR_REG_0__SCAN_IN), .Z(n10549) );
  NAND2_X1 U13208 ( .A1(P2_U3088), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n10548) );
  OAI211_X1 U13209 ( .C1(n15746), .C2(n15493), .A(n10549), .B(n10548), .ZN(
        P2_U3214) );
  INV_X1 U13210 ( .A(n10550), .ZN(n10552) );
  AOI21_X1 U13211 ( .B1(n10552), .B2(n12878), .A(n10551), .ZN(n10557) );
  NOR2_X1 U13212 ( .A1(n10553), .A2(P2_U3088), .ZN(n10661) );
  INV_X1 U13213 ( .A(n10661), .ZN(n10578) );
  AOI22_X1 U13214 ( .A1(n10578), .A2(P2_REG3_REG_0__SCAN_IN), .B1(n14146), 
        .B2(n10746), .ZN(n10556) );
  NOR2_X1 U13215 ( .A1(n10554), .A2(n14325), .ZN(n10685) );
  NAND2_X1 U13216 ( .A1(n14131), .A2(n10685), .ZN(n10555) );
  OAI211_X1 U13217 ( .C1(n10557), .C2(n14148), .A(n10556), .B(n10555), .ZN(
        P2_U3204) );
  OAI21_X1 U13218 ( .B1(n10560), .B2(n10559), .A(n10558), .ZN(n10569) );
  INV_X1 U13219 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10563) );
  NAND2_X1 U13220 ( .A1(n15263), .A2(n10561), .ZN(n10562) );
  NAND2_X1 U13221 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n11212) );
  OAI211_X1 U13222 ( .C1(n15271), .C2(n10563), .A(n10562), .B(n11212), .ZN(
        n10568) );
  AOI211_X1 U13223 ( .C1(n10566), .C2(n10565), .A(n10564), .B(n15266), .ZN(
        n10567) );
  AOI211_X1 U13224 ( .C1(n15260), .C2(n10569), .A(n10568), .B(n10567), .ZN(
        n10570) );
  INV_X1 U13225 ( .A(n10570), .ZN(P1_U3248) );
  INV_X1 U13226 ( .A(n13640), .ZN(n13648) );
  OAI222_X1 U13227 ( .A1(n13382), .A2(n10572), .B1(n12850), .B2(n10571), .C1(
        n13648), .C2(P3_U3151), .ZN(P3_U3279) );
  XNOR2_X1 U13228 ( .A(n10574), .B(n10573), .ZN(n10575) );
  NAND2_X1 U13229 ( .A1(n10575), .A2(n14103), .ZN(n10580) );
  OAI22_X1 U13230 ( .A1(n10577), .A2(n14325), .B1(n10576), .B2(n14323), .ZN(
        n10750) );
  AOI22_X1 U13231 ( .A1(n10578), .A2(P2_REG3_REG_1__SCAN_IN), .B1(n10750), 
        .B2(n14131), .ZN(n10579) );
  OAI211_X1 U13232 ( .C1(n15502), .C2(n14102), .A(n10580), .B(n10579), .ZN(
        P2_U3194) );
  INV_X1 U13233 ( .A(n10581), .ZN(n10584) );
  INV_X1 U13234 ( .A(n15433), .ZN(n10582) );
  OAI222_X1 U13235 ( .A1(n12959), .A2(n10583), .B1(n14531), .B2(n10584), .C1(
        P2_U3088), .C2(n10582), .ZN(P2_U3317) );
  INV_X1 U13236 ( .A(n11054), .ZN(n11051) );
  OAI222_X1 U13237 ( .A1(n12476), .A2(n10585), .B1(n13377), .B2(n10584), .C1(
        P1_U3086), .C2(n11051), .ZN(P1_U3345) );
  INV_X1 U13238 ( .A(n10697), .ZN(n10586) );
  NAND2_X1 U13239 ( .A1(n14663), .A2(n10586), .ZN(n10588) );
  NAND2_X1 U13240 ( .A1(n10590), .A2(n10821), .ZN(n10587) );
  AND2_X1 U13241 ( .A1(n10588), .A2(n10587), .ZN(n10595) );
  NAND2_X1 U13242 ( .A1(n6680), .A2(n10590), .ZN(n10592) );
  NAND2_X1 U13243 ( .A1(n14663), .A2(n10821), .ZN(n10591) );
  NAND2_X1 U13244 ( .A1(n10592), .A2(n10591), .ZN(n10593) );
  NAND2_X1 U13245 ( .A1(n10595), .A2(n10594), .ZN(n10691) );
  INV_X1 U13246 ( .A(n10594), .ZN(n10597) );
  NAND2_X1 U13247 ( .A1(n10597), .A2(n10596), .ZN(n10598) );
  NAND2_X1 U13248 ( .A1(n10691), .A2(n10598), .ZN(n10602) );
  AOI21_X1 U13249 ( .B1(n10602), .B2(n10601), .A(n10693), .ZN(n10607) );
  INV_X1 U13250 ( .A(n14587), .ZN(n15206) );
  AND2_X1 U13251 ( .A1(n15183), .A2(n14975), .ZN(n14615) );
  AOI22_X1 U13252 ( .A1(n14615), .A2(n14662), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n10701), .ZN(n10604) );
  OAI21_X1 U13253 ( .B1(n10603), .B2(n15206), .A(n10604), .ZN(n10605) );
  AOI21_X1 U13254 ( .B1(n15218), .B2(n10590), .A(n10605), .ZN(n10606) );
  OAI21_X1 U13255 ( .B1(n10607), .B2(n15212), .A(n10606), .ZN(P1_U3222) );
  INV_X1 U13256 ( .A(n14035), .ZN(n10608) );
  NOR2_X1 U13257 ( .A1(n10608), .A2(n9348), .ZN(n10610) );
  INV_X1 U13258 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10609) );
  NOR2_X1 U13259 ( .A1(n10628), .A2(n10609), .ZN(P3_U3262) );
  INV_X1 U13260 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10611) );
  NOR2_X1 U13261 ( .A1(n10628), .A2(n10611), .ZN(P3_U3261) );
  INV_X1 U13262 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10612) );
  NOR2_X1 U13263 ( .A1(n10610), .A2(n10612), .ZN(P3_U3260) );
  INV_X1 U13264 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10613) );
  NOR2_X1 U13265 ( .A1(n10628), .A2(n10613), .ZN(P3_U3259) );
  INV_X1 U13266 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10614) );
  NOR2_X1 U13267 ( .A1(n10610), .A2(n10614), .ZN(P3_U3258) );
  INV_X1 U13268 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10615) );
  NOR2_X1 U13269 ( .A1(n10628), .A2(n10615), .ZN(P3_U3257) );
  INV_X1 U13270 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10616) );
  NOR2_X1 U13271 ( .A1(n10628), .A2(n10616), .ZN(P3_U3256) );
  INV_X1 U13272 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10617) );
  NOR2_X1 U13273 ( .A1(n10628), .A2(n10617), .ZN(P3_U3255) );
  INV_X1 U13274 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10618) );
  NOR2_X1 U13275 ( .A1(n10628), .A2(n10618), .ZN(P3_U3254) );
  INV_X1 U13276 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n10619) );
  NOR2_X1 U13277 ( .A1(n10628), .A2(n10619), .ZN(P3_U3253) );
  INV_X1 U13278 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10620) );
  NOR2_X1 U13279 ( .A1(n10628), .A2(n10620), .ZN(P3_U3263) );
  INV_X1 U13280 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10621) );
  NOR2_X1 U13281 ( .A1(n10628), .A2(n10621), .ZN(P3_U3252) );
  INV_X1 U13282 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10622) );
  NOR2_X1 U13283 ( .A1(n10628), .A2(n10622), .ZN(P3_U3251) );
  INV_X1 U13284 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10623) );
  NOR2_X1 U13285 ( .A1(n10628), .A2(n10623), .ZN(P3_U3250) );
  INV_X1 U13286 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10624) );
  NOR2_X1 U13287 ( .A1(n10628), .A2(n10624), .ZN(P3_U3249) );
  INV_X1 U13288 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10625) );
  NOR2_X1 U13289 ( .A1(n10628), .A2(n10625), .ZN(P3_U3248) );
  INV_X1 U13290 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10626) );
  NOR2_X1 U13291 ( .A1(n10628), .A2(n10626), .ZN(P3_U3247) );
  INV_X1 U13292 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10627) );
  NOR2_X1 U13293 ( .A1(n10628), .A2(n10627), .ZN(P3_U3246) );
  INV_X1 U13294 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10629) );
  NOR2_X1 U13295 ( .A1(n10610), .A2(n10629), .ZN(P3_U3245) );
  INV_X1 U13296 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10630) );
  NOR2_X1 U13297 ( .A1(n10610), .A2(n10630), .ZN(P3_U3244) );
  INV_X1 U13298 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10631) );
  NOR2_X1 U13299 ( .A1(n10610), .A2(n10631), .ZN(P3_U3243) );
  INV_X1 U13300 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n10632) );
  NOR2_X1 U13301 ( .A1(n10610), .A2(n10632), .ZN(P3_U3234) );
  INV_X1 U13302 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10633) );
  NOR2_X1 U13303 ( .A1(n10610), .A2(n10633), .ZN(P3_U3241) );
  INV_X1 U13304 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10634) );
  NOR2_X1 U13305 ( .A1(n10610), .A2(n10634), .ZN(P3_U3242) );
  INV_X1 U13306 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10635) );
  NOR2_X1 U13307 ( .A1(n10610), .A2(n10635), .ZN(P3_U3239) );
  INV_X1 U13308 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10636) );
  NOR2_X1 U13309 ( .A1(n10610), .A2(n10636), .ZN(P3_U3235) );
  INV_X1 U13310 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10637) );
  NOR2_X1 U13311 ( .A1(n10610), .A2(n10637), .ZN(P3_U3237) );
  INV_X1 U13312 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10638) );
  NOR2_X1 U13313 ( .A1(n10628), .A2(n10638), .ZN(P3_U3240) );
  INV_X1 U13314 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10639) );
  NOR2_X1 U13315 ( .A1(n10628), .A2(n10639), .ZN(P3_U3238) );
  INV_X1 U13316 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10640) );
  NOR2_X1 U13317 ( .A1(n10628), .A2(n10640), .ZN(P3_U3236) );
  MUX2_X1 U13318 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10643), .S(n10727), .Z(
        n10644) );
  OAI21_X1 U13319 ( .B1(n10645), .B2(n10644), .A(n10726), .ZN(n10656) );
  NOR2_X1 U13320 ( .A1(n10646), .A2(n11487), .ZN(n10648) );
  MUX2_X1 U13321 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n11609), .S(n10727), .Z(
        n10647) );
  OAI21_X1 U13322 ( .B1(n10649), .B2(n10648), .A(n10647), .ZN(n10723) );
  INV_X1 U13323 ( .A(n10723), .ZN(n10651) );
  NOR3_X1 U13324 ( .A1(n10649), .A2(n10648), .A3(n10647), .ZN(n10650) );
  NOR3_X1 U13325 ( .A1(n10651), .A2(n10650), .A3(n15266), .ZN(n10655) );
  AND2_X1 U13326 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n11929) );
  AOI21_X1 U13327 ( .B1(n14737), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n11929), .ZN(
        n10652) );
  OAI21_X1 U13328 ( .B1(n10653), .B2(n14757), .A(n10652), .ZN(n10654) );
  AOI211_X1 U13329 ( .C1(n10656), .C2(n15260), .A(n10655), .B(n10654), .ZN(
        n10657) );
  INV_X1 U13330 ( .A(n10657), .ZN(P1_U3251) );
  XOR2_X1 U13331 ( .A(n10659), .B(n10658), .Z(n10664) );
  INV_X1 U13332 ( .A(n14131), .ZN(n14096) );
  AOI22_X1 U13333 ( .A1(n14368), .A2(n14170), .B1(n14167), .B2(n14369), .ZN(
        n10810) );
  INV_X1 U13334 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10660) );
  OAI22_X1 U13335 ( .A1(n14096), .A2(n10810), .B1(n10661), .B2(n10660), .ZN(
        n10662) );
  AOI21_X1 U13336 ( .B1(n10812), .B2(n14146), .A(n10662), .ZN(n10663) );
  OAI21_X1 U13337 ( .B1(n10664), .B2(n14148), .A(n10663), .ZN(P2_U3209) );
  NAND2_X1 U13338 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14671) );
  MUX2_X1 U13339 ( .A(n14671), .B(n10665), .S(n10214), .Z(n10669) );
  NAND2_X1 U13340 ( .A1(n10667), .A2(n10666), .ZN(n10668) );
  OAI211_X1 U13341 ( .C1(n10669), .C2(n12993), .A(P1_U4016), .B(n10668), .ZN(
        n14693) );
  XOR2_X1 U13342 ( .A(n10671), .B(n10670), .Z(n10679) );
  NAND2_X1 U13343 ( .A1(n14737), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n10672) );
  NAND2_X1 U13344 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n11335) );
  OAI211_X1 U13345 ( .C1(n14757), .C2(n10673), .A(n10672), .B(n11335), .ZN(
        n10678) );
  AOI211_X1 U13346 ( .C1(n10676), .C2(n10675), .A(n10674), .B(n14759), .ZN(
        n10677) );
  AOI211_X1 U13347 ( .C1(n14762), .C2(n10679), .A(n10678), .B(n10677), .ZN(
        n10680) );
  NAND2_X1 U13348 ( .A1(n14693), .A2(n10680), .ZN(P1_U3247) );
  INV_X1 U13349 ( .A(n10681), .ZN(n10683) );
  INV_X1 U13350 ( .A(n11536), .ZN(n11306) );
  OAI222_X1 U13351 ( .A1(n12959), .A2(n10682), .B1(n14531), .B2(n10683), .C1(
        P2_U3088), .C2(n11306), .ZN(P2_U3316) );
  INV_X1 U13352 ( .A(n11420), .ZN(n11415) );
  OAI222_X1 U13353 ( .A1(n12476), .A2(n10684), .B1(n13377), .B2(n10683), .C1(
        P1_U3086), .C2(n11415), .ZN(P1_U3344) );
  AOI21_X1 U13354 ( .B1(n14395), .B2(n10234), .A(n10716), .ZN(n10686) );
  NOR2_X1 U13355 ( .A1(n10686), .A2(n10685), .ZN(n10711) );
  OAI211_X1 U13356 ( .C1(n10716), .C2(n14434), .A(n10711), .B(n10712), .ZN(
        n11155) );
  NAND2_X1 U13357 ( .A1(n11155), .A2(n15550), .ZN(n10687) );
  OAI21_X1 U13358 ( .B1(n15550), .B2(n10545), .A(n10687), .ZN(P2_U3499) );
  INV_X1 U13359 ( .A(n10688), .ZN(n10690) );
  INV_X1 U13360 ( .A(SI_17_), .ZN(n10689) );
  OAI222_X1 U13361 ( .A1(n13649), .A2(P3_U3151), .B1(n12850), .B2(n10690), 
        .C1(n10689), .C2(n13382), .ZN(P3_U3278) );
  INV_X1 U13362 ( .A(n10691), .ZN(n10692) );
  NAND2_X1 U13363 ( .A1(n14662), .A2(n10821), .ZN(n10695) );
  NAND2_X1 U13364 ( .A1(n6680), .A2(n12589), .ZN(n10694) );
  NAND2_X1 U13365 ( .A1(n10695), .A2(n10694), .ZN(n10696) );
  XNOR2_X1 U13366 ( .A(n10696), .B(n13115), .ZN(n10819) );
  OAI22_X1 U13367 ( .A1(n7742), .A2(n13112), .B1(n15301), .B2(n6681), .ZN(
        n10818) );
  XNOR2_X1 U13368 ( .A(n10819), .B(n10818), .ZN(n10698) );
  NOR2_X1 U13369 ( .A1(n10699), .A2(n10698), .ZN(n10820) );
  AOI21_X1 U13370 ( .B1(n10699), .B2(n10698), .A(n10820), .ZN(n10704) );
  INV_X1 U13371 ( .A(n14661), .ZN(n10700) );
  OAI22_X1 U13372 ( .A1(n6865), .A2(n14869), .B1(n10700), .B2(n14871), .ZN(
        n11584) );
  AOI22_X1 U13373 ( .A1(n11584), .A2(n15183), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n10701), .ZN(n10703) );
  NAND2_X1 U13374 ( .A1(n15218), .A2(n12589), .ZN(n10702) );
  OAI211_X1 U13375 ( .C1(n10704), .C2(n15212), .A(n10703), .B(n10702), .ZN(
        P1_U3237) );
  INV_X1 U13376 ( .A(n10705), .ZN(n10708) );
  INV_X1 U13377 ( .A(n10706), .ZN(n10707) );
  NAND4_X1 U13378 ( .A1(n10708), .A2(n10707), .A3(n15512), .A4(n15511), .ZN(
        n10709) );
  NAND2_X1 U13379 ( .A1(n11007), .A2(n10710), .ZN(n10997) );
  NOR2_X1 U13380 ( .A1(n6677), .A2(n10997), .ZN(n14295) );
  INV_X1 U13381 ( .A(n14295), .ZN(n14381) );
  OAI21_X1 U13382 ( .B1(n8741), .B2(n10712), .A(n10711), .ZN(n10713) );
  NAND2_X1 U13383 ( .A1(n10713), .A2(n14397), .ZN(n10715) );
  INV_X2 U13384 ( .A(n14387), .ZN(n15499) );
  AOI22_X1 U13385 ( .A1(n6677), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(n15499), .ZN(n10714) );
  OAI211_X1 U13386 ( .C1(n10716), .C2(n14381), .A(n10715), .B(n10714), .ZN(
        P2_U3265) );
  NAND2_X1 U13387 ( .A1(n9273), .A2(P3_U3897), .ZN(n10717) );
  OAI21_X1 U13388 ( .B1(n6678), .B2(n10718), .A(n10717), .ZN(P3_U3493) );
  NAND2_X1 U13389 ( .A1(n6679), .A2(n6678), .ZN(n10719) );
  OAI21_X1 U13390 ( .B1(n6678), .B2(n10720), .A(n10719), .ZN(P3_U3494) );
  NAND2_X1 U13391 ( .A1(n10727), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10722) );
  MUX2_X1 U13392 ( .A(n11439), .B(P1_REG2_REG_9__SCAN_IN), .S(n10909), .Z(
        n10721) );
  NAND3_X1 U13393 ( .A1(n10723), .A2(n10722), .A3(n10721), .ZN(n10724) );
  NAND2_X1 U13394 ( .A1(n10724), .A2(n14762), .ZN(n10735) );
  MUX2_X1 U13395 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10725), .S(n10909), .Z(
        n10729) );
  OAI21_X1 U13396 ( .B1(n10727), .B2(P1_REG1_REG_8__SCAN_IN), .A(n10726), .ZN(
        n10728) );
  NAND2_X1 U13397 ( .A1(n10728), .A2(n10729), .ZN(n10908) );
  OAI21_X1 U13398 ( .B1(n10729), .B2(n10728), .A(n10908), .ZN(n10730) );
  NAND2_X1 U13399 ( .A1(n10730), .A2(n15260), .ZN(n10734) );
  NAND2_X1 U13400 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n12096) );
  INV_X1 U13401 ( .A(n12096), .ZN(n10732) );
  NOR2_X1 U13402 ( .A1(n14757), .A2(n10912), .ZN(n10731) );
  AOI211_X1 U13403 ( .C1(n14737), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n10732), .B(
        n10731), .ZN(n10733) );
  OAI211_X1 U13404 ( .C1(n10916), .C2(n10735), .A(n10734), .B(n10733), .ZN(
        P1_U3252) );
  INV_X1 U13405 ( .A(n10736), .ZN(n10763) );
  AOI22_X1 U13406 ( .A1(n11712), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n12964), .ZN(n10737) );
  OAI21_X1 U13407 ( .B1(n10763), .B2(n13377), .A(n10737), .ZN(P1_U3343) );
  INV_X1 U13408 ( .A(n13664), .ZN(n13672) );
  OAI222_X1 U13409 ( .A1(P3_U3151), .A2(n13672), .B1(n13382), .B2(n10739), 
        .C1(n12850), .C2(n10738), .ZN(P3_U3277) );
  NAND2_X1 U13410 ( .A1(n13532), .A2(P3_DATAO_REG_21__SCAN_IN), .ZN(n10740) );
  OAI21_X1 U13411 ( .B1(n13801), .B2(n13532), .A(n10740), .ZN(P3_U3512) );
  NAND2_X1 U13412 ( .A1(n11949), .A2(n6678), .ZN(n10741) );
  OAI21_X1 U13413 ( .B1(n6678), .B2(n10742), .A(n10741), .ZN(P3_U3496) );
  NAND2_X1 U13414 ( .A1(n10743), .A2(n10749), .ZN(n10744) );
  NAND2_X1 U13415 ( .A1(n10745), .A2(n10744), .ZN(n15495) );
  AOI21_X1 U13416 ( .B1(n10753), .B2(n10746), .A(n12878), .ZN(n10747) );
  AND2_X1 U13417 ( .A1(n10807), .A2(n10747), .ZN(n15497) );
  XNOR2_X1 U13418 ( .A(n10749), .B(n10748), .ZN(n10751) );
  AOI21_X1 U13419 ( .B1(n10751), .B2(n14358), .A(n10750), .ZN(n15507) );
  INV_X1 U13420 ( .A(n15507), .ZN(n10752) );
  AOI211_X1 U13421 ( .C1(n15520), .C2(n15495), .A(n15497), .B(n10752), .ZN(
        n11471) );
  INV_X1 U13422 ( .A(n14472), .ZN(n14407) );
  AOI22_X1 U13423 ( .A1(n14407), .A2(n10753), .B1(n15548), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n10754) );
  OAI21_X1 U13424 ( .B1(n11471), .B2(n15548), .A(n10754), .ZN(P2_U3500) );
  NAND2_X1 U13425 ( .A1(n13878), .A2(n6678), .ZN(n10755) );
  OAI21_X1 U13426 ( .B1(n6678), .B2(n10756), .A(n10755), .ZN(P3_U3506) );
  NAND2_X1 U13427 ( .A1(n8859), .A2(n6678), .ZN(n10757) );
  OAI21_X1 U13428 ( .B1(n6678), .B2(n10758), .A(n10757), .ZN(P3_U3495) );
  NAND2_X1 U13429 ( .A1(n13879), .A2(n6678), .ZN(n10759) );
  OAI21_X1 U13430 ( .B1(n6678), .B2(n10760), .A(n10759), .ZN(P3_U3504) );
  NAND2_X1 U13431 ( .A1(n13842), .A2(n6678), .ZN(n10761) );
  OAI21_X1 U13432 ( .B1(n6678), .B2(n10762), .A(n10761), .ZN(P3_U3509) );
  INV_X1 U13433 ( .A(n11975), .ZN(n11540) );
  OAI222_X1 U13434 ( .A1(n12959), .A2(n10764), .B1(n14531), .B2(n10763), .C1(
        n11540), .C2(P2_U3088), .ZN(P2_U3315) );
  NAND2_X1 U13435 ( .A1(n10765), .A2(P3_U3897), .ZN(n10766) );
  OAI21_X1 U13436 ( .B1(n6678), .B2(n10767), .A(n10766), .ZN(P3_U3498) );
  XNOR2_X1 U13437 ( .A(n10768), .B(n10771), .ZN(n10775) );
  OAI21_X1 U13438 ( .B1(n10771), .B2(n10770), .A(n10769), .ZN(n10772) );
  INV_X1 U13439 ( .A(n11145), .ZN(n14980) );
  NAND2_X1 U13440 ( .A1(n10772), .A2(n14980), .ZN(n10774) );
  AOI22_X1 U13441 ( .A1(n14975), .A2(n14660), .B1(n14662), .B2(n14974), .ZN(
        n10773) );
  OAI211_X1 U13442 ( .C1(n15286), .C2(n10775), .A(n10774), .B(n10773), .ZN(
        n11310) );
  INV_X1 U13443 ( .A(n11310), .ZN(n10777) );
  AOI21_X1 U13444 ( .B1(n11589), .B2(n12593), .A(n14958), .ZN(n10776) );
  NAND2_X1 U13445 ( .A1(n10776), .A2(n10836), .ZN(n11315) );
  NAND2_X1 U13446 ( .A1(n10777), .A2(n11315), .ZN(n10782) );
  OAI22_X1 U13447 ( .A1(n15089), .A2(n7755), .B1(n15324), .B2(n7745), .ZN(
        n10778) );
  AOI21_X1 U13448 ( .B1(n10782), .B2(n15324), .A(n10778), .ZN(n10779) );
  INV_X1 U13449 ( .A(n10779), .ZN(P1_U3468) );
  INV_X1 U13450 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10780) );
  OAI22_X1 U13451 ( .A1(n15046), .A2(n7755), .B1(n15332), .B2(n10780), .ZN(
        n10781) );
  AOI21_X1 U13452 ( .B1(n10782), .B2(n15332), .A(n10781), .ZN(n10783) );
  INV_X1 U13453 ( .A(n10783), .ZN(P1_U3531) );
  OAI222_X1 U13454 ( .A1(n12850), .A2(n10785), .B1(n13382), .B2(n10784), .C1(
        P3_U3151), .C2(n13679), .ZN(P3_U3276) );
  NAND2_X1 U13455 ( .A1(n12923), .A2(n6678), .ZN(n10786) );
  OAI21_X1 U13456 ( .B1(P3_U3897), .B2(n10787), .A(n10786), .ZN(P3_U3510) );
  NAND2_X1 U13457 ( .A1(n13483), .A2(P3_U3897), .ZN(n10788) );
  OAI21_X1 U13458 ( .B1(n6678), .B2(n10789), .A(n10788), .ZN(P3_U3503) );
  NAND2_X1 U13459 ( .A1(n13852), .A2(n6678), .ZN(n10790) );
  OAI21_X1 U13460 ( .B1(n6678), .B2(n10791), .A(n10790), .ZN(P3_U3508) );
  OAI21_X1 U13461 ( .B1(n10794), .B2(n10793), .A(n10792), .ZN(n10801) );
  NAND2_X1 U13462 ( .A1(n14165), .A2(n14369), .ZN(n10796) );
  NAND2_X1 U13463 ( .A1(n14167), .A2(n14368), .ZN(n10795) );
  AND2_X1 U13464 ( .A1(n10796), .A2(n10795), .ZN(n11001) );
  INV_X1 U13465 ( .A(n11001), .ZN(n10797) );
  AOI22_X1 U13466 ( .A1(n14131), .A2(n10797), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10799) );
  NAND2_X1 U13467 ( .A1(n14146), .A2(n11019), .ZN(n10798) );
  OAI211_X1 U13468 ( .C1(n14140), .C2(n11009), .A(n10799), .B(n10798), .ZN(
        n10800) );
  AOI21_X1 U13469 ( .B1(n10801), .B2(n14103), .A(n10800), .ZN(n10802) );
  INV_X1 U13470 ( .A(n10802), .ZN(P2_U3202) );
  NAND2_X1 U13471 ( .A1(n13812), .A2(n6678), .ZN(n10803) );
  OAI21_X1 U13472 ( .B1(P3_U3897), .B2(n10804), .A(n10803), .ZN(P3_U3511) );
  OAI21_X1 U13473 ( .B1(n10806), .B2(n10809), .A(n10805), .ZN(n11042) );
  AOI211_X1 U13474 ( .C1(n10812), .C2(n10807), .A(n12878), .B(n10848), .ZN(
        n11038) );
  XNOR2_X1 U13475 ( .A(n10809), .B(n10808), .ZN(n10811) );
  OAI21_X1 U13476 ( .B1(n10811), .B2(n14395), .A(n10810), .ZN(n11037) );
  AOI211_X1 U13477 ( .C1(n15520), .C2(n11042), .A(n11038), .B(n11037), .ZN(
        n11475) );
  AOI22_X1 U13478 ( .A1(n14407), .A2(n10812), .B1(n15548), .B2(
        P2_REG1_REG_2__SCAN_IN), .ZN(n10813) );
  OAI21_X1 U13479 ( .B1(n11475), .B2(n15548), .A(n10813), .ZN(P2_U3501) );
  INV_X1 U13480 ( .A(n12217), .ZN(n11983) );
  INV_X1 U13481 ( .A(n10814), .ZN(n10816) );
  INV_X1 U13482 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10815) );
  OAI222_X1 U13483 ( .A1(P2_U3088), .A2(n11983), .B1(n12957), .B2(n10816), 
        .C1(n10815), .C2(n12959), .ZN(P2_U3314) );
  OAI222_X1 U13484 ( .A1(n12476), .A2(n10817), .B1(n13377), .B2(n10816), .C1(
        n11756), .C2(P1_U3086), .ZN(P1_U3342) );
  AOI22_X1 U13485 ( .A1(n14661), .A2(n13068), .B1(n13103), .B2(n12593), .ZN(
        n11190) );
  AOI22_X1 U13486 ( .A1(n14661), .A2(n13103), .B1(n13102), .B2(n12593), .ZN(
        n10822) );
  XNOR2_X1 U13487 ( .A(n10822), .B(n13115), .ZN(n11189) );
  OAI211_X1 U13488 ( .C1(n10824), .C2(n10823), .A(n11193), .B(n15179), .ZN(
        n10832) );
  INV_X1 U13489 ( .A(n10825), .ZN(n10826) );
  NAND2_X1 U13490 ( .A1(n10827), .A2(n10826), .ZN(n10828) );
  INV_X1 U13491 ( .A(n15222), .ZN(n14636) );
  MUX2_X1 U13492 ( .A(n14636), .B(P1_U3086), .S(P1_REG3_REG_3__SCAN_IN), .Z(
        n10830) );
  OAI22_X1 U13493 ( .A1(n11197), .A2(n15205), .B1(n15206), .B2(n7742), .ZN(
        n10829) );
  AOI211_X1 U13494 ( .C1(n15218), .C2(n12593), .A(n10830), .B(n10829), .ZN(
        n10831) );
  NAND2_X1 U13495 ( .A1(n10832), .A2(n10831), .ZN(P1_U3218) );
  XNOR2_X1 U13496 ( .A(n10833), .B(n12780), .ZN(n11265) );
  OAI21_X1 U13497 ( .B1(n10835), .B2(n12780), .A(n10834), .ZN(n11263) );
  AOI211_X1 U13498 ( .C1(n12599), .C2(n10836), .A(n14958), .B(n10926), .ZN(
        n11256) );
  NAND2_X1 U13499 ( .A1(n14661), .A2(n14974), .ZN(n10838) );
  NAND2_X1 U13500 ( .A1(n14659), .A2(n14975), .ZN(n10837) );
  NAND2_X1 U13501 ( .A1(n10838), .A2(n10837), .ZN(n11333) );
  AOI211_X1 U13502 ( .C1(n11263), .C2(n15321), .A(n11256), .B(n11333), .ZN(
        n10839) );
  OAI21_X1 U13503 ( .B1(n15286), .B2(n11265), .A(n10839), .ZN(n10844) );
  OAI22_X1 U13504 ( .A1(n15089), .A2(n11261), .B1(n15324), .B2(n7762), .ZN(
        n10840) );
  AOI21_X1 U13505 ( .B1(n10844), .B2(n15324), .A(n10840), .ZN(n10841) );
  INV_X1 U13506 ( .A(n10841), .ZN(P1_U3471) );
  INV_X1 U13507 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10842) );
  OAI22_X1 U13508 ( .A1(n15046), .A2(n11261), .B1(n15332), .B2(n10842), .ZN(
        n10843) );
  AOI21_X1 U13509 ( .B1(n10844), .B2(n15332), .A(n10843), .ZN(n10845) );
  INV_X1 U13510 ( .A(n10845), .ZN(P1_U3532) );
  OAI21_X1 U13511 ( .B1(n10847), .B2(n10851), .A(n10846), .ZN(n11034) );
  INV_X1 U13512 ( .A(n10848), .ZN(n10849) );
  AOI211_X1 U13513 ( .C1(n10905), .C2(n10849), .A(n12878), .B(n11004), .ZN(
        n11029) );
  XNOR2_X1 U13514 ( .A(n10851), .B(n10850), .ZN(n10852) );
  AOI22_X1 U13515 ( .A1(n14368), .A2(n14169), .B1(n14166), .B2(n14369), .ZN(
        n10896) );
  OAI21_X1 U13516 ( .B1(n10852), .B2(n14395), .A(n10896), .ZN(n11028) );
  AOI211_X1 U13517 ( .C1(n15520), .C2(n11034), .A(n11029), .B(n11028), .ZN(
        n11467) );
  AOI22_X1 U13518 ( .A1(n14407), .A2(n10905), .B1(n15548), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n10853) );
  OAI21_X1 U13519 ( .B1(n11467), .B2(n15548), .A(n10853), .ZN(P2_U3502) );
  OR2_X1 U13520 ( .A1(n10855), .A2(P3_U3151), .ZN(n13359) );
  INV_X1 U13521 ( .A(n13359), .ZN(n10854) );
  OR2_X1 U13522 ( .A1(n11118), .A2(n10854), .ZN(n10868) );
  NAND2_X1 U13523 ( .A1(n13305), .A2(n10855), .ZN(n10857) );
  NAND2_X1 U13524 ( .A1(n10868), .A2(n10866), .ZN(n10869) );
  MUX2_X1 U13525 ( .A(n13532), .B(n10869), .S(n13354), .Z(n15671) );
  AND2_X1 U13526 ( .A1(P3_U3897), .A2(n13354), .ZN(n15666) );
  INV_X1 U13527 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10859) );
  INV_X1 U13528 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10858) );
  MUX2_X1 U13529 ( .A(n10859), .B(n10858), .S(n13667), .Z(n11223) );
  MUX2_X1 U13530 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n13667), .Z(n10860) );
  NOR2_X1 U13531 ( .A1(n10860), .A2(n10881), .ZN(n10950) );
  AOI21_X1 U13532 ( .B1(n10860), .B2(n10881), .A(n10950), .ZN(n10861) );
  NAND2_X1 U13533 ( .A1(n10861), .A2(n11217), .ZN(n10957) );
  OAI21_X1 U13534 ( .B1(n11217), .B2(n10861), .A(n10957), .ZN(n10879) );
  NAND2_X1 U13535 ( .A1(n10943), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10862) );
  NOR2_X1 U13536 ( .A1(n10863), .A2(n11678), .ZN(n10942) );
  AND2_X1 U13537 ( .A1(n10863), .A2(n11678), .ZN(n10865) );
  INV_X1 U13538 ( .A(n15681), .ZN(n13655) );
  OAI21_X1 U13539 ( .B1(n10942), .B2(n10865), .A(n13655), .ZN(n10877) );
  INV_X1 U13540 ( .A(n10866), .ZN(n10867) );
  AOI22_X1 U13541 ( .A1(n15674), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10876) );
  OR2_X1 U13542 ( .A1(n10869), .A2(n13590), .ZN(n15583) );
  INV_X1 U13543 ( .A(n11218), .ZN(n10939) );
  OR2_X1 U13544 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10939), .ZN(n10870) );
  OAI21_X1 U13545 ( .B1(n10881), .B2(n11218), .A(n10870), .ZN(n10872) );
  INV_X1 U13546 ( .A(n10872), .ZN(n10873) );
  OAI21_X1 U13547 ( .B1(n10873), .B2(P3_REG1_REG_1__SCAN_IN), .A(n10938), .ZN(
        n10874) );
  NAND2_X1 U13548 ( .A1(n15677), .A2(n10874), .ZN(n10875) );
  NAND3_X1 U13549 ( .A1(n10877), .A2(n10876), .A3(n10875), .ZN(n10878) );
  AOI21_X1 U13550 ( .B1(n15666), .B2(n10879), .A(n10878), .ZN(n10880) );
  OAI21_X1 U13551 ( .B1(n10881), .B2(n15671), .A(n10880), .ZN(P3_U3183) );
  NAND2_X1 U13552 ( .A1(n9301), .A2(P3_U3897), .ZN(n10882) );
  OAI21_X1 U13553 ( .B1(n6678), .B2(n10883), .A(n10882), .ZN(P3_U3513) );
  OAI21_X1 U13554 ( .B1(n10886), .B2(n10885), .A(n10884), .ZN(n10887) );
  NAND2_X1 U13555 ( .A1(n10887), .A2(n14103), .ZN(n10894) );
  INV_X1 U13556 ( .A(n14140), .ZN(n14107) );
  NAND2_X1 U13557 ( .A1(n14164), .A2(n14369), .ZN(n10889) );
  NAND2_X1 U13558 ( .A1(n14166), .A2(n14368), .ZN(n10888) );
  NAND2_X1 U13559 ( .A1(n10889), .A2(n10888), .ZN(n11071) );
  NAND2_X1 U13560 ( .A1(n14131), .A2(n11071), .ZN(n10890) );
  OAI21_X1 U13561 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n10891), .A(n10890), .ZN(
        n10892) );
  AOI21_X1 U13562 ( .B1(n11125), .B2(n14107), .A(n10892), .ZN(n10893) );
  OAI211_X1 U13563 ( .C1(n11127), .C2(n14102), .A(n10894), .B(n10893), .ZN(
        P2_U3199) );
  MUX2_X1 U13564 ( .A(P2_STATE_REG_SCAN_IN), .B(n14140), .S(n11030), .Z(n10895) );
  OAI21_X1 U13565 ( .B1(n10896), .B2(n14096), .A(n10895), .ZN(n10904) );
  NAND2_X1 U13566 ( .A1(n10898), .A2(n10897), .ZN(n10902) );
  INV_X1 U13567 ( .A(n10899), .ZN(n10900) );
  AOI211_X1 U13568 ( .C1(n10902), .C2(n10901), .A(n14148), .B(n10900), .ZN(
        n10903) );
  AOI211_X1 U13569 ( .C1(n10905), .C2(n14146), .A(n10904), .B(n10903), .ZN(
        n10906) );
  INV_X1 U13570 ( .A(n10906), .ZN(P2_U3190) );
  INV_X1 U13571 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10907) );
  MUX2_X1 U13572 ( .A(n10907), .B(P1_REG1_REG_10__SCAN_IN), .S(n11054), .Z(
        n10911) );
  OAI21_X1 U13573 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n10909), .A(n10908), .ZN(
        n10910) );
  NOR2_X1 U13574 ( .A1(n10910), .A2(n10911), .ZN(n11053) );
  AOI211_X1 U13575 ( .C1(n10911), .C2(n10910), .A(n14759), .B(n11053), .ZN(
        n10923) );
  NOR2_X1 U13576 ( .A1(n10912), .A2(n11439), .ZN(n10915) );
  MUX2_X1 U13577 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n10913), .S(n11054), .Z(
        n10914) );
  OAI21_X1 U13578 ( .B1(n10916), .B2(n10915), .A(n10914), .ZN(n11050) );
  OR3_X1 U13579 ( .A1(n10916), .A2(n10915), .A3(n10914), .ZN(n10917) );
  NAND3_X1 U13580 ( .A1(n11050), .A2(n14762), .A3(n10917), .ZN(n10921) );
  NOR2_X1 U13581 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10918), .ZN(n10919) );
  AOI21_X1 U13582 ( .B1(n14737), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n10919), 
        .ZN(n10920) );
  OAI211_X1 U13583 ( .C1(n14757), .C2(n11051), .A(n10921), .B(n10920), .ZN(
        n10922) );
  OR2_X1 U13584 ( .A1(n10923), .A2(n10922), .ZN(P1_U3253) );
  OAI21_X1 U13585 ( .B1(n10925), .B2(n12781), .A(n10924), .ZN(n11146) );
  OAI21_X1 U13586 ( .B1(n10926), .B2(n11148), .A(n15049), .ZN(n10927) );
  NOR2_X1 U13587 ( .A1(n10927), .A2(n11549), .ZN(n11151) );
  XNOR2_X1 U13588 ( .A(n10928), .B(n12781), .ZN(n10932) );
  NAND2_X1 U13589 ( .A1(n14660), .A2(n14974), .ZN(n10930) );
  NAND2_X1 U13590 ( .A1(n14658), .A2(n14975), .ZN(n10929) );
  NAND2_X1 U13591 ( .A1(n10930), .A2(n10929), .ZN(n11210) );
  INV_X1 U13592 ( .A(n11210), .ZN(n10931) );
  OAI21_X1 U13593 ( .B1(n10932), .B2(n15286), .A(n10931), .ZN(n11144) );
  AOI211_X1 U13594 ( .C1(n11146), .C2(n15321), .A(n11151), .B(n11144), .ZN(
        n10937) );
  INV_X1 U13595 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10933) );
  OAI22_X1 U13596 ( .A1(n15089), .A2(n11148), .B1(n15324), .B2(n10933), .ZN(
        n10934) );
  INV_X1 U13597 ( .A(n10934), .ZN(n10935) );
  OAI21_X1 U13598 ( .B1(n10937), .B2(n10226), .A(n10935), .ZN(P1_U3474) );
  INV_X1 U13599 ( .A(n15046), .ZN(n12189) );
  AOI22_X1 U13600 ( .A1(n12189), .A2(n12608), .B1(n15330), .B2(
        P1_REG1_REG_5__SCAN_IN), .ZN(n10936) );
  OAI21_X1 U13601 ( .B1(n10937), .B2(n15330), .A(n10936), .ZN(P1_U3533) );
  INV_X1 U13602 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n11899) );
  MUX2_X1 U13603 ( .A(n11899), .B(P3_REG1_REG_2__SCAN_IN), .S(n11900), .Z(
        n10941) );
  NAND2_X1 U13604 ( .A1(n10941), .A2(n10940), .ZN(n11898) );
  OAI21_X1 U13605 ( .B1(n10941), .B2(n10940), .A(n11898), .ZN(n10949) );
  INV_X1 U13606 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10951) );
  XNOR2_X1 U13607 ( .A(n11900), .B(n10951), .ZN(n10945) );
  AOI21_X1 U13608 ( .B1(P3_REG2_REG_0__SCAN_IN), .B2(n10943), .A(n10942), .ZN(
        n10944) );
  NOR2_X1 U13609 ( .A1(n10944), .A2(n10945), .ZN(n11834) );
  AOI21_X1 U13610 ( .B1(n10945), .B2(n10944), .A(n11834), .ZN(n10946) );
  NOR2_X1 U13611 ( .A1(n15681), .A2(n10946), .ZN(n10948) );
  INV_X1 U13612 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n11187) );
  OAI22_X1 U13613 ( .A1(n15591), .A2(n9616), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11187), .ZN(n10947) );
  AOI211_X1 U13614 ( .C1(n15677), .C2(n10949), .A(n10948), .B(n10947), .ZN(
        n10960) );
  INV_X1 U13615 ( .A(n10950), .ZN(n10956) );
  MUX2_X1 U13616 ( .A(n10951), .B(n11899), .S(n13667), .Z(n10952) );
  NAND2_X1 U13617 ( .A1(n10952), .A2(n11900), .ZN(n11850) );
  INV_X1 U13618 ( .A(n10952), .ZN(n10953) );
  NAND2_X1 U13619 ( .A1(n10953), .A2(n11835), .ZN(n10954) );
  NAND2_X1 U13620 ( .A1(n11850), .A2(n10954), .ZN(n10955) );
  AND3_X1 U13621 ( .A1(n10957), .A2(n10956), .A3(n10955), .ZN(n10958) );
  OAI21_X1 U13622 ( .B1(n15557), .B2(n10958), .A(n15666), .ZN(n10959) );
  OAI211_X1 U13623 ( .C1(n15671), .C2(n11835), .A(n10960), .B(n10959), .ZN(
        P3_U3184) );
  INV_X1 U13624 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10961) );
  MUX2_X1 U13625 ( .A(n10961), .B(P2_REG1_REG_9__SCAN_IN), .S(n11295), .Z(
        n10976) );
  INV_X1 U13626 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10962) );
  AND2_X1 U13627 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n15335) );
  NAND2_X1 U13628 ( .A1(n15336), .A2(n15335), .ZN(n15334) );
  NAND2_X1 U13629 ( .A1(n15344), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10963) );
  NAND2_X1 U13630 ( .A1(n15334), .A2(n10963), .ZN(n14177) );
  INV_X1 U13631 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10964) );
  MUX2_X1 U13632 ( .A(n10964), .B(P2_REG1_REG_2__SCAN_IN), .S(n10978), .Z(
        n14178) );
  NAND2_X1 U13633 ( .A1(n14177), .A2(n14178), .ZN(n14176) );
  INV_X1 U13634 ( .A(n10978), .ZN(n14175) );
  NAND2_X1 U13635 ( .A1(n14175), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10965) );
  NAND2_X1 U13636 ( .A1(n14176), .A2(n10965), .ZN(n15348) );
  INV_X1 U13637 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10966) );
  MUX2_X1 U13638 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n10966), .S(n15356), .Z(
        n15349) );
  NAND2_X1 U13639 ( .A1(n15348), .A2(n15349), .ZN(n15347) );
  NAND2_X1 U13640 ( .A1(n15356), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10967) );
  NAND2_X1 U13641 ( .A1(n15347), .A2(n10967), .ZN(n15361) );
  INV_X1 U13642 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10968) );
  MUX2_X1 U13643 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n10968), .S(n15369), .Z(
        n15362) );
  NAND2_X1 U13644 ( .A1(n15361), .A2(n15362), .ZN(n15360) );
  NAND2_X1 U13645 ( .A1(n15369), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10969) );
  NAND2_X1 U13646 ( .A1(n15360), .A2(n10969), .ZN(n15374) );
  INV_X1 U13647 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n11077) );
  MUX2_X1 U13648 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n11077), .S(n15382), .Z(
        n15375) );
  NAND2_X1 U13649 ( .A1(n15374), .A2(n15375), .ZN(n15373) );
  NAND2_X1 U13650 ( .A1(n15382), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10970) );
  NAND2_X1 U13651 ( .A1(n15373), .A2(n10970), .ZN(n15386) );
  INV_X1 U13652 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n11690) );
  MUX2_X1 U13653 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n11690), .S(n15394), .Z(
        n15387) );
  NAND2_X1 U13654 ( .A1(n15386), .A2(n15387), .ZN(n15385) );
  NAND2_X1 U13655 ( .A1(n15394), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n10971) );
  NAND2_X1 U13656 ( .A1(n15385), .A2(n10971), .ZN(n15399) );
  INV_X1 U13657 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n15544) );
  MUX2_X1 U13658 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n15544), .S(n15407), .Z(
        n15400) );
  NAND2_X1 U13659 ( .A1(n15399), .A2(n15400), .ZN(n15398) );
  NAND2_X1 U13660 ( .A1(n15407), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10972) );
  NAND2_X1 U13661 ( .A1(n15398), .A2(n10972), .ZN(n15415) );
  INV_X1 U13662 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n15546) );
  MUX2_X1 U13663 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n15546), .S(n10984), .Z(
        n15416) );
  NAND2_X1 U13664 ( .A1(n15415), .A2(n15416), .ZN(n15414) );
  NAND2_X1 U13665 ( .A1(n10984), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10973) );
  NAND2_X1 U13666 ( .A1(n15414), .A2(n10973), .ZN(n10975) );
  OR2_X1 U13667 ( .A1(n10975), .A2(n10976), .ZN(n11297) );
  INV_X1 U13668 ( .A(n11297), .ZN(n10974) );
  AOI21_X1 U13669 ( .B1(n10976), .B2(n10975), .A(n10974), .ZN(n10994) );
  INV_X1 U13670 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10977) );
  AND3_X1 U13671 ( .A1(n15338), .A2(P2_IR_REG_0__SCAN_IN), .A3(
        P2_REG2_REG_0__SCAN_IN), .ZN(n15339) );
  INV_X1 U13672 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10979) );
  MUX2_X1 U13673 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10979), .S(n10978), .Z(
        n14172) );
  AOI21_X1 U13674 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n14175), .A(n14171), .ZN(
        n15353) );
  INV_X1 U13675 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10980) );
  MUX2_X1 U13676 ( .A(n10980), .B(P2_REG2_REG_3__SCAN_IN), .S(n15356), .Z(
        n15352) );
  AOI21_X1 U13677 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(n15356), .A(n15351), .ZN(
        n15366) );
  INV_X1 U13678 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10981) );
  MUX2_X1 U13679 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n10981), .S(n15369), .Z(
        n10982) );
  INV_X1 U13680 ( .A(n10982), .ZN(n15365) );
  INV_X1 U13681 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10983) );
  MUX2_X1 U13682 ( .A(n10983), .B(P2_REG2_REG_5__SCAN_IN), .S(n15382), .Z(
        n15378) );
  XNOR2_X1 U13683 ( .A(n15394), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n15390) );
  XNOR2_X1 U13684 ( .A(n15407), .B(P2_REG2_REG_7__SCAN_IN), .ZN(n15403) );
  XNOR2_X1 U13685 ( .A(n10984), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n15412) );
  INV_X1 U13686 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10985) );
  MUX2_X1 U13687 ( .A(n10985), .B(P2_REG2_REG_9__SCAN_IN), .S(n11295), .Z(
        n10986) );
  INV_X1 U13688 ( .A(n10986), .ZN(n10987) );
  OAI21_X1 U13689 ( .B1(n10988), .B2(n10987), .A(n11290), .ZN(n10992) );
  NAND2_X1 U13690 ( .A1(n15333), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n10989) );
  NAND2_X1 U13691 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n11452) );
  OAI211_X1 U13692 ( .C1(n15489), .C2(n10990), .A(n10989), .B(n11452), .ZN(
        n10991) );
  AOI21_X1 U13693 ( .B1(n10992), .B2(n15478), .A(n10991), .ZN(n10993) );
  OAI21_X1 U13694 ( .B1(n10994), .B2(n15465), .A(n10993), .ZN(P2_U3223) );
  OAI21_X1 U13695 ( .B1(n10996), .B2(n10999), .A(n10995), .ZN(n11018) );
  INV_X1 U13696 ( .A(n11018), .ZN(n11013) );
  NAND2_X1 U13697 ( .A1(n10234), .A2(n10997), .ZN(n10998) );
  NAND2_X1 U13698 ( .A1(n14397), .A2(n10998), .ZN(n14362) );
  XNOR2_X1 U13699 ( .A(n11000), .B(n10999), .ZN(n11002) );
  OAI21_X1 U13700 ( .B1(n11002), .B2(n14395), .A(n11001), .ZN(n11016) );
  INV_X1 U13701 ( .A(n11016), .ZN(n11003) );
  MUX2_X1 U13702 ( .A(n10981), .B(n11003), .S(n14397), .Z(n11012) );
  INV_X1 U13703 ( .A(n11004), .ZN(n11006) );
  INV_X1 U13704 ( .A(n11073), .ZN(n11005) );
  AOI211_X1 U13705 ( .C1(n11019), .C2(n11006), .A(n12878), .B(n11005), .ZN(
        n11017) );
  OAI22_X1 U13706 ( .A1(n15503), .A2(n11459), .B1(n11009), .B2(n14387), .ZN(
        n11010) );
  AOI21_X1 U13707 ( .B1(n11017), .B2(n15498), .A(n11010), .ZN(n11011) );
  OAI211_X1 U13708 ( .C1(n11013), .C2(n14362), .A(n11012), .B(n11011), .ZN(
        P2_U3261) );
  NAND2_X1 U13709 ( .A1(n6684), .A2(n6678), .ZN(n11014) );
  OAI21_X1 U13710 ( .B1(n6678), .B2(n11015), .A(n11014), .ZN(P3_U3514) );
  AOI211_X1 U13711 ( .C1(n15520), .C2(n11018), .A(n11017), .B(n11016), .ZN(
        n11462) );
  AOI22_X1 U13712 ( .A1(n14407), .A2(n11019), .B1(n15548), .B2(
        P2_REG1_REG_4__SCAN_IN), .ZN(n11020) );
  OAI21_X1 U13713 ( .B1(n11462), .B2(n15548), .A(n11020), .ZN(P2_U3503) );
  INV_X1 U13714 ( .A(n11021), .ZN(n11024) );
  INV_X1 U13715 ( .A(n15457), .ZN(n11022) );
  OAI222_X1 U13716 ( .A1(n12959), .A2(n11023), .B1(n12957), .B2(n11024), .C1(
        n11022), .C2(P2_U3088), .ZN(P2_U3311) );
  INV_X1 U13717 ( .A(n14716), .ZN(n14721) );
  OAI222_X1 U13718 ( .A1(n12476), .A2(n11025), .B1(n13377), .B2(n11024), .C1(
        n14721), .C2(P1_U3086), .ZN(P1_U3339) );
  OAI222_X1 U13719 ( .A1(n12850), .A2(n11027), .B1(n13382), .B2(n11026), .C1(
        P3_U3151), .C2(n11159), .ZN(P3_U3275) );
  INV_X1 U13720 ( .A(n11028), .ZN(n11036) );
  INV_X1 U13721 ( .A(n14362), .ZN(n15496) );
  NAND2_X1 U13722 ( .A1(n11029), .A2(n15498), .ZN(n11032) );
  AOI22_X1 U13723 ( .A1(n6677), .A2(P2_REG2_REG_3__SCAN_IN), .B1(n15499), .B2(
        n11030), .ZN(n11031) );
  OAI211_X1 U13724 ( .C1(n11464), .C2(n15503), .A(n11032), .B(n11031), .ZN(
        n11033) );
  AOI21_X1 U13725 ( .B1(n15496), .B2(n11034), .A(n11033), .ZN(n11035) );
  OAI21_X1 U13726 ( .B1(n11036), .B2(n6677), .A(n11035), .ZN(P2_U3262) );
  INV_X1 U13727 ( .A(n11037), .ZN(n11044) );
  NAND2_X1 U13728 ( .A1(n11038), .A2(n15498), .ZN(n11040) );
  AOI22_X1 U13729 ( .A1(n6677), .A2(P2_REG2_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(n15499), .ZN(n11039) );
  OAI211_X1 U13730 ( .C1(n8299), .C2(n15503), .A(n11040), .B(n11039), .ZN(
        n11041) );
  AOI21_X1 U13731 ( .B1(n15496), .B2(n11042), .A(n11041), .ZN(n11043) );
  OAI21_X1 U13732 ( .B1(n11044), .B2(n6677), .A(n11043), .ZN(P2_U3263) );
  INV_X1 U13733 ( .A(n11045), .ZN(n11047) );
  INV_X1 U13734 ( .A(n14184), .ZN(n12214) );
  OAI222_X1 U13735 ( .A1(n12959), .A2(n11046), .B1(n12957), .B2(n11047), .C1(
        n12214), .C2(P2_U3088), .ZN(P2_U3313) );
  INV_X1 U13736 ( .A(n14695), .ZN(n14705) );
  OAI222_X1 U13737 ( .A1(n12476), .A2(n11048), .B1(n13377), .B2(n11047), .C1(
        n14705), .C2(P1_U3086), .ZN(P1_U3341) );
  NAND2_X1 U13738 ( .A1(n11420), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n11049) );
  OAI21_X1 U13739 ( .B1(n11420), .B2(P1_REG2_REG_11__SCAN_IN), .A(n11049), 
        .ZN(n11411) );
  OAI21_X1 U13740 ( .B1(n10913), .B2(n11051), .A(n11050), .ZN(n11412) );
  XOR2_X1 U13741 ( .A(n11411), .B(n11412), .Z(n11062) );
  MUX2_X1 U13742 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n11052), .S(n11420), .Z(
        n11056) );
  OAI21_X1 U13743 ( .B1(n11056), .B2(n11055), .A(n11419), .ZN(n11057) );
  NAND2_X1 U13744 ( .A1(n11057), .A2(n15260), .ZN(n11061) );
  NAND2_X1 U13745 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n15219)
         );
  INV_X1 U13746 ( .A(n15219), .ZN(n11059) );
  NOR2_X1 U13747 ( .A1(n14757), .A2(n11415), .ZN(n11058) );
  AOI211_X1 U13748 ( .C1(n14737), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n11059), 
        .B(n11058), .ZN(n11060) );
  OAI211_X1 U13749 ( .C1(n11062), .C2(n15266), .A(n11061), .B(n11060), .ZN(
        P1_U3254) );
  INV_X1 U13750 ( .A(n11063), .ZN(n11066) );
  INV_X1 U13751 ( .A(n14733), .ZN(n14736) );
  OAI222_X1 U13752 ( .A1(n12476), .A2(n11064), .B1(n13377), .B2(n11066), .C1(
        n14736), .C2(P1_U3086), .ZN(P1_U3338) );
  INV_X1 U13753 ( .A(n15471), .ZN(n11065) );
  OAI222_X1 U13754 ( .A1(n12959), .A2(n11067), .B1(n12957), .B2(n11066), .C1(
        n11065), .C2(P2_U3088), .ZN(P2_U3310) );
  XNOR2_X1 U13755 ( .A(n11068), .B(n11070), .ZN(n11128) );
  XNOR2_X1 U13756 ( .A(n11069), .B(n11070), .ZN(n11072) );
  AOI21_X1 U13757 ( .B1(n11072), .B2(n14358), .A(n11071), .ZN(n11133) );
  AOI211_X1 U13758 ( .C1(n11074), .C2(n11073), .A(n12878), .B(n11324), .ZN(
        n11131) );
  AOI21_X1 U13759 ( .B1(n15532), .B2(n11074), .A(n11131), .ZN(n11075) );
  OAI211_X1 U13760 ( .C1(n11128), .C2(n14478), .A(n11133), .B(n11075), .ZN(
        n11134) );
  NAND2_X1 U13761 ( .A1(n11134), .A2(n15550), .ZN(n11076) );
  OAI21_X1 U13762 ( .B1(n15550), .B2(n11077), .A(n11076), .ZN(P2_U3504) );
  INV_X1 U13763 ( .A(n11078), .ZN(n11080) );
  OAI222_X1 U13764 ( .A1(n12959), .A2(n11079), .B1(n12957), .B2(n11080), .C1(
        n15437), .C2(P2_U3088), .ZN(P2_U3312) );
  INV_X1 U13765 ( .A(n15262), .ZN(n14707) );
  OAI222_X1 U13766 ( .A1(n12476), .A2(n11081), .B1(n13377), .B2(n11080), .C1(
        n14707), .C2(P1_U3086), .ZN(P1_U3340) );
  NAND2_X1 U13767 ( .A1(n13536), .A2(n11368), .ZN(n13168) );
  INV_X1 U13768 ( .A(n13168), .ZN(n11082) );
  NOR2_X1 U13769 ( .A1(n11083), .A2(n11082), .ZN(n13318) );
  INV_X1 U13770 ( .A(n11084), .ZN(n11106) );
  NOR3_X1 U13771 ( .A1(n13318), .A2(n15731), .A3(n11106), .ZN(n11085) );
  AOI21_X1 U13772 ( .B1(n13877), .B2(n13535), .A(n11085), .ZN(n11371) );
  OAI22_X1 U13773 ( .A1(n13983), .A2(n11368), .B1(n15741), .B2(n10858), .ZN(
        n11086) );
  INV_X1 U13774 ( .A(n11086), .ZN(n11087) );
  OAI21_X1 U13775 ( .B1(n11371), .B2(n15739), .A(n11087), .ZN(P3_U3459) );
  INV_X1 U13776 ( .A(n11088), .ZN(n15518) );
  OAI211_X1 U13777 ( .C1(n11091), .C2(n11090), .A(n11089), .B(n14103), .ZN(
        n11098) );
  OAI22_X1 U13778 ( .A1(n11093), .A2(n14325), .B1(n11092), .B2(n14323), .ZN(
        n11267) );
  INV_X1 U13779 ( .A(n11267), .ZN(n11095) );
  OAI22_X1 U13780 ( .A1(n11095), .A2(n14096), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11094), .ZN(n11096) );
  AOI21_X1 U13781 ( .B1(n11272), .B2(n14107), .A(n11096), .ZN(n11097) );
  OAI211_X1 U13782 ( .C1(n15518), .C2(n14102), .A(n11098), .B(n11097), .ZN(
        P2_U3185) );
  OAI222_X1 U13783 ( .A1(n12850), .A2(n11100), .B1(n13382), .B2(n11099), .C1(
        P3_U3151), .C2(n11160), .ZN(P3_U3274) );
  NAND2_X1 U13784 ( .A1(n11120), .A2(n11109), .ZN(n11104) );
  OR2_X1 U13785 ( .A1(n11115), .A2(n11110), .ZN(n11102) );
  NAND4_X1 U13786 ( .A1(n11104), .A2(n11103), .A3(n11102), .A4(n11101), .ZN(
        n11105) );
  NAND2_X1 U13787 ( .A1(n11105), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11108) );
  NAND2_X1 U13788 ( .A1(n11118), .A2(n11106), .ZN(n13355) );
  OR2_X1 U13789 ( .A1(n11115), .A2(n13355), .ZN(n11107) );
  AND2_X1 U13790 ( .A1(n11278), .A2(n14035), .ZN(n11188) );
  INV_X1 U13791 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n11367) );
  INV_X1 U13792 ( .A(n13318), .ZN(n11123) );
  NAND2_X1 U13793 ( .A1(n11109), .A2(n15719), .ZN(n11113) );
  INV_X1 U13794 ( .A(n11110), .ZN(n11111) );
  NAND2_X1 U13795 ( .A1(n11115), .A2(n11111), .ZN(n11112) );
  OAI21_X1 U13796 ( .B1(n11120), .B2(n11113), .A(n11112), .ZN(n11114) );
  AND2_X1 U13797 ( .A1(n11118), .A2(n13347), .ZN(n11116) );
  NAND2_X1 U13798 ( .A1(n11116), .A2(n11115), .ZN(n11172) );
  NOR2_X1 U13799 ( .A1(n15719), .A2(n15698), .ZN(n11117) );
  NAND2_X1 U13800 ( .A1(n11118), .A2(n15731), .ZN(n11119) );
  OR2_X1 U13801 ( .A1(n11120), .A2(n11119), .ZN(n11121) );
  INV_X1 U13802 ( .A(n13520), .ZN(n13501) );
  OAI22_X1 U13803 ( .A1(n15691), .A2(n13514), .B1(n13501), .B2(n11368), .ZN(
        n11122) );
  AOI21_X1 U13804 ( .B1(n11123), .B2(n13492), .A(n11122), .ZN(n11124) );
  OAI21_X1 U13805 ( .B1(n11188), .B2(n11367), .A(n11124), .ZN(P3_U3172) );
  AOI22_X1 U13806 ( .A1(n6677), .A2(P2_REG2_REG_5__SCAN_IN), .B1(n11125), .B2(
        n15499), .ZN(n11126) );
  OAI21_X1 U13807 ( .B1(n15503), .B2(n11127), .A(n11126), .ZN(n11130) );
  NOR2_X1 U13808 ( .A1(n11128), .A2(n14362), .ZN(n11129) );
  AOI211_X1 U13809 ( .C1(n11131), .C2(n15498), .A(n11130), .B(n11129), .ZN(
        n11132) );
  OAI21_X1 U13810 ( .B1(n6677), .B2(n11133), .A(n11132), .ZN(P2_U3260) );
  INV_X1 U13811 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n11136) );
  NAND2_X1 U13812 ( .A1(n11134), .A2(n15543), .ZN(n11135) );
  OAI21_X1 U13813 ( .B1(n15543), .B2(n11136), .A(n11135), .ZN(P2_U3445) );
  INV_X1 U13814 ( .A(n11137), .ZN(n11138) );
  NAND3_X1 U13815 ( .A1(n11140), .A2(n11139), .A3(n11138), .ZN(n14784) );
  INV_X1 U13816 ( .A(n11141), .ZN(n11143) );
  INV_X2 U13817 ( .A(n14913), .ZN(n14962) );
  INV_X1 U13818 ( .A(n11144), .ZN(n11154) );
  NOR2_X2 U13819 ( .A1(n14962), .A2(n11145), .ZN(n15279) );
  NAND2_X1 U13820 ( .A1(n11146), .A2(n15279), .ZN(n11153) );
  NOR2_X2 U13821 ( .A1(n14962), .A2(n15275), .ZN(n14944) );
  OAI22_X1 U13822 ( .A1(n14913), .A2(n7783), .B1(n11213), .B2(n14982), .ZN(
        n11150) );
  NOR2_X1 U13823 ( .A1(n15273), .A2(n8213), .ZN(n11147) );
  NOR2_X1 U13824 ( .A1(n14949), .A2(n11148), .ZN(n11149) );
  AOI211_X1 U13825 ( .C1(n11151), .C2(n14944), .A(n11150), .B(n11149), .ZN(
        n11152) );
  OAI211_X1 U13826 ( .C1(n14962), .C2(n11154), .A(n11153), .B(n11152), .ZN(
        P1_U3288) );
  INV_X1 U13827 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n11157) );
  NAND2_X1 U13828 ( .A1(n11155), .A2(n15543), .ZN(n11156) );
  OAI21_X1 U13829 ( .B1(n15543), .B2(n11157), .A(n11156), .ZN(P2_U3430) );
  AND2_X4 U13830 ( .A1(n11164), .A2(n11163), .ZN(n12970) );
  NOR3_X1 U13831 ( .A1(n15691), .A2(n11173), .A3(n11573), .ZN(n11165) );
  INV_X1 U13832 ( .A(n11673), .ZN(n11167) );
  OAI21_X1 U13833 ( .B1(n11167), .B2(n11573), .A(n11166), .ZN(n11168) );
  INV_X1 U13834 ( .A(n11169), .ZN(n13320) );
  INV_X1 U13835 ( .A(n13320), .ZN(n11679) );
  NAND3_X1 U13836 ( .A1(n11679), .A2(n11573), .A3(n13172), .ZN(n11170) );
  OAI211_X1 U13837 ( .C1(n6818), .C2(n11673), .A(n11180), .B(n11170), .ZN(
        n11171) );
  NAND2_X1 U13838 ( .A1(n11171), .A2(n13492), .ZN(n11176) );
  INV_X1 U13839 ( .A(n9273), .ZN(n11285) );
  OAI22_X1 U13840 ( .A1(n11285), .A2(n13514), .B1(n13501), .B2(n11173), .ZN(
        n11174) );
  AOI21_X1 U13841 ( .B1(n13516), .B2(n13536), .A(n11174), .ZN(n11175) );
  OAI211_X1 U13842 ( .C1(n11188), .C2(n11177), .A(n11176), .B(n11175), .ZN(
        P3_U3162) );
  XNOR2_X1 U13843 ( .A(n11178), .B(n13364), .ZN(n11279) );
  XNOR2_X1 U13844 ( .A(n11279), .B(n9273), .ZN(n11182) );
  NAND2_X1 U13845 ( .A1(n11180), .A2(n7154), .ZN(n11181) );
  OAI21_X1 U13846 ( .B1(n11182), .B2(n11181), .A(n11281), .ZN(n11183) );
  NAND2_X1 U13847 ( .A1(n11183), .A2(n13492), .ZN(n11186) );
  OAI22_X1 U13848 ( .A1(n8839), .A2(n13514), .B1(n13501), .B2(n15697), .ZN(
        n11184) );
  AOI21_X1 U13849 ( .B1(n13516), .B2(n13535), .A(n11184), .ZN(n11185) );
  OAI211_X1 U13850 ( .C1(n11188), .C2(n11187), .A(n11186), .B(n11185), .ZN(
        P3_U3177) );
  NAND2_X1 U13851 ( .A1(n12599), .A2(n13103), .ZN(n11195) );
  NAND2_X1 U13852 ( .A1(n14660), .A2(n13068), .ZN(n11194) );
  NAND2_X1 U13853 ( .A1(n11195), .A2(n11194), .ZN(n11200) );
  INV_X1 U13854 ( .A(n11200), .ZN(n11196) );
  OAI22_X1 U13855 ( .A1(n11261), .A2(n13111), .B1(n11197), .B2(n6681), .ZN(
        n11198) );
  XNOR2_X1 U13856 ( .A(n11198), .B(n13115), .ZN(n11338) );
  NAND2_X1 U13857 ( .A1(n12608), .A2(n13102), .ZN(n11202) );
  NAND2_X1 U13858 ( .A1(n14659), .A2(n13103), .ZN(n11201) );
  NAND2_X1 U13859 ( .A1(n11202), .A2(n11201), .ZN(n11203) );
  XNOR2_X1 U13860 ( .A(n11203), .B(n13115), .ZN(n11207) );
  NAND2_X1 U13861 ( .A1(n12608), .A2(n13103), .ZN(n11205) );
  NAND2_X1 U13862 ( .A1(n14659), .A2(n13068), .ZN(n11204) );
  NAND2_X1 U13863 ( .A1(n11205), .A2(n11204), .ZN(n11206) );
  NOR2_X1 U13864 ( .A1(n11207), .A2(n11206), .ZN(n11344) );
  INV_X1 U13865 ( .A(n11344), .ZN(n11208) );
  NAND2_X1 U13866 ( .A1(n11207), .A2(n11206), .ZN(n11343) );
  NAND2_X1 U13867 ( .A1(n11208), .A2(n11343), .ZN(n11209) );
  XNOR2_X1 U13868 ( .A(n11345), .B(n11209), .ZN(n11216) );
  NAND2_X1 U13869 ( .A1(n15183), .A2(n11210), .ZN(n11211) );
  OAI211_X1 U13870 ( .C1(n15222), .C2(n11213), .A(n11212), .B(n11211), .ZN(
        n11214) );
  AOI21_X1 U13871 ( .B1(n15218), .B2(n12608), .A(n11214), .ZN(n11215) );
  OAI21_X1 U13872 ( .B1(n11216), .B2(n15212), .A(n11215), .ZN(P1_U3227) );
  NOR3_X1 U13873 ( .A1(n13655), .A2(n15677), .A3(n15666), .ZN(n11227) );
  AND2_X1 U13874 ( .A1(n15677), .A2(n11218), .ZN(n11221) );
  OAI22_X1 U13875 ( .A1(n15591), .A2(n11219), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11367), .ZN(n11220) );
  AOI211_X1 U13876 ( .C1(n11222), .C2(n13655), .A(n11221), .B(n11220), .ZN(
        n11226) );
  OR2_X1 U13877 ( .A1(n15595), .A2(n11223), .ZN(n11224) );
  OAI211_X1 U13878 ( .C1(n11227), .C2(n7267), .A(n11226), .B(n11225), .ZN(
        P3_U3182) );
  INV_X1 U13879 ( .A(n11327), .ZN(n11231) );
  OAI22_X1 U13880 ( .A1(n11229), .A2(n14325), .B1(n11228), .B2(n14323), .ZN(
        n11322) );
  AOI22_X1 U13881 ( .A1(n11322), .A2(n14131), .B1(P2_REG3_REG_6__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11230) );
  OAI21_X1 U13882 ( .B1(n11231), .B2(n14140), .A(n11230), .ZN(n11237) );
  INV_X1 U13883 ( .A(n11232), .ZN(n11233) );
  AOI211_X1 U13884 ( .C1(n11235), .C2(n11234), .A(n14148), .B(n11233), .ZN(
        n11236) );
  AOI211_X1 U13885 ( .C1(n11685), .C2(n14146), .A(n11237), .B(n11236), .ZN(
        n11238) );
  INV_X1 U13886 ( .A(n11238), .ZN(P2_U3211) );
  INV_X1 U13887 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n11239) );
  OAI22_X1 U13888 ( .A1(n14033), .A2(n11368), .B1(n15734), .B2(n11239), .ZN(
        n11240) );
  INV_X1 U13889 ( .A(n11240), .ZN(n11241) );
  OAI21_X1 U13890 ( .B1(n11371), .B2(n15732), .A(n11241), .ZN(P3_U3390) );
  NAND2_X1 U13891 ( .A1(n11243), .A2(n11242), .ZN(n11245) );
  XOR2_X1 U13892 ( .A(n11245), .B(n11244), .Z(n11250) );
  AOI22_X1 U13893 ( .A1(n14109), .A2(n14163), .B1(n14108), .B2(n14161), .ZN(
        n11246) );
  NAND2_X1 U13894 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n15421) );
  OAI211_X1 U13895 ( .C1(n11247), .C2(n14140), .A(n11246), .B(n15421), .ZN(
        n11248) );
  AOI21_X1 U13896 ( .B1(n15523), .B2(n14146), .A(n11248), .ZN(n11249) );
  OAI21_X1 U13897 ( .B1(n11250), .B2(n14148), .A(n11249), .ZN(P2_U3193) );
  NOR2_X1 U13898 ( .A1(n14049), .A2(SI_22_), .ZN(n11251) );
  AOI21_X1 U13899 ( .B1(n11252), .B2(P3_STATE_REG_SCAN_IN), .A(n11251), .ZN(
        n11253) );
  OAI21_X1 U13900 ( .B1(n11254), .B2(n12850), .A(n11253), .ZN(n11255) );
  INV_X1 U13901 ( .A(n11255), .ZN(P3_U3273) );
  NAND2_X1 U13902 ( .A1(n14913), .A2(n6966), .ZN(n14969) );
  NAND2_X1 U13903 ( .A1(n11256), .A2(n14944), .ZN(n11260) );
  INV_X1 U13904 ( .A(n11336), .ZN(n11258) );
  MUX2_X1 U13905 ( .A(n11333), .B(P1_REG2_REG_4__SCAN_IN), .S(n14962), .Z(
        n11257) );
  AOI21_X1 U13906 ( .B1(n15277), .B2(n11258), .A(n11257), .ZN(n11259) );
  OAI211_X1 U13907 ( .C1(n11261), .C2(n14949), .A(n11260), .B(n11259), .ZN(
        n11262) );
  AOI21_X1 U13908 ( .B1(n11263), .B2(n15279), .A(n11262), .ZN(n11264) );
  OAI21_X1 U13909 ( .B1(n11265), .B2(n14969), .A(n11264), .ZN(P1_U3289) );
  XNOR2_X1 U13910 ( .A(n11266), .B(n11269), .ZN(n11268) );
  AOI21_X1 U13911 ( .B1(n11268), .B2(n14358), .A(n11267), .ZN(n15517) );
  XNOR2_X1 U13912 ( .A(n11270), .B(n11269), .ZN(n15521) );
  NAND2_X1 U13913 ( .A1(n15521), .A2(n15496), .ZN(n11277) );
  INV_X1 U13914 ( .A(n11271), .ZN(n11325) );
  OAI211_X1 U13915 ( .C1(n11325), .C2(n15518), .A(n14398), .B(n11380), .ZN(
        n15516) );
  INV_X1 U13916 ( .A(n15516), .ZN(n11275) );
  AOI22_X1 U13917 ( .A1(n6677), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n11272), .B2(
        n15499), .ZN(n11273) );
  OAI21_X1 U13918 ( .B1(n15518), .B2(n15503), .A(n11273), .ZN(n11274) );
  AOI21_X1 U13919 ( .B1(n11275), .B2(n15498), .A(n11274), .ZN(n11276) );
  OAI211_X1 U13920 ( .C1(n6677), .C2(n15517), .A(n11277), .B(n11276), .ZN(
        P2_U3258) );
  NAND2_X1 U13921 ( .A1(n11285), .A2(n11279), .ZN(n11280) );
  AND2_X1 U13922 ( .A1(n11281), .A2(n11280), .ZN(n11283) );
  XNOR2_X1 U13923 ( .A(n12970), .B(n11287), .ZN(n11570) );
  XNOR2_X1 U13924 ( .A(n11570), .B(n8839), .ZN(n11282) );
  OAI211_X1 U13925 ( .C1(n11283), .C2(n11282), .A(n13492), .B(n11572), .ZN(
        n11289) );
  NOR2_X1 U13926 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11284), .ZN(n15553) );
  OAI22_X1 U13927 ( .A1(n11285), .A2(n13495), .B1(n11696), .B2(n13514), .ZN(
        n11286) );
  AOI211_X1 U13928 ( .C1(n11287), .C2(n13520), .A(n15553), .B(n11286), .ZN(
        n11288) );
  OAI211_X1 U13929 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n13518), .A(n11289), .B(
        n11288), .ZN(P3_U3158) );
  XNOR2_X1 U13930 ( .A(n15433), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n15430) );
  INV_X1 U13931 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11291) );
  MUX2_X1 U13932 ( .A(n11291), .B(P2_REG2_REG_11__SCAN_IN), .S(n11536), .Z(
        n11292) );
  INV_X1 U13933 ( .A(n11292), .ZN(n11293) );
  OAI21_X1 U13934 ( .B1(n11294), .B2(n11293), .A(n11535), .ZN(n11308) );
  OR2_X1 U13935 ( .A1(n11295), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n11296) );
  NAND2_X1 U13936 ( .A1(n11297), .A2(n11296), .ZN(n15426) );
  INV_X1 U13937 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n11298) );
  MUX2_X1 U13938 ( .A(n11298), .B(P2_REG1_REG_10__SCAN_IN), .S(n15433), .Z(
        n15427) );
  OR2_X1 U13939 ( .A1(n15426), .A2(n15427), .ZN(n15424) );
  NAND2_X1 U13940 ( .A1(n15433), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n11299) );
  NAND2_X1 U13941 ( .A1(n15424), .A2(n11299), .ZN(n11302) );
  INV_X1 U13942 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n11300) );
  MUX2_X1 U13943 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n11300), .S(n11536), .Z(
        n11301) );
  NAND2_X1 U13944 ( .A1(n11302), .A2(n11301), .ZN(n11529) );
  OAI211_X1 U13945 ( .C1(n11302), .C2(n11301), .A(n11529), .B(n15484), .ZN(
        n11305) );
  NOR2_X1 U13946 ( .A1(n11303), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11750) );
  AOI21_X1 U13947 ( .B1(n15333), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n11750), 
        .ZN(n11304) );
  OAI211_X1 U13948 ( .C1(n15489), .C2(n11306), .A(n11305), .B(n11304), .ZN(
        n11307) );
  AOI21_X1 U13949 ( .B1(n11308), .B2(n15478), .A(n11307), .ZN(n11309) );
  INV_X1 U13950 ( .A(n11309), .ZN(P2_U3225) );
  MUX2_X1 U13951 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n11310), .S(n14913), .Z(
        n11311) );
  INV_X1 U13952 ( .A(n11311), .ZN(n11314) );
  AOI22_X1 U13953 ( .A1(n14992), .A2(n12593), .B1(n15277), .B2(n11312), .ZN(
        n11313) );
  OAI211_X1 U13954 ( .C1(n14988), .C2(n11315), .A(n11314), .B(n11313), .ZN(
        P1_U3290) );
  XNOR2_X1 U13955 ( .A(n11316), .B(n11317), .ZN(n11323) );
  NAND2_X1 U13956 ( .A1(n11318), .A2(n11317), .ZN(n11319) );
  NAND2_X1 U13957 ( .A1(n11320), .A2(n11319), .ZN(n11688) );
  NOR2_X1 U13958 ( .A1(n11688), .A2(n10234), .ZN(n11321) );
  AOI211_X1 U13959 ( .C1(n14358), .C2(n11323), .A(n11322), .B(n11321), .ZN(
        n11687) );
  INV_X1 U13960 ( .A(n11324), .ZN(n11326) );
  AOI211_X1 U13961 ( .C1(n11685), .C2(n11326), .A(n12878), .B(n11325), .ZN(
        n11684) );
  AOI22_X1 U13962 ( .A1(n6677), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n11327), .B2(
        n15499), .ZN(n11328) );
  OAI21_X1 U13963 ( .B1(n11329), .B2(n15503), .A(n11328), .ZN(n11331) );
  NOR2_X1 U13964 ( .A1(n11688), .A2(n14381), .ZN(n11330) );
  AOI211_X1 U13965 ( .C1(n11684), .C2(n15498), .A(n11331), .B(n11330), .ZN(
        n11332) );
  OAI21_X1 U13966 ( .B1(n11687), .B2(n6677), .A(n11332), .ZN(P2_U3259) );
  NAND2_X1 U13967 ( .A1(n15183), .A2(n11333), .ZN(n11334) );
  OAI211_X1 U13968 ( .C1(n15222), .C2(n11336), .A(n11335), .B(n11334), .ZN(
        n11341) );
  XNOR2_X1 U13969 ( .A(n11337), .B(n11338), .ZN(n11339) );
  NOR2_X1 U13970 ( .A1(n11339), .A2(n15212), .ZN(n11340) );
  AOI211_X1 U13971 ( .C1(n15218), .C2(n12599), .A(n11341), .B(n11340), .ZN(
        n11342) );
  INV_X1 U13972 ( .A(n11342), .ZN(P1_U3230) );
  INV_X1 U13973 ( .A(n14627), .ZN(n14584) );
  NAND2_X1 U13974 ( .A1(n12611), .A2(n15224), .ZN(n15306) );
  OAI22_X1 U13975 ( .A1(n11548), .A2(n13111), .B1(n11346), .B2(n6681), .ZN(
        n11347) );
  XNOR2_X1 U13976 ( .A(n11347), .B(n13115), .ZN(n11635) );
  AND2_X1 U13977 ( .A1(n13068), .A2(n14658), .ZN(n11348) );
  AOI21_X1 U13978 ( .B1(n12611), .B2(n13103), .A(n11348), .ZN(n11636) );
  XNOR2_X1 U13979 ( .A(n11635), .B(n11636), .ZN(n11349) );
  OAI211_X1 U13980 ( .C1(n11350), .C2(n11349), .A(n11638), .B(n15179), .ZN(
        n11357) );
  INV_X1 U13981 ( .A(n11351), .ZN(n11550) );
  INV_X1 U13982 ( .A(n15183), .ZN(n14633) );
  NAND2_X1 U13983 ( .A1(n14659), .A2(n14974), .ZN(n11353) );
  NAND2_X1 U13984 ( .A1(n14657), .A2(n14975), .ZN(n11352) );
  AND2_X1 U13985 ( .A1(n11353), .A2(n11352), .ZN(n15307) );
  INV_X1 U13986 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n11354) );
  OAI22_X1 U13987 ( .A1(n14633), .A2(n15307), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11354), .ZN(n11355) );
  AOI21_X1 U13988 ( .B1(n11550), .B2(n14636), .A(n11355), .ZN(n11356) );
  OAI211_X1 U13989 ( .C1(n14584), .C2(n15306), .A(n11357), .B(n11356), .ZN(
        P1_U3239) );
  NAND2_X1 U13990 ( .A1(n11359), .A2(n11358), .ZN(n11362) );
  NAND2_X1 U13991 ( .A1(n14034), .A2(n11360), .ZN(n11361) );
  NAND2_X1 U13992 ( .A1(n11364), .A2(n11363), .ZN(n11366) );
  INV_X1 U13993 ( .A(n15703), .ZN(n13869) );
  OR2_X1 U13994 ( .A1(n15719), .A2(n11501), .ZN(n11365) );
  OAI22_X1 U13995 ( .A1(n13913), .A2(n11368), .B1(n13914), .B2(n11367), .ZN(
        n11369) );
  AOI21_X1 U13996 ( .B1(n13869), .B2(P3_REG2_REG_0__SCAN_IN), .A(n11369), .ZN(
        n11370) );
  OAI21_X1 U13997 ( .B1(n11371), .B2(n13921), .A(n11370), .ZN(P3_U3233) );
  XNOR2_X1 U13998 ( .A(n11372), .B(n11375), .ZN(n15528) );
  INV_X1 U13999 ( .A(n10234), .ZN(n14366) );
  OAI21_X1 U14000 ( .B1(n11375), .B2(n11374), .A(n11373), .ZN(n11376) );
  NAND2_X1 U14001 ( .A1(n11376), .A2(n14358), .ZN(n11378) );
  AOI22_X1 U14002 ( .A1(n14368), .A2(n14163), .B1(n14161), .B2(n14369), .ZN(
        n11377) );
  NAND2_X1 U14003 ( .A1(n11378), .A2(n11377), .ZN(n11379) );
  AOI21_X1 U14004 ( .B1(n15528), .B2(n14366), .A(n11379), .ZN(n15530) );
  NAND2_X1 U14005 ( .A1(n11380), .A2(n15523), .ZN(n11381) );
  NAND2_X1 U14006 ( .A1(n11381), .A2(n14398), .ZN(n11382) );
  OR2_X1 U14007 ( .A1(n11739), .A2(n11382), .ZN(n15524) );
  AOI22_X1 U14008 ( .A1(n6677), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n11383), .B2(
        n15499), .ZN(n11385) );
  INV_X1 U14009 ( .A(n15503), .ZN(n14389) );
  NAND2_X1 U14010 ( .A1(n15523), .A2(n14389), .ZN(n11384) );
  OAI211_X1 U14011 ( .C1(n15524), .C2(n14214), .A(n11385), .B(n11384), .ZN(
        n11386) );
  AOI21_X1 U14012 ( .B1(n15528), .B2(n14295), .A(n11386), .ZN(n11387) );
  OAI21_X1 U14013 ( .B1(n15530), .B2(n6677), .A(n11387), .ZN(P2_U3257) );
  INV_X1 U14014 ( .A(n11388), .ZN(n11390) );
  INV_X1 U14015 ( .A(n14751), .ZN(n14740) );
  OAI222_X1 U14016 ( .A1(n12476), .A2(n11389), .B1(n13377), .B2(n11390), .C1(
        P1_U3086), .C2(n14740), .ZN(P1_U3337) );
  OAI222_X1 U14017 ( .A1(n12959), .A2(n11391), .B1(n12957), .B2(n11390), .C1(
        P2_U3088), .C2(n15488), .ZN(P2_U3309) );
  OAI21_X1 U14018 ( .B1(n11393), .B2(n9280), .A(n11392), .ZN(n11822) );
  AND2_X1 U14019 ( .A1(n11395), .A2(n11394), .ZN(n11398) );
  OAI211_X1 U14020 ( .C1(n11398), .C2(n11397), .A(n11396), .B(n13874), .ZN(
        n11400) );
  AOI22_X1 U14021 ( .A1(n13880), .A2(n6679), .B1(n11949), .B2(n13877), .ZN(
        n11399) );
  NAND2_X1 U14022 ( .A1(n11400), .A2(n11399), .ZN(n11819) );
  AOI21_X1 U14023 ( .B1(n15724), .B2(n11822), .A(n11819), .ZN(n11405) );
  OAI22_X1 U14024 ( .A1(n14033), .A2(n11818), .B1(n15734), .B2(n8842), .ZN(
        n11401) );
  INV_X1 U14025 ( .A(n11401), .ZN(n11402) );
  OAI21_X1 U14026 ( .B1(n11405), .B2(n15732), .A(n11402), .ZN(P3_U3402) );
  OAI22_X1 U14027 ( .A1(n13983), .A2(n11818), .B1(n15741), .B2(n11856), .ZN(
        n11403) );
  INV_X1 U14028 ( .A(n11403), .ZN(n11404) );
  OAI21_X1 U14029 ( .B1(n11405), .B2(n15739), .A(n11404), .ZN(P3_U3463) );
  NAND2_X1 U14030 ( .A1(n11406), .A2(n14037), .ZN(n11407) );
  OAI211_X1 U14031 ( .C1(n11408), .C2(n13382), .A(n11407), .B(n13359), .ZN(
        P3_U3272) );
  INV_X1 U14032 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n11409) );
  NAND2_X1 U14033 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n12455)
         );
  OAI21_X1 U14034 ( .B1(n15271), .B2(n11409), .A(n12455), .ZN(n11427) );
  NOR2_X1 U14035 ( .A1(n11712), .A2(n12144), .ZN(n11410) );
  AOI21_X1 U14036 ( .B1(n11712), .B2(n12144), .A(n11410), .ZN(n11417) );
  INV_X1 U14037 ( .A(n11411), .ZN(n11413) );
  NAND2_X1 U14038 ( .A1(n11413), .A2(n11412), .ZN(n11414) );
  OAI21_X1 U14039 ( .B1(n11415), .B2(n7869), .A(n11414), .ZN(n11416) );
  NOR2_X1 U14040 ( .A1(n11417), .A2(n11416), .ZN(n11718) );
  AOI21_X1 U14041 ( .B1(n11417), .B2(n11416), .A(n11718), .ZN(n11425) );
  NAND2_X1 U14042 ( .A1(n11712), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n11418) );
  OAI21_X1 U14043 ( .B1(n11712), .B2(P1_REG1_REG_12__SCAN_IN), .A(n11418), 
        .ZN(n11423) );
  INV_X1 U14044 ( .A(n11715), .ZN(n11421) );
  AOI21_X1 U14045 ( .B1(n11423), .B2(n11422), .A(n11421), .ZN(n11424) );
  OAI22_X1 U14046 ( .A1(n15266), .A2(n11425), .B1(n11424), .B2(n14759), .ZN(
        n11426) );
  AOI211_X1 U14047 ( .C1(n11712), .C2(n15263), .A(n11427), .B(n11426), .ZN(
        n11428) );
  INV_X1 U14048 ( .A(n11428), .ZN(P1_U3255) );
  INV_X1 U14049 ( .A(n11429), .ZN(n11430) );
  AOI21_X1 U14050 ( .B1(n12788), .B2(n11431), .A(n11430), .ZN(n11437) );
  OAI21_X1 U14051 ( .B1(n12788), .B2(n11433), .A(n11432), .ZN(n11434) );
  NAND2_X1 U14052 ( .A1(n11434), .A2(n14980), .ZN(n11436) );
  AOI22_X1 U14053 ( .A1(n14974), .A2(n14656), .B1(n14654), .B2(n14975), .ZN(
        n11435) );
  OAI211_X1 U14054 ( .C1(n15286), .C2(n11437), .A(n11436), .B(n11435), .ZN(
        n11512) );
  INV_X1 U14055 ( .A(n11512), .ZN(n11443) );
  XNOR2_X1 U14056 ( .A(n11606), .B(n12093), .ZN(n11438) );
  NOR2_X1 U14057 ( .A1(n11438), .A2(n14958), .ZN(n11511) );
  NOR2_X1 U14058 ( .A1(n12093), .A2(n14949), .ZN(n11441) );
  OAI22_X1 U14059 ( .A1(n14913), .A2(n11439), .B1(n12099), .B2(n14982), .ZN(
        n11440) );
  AOI211_X1 U14060 ( .C1(n11511), .C2(n14944), .A(n11441), .B(n11440), .ZN(
        n11442) );
  OAI21_X1 U14061 ( .B1(n11443), .B2(n14962), .A(n11442), .ZN(P1_U3284) );
  NAND2_X1 U14062 ( .A1(n13299), .A2(n6678), .ZN(n11444) );
  OAI21_X1 U14063 ( .B1(P3_U3897), .B2(n11445), .A(n11444), .ZN(P3_U3518) );
  INV_X1 U14064 ( .A(n11446), .ZN(n11447) );
  AOI21_X1 U14065 ( .B1(n11449), .B2(n11448), .A(n11447), .ZN(n11457) );
  INV_X1 U14066 ( .A(n11742), .ZN(n11454) );
  NAND2_X1 U14067 ( .A1(n14160), .A2(n14369), .ZN(n11451) );
  NAND2_X1 U14068 ( .A1(n14162), .A2(n14368), .ZN(n11450) );
  NAND2_X1 U14069 ( .A1(n11451), .A2(n11450), .ZN(n11736) );
  NAND2_X1 U14070 ( .A1(n14131), .A2(n11736), .ZN(n11453) );
  OAI211_X1 U14071 ( .C1(n14140), .C2(n11454), .A(n11453), .B(n11452), .ZN(
        n11455) );
  AOI21_X1 U14072 ( .B1(n11995), .B2(n14146), .A(n11455), .ZN(n11456) );
  OAI21_X1 U14073 ( .B1(n11457), .B2(n14148), .A(n11456), .ZN(P2_U3203) );
  INV_X1 U14074 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n11458) );
  OAI22_X1 U14075 ( .A1(n14517), .A2(n11459), .B1(n15543), .B2(n11458), .ZN(
        n11460) );
  INV_X1 U14076 ( .A(n11460), .ZN(n11461) );
  OAI21_X1 U14077 ( .B1(n11462), .B2(n15541), .A(n11461), .ZN(P2_U3442) );
  INV_X1 U14078 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n11463) );
  OAI22_X1 U14079 ( .A1(n14517), .A2(n11464), .B1(n15543), .B2(n11463), .ZN(
        n11465) );
  INV_X1 U14080 ( .A(n11465), .ZN(n11466) );
  OAI21_X1 U14081 ( .B1(n11467), .B2(n15541), .A(n11466), .ZN(P2_U3439) );
  INV_X1 U14082 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n11468) );
  OAI22_X1 U14083 ( .A1(n14517), .A2(n15502), .B1(n15543), .B2(n11468), .ZN(
        n11469) );
  INV_X1 U14084 ( .A(n11469), .ZN(n11470) );
  OAI21_X1 U14085 ( .B1(n11471), .B2(n15541), .A(n11470), .ZN(P2_U3433) );
  INV_X1 U14086 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n11472) );
  OAI22_X1 U14087 ( .A1(n14517), .A2(n8299), .B1(n15543), .B2(n11472), .ZN(
        n11473) );
  INV_X1 U14088 ( .A(n11473), .ZN(n11474) );
  OAI21_X1 U14089 ( .B1(n11475), .B2(n15541), .A(n11474), .ZN(P2_U3436) );
  INV_X1 U14090 ( .A(n11547), .ZN(n11477) );
  OAI211_X1 U14091 ( .C1(n11477), .C2(n11476), .A(n15049), .B(n11605), .ZN(
        n15313) );
  XNOR2_X1 U14092 ( .A(n11478), .B(n12784), .ZN(n11485) );
  OAI21_X1 U14093 ( .B1(n11479), .B2(n11481), .A(n11480), .ZN(n11482) );
  NAND2_X1 U14094 ( .A1(n11482), .A2(n14980), .ZN(n11484) );
  AOI22_X1 U14095 ( .A1(n14974), .A2(n14658), .B1(n14656), .B2(n14975), .ZN(
        n11483) );
  OAI211_X1 U14096 ( .C1(n15286), .C2(n11485), .A(n11484), .B(n11483), .ZN(
        n15314) );
  INV_X1 U14097 ( .A(n15314), .ZN(n11486) );
  MUX2_X1 U14098 ( .A(n11487), .B(n11486), .S(n14913), .Z(n11490) );
  INV_X1 U14099 ( .A(n11643), .ZN(n11488) );
  AOI22_X1 U14100 ( .A1(n14992), .A2(n12620), .B1(n11488), .B2(n15277), .ZN(
        n11489) );
  OAI211_X1 U14101 ( .C1(n14988), .C2(n15313), .A(n11490), .B(n11489), .ZN(
        P1_U3286) );
  INV_X1 U14102 ( .A(n13319), .ZN(n11496) );
  XNOR2_X1 U14103 ( .A(n11491), .B(n11496), .ZN(n11500) );
  AOI22_X1 U14104 ( .A1(n8859), .A2(n13877), .B1(n13880), .B2(n9273), .ZN(
        n11499) );
  AND2_X1 U14105 ( .A1(n11493), .A2(n11492), .ZN(n11494) );
  INV_X1 U14106 ( .A(n11494), .ZN(n11497) );
  OR2_X1 U14107 ( .A1(n11494), .A2(n13319), .ZN(n11495) );
  OAI211_X1 U14108 ( .C1(n11497), .C2(n11496), .A(n13874), .B(n11495), .ZN(
        n11498) );
  OAI211_X1 U14109 ( .C1(n11500), .C2(n13728), .A(n11499), .B(n11498), .ZN(
        n15714) );
  INV_X1 U14110 ( .A(n15714), .ZN(n11505) );
  INV_X1 U14111 ( .A(n11500), .ZN(n15717) );
  AND2_X1 U14112 ( .A1(n13173), .A2(n11501), .ZN(n15699) );
  NAND2_X1 U14113 ( .A1(n15703), .A2(n15699), .ZN(n11681) );
  INV_X1 U14114 ( .A(n11681), .ZN(n13733) );
  NOR2_X1 U14115 ( .A1(n15703), .A2(n11852), .ZN(n11503) );
  OAI22_X1 U14116 ( .A1(n13913), .A2(n15713), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(n13914), .ZN(n11502) );
  AOI211_X1 U14117 ( .C1(n15717), .C2(n13733), .A(n11503), .B(n11502), .ZN(
        n11504) );
  OAI21_X1 U14118 ( .B1(n11505), .B2(n13921), .A(n11504), .ZN(P3_U3230) );
  INV_X1 U14119 ( .A(P3_DATAO_REG_29__SCAN_IN), .ZN(n11508) );
  INV_X1 U14120 ( .A(n13702), .ZN(n11506) );
  NAND2_X1 U14121 ( .A1(n11506), .A2(n6678), .ZN(n11507) );
  OAI21_X1 U14122 ( .B1(P3_U3897), .B2(n11508), .A(n11507), .ZN(P3_U3520) );
  INV_X1 U14123 ( .A(n13153), .ZN(n13158) );
  NAND2_X1 U14124 ( .A1(n13158), .A2(n6678), .ZN(n11509) );
  OAI21_X1 U14125 ( .B1(n6678), .B2(n11510), .A(n11509), .ZN(P3_U3521) );
  NOR2_X1 U14126 ( .A1(n11512), .A2(n11511), .ZN(n11517) );
  AOI22_X1 U14127 ( .A1(n12632), .A2(n12189), .B1(n15330), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n11513) );
  OAI21_X1 U14128 ( .B1(n11517), .B2(n15330), .A(n11513), .ZN(P1_U3537) );
  INV_X1 U14129 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n11514) );
  OAI22_X1 U14130 ( .A1(n12093), .A2(n15089), .B1(n15324), .B2(n11514), .ZN(
        n11515) );
  INV_X1 U14131 ( .A(n11515), .ZN(n11516) );
  OAI21_X1 U14132 ( .B1(n11517), .B2(n10226), .A(n11516), .ZN(P1_U3486) );
  INV_X1 U14133 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n11522) );
  NAND2_X1 U14134 ( .A1(n9266), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n11520) );
  INV_X1 U14135 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n11518) );
  OR2_X1 U14136 ( .A1(n8860), .A2(n11518), .ZN(n11519) );
  OAI211_X1 U14137 ( .C1(n11522), .C2(n11521), .A(n11520), .B(n11519), .ZN(
        n11523) );
  INV_X1 U14138 ( .A(n11523), .ZN(n11524) );
  AND2_X1 U14139 ( .A1(n11525), .A2(n11524), .ZN(n13684) );
  INV_X1 U14140 ( .A(n13684), .ZN(n13157) );
  NAND2_X1 U14141 ( .A1(n13157), .A2(n6678), .ZN(n11526) );
  OAI21_X1 U14142 ( .B1(P3_U3897), .B2(n11527), .A(n11526), .ZN(P3_U3522) );
  INV_X1 U14143 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n15165) );
  MUX2_X1 U14144 ( .A(n15165), .B(P2_REG1_REG_12__SCAN_IN), .S(n11975), .Z(
        n11532) );
  NAND2_X1 U14145 ( .A1(n11536), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n11528) );
  NAND2_X1 U14146 ( .A1(n11529), .A2(n11528), .ZN(n11531) );
  INV_X1 U14147 ( .A(n11977), .ZN(n11530) );
  AOI21_X1 U14148 ( .B1(n11532), .B2(n11531), .A(n11530), .ZN(n11544) );
  INV_X1 U14149 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11533) );
  MUX2_X1 U14150 ( .A(n11533), .B(P2_REG2_REG_12__SCAN_IN), .S(n11975), .Z(
        n11534) );
  INV_X1 U14151 ( .A(n11534), .ZN(n11538) );
  OAI21_X1 U14152 ( .B1(n11538), .B2(n11537), .A(n11971), .ZN(n11539) );
  NAND2_X1 U14153 ( .A1(n11539), .A2(n15478), .ZN(n11543) );
  NAND2_X1 U14154 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n12017)
         );
  OAI21_X1 U14155 ( .B1(n15489), .B2(n11540), .A(n12017), .ZN(n11541) );
  AOI21_X1 U14156 ( .B1(n15333), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n11541), 
        .ZN(n11542) );
  OAI211_X1 U14157 ( .C1(n11544), .C2(n15465), .A(n11543), .B(n11542), .ZN(
        P2_U3226) );
  OAI21_X1 U14158 ( .B1(n11546), .B2(n11552), .A(n11545), .ZN(n15311) );
  OAI211_X1 U14159 ( .C1(n11549), .C2(n11548), .A(n15049), .B(n11547), .ZN(
        n15308) );
  AOI22_X1 U14160 ( .A1(n14992), .A2(n12611), .B1(n11550), .B2(n15277), .ZN(
        n11551) );
  OAI21_X1 U14161 ( .B1(n15308), .B2(n14988), .A(n11551), .ZN(n11558) );
  XNOR2_X1 U14162 ( .A(n11553), .B(n11552), .ZN(n11554) );
  NOR2_X1 U14163 ( .A1(n11554), .A2(n15286), .ZN(n15310) );
  INV_X1 U14164 ( .A(n15310), .ZN(n11555) );
  NAND2_X1 U14165 ( .A1(n11555), .A2(n15307), .ZN(n11556) );
  MUX2_X1 U14166 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n11556), .S(n14913), .Z(
        n11557) );
  AOI211_X1 U14167 ( .C1(n15279), .C2(n15311), .A(n11558), .B(n11557), .ZN(
        n11559) );
  INV_X1 U14168 ( .A(n11559), .ZN(P1_U3287) );
  NOR2_X1 U14169 ( .A1(n7742), .A2(n14871), .ZN(n15292) );
  OAI21_X1 U14170 ( .B1(n12775), .B2(n10603), .A(n6966), .ZN(n11562) );
  AOI21_X1 U14171 ( .B1(n12578), .B2(n10590), .A(n11590), .ZN(n11565) );
  XNOR2_X1 U14172 ( .A(n11565), .B(n6865), .ZN(n11560) );
  AOI21_X1 U14173 ( .B1(n11560), .B2(n6966), .A(n14664), .ZN(n11561) );
  AOI21_X1 U14174 ( .B1(n14869), .B2(n11562), .A(n11561), .ZN(n15296) );
  AOI211_X1 U14175 ( .C1(n15277), .C2(P1_REG3_REG_1__SCAN_IN), .A(n15292), .B(
        n15296), .ZN(n11569) );
  OAI21_X1 U14176 ( .B1(n12775), .B2(n11564), .A(n11563), .ZN(n15298) );
  OAI22_X1 U14177 ( .A1(n14949), .A2(n15295), .B1(n14673), .B2(n14913), .ZN(
        n11567) );
  NAND2_X1 U14178 ( .A1(n11565), .A2(n15049), .ZN(n15294) );
  NOR2_X1 U14179 ( .A1(n14988), .A2(n15294), .ZN(n11566) );
  AOI211_X1 U14180 ( .C1(n15279), .C2(n15298), .A(n11567), .B(n11566), .ZN(
        n11568) );
  OAI21_X1 U14181 ( .B1(n11569), .B2(n14962), .A(n11568), .ZN(P1_U3292) );
  XNOR2_X1 U14182 ( .A(n11573), .B(n11578), .ZN(n11574) );
  NAND2_X1 U14183 ( .A1(n11574), .A2(n11696), .ZN(n11654) );
  OAI21_X1 U14184 ( .B1(n11574), .B2(n11696), .A(n11654), .ZN(n11651) );
  OR2_X1 U14185 ( .A1(n11653), .A2(n11651), .ZN(n11650) );
  INV_X1 U14186 ( .A(n11650), .ZN(n11575) );
  AOI21_X1 U14187 ( .B1(n11653), .B2(n11651), .A(n11575), .ZN(n11582) );
  NOR2_X1 U14188 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11576), .ZN(n15569) );
  OAI22_X1 U14189 ( .A1(n8839), .A2(n13495), .B1(n12007), .B2(n13514), .ZN(
        n11577) );
  AOI211_X1 U14190 ( .C1(n11578), .C2(n13520), .A(n15569), .B(n11577), .ZN(
        n11581) );
  INV_X1 U14191 ( .A(n13518), .ZN(n13498) );
  INV_X1 U14192 ( .A(n11817), .ZN(n11579) );
  NAND2_X1 U14193 ( .A1(n13498), .A2(n11579), .ZN(n11580) );
  OAI211_X1 U14194 ( .C1(n11582), .C2(n13523), .A(n11581), .B(n11580), .ZN(
        P3_U3170) );
  XNOR2_X1 U14195 ( .A(n12587), .B(n11583), .ZN(n11586) );
  INV_X1 U14196 ( .A(n11584), .ZN(n11585) );
  OAI21_X1 U14197 ( .B1(n11586), .B2(n15286), .A(n11585), .ZN(n15302) );
  INV_X1 U14198 ( .A(n15302), .ZN(n11595) );
  OAI21_X1 U14199 ( .B1(n11588), .B2(n12587), .A(n11587), .ZN(n15304) );
  OAI211_X1 U14200 ( .C1(n11590), .C2(n15301), .A(n11589), .B(n15049), .ZN(
        n15300) );
  OAI22_X1 U14201 ( .A1(n14913), .A2(n7730), .B1(n14679), .B2(n14982), .ZN(
        n11591) );
  AOI21_X1 U14202 ( .B1(n14992), .B2(n12589), .A(n11591), .ZN(n11592) );
  OAI21_X1 U14203 ( .B1(n14988), .B2(n15300), .A(n11592), .ZN(n11593) );
  AOI21_X1 U14204 ( .B1(n15279), .B2(n15304), .A(n11593), .ZN(n11594) );
  OAI21_X1 U14205 ( .B1(n14962), .B2(n11595), .A(n11594), .ZN(P1_U3291) );
  INV_X1 U14206 ( .A(n11596), .ZN(n12956) );
  OAI222_X1 U14207 ( .A1(n12476), .A2(n11597), .B1(n13377), .B2(n12956), .C1(
        P1_U3086), .C2(n14764), .ZN(P1_U3336) );
  XNOR2_X1 U14208 ( .A(n11598), .B(n11599), .ZN(n15322) );
  INV_X1 U14209 ( .A(n15322), .ZN(n11614) );
  INV_X1 U14210 ( .A(n15279), .ZN(n14862) );
  NAND2_X1 U14211 ( .A1(n11600), .A2(n11599), .ZN(n11601) );
  NAND3_X1 U14212 ( .A1(n11602), .A2(n6966), .A3(n11601), .ZN(n11604) );
  AOI22_X1 U14213 ( .A1(n14974), .A2(n14657), .B1(n14655), .B2(n14975), .ZN(
        n11603) );
  NAND2_X1 U14214 ( .A1(n11604), .A2(n11603), .ZN(n15320) );
  INV_X1 U14215 ( .A(n12623), .ZN(n15318) );
  INV_X1 U14216 ( .A(n11605), .ZN(n11608) );
  INV_X1 U14217 ( .A(n11606), .ZN(n11607) );
  OAI211_X1 U14218 ( .C1(n15318), .C2(n11608), .A(n11607), .B(n15049), .ZN(
        n15316) );
  OAI22_X1 U14219 ( .A1(n14913), .A2(n11609), .B1(n11932), .B2(n14982), .ZN(
        n11610) );
  AOI21_X1 U14220 ( .B1(n12623), .B2(n14992), .A(n11610), .ZN(n11611) );
  OAI21_X1 U14221 ( .B1(n15316), .B2(n14988), .A(n11611), .ZN(n11612) );
  AOI21_X1 U14222 ( .B1(n15320), .B2(n14913), .A(n11612), .ZN(n11613) );
  OAI21_X1 U14223 ( .B1(n11614), .B2(n14862), .A(n11613), .ZN(P1_U3285) );
  XNOR2_X1 U14224 ( .A(n11616), .B(n11615), .ZN(n11621) );
  INV_X1 U14225 ( .A(n11785), .ZN(n11618) );
  AOI22_X1 U14226 ( .A1(n14109), .A2(n14161), .B1(n14108), .B2(n14159), .ZN(
        n11617) );
  NAND2_X1 U14227 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n15434)
         );
  OAI211_X1 U14228 ( .C1(n11618), .C2(n14140), .A(n11617), .B(n15434), .ZN(
        n11619) );
  AOI21_X1 U14229 ( .B1(n15533), .B2(n14146), .A(n11619), .ZN(n11620) );
  OAI21_X1 U14230 ( .B1(n11621), .B2(n14148), .A(n11620), .ZN(P2_U3189) );
  OAI21_X1 U14231 ( .B1(n11623), .B2(n12789), .A(n11622), .ZN(n11670) );
  OAI211_X1 U14232 ( .C1(n6814), .C2(n11625), .A(n6966), .B(n11624), .ZN(
        n11663) );
  AOI21_X1 U14233 ( .B1(n11626), .B2(n12641), .A(n14958), .ZN(n11629) );
  NAND2_X1 U14234 ( .A1(n14655), .A2(n14974), .ZN(n11628) );
  NAND2_X1 U14235 ( .A1(n14653), .A2(n14975), .ZN(n11627) );
  NAND2_X1 U14236 ( .A1(n11628), .A2(n11627), .ZN(n15182) );
  AOI21_X1 U14237 ( .B1(n11629), .B2(n11804), .A(n15182), .ZN(n11667) );
  NAND2_X1 U14238 ( .A1(n11663), .A2(n11667), .ZN(n11630) );
  AOI21_X1 U14239 ( .B1(n11670), .B2(n15321), .A(n11630), .ZN(n11634) );
  AOI22_X1 U14240 ( .A1(n12641), .A2(n12189), .B1(n15330), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n11631) );
  OAI21_X1 U14241 ( .B1(n11634), .B2(n15330), .A(n11631), .ZN(P1_U3538) );
  INV_X1 U14242 ( .A(n12641), .ZN(n15187) );
  OAI22_X1 U14243 ( .A1(n15187), .A2(n15089), .B1(n15324), .B2(n7850), .ZN(
        n11632) );
  INV_X1 U14244 ( .A(n11632), .ZN(n11633) );
  OAI21_X1 U14245 ( .B1(n11634), .B2(n10226), .A(n11633), .ZN(P1_U3489) );
  NAND2_X1 U14246 ( .A1(n12620), .A2(n15224), .ZN(n15312) );
  INV_X1 U14247 ( .A(n11635), .ZN(n11637) );
  AND2_X1 U14248 ( .A1(n13068), .A2(n14657), .ZN(n11639) );
  AOI21_X1 U14249 ( .B1(n12620), .B2(n13103), .A(n11639), .ZN(n11923) );
  AOI22_X1 U14250 ( .A1(n12620), .A2(n13102), .B1(n13103), .B2(n14657), .ZN(
        n11640) );
  XNOR2_X1 U14251 ( .A(n11640), .B(n13115), .ZN(n11922) );
  XOR2_X1 U14252 ( .A(n11923), .B(n11922), .Z(n11641) );
  OAI211_X1 U14253 ( .C1(n11642), .C2(n11641), .A(n11926), .B(n15179), .ZN(
        n11649) );
  NOR2_X1 U14254 ( .A1(n15222), .A2(n11643), .ZN(n11647) );
  OAI21_X1 U14255 ( .B1(n15205), .B2(n11645), .A(n11644), .ZN(n11646) );
  AOI211_X1 U14256 ( .C1(n14587), .C2(n14658), .A(n11647), .B(n11646), .ZN(
        n11648) );
  OAI211_X1 U14257 ( .C1(n14584), .C2(n15312), .A(n11649), .B(n11648), .ZN(
        P1_U3213) );
  XNOR2_X1 U14258 ( .A(n11795), .B(n13364), .ZN(n11950) );
  XNOR2_X1 U14259 ( .A(n11950), .B(n12007), .ZN(n11657) );
  NAND2_X1 U14260 ( .A1(n11650), .A2(n11654), .ZN(n11656) );
  INV_X1 U14261 ( .A(n11657), .ZN(n11655) );
  OR2_X1 U14262 ( .A1(n11651), .A2(n11655), .ZN(n11652) );
  OAI21_X1 U14263 ( .B1(n11657), .B2(n11656), .A(n11952), .ZN(n11658) );
  NAND2_X1 U14264 ( .A1(n11658), .A2(n13492), .ZN(n11662) );
  NOR2_X1 U14265 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8862), .ZN(n15589) );
  OAI22_X1 U14266 ( .A1(n11696), .A2(n13495), .B1(n12028), .B2(n13514), .ZN(
        n11659) );
  AOI211_X1 U14267 ( .C1(n11660), .C2(n13520), .A(n15589), .B(n11659), .ZN(
        n11661) );
  OAI211_X1 U14268 ( .C1(n11699), .C2(n13518), .A(n11662), .B(n11661), .ZN(
        P3_U3167) );
  NOR2_X1 U14269 ( .A1(n11663), .A2(n14962), .ZN(n11669) );
  INV_X1 U14270 ( .A(n15190), .ZN(n11664) );
  AOI22_X1 U14271 ( .A1(n14962), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n11664), 
        .B2(n15277), .ZN(n11666) );
  NAND2_X1 U14272 ( .A1(n12641), .A2(n14992), .ZN(n11665) );
  OAI211_X1 U14273 ( .C1(n11667), .C2(n14988), .A(n11666), .B(n11665), .ZN(
        n11668) );
  AOI211_X1 U14274 ( .C1(n11670), .C2(n15279), .A(n11669), .B(n11668), .ZN(
        n11671) );
  INV_X1 U14275 ( .A(n11671), .ZN(P1_U3283) );
  AND2_X1 U14276 ( .A1(n11672), .A2(n15731), .ZN(n15706) );
  XNOR2_X1 U14277 ( .A(n11679), .B(n11673), .ZN(n11674) );
  NAND2_X1 U14278 ( .A1(n11674), .A2(n13874), .ZN(n11676) );
  AOI22_X1 U14279 ( .A1(n13877), .A2(n9273), .B1(n13536), .B2(n13880), .ZN(
        n11675) );
  NAND2_X1 U14280 ( .A1(n11676), .A2(n11675), .ZN(n15705) );
  AOI21_X1 U14281 ( .B1(n15706), .B2(n15698), .A(n15705), .ZN(n11677) );
  MUX2_X1 U14282 ( .A(n11678), .B(n11677), .S(n15703), .Z(n11683) );
  XNOR2_X1 U14283 ( .A(n13172), .B(n11679), .ZN(n15707) );
  NAND2_X1 U14284 ( .A1(n15703), .A2(n15693), .ZN(n11680) );
  AOI22_X1 U14285 ( .A1(n15707), .A2(n13919), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15702), .ZN(n11682) );
  NAND2_X1 U14286 ( .A1(n11683), .A2(n11682), .ZN(P3_U3232) );
  AOI21_X1 U14287 ( .B1(n15532), .B2(n11685), .A(n11684), .ZN(n11686) );
  OAI211_X1 U14288 ( .C1(n14434), .C2(n11688), .A(n11687), .B(n11686), .ZN(
        n11704) );
  NAND2_X1 U14289 ( .A1(n11704), .A2(n15550), .ZN(n11689) );
  OAI21_X1 U14290 ( .B1(n15550), .B2(n11690), .A(n11689), .ZN(P2_U3505) );
  INV_X1 U14291 ( .A(n11692), .ZN(n11693) );
  AOI21_X1 U14292 ( .B1(n13316), .B2(n11694), .A(n11693), .ZN(n11695) );
  OAI222_X1 U14293 ( .A1(n15689), .A2(n12028), .B1(n15690), .B2(n11696), .C1(
        n15696), .C2(n11695), .ZN(n11790) );
  INV_X1 U14294 ( .A(n11790), .ZN(n11703) );
  OAI21_X1 U14295 ( .B1(n11698), .B2(n13316), .A(n11697), .ZN(n11791) );
  NOR2_X1 U14296 ( .A1(n15703), .A2(n11862), .ZN(n11701) );
  OAI22_X1 U14297 ( .A1(n13913), .A2(n11795), .B1(n11699), .B2(n13914), .ZN(
        n11700) );
  AOI211_X1 U14298 ( .C1(n11791), .C2(n13919), .A(n11701), .B(n11700), .ZN(
        n11702) );
  OAI21_X1 U14299 ( .B1(n11703), .B2(n13921), .A(n11702), .ZN(P3_U3228) );
  INV_X1 U14300 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n11706) );
  NAND2_X1 U14301 ( .A1(n11704), .A2(n15543), .ZN(n11705) );
  OAI21_X1 U14302 ( .B1(n15543), .B2(n11706), .A(n11705), .ZN(P2_U3448) );
  INV_X1 U14303 ( .A(n11707), .ZN(n13124) );
  OAI222_X1 U14304 ( .A1(n12959), .A2(n11709), .B1(P2_U3088), .B2(n11708), 
        .C1(n14531), .C2(n13124), .ZN(P2_U3307) );
  NAND2_X1 U14305 ( .A1(n11756), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n11710) );
  OAI21_X1 U14306 ( .B1(n11756), .B2(P1_REG1_REG_13__SCAN_IN), .A(n11710), 
        .ZN(n11711) );
  INV_X1 U14307 ( .A(n11711), .ZN(n11717) );
  INV_X1 U14308 ( .A(n11712), .ZN(n11719) );
  NAND2_X1 U14309 ( .A1(n11719), .A2(n11713), .ZN(n11714) );
  NAND2_X1 U14310 ( .A1(n11715), .A2(n11714), .ZN(n11716) );
  AOI211_X1 U14311 ( .C1(n11717), .C2(n11716), .A(n11758), .B(n14759), .ZN(
        n11727) );
  NOR2_X1 U14312 ( .A1(n11721), .A2(n11722), .ZN(n11720) );
  AOI211_X1 U14313 ( .C1(n11721), .C2(n11722), .A(n11720), .B(n11723), .ZN(
        n11725) );
  NOR2_X1 U14314 ( .A1(n11756), .A2(n11722), .ZN(n11768) );
  INV_X1 U14315 ( .A(n11723), .ZN(n11724) );
  NOR3_X1 U14316 ( .A1(n15266), .A2(n11725), .A3(n11770), .ZN(n11726) );
  NOR2_X1 U14317 ( .A1(n11727), .A2(n11726), .ZN(n11730) );
  NAND2_X1 U14318 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n12542)
         );
  INV_X1 U14319 ( .A(n12542), .ZN(n11728) );
  AOI21_X1 U14320 ( .B1(n14737), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n11728), 
        .ZN(n11729) );
  OAI211_X1 U14321 ( .C1(n11756), .C2(n14757), .A(n11730), .B(n11729), .ZN(
        P1_U3256) );
  XNOR2_X1 U14322 ( .A(n11732), .B(n11731), .ZN(n11987) );
  OAI21_X1 U14323 ( .B1(n11735), .B2(n11734), .A(n11733), .ZN(n11737) );
  AOI21_X1 U14324 ( .B1(n11737), .B2(n14358), .A(n11736), .ZN(n11738) );
  OAI21_X1 U14325 ( .B1(n11987), .B2(n10234), .A(n11738), .ZN(n11988) );
  NAND2_X1 U14326 ( .A1(n11988), .A2(n14397), .ZN(n11746) );
  INV_X1 U14327 ( .A(n11739), .ZN(n11741) );
  INV_X1 U14328 ( .A(n11782), .ZN(n11740) );
  AOI211_X1 U14329 ( .C1(n11995), .C2(n11741), .A(n12878), .B(n11740), .ZN(
        n11989) );
  AOI22_X1 U14330 ( .A1(n6677), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n11742), .B2(
        n15499), .ZN(n11743) );
  OAI21_X1 U14331 ( .B1(n11992), .B2(n15503), .A(n11743), .ZN(n11744) );
  AOI21_X1 U14332 ( .B1(n11989), .B2(n15498), .A(n11744), .ZN(n11745) );
  OAI211_X1 U14333 ( .C1(n11987), .C2(n14381), .A(n11746), .B(n11745), .ZN(
        P2_U3256) );
  XNOR2_X1 U14334 ( .A(n11748), .B(n11747), .ZN(n11753) );
  OAI22_X1 U14335 ( .A1(n12108), .A2(n14143), .B1(n14142), .B2(n12107), .ZN(
        n11749) );
  AOI211_X1 U14336 ( .C1(n14107), .C2(n12114), .A(n11750), .B(n11749), .ZN(
        n11752) );
  NAND2_X1 U14337 ( .A1(n12257), .A2(n14146), .ZN(n11751) );
  OAI211_X1 U14338 ( .C1(n11753), .C2(n14148), .A(n11752), .B(n11751), .ZN(
        P2_U3208) );
  NAND2_X1 U14339 ( .A1(n14695), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n11754) );
  OAI21_X1 U14340 ( .B1(n14695), .B2(P1_REG1_REG_14__SCAN_IN), .A(n11754), 
        .ZN(n11760) );
  INV_X1 U14341 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11755) );
  NOR2_X1 U14342 ( .A1(n11756), .A2(n11755), .ZN(n11757) );
  AOI21_X1 U14343 ( .B1(n11760), .B2(n11759), .A(n14694), .ZN(n11773) );
  NAND2_X1 U14344 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n15176)
         );
  INV_X1 U14345 ( .A(n15176), .ZN(n11762) );
  NOR2_X1 U14346 ( .A1(n14757), .A2(n14705), .ZN(n11761) );
  AOI211_X1 U14347 ( .C1(n14737), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n11762), 
        .B(n11761), .ZN(n11772) );
  NAND2_X1 U14348 ( .A1(n14695), .A2(n11763), .ZN(n11765) );
  INV_X1 U14349 ( .A(n11768), .ZN(n11764) );
  OAI211_X1 U14350 ( .C1(n14695), .C2(n11763), .A(n11765), .B(n11764), .ZN(
        n11769) );
  NAND2_X1 U14351 ( .A1(n14695), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11767) );
  NAND2_X1 U14352 ( .A1(n14705), .A2(n11763), .ZN(n11766) );
  OAI211_X1 U14353 ( .C1(n11770), .C2(n11768), .A(n11767), .B(n11766), .ZN(
        n14704) );
  OAI211_X1 U14354 ( .C1(n11770), .C2(n11769), .A(n14762), .B(n14704), .ZN(
        n11771) );
  OAI211_X1 U14355 ( .C1(n11773), .C2(n14759), .A(n11772), .B(n11771), .ZN(
        P1_U3257) );
  XNOR2_X1 U14356 ( .A(n11774), .B(n11777), .ZN(n15538) );
  OAI21_X1 U14357 ( .B1(n11777), .B2(n11776), .A(n11775), .ZN(n11778) );
  NAND2_X1 U14358 ( .A1(n11778), .A2(n14358), .ZN(n11780) );
  AOI22_X1 U14359 ( .A1(n14368), .A2(n14161), .B1(n14159), .B2(n14369), .ZN(
        n11779) );
  NAND2_X1 U14360 ( .A1(n11780), .A2(n11779), .ZN(n11781) );
  AOI21_X1 U14361 ( .B1(n15538), .B2(n14366), .A(n11781), .ZN(n15540) );
  AOI21_X1 U14362 ( .B1(n11782), .B2(n15533), .A(n12878), .ZN(n11784) );
  NAND2_X1 U14363 ( .A1(n11784), .A2(n12113), .ZN(n15535) );
  AOI22_X1 U14364 ( .A1(n6677), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n11785), 
        .B2(n15499), .ZN(n11787) );
  NAND2_X1 U14365 ( .A1(n15533), .A2(n14389), .ZN(n11786) );
  OAI211_X1 U14366 ( .C1(n15535), .C2(n14214), .A(n11787), .B(n11786), .ZN(
        n11788) );
  AOI21_X1 U14367 ( .B1(n15538), .B2(n14295), .A(n11788), .ZN(n11789) );
  OAI21_X1 U14368 ( .B1(n15540), .B2(n6677), .A(n11789), .ZN(P2_U3255) );
  AOI21_X1 U14369 ( .B1(n15724), .B2(n11791), .A(n11790), .ZN(n11798) );
  INV_X1 U14370 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n11792) );
  OAI22_X1 U14371 ( .A1(n14033), .A2(n11795), .B1(n15734), .B2(n11792), .ZN(
        n11793) );
  INV_X1 U14372 ( .A(n11793), .ZN(n11794) );
  OAI21_X1 U14373 ( .B1(n11798), .B2(n15732), .A(n11794), .ZN(P3_U3405) );
  OAI22_X1 U14374 ( .A1(n13983), .A2(n11795), .B1(n15741), .B2(n15601), .ZN(
        n11796) );
  INV_X1 U14375 ( .A(n11796), .ZN(n11797) );
  OAI21_X1 U14376 ( .B1(n11798), .B2(n15739), .A(n11797), .ZN(P3_U3464) );
  XNOR2_X1 U14377 ( .A(n11800), .B(n11799), .ZN(n11801) );
  OAI222_X1 U14378 ( .A1(n14871), .A2(n15204), .B1(n14869), .B2(n15207), .C1(
        n11801), .C2(n15286), .ZN(n11961) );
  INV_X1 U14379 ( .A(n11961), .ZN(n11812) );
  OAI21_X1 U14380 ( .B1(n11803), .B2(n12790), .A(n11802), .ZN(n11963) );
  NAND2_X1 U14381 ( .A1(n11804), .A2(n15217), .ZN(n11805) );
  NAND2_X1 U14382 ( .A1(n11805), .A2(n15049), .ZN(n11806) );
  NOR2_X1 U14383 ( .A1(n12135), .A2(n11806), .ZN(n11962) );
  NAND2_X1 U14384 ( .A1(n11962), .A2(n14944), .ZN(n11809) );
  INV_X1 U14385 ( .A(n15221), .ZN(n11807) );
  AOI22_X1 U14386 ( .A1(n14962), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n11807), 
        .B2(n15277), .ZN(n11808) );
  OAI211_X1 U14387 ( .C1(n7139), .C2(n14949), .A(n11809), .B(n11808), .ZN(
        n11810) );
  AOI21_X1 U14388 ( .B1(n11963), .B2(n15279), .A(n11810), .ZN(n11811) );
  OAI21_X1 U14389 ( .B1(n14962), .B2(n11812), .A(n11811), .ZN(P1_U3282) );
  INV_X1 U14390 ( .A(n11813), .ZN(n11815) );
  OAI222_X1 U14391 ( .A1(n12959), .A2(n11814), .B1(n12957), .B2(n11815), .C1(
        n8697), .C2(P2_U3088), .ZN(P2_U3306) );
  OAI222_X1 U14392 ( .A1(n12476), .A2(n11816), .B1(n13377), .B2(n11815), .C1(
        P1_U3086), .C2(n12813), .ZN(P1_U3334) );
  OAI22_X1 U14393 ( .A1(n13913), .A2(n11818), .B1(n11817), .B2(n13914), .ZN(
        n11821) );
  MUX2_X1 U14394 ( .A(n11819), .B(P3_REG2_REG_4__SCAN_IN), .S(n13869), .Z(
        n11820) );
  AOI211_X1 U14395 ( .C1(n13919), .C2(n11822), .A(n11821), .B(n11820), .ZN(
        n11823) );
  INV_X1 U14396 ( .A(n11823), .ZN(P3_U3229) );
  OAI211_X1 U14397 ( .C1(n11825), .C2(n12023), .A(n11824), .B(n13874), .ZN(
        n11827) );
  AOI22_X1 U14398 ( .A1(n13534), .A2(n13880), .B1(n13877), .B2(n13533), .ZN(
        n11826) );
  NAND2_X1 U14399 ( .A1(n11827), .A2(n11826), .ZN(n11940) );
  INV_X1 U14400 ( .A(n11940), .ZN(n11833) );
  OAI21_X1 U14401 ( .B1(n11829), .B2(n13317), .A(n11828), .ZN(n11941) );
  NOR2_X1 U14402 ( .A1(n15703), .A2(n11874), .ZN(n11831) );
  OAI22_X1 U14403 ( .A1(n13913), .A2(n11945), .B1(n12033), .B2(n13914), .ZN(
        n11830) );
  AOI211_X1 U14404 ( .C1(n11941), .C2(n13919), .A(n11831), .B(n11830), .ZN(
        n11832) );
  OAI21_X1 U14405 ( .B1(n11833), .B2(n13921), .A(n11832), .ZN(P3_U3226) );
  XNOR2_X1 U14406 ( .A(n11836), .B(n15561), .ZN(n15552) );
  NOR2_X1 U14407 ( .A1(n15552), .A2(n11852), .ZN(n15551) );
  INV_X1 U14408 ( .A(n11836), .ZN(n11837) );
  INV_X1 U14409 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11857) );
  XNOR2_X1 U14410 ( .A(n15578), .B(n11857), .ZN(n15568) );
  INV_X1 U14411 ( .A(n11839), .ZN(n11840) );
  NOR2_X1 U14412 ( .A1(n15588), .A2(n11862), .ZN(n15587) );
  NAND2_X1 U14413 ( .A1(P3_REG2_REG_6__SCAN_IN), .A2(n15615), .ZN(n11841) );
  OAI21_X1 U14414 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n15615), .A(n11841), .ZN(
        n15608) );
  NAND2_X1 U14415 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n15649), .ZN(n11844) );
  OAI21_X1 U14416 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n15649), .A(n11844), .ZN(
        n15643) );
  NOR2_X1 U14417 ( .A1(n11910), .A2(n11845), .ZN(n11846) );
  INV_X1 U14418 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n15661) );
  NAND2_X1 U14419 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n12262), .ZN(n11847) );
  OAI21_X1 U14420 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n12262), .A(n11847), 
        .ZN(n11848) );
  AOI21_X1 U14421 ( .B1(n11849), .B2(n11848), .A(n12260), .ZN(n11920) );
  INV_X1 U14422 ( .A(n11850), .ZN(n15556) );
  INV_X1 U14423 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n11851) );
  MUX2_X1 U14425 ( .A(n11852), .B(n11851), .S(n13629), .Z(n11853) );
  NAND2_X1 U14426 ( .A1(n11853), .A2(n15561), .ZN(n15572) );
  INV_X1 U14427 ( .A(n11853), .ZN(n11854) );
  NAND2_X1 U14428 ( .A1(n11854), .A2(n11902), .ZN(n11855) );
  AND2_X1 U14429 ( .A1(n15572), .A2(n11855), .ZN(n15555) );
  OAI21_X1 U14430 ( .B1(n15557), .B2(n15556), .A(n15555), .ZN(n15573) );
  MUX2_X1 U14431 ( .A(n11857), .B(n11856), .S(n13667), .Z(n11858) );
  NAND2_X1 U14432 ( .A1(n11858), .A2(n15578), .ZN(n11861) );
  INV_X1 U14433 ( .A(n11858), .ZN(n11859) );
  NAND2_X1 U14434 ( .A1(n11859), .A2(n11903), .ZN(n11860) );
  NAND2_X1 U14435 ( .A1(n11861), .A2(n11860), .ZN(n15571) );
  INV_X1 U14436 ( .A(n11861), .ZN(n15593) );
  MUX2_X1 U14437 ( .A(n11862), .B(n15601), .S(n13667), .Z(n11863) );
  NAND2_X1 U14438 ( .A1(n11863), .A2(n15599), .ZN(n15611) );
  INV_X1 U14439 ( .A(n11863), .ZN(n11865) );
  NAND2_X1 U14440 ( .A1(n11865), .A2(n11864), .ZN(n11866) );
  AND2_X1 U14441 ( .A1(n15611), .A2(n11866), .ZN(n15592) );
  OAI21_X1 U14442 ( .B1(n15594), .B2(n15593), .A(n15592), .ZN(n15612) );
  MUX2_X1 U14443 ( .A(n11868), .B(n11867), .S(n13629), .Z(n11869) );
  NAND2_X1 U14444 ( .A1(n11869), .A2(n11897), .ZN(n11872) );
  INV_X1 U14445 ( .A(n11869), .ZN(n11870) );
  NAND2_X1 U14446 ( .A1(n11870), .A2(n15615), .ZN(n11871) );
  NAND2_X1 U14447 ( .A1(n11872), .A2(n11871), .ZN(n15610) );
  AOI21_X1 U14448 ( .B1(n15612), .B2(n15611), .A(n15610), .ZN(n15629) );
  INV_X1 U14449 ( .A(n11872), .ZN(n15628) );
  MUX2_X1 U14450 ( .A(n11874), .B(n11873), .S(n13629), .Z(n11876) );
  NAND2_X1 U14451 ( .A1(n11876), .A2(n11875), .ZN(n15645) );
  INV_X1 U14452 ( .A(n11876), .ZN(n11877) );
  NAND2_X1 U14453 ( .A1(n11877), .A2(n15633), .ZN(n11878) );
  AND2_X1 U14454 ( .A1(n15645), .A2(n11878), .ZN(n15627) );
  OAI21_X1 U14455 ( .B1(n15629), .B2(n15628), .A(n15627), .ZN(n15646) );
  MUX2_X1 U14456 ( .A(n12161), .B(n11879), .S(n13629), .Z(n11880) );
  NAND2_X1 U14457 ( .A1(n11880), .A2(n11896), .ZN(n11883) );
  INV_X1 U14458 ( .A(n11880), .ZN(n11881) );
  NAND2_X1 U14459 ( .A1(n11881), .A2(n15649), .ZN(n11882) );
  NAND2_X1 U14460 ( .A1(n11883), .A2(n11882), .ZN(n15644) );
  INV_X1 U14461 ( .A(n11883), .ZN(n15664) );
  MUX2_X1 U14462 ( .A(n15661), .B(n11884), .S(n13629), .Z(n11885) );
  NAND2_X1 U14463 ( .A1(n11885), .A2(n11910), .ZN(n11893) );
  INV_X1 U14464 ( .A(n11885), .ZN(n11886) );
  NAND2_X1 U14465 ( .A1(n11886), .A2(n15670), .ZN(n11887) );
  AND2_X1 U14466 ( .A1(n11893), .A2(n11887), .ZN(n15663) );
  OAI21_X1 U14467 ( .B1(n15665), .B2(n15664), .A(n15663), .ZN(n15662) );
  MUX2_X1 U14468 ( .A(n12395), .B(n11888), .S(n13629), .Z(n11889) );
  NAND2_X1 U14469 ( .A1(n11889), .A2(n11895), .ZN(n12268) );
  INV_X1 U14470 ( .A(n11889), .ZN(n11890) );
  NAND2_X1 U14471 ( .A1(n11890), .A2(n12262), .ZN(n11891) );
  NAND2_X1 U14472 ( .A1(n12268), .A2(n11891), .ZN(n11892) );
  AOI21_X1 U14473 ( .B1(n15662), .B2(n11893), .A(n11892), .ZN(n12270) );
  AND3_X1 U14474 ( .A1(n15662), .A2(n11893), .A3(n11892), .ZN(n11894) );
  OAI21_X1 U14475 ( .B1(n12270), .B2(n11894), .A(n15666), .ZN(n11919) );
  AOI22_X1 U14476 ( .A1(n11895), .A2(n11888), .B1(P3_REG1_REG_10__SCAN_IN), 
        .B2(n12262), .ZN(n11913) );
  NAND2_X1 U14477 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n15649), .ZN(n11908) );
  AOI22_X1 U14478 ( .A1(n11896), .A2(n11879), .B1(P3_REG1_REG_8__SCAN_IN), 
        .B2(n15649), .ZN(n15653) );
  NAND2_X1 U14479 ( .A1(P3_REG1_REG_6__SCAN_IN), .A2(n15615), .ZN(n11905) );
  AOI22_X1 U14480 ( .A1(n11897), .A2(n11867), .B1(P3_REG1_REG_6__SCAN_IN), 
        .B2(n15615), .ZN(n15619) );
  OAI21_X1 U14481 ( .B1(n11900), .B2(n11899), .A(n11898), .ZN(n11901) );
  MUX2_X1 U14482 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n11856), .S(n15578), .Z(
        n15580) );
  XNOR2_X1 U14483 ( .A(n11904), .B(n15599), .ZN(n15602) );
  OAI22_X1 U14484 ( .A1(n15602), .A2(n15601), .B1(n15599), .B2(n11904), .ZN(
        n15620) );
  NAND2_X1 U14485 ( .A1(n15633), .A2(n11906), .ZN(n11907) );
  NAND2_X1 U14486 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n15637), .ZN(n15636) );
  NAND2_X1 U14487 ( .A1(n11907), .A2(n15636), .ZN(n15654) );
  NAND2_X1 U14488 ( .A1(n15670), .A2(n11909), .ZN(n11911) );
  XNOR2_X1 U14489 ( .A(n11910), .B(n11909), .ZN(n15676) );
  NAND2_X1 U14490 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n15676), .ZN(n15675) );
  NAND2_X1 U14491 ( .A1(n11911), .A2(n15675), .ZN(n11912) );
  OAI21_X1 U14492 ( .B1(n11913), .B2(n11912), .A(n12263), .ZN(n11917) );
  NOR2_X1 U14493 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11914), .ZN(n12359) );
  AOI21_X1 U14494 ( .B1(n15674), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n12359), 
        .ZN(n11915) );
  OAI21_X1 U14495 ( .B1(n15671), .B2(n12262), .A(n11915), .ZN(n11916) );
  AOI21_X1 U14496 ( .B1(n11917), .B2(n15677), .A(n11916), .ZN(n11918) );
  OAI211_X1 U14497 ( .C1(n11920), .C2(n15681), .A(n11919), .B(n11918), .ZN(
        P3_U3192) );
  AOI22_X1 U14498 ( .A1(n12623), .A2(n13102), .B1(n13103), .B2(n14656), .ZN(
        n11921) );
  XNOR2_X1 U14499 ( .A(n11921), .B(n13115), .ZN(n12087) );
  AOI22_X1 U14500 ( .A1(n12623), .A2(n13103), .B1(n13068), .B2(n14656), .ZN(
        n12088) );
  XNOR2_X1 U14501 ( .A(n12087), .B(n12088), .ZN(n11928) );
  INV_X1 U14502 ( .A(n11922), .ZN(n11925) );
  INV_X1 U14503 ( .A(n11923), .ZN(n11924) );
  NOR2_X1 U14504 ( .A1(n11927), .A2(n11928), .ZN(n12086) );
  AOI21_X1 U14505 ( .B1(n11928), .B2(n11927), .A(n12086), .ZN(n11935) );
  AOI21_X1 U14506 ( .B1(n14615), .B2(n14655), .A(n11929), .ZN(n11931) );
  NAND2_X1 U14507 ( .A1(n14587), .A2(n14657), .ZN(n11930) );
  OAI211_X1 U14508 ( .C1(n15222), .C2(n11932), .A(n11931), .B(n11930), .ZN(
        n11933) );
  AOI21_X1 U14509 ( .B1(n12623), .B2(n15218), .A(n11933), .ZN(n11934) );
  OAI21_X1 U14510 ( .B1(n11935), .B2(n15212), .A(n11934), .ZN(P1_U3221) );
  INV_X1 U14511 ( .A(n11936), .ZN(n11938) );
  OAI222_X1 U14512 ( .A1(P3_U3151), .A2(n11939), .B1(n12850), .B2(n11938), 
        .C1(n11937), .C2(n13382), .ZN(P3_U3271) );
  AOI21_X1 U14513 ( .B1(n15724), .B2(n11941), .A(n11940), .ZN(n11948) );
  INV_X1 U14514 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n11942) );
  OAI22_X1 U14515 ( .A1(n14033), .A2(n11945), .B1(n15734), .B2(n11942), .ZN(
        n11943) );
  INV_X1 U14516 ( .A(n11943), .ZN(n11944) );
  OAI21_X1 U14517 ( .B1(n11948), .B2(n15732), .A(n11944), .ZN(P3_U3411) );
  OAI22_X1 U14518 ( .A1(n13983), .A2(n11945), .B1(n15741), .B2(n11873), .ZN(
        n11946) );
  INV_X1 U14519 ( .A(n11946), .ZN(n11947) );
  OAI21_X1 U14520 ( .B1(n11948), .B2(n15739), .A(n11947), .ZN(P3_U3466) );
  XNOR2_X1 U14521 ( .A(n11958), .B(n13364), .ZN(n12024) );
  XNOR2_X1 U14522 ( .A(n12028), .B(n12024), .ZN(n11954) );
  NAND2_X1 U14523 ( .A1(n11952), .A2(n11951), .ZN(n11953) );
  AOI211_X1 U14524 ( .C1(n11954), .C2(n11953), .A(n13523), .B(n12025), .ZN(
        n11955) );
  INV_X1 U14525 ( .A(n11955), .ZN(n11960) );
  INV_X1 U14526 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n11956) );
  NOR2_X1 U14527 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11956), .ZN(n15617) );
  OAI22_X1 U14528 ( .A1(n12007), .A2(n13495), .B1(n12155), .B2(n13514), .ZN(
        n11957) );
  AOI211_X1 U14529 ( .C1(n11958), .C2(n13520), .A(n15617), .B(n11957), .ZN(
        n11959) );
  OAI211_X1 U14530 ( .C1(n12003), .C2(n13518), .A(n11960), .B(n11959), .ZN(
        P3_U3179) );
  AOI211_X1 U14531 ( .C1(n15321), .C2(n11963), .A(n11962), .B(n11961), .ZN(
        n11968) );
  AOI22_X1 U14532 ( .A1(n15217), .A2(n12189), .B1(n15330), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n11964) );
  OAI21_X1 U14533 ( .B1(n11968), .B2(n15330), .A(n11964), .ZN(P1_U3539) );
  INV_X1 U14534 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n11965) );
  OAI22_X1 U14535 ( .A1(n7139), .A2(n15089), .B1(n15324), .B2(n11965), .ZN(
        n11966) );
  INV_X1 U14536 ( .A(n11966), .ZN(n11967) );
  OAI21_X1 U14537 ( .B1(n11968), .B2(n10226), .A(n11967), .ZN(P1_U3492) );
  INV_X1 U14538 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11969) );
  MUX2_X1 U14539 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n11969), .S(n12217), .Z(
        n11970) );
  INV_X1 U14540 ( .A(n11970), .ZN(n11973) );
  NOR2_X1 U14541 ( .A1(n11972), .A2(n11973), .ZN(n12210) );
  AOI211_X1 U14542 ( .C1(n11973), .C2(n11972), .A(n15461), .B(n12210), .ZN(
        n11986) );
  INV_X1 U14543 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11974) );
  MUX2_X1 U14544 ( .A(n11974), .B(P2_REG1_REG_13__SCAN_IN), .S(n12217), .Z(
        n11980) );
  OR2_X1 U14545 ( .A1(n11975), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n11976) );
  NAND2_X1 U14546 ( .A1(n11977), .A2(n11976), .ZN(n11979) );
  INV_X1 U14547 ( .A(n12219), .ZN(n11978) );
  AOI211_X1 U14548 ( .C1(n11980), .C2(n11979), .A(n15465), .B(n11978), .ZN(
        n11985) );
  NAND2_X1 U14549 ( .A1(n15333), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n11982) );
  NAND2_X1 U14550 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n11981)
         );
  OAI211_X1 U14551 ( .C1(n15489), .C2(n11983), .A(n11982), .B(n11981), .ZN(
        n11984) );
  OR3_X1 U14552 ( .A1(n11986), .A2(n11985), .A3(n11984), .ZN(P2_U3227) );
  INV_X1 U14553 ( .A(n11987), .ZN(n11990) );
  INV_X1 U14554 ( .A(n14434), .ZN(n15537) );
  AOI211_X1 U14555 ( .C1(n11990), .C2(n15537), .A(n11989), .B(n11988), .ZN(
        n11997) );
  INV_X1 U14556 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11991) );
  OAI22_X1 U14557 ( .A1(n11992), .A2(n14517), .B1(n15543), .B2(n11991), .ZN(
        n11993) );
  INV_X1 U14558 ( .A(n11993), .ZN(n11994) );
  OAI21_X1 U14559 ( .B1(n11997), .B2(n15541), .A(n11994), .ZN(P2_U3457) );
  AOI22_X1 U14560 ( .A1(n11995), .A2(n14407), .B1(n15548), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n11996) );
  OAI21_X1 U14561 ( .B1(n11997), .B2(n15548), .A(n11996), .ZN(P2_U3508) );
  INV_X1 U14562 ( .A(n11998), .ZN(n11999) );
  OAI222_X1 U14563 ( .A1(n12959), .A2(n12000), .B1(n12957), .B2(n11999), .C1(
        n8713), .C2(P2_U3088), .ZN(P2_U3305) );
  OAI21_X1 U14564 ( .B1(n12002), .B2(n13322), .A(n12001), .ZN(n15723) );
  OAI22_X1 U14565 ( .A1(n13913), .A2(n15720), .B1(n12003), .B2(n13914), .ZN(
        n12012) );
  OAI211_X1 U14566 ( .C1(n12006), .C2(n12005), .A(n12004), .B(n13874), .ZN(
        n12010) );
  OAI22_X1 U14567 ( .A1(n12007), .A2(n15690), .B1(n12155), .B2(n15689), .ZN(
        n12008) );
  INV_X1 U14568 ( .A(n12008), .ZN(n12009) );
  NAND2_X1 U14569 ( .A1(n12010), .A2(n12009), .ZN(n15721) );
  MUX2_X1 U14570 ( .A(n15721), .B(P3_REG2_REG_6__SCAN_IN), .S(n13869), .Z(
        n12011) );
  AOI211_X1 U14571 ( .C1(n13919), .C2(n15723), .A(n12012), .B(n12011), .ZN(
        n12013) );
  INV_X1 U14572 ( .A(n12013), .ZN(P3_U3227) );
  INV_X1 U14573 ( .A(n12063), .ZN(n12015) );
  AOI21_X1 U14574 ( .B1(n12014), .B2(n12016), .A(n12015), .ZN(n12022) );
  INV_X1 U14575 ( .A(n12050), .ZN(n12019) );
  AOI22_X1 U14576 ( .A1(n14109), .A2(n14159), .B1(n14108), .B2(n14157), .ZN(
        n12018) );
  OAI211_X1 U14577 ( .C1(n12019), .C2(n14140), .A(n12018), .B(n12017), .ZN(
        n12020) );
  AOI21_X1 U14578 ( .B1(n12051), .B2(n14146), .A(n12020), .ZN(n12021) );
  OAI21_X1 U14579 ( .B1(n12022), .B2(n14148), .A(n12021), .ZN(P2_U3196) );
  XNOR2_X1 U14580 ( .A(n12023), .B(n11573), .ZN(n12126) );
  INV_X1 U14581 ( .A(n12024), .ZN(n12026) );
  XOR2_X1 U14582 ( .A(n12126), .B(n12128), .Z(n12027) );
  NAND2_X1 U14583 ( .A1(n12027), .A2(n13492), .ZN(n12032) );
  AND2_X1 U14584 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n15635) );
  OAI22_X1 U14585 ( .A1(n12304), .A2(n13514), .B1(n12028), .B2(n13495), .ZN(
        n12029) );
  AOI211_X1 U14586 ( .C1(n12030), .C2(n13520), .A(n15635), .B(n12029), .ZN(
        n12031) );
  OAI211_X1 U14587 ( .C1(n12033), .C2(n13518), .A(n12032), .B(n12031), .ZN(
        P3_U3153) );
  INV_X1 U14588 ( .A(n12058), .ZN(n12035) );
  NAND2_X1 U14589 ( .A1(n12964), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n12034) );
  OAI211_X1 U14590 ( .C1(n12035), .C2(n13377), .A(n12034), .B(n12846), .ZN(
        P1_U3332) );
  INV_X1 U14591 ( .A(n12036), .ZN(n12039) );
  OAI222_X1 U14592 ( .A1(n12850), .A2(n12039), .B1(n13382), .B2(n12038), .C1(
        P3_U3151), .C2(n12037), .ZN(P3_U3270) );
  XNOR2_X1 U14593 ( .A(n12040), .B(n12041), .ZN(n12047) );
  XNOR2_X1 U14594 ( .A(n12042), .B(n12041), .ZN(n12045) );
  OAI22_X1 U14595 ( .A1(n12043), .A2(n14323), .B1(n12314), .B2(n14325), .ZN(
        n12044) );
  AOI21_X1 U14596 ( .B1(n12045), .B2(n14358), .A(n12044), .ZN(n12046) );
  OAI21_X1 U14597 ( .B1(n12047), .B2(n10234), .A(n12046), .ZN(n15162) );
  INV_X1 U14598 ( .A(n15162), .ZN(n12056) );
  INV_X1 U14599 ( .A(n12047), .ZN(n15164) );
  INV_X1 U14600 ( .A(n12051), .ZN(n15161) );
  INV_X1 U14601 ( .A(n12048), .ZN(n12112) );
  INV_X1 U14602 ( .A(n12078), .ZN(n12049) );
  OAI211_X1 U14603 ( .C1(n15161), .C2(n12112), .A(n12049), .B(n14398), .ZN(
        n15160) );
  AOI22_X1 U14604 ( .A1(n6677), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n12050), 
        .B2(n15499), .ZN(n12053) );
  NAND2_X1 U14605 ( .A1(n12051), .A2(n14389), .ZN(n12052) );
  OAI211_X1 U14606 ( .C1(n15160), .C2(n14214), .A(n12053), .B(n12052), .ZN(
        n12054) );
  AOI21_X1 U14607 ( .B1(n15164), .B2(n14295), .A(n12054), .ZN(n12055) );
  OAI21_X1 U14608 ( .B1(n12056), .B2(n6677), .A(n12055), .ZN(P2_U3253) );
  NAND2_X1 U14609 ( .A1(n12058), .A2(n12057), .ZN(n12060) );
  OAI211_X1 U14610 ( .C1(n12061), .C2(n12959), .A(n12060), .B(n12059), .ZN(
        P2_U3304) );
  NAND2_X1 U14611 ( .A1(n12063), .A2(n12062), .ZN(n12065) );
  XNOR2_X1 U14612 ( .A(n12065), .B(n12064), .ZN(n12072) );
  INV_X1 U14613 ( .A(n12079), .ZN(n12069) );
  NAND2_X1 U14614 ( .A1(n14156), .A2(n14369), .ZN(n12067) );
  NAND2_X1 U14615 ( .A1(n14158), .A2(n14368), .ZN(n12066) );
  NAND2_X1 U14616 ( .A1(n12067), .A2(n12066), .ZN(n12076) );
  AOI22_X1 U14617 ( .A1(n14131), .A2(n12076), .B1(P2_REG3_REG_13__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12068) );
  OAI21_X1 U14618 ( .B1(n12069), .B2(n14140), .A(n12068), .ZN(n12070) );
  AOI21_X1 U14619 ( .B1(n12080), .B2(n14146), .A(n12070), .ZN(n12071) );
  OAI21_X1 U14620 ( .B1(n12072), .B2(n14148), .A(n12071), .ZN(P2_U3206) );
  XNOR2_X1 U14621 ( .A(n12073), .B(n12075), .ZN(n12242) );
  XOR2_X1 U14622 ( .A(n12075), .B(n12074), .Z(n12077) );
  AOI21_X1 U14623 ( .B1(n12077), .B2(n14358), .A(n12076), .ZN(n12241) );
  INV_X1 U14624 ( .A(n12241), .ZN(n12084) );
  OAI211_X1 U14625 ( .C1(n12246), .C2(n12078), .A(n14398), .B(n12317), .ZN(
        n12240) );
  AOI22_X1 U14626 ( .A1(n6677), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n12079), 
        .B2(n15499), .ZN(n12082) );
  NAND2_X1 U14627 ( .A1(n12080), .A2(n14389), .ZN(n12081) );
  OAI211_X1 U14628 ( .C1(n12240), .C2(n14214), .A(n12082), .B(n12081), .ZN(
        n12083) );
  AOI21_X1 U14629 ( .B1(n12084), .B2(n14397), .A(n12083), .ZN(n12085) );
  OAI21_X1 U14630 ( .B1(n14362), .B2(n12242), .A(n12085), .ZN(P2_U3252) );
  NAND2_X1 U14631 ( .A1(n12632), .A2(n13102), .ZN(n12090) );
  NAND2_X1 U14632 ( .A1(n14655), .A2(n13103), .ZN(n12089) );
  NAND2_X1 U14633 ( .A1(n12090), .A2(n12089), .ZN(n12091) );
  XNOR2_X1 U14634 ( .A(n12091), .B(n13115), .ZN(n12426) );
  OAI22_X1 U14635 ( .A1(n12093), .A2(n6681), .B1(n12092), .B2(n13112), .ZN(
        n12425) );
  XNOR2_X1 U14636 ( .A(n12426), .B(n12425), .ZN(n12094) );
  AOI21_X1 U14637 ( .B1(n12095), .B2(n12094), .A(n12428), .ZN(n12102) );
  OAI21_X1 U14638 ( .B1(n15205), .B2(n15207), .A(n12096), .ZN(n12097) );
  AOI21_X1 U14639 ( .B1(n14587), .B2(n14656), .A(n12097), .ZN(n12098) );
  OAI21_X1 U14640 ( .B1(n12099), .B2(n15222), .A(n12098), .ZN(n12100) );
  AOI21_X1 U14641 ( .B1(n15218), .B2(n12632), .A(n12100), .ZN(n12101) );
  OAI21_X1 U14642 ( .B1(n12102), .B2(n15212), .A(n12101), .ZN(P1_U3231) );
  XOR2_X1 U14643 ( .A(n12105), .B(n12103), .Z(n12250) );
  OAI21_X1 U14644 ( .B1(n12106), .B2(n12105), .A(n12104), .ZN(n12110) );
  OAI22_X1 U14645 ( .A1(n12108), .A2(n14323), .B1(n12107), .B2(n14325), .ZN(
        n12109) );
  AOI21_X1 U14646 ( .B1(n12110), .B2(n14358), .A(n12109), .ZN(n12111) );
  OAI21_X1 U14647 ( .B1(n12250), .B2(n10234), .A(n12111), .ZN(n12251) );
  NAND2_X1 U14648 ( .A1(n12251), .A2(n14397), .ZN(n12119) );
  AOI211_X1 U14649 ( .C1(n12257), .C2(n12113), .A(n12878), .B(n12112), .ZN(
        n12252) );
  INV_X1 U14650 ( .A(n12257), .ZN(n12116) );
  AOI22_X1 U14651 ( .A1(n6677), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n12114), 
        .B2(n15499), .ZN(n12115) );
  OAI21_X1 U14652 ( .B1(n12116), .B2(n15503), .A(n12115), .ZN(n12117) );
  AOI21_X1 U14653 ( .B1(n12252), .B2(n15498), .A(n12117), .ZN(n12118) );
  OAI211_X1 U14654 ( .C1(n12250), .C2(n14381), .A(n12119), .B(n12118), .ZN(
        P2_U3254) );
  INV_X1 U14655 ( .A(n12120), .ZN(n12124) );
  OAI222_X1 U14656 ( .A1(n12959), .A2(n12122), .B1(n12957), .B2(n12124), .C1(
        P2_U3088), .C2(n12121), .ZN(P2_U3303) );
  OAI222_X1 U14657 ( .A1(n12476), .A2(n12125), .B1(n13377), .B2(n12124), .C1(
        P1_U3086), .C2(n12123), .ZN(P1_U3331) );
  INV_X1 U14658 ( .A(n12126), .ZN(n12127) );
  XNOR2_X1 U14659 ( .A(n13364), .B(n12159), .ZN(n12296) );
  XNOR2_X1 U14660 ( .A(n12296), .B(n13533), .ZN(n12299) );
  XNOR2_X1 U14661 ( .A(n12300), .B(n12299), .ZN(n12134) );
  NOR2_X1 U14662 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12129), .ZN(n15651) );
  AOI21_X1 U14663 ( .B1(n13520), .B2(n12159), .A(n15651), .ZN(n12131) );
  INV_X1 U14664 ( .A(n13514), .ZN(n13482) );
  NAND2_X1 U14665 ( .A1(n13482), .A2(n13531), .ZN(n12130) );
  OAI211_X1 U14666 ( .C1(n12155), .C2(n13495), .A(n12131), .B(n12130), .ZN(
        n12132) );
  AOI21_X1 U14667 ( .B1(n13498), .B2(n12158), .A(n12132), .ZN(n12133) );
  OAI21_X1 U14668 ( .B1(n12134), .B2(n13523), .A(n12133), .ZN(P3_U3161) );
  OAI211_X1 U14669 ( .C1(n15117), .C2(n12135), .A(n15049), .B(n12179), .ZN(
        n15116) );
  XNOR2_X1 U14670 ( .A(n12136), .B(n12791), .ZN(n12143) );
  OAI21_X1 U14671 ( .B1(n12139), .B2(n12138), .A(n12137), .ZN(n12140) );
  NAND2_X1 U14672 ( .A1(n12140), .A2(n14980), .ZN(n12142) );
  AOI22_X1 U14673 ( .A1(n14975), .A2(n14651), .B1(n14653), .B2(n14974), .ZN(
        n12141) );
  OAI211_X1 U14674 ( .C1(n15286), .C2(n12143), .A(n12142), .B(n12141), .ZN(
        n15118) );
  NAND2_X1 U14675 ( .A1(n15118), .A2(n14913), .ZN(n12147) );
  OAI22_X1 U14676 ( .A1(n14913), .A2(n12144), .B1(n12454), .B2(n14982), .ZN(
        n12145) );
  AOI21_X1 U14677 ( .B1(n12653), .B2(n14992), .A(n12145), .ZN(n12146) );
  OAI211_X1 U14678 ( .C1(n14988), .C2(n15116), .A(n12147), .B(n12146), .ZN(
        P1_U3281) );
  INV_X1 U14679 ( .A(n12148), .ZN(n12151) );
  OAI222_X1 U14680 ( .A1(n12850), .A2(n12151), .B1(n13382), .B2(n12150), .C1(
        P3_U3151), .C2(n12149), .ZN(P3_U3269) );
  AOI21_X1 U14681 ( .B1(n13326), .B2(n12153), .A(n12152), .ZN(n12154) );
  OAI222_X1 U14682 ( .A1(n15689), .A2(n12357), .B1(n15690), .B2(n12155), .C1(
        n15696), .C2(n12154), .ZN(n12194) );
  INV_X1 U14683 ( .A(n12194), .ZN(n12164) );
  OAI21_X1 U14684 ( .B1(n12157), .B2(n13326), .A(n12156), .ZN(n12195) );
  AOI22_X1 U14685 ( .A1(n13901), .A2(n12159), .B1(n15702), .B2(n12158), .ZN(
        n12160) );
  OAI21_X1 U14686 ( .B1(n12161), .B2(n15703), .A(n12160), .ZN(n12162) );
  AOI21_X1 U14687 ( .B1(n12195), .B2(n13919), .A(n12162), .ZN(n12163) );
  OAI21_X1 U14688 ( .B1(n12164), .B2(n13921), .A(n12163), .ZN(P3_U3225) );
  INV_X1 U14689 ( .A(n12165), .ZN(n12573) );
  OAI222_X1 U14690 ( .A1(n12959), .A2(n12167), .B1(n12957), .B2(n12573), .C1(
        P2_U3088), .C2(n12166), .ZN(P2_U3302) );
  INV_X1 U14691 ( .A(n12168), .ZN(n12545) );
  OR2_X1 U14692 ( .A1(n12999), .A2(n14871), .ZN(n12170) );
  NAND2_X1 U14693 ( .A1(n14652), .A2(n14974), .ZN(n12169) );
  AND2_X1 U14694 ( .A1(n12170), .A2(n12169), .ZN(n12543) );
  INV_X1 U14695 ( .A(n12543), .ZN(n12174) );
  XNOR2_X1 U14696 ( .A(n12171), .B(n12178), .ZN(n12172) );
  NAND2_X1 U14697 ( .A1(n12172), .A2(n6966), .ZN(n12186) );
  INV_X1 U14698 ( .A(n12186), .ZN(n12173) );
  AOI211_X1 U14699 ( .C1(n15277), .C2(n12545), .A(n12174), .B(n12173), .ZN(
        n12184) );
  INV_X1 U14700 ( .A(n12175), .ZN(n12176) );
  OAI21_X1 U14701 ( .B1(n12178), .B2(n12177), .A(n12176), .ZN(n12188) );
  AOI21_X1 U14702 ( .B1(n12179), .B2(n12662), .A(n14958), .ZN(n12180) );
  NAND2_X1 U14703 ( .A1(n12180), .A2(n12227), .ZN(n12185) );
  AOI22_X1 U14704 ( .A1(n12662), .A2(n14992), .B1(n14962), .B2(
        P1_REG2_REG_13__SCAN_IN), .ZN(n12181) );
  OAI21_X1 U14705 ( .B1(n12185), .B2(n14988), .A(n12181), .ZN(n12182) );
  AOI21_X1 U14706 ( .B1(n12188), .B2(n15279), .A(n12182), .ZN(n12183) );
  OAI21_X1 U14707 ( .B1(n14962), .B2(n12184), .A(n12183), .ZN(P1_U3280) );
  NAND3_X1 U14708 ( .A1(n12186), .A2(n12543), .A3(n12185), .ZN(n12187) );
  AOI21_X1 U14709 ( .B1(n12188), .B2(n15321), .A(n12187), .ZN(n12193) );
  AOI22_X1 U14710 ( .A1(n12662), .A2(n12189), .B1(n15330), .B2(
        P1_REG1_REG_13__SCAN_IN), .ZN(n12190) );
  OAI21_X1 U14711 ( .B1(n12193), .B2(n15330), .A(n12190), .ZN(P1_U3541) );
  OAI22_X1 U14712 ( .A1(n12663), .A2(n15089), .B1(n15324), .B2(n7898), .ZN(
        n12191) );
  INV_X1 U14713 ( .A(n12191), .ZN(n12192) );
  OAI21_X1 U14714 ( .B1(n12193), .B2(n10226), .A(n12192), .ZN(P1_U3498) );
  AOI21_X1 U14715 ( .B1(n15724), .B2(n12195), .A(n12194), .ZN(n12201) );
  OAI22_X1 U14716 ( .A1(n13983), .A2(n13210), .B1(n15741), .B2(n11879), .ZN(
        n12196) );
  INV_X1 U14717 ( .A(n12196), .ZN(n12197) );
  OAI21_X1 U14718 ( .B1(n12201), .B2(n15739), .A(n12197), .ZN(P3_U3467) );
  INV_X1 U14719 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n12198) );
  OAI22_X1 U14720 ( .A1(n14033), .A2(n13210), .B1(n15734), .B2(n12198), .ZN(
        n12199) );
  INV_X1 U14721 ( .A(n12199), .ZN(n12200) );
  OAI21_X1 U14722 ( .B1(n12201), .B2(n15732), .A(n12200), .ZN(P3_U3414) );
  OAI21_X1 U14723 ( .B1(n12204), .B2(n12203), .A(n12202), .ZN(n12205) );
  NAND2_X1 U14724 ( .A1(n12205), .A2(n14103), .ZN(n12209) );
  NAND2_X1 U14725 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n12213)
         );
  INV_X1 U14726 ( .A(n12213), .ZN(n12207) );
  OAI22_X1 U14727 ( .A1(n12485), .A2(n14142), .B1(n14143), .B2(n12314), .ZN(
        n12206) );
  AOI211_X1 U14728 ( .C1(n12320), .C2(n14107), .A(n12207), .B(n12206), .ZN(
        n12208) );
  OAI211_X1 U14729 ( .C1(n12363), .C2(n14102), .A(n12209), .B(n12208), .ZN(
        P2_U3187) );
  NOR2_X1 U14730 ( .A1(n12211), .A2(n12214), .ZN(n14191) );
  OAI21_X1 U14731 ( .B1(n12212), .B2(P2_REG2_REG_14__SCAN_IN), .A(n15478), 
        .ZN(n12225) );
  OAI21_X1 U14732 ( .B1(n15489), .B2(n12214), .A(n12213), .ZN(n12215) );
  AOI21_X1 U14733 ( .B1(n15333), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n12215), 
        .ZN(n12224) );
  INV_X1 U14734 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n12216) );
  XNOR2_X1 U14735 ( .A(n14184), .B(n12216), .ZN(n12222) );
  NAND2_X1 U14736 ( .A1(n12217), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n12218) );
  NAND2_X1 U14737 ( .A1(n12219), .A2(n12218), .ZN(n12221) );
  INV_X1 U14738 ( .A(n14183), .ZN(n12220) );
  OAI211_X1 U14739 ( .C1(n12222), .C2(n12221), .A(n12220), .B(n15484), .ZN(
        n12223) );
  OAI211_X1 U14740 ( .C1(n14190), .C2(n12225), .A(n12224), .B(n12223), .ZN(
        P2_U3228) );
  OAI21_X1 U14741 ( .B1(n6801), .B2(n12795), .A(n12226), .ZN(n15228) );
  AOI21_X1 U14742 ( .B1(n15225), .B2(n12227), .A(n14958), .ZN(n12229) );
  INV_X1 U14743 ( .A(n12228), .ZN(n12419) );
  NAND2_X1 U14744 ( .A1(n12229), .A2(n12419), .ZN(n15226) );
  INV_X1 U14745 ( .A(n15226), .ZN(n12236) );
  OR2_X1 U14746 ( .A1(n15192), .A2(n14871), .ZN(n12231) );
  NAND2_X1 U14747 ( .A1(n14651), .A2(n14974), .ZN(n12230) );
  NAND2_X1 U14748 ( .A1(n12231), .A2(n12230), .ZN(n15223) );
  OAI22_X1 U14749 ( .A1(n14913), .A2(n11763), .B1(n15178), .B2(n14982), .ZN(
        n12232) );
  AOI21_X1 U14750 ( .B1(n14913), .B2(n15223), .A(n12232), .ZN(n12233) );
  OAI21_X1 U14751 ( .B1(n12234), .B2(n14949), .A(n12233), .ZN(n12235) );
  AOI21_X1 U14752 ( .B1(n12236), .B2(n14944), .A(n12235), .ZN(n12239) );
  XNOR2_X1 U14753 ( .A(n12237), .B(n12795), .ZN(n15230) );
  INV_X1 U14754 ( .A(n14969), .ZN(n15280) );
  NAND2_X1 U14755 ( .A1(n15230), .A2(n15280), .ZN(n12238) );
  OAI211_X1 U14756 ( .C1(n15228), .C2(n14862), .A(n12239), .B(n12238), .ZN(
        P1_U3279) );
  OAI211_X1 U14757 ( .C1(n12242), .C2(n14478), .A(n12241), .B(n12240), .ZN(
        n12248) );
  OAI22_X1 U14758 ( .A1(n12246), .A2(n14472), .B1(n15550), .B2(n11974), .ZN(
        n12243) );
  AOI21_X1 U14759 ( .B1(n12248), .B2(n15550), .A(n12243), .ZN(n12244) );
  INV_X1 U14760 ( .A(n12244), .ZN(P2_U3512) );
  INV_X1 U14761 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n12245) );
  OAI22_X1 U14762 ( .A1(n12246), .A2(n14517), .B1(n15543), .B2(n12245), .ZN(
        n12247) );
  AOI21_X1 U14763 ( .B1(n12248), .B2(n15543), .A(n12247), .ZN(n12249) );
  INV_X1 U14764 ( .A(n12249), .ZN(P2_U3469) );
  INV_X1 U14765 ( .A(n12250), .ZN(n12253) );
  AOI211_X1 U14766 ( .C1(n15537), .C2(n12253), .A(n12252), .B(n12251), .ZN(
        n12259) );
  AOI22_X1 U14767 ( .A1(n12257), .A2(n14407), .B1(n15548), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n12254) );
  OAI21_X1 U14768 ( .B1(n12259), .B2(n15548), .A(n12254), .ZN(P2_U3510) );
  INV_X1 U14769 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n12255) );
  NOR2_X1 U14770 ( .A1(n15543), .A2(n12255), .ZN(n12256) );
  AOI21_X1 U14771 ( .B1(n12257), .B2(n10162), .A(n12256), .ZN(n12258) );
  OAI21_X1 U14772 ( .B1(n12259), .B2(n15541), .A(n12258), .ZN(P2_U3463) );
  AOI21_X1 U14773 ( .B1(n12528), .B2(n12261), .A(n12329), .ZN(n12278) );
  NAND2_X1 U14774 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n12262), .ZN(n12264) );
  NAND2_X1 U14775 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n12265), .ZN(n12333) );
  OAI21_X1 U14776 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n12265), .A(n12333), 
        .ZN(n12276) );
  NOR2_X1 U14777 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12266), .ZN(n12509) );
  AOI21_X1 U14778 ( .B1(n15674), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n12509), 
        .ZN(n12267) );
  OAI21_X1 U14779 ( .B1(n15671), .B2(n12339), .A(n12267), .ZN(n12275) );
  INV_X1 U14780 ( .A(n12268), .ZN(n12269) );
  NOR2_X1 U14781 ( .A1(n12270), .A2(n12269), .ZN(n12272) );
  MUX2_X1 U14782 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n13629), .Z(n12340) );
  XNOR2_X1 U14783 ( .A(n12340), .B(n12339), .ZN(n12271) );
  AOI21_X1 U14784 ( .B1(n12272), .B2(n12271), .A(n12342), .ZN(n12273) );
  NOR2_X1 U14785 ( .A1(n12273), .A2(n15595), .ZN(n12274) );
  AOI211_X1 U14786 ( .C1(n15677), .C2(n12276), .A(n12275), .B(n12274), .ZN(
        n12277) );
  OAI21_X1 U14787 ( .B1(n12278), .B2(n15681), .A(n12277), .ZN(P3_U3193) );
  INV_X1 U14788 ( .A(n13323), .ZN(n13214) );
  XNOR2_X1 U14789 ( .A(n12279), .B(n13214), .ZN(n12288) );
  INV_X1 U14790 ( .A(n12288), .ZN(n12286) );
  OAI211_X1 U14791 ( .C1(n6813), .C2(n13323), .A(n12280), .B(n13874), .ZN(
        n12282) );
  AOI22_X1 U14792 ( .A1(n13530), .A2(n13877), .B1(n13880), .B2(n13533), .ZN(
        n12281) );
  NAND2_X1 U14793 ( .A1(n12282), .A2(n12281), .ZN(n12287) );
  NOR2_X1 U14794 ( .A1(n15703), .A2(n15661), .ZN(n12284) );
  OAI22_X1 U14795 ( .A1(n13913), .A2(n12295), .B1(n12308), .B2(n13914), .ZN(
        n12283) );
  AOI211_X1 U14796 ( .C1(n12287), .C2(n15703), .A(n12284), .B(n12283), .ZN(
        n12285) );
  OAI21_X1 U14797 ( .B1(n13905), .B2(n12286), .A(n12285), .ZN(P3_U3224) );
  AOI21_X1 U14798 ( .B1(n12288), .B2(n15724), .A(n12287), .ZN(n12294) );
  OAI22_X1 U14799 ( .A1(n13983), .A2(n12295), .B1(n15741), .B2(n11884), .ZN(
        n12289) );
  INV_X1 U14800 ( .A(n12289), .ZN(n12290) );
  OAI21_X1 U14801 ( .B1(n12294), .B2(n15739), .A(n12290), .ZN(P3_U3468) );
  INV_X1 U14802 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n12291) );
  OAI22_X1 U14803 ( .A1(n14033), .A2(n12295), .B1(n15734), .B2(n12291), .ZN(
        n12292) );
  INV_X1 U14804 ( .A(n12292), .ZN(n12293) );
  OAI21_X1 U14805 ( .B1(n12294), .B2(n15732), .A(n12293), .ZN(P3_U3417) );
  XNOR2_X1 U14806 ( .A(n12295), .B(n13364), .ZN(n12350) );
  XNOR2_X1 U14807 ( .A(n12357), .B(n12350), .ZN(n12302) );
  INV_X1 U14808 ( .A(n12296), .ZN(n12297) );
  NAND2_X1 U14809 ( .A1(n12301), .A2(n12302), .ZN(n12354) );
  OAI21_X1 U14810 ( .B1(n12302), .B2(n12301), .A(n12354), .ZN(n12303) );
  NAND2_X1 U14811 ( .A1(n12303), .A2(n13492), .ZN(n12307) );
  NOR2_X1 U14812 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8931), .ZN(n15673) );
  OAI22_X1 U14813 ( .A1(n12304), .A2(n13495), .B1(n12526), .B2(n13514), .ZN(
        n12305) );
  AOI211_X1 U14814 ( .C1(n9286), .C2(n13520), .A(n15673), .B(n12305), .ZN(
        n12306) );
  OAI211_X1 U14815 ( .C1(n12308), .C2(n13518), .A(n12307), .B(n12306), .ZN(
        P3_U3171) );
  INV_X1 U14816 ( .A(n12309), .ZN(n12311) );
  OAI222_X1 U14817 ( .A1(P3_U3151), .A2(n13629), .B1(n12850), .B2(n12311), 
        .C1(n12310), .C2(n13382), .ZN(P3_U3268) );
  XNOR2_X1 U14818 ( .A(n12312), .B(n12315), .ZN(n12313) );
  OAI222_X1 U14819 ( .A1(n14323), .A2(n12314), .B1(n14325), .B2(n12485), .C1(
        n12313), .C2(n14395), .ZN(n12364) );
  INV_X1 U14820 ( .A(n12364), .ZN(n12326) );
  XOR2_X1 U14821 ( .A(n12316), .B(n12315), .Z(n12366) );
  AOI21_X1 U14822 ( .B1(n12321), .B2(n12317), .A(n12878), .ZN(n12319) );
  INV_X1 U14823 ( .A(n12318), .ZN(n12377) );
  NAND2_X1 U14824 ( .A1(n12319), .A2(n12377), .ZN(n12362) );
  AOI22_X1 U14825 ( .A1(n6677), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n12320), 
        .B2(n15499), .ZN(n12323) );
  NAND2_X1 U14826 ( .A1(n12321), .A2(n14389), .ZN(n12322) );
  OAI211_X1 U14827 ( .C1(n12362), .C2(n14214), .A(n12323), .B(n12322), .ZN(
        n12324) );
  AOI21_X1 U14828 ( .B1(n12366), .B2(n15496), .A(n12324), .ZN(n12325) );
  OAI21_X1 U14829 ( .B1(n6677), .B2(n12326), .A(n12325), .ZN(P2_U3251) );
  AOI22_X1 U14830 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n13545), .B1(n13540), 
        .B2(n13916), .ZN(n12330) );
  AOI21_X1 U14831 ( .B1(n12331), .B2(n12330), .A(n13537), .ZN(n12349) );
  AOI22_X1 U14832 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n13540), .B1(n13545), 
        .B2(n8989), .ZN(n12336) );
  NAND2_X1 U14833 ( .A1(n12339), .A2(n12332), .ZN(n12334) );
  NAND2_X1 U14834 ( .A1(n12334), .A2(n12333), .ZN(n12335) );
  NAND2_X1 U14835 ( .A1(n12336), .A2(n12335), .ZN(n13544) );
  OAI21_X1 U14836 ( .B1(n12336), .B2(n12335), .A(n13544), .ZN(n12347) );
  INV_X1 U14837 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n12337) );
  NOR2_X1 U14838 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12337), .ZN(n13421) );
  AOI21_X1 U14839 ( .B1(n15674), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n13421), 
        .ZN(n12338) );
  OAI21_X1 U14840 ( .B1(n15671), .B2(n13540), .A(n12338), .ZN(n12346) );
  MUX2_X1 U14841 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n13629), .Z(n13541) );
  XNOR2_X1 U14842 ( .A(n13541), .B(n13540), .ZN(n12344) );
  NOR2_X1 U14843 ( .A1(n12340), .A2(n12339), .ZN(n12341) );
  OR2_X1 U14844 ( .A1(n12342), .A2(n12341), .ZN(n12343) );
  NOR3_X1 U14845 ( .A1(n12342), .A2(n12341), .A3(n12344), .ZN(n13539) );
  AOI211_X1 U14846 ( .C1(n12344), .C2(n12343), .A(n15595), .B(n13539), .ZN(
        n12345) );
  AOI211_X1 U14847 ( .C1(n15677), .C2(n12347), .A(n12346), .B(n12345), .ZN(
        n12348) );
  OAI21_X1 U14848 ( .B1(n12349), .B2(n15681), .A(n12348), .ZN(P3_U3194) );
  INV_X1 U14849 ( .A(n12350), .ZN(n12351) );
  NAND2_X1 U14850 ( .A1(n12351), .A2(n12357), .ZN(n12352) );
  AND2_X1 U14851 ( .A1(n12354), .A2(n12352), .ZN(n12356) );
  XNOR2_X1 U14852 ( .A(n12970), .B(n15730), .ZN(n12504) );
  XNOR2_X1 U14853 ( .A(n12504), .B(n12526), .ZN(n12355) );
  OAI211_X1 U14854 ( .C1(n12356), .C2(n12355), .A(n13492), .B(n12506), .ZN(
        n12361) );
  OAI22_X1 U14855 ( .A1(n12357), .A2(n13495), .B1(n13909), .B2(n13514), .ZN(
        n12358) );
  AOI211_X1 U14856 ( .C1(n15730), .C2(n13520), .A(n12359), .B(n12358), .ZN(
        n12360) );
  OAI211_X1 U14857 ( .C1(n12396), .C2(n13518), .A(n12361), .B(n12360), .ZN(
        P3_U3157) );
  OAI21_X1 U14858 ( .B1(n12363), .B2(n15525), .A(n12362), .ZN(n12365) );
  AOI211_X1 U14859 ( .C1(n12366), .C2(n15520), .A(n12365), .B(n12364), .ZN(
        n12369) );
  NAND2_X1 U14860 ( .A1(n15548), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n12367) );
  OAI21_X1 U14861 ( .B1(n12369), .B2(n15548), .A(n12367), .ZN(P2_U3513) );
  NAND2_X1 U14862 ( .A1(n15541), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n12368) );
  OAI21_X1 U14863 ( .B1(n12369), .B2(n15541), .A(n12368), .ZN(P2_U3472) );
  XNOR2_X1 U14864 ( .A(n12370), .B(n12374), .ZN(n14479) );
  INV_X1 U14865 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n12372) );
  INV_X1 U14866 ( .A(n12371), .ZN(n12404) );
  OAI22_X1 U14867 ( .A1(n14397), .A2(n12372), .B1(n12404), .B2(n14387), .ZN(
        n12373) );
  AOI21_X1 U14868 ( .B1(n12409), .B2(n14389), .A(n12373), .ZN(n12383) );
  XNOR2_X1 U14869 ( .A(n12375), .B(n7233), .ZN(n12376) );
  NAND2_X1 U14870 ( .A1(n12376), .A2(n14358), .ZN(n12379) );
  OAI21_X1 U14871 ( .B1(n12379), .B2(n6677), .A(n14214), .ZN(n12381) );
  XNOR2_X1 U14872 ( .A(n12409), .B(n12377), .ZN(n12380) );
  AOI22_X1 U14873 ( .A1(n14154), .A2(n14369), .B1(n14156), .B2(n14368), .ZN(
        n12378) );
  OAI211_X1 U14874 ( .C1(n12878), .C2(n12380), .A(n12379), .B(n12378), .ZN(
        n14480) );
  NAND2_X1 U14875 ( .A1(n12381), .A2(n14480), .ZN(n12382) );
  OAI211_X1 U14876 ( .C1(n14479), .C2(n14362), .A(n12383), .B(n12382), .ZN(
        P2_U3250) );
  INV_X1 U14877 ( .A(n12384), .ZN(n12388) );
  OAI222_X1 U14878 ( .A1(P2_U3088), .A2(n12386), .B1(n12957), .B2(n12388), 
        .C1(n12385), .C2(n12959), .ZN(P2_U3301) );
  OAI222_X1 U14879 ( .A1(n12476), .A2(n12389), .B1(n13377), .B2(n12388), .C1(
        n12387), .C2(P1_U3086), .ZN(P1_U3329) );
  XNOR2_X1 U14880 ( .A(n12390), .B(n13220), .ZN(n15727) );
  OAI21_X1 U14881 ( .B1(n12391), .B2(n13220), .A(n13874), .ZN(n12394) );
  AOI22_X1 U14882 ( .A1(n13880), .A2(n13531), .B1(n13529), .B2(n13877), .ZN(
        n12393) );
  OAI21_X1 U14883 ( .B1(n12394), .B2(n12392), .A(n12393), .ZN(n15728) );
  NOR2_X1 U14884 ( .A1(n15703), .A2(n12395), .ZN(n12399) );
  OAI22_X1 U14885 ( .A1(n13913), .A2(n12397), .B1(n12396), .B2(n13914), .ZN(
        n12398) );
  AOI211_X1 U14886 ( .C1(n15728), .C2(n15703), .A(n12399), .B(n12398), .ZN(
        n12400) );
  OAI21_X1 U14887 ( .B1(n13905), .B2(n15727), .A(n12400), .ZN(P3_U3223) );
  XNOR2_X1 U14888 ( .A(n12402), .B(n12401), .ZN(n12411) );
  OAI22_X1 U14889 ( .A1(n14140), .A2(n12404), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12403), .ZN(n12408) );
  OAI22_X1 U14890 ( .A1(n12406), .A2(n14143), .B1(n14142), .B2(n12405), .ZN(
        n12407) );
  AOI211_X1 U14891 ( .C1(n12409), .C2(n14146), .A(n12408), .B(n12407), .ZN(
        n12410) );
  OAI21_X1 U14892 ( .B1(n12411), .B2(n14148), .A(n12410), .ZN(P2_U3213) );
  XNOR2_X1 U14893 ( .A(n12412), .B(n12413), .ZN(n12516) );
  XNOR2_X1 U14894 ( .A(n12414), .B(n12413), .ZN(n12518) );
  NAND2_X1 U14895 ( .A1(n12518), .A2(n15279), .ZN(n12424) );
  OR2_X1 U14896 ( .A1(n14579), .A2(n14871), .ZN(n12416) );
  OR2_X1 U14897 ( .A1(n12999), .A2(n14869), .ZN(n12415) );
  AND2_X1 U14898 ( .A1(n12416), .A2(n12415), .ZN(n14634) );
  INV_X1 U14899 ( .A(n12417), .ZN(n14637) );
  AOI22_X1 U14900 ( .A1(n14962), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n14637), 
        .B2(n15277), .ZN(n12418) );
  OAI21_X1 U14901 ( .B1(n14962), .B2(n14634), .A(n12418), .ZN(n12422) );
  NAND2_X1 U14902 ( .A1(n13009), .A2(n12419), .ZN(n12420) );
  NAND3_X1 U14903 ( .A1(n12465), .A2(n15049), .A3(n12420), .ZN(n12515) );
  NOR2_X1 U14904 ( .A1(n12515), .A2(n14988), .ZN(n12421) );
  AOI211_X1 U14905 ( .C1(n14992), .C2(n13009), .A(n12422), .B(n12421), .ZN(
        n12423) );
  OAI211_X1 U14906 ( .C1(n12516), .C2(n14969), .A(n12424), .B(n12423), .ZN(
        P1_U3278) );
  NOR2_X1 U14907 ( .A1(n12426), .A2(n12425), .ZN(n12427) );
  NAND2_X1 U14908 ( .A1(n12641), .A2(n13102), .ZN(n12430) );
  NAND2_X1 U14909 ( .A1(n14654), .A2(n13103), .ZN(n12429) );
  NAND2_X1 U14910 ( .A1(n12430), .A2(n12429), .ZN(n12431) );
  XNOR2_X1 U14911 ( .A(n12431), .B(n13115), .ZN(n12439) );
  AND2_X1 U14912 ( .A1(n13068), .A2(n14654), .ZN(n12432) );
  AOI21_X1 U14913 ( .B1(n12641), .B2(n13103), .A(n12432), .ZN(n12437) );
  XNOR2_X1 U14914 ( .A(n12439), .B(n12437), .ZN(n15180) );
  NAND2_X1 U14915 ( .A1(n15217), .A2(n13102), .ZN(n12434) );
  NAND2_X1 U14916 ( .A1(n14653), .A2(n13103), .ZN(n12433) );
  NAND2_X1 U14917 ( .A1(n12434), .A2(n12433), .ZN(n12435) );
  XNOR2_X1 U14918 ( .A(n12435), .B(n13115), .ZN(n12441) );
  AND2_X1 U14919 ( .A1(n13068), .A2(n14653), .ZN(n12436) );
  AOI21_X1 U14920 ( .B1(n15217), .B2(n13103), .A(n12436), .ZN(n12442) );
  XNOR2_X1 U14921 ( .A(n12441), .B(n12442), .ZN(n15208) );
  INV_X1 U14922 ( .A(n12437), .ZN(n12438) );
  NAND2_X1 U14923 ( .A1(n12439), .A2(n12438), .ZN(n15209) );
  AND2_X1 U14924 ( .A1(n15208), .A2(n15209), .ZN(n12440) );
  NAND2_X1 U14925 ( .A1(n15210), .A2(n12440), .ZN(n15213) );
  INV_X1 U14926 ( .A(n12441), .ZN(n12443) );
  NAND2_X1 U14927 ( .A1(n12443), .A2(n12442), .ZN(n12444) );
  AND2_X1 U14928 ( .A1(n13068), .A2(n14652), .ZN(n12445) );
  AOI21_X1 U14929 ( .B1(n12653), .B2(n13103), .A(n12445), .ZN(n12535) );
  NAND2_X1 U14930 ( .A1(n12653), .A2(n13102), .ZN(n12447) );
  NAND2_X1 U14931 ( .A1(n14652), .A2(n13103), .ZN(n12446) );
  NAND2_X1 U14932 ( .A1(n12447), .A2(n12446), .ZN(n12448) );
  XNOR2_X1 U14933 ( .A(n12448), .B(n13115), .ZN(n12537) );
  XOR2_X1 U14934 ( .A(n12535), .B(n12537), .Z(n12450) );
  AOI21_X1 U14935 ( .B1(n12449), .B2(n12450), .A(n15212), .ZN(n12453) );
  INV_X1 U14936 ( .A(n12450), .ZN(n12451) );
  NAND2_X1 U14937 ( .A1(n12453), .A2(n12539), .ZN(n12459) );
  NOR2_X1 U14938 ( .A1(n15222), .A2(n12454), .ZN(n12457) );
  OAI21_X1 U14939 ( .B1(n15205), .B2(n15168), .A(n12455), .ZN(n12456) );
  AOI211_X1 U14940 ( .C1(n14587), .C2(n14653), .A(n12457), .B(n12456), .ZN(
        n12458) );
  OAI211_X1 U14941 ( .C1(n15117), .C2(n15186), .A(n12459), .B(n12458), .ZN(
        P1_U3224) );
  INV_X1 U14942 ( .A(n12460), .ZN(n12461) );
  AOI21_X1 U14943 ( .B1(n12798), .B2(n12462), .A(n12461), .ZN(n15072) );
  OAI21_X1 U14944 ( .B1(n12464), .B2(n12798), .A(n12463), .ZN(n15067) );
  NAND2_X1 U14945 ( .A1(n15067), .A2(n15279), .ZN(n12473) );
  AOI211_X1 U14946 ( .C1(n15200), .C2(n12465), .A(n14958), .B(n6798), .ZN(
        n15068) );
  AOI22_X1 U14947 ( .A1(n14962), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n12466), 
        .B2(n15277), .ZN(n12470) );
  OR2_X1 U14948 ( .A1(n15192), .A2(n14869), .ZN(n12468) );
  NAND2_X1 U14949 ( .A1(n14973), .A2(n14975), .ZN(n12467) );
  NAND2_X1 U14950 ( .A1(n12468), .A2(n12467), .ZN(n15069) );
  NAND2_X1 U14951 ( .A1(n14913), .A2(n15069), .ZN(n12469) );
  OAI211_X1 U14952 ( .C1(n13017), .C2(n14949), .A(n12470), .B(n12469), .ZN(
        n12471) );
  AOI21_X1 U14953 ( .B1(n15068), .B2(n14944), .A(n12471), .ZN(n12472) );
  OAI211_X1 U14954 ( .C1(n15072), .C2(n14969), .A(n12473), .B(n12472), .ZN(
        P1_U3277) );
  INV_X1 U14955 ( .A(n12474), .ZN(n12478) );
  OAI222_X1 U14956 ( .A1(n12476), .A2(n12475), .B1(n13377), .B2(n12478), .C1(
        n10214), .C2(P1_U3086), .ZN(P1_U3328) );
  OAI222_X1 U14957 ( .A1(n12959), .A2(n12479), .B1(n12957), .B2(n12478), .C1(
        n12477), .C2(P2_U3088), .ZN(P2_U3300) );
  OAI21_X1 U14958 ( .B1(n7283), .B2(n12481), .A(n12480), .ZN(n14477) );
  XNOR2_X1 U14959 ( .A(n12483), .B(n12482), .ZN(n12484) );
  OAI222_X1 U14960 ( .A1(n14325), .A2(n14129), .B1(n14323), .B2(n12485), .C1(
        n12484), .C2(n14395), .ZN(n14473) );
  NAND2_X1 U14961 ( .A1(n14473), .A2(n14397), .ZN(n12493) );
  INV_X1 U14962 ( .A(n12564), .ZN(n12486) );
  AOI211_X1 U14963 ( .C1(n14475), .C2(n12487), .A(n12878), .B(n12486), .ZN(
        n14474) );
  INV_X1 U14964 ( .A(n14475), .ZN(n12488) );
  NOR2_X1 U14965 ( .A1(n12488), .A2(n15503), .ZN(n12491) );
  OAI22_X1 U14966 ( .A1(n14397), .A2(n12489), .B1(n12500), .B2(n14387), .ZN(
        n12490) );
  AOI211_X1 U14967 ( .C1(n14474), .C2(n15498), .A(n12491), .B(n12490), .ZN(
        n12492) );
  OAI211_X1 U14968 ( .C1(n14477), .C2(n14362), .A(n12493), .B(n12492), .ZN(
        P2_U3249) );
  INV_X1 U14969 ( .A(n12494), .ZN(n12994) );
  AOI21_X1 U14970 ( .B1(n14525), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n12495), 
        .ZN(n12496) );
  OAI21_X1 U14971 ( .B1(n12994), .B2(n14531), .A(n12496), .ZN(P2_U3299) );
  AOI21_X1 U14972 ( .B1(n12498), .B2(n12497), .A(n14091), .ZN(n12503) );
  AOI22_X1 U14973 ( .A1(n14109), .A2(n14155), .B1(n14108), .B2(n14153), .ZN(
        n12499) );
  NAND2_X1 U14974 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n15458)
         );
  OAI211_X1 U14975 ( .C1(n14140), .C2(n12500), .A(n12499), .B(n15458), .ZN(
        n12501) );
  AOI21_X1 U14976 ( .B1(n14475), .B2(n14146), .A(n12501), .ZN(n12502) );
  OAI21_X1 U14977 ( .B1(n12503), .B2(n14148), .A(n12502), .ZN(P2_U3198) );
  INV_X1 U14978 ( .A(n12504), .ZN(n12505) );
  XNOR2_X1 U14979 ( .A(n15150), .B(n13364), .ZN(n12507) );
  NAND2_X1 U14980 ( .A1(n7174), .A2(n12896), .ZN(n12508) );
  XNOR2_X1 U14981 ( .A(n12508), .B(n13909), .ZN(n12514) );
  AOI21_X1 U14982 ( .B1(n13483), .B2(n13482), .A(n12509), .ZN(n12511) );
  NAND2_X1 U14983 ( .A1(n13530), .A2(n13516), .ZN(n12510) );
  OAI211_X1 U14984 ( .C1(n13518), .C2(n12527), .A(n12511), .B(n12510), .ZN(
        n12512) );
  AOI21_X1 U14985 ( .B1(n12530), .B2(n13520), .A(n12512), .ZN(n12513) );
  OAI21_X1 U14986 ( .B1(n12514), .B2(n13523), .A(n12513), .ZN(P3_U3176) );
  INV_X1 U14987 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n12519) );
  OAI211_X1 U14988 ( .C1(n12516), .C2(n15286), .A(n14634), .B(n12515), .ZN(
        n12517) );
  AOI21_X1 U14989 ( .B1(n12518), .B2(n15321), .A(n12517), .ZN(n12521) );
  MUX2_X1 U14990 ( .A(n12519), .B(n12521), .S(n15324), .Z(n12520) );
  OAI21_X1 U14991 ( .B1(n8211), .B2(n15089), .A(n12520), .ZN(P1_U3504) );
  MUX2_X1 U14992 ( .A(n15258), .B(n12521), .S(n15332), .Z(n12522) );
  OAI21_X1 U14993 ( .B1(n8211), .B2(n15046), .A(n12522), .ZN(P1_U3543) );
  XOR2_X1 U14994 ( .A(n13327), .B(n12523), .Z(n15151) );
  XNOR2_X1 U14995 ( .A(n12524), .B(n13327), .ZN(n12525) );
  OAI222_X1 U14996 ( .A1(n15689), .A2(n13897), .B1(n15690), .B2(n12526), .C1(
        n12525), .C2(n15696), .ZN(n15153) );
  NAND2_X1 U14997 ( .A1(n15153), .A2(n15703), .ZN(n12532) );
  OAI22_X1 U14998 ( .A1(n15703), .A2(n12528), .B1(n12527), .B2(n13914), .ZN(
        n12529) );
  AOI21_X1 U14999 ( .B1(n12530), .B2(n13901), .A(n12529), .ZN(n12531) );
  OAI211_X1 U15000 ( .C1(n13905), .C2(n15151), .A(n12532), .B(n12531), .ZN(
        P3_U3222) );
  OAI22_X1 U15001 ( .A1(n12663), .A2(n13111), .B1(n15168), .B2(n6681), .ZN(
        n12533) );
  XNOR2_X1 U15002 ( .A(n12533), .B(n13115), .ZN(n13001) );
  AND2_X1 U15003 ( .A1(n13068), .A2(n14651), .ZN(n12534) );
  AOI21_X1 U15004 ( .B1(n12662), .B2(n13103), .A(n12534), .ZN(n13002) );
  XNOR2_X1 U15005 ( .A(n13001), .B(n13002), .ZN(n12541) );
  INV_X1 U15006 ( .A(n12535), .ZN(n12536) );
  NAND2_X1 U15007 ( .A1(n12537), .A2(n12536), .ZN(n12538) );
  OAI211_X1 U15008 ( .C1(n12541), .C2(n12540), .A(n13005), .B(n15179), .ZN(
        n12547) );
  OAI21_X1 U15009 ( .B1(n12543), .B2(n14633), .A(n12542), .ZN(n12544) );
  AOI21_X1 U15010 ( .B1(n12545), .B2(n14636), .A(n12544), .ZN(n12546) );
  OAI211_X1 U15011 ( .C1(n12663), .C2(n15186), .A(n12547), .B(n12546), .ZN(
        P1_U3234) );
  AOI21_X1 U15012 ( .B1(n12548), .B2(n12553), .A(n15286), .ZN(n12552) );
  OAI22_X1 U15013 ( .A1(n12549), .A2(n14871), .B1(n14579), .B2(n14869), .ZN(
        n12550) );
  AOI21_X1 U15014 ( .B1(n12552), .B2(n12551), .A(n12550), .ZN(n15065) );
  XNOR2_X1 U15015 ( .A(n12554), .B(n12553), .ZN(n15062) );
  NAND2_X1 U15016 ( .A1(n15062), .A2(n15279), .ZN(n12559) );
  OAI22_X1 U15017 ( .A1(n14913), .A2(n14722), .B1(n12555), .B2(n14982), .ZN(
        n12557) );
  OAI211_X1 U15018 ( .C1(n6798), .C2(n13022), .A(n14985), .B(n15049), .ZN(
        n15063) );
  NOR2_X1 U15019 ( .A1(n15063), .A2(n14988), .ZN(n12556) );
  AOI211_X1 U15020 ( .C1(n14992), .C2(n14573), .A(n12557), .B(n12556), .ZN(
        n12558) );
  OAI211_X1 U15021 ( .C1(n14962), .C2(n15065), .A(n12559), .B(n12558), .ZN(
        P1_U3276) );
  XOR2_X1 U15022 ( .A(n12560), .B(n12561), .Z(n14469) );
  INV_X1 U15023 ( .A(n14469), .ZN(n12571) );
  XNOR2_X1 U15024 ( .A(n12562), .B(n12561), .ZN(n12563) );
  AOI22_X1 U15025 ( .A1(n14367), .A2(n14369), .B1(n14368), .B2(n14154), .ZN(
        n14097) );
  OAI21_X1 U15026 ( .B1(n12563), .B2(n14395), .A(n14097), .ZN(n14467) );
  AOI211_X1 U15027 ( .C1(n12565), .C2(n12564), .A(n12878), .B(n6800), .ZN(
        n14468) );
  NAND2_X1 U15028 ( .A1(n14468), .A2(n15498), .ZN(n12568) );
  INV_X1 U15029 ( .A(n12566), .ZN(n14099) );
  AOI22_X1 U15030 ( .A1(n6677), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n14099), 
        .B2(n15499), .ZN(n12567) );
  OAI211_X1 U15031 ( .C1(n14518), .C2(n15503), .A(n12568), .B(n12567), .ZN(
        n12569) );
  AOI21_X1 U15032 ( .B1(n14467), .B2(n14397), .A(n12569), .ZN(n12570) );
  OAI21_X1 U15033 ( .B1(n12571), .B2(n14362), .A(n12570), .ZN(P2_U3248) );
  OAI222_X1 U15034 ( .A1(n13374), .A2(n12574), .B1(n13377), .B2(n12573), .C1(
        P1_U3086), .C2(n12572), .ZN(P1_U3330) );
  OR2_X1 U15035 ( .A1(n14663), .A2(n14664), .ZN(n12584) );
  NAND2_X1 U15036 ( .A1(n12764), .A2(n12578), .ZN(n12581) );
  NAND2_X1 U15037 ( .A1(n12578), .A2(n12577), .ZN(n12582) );
  AND2_X1 U15038 ( .A1(n12769), .A2(n15274), .ZN(n12583) );
  NAND3_X1 U15039 ( .A1(n14663), .A2(n12583), .A3(n6682), .ZN(n12580) );
  OAI211_X1 U15040 ( .C1(n14663), .C2(n12582), .A(n15295), .B(n6682), .ZN(
        n12586) );
  NOR2_X1 U15041 ( .A1(n12584), .A2(n12583), .ZN(n12585) );
  NAND2_X1 U15042 ( .A1(n12588), .A2(n8157), .ZN(n12592) );
  MUX2_X1 U15043 ( .A(n14662), .B(n12589), .S(n12764), .Z(n12590) );
  OAI21_X1 U15044 ( .B1(n7742), .B2(n15301), .A(n12590), .ZN(n12591) );
  NAND3_X1 U15045 ( .A1(n12592), .A2(n12778), .A3(n12591), .ZN(n12598) );
  AND2_X1 U15046 ( .A1(n14661), .A2(n12764), .ZN(n12595) );
  NOR2_X1 U15047 ( .A1(n14661), .A2(n12764), .ZN(n12594) );
  MUX2_X1 U15048 ( .A(n12595), .B(n12594), .S(n12593), .Z(n12596) );
  INV_X1 U15049 ( .A(n12596), .ZN(n12597) );
  NAND2_X1 U15050 ( .A1(n12598), .A2(n12597), .ZN(n12602) );
  MUX2_X1 U15051 ( .A(n14660), .B(n12599), .S(n6683), .Z(n12603) );
  NAND2_X1 U15052 ( .A1(n12602), .A2(n12603), .ZN(n12601) );
  MUX2_X1 U15053 ( .A(n14660), .B(n12599), .S(n12764), .Z(n12600) );
  NAND2_X1 U15054 ( .A1(n12601), .A2(n12600), .ZN(n12607) );
  INV_X1 U15055 ( .A(n12602), .ZN(n12605) );
  INV_X1 U15056 ( .A(n12603), .ZN(n12604) );
  MUX2_X1 U15057 ( .A(n14659), .B(n12608), .S(n12764), .Z(n12610) );
  MUX2_X1 U15058 ( .A(n14659), .B(n12608), .S(n6682), .Z(n12609) );
  MUX2_X1 U15059 ( .A(n14658), .B(n12611), .S(n6682), .Z(n12615) );
  NAND2_X1 U15060 ( .A1(n12614), .A2(n12615), .ZN(n12613) );
  MUX2_X1 U15061 ( .A(n14658), .B(n12611), .S(n12764), .Z(n12612) );
  NAND2_X1 U15062 ( .A1(n12613), .A2(n12612), .ZN(n12619) );
  INV_X1 U15063 ( .A(n12614), .ZN(n12617) );
  INV_X1 U15064 ( .A(n12615), .ZN(n12616) );
  NAND2_X1 U15065 ( .A1(n12617), .A2(n12616), .ZN(n12618) );
  MUX2_X1 U15066 ( .A(n14657), .B(n12620), .S(n12764), .Z(n12622) );
  MUX2_X1 U15067 ( .A(n14657), .B(n12620), .S(n6683), .Z(n12621) );
  MUX2_X1 U15068 ( .A(n14656), .B(n12623), .S(n6683), .Z(n12627) );
  NAND2_X1 U15069 ( .A1(n12626), .A2(n12627), .ZN(n12625) );
  MUX2_X1 U15070 ( .A(n14656), .B(n12623), .S(n12764), .Z(n12624) );
  NAND2_X1 U15071 ( .A1(n12625), .A2(n12624), .ZN(n12631) );
  INV_X1 U15072 ( .A(n12626), .ZN(n12629) );
  INV_X1 U15073 ( .A(n12627), .ZN(n12628) );
  NAND2_X1 U15074 ( .A1(n12629), .A2(n12628), .ZN(n12630) );
  NAND2_X1 U15075 ( .A1(n12631), .A2(n12630), .ZN(n12635) );
  MUX2_X1 U15076 ( .A(n14655), .B(n12632), .S(n12764), .Z(n12636) );
  NAND2_X1 U15077 ( .A1(n12635), .A2(n12636), .ZN(n12634) );
  MUX2_X1 U15078 ( .A(n14655), .B(n12632), .S(n6683), .Z(n12633) );
  NAND2_X1 U15079 ( .A1(n12634), .A2(n12633), .ZN(n12640) );
  INV_X1 U15080 ( .A(n12635), .ZN(n12638) );
  INV_X1 U15081 ( .A(n12636), .ZN(n12637) );
  NAND2_X1 U15082 ( .A1(n12638), .A2(n12637), .ZN(n12639) );
  MUX2_X1 U15083 ( .A(n14654), .B(n12641), .S(n6683), .Z(n12643) );
  MUX2_X1 U15084 ( .A(n14654), .B(n12641), .S(n12764), .Z(n12642) );
  INV_X1 U15085 ( .A(n12643), .ZN(n12644) );
  MUX2_X1 U15086 ( .A(n14653), .B(n15217), .S(n12764), .Z(n12648) );
  NAND2_X1 U15087 ( .A1(n12647), .A2(n12648), .ZN(n12646) );
  MUX2_X1 U15088 ( .A(n14653), .B(n15217), .S(n6682), .Z(n12645) );
  NAND2_X1 U15089 ( .A1(n12646), .A2(n12645), .ZN(n12652) );
  INV_X1 U15090 ( .A(n12647), .ZN(n12650) );
  INV_X1 U15091 ( .A(n12648), .ZN(n12649) );
  NAND2_X1 U15092 ( .A1(n12650), .A2(n12649), .ZN(n12651) );
  NAND2_X1 U15093 ( .A1(n12652), .A2(n12651), .ZN(n12656) );
  MUX2_X1 U15094 ( .A(n14652), .B(n12653), .S(n6682), .Z(n12657) );
  NAND2_X1 U15095 ( .A1(n12656), .A2(n12657), .ZN(n12655) );
  MUX2_X1 U15096 ( .A(n14652), .B(n12653), .S(n12764), .Z(n12654) );
  NAND2_X1 U15097 ( .A1(n12655), .A2(n12654), .ZN(n12661) );
  INV_X1 U15098 ( .A(n12656), .ZN(n12659) );
  INV_X1 U15099 ( .A(n12657), .ZN(n12658) );
  NAND2_X1 U15100 ( .A1(n12659), .A2(n12658), .ZN(n12660) );
  MUX2_X1 U15101 ( .A(n14651), .B(n12662), .S(n12764), .Z(n12665) );
  MUX2_X1 U15102 ( .A(n15168), .B(n12663), .S(n6682), .Z(n12664) );
  AOI21_X1 U15103 ( .B1(n12675), .B2(n12666), .A(n6682), .ZN(n12667) );
  AND2_X1 U15104 ( .A1(n12670), .A2(n12669), .ZN(n12671) );
  OAI22_X1 U15105 ( .A1(n12672), .A2(n7543), .B1(n12764), .B2(n12671), .ZN(
        n12678) );
  MUX2_X1 U15106 ( .A(n14973), .B(n14573), .S(n12764), .Z(n12684) );
  OR2_X1 U15107 ( .A1(n12684), .A2(n12673), .ZN(n12674) );
  INV_X1 U15108 ( .A(n12675), .ZN(n12676) );
  MUX2_X1 U15109 ( .A(n14579), .B(n13017), .S(n12764), .Z(n12681) );
  MUX2_X1 U15110 ( .A(n14649), .B(n15200), .S(n6683), .Z(n12680) );
  AOI22_X1 U15111 ( .A1(n12676), .A2(n6683), .B1(n12681), .B2(n12680), .ZN(
        n12677) );
  NAND3_X1 U15112 ( .A1(n12678), .A2(n12679), .A3(n12677), .ZN(n12690) );
  INV_X1 U15113 ( .A(n12679), .ZN(n12682) );
  NAND3_X1 U15114 ( .A1(n14972), .A2(n12684), .A3(n12683), .ZN(n12688) );
  MUX2_X1 U15115 ( .A(n14648), .B(n14991), .S(n12764), .Z(n12686) );
  NAND2_X1 U15116 ( .A1(n12686), .A2(n12685), .ZN(n12687) );
  MUX2_X1 U15117 ( .A(n12692), .B(n12691), .S(n6682), .Z(n12693) );
  NAND2_X1 U15118 ( .A1(n12694), .A2(n12693), .ZN(n12697) );
  MUX2_X1 U15119 ( .A(n14647), .B(n15048), .S(n12764), .Z(n12698) );
  NAND2_X1 U15120 ( .A1(n12697), .A2(n12698), .ZN(n12696) );
  MUX2_X1 U15121 ( .A(n14647), .B(n15048), .S(n6682), .Z(n12695) );
  NAND2_X1 U15122 ( .A1(n12696), .A2(n12695), .ZN(n12702) );
  INV_X1 U15123 ( .A(n12697), .ZN(n12700) );
  INV_X1 U15124 ( .A(n12698), .ZN(n12699) );
  NAND2_X1 U15125 ( .A1(n12700), .A2(n12699), .ZN(n12701) );
  MUX2_X1 U15126 ( .A(n14646), .B(n14928), .S(n6683), .Z(n12704) );
  MUX2_X1 U15127 ( .A(n14646), .B(n14928), .S(n12764), .Z(n12703) );
  INV_X1 U15128 ( .A(n12704), .ZN(n12705) );
  INV_X1 U15129 ( .A(n12709), .ZN(n12707) );
  MUX2_X1 U15130 ( .A(n15035), .B(n14888), .S(n6682), .Z(n12708) );
  INV_X1 U15131 ( .A(n12708), .ZN(n12706) );
  NAND2_X1 U15132 ( .A1(n12709), .A2(n12708), .ZN(n12711) );
  MUX2_X1 U15133 ( .A(n15035), .B(n14888), .S(n12764), .Z(n12710) );
  NAND2_X1 U15134 ( .A1(n12711), .A2(n12710), .ZN(n12712) );
  MUX2_X1 U15135 ( .A(n14645), .B(n14898), .S(n6683), .Z(n12715) );
  MUX2_X1 U15136 ( .A(n14645), .B(n14898), .S(n12764), .Z(n12714) );
  INV_X1 U15137 ( .A(n12715), .ZN(n12716) );
  MUX2_X1 U15138 ( .A(n14887), .B(n14883), .S(n12764), .Z(n12720) );
  NAND2_X1 U15139 ( .A1(n12719), .A2(n12720), .ZN(n12718) );
  MUX2_X1 U15140 ( .A(n14887), .B(n14883), .S(n6682), .Z(n12717) );
  NAND2_X1 U15141 ( .A1(n12718), .A2(n12717), .ZN(n12724) );
  INV_X1 U15142 ( .A(n12719), .ZN(n12722) );
  INV_X1 U15143 ( .A(n12720), .ZN(n12721) );
  MUX2_X1 U15144 ( .A(n14644), .B(n15017), .S(n6683), .Z(n12726) );
  MUX2_X1 U15145 ( .A(n14644), .B(n15017), .S(n12764), .Z(n12725) );
  INV_X1 U15146 ( .A(n12726), .ZN(n12727) );
  MUX2_X1 U15147 ( .A(n14622), .B(n14643), .S(n6683), .Z(n12731) );
  NAND2_X1 U15148 ( .A1(n12730), .A2(n12731), .ZN(n12729) );
  MUX2_X1 U15149 ( .A(n14643), .B(n14622), .S(n6682), .Z(n12728) );
  NAND2_X1 U15150 ( .A1(n12729), .A2(n12728), .ZN(n12735) );
  INV_X1 U15151 ( .A(n12730), .ZN(n12733) );
  INV_X1 U15152 ( .A(n12731), .ZN(n12732) );
  NAND2_X1 U15153 ( .A1(n12733), .A2(n12732), .ZN(n12734) );
  MUX2_X1 U15154 ( .A(n14803), .B(n14537), .S(n6683), .Z(n12737) );
  MUX2_X1 U15155 ( .A(n14803), .B(n14537), .S(n12764), .Z(n12736) );
  INV_X1 U15156 ( .A(n12737), .ZN(n12738) );
  MUX2_X1 U15157 ( .A(n14642), .B(n15004), .S(n12764), .Z(n12742) );
  NAND2_X1 U15158 ( .A1(n12741), .A2(n12742), .ZN(n12740) );
  MUX2_X1 U15159 ( .A(n14642), .B(n15004), .S(n6682), .Z(n12739) );
  NAND2_X1 U15160 ( .A1(n12740), .A2(n12739), .ZN(n12746) );
  INV_X1 U15161 ( .A(n12741), .ZN(n12744) );
  INV_X1 U15162 ( .A(n12742), .ZN(n12743) );
  NAND2_X1 U15163 ( .A1(n12744), .A2(n12743), .ZN(n12745) );
  MUX2_X1 U15164 ( .A(n14802), .B(n12747), .S(n6683), .Z(n12749) );
  MUX2_X1 U15165 ( .A(n14802), .B(n12747), .S(n12764), .Z(n12748) );
  INV_X1 U15166 ( .A(n12749), .ZN(n12750) );
  NAND2_X1 U15167 ( .A1(n12960), .A2(n12766), .ZN(n12753) );
  NAND2_X1 U15168 ( .A1(n12751), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12752) );
  INV_X1 U15169 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n12757) );
  NAND2_X1 U15170 ( .A1(n7763), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n12756) );
  NAND2_X1 U15171 ( .A1(n12754), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n12755) );
  OAI211_X1 U15172 ( .C1(n12758), .C2(n12757), .A(n12756), .B(n12755), .ZN(
        n14773) );
  INV_X1 U15173 ( .A(n12759), .ZN(n12760) );
  AOI22_X1 U15174 ( .A1(n14773), .A2(n12764), .B1(n12760), .B2(n12813), .ZN(
        n12761) );
  OAI22_X1 U15175 ( .A1(n15079), .A2(n12764), .B1(n12762), .B2(n12761), .ZN(
        n12824) );
  INV_X1 U15176 ( .A(n12762), .ZN(n14641) );
  OAI21_X1 U15177 ( .B1(n14773), .B2(n12763), .A(n14641), .ZN(n12765) );
  MUX2_X1 U15178 ( .A(n12765), .B(n15079), .S(n12764), .Z(n12825) );
  NOR2_X1 U15179 ( .A1(n12824), .A2(n12825), .ZN(n12828) );
  INV_X1 U15180 ( .A(n12828), .ZN(n12774) );
  NAND2_X1 U15181 ( .A1(n14521), .A2(n12766), .ZN(n12768) );
  NAND2_X1 U15182 ( .A1(n12751), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n12767) );
  XNOR2_X1 U15183 ( .A(n14774), .B(n14773), .ZN(n12814) );
  OR2_X1 U15184 ( .A1(n12769), .A2(n14764), .ZN(n12773) );
  NAND2_X1 U15185 ( .A1(n12771), .A2(n12770), .ZN(n12772) );
  AND2_X1 U15186 ( .A1(n12773), .A2(n12772), .ZN(n12815) );
  INV_X1 U15187 ( .A(n12775), .ZN(n12779) );
  NAND2_X1 U15188 ( .A1(n14664), .A2(n15274), .ZN(n12776) );
  AND2_X1 U15189 ( .A1(n12777), .A2(n12776), .ZN(n15285) );
  NAND4_X1 U15190 ( .A1(n12779), .A2(n15285), .A3(n12778), .A4(n8157), .ZN(
        n12782) );
  NOR3_X1 U15191 ( .A1(n12782), .A2(n12781), .A3(n12780), .ZN(n12786) );
  NAND4_X1 U15192 ( .A1(n12786), .A2(n12785), .A3(n12784), .A4(n12783), .ZN(
        n12787) );
  NOR4_X1 U15193 ( .A1(n12790), .A2(n12789), .A3(n12788), .A4(n12787), .ZN(
        n12793) );
  NAND4_X1 U15194 ( .A1(n12794), .A2(n12793), .A3(n12792), .A4(n12791), .ZN(
        n12796) );
  NOR4_X1 U15195 ( .A1(n12798), .A2(n12797), .A3(n12796), .A4(n12795), .ZN(
        n12799) );
  NAND3_X1 U15196 ( .A1(n14953), .A2(n12799), .A3(n14972), .ZN(n12800) );
  NOR4_X1 U15197 ( .A1(n12801), .A2(n14907), .A3(n12800), .A4(n14934), .ZN(
        n12804) );
  NAND4_X1 U15198 ( .A1(n12804), .A2(n12803), .A3(n14850), .A4(n12802), .ZN(
        n12805) );
  NOR4_X1 U15199 ( .A1(n14809), .A2(n12807), .A3(n12806), .A4(n12805), .ZN(
        n12810) );
  XNOR2_X1 U15200 ( .A(n7145), .B(n14641), .ZN(n12809) );
  NAND4_X1 U15201 ( .A1(n12814), .A2(n12810), .A3(n12809), .A4(n12808), .ZN(
        n12811) );
  XNOR2_X1 U15202 ( .A(n12811), .B(n14764), .ZN(n12832) );
  NAND2_X1 U15203 ( .A1(n12813), .A2(n12812), .ZN(n12831) );
  INV_X1 U15204 ( .A(n12814), .ZN(n12816) );
  INV_X1 U15205 ( .A(n12815), .ZN(n12819) );
  AND2_X1 U15206 ( .A1(n12819), .A2(n12831), .ZN(n12823) );
  NAND2_X1 U15207 ( .A1(n12816), .A2(n12823), .ZN(n12820) );
  MUX2_X1 U15208 ( .A(n14773), .B(n14774), .S(n6682), .Z(n12818) );
  NOR2_X1 U15209 ( .A1(n14774), .A2(n14773), .ZN(n12817) );
  NOR2_X1 U15210 ( .A1(n12818), .A2(n12817), .ZN(n12821) );
  MUX2_X1 U15211 ( .A(n12820), .B(n12819), .S(n12821), .Z(n12830) );
  INV_X1 U15212 ( .A(n12821), .ZN(n12822) );
  INV_X1 U15213 ( .A(n12824), .ZN(n12827) );
  INV_X1 U15214 ( .A(n12825), .ZN(n12826) );
  NOR2_X1 U15215 ( .A1(n12827), .A2(n12826), .ZN(n12835) );
  AOI22_X1 U15216 ( .A1(n12834), .A2(n12828), .B1(n7602), .B2(n12835), .ZN(
        n12829) );
  OAI211_X1 U15217 ( .C1(n12832), .C2(n12831), .A(n12830), .B(n12829), .ZN(
        n12833) );
  INV_X1 U15218 ( .A(n12833), .ZN(n12839) );
  INV_X1 U15219 ( .A(n12834), .ZN(n12836) );
  NOR2_X1 U15220 ( .A1(n12836), .A2(n12835), .ZN(n12837) );
  OAI211_X1 U15221 ( .C1(n12841), .C2(n12840), .A(n12839), .B(n12838), .ZN(
        n12842) );
  INV_X1 U15222 ( .A(n12842), .ZN(n12847) );
  NOR3_X1 U15223 ( .A1(n12843), .A2(n10214), .A3(n14869), .ZN(n12845) );
  OAI21_X1 U15224 ( .B1(n12846), .B2(n15097), .A(P1_B_REG_SCAN_IN), .ZN(n12844) );
  OAI22_X1 U15225 ( .A1(n12847), .A2(n12846), .B1(n12845), .B2(n12844), .ZN(
        P1_U3242) );
  INV_X1 U15226 ( .A(n12848), .ZN(n12849) );
  OAI222_X1 U15227 ( .A1(n14049), .A2(n12851), .B1(P3_U3151), .B2(n13354), 
        .C1(n12850), .C2(n12849), .ZN(P3_U3267) );
  INV_X1 U15228 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n12852) );
  OAI22_X1 U15229 ( .A1(n12853), .A2(n15503), .B1(n14397), .B2(n12852), .ZN(
        n12855) );
  AND2_X1 U15230 ( .A1(n12859), .A2(n12858), .ZN(n12860) );
  XNOR2_X1 U15231 ( .A(n14306), .B(n12882), .ZN(n12863) );
  NOR2_X1 U15232 ( .A1(n14326), .A2(n14398), .ZN(n14058) );
  INV_X1 U15233 ( .A(n12862), .ZN(n12864) );
  XNOR2_X1 U15234 ( .A(n14430), .B(n12877), .ZN(n12867) );
  NAND2_X1 U15235 ( .A1(n14151), .A2(n12878), .ZN(n12866) );
  NOR2_X1 U15236 ( .A1(n12867), .A2(n12866), .ZN(n12868) );
  AOI21_X1 U15237 ( .B1(n12867), .B2(n12866), .A(n12868), .ZN(n14105) );
  INV_X1 U15238 ( .A(n12868), .ZN(n12869) );
  XNOR2_X1 U15239 ( .A(n14085), .B(n12877), .ZN(n12871) );
  NAND2_X1 U15240 ( .A1(n14254), .A2(n12878), .ZN(n12870) );
  NOR2_X1 U15241 ( .A1(n12871), .A2(n12870), .ZN(n12872) );
  AOI21_X1 U15242 ( .B1(n12871), .B2(n12870), .A(n12872), .ZN(n14083) );
  INV_X1 U15243 ( .A(n12872), .ZN(n12873) );
  NAND2_X1 U15244 ( .A1(n14229), .A2(n12878), .ZN(n12875) );
  XNOR2_X1 U15245 ( .A(n14420), .B(n12882), .ZN(n12874) );
  XOR2_X1 U15246 ( .A(n12875), .B(n12874), .Z(n14137) );
  INV_X1 U15247 ( .A(n12874), .ZN(n12876) );
  XNOR2_X1 U15248 ( .A(n14415), .B(n12877), .ZN(n12880) );
  NAND2_X1 U15249 ( .A1(n14255), .A2(n12878), .ZN(n12879) );
  NOR2_X1 U15250 ( .A1(n12880), .A2(n12879), .ZN(n12881) );
  AOI21_X1 U15251 ( .B1(n12880), .B2(n12879), .A(n12881), .ZN(n14051) );
  NAND2_X1 U15252 ( .A1(n14228), .A2(n12878), .ZN(n12883) );
  XNOR2_X1 U15253 ( .A(n12883), .B(n12882), .ZN(n12884) );
  XNOR2_X1 U15254 ( .A(n12892), .B(n12884), .ZN(n12885) );
  XNOR2_X1 U15255 ( .A(n12886), .B(n12885), .ZN(n12894) );
  INV_X1 U15256 ( .A(n12887), .ZN(n12890) );
  AOI22_X1 U15257 ( .A1(n14131), .A2(n12888), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12889) );
  OAI21_X1 U15258 ( .B1(n12890), .B2(n14140), .A(n12889), .ZN(n12891) );
  AOI21_X1 U15259 ( .B1(n12892), .B2(n14146), .A(n12891), .ZN(n12893) );
  OAI21_X1 U15260 ( .B1(n12894), .B2(n14148), .A(n12893), .ZN(P2_U3192) );
  XNOR2_X1 U15261 ( .A(n13715), .B(n11573), .ZN(n12895) );
  NOR2_X1 U15262 ( .A1(n12895), .A2(n13526), .ZN(n12973) );
  AOI21_X1 U15263 ( .B1(n12895), .B2(n13526), .A(n12973), .ZN(n12981) );
  XNOR2_X1 U15264 ( .A(n12970), .B(n12897), .ZN(n12898) );
  NOR2_X1 U15265 ( .A1(n13483), .A2(n12898), .ZN(n12899) );
  AOI21_X1 U15266 ( .B1(n12898), .B2(n13483), .A(n12899), .ZN(n13419) );
  NAND2_X1 U15267 ( .A1(n13418), .A2(n13419), .ZN(n13417) );
  INV_X1 U15268 ( .A(n12899), .ZN(n12900) );
  NAND2_X1 U15269 ( .A1(n13417), .A2(n12900), .ZN(n13481) );
  XNOR2_X1 U15270 ( .A(n15142), .B(n11573), .ZN(n12901) );
  NOR2_X1 U15271 ( .A1(n12901), .A2(n13879), .ZN(n13477) );
  NAND2_X1 U15272 ( .A1(n12901), .A2(n13879), .ZN(n13478) );
  XNOR2_X1 U15273 ( .A(n14032), .B(n13364), .ZN(n12902) );
  XNOR2_X1 U15274 ( .A(n12902), .B(n13896), .ZN(n13384) );
  NAND2_X1 U15275 ( .A1(n12902), .A2(n13528), .ZN(n12903) );
  XNOR2_X1 U15276 ( .A(n13521), .B(n12970), .ZN(n13511) );
  NAND2_X1 U15277 ( .A1(n13511), .A2(n13878), .ZN(n12904) );
  XNOR2_X1 U15278 ( .A(n13971), .B(n11573), .ZN(n12906) );
  XNOR2_X1 U15279 ( .A(n12906), .B(n13843), .ZN(n13439) );
  NAND2_X1 U15280 ( .A1(n13440), .A2(n13439), .ZN(n12909) );
  INV_X1 U15281 ( .A(n12906), .ZN(n12907) );
  NAND2_X1 U15282 ( .A1(n12907), .A2(n13843), .ZN(n12908) );
  NAND2_X1 U15283 ( .A1(n12909), .A2(n12908), .ZN(n13447) );
  XNOR2_X1 U15284 ( .A(n13967), .B(n11573), .ZN(n12910) );
  XNOR2_X1 U15285 ( .A(n12910), .B(n13852), .ZN(n13448) );
  NAND2_X1 U15286 ( .A1(n13447), .A2(n13448), .ZN(n12913) );
  INV_X1 U15287 ( .A(n12910), .ZN(n12911) );
  NAND2_X1 U15288 ( .A1(n12911), .A2(n13852), .ZN(n12912) );
  XNOR2_X1 U15289 ( .A(n13960), .B(n13364), .ZN(n12914) );
  XNOR2_X1 U15290 ( .A(n12914), .B(n13842), .ZN(n13503) );
  INV_X1 U15291 ( .A(n12914), .ZN(n12915) );
  XNOR2_X1 U15292 ( .A(n13817), .B(n11573), .ZN(n12922) );
  XNOR2_X1 U15293 ( .A(n12922), .B(n12923), .ZN(n13466) );
  XNOR2_X1 U15294 ( .A(n13804), .B(n13364), .ZN(n12917) );
  INV_X1 U15295 ( .A(n12917), .ZN(n12916) );
  NAND2_X1 U15296 ( .A1(n12916), .A2(n13812), .ZN(n12925) );
  INV_X1 U15297 ( .A(n12925), .ZN(n12918) );
  XNOR2_X1 U15298 ( .A(n12917), .B(n13812), .ZN(n13469) );
  XNOR2_X1 U15299 ( .A(n13414), .B(n11573), .ZN(n12920) );
  NAND2_X1 U15300 ( .A1(n12920), .A2(n13801), .ZN(n12930) );
  OAI21_X1 U15301 ( .B1(n12920), .B2(n13801), .A(n12930), .ZN(n13410) );
  INV_X1 U15302 ( .A(n13410), .ZN(n12928) );
  INV_X1 U15303 ( .A(n12921), .ZN(n12927) );
  INV_X1 U15304 ( .A(n12922), .ZN(n12924) );
  NAND2_X1 U15305 ( .A1(n12924), .A2(n12923), .ZN(n13467) );
  AND2_X1 U15306 ( .A1(n13467), .A2(n12925), .ZN(n12926) );
  NAND2_X1 U15307 ( .A1(n13406), .A2(n12929), .ZN(n13407) );
  NAND2_X1 U15308 ( .A1(n13407), .A2(n12930), .ZN(n12933) );
  XNOR2_X1 U15309 ( .A(n12931), .B(n13364), .ZN(n12932) );
  NAND2_X1 U15310 ( .A1(n12933), .A2(n12932), .ZN(n12937) );
  OR2_X1 U15311 ( .A1(n12933), .A2(n12932), .ZN(n13489) );
  NAND2_X1 U15312 ( .A1(n12934), .A2(n13489), .ZN(n13490) );
  NAND2_X1 U15313 ( .A1(n13490), .A2(n12937), .ZN(n12941) );
  XNOR2_X1 U15314 ( .A(n13766), .B(n11573), .ZN(n12940) );
  INV_X1 U15315 ( .A(n12940), .ZN(n12936) );
  NOR2_X1 U15316 ( .A1(n9301), .A2(n12936), .ZN(n12935) );
  NAND2_X1 U15317 ( .A1(n12935), .A2(n13489), .ZN(n12939) );
  NAND2_X1 U15318 ( .A1(n13392), .A2(n13455), .ZN(n12945) );
  XNOR2_X1 U15319 ( .A(n13937), .B(n13364), .ZN(n12942) );
  NAND2_X1 U15320 ( .A1(n12942), .A2(n13723), .ZN(n13429) );
  INV_X1 U15321 ( .A(n12942), .ZN(n12943) );
  NAND2_X1 U15322 ( .A1(n12943), .A2(n13763), .ZN(n12944) );
  NAND2_X1 U15323 ( .A1(n12945), .A2(n13456), .ZN(n13428) );
  NAND2_X1 U15324 ( .A1(n13428), .A2(n13429), .ZN(n12949) );
  XNOR2_X1 U15325 ( .A(n13427), .B(n11573), .ZN(n12946) );
  NAND2_X1 U15326 ( .A1(n12946), .A2(n13750), .ZN(n12977) );
  INV_X1 U15327 ( .A(n12946), .ZN(n12947) );
  NAND2_X1 U15328 ( .A1(n12947), .A2(n13527), .ZN(n12948) );
  OAI21_X1 U15329 ( .B1(n12981), .B2(n12950), .A(n12974), .ZN(n12951) );
  NAND2_X1 U15330 ( .A1(n12951), .A2(n13492), .ZN(n12955) );
  AOI22_X1 U15331 ( .A1(n13527), .A2(n13516), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12952) );
  OAI21_X1 U15332 ( .B1(n13703), .B2(n13514), .A(n12952), .ZN(n12953) );
  AOI21_X1 U15333 ( .B1(n13713), .B2(n13498), .A(n12953), .ZN(n12954) );
  OAI211_X1 U15334 ( .C1(n13715), .C2(n13501), .A(n12955), .B(n12954), .ZN(
        P3_U3180) );
  OAI222_X1 U15335 ( .A1(n12959), .A2(n12958), .B1(n12957), .B2(n12956), .C1(
        n14201), .C2(P2_U3088), .ZN(P2_U3308) );
  INV_X1 U15336 ( .A(n12960), .ZN(n12969) );
  OAI222_X1 U15337 ( .A1(n14531), .A2(n12969), .B1(P2_U3088), .B2(n7310), .C1(
        n13139), .C2(n12959), .ZN(P2_U3297) );
  NAND3_X1 U15338 ( .A1(n12962), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n12967) );
  NAND2_X1 U15339 ( .A1(n14521), .A2(n12963), .ZN(n12966) );
  NAND2_X1 U15340 ( .A1(n12964), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n12965) );
  OAI211_X1 U15341 ( .C1(n12961), .C2(n12967), .A(n12966), .B(n12965), .ZN(
        P1_U3324) );
  INV_X1 U15342 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n13140) );
  XNOR2_X1 U15343 ( .A(n12971), .B(n12970), .ZN(n12972) );
  NOR2_X1 U15344 ( .A1(n12972), .A2(n13299), .ZN(n13361) );
  AOI21_X1 U15345 ( .B1(n12972), .B2(n13299), .A(n13361), .ZN(n12980) );
  INV_X1 U15346 ( .A(n12973), .ZN(n12975) );
  INV_X1 U15347 ( .A(n12980), .ZN(n12976) );
  AND2_X1 U15348 ( .A1(n12977), .A2(n12979), .ZN(n12978) );
  NAND2_X1 U15349 ( .A1(n13432), .A2(n12978), .ZN(n12985) );
  INV_X1 U15350 ( .A(n12979), .ZN(n12983) );
  AND2_X1 U15351 ( .A1(n12981), .A2(n12980), .ZN(n12982) );
  NAND2_X1 U15352 ( .A1(n12985), .A2(n12984), .ZN(n13363) );
  NAND2_X1 U15353 ( .A1(n12986), .A2(n13363), .ZN(n12987) );
  NAND2_X1 U15354 ( .A1(n12987), .A2(n13492), .ZN(n12992) );
  INV_X1 U15355 ( .A(n13127), .ZN(n12989) );
  AOI22_X1 U15356 ( .A1(n13526), .A2(n13516), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12988) );
  OAI21_X1 U15357 ( .B1(n12989), .B2(n13518), .A(n12988), .ZN(n12990) );
  AOI21_X1 U15358 ( .B1(n13525), .B2(n13482), .A(n12990), .ZN(n12991) );
  OAI211_X1 U15359 ( .C1(n13300), .C2(n13501), .A(n12992), .B(n12991), .ZN(
        P3_U3154) );
  OAI222_X1 U15360 ( .A1(n13374), .A2(n12995), .B1(n13377), .B2(n12994), .C1(
        P1_U3086), .C2(n12993), .ZN(P1_U3327) );
  NAND2_X1 U15361 ( .A1(n15225), .A2(n13102), .ZN(n12997) );
  OR2_X1 U15362 ( .A1(n12999), .A2(n6681), .ZN(n12996) );
  NAND2_X1 U15363 ( .A1(n12997), .A2(n12996), .ZN(n12998) );
  XNOR2_X1 U15364 ( .A(n12998), .B(n6706), .ZN(n13007) );
  NOR2_X1 U15365 ( .A1(n12999), .A2(n13112), .ZN(n13000) );
  AOI21_X1 U15366 ( .B1(n15225), .B2(n13103), .A(n13000), .ZN(n13006) );
  XNOR2_X1 U15367 ( .A(n13007), .B(n13006), .ZN(n15169) );
  INV_X1 U15368 ( .A(n13001), .ZN(n13003) );
  NOR2_X1 U15369 ( .A1(n13003), .A2(n13002), .ZN(n15170) );
  NOR2_X1 U15370 ( .A1(n15169), .A2(n15170), .ZN(n13004) );
  NAND2_X1 U15371 ( .A1(n13007), .A2(n13006), .ZN(n13008) );
  NAND2_X1 U15372 ( .A1(n13009), .A2(n13102), .ZN(n13011) );
  OR2_X1 U15373 ( .A1(n15192), .A2(n6681), .ZN(n13010) );
  NAND2_X1 U15374 ( .A1(n13011), .A2(n13010), .ZN(n13012) );
  XNOR2_X1 U15375 ( .A(n13012), .B(n6706), .ZN(n13014) );
  INV_X1 U15376 ( .A(n13014), .ZN(n13013) );
  XNOR2_X1 U15377 ( .A(n13015), .B(n13013), .ZN(n14632) );
  OAI22_X1 U15378 ( .A1(n8211), .A2(n6681), .B1(n15192), .B2(n13112), .ZN(
        n14631) );
  NOR2_X1 U15379 ( .A1(n13015), .A2(n13014), .ZN(n15194) );
  OAI22_X1 U15380 ( .A1(n13017), .A2(n13111), .B1(n14579), .B2(n6681), .ZN(
        n13016) );
  XNOR2_X1 U15381 ( .A(n13016), .B(n13115), .ZN(n13020) );
  OAI22_X1 U15382 ( .A1(n13017), .A2(n6681), .B1(n14579), .B2(n13112), .ZN(
        n13019) );
  XNOR2_X1 U15383 ( .A(n13020), .B(n13019), .ZN(n15193) );
  OR2_X1 U15384 ( .A1(n13020), .A2(n13019), .ZN(n13021) );
  OAI22_X1 U15385 ( .A1(n13022), .A2(n6681), .B1(n15191), .B2(n13112), .ZN(
        n13027) );
  NAND2_X1 U15386 ( .A1(n14573), .A2(n13102), .ZN(n13024) );
  NAND2_X1 U15387 ( .A1(n14973), .A2(n13103), .ZN(n13023) );
  NAND2_X1 U15388 ( .A1(n13024), .A2(n13023), .ZN(n13025) );
  XNOR2_X1 U15389 ( .A(n13025), .B(n13115), .ZN(n13026) );
  XOR2_X1 U15390 ( .A(n13027), .B(n13026), .Z(n14576) );
  INV_X1 U15391 ( .A(n13026), .ZN(n13029) );
  INV_X1 U15392 ( .A(n13027), .ZN(n13028) );
  NAND2_X1 U15393 ( .A1(n14991), .A2(n13102), .ZN(n13031) );
  NAND2_X1 U15394 ( .A1(n14648), .A2(n13103), .ZN(n13030) );
  NAND2_X1 U15395 ( .A1(n13031), .A2(n13030), .ZN(n13032) );
  XNOR2_X1 U15396 ( .A(n13032), .B(n13115), .ZN(n13033) );
  AOI22_X1 U15397 ( .A1(n14991), .A2(n13103), .B1(n13068), .B2(n14648), .ZN(
        n13034) );
  XNOR2_X1 U15398 ( .A(n13033), .B(n13034), .ZN(n14612) );
  NAND2_X1 U15399 ( .A1(n14613), .A2(n14612), .ZN(n13037) );
  INV_X1 U15400 ( .A(n13033), .ZN(n13035) );
  NAND2_X1 U15401 ( .A1(n13035), .A2(n13034), .ZN(n13036) );
  NAND2_X1 U15402 ( .A1(n13037), .A2(n13036), .ZN(n14546) );
  NOR2_X1 U15403 ( .A1(n14597), .A2(n13112), .ZN(n13038) );
  AOI21_X1 U15404 ( .B1(n14965), .B2(n13103), .A(n13038), .ZN(n13044) );
  NAND2_X1 U15405 ( .A1(n14965), .A2(n13102), .ZN(n13040) );
  OR2_X1 U15406 ( .A1(n14597), .A2(n6681), .ZN(n13039) );
  NAND2_X1 U15407 ( .A1(n13040), .A2(n13039), .ZN(n13041) );
  XNOR2_X1 U15408 ( .A(n13041), .B(n13115), .ZN(n13043) );
  XOR2_X1 U15409 ( .A(n13044), .B(n13043), .Z(n14547) );
  INV_X1 U15410 ( .A(n14547), .ZN(n13042) );
  INV_X1 U15411 ( .A(n13043), .ZN(n13045) );
  OR2_X1 U15412 ( .A1(n13045), .A2(n13044), .ZN(n13046) );
  AND2_X1 U15413 ( .A1(n14647), .A2(n13068), .ZN(n13047) );
  AOI21_X1 U15414 ( .B1(n15048), .B2(n13103), .A(n13047), .ZN(n13050) );
  AOI22_X1 U15415 ( .A1(n15048), .A2(n13102), .B1(n13103), .B2(n14647), .ZN(
        n13048) );
  XNOR2_X1 U15416 ( .A(n13048), .B(n13115), .ZN(n13049) );
  XOR2_X1 U15417 ( .A(n13050), .B(n13049), .Z(n14594) );
  INV_X1 U15418 ( .A(n13049), .ZN(n13052) );
  INV_X1 U15419 ( .A(n13050), .ZN(n13051) );
  NAND2_X1 U15420 ( .A1(n13052), .A2(n13051), .ZN(n13053) );
  OAI22_X1 U15421 ( .A1(n15090), .A2(n13111), .B1(n14596), .B2(n6681), .ZN(
        n13054) );
  XNOR2_X1 U15422 ( .A(n13054), .B(n13115), .ZN(n13055) );
  OAI22_X1 U15423 ( .A1(n15090), .A2(n6681), .B1(n14596), .B2(n13112), .ZN(
        n13056) );
  XNOR2_X1 U15424 ( .A(n13055), .B(n13056), .ZN(n14558) );
  INV_X1 U15425 ( .A(n13055), .ZN(n13058) );
  INV_X1 U15426 ( .A(n13056), .ZN(n13057) );
  NAND2_X1 U15427 ( .A1(n13058), .A2(n13057), .ZN(n13059) );
  AND2_X1 U15428 ( .A1(n13068), .A2(n14888), .ZN(n13060) );
  AOI21_X1 U15429 ( .B1(n15035), .B2(n13103), .A(n13060), .ZN(n13062) );
  AOI22_X1 U15430 ( .A1(n15035), .A2(n13102), .B1(n13103), .B2(n14888), .ZN(
        n13061) );
  XNOR2_X1 U15431 ( .A(n13061), .B(n13115), .ZN(n13063) );
  XOR2_X1 U15432 ( .A(n13062), .B(n13063), .Z(n14604) );
  NAND2_X1 U15433 ( .A1(n13063), .A2(n13062), .ZN(n13064) );
  NAND2_X1 U15434 ( .A1(n14898), .A2(n13102), .ZN(n13066) );
  NAND2_X1 U15435 ( .A1(n14645), .A2(n13103), .ZN(n13065) );
  NAND2_X1 U15436 ( .A1(n13066), .A2(n13065), .ZN(n13067) );
  XNOR2_X1 U15437 ( .A(n13067), .B(n13115), .ZN(n13069) );
  AOI22_X1 U15438 ( .A1(n14898), .A2(n13103), .B1(n13068), .B2(n14645), .ZN(
        n13070) );
  XNOR2_X1 U15439 ( .A(n13069), .B(n13070), .ZN(n14540) );
  INV_X1 U15440 ( .A(n13069), .ZN(n13071) );
  OAI22_X1 U15441 ( .A1(n14880), .A2(n6681), .B1(n13072), .B2(n13112), .ZN(
        n13077) );
  NAND2_X1 U15442 ( .A1(n14883), .A2(n13102), .ZN(n13074) );
  NAND2_X1 U15443 ( .A1(n14887), .A2(n13103), .ZN(n13073) );
  NAND2_X1 U15444 ( .A1(n13074), .A2(n13073), .ZN(n13075) );
  XNOR2_X1 U15445 ( .A(n13075), .B(n13115), .ZN(n13076) );
  XOR2_X1 U15446 ( .A(n13077), .B(n13076), .Z(n14586) );
  NAND2_X1 U15447 ( .A1(n14585), .A2(n14586), .ZN(n13081) );
  INV_X1 U15448 ( .A(n13076), .ZN(n13079) );
  INV_X1 U15449 ( .A(n13077), .ZN(n13078) );
  NAND2_X1 U15450 ( .A1(n13079), .A2(n13078), .ZN(n13080) );
  NAND2_X1 U15451 ( .A1(n13081), .A2(n13080), .ZN(n14565) );
  OAI22_X1 U15452 ( .A1(n14859), .A2(n6681), .B1(n14872), .B2(n13112), .ZN(
        n13086) );
  NAND2_X1 U15453 ( .A1(n15017), .A2(n13102), .ZN(n13083) );
  NAND2_X1 U15454 ( .A1(n14644), .A2(n13103), .ZN(n13082) );
  NAND2_X1 U15455 ( .A1(n13083), .A2(n13082), .ZN(n13084) );
  XNOR2_X1 U15456 ( .A(n13084), .B(n13115), .ZN(n13085) );
  XOR2_X1 U15457 ( .A(n13086), .B(n13085), .Z(n14566) );
  NAND2_X1 U15458 ( .A1(n14565), .A2(n14566), .ZN(n13090) );
  INV_X1 U15459 ( .A(n13085), .ZN(n13088) );
  INV_X1 U15460 ( .A(n13086), .ZN(n13087) );
  NAND2_X1 U15461 ( .A1(n13088), .A2(n13087), .ZN(n13089) );
  NAND2_X1 U15462 ( .A1(n13090), .A2(n13089), .ZN(n14620) );
  OAI22_X1 U15463 ( .A1(n14841), .A2(n6681), .B1(n13091), .B2(n13112), .ZN(
        n13096) );
  NAND2_X1 U15464 ( .A1(n14622), .A2(n13102), .ZN(n13093) );
  NAND2_X1 U15465 ( .A1(n14643), .A2(n13103), .ZN(n13092) );
  NAND2_X1 U15466 ( .A1(n13093), .A2(n13092), .ZN(n13094) );
  XNOR2_X1 U15467 ( .A(n13094), .B(n13115), .ZN(n13095) );
  XOR2_X1 U15468 ( .A(n13096), .B(n13095), .Z(n14621) );
  INV_X1 U15469 ( .A(n13095), .ZN(n13098) );
  INV_X1 U15470 ( .A(n13096), .ZN(n13097) );
  NAND2_X1 U15471 ( .A1(n13098), .A2(n13097), .ZN(n13099) );
  OAI22_X1 U15472 ( .A1(n14826), .A2(n6681), .B1(n13101), .B2(n13112), .ZN(
        n13108) );
  NAND2_X1 U15473 ( .A1(n14537), .A2(n13102), .ZN(n13105) );
  NAND2_X1 U15474 ( .A1(n14803), .A2(n13103), .ZN(n13104) );
  NAND2_X1 U15475 ( .A1(n13105), .A2(n13104), .ZN(n13106) );
  XNOR2_X1 U15476 ( .A(n13106), .B(n13115), .ZN(n13107) );
  XOR2_X1 U15477 ( .A(n13108), .B(n13107), .Z(n14533) );
  INV_X1 U15478 ( .A(n13107), .ZN(n13110) );
  INV_X1 U15479 ( .A(n13108), .ZN(n13109) );
  OAI22_X1 U15480 ( .A1(n14817), .A2(n13111), .B1(n13113), .B2(n6681), .ZN(
        n13118) );
  OAI22_X1 U15481 ( .A1(n14817), .A2(n6681), .B1(n13113), .B2(n13112), .ZN(
        n13116) );
  XNOR2_X1 U15482 ( .A(n13116), .B(n13115), .ZN(n13117) );
  XOR2_X1 U15483 ( .A(n13118), .B(n13117), .Z(n13119) );
  AOI22_X1 U15484 ( .A1(n14587), .A2(n14803), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13121) );
  NAND2_X1 U15485 ( .A1(n14615), .A2(n14802), .ZN(n13120) );
  OAI211_X1 U15486 ( .C1(n15222), .C2(n14813), .A(n13121), .B(n13120), .ZN(
        n13122) );
  AOI21_X1 U15487 ( .B1(n15004), .B2(n15218), .A(n13122), .ZN(n13123) );
  INV_X1 U15488 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n13125) );
  OAI222_X1 U15489 ( .A1(n13374), .A2(n13125), .B1(n13377), .B2(n13124), .C1(
        n8213), .C2(P1_U3086), .ZN(P1_U3335) );
  INV_X1 U15490 ( .A(n13126), .ZN(n13130) );
  AOI22_X1 U15491 ( .A1(n13127), .A2(n15702), .B1(n13869), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n13128) );
  OAI21_X1 U15492 ( .B1(n13300), .B2(n13913), .A(n13128), .ZN(n13129) );
  AOI21_X1 U15493 ( .B1(n13130), .B2(n13733), .A(n13129), .ZN(n13131) );
  OAI21_X1 U15494 ( .B1(n13132), .B2(n13921), .A(n13131), .ZN(P3_U3206) );
  INV_X1 U15495 ( .A(n13134), .ZN(n13135) );
  NAND2_X1 U15496 ( .A1(n13375), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13137) );
  NAND2_X1 U15497 ( .A1(n13139), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13142) );
  NAND2_X1 U15498 ( .A1(n13140), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13141) );
  NAND2_X1 U15499 ( .A1(n13142), .A2(n13141), .ZN(n13147) );
  OAI21_X1 U15500 ( .B1(n13148), .B2(n13147), .A(n13142), .ZN(n13144) );
  XNOR2_X1 U15501 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n13143) );
  XNOR2_X1 U15502 ( .A(n13144), .B(n13143), .ZN(n14038) );
  NAND2_X1 U15503 ( .A1(n14038), .A2(n13149), .ZN(n13146) );
  OR2_X1 U15504 ( .A1(n13150), .A2(n14044), .ZN(n13145) );
  OR2_X1 U15505 ( .A1(n13159), .A2(n13684), .ZN(n13155) );
  XNOR2_X1 U15506 ( .A(n13148), .B(n13147), .ZN(n13378) );
  NAND2_X1 U15507 ( .A1(n13378), .A2(n13149), .ZN(n13152) );
  OR2_X1 U15508 ( .A1(n13150), .A2(n13381), .ZN(n13151) );
  NAND2_X1 U15509 ( .A1(n13924), .A2(n13153), .ZN(n13154) );
  NAND2_X1 U15510 ( .A1(n13155), .A2(n13154), .ZN(n13341) );
  OAI21_X1 U15511 ( .B1(n13989), .B2(n13157), .A(n13306), .ZN(n13156) );
  NOR2_X1 U15512 ( .A1(n13341), .A2(n13156), .ZN(n13163) );
  NOR2_X1 U15513 ( .A1(n13986), .A2(n13157), .ZN(n13342) );
  INV_X1 U15514 ( .A(n13342), .ZN(n13161) );
  NAND2_X1 U15515 ( .A1(n13340), .A2(n13159), .ZN(n13160) );
  XNOR2_X1 U15516 ( .A(n13165), .B(n13679), .ZN(n13353) );
  INV_X1 U15517 ( .A(n13166), .ZN(n13352) );
  NAND2_X1 U15518 ( .A1(n13168), .A2(n13173), .ZN(n13167) );
  NAND2_X1 U15519 ( .A1(n13167), .A2(n13267), .ZN(n13170) );
  NAND3_X1 U15520 ( .A1(n13168), .A2(n13176), .A3(n13356), .ZN(n13169) );
  NAND2_X1 U15521 ( .A1(n13170), .A2(n13169), .ZN(n13171) );
  OAI21_X1 U15522 ( .B1(n13173), .B2(n13172), .A(n13171), .ZN(n13175) );
  NOR2_X1 U15523 ( .A1(n13176), .A2(n13305), .ZN(n13177) );
  NOR2_X1 U15524 ( .A1(n13178), .A2(n13177), .ZN(n13181) );
  AOI21_X1 U15525 ( .B1(n13189), .B2(n13179), .A(n13305), .ZN(n13180) );
  AOI21_X1 U15526 ( .B1(n13182), .B2(n13181), .A(n13180), .ZN(n13187) );
  INV_X1 U15527 ( .A(n13184), .ZN(n13186) );
  NAND2_X1 U15528 ( .A1(n9273), .A2(n15697), .ZN(n13183) );
  AND2_X1 U15529 ( .A1(n13184), .A2(n13183), .ZN(n13185) );
  OAI211_X1 U15530 ( .C1(n13189), .C2(n13267), .A(n13188), .B(n9280), .ZN(
        n13190) );
  NAND2_X1 U15531 ( .A1(n13190), .A2(n13316), .ZN(n13199) );
  NAND2_X1 U15532 ( .A1(n13202), .A2(n13191), .ZN(n13194) );
  NAND2_X1 U15533 ( .A1(n13194), .A2(n13305), .ZN(n13198) );
  INV_X1 U15534 ( .A(n13192), .ZN(n13196) );
  NOR2_X1 U15535 ( .A1(n13194), .A2(n13193), .ZN(n13195) );
  MUX2_X1 U15536 ( .A(n13196), .B(n13195), .S(n13305), .Z(n13197) );
  AOI21_X1 U15537 ( .B1(n13199), .B2(n13198), .A(n13197), .ZN(n13205) );
  AOI21_X1 U15538 ( .B1(n13200), .B2(n13201), .A(n13305), .ZN(n13204) );
  MUX2_X1 U15539 ( .A(n13202), .B(n13201), .S(n13305), .Z(n13203) );
  OAI211_X1 U15540 ( .C1(n13205), .C2(n13204), .A(n13317), .B(n13203), .ZN(
        n13209) );
  MUX2_X1 U15541 ( .A(n13207), .B(n13206), .S(n13305), .Z(n13208) );
  NAND3_X1 U15542 ( .A1(n13209), .A2(n13326), .A3(n13208), .ZN(n13215) );
  NAND2_X1 U15543 ( .A1(n13533), .A2(n13210), .ZN(n13211) );
  MUX2_X1 U15544 ( .A(n13212), .B(n13211), .S(n13305), .Z(n13213) );
  NAND3_X1 U15545 ( .A1(n13215), .A2(n13214), .A3(n13213), .ZN(n13219) );
  MUX2_X1 U15546 ( .A(n13217), .B(n13216), .S(n13305), .Z(n13218) );
  NAND2_X1 U15547 ( .A1(n13219), .A2(n13218), .ZN(n13225) );
  INV_X1 U15548 ( .A(n13220), .ZN(n13321) );
  MUX2_X1 U15549 ( .A(n13222), .B(n13221), .S(n13305), .Z(n13223) );
  NAND2_X1 U15550 ( .A1(n13223), .A2(n13327), .ZN(n13224) );
  AOI21_X1 U15551 ( .B1(n13225), .B2(n13321), .A(n13224), .ZN(n13235) );
  NAND2_X1 U15552 ( .A1(n13232), .A2(n13226), .ZN(n13229) );
  NAND2_X1 U15553 ( .A1(n13231), .A2(n13227), .ZN(n13228) );
  MUX2_X1 U15554 ( .A(n13229), .B(n13228), .S(n13267), .Z(n13234) );
  INV_X1 U15555 ( .A(n13230), .ZN(n13244) );
  OR2_X1 U15556 ( .A1(n13236), .A2(n13244), .ZN(n13891) );
  INV_X1 U15557 ( .A(n13891), .ZN(n13893) );
  MUX2_X1 U15558 ( .A(n13232), .B(n13231), .S(n13305), .Z(n13233) );
  AND2_X1 U15559 ( .A1(n13236), .A2(n13267), .ZN(n13237) );
  NOR2_X1 U15560 ( .A1(n13883), .A2(n13237), .ZN(n13238) );
  NAND2_X1 U15561 ( .A1(n14032), .A2(n13528), .ZN(n13239) );
  INV_X1 U15562 ( .A(n13865), .ZN(n13861) );
  AOI21_X1 U15563 ( .B1(n13245), .B2(n13239), .A(n13861), .ZN(n13242) );
  NAND2_X1 U15564 ( .A1(n13252), .A2(n13240), .ZN(n13241) );
  NAND2_X1 U15565 ( .A1(n13896), .A2(n13305), .ZN(n13243) );
  OAI22_X1 U15566 ( .A1(n13245), .A2(n13244), .B1(n14032), .B2(n13243), .ZN(
        n13246) );
  NAND2_X1 U15567 ( .A1(n13246), .A2(n13865), .ZN(n13248) );
  INV_X1 U15568 ( .A(n13251), .ZN(n13247) );
  AOI21_X1 U15569 ( .B1(n13249), .B2(n13248), .A(n13247), .ZN(n13254) );
  AOI21_X1 U15570 ( .B1(n13251), .B2(n13250), .A(n13267), .ZN(n13253) );
  OAI22_X1 U15571 ( .A1(n13254), .A2(n13253), .B1(n13267), .B2(n13252), .ZN(
        n13261) );
  INV_X1 U15572 ( .A(n13255), .ZN(n13260) );
  INV_X1 U15573 ( .A(n13262), .ZN(n13259) );
  AND2_X1 U15574 ( .A1(n13256), .A2(n13305), .ZN(n13257) );
  OAI211_X1 U15575 ( .C1(n13259), .C2(n13258), .A(n13268), .B(n13257), .ZN(
        n13264) );
  AOI22_X1 U15576 ( .A1(n13261), .A2(n13847), .B1(n13260), .B2(n13264), .ZN(
        n13266) );
  NAND3_X1 U15577 ( .A1(n13269), .A2(n13267), .A3(n13262), .ZN(n13263) );
  NAND2_X1 U15578 ( .A1(n13264), .A2(n13263), .ZN(n13265) );
  OAI21_X1 U15579 ( .B1(n13266), .B2(n13831), .A(n13265), .ZN(n13271) );
  INV_X1 U15580 ( .A(n13798), .ZN(n13802) );
  MUX2_X1 U15581 ( .A(n13269), .B(n13268), .S(n13267), .Z(n13270) );
  MUX2_X1 U15582 ( .A(n13273), .B(n13272), .S(n13305), .Z(n13274) );
  MUX2_X1 U15583 ( .A(n13737), .B(n13736), .S(n13305), .Z(n13275) );
  NAND3_X1 U15584 ( .A1(n13276), .A2(n13773), .A3(n13275), .ZN(n13278) );
  MUX2_X1 U15585 ( .A(n13739), .B(n13757), .S(n13305), .Z(n13277) );
  NAND3_X1 U15586 ( .A1(n13278), .A2(n13760), .A3(n13277), .ZN(n13280) );
  NAND3_X1 U15587 ( .A1(n13766), .A2(n13776), .A3(n13305), .ZN(n13279) );
  AOI21_X1 U15588 ( .B1(n13280), .B2(n13279), .A(n13746), .ZN(n13286) );
  INV_X1 U15589 ( .A(n13746), .ZN(n13284) );
  XNOR2_X1 U15590 ( .A(n13281), .B(n13305), .ZN(n13282) );
  AOI21_X1 U15591 ( .B1(n13284), .B2(n13283), .A(n13282), .ZN(n13285) );
  NOR2_X1 U15592 ( .A1(n13335), .A2(n13287), .ZN(n13289) );
  AOI21_X1 U15593 ( .B1(n13294), .B2(n13289), .A(n13288), .ZN(n13296) );
  INV_X1 U15594 ( .A(n13290), .ZN(n13291) );
  NOR2_X1 U15595 ( .A1(n13335), .A2(n13291), .ZN(n13293) );
  AOI21_X1 U15596 ( .B1(n13294), .B2(n13293), .A(n13292), .ZN(n13295) );
  NAND2_X1 U15597 ( .A1(n13300), .A2(n13299), .ZN(n13301) );
  AOI21_X1 U15598 ( .B1(n13308), .B2(n13301), .A(n9317), .ZN(n13302) );
  NAND2_X1 U15599 ( .A1(n13700), .A2(n13305), .ZN(n13307) );
  OAI21_X1 U15600 ( .B1(n13308), .B2(n13307), .A(n13306), .ZN(n13311) );
  INV_X1 U15601 ( .A(n13340), .ZN(n13309) );
  OAI211_X1 U15602 ( .C1(n13312), .C2(n13311), .A(n13310), .B(n13309), .ZN(
        n13314) );
  INV_X1 U15603 ( .A(n13341), .ZN(n13313) );
  NAND4_X1 U15604 ( .A1(n13318), .A2(n13317), .A3(n9280), .A4(n13316), .ZN(
        n13325) );
  NAND4_X1 U15605 ( .A1(n13322), .A2(n13321), .A3(n13320), .A4(n13319), .ZN(
        n13324) );
  NOR3_X1 U15606 ( .A1(n13325), .A2(n13324), .A3(n13323), .ZN(n13328) );
  NAND4_X1 U15607 ( .A1(n13328), .A2(n15687), .A3(n13327), .A4(n13326), .ZN(
        n13329) );
  NOR4_X1 U15608 ( .A1(n13861), .A2(n13329), .A3(n13906), .A4(n13891), .ZN(
        n13330) );
  NAND4_X1 U15609 ( .A1(n9106), .A2(n13857), .A3(n13330), .A4(n9038), .ZN(
        n13331) );
  NOR4_X1 U15610 ( .A1(n13798), .A2(n13332), .A3(n13815), .A4(n13331), .ZN(
        n13333) );
  NAND4_X1 U15611 ( .A1(n13760), .A2(n13786), .A3(n13773), .A4(n13333), .ZN(
        n13334) );
  NOR4_X1 U15612 ( .A1(n13335), .A2(n13746), .A3(n13721), .A4(n13334), .ZN(
        n13337) );
  NAND4_X1 U15613 ( .A1(n13338), .A2(n13700), .A3(n13337), .A4(n13336), .ZN(
        n13339) );
  XNOR2_X1 U15614 ( .A(n13343), .B(n13666), .ZN(n13344) );
  OAI22_X1 U15615 ( .A1(n13348), .A2(n15698), .B1(n13345), .B2(n13344), .ZN(
        n13346) );
  NAND2_X1 U15616 ( .A1(n13348), .A2(n13347), .ZN(n13349) );
  NOR3_X1 U15617 ( .A1(n13355), .A2(n13590), .A3(n13354), .ZN(n13358) );
  OAI21_X1 U15618 ( .B1(n13359), .B2(n13356), .A(P3_B_REG_SCAN_IN), .ZN(n13357) );
  OAI22_X1 U15619 ( .A1(n13360), .A2(n13359), .B1(n13358), .B2(n13357), .ZN(
        P3_U3296) );
  INV_X1 U15620 ( .A(n13361), .ZN(n13362) );
  NAND2_X1 U15621 ( .A1(n13363), .A2(n13362), .ZN(n13366) );
  XOR2_X1 U15622 ( .A(n13364), .B(n13700), .Z(n13365) );
  XNOR2_X1 U15623 ( .A(n13366), .B(n13365), .ZN(n13372) );
  OAI22_X1 U15624 ( .A1(n13703), .A2(n13495), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13367), .ZN(n13370) );
  INV_X1 U15625 ( .A(n13708), .ZN(n13368) );
  OAI22_X1 U15626 ( .A1(n13702), .A2(n13514), .B1(n13368), .B2(n13518), .ZN(
        n13369) );
  AOI211_X1 U15627 ( .C1(n13707), .C2(n13520), .A(n13370), .B(n13369), .ZN(
        n13371) );
  OAI21_X1 U15628 ( .B1(n13372), .B2(n13523), .A(n13371), .ZN(P3_U3160) );
  INV_X1 U15629 ( .A(n13373), .ZN(n14530) );
  OAI222_X1 U15630 ( .A1(n13377), .A2(n14530), .B1(P1_U3086), .B2(n13376), 
        .C1(n13375), .C2(n13374), .ZN(P1_U3326) );
  INV_X1 U15631 ( .A(n13378), .ZN(n13380) );
  OAI222_X1 U15632 ( .A1(n13382), .A2(n13381), .B1(n12850), .B2(n13380), .C1(
        n13379), .C2(P3_U3151), .ZN(P3_U3265) );
  OAI211_X1 U15633 ( .C1(n13385), .C2(n13384), .A(n13383), .B(n13492), .ZN(
        n13391) );
  INV_X1 U15634 ( .A(n13885), .ZN(n13389) );
  NOR2_X1 U15635 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13386), .ZN(n13575) );
  AOI21_X1 U15636 ( .B1(n13482), .B2(n13878), .A(n13575), .ZN(n13387) );
  OAI21_X1 U15637 ( .B1(n7491), .B2(n13495), .A(n13387), .ZN(n13388) );
  AOI21_X1 U15638 ( .B1(n13498), .B2(n13389), .A(n13388), .ZN(n13390) );
  OAI211_X1 U15639 ( .C1(n13501), .C2(n14032), .A(n13391), .B(n13390), .ZN(
        P3_U3155) );
  INV_X1 U15640 ( .A(n13392), .ZN(n13458) );
  AOI21_X1 U15641 ( .B1(n6684), .B2(n13393), .A(n13458), .ZN(n13398) );
  AOI22_X1 U15642 ( .A1(n9301), .A2(n13516), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13395) );
  NAND2_X1 U15643 ( .A1(n13498), .A2(n13767), .ZN(n13394) );
  OAI211_X1 U15644 ( .C1(n13723), .C2(n13514), .A(n13395), .B(n13394), .ZN(
        n13396) );
  AOI21_X1 U15645 ( .B1(n13766), .B2(n13520), .A(n13396), .ZN(n13397) );
  OAI21_X1 U15646 ( .B1(n13398), .B2(n13523), .A(n13397), .ZN(P3_U3156) );
  XNOR2_X1 U15647 ( .A(n13399), .B(n13466), .ZN(n13404) );
  NAND2_X1 U15648 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13678)
         );
  OAI21_X1 U15649 ( .B1(n13789), .B2(n13514), .A(n13678), .ZN(n13400) );
  AOI21_X1 U15650 ( .B1(n13516), .B2(n13842), .A(n13400), .ZN(n13401) );
  OAI21_X1 U15651 ( .B1(n13818), .B2(n13518), .A(n13401), .ZN(n13402) );
  AOI21_X1 U15652 ( .B1(n13817), .B2(n13520), .A(n13402), .ZN(n13403) );
  OAI21_X1 U15653 ( .B1(n13404), .B2(n13523), .A(n13403), .ZN(P3_U3159) );
  NAND2_X1 U15654 ( .A1(n13406), .A2(n13405), .ZN(n13409) );
  INV_X1 U15655 ( .A(n13407), .ZN(n13408) );
  AOI21_X1 U15656 ( .B1(n13410), .B2(n13409), .A(n13408), .ZN(n13416) );
  NAND2_X1 U15657 ( .A1(n13498), .A2(n13790), .ZN(n13412) );
  AOI22_X1 U15658 ( .A1(n13812), .A2(n13516), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13411) );
  OAI211_X1 U15659 ( .C1(n13788), .C2(n13514), .A(n13412), .B(n13411), .ZN(
        n13413) );
  AOI21_X1 U15660 ( .B1(n13414), .B2(n13520), .A(n13413), .ZN(n13415) );
  OAI21_X1 U15661 ( .B1(n13416), .B2(n13523), .A(n13415), .ZN(P3_U3163) );
  OAI21_X1 U15662 ( .B1(n13419), .B2(n13418), .A(n13417), .ZN(n13420) );
  NAND2_X1 U15663 ( .A1(n13420), .A2(n13492), .ZN(n13426) );
  AOI21_X1 U15664 ( .B1(n13482), .B2(n13879), .A(n13421), .ZN(n13423) );
  NAND2_X1 U15665 ( .A1(n13516), .A2(n13529), .ZN(n13422) );
  OAI211_X1 U15666 ( .C1(n13518), .C2(n13915), .A(n13423), .B(n13422), .ZN(
        n13424) );
  INV_X1 U15667 ( .A(n13424), .ZN(n13425) );
  OAI211_X1 U15668 ( .C1(n15146), .C2(n13501), .A(n13426), .B(n13425), .ZN(
        P3_U3164) );
  INV_X1 U15669 ( .A(n13428), .ZN(n13459) );
  INV_X1 U15670 ( .A(n13429), .ZN(n13431) );
  NOR3_X1 U15671 ( .A1(n13459), .A2(n13431), .A3(n13430), .ZN(n13434) );
  INV_X1 U15672 ( .A(n13432), .ZN(n13433) );
  OAI21_X1 U15673 ( .B1(n13434), .B2(n13433), .A(n13492), .ZN(n13438) );
  AOI22_X1 U15674 ( .A1(n13763), .A2(n13516), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13435) );
  OAI21_X1 U15675 ( .B1(n13724), .B2(n13514), .A(n13435), .ZN(n13436) );
  AOI21_X1 U15676 ( .B1(n13730), .B2(n13498), .A(n13436), .ZN(n13437) );
  OAI211_X1 U15677 ( .C1(n13997), .C2(n13501), .A(n13438), .B(n13437), .ZN(
        P3_U3165) );
  XNOR2_X1 U15678 ( .A(n13440), .B(n13439), .ZN(n13446) );
  NOR2_X1 U15679 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13441), .ZN(n13622) );
  NOR2_X1 U15680 ( .A1(n13828), .A2(n13514), .ZN(n13442) );
  AOI211_X1 U15681 ( .C1(n13516), .C2(n13878), .A(n13622), .B(n13442), .ZN(
        n13443) );
  OAI21_X1 U15682 ( .B1(n6707), .B2(n13518), .A(n13443), .ZN(n13444) );
  AOI21_X1 U15683 ( .B1(n13971), .B2(n13520), .A(n13444), .ZN(n13445) );
  OAI21_X1 U15684 ( .B1(n13446), .B2(n13523), .A(n13445), .ZN(P3_U3166) );
  XNOR2_X1 U15685 ( .A(n13447), .B(n13448), .ZN(n13454) );
  NAND2_X1 U15686 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n15131)
         );
  OAI21_X1 U15687 ( .B1(n13449), .B2(n13514), .A(n15131), .ZN(n13450) );
  AOI21_X1 U15688 ( .B1(n13516), .B2(n13843), .A(n13450), .ZN(n13451) );
  OAI21_X1 U15689 ( .B1(n13845), .B2(n13518), .A(n13451), .ZN(n13452) );
  AOI21_X1 U15690 ( .B1(n13967), .B2(n13520), .A(n13452), .ZN(n13453) );
  OAI21_X1 U15691 ( .B1(n13454), .B2(n13523), .A(n13453), .ZN(P3_U3168) );
  INV_X1 U15692 ( .A(n13937), .ZN(n13465) );
  INV_X1 U15693 ( .A(n13455), .ZN(n13457) );
  NOR3_X1 U15694 ( .A1(n13458), .A2(n13457), .A3(n13456), .ZN(n13460) );
  OAI21_X1 U15695 ( .B1(n13460), .B2(n13459), .A(n13492), .ZN(n13464) );
  AOI22_X1 U15696 ( .A1(n6684), .A2(n13516), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13461) );
  OAI21_X1 U15697 ( .B1(n13750), .B2(n13514), .A(n13461), .ZN(n13462) );
  AOI21_X1 U15698 ( .B1(n13751), .B2(n13498), .A(n13462), .ZN(n13463) );
  OAI211_X1 U15699 ( .C1(n13465), .C2(n13501), .A(n13464), .B(n13463), .ZN(
        P3_U3169) );
  NAND2_X1 U15700 ( .A1(n13399), .A2(n13466), .ZN(n13468) );
  NAND2_X1 U15701 ( .A1(n13468), .A2(n13467), .ZN(n13470) );
  XNOR2_X1 U15702 ( .A(n13470), .B(n13469), .ZN(n13476) );
  NOR2_X1 U15703 ( .A1(n13827), .A2(n13495), .ZN(n13473) );
  OAI22_X1 U15704 ( .A1(n13801), .A2(n13514), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13471), .ZN(n13472) );
  AOI211_X1 U15705 ( .C1(n13805), .C2(n13498), .A(n13473), .B(n13472), .ZN(
        n13475) );
  NAND2_X1 U15706 ( .A1(n13804), .A2(n13520), .ZN(n13474) );
  OAI211_X1 U15707 ( .C1(n13476), .C2(n13523), .A(n13475), .B(n13474), .ZN(
        P3_U3173) );
  INV_X1 U15708 ( .A(n13477), .ZN(n13479) );
  NAND2_X1 U15709 ( .A1(n13479), .A2(n13478), .ZN(n13480) );
  XNOR2_X1 U15710 ( .A(n13481), .B(n13480), .ZN(n13488) );
  INV_X1 U15711 ( .A(n15142), .ZN(n13902) );
  NOR2_X1 U15712 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9013), .ZN(n13548) );
  AOI21_X1 U15713 ( .B1(n13528), .B2(n13482), .A(n13548), .ZN(n13485) );
  NAND2_X1 U15714 ( .A1(n13483), .A2(n13516), .ZN(n13484) );
  OAI211_X1 U15715 ( .C1(n13518), .C2(n13898), .A(n13485), .B(n13484), .ZN(
        n13486) );
  AOI21_X1 U15716 ( .B1(n13902), .B2(n13520), .A(n13486), .ZN(n13487) );
  OAI21_X1 U15717 ( .B1(n13488), .B2(n13523), .A(n13487), .ZN(P3_U3174) );
  AND2_X1 U15718 ( .A1(n12937), .A2(n13489), .ZN(n13491) );
  OAI21_X1 U15719 ( .B1(n13491), .B2(n13788), .A(n13490), .ZN(n13493) );
  NAND2_X1 U15720 ( .A1(n13493), .A2(n13492), .ZN(n13500) );
  OAI22_X1 U15721 ( .A1(n13801), .A2(n13495), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13494), .ZN(n13497) );
  NOR2_X1 U15722 ( .A1(n13776), .A2(n13514), .ZN(n13496) );
  AOI211_X1 U15723 ( .C1(n13777), .C2(n13498), .A(n13497), .B(n13496), .ZN(
        n13499) );
  OAI211_X1 U15724 ( .C1(n14006), .C2(n13501), .A(n13500), .B(n13499), .ZN(
        P3_U3175) );
  XNOR2_X1 U15725 ( .A(n13502), .B(n13503), .ZN(n13508) );
  NAND2_X1 U15726 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13636)
         );
  OAI21_X1 U15727 ( .B1(n13827), .B2(n13514), .A(n13636), .ZN(n13504) );
  AOI21_X1 U15728 ( .B1(n13516), .B2(n13852), .A(n13504), .ZN(n13505) );
  OAI21_X1 U15729 ( .B1(n13829), .B2(n13518), .A(n13505), .ZN(n13506) );
  AOI21_X1 U15730 ( .B1(n13960), .B2(n13520), .A(n13506), .ZN(n13507) );
  OAI21_X1 U15731 ( .B1(n13508), .B2(n13523), .A(n13507), .ZN(P3_U3178) );
  XNOR2_X1 U15732 ( .A(n13511), .B(n13510), .ZN(n13512) );
  XNOR2_X1 U15733 ( .A(n13509), .B(n13512), .ZN(n13524) );
  NOR2_X1 U15734 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13513), .ZN(n13588) );
  NOR2_X1 U15735 ( .A1(n13864), .A2(n13514), .ZN(n13515) );
  AOI211_X1 U15736 ( .C1(n13516), .C2(n13528), .A(n13588), .B(n13515), .ZN(
        n13517) );
  OAI21_X1 U15737 ( .B1(n13867), .B2(n13518), .A(n13517), .ZN(n13519) );
  AOI21_X1 U15738 ( .B1(n13521), .B2(n13520), .A(n13519), .ZN(n13522) );
  OAI21_X1 U15739 ( .B1(n13524), .B2(n13523), .A(n13522), .ZN(P3_U3181) );
  MUX2_X1 U15740 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n13525), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U15741 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n13526), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U15742 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n13527), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U15743 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n13763), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U15744 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n13843), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U15745 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n13528), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U15746 ( .A(n13529), .B(P3_DATAO_REG_11__SCAN_IN), .S(n13532), .Z(
        P3_U3502) );
  MUX2_X1 U15747 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n13530), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U15748 ( .A(n13531), .B(P3_DATAO_REG_9__SCAN_IN), .S(n13532), .Z(
        P3_U3500) );
  MUX2_X1 U15749 ( .A(n13533), .B(P3_DATAO_REG_8__SCAN_IN), .S(n13532), .Z(
        P3_U3499) );
  MUX2_X1 U15750 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n13534), .S(n6678), .Z(
        P3_U3497) );
  MUX2_X1 U15751 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n13535), .S(n6678), .Z(
        P3_U3492) );
  MUX2_X1 U15752 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n13536), .S(n6678), .Z(
        P3_U3491) );
  INV_X1 U15753 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n13899) );
  INV_X1 U15754 ( .A(n13560), .ZN(n13566) );
  XNOR2_X1 U15755 ( .A(n13555), .B(n13566), .ZN(n13538) );
  AOI21_X1 U15756 ( .B1(n13899), .B2(n13538), .A(n13556), .ZN(n13554) );
  AOI21_X1 U15757 ( .B1(n13541), .B2(n13540), .A(n13539), .ZN(n13543) );
  MUX2_X1 U15758 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n13629), .Z(n13565) );
  XNOR2_X1 U15759 ( .A(n13565), .B(n13566), .ZN(n13542) );
  NAND2_X1 U15760 ( .A1(n13543), .A2(n13542), .ZN(n13572) );
  OAI21_X1 U15761 ( .B1(n13543), .B2(n13542), .A(n13572), .ZN(n13552) );
  OAI21_X1 U15762 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n13546), .A(n13561), 
        .ZN(n13547) );
  NAND2_X1 U15763 ( .A1(n13547), .A2(n15677), .ZN(n13550) );
  AOI21_X1 U15764 ( .B1(n15674), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n13548), 
        .ZN(n13549) );
  OAI211_X1 U15765 ( .C1(n15671), .C2(n13560), .A(n13550), .B(n13549), .ZN(
        n13551) );
  AOI21_X1 U15766 ( .B1(n13552), .B2(n15666), .A(n13551), .ZN(n13553) );
  OAI21_X1 U15767 ( .B1(n13554), .B2(n15681), .A(n13553), .ZN(P3_U3195) );
  NOR2_X1 U15768 ( .A1(n13566), .A2(n13555), .ZN(n13557) );
  NAND2_X1 U15769 ( .A1(n13583), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n13591) );
  OAI21_X1 U15770 ( .B1(P3_REG2_REG_14__SCAN_IN), .B2(n13583), .A(n13591), 
        .ZN(n13568) );
  AOI21_X1 U15771 ( .B1(n13558), .B2(n13568), .A(n13582), .ZN(n13581) );
  NAND2_X1 U15772 ( .A1(n13560), .A2(n13559), .ZN(n13562) );
  NAND2_X1 U15773 ( .A1(n13562), .A2(n13561), .ZN(n13564) );
  NAND2_X1 U15774 ( .A1(n13583), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n13592) );
  OR2_X1 U15775 ( .A1(n13583), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n13563) );
  AND2_X1 U15776 ( .A1(n13592), .A2(n13563), .ZN(n13570) );
  OAI21_X1 U15777 ( .B1(n13564), .B2(n13570), .A(n13586), .ZN(n13579) );
  INV_X1 U15778 ( .A(n13565), .ZN(n13567) );
  NAND2_X1 U15779 ( .A1(n13567), .A2(n13566), .ZN(n13571) );
  AND2_X1 U15780 ( .A1(n13572), .A2(n13571), .ZN(n13574) );
  INV_X1 U15781 ( .A(n13568), .ZN(n13569) );
  MUX2_X1 U15782 ( .A(n13570), .B(n13569), .S(n13590), .Z(n13573) );
  NAND3_X1 U15783 ( .A1(n13572), .A2(n13573), .A3(n13571), .ZN(n13594) );
  OAI211_X1 U15784 ( .C1(n13574), .C2(n13573), .A(n15666), .B(n13594), .ZN(
        n13577) );
  AOI21_X1 U15785 ( .B1(n15674), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n13575), 
        .ZN(n13576) );
  OAI211_X1 U15786 ( .C1(n15671), .C2(n13583), .A(n13577), .B(n13576), .ZN(
        n13578) );
  AOI21_X1 U15787 ( .B1(n15677), .B2(n13579), .A(n13578), .ZN(n13580) );
  OAI21_X1 U15788 ( .B1(n13581), .B2(n15681), .A(n13580), .ZN(P3_U3196) );
  AOI21_X1 U15789 ( .B1(n13585), .B2(n13584), .A(n13604), .ZN(n13602) );
  XNOR2_X1 U15790 ( .A(n13610), .B(n13615), .ZN(n13587) );
  NAND2_X1 U15791 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n13587), .ZN(n13617) );
  OAI21_X1 U15792 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n13587), .A(n13617), 
        .ZN(n13600) );
  AOI21_X1 U15793 ( .B1(n15674), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n13588), 
        .ZN(n13589) );
  OAI21_X1 U15794 ( .B1(n15671), .B2(n13616), .A(n13589), .ZN(n13599) );
  MUX2_X1 U15795 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n13629), .Z(n13596) );
  MUX2_X1 U15796 ( .A(n13592), .B(n13591), .S(n13590), .Z(n13593) );
  NAND2_X1 U15797 ( .A1(n13594), .A2(n13593), .ZN(n13608) );
  XNOR2_X1 U15798 ( .A(n13608), .B(n13616), .ZN(n13595) );
  AOI21_X1 U15799 ( .B1(n13596), .B2(n13595), .A(n13609), .ZN(n13597) );
  NOR2_X1 U15800 ( .A1(n13597), .A2(n15595), .ZN(n13598) );
  AOI211_X1 U15801 ( .C1(n15677), .C2(n13600), .A(n13599), .B(n13598), .ZN(
        n13601) );
  OAI21_X1 U15802 ( .B1(n13602), .B2(n15681), .A(n13601), .ZN(P3_U3197) );
  NOR2_X1 U15803 ( .A1(n13610), .A2(n13603), .ZN(n13605) );
  AOI22_X1 U15804 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n13640), .B1(n13648), 
        .B2(n13854), .ZN(n13606) );
  AOI21_X1 U15805 ( .B1(n13607), .B2(n13606), .A(n6738), .ZN(n13628) );
  INV_X1 U15806 ( .A(n13608), .ZN(n13611) );
  AOI21_X1 U15807 ( .B1(n13611), .B2(n13610), .A(n13609), .ZN(n13632) );
  MUX2_X1 U15808 ( .A(n13854), .B(n13639), .S(n13667), .Z(n13612) );
  NOR2_X1 U15809 ( .A1(n13612), .A2(n13640), .ZN(n13631) );
  INV_X1 U15810 ( .A(n13631), .ZN(n13613) );
  NAND2_X1 U15811 ( .A1(n13612), .A2(n13640), .ZN(n13630) );
  NAND2_X1 U15812 ( .A1(n13613), .A2(n13630), .ZN(n13614) );
  XNOR2_X1 U15813 ( .A(n13632), .B(n13614), .ZN(n13626) );
  AOI22_X1 U15814 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n13648), .B1(n13640), 
        .B2(n13639), .ZN(n13620) );
  NAND2_X1 U15815 ( .A1(n13616), .A2(n13615), .ZN(n13618) );
  NAND2_X1 U15816 ( .A1(n13620), .A2(n13619), .ZN(n13638) );
  OAI21_X1 U15817 ( .B1(n13620), .B2(n13619), .A(n13638), .ZN(n13621) );
  NAND2_X1 U15818 ( .A1(n13621), .A2(n15677), .ZN(n13624) );
  AOI21_X1 U15819 ( .B1(n15674), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n13622), 
        .ZN(n13623) );
  OAI211_X1 U15820 ( .C1(n15671), .C2(n13648), .A(n13624), .B(n13623), .ZN(
        n13625) );
  AOI21_X1 U15821 ( .B1(n13626), .B2(n15666), .A(n13625), .ZN(n13627) );
  OAI21_X1 U15822 ( .B1(n13628), .B2(n15681), .A(n13627), .ZN(P3_U3198) );
  MUX2_X1 U15823 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n13629), .Z(n13635) );
  MUX2_X1 U15824 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n13629), .Z(n13633) );
  OAI21_X1 U15825 ( .B1(n13632), .B2(n13631), .A(n13630), .ZN(n15135) );
  XNOR2_X1 U15826 ( .A(n13633), .B(n13649), .ZN(n15136) );
  NOR2_X1 U15827 ( .A1(n15135), .A2(n15136), .ZN(n15134) );
  XNOR2_X1 U15828 ( .A(n13665), .B(n13664), .ZN(n13634) );
  NOR2_X1 U15829 ( .A1(n13634), .A2(n13635), .ZN(n13663) );
  AOI21_X1 U15830 ( .B1(n13635), .B2(n13634), .A(n13663), .ZN(n13659) );
  INV_X1 U15831 ( .A(n15671), .ZN(n15600) );
  INV_X1 U15832 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n13637) );
  OAI21_X1 U15833 ( .B1(n15591), .B2(n13637), .A(n13636), .ZN(n13647) );
  NAND2_X1 U15834 ( .A1(n13641), .A2(n13649), .ZN(n13643) );
  NAND2_X1 U15835 ( .A1(P3_REG1_REG_17__SCAN_IN), .A2(n15129), .ZN(n15128) );
  INV_X1 U15836 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13965) );
  XNOR2_X1 U15837 ( .A(n13664), .B(n13965), .ZN(n13642) );
  INV_X1 U15838 ( .A(n13671), .ZN(n13645) );
  NAND3_X1 U15839 ( .A1(n13643), .A2(n15128), .A3(n13642), .ZN(n13644) );
  AOI21_X1 U15840 ( .B1(n13645), .B2(n13644), .A(n15583), .ZN(n13646) );
  AOI211_X1 U15841 ( .C1(n15600), .C2(n13664), .A(n13647), .B(n13646), .ZN(
        n13658) );
  OR2_X1 U15842 ( .A1(n13650), .A2(n15130), .ZN(n13653) );
  INV_X1 U15843 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13830) );
  OR2_X1 U15844 ( .A1(n13664), .A2(n13830), .ZN(n13660) );
  NAND2_X1 U15845 ( .A1(n13664), .A2(n13830), .ZN(n13651) );
  NAND2_X1 U15846 ( .A1(n13660), .A2(n13651), .ZN(n13652) );
  AND3_X1 U15847 ( .A1(n13654), .A2(n13653), .A3(n13652), .ZN(n13656) );
  OAI21_X1 U15848 ( .B1(n13661), .B2(n13656), .A(n13655), .ZN(n13657) );
  OAI211_X1 U15849 ( .C1(n13659), .C2(n15595), .A(n13658), .B(n13657), .ZN(
        P3_U3200) );
  XNOR2_X1 U15850 ( .A(n13666), .B(n13819), .ZN(n13668) );
  INV_X1 U15851 ( .A(n13668), .ZN(n13662) );
  AOI21_X1 U15852 ( .B1(n13665), .B2(n13664), .A(n13663), .ZN(n13670) );
  XNOR2_X1 U15853 ( .A(n13666), .B(n13958), .ZN(n13673) );
  MUX2_X1 U15854 ( .A(n13668), .B(n13673), .S(n13667), .Z(n13669) );
  XNOR2_X1 U15855 ( .A(n13670), .B(n13669), .ZN(n13681) );
  INV_X1 U15856 ( .A(n13673), .ZN(n13674) );
  XNOR2_X1 U15857 ( .A(n13675), .B(n13674), .ZN(n13676) );
  NAND2_X1 U15858 ( .A1(n15674), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n13677) );
  OAI211_X1 U15859 ( .C1(n15671), .C2(n13679), .A(n13678), .B(n13677), .ZN(
        n13680) );
  NAND2_X1 U15860 ( .A1(n13690), .A2(n15702), .ZN(n13685) );
  AOI21_X1 U15861 ( .B1(n13685), .B2(n13984), .A(n13869), .ZN(n13687) );
  AOI21_X1 U15862 ( .B1(n13869), .B2(P3_REG2_REG_31__SCAN_IN), .A(n13687), 
        .ZN(n13686) );
  OAI21_X1 U15863 ( .B1(n13986), .B2(n13913), .A(n13686), .ZN(P3_U3202) );
  AOI21_X1 U15864 ( .B1(n13869), .B2(P3_REG2_REG_30__SCAN_IN), .A(n13687), 
        .ZN(n13688) );
  OAI21_X1 U15865 ( .B1(n13989), .B2(n13913), .A(n13688), .ZN(P3_U3203) );
  INV_X1 U15866 ( .A(n13689), .ZN(n13694) );
  AOI22_X1 U15867 ( .A1(n13690), .A2(n15702), .B1(P3_REG2_REG_29__SCAN_IN), 
        .B2(n13921), .ZN(n13691) );
  OAI21_X1 U15868 ( .B1(n13692), .B2(n13913), .A(n13691), .ZN(n13693) );
  AOI21_X1 U15869 ( .B1(n13694), .B2(n13919), .A(n13693), .ZN(n13695) );
  OAI21_X1 U15870 ( .B1(n13696), .B2(n13921), .A(n13695), .ZN(P3_U3204) );
  NOR2_X1 U15871 ( .A1(n13698), .A2(n13697), .ZN(n13699) );
  AOI21_X1 U15872 ( .B1(n13701), .B2(n13700), .A(n15696), .ZN(n13706) );
  OAI22_X1 U15873 ( .A1(n13703), .A2(n15690), .B1(n13702), .B2(n15689), .ZN(
        n13704) );
  INV_X1 U15874 ( .A(n13928), .ZN(n13711) );
  INV_X1 U15875 ( .A(n13707), .ZN(n13993) );
  AOI22_X1 U15876 ( .A1(n13708), .A2(n15702), .B1(n13869), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n13709) );
  OAI21_X1 U15877 ( .B1(n13993), .B2(n13913), .A(n13709), .ZN(n13710) );
  AOI21_X1 U15878 ( .B1(n13711), .B2(n15703), .A(n13710), .ZN(n13712) );
  OAI21_X1 U15879 ( .B1(n13905), .B2(n13929), .A(n13712), .ZN(P3_U3205) );
  AOI22_X1 U15880 ( .A1(n13713), .A2(n15702), .B1(n13869), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n13714) );
  OAI21_X1 U15881 ( .B1(n13715), .B2(n13913), .A(n13714), .ZN(n13716) );
  AOI21_X1 U15882 ( .B1(n13717), .B2(n13733), .A(n13716), .ZN(n13718) );
  OAI21_X1 U15883 ( .B1(n6735), .B2(n13921), .A(n13718), .ZN(P3_U3207) );
  XNOR2_X1 U15884 ( .A(n13719), .B(n13721), .ZN(n13729) );
  OAI211_X1 U15885 ( .C1(n13722), .C2(n13721), .A(n13720), .B(n13874), .ZN(
        n13727) );
  OAI22_X1 U15886 ( .A1(n13724), .A2(n15689), .B1(n13723), .B2(n15690), .ZN(
        n13725) );
  INV_X1 U15887 ( .A(n13725), .ZN(n13726) );
  OAI211_X1 U15888 ( .C1(n13728), .C2(n13729), .A(n13727), .B(n13726), .ZN(
        n13932) );
  INV_X1 U15889 ( .A(n13932), .ZN(n13735) );
  INV_X1 U15890 ( .A(n13729), .ZN(n13933) );
  AOI22_X1 U15891 ( .A1(n13730), .A2(n15702), .B1(n13869), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n13731) );
  OAI21_X1 U15892 ( .B1(n13997), .B2(n13913), .A(n13731), .ZN(n13732) );
  AOI21_X1 U15893 ( .B1(n13933), .B2(n13733), .A(n13732), .ZN(n13734) );
  OAI21_X1 U15894 ( .B1(n13735), .B2(n13869), .A(n13734), .ZN(P3_U3208) );
  NAND2_X1 U15895 ( .A1(n13782), .A2(n13736), .ZN(n13738) );
  NAND2_X1 U15896 ( .A1(n13738), .A2(n13737), .ZN(n13772) );
  NAND2_X1 U15897 ( .A1(n13772), .A2(n13739), .ZN(n13758) );
  NAND2_X1 U15898 ( .A1(n13758), .A2(n13740), .ZN(n13742) );
  NOR2_X1 U15899 ( .A1(n13744), .A2(n13746), .ZN(n13743) );
  AOI21_X1 U15900 ( .B1(n13746), .B2(n13744), .A(n13743), .ZN(n13939) );
  OAI211_X1 U15901 ( .C1(n10168), .C2(n13746), .A(n13745), .B(n13874), .ZN(
        n13749) );
  NAND2_X1 U15902 ( .A1(n6684), .A2(n13880), .ZN(n13748) );
  OAI211_X1 U15903 ( .C1(n13750), .C2(n15689), .A(n13749), .B(n13748), .ZN(
        n13936) );
  NAND2_X1 U15904 ( .A1(n13936), .A2(n15703), .ZN(n13756) );
  INV_X1 U15905 ( .A(n13751), .ZN(n13753) );
  INV_X1 U15906 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n13752) );
  OAI22_X1 U15907 ( .A1(n13753), .A2(n13914), .B1(n15703), .B2(n13752), .ZN(
        n13754) );
  AOI21_X1 U15908 ( .B1(n13937), .B2(n13901), .A(n13754), .ZN(n13755) );
  OAI211_X1 U15909 ( .C1(n13905), .C2(n13939), .A(n13756), .B(n13755), .ZN(
        P3_U3209) );
  NAND2_X1 U15910 ( .A1(n13758), .A2(n13757), .ZN(n13759) );
  XOR2_X1 U15911 ( .A(n13760), .B(n13759), .Z(n13941) );
  INV_X1 U15912 ( .A(n13941), .ZN(n13771) );
  OAI211_X1 U15913 ( .C1(n13762), .C2(n9305), .A(n13761), .B(n13874), .ZN(
        n13765) );
  AOI22_X1 U15914 ( .A1(n13763), .A2(n13877), .B1(n13880), .B2(n9301), .ZN(
        n13764) );
  NAND2_X1 U15915 ( .A1(n13765), .A2(n13764), .ZN(n13940) );
  INV_X1 U15916 ( .A(n13766), .ZN(n14002) );
  AOI22_X1 U15917 ( .A1(n13869), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n13767), 
        .B2(n15702), .ZN(n13768) );
  OAI21_X1 U15918 ( .B1(n14002), .B2(n13913), .A(n13768), .ZN(n13769) );
  AOI21_X1 U15919 ( .B1(n13940), .B2(n15703), .A(n13769), .ZN(n13770) );
  OAI21_X1 U15920 ( .B1(n13905), .B2(n13771), .A(n13770), .ZN(P3_U3210) );
  XOR2_X1 U15921 ( .A(n13773), .B(n13772), .Z(n13945) );
  INV_X1 U15922 ( .A(n13945), .ZN(n13781) );
  XNOR2_X1 U15923 ( .A(n13774), .B(n13773), .ZN(n13775) );
  OAI222_X1 U15924 ( .A1(n15690), .A2(n13801), .B1(n15689), .B2(n13776), .C1(
        n15696), .C2(n13775), .ZN(n13944) );
  AOI22_X1 U15925 ( .A1(n13869), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n15702), 
        .B2(n13777), .ZN(n13778) );
  OAI21_X1 U15926 ( .B1(n14006), .B2(n13913), .A(n13778), .ZN(n13779) );
  AOI21_X1 U15927 ( .B1(n13944), .B2(n15703), .A(n13779), .ZN(n13780) );
  OAI21_X1 U15928 ( .B1(n13905), .B2(n13781), .A(n13780), .ZN(P3_U3211) );
  XOR2_X1 U15929 ( .A(n13786), .B(n13782), .Z(n13949) );
  INV_X1 U15930 ( .A(n13949), .ZN(n13794) );
  AOI21_X1 U15931 ( .B1(n13786), .B2(n13785), .A(n13784), .ZN(n13787) );
  OAI222_X1 U15932 ( .A1(n15690), .A2(n13789), .B1(n15689), .B2(n13788), .C1(
        n15696), .C2(n13787), .ZN(n13948) );
  AOI22_X1 U15933 ( .A1(n13869), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15702), 
        .B2(n13790), .ZN(n13791) );
  OAI21_X1 U15934 ( .B1(n14010), .B2(n13913), .A(n13791), .ZN(n13792) );
  AOI21_X1 U15935 ( .B1(n13948), .B2(n15703), .A(n13792), .ZN(n13793) );
  OAI21_X1 U15936 ( .B1(n13905), .B2(n13794), .A(n13793), .ZN(P3_U3212) );
  NOR2_X1 U15937 ( .A1(n13824), .A2(n13796), .ZN(n13811) );
  NAND2_X1 U15938 ( .A1(n13811), .A2(n13815), .ZN(n13810) );
  NAND2_X1 U15939 ( .A1(n13810), .A2(n13797), .ZN(n13799) );
  XNOR2_X1 U15940 ( .A(n13799), .B(n13798), .ZN(n13800) );
  OAI222_X1 U15941 ( .A1(n15689), .A2(n13801), .B1(n15690), .B2(n13827), .C1(
        n13800), .C2(n15696), .ZN(n13952) );
  INV_X1 U15942 ( .A(n13952), .ZN(n13809) );
  XNOR2_X1 U15943 ( .A(n13803), .B(n13802), .ZN(n13953) );
  INV_X1 U15944 ( .A(n13804), .ZN(n14014) );
  AOI22_X1 U15945 ( .A1(n13869), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15702), 
        .B2(n13805), .ZN(n13806) );
  OAI21_X1 U15946 ( .B1(n14014), .B2(n13913), .A(n13806), .ZN(n13807) );
  AOI21_X1 U15947 ( .B1(n13953), .B2(n13919), .A(n13807), .ZN(n13808) );
  OAI21_X1 U15948 ( .B1(n13809), .B2(n13869), .A(n13808), .ZN(P3_U3213) );
  OAI211_X1 U15949 ( .C1(n13811), .C2(n13815), .A(n13810), .B(n13874), .ZN(
        n13814) );
  AOI22_X1 U15950 ( .A1(n13812), .A2(n13877), .B1(n13880), .B2(n13842), .ZN(
        n13813) );
  NAND2_X1 U15951 ( .A1(n13814), .A2(n13813), .ZN(n13956) );
  INV_X1 U15952 ( .A(n13956), .ZN(n13823) );
  XNOR2_X1 U15953 ( .A(n13816), .B(n13815), .ZN(n13957) );
  INV_X1 U15954 ( .A(n13817), .ZN(n14018) );
  NOR2_X1 U15955 ( .A1(n14018), .A2(n13913), .ZN(n13821) );
  OAI22_X1 U15956 ( .A1(n15703), .A2(n13819), .B1(n13818), .B2(n13914), .ZN(
        n13820) );
  AOI211_X1 U15957 ( .C1(n13957), .C2(n13919), .A(n13821), .B(n13820), .ZN(
        n13822) );
  OAI21_X1 U15958 ( .B1(n13823), .B2(n13869), .A(n13822), .ZN(P3_U3214) );
  AOI21_X1 U15959 ( .B1(n9106), .B2(n13825), .A(n13824), .ZN(n13826) );
  OAI222_X1 U15960 ( .A1(n15690), .A2(n13828), .B1(n15689), .B2(n13827), .C1(
        n15696), .C2(n13826), .ZN(n13962) );
  INV_X1 U15961 ( .A(n13962), .ZN(n13837) );
  OAI22_X1 U15962 ( .A1(n15703), .A2(n13830), .B1(n13829), .B2(n13914), .ZN(
        n13835) );
  INV_X1 U15963 ( .A(n13963), .ZN(n13833) );
  AND2_X1 U15964 ( .A1(n13832), .A2(n13831), .ZN(n13961) );
  NOR3_X1 U15965 ( .A1(n13833), .A2(n13961), .A3(n13905), .ZN(n13834) );
  AOI211_X1 U15966 ( .C1(n13901), .C2(n13960), .A(n13835), .B(n13834), .ZN(
        n13836) );
  OAI21_X1 U15967 ( .B1(n13837), .B2(n13921), .A(n13836), .ZN(P3_U3215) );
  NAND2_X1 U15968 ( .A1(n13851), .A2(n13838), .ZN(n13840) );
  NAND2_X1 U15969 ( .A1(n13840), .A2(n13839), .ZN(n13841) );
  XNOR2_X1 U15970 ( .A(n13841), .B(n13847), .ZN(n13844) );
  AOI222_X1 U15971 ( .A1(n13874), .A2(n13844), .B1(n13843), .B2(n13880), .C1(
        n13842), .C2(n13877), .ZN(n13970) );
  OAI22_X1 U15972 ( .A1(n15703), .A2(n15127), .B1(n13845), .B2(n13914), .ZN(
        n13846) );
  AOI21_X1 U15973 ( .B1(n13967), .B2(n13901), .A(n13846), .ZN(n13850) );
  XNOR2_X1 U15974 ( .A(n13848), .B(n13847), .ZN(n13968) );
  NAND2_X1 U15975 ( .A1(n13968), .A2(n13919), .ZN(n13849) );
  OAI211_X1 U15976 ( .C1(n13970), .C2(n13869), .A(n13850), .B(n13849), .ZN(
        P3_U3216) );
  XNOR2_X1 U15977 ( .A(n13851), .B(n13857), .ZN(n13853) );
  AOI222_X1 U15978 ( .A1(n13874), .A2(n13853), .B1(n13878), .B2(n13880), .C1(
        n13852), .C2(n13877), .ZN(n13974) );
  OAI22_X1 U15979 ( .A1(n15703), .A2(n13854), .B1(n6707), .B2(n13914), .ZN(
        n13855) );
  AOI21_X1 U15980 ( .B1(n13971), .B2(n13901), .A(n13855), .ZN(n13860) );
  OAI21_X1 U15981 ( .B1(n13858), .B2(n13857), .A(n13856), .ZN(n13972) );
  NAND2_X1 U15982 ( .A1(n13972), .A2(n13919), .ZN(n13859) );
  OAI211_X1 U15983 ( .C1(n13974), .C2(n13869), .A(n13860), .B(n13859), .ZN(
        P3_U3217) );
  XNOR2_X1 U15984 ( .A(n13862), .B(n13861), .ZN(n13863) );
  OAI222_X1 U15985 ( .A1(n15690), .A2(n13896), .B1(n15689), .B2(n13864), .C1(
        n13863), .C2(n15696), .ZN(n13975) );
  INV_X1 U15986 ( .A(n13975), .ZN(n13873) );
  XNOR2_X1 U15987 ( .A(n13866), .B(n13865), .ZN(n13976) );
  INV_X1 U15988 ( .A(n13867), .ZN(n13868) );
  AOI22_X1 U15989 ( .A1(n13869), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15702), 
        .B2(n13868), .ZN(n13870) );
  OAI21_X1 U15990 ( .B1(n14028), .B2(n13913), .A(n13870), .ZN(n13871) );
  AOI21_X1 U15991 ( .B1(n13976), .B2(n13919), .A(n13871), .ZN(n13872) );
  OAI21_X1 U15992 ( .B1(n13873), .B2(n13921), .A(n13872), .ZN(P3_U3218) );
  OAI211_X1 U15993 ( .C1(n13876), .C2(n13883), .A(n13875), .B(n13874), .ZN(
        n13882) );
  AOI22_X1 U15994 ( .A1(n13880), .A2(n13879), .B1(n13878), .B2(n13877), .ZN(
        n13881) );
  NAND2_X1 U15995 ( .A1(n13882), .A2(n13881), .ZN(n13979) );
  INV_X1 U15996 ( .A(n13979), .ZN(n13890) );
  XNOR2_X1 U15997 ( .A(n13884), .B(n13883), .ZN(n13980) );
  NOR2_X1 U15998 ( .A1(n14032), .A2(n13913), .ZN(n13888) );
  INV_X1 U15999 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n13886) );
  OAI22_X1 U16000 ( .A1(n15703), .A2(n13886), .B1(n13885), .B2(n13914), .ZN(
        n13887) );
  AOI211_X1 U16001 ( .C1(n13980), .C2(n13919), .A(n13888), .B(n13887), .ZN(
        n13889) );
  OAI21_X1 U16002 ( .B1(n13890), .B2(n13921), .A(n13889), .ZN(P3_U3219) );
  XNOR2_X1 U16003 ( .A(n13892), .B(n13891), .ZN(n15143) );
  XNOR2_X1 U16004 ( .A(n13894), .B(n13893), .ZN(n13895) );
  OAI222_X1 U16005 ( .A1(n15690), .A2(n13897), .B1(n15689), .B2(n13896), .C1(
        n13895), .C2(n15696), .ZN(n15145) );
  NAND2_X1 U16006 ( .A1(n15145), .A2(n15703), .ZN(n13904) );
  OAI22_X1 U16007 ( .A1(n15703), .A2(n13899), .B1(n13898), .B2(n13914), .ZN(
        n13900) );
  AOI21_X1 U16008 ( .B1(n13902), .B2(n13901), .A(n13900), .ZN(n13903) );
  OAI211_X1 U16009 ( .C1(n13905), .C2(n15143), .A(n13904), .B(n13903), .ZN(
        P3_U3220) );
  XNOR2_X1 U16010 ( .A(n13907), .B(n13906), .ZN(n13908) );
  OAI222_X1 U16011 ( .A1(n15689), .A2(n7491), .B1(n15690), .B2(n13909), .C1(
        n13908), .C2(n15696), .ZN(n15147) );
  INV_X1 U16012 ( .A(n15147), .ZN(n13922) );
  OAI21_X1 U16013 ( .B1(n13912), .B2(n13911), .A(n13910), .ZN(n15149) );
  NOR2_X1 U16014 ( .A1(n13913), .A2(n15146), .ZN(n13918) );
  OAI22_X1 U16015 ( .A1(n15703), .A2(n13916), .B1(n13915), .B2(n13914), .ZN(
        n13917) );
  AOI211_X1 U16016 ( .C1(n15149), .C2(n13919), .A(n13918), .B(n13917), .ZN(
        n13920) );
  OAI21_X1 U16017 ( .B1(n13922), .B2(n13921), .A(n13920), .ZN(P3_U3221) );
  NOR2_X1 U16018 ( .A1(n13984), .A2(n15739), .ZN(n13925) );
  AOI21_X1 U16019 ( .B1(P3_REG1_REG_31__SCAN_IN), .B2(n15739), .A(n13925), 
        .ZN(n13923) );
  OAI21_X1 U16020 ( .B1(n13986), .B2(n13983), .A(n13923), .ZN(P3_U3490) );
  NAND2_X1 U16021 ( .A1(n13924), .A2(n10189), .ZN(n13927) );
  INV_X1 U16022 ( .A(n13925), .ZN(n13926) );
  OAI211_X1 U16023 ( .C1(n15741), .C2(n9324), .A(n13927), .B(n13926), .ZN(
        P3_U3489) );
  OAI21_X1 U16024 ( .B1(n15726), .B2(n13929), .A(n13928), .ZN(n13990) );
  MUX2_X1 U16025 ( .A(P3_REG1_REG_28__SCAN_IN), .B(n13990), .S(n15741), .Z(
        n13930) );
  INV_X1 U16026 ( .A(n13930), .ZN(n13931) );
  OAI21_X1 U16027 ( .B1(n13993), .B2(n13983), .A(n13931), .ZN(P3_U3487) );
  AOI21_X1 U16028 ( .B1(n15716), .B2(n13933), .A(n13932), .ZN(n13994) );
  MUX2_X1 U16029 ( .A(n13934), .B(n13994), .S(n15741), .Z(n13935) );
  OAI21_X1 U16030 ( .B1(n13997), .B2(n13983), .A(n13935), .ZN(P3_U3484) );
  AOI21_X1 U16031 ( .B1(n15731), .B2(n13937), .A(n13936), .ZN(n13938) );
  OAI21_X1 U16032 ( .B1(n15726), .B2(n13939), .A(n13938), .ZN(n13998) );
  MUX2_X1 U16033 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n13998), .S(n15741), .Z(
        P3_U3483) );
  AOI21_X1 U16034 ( .B1(n13941), .B2(n15724), .A(n13940), .ZN(n13999) );
  MUX2_X1 U16035 ( .A(n13942), .B(n13999), .S(n15741), .Z(n13943) );
  OAI21_X1 U16036 ( .B1(n14002), .B2(n13983), .A(n13943), .ZN(P3_U3482) );
  INV_X1 U16037 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13946) );
  AOI21_X1 U16038 ( .B1(n15724), .B2(n13945), .A(n13944), .ZN(n14003) );
  MUX2_X1 U16039 ( .A(n13946), .B(n14003), .S(n15741), .Z(n13947) );
  OAI21_X1 U16040 ( .B1(n14006), .B2(n13983), .A(n13947), .ZN(P3_U3481) );
  INV_X1 U16041 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13950) );
  AOI21_X1 U16042 ( .B1(n15724), .B2(n13949), .A(n13948), .ZN(n14007) );
  MUX2_X1 U16043 ( .A(n13950), .B(n14007), .S(n15741), .Z(n13951) );
  OAI21_X1 U16044 ( .B1(n14010), .B2(n13983), .A(n13951), .ZN(P3_U3480) );
  AOI21_X1 U16045 ( .B1(n13953), .B2(n15724), .A(n13952), .ZN(n14011) );
  MUX2_X1 U16046 ( .A(n13954), .B(n14011), .S(n15741), .Z(n13955) );
  OAI21_X1 U16047 ( .B1(n14014), .B2(n13983), .A(n13955), .ZN(P3_U3479) );
  AOI21_X1 U16048 ( .B1(n15724), .B2(n13957), .A(n13956), .ZN(n14015) );
  MUX2_X1 U16049 ( .A(n13958), .B(n14015), .S(n15741), .Z(n13959) );
  OAI21_X1 U16050 ( .B1(n14018), .B2(n13983), .A(n13959), .ZN(P3_U3478) );
  INV_X1 U16051 ( .A(n13960), .ZN(n14022) );
  NOR2_X1 U16052 ( .A1(n13961), .A2(n15726), .ZN(n13964) );
  AOI21_X1 U16053 ( .B1(n13964), .B2(n13963), .A(n13962), .ZN(n14019) );
  MUX2_X1 U16054 ( .A(n13965), .B(n14019), .S(n15741), .Z(n13966) );
  OAI21_X1 U16055 ( .B1(n14022), .B2(n13983), .A(n13966), .ZN(P3_U3477) );
  AOI22_X1 U16056 ( .A1(n13968), .A2(n15724), .B1(n15731), .B2(n13967), .ZN(
        n13969) );
  NAND2_X1 U16057 ( .A1(n13970), .A2(n13969), .ZN(n14023) );
  MUX2_X1 U16058 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n14023), .S(n15741), .Z(
        P3_U3476) );
  AOI22_X1 U16059 ( .A1(n13972), .A2(n15724), .B1(n15731), .B2(n13971), .ZN(
        n13973) );
  NAND2_X1 U16060 ( .A1(n13974), .A2(n13973), .ZN(n14024) );
  MUX2_X1 U16061 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n14024), .S(n15741), .Z(
        P3_U3475) );
  AOI21_X1 U16062 ( .B1(n13976), .B2(n15724), .A(n13975), .ZN(n14025) );
  MUX2_X1 U16063 ( .A(n13977), .B(n14025), .S(n15741), .Z(n13978) );
  OAI21_X1 U16064 ( .B1(n14028), .B2(n13983), .A(n13978), .ZN(P3_U3474) );
  AOI21_X1 U16065 ( .B1(n13980), .B2(n15724), .A(n13979), .ZN(n14029) );
  MUX2_X1 U16066 ( .A(n13981), .B(n14029), .S(n15741), .Z(n13982) );
  OAI21_X1 U16067 ( .B1(n13983), .B2(n14032), .A(n13982), .ZN(P3_U3473) );
  NOR2_X1 U16068 ( .A1(n13984), .A2(n15732), .ZN(n13987) );
  AOI21_X1 U16069 ( .B1(P3_REG0_REG_31__SCAN_IN), .B2(n15732), .A(n13987), 
        .ZN(n13985) );
  OAI21_X1 U16070 ( .B1(n13986), .B2(n14033), .A(n13985), .ZN(P3_U3458) );
  AOI21_X1 U16071 ( .B1(P3_REG0_REG_30__SCAN_IN), .B2(n15732), .A(n13987), 
        .ZN(n13988) );
  OAI21_X1 U16072 ( .B1(n13989), .B2(n14033), .A(n13988), .ZN(P3_U3457) );
  MUX2_X1 U16073 ( .A(P3_REG0_REG_28__SCAN_IN), .B(n13990), .S(n15734), .Z(
        n13991) );
  INV_X1 U16074 ( .A(n13991), .ZN(n13992) );
  OAI21_X1 U16075 ( .B1(n13993), .B2(n14033), .A(n13992), .ZN(P3_U3455) );
  INV_X1 U16076 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13995) );
  MUX2_X1 U16077 ( .A(n13995), .B(n13994), .S(n15734), .Z(n13996) );
  OAI21_X1 U16078 ( .B1(n13997), .B2(n14033), .A(n13996), .ZN(P3_U3452) );
  MUX2_X1 U16079 ( .A(P3_REG0_REG_24__SCAN_IN), .B(n13998), .S(n15734), .Z(
        P3_U3451) );
  INV_X1 U16080 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n14000) );
  MUX2_X1 U16081 ( .A(n14000), .B(n13999), .S(n15734), .Z(n14001) );
  OAI21_X1 U16082 ( .B1(n14002), .B2(n14033), .A(n14001), .ZN(P3_U3450) );
  INV_X1 U16083 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n14004) );
  MUX2_X1 U16084 ( .A(n14004), .B(n14003), .S(n15734), .Z(n14005) );
  OAI21_X1 U16085 ( .B1(n14006), .B2(n14033), .A(n14005), .ZN(P3_U3449) );
  INV_X1 U16086 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n14008) );
  MUX2_X1 U16087 ( .A(n14008), .B(n14007), .S(n15734), .Z(n14009) );
  OAI21_X1 U16088 ( .B1(n14010), .B2(n14033), .A(n14009), .ZN(P3_U3448) );
  INV_X1 U16089 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n14012) );
  MUX2_X1 U16090 ( .A(n14012), .B(n14011), .S(n15734), .Z(n14013) );
  OAI21_X1 U16091 ( .B1(n14014), .B2(n14033), .A(n14013), .ZN(P3_U3447) );
  INV_X1 U16092 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n14016) );
  MUX2_X1 U16093 ( .A(n14016), .B(n14015), .S(n15734), .Z(n14017) );
  OAI21_X1 U16094 ( .B1(n14018), .B2(n14033), .A(n14017), .ZN(P3_U3446) );
  INV_X1 U16095 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n14020) );
  MUX2_X1 U16096 ( .A(n14020), .B(n14019), .S(n15734), .Z(n14021) );
  OAI21_X1 U16097 ( .B1(n14022), .B2(n14033), .A(n14021), .ZN(P3_U3444) );
  MUX2_X1 U16098 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n14023), .S(n15734), .Z(
        P3_U3441) );
  MUX2_X1 U16099 ( .A(P3_REG0_REG_16__SCAN_IN), .B(n14024), .S(n15734), .Z(
        P3_U3438) );
  INV_X1 U16100 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n14026) );
  MUX2_X1 U16101 ( .A(n14026), .B(n14025), .S(n15734), .Z(n14027) );
  OAI21_X1 U16102 ( .B1(n14028), .B2(n14033), .A(n14027), .ZN(P3_U3435) );
  MUX2_X1 U16103 ( .A(n14030), .B(n14029), .S(n15734), .Z(n14031) );
  OAI21_X1 U16104 ( .B1(n14033), .B2(n14032), .A(n14031), .ZN(P3_U3432) );
  MUX2_X1 U16105 ( .A(P3_D_REG_1__SCAN_IN), .B(n14034), .S(n14035), .Z(
        P3_U3377) );
  MUX2_X1 U16106 ( .A(P3_D_REG_0__SCAN_IN), .B(n14036), .S(n14035), .Z(
        P3_U3376) );
  NAND2_X1 U16107 ( .A1(n14038), .A2(n14037), .ZN(n14043) );
  INV_X1 U16108 ( .A(n14039), .ZN(n14041) );
  OR4_X1 U16109 ( .A1(n14041), .A2(P3_IR_REG_30__SCAN_IN), .A3(n14040), .A4(
        P3_U3151), .ZN(n14042) );
  OAI211_X1 U16110 ( .C1(n14044), .C2(n14049), .A(n14043), .B(n14042), .ZN(
        P3_U3264) );
  INV_X1 U16111 ( .A(n14045), .ZN(n14047) );
  OAI222_X1 U16112 ( .A1(n14049), .A2(n14048), .B1(n12850), .B2(n14047), .C1(
        n14046), .C2(P3_U3151), .ZN(P3_U3266) );
  AOI22_X1 U16113 ( .A1(n14107), .A2(n14233), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14055) );
  AOI22_X1 U16114 ( .A1(n14108), .A2(n14228), .B1(n14109), .B2(n14229), .ZN(
        n14054) );
  NAND2_X1 U16115 ( .A1(n14415), .A2(n14146), .ZN(n14053) );
  NAND4_X1 U16116 ( .A1(n14056), .A2(n14055), .A3(n14054), .A4(n14053), .ZN(
        P2_U3186) );
  OAI211_X1 U16117 ( .C1(n14059), .C2(n14058), .A(n14057), .B(n14103), .ZN(
        n14064) );
  AND2_X1 U16118 ( .A1(n14151), .A2(n14369), .ZN(n14060) );
  AOI21_X1 U16119 ( .B1(n14335), .B2(n14368), .A(n14060), .ZN(n14304) );
  INV_X1 U16120 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n14061) );
  OAI22_X1 U16121 ( .A1(n14304), .A2(n14096), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14061), .ZN(n14062) );
  AOI21_X1 U16122 ( .B1(n14309), .B2(n14107), .A(n14062), .ZN(n14063) );
  OAI211_X1 U16123 ( .C1(n7227), .C2(n14102), .A(n14064), .B(n14063), .ZN(
        P2_U3188) );
  INV_X1 U16124 ( .A(n14375), .ZN(n14509) );
  OAI21_X1 U16125 ( .B1(n14067), .B2(n14066), .A(n14065), .ZN(n14068) );
  NAND2_X1 U16126 ( .A1(n14068), .A2(n14103), .ZN(n14074) );
  INV_X1 U16127 ( .A(n14069), .ZN(n14376) );
  OAI22_X1 U16128 ( .A1(n14071), .A2(n14143), .B1(n14142), .B2(n14070), .ZN(
        n14072) );
  AOI211_X1 U16129 ( .C1(n14107), .C2(n14376), .A(n6819), .B(n14072), .ZN(
        n14073) );
  OAI211_X1 U16130 ( .C1(n14509), .C2(n14102), .A(n14074), .B(n14073), .ZN(
        P2_U3191) );
  OAI211_X1 U16131 ( .C1(n14077), .C2(n14076), .A(n14075), .B(n14103), .ZN(
        n14081) );
  AOI22_X1 U16132 ( .A1(n14339), .A2(n14107), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14080) );
  AOI22_X1 U16133 ( .A1(n14335), .A2(n14108), .B1(n14109), .B2(n14370), .ZN(
        n14079) );
  NAND2_X1 U16134 ( .A1(n14338), .A2(n14146), .ZN(n14078) );
  NAND4_X1 U16135 ( .A1(n14081), .A2(n14080), .A3(n14079), .A4(n14078), .ZN(
        P2_U3195) );
  OAI211_X1 U16136 ( .C1(n14084), .C2(n14083), .A(n14082), .B(n14103), .ZN(
        n14089) );
  AOI22_X1 U16137 ( .A1(n14107), .A2(n14272), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14088) );
  AOI22_X1 U16138 ( .A1(n14109), .A2(n14151), .B1(n14108), .B2(n14229), .ZN(
        n14087) );
  NAND2_X1 U16139 ( .A1(n14085), .A2(n14146), .ZN(n14086) );
  NAND4_X1 U16140 ( .A1(n14089), .A2(n14088), .A3(n14087), .A4(n14086), .ZN(
        P2_U3197) );
  AND2_X1 U16141 ( .A1(n14090), .A2(n14125), .ZN(n14094) );
  NAND2_X1 U16142 ( .A1(n7244), .A2(n14092), .ZN(n14093) );
  NAND2_X1 U16143 ( .A1(n14093), .A2(n14094), .ZN(n14126) );
  OAI21_X1 U16144 ( .B1(n14094), .B2(n14093), .A(n14126), .ZN(n14095) );
  NAND2_X1 U16145 ( .A1(n14095), .A2(n14103), .ZN(n14101) );
  NAND2_X1 U16146 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n15472)
         );
  OAI21_X1 U16147 ( .B1(n14097), .B2(n14096), .A(n15472), .ZN(n14098) );
  AOI21_X1 U16148 ( .B1(n14099), .B2(n14107), .A(n14098), .ZN(n14100) );
  OAI211_X1 U16149 ( .C1(n14518), .C2(n14102), .A(n14101), .B(n14100), .ZN(
        P2_U3200) );
  OAI211_X1 U16150 ( .C1(n14106), .C2(n14105), .A(n14104), .B(n14103), .ZN(
        n14113) );
  AOI22_X1 U16151 ( .A1(n14107), .A2(n14290), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14112) );
  AOI22_X1 U16152 ( .A1(n14152), .A2(n14109), .B1(n14108), .B2(n14254), .ZN(
        n14111) );
  NAND2_X1 U16153 ( .A1(n14430), .A2(n14146), .ZN(n14110) );
  NAND4_X1 U16154 ( .A1(n14113), .A2(n14112), .A3(n14111), .A4(n14110), .ZN(
        P2_U3201) );
  INV_X1 U16155 ( .A(n14114), .ZN(n14116) );
  NAND2_X1 U16156 ( .A1(n14116), .A2(n14115), .ZN(n14117) );
  XNOR2_X1 U16157 ( .A(n14118), .B(n14117), .ZN(n14124) );
  INV_X1 U16158 ( .A(n14350), .ZN(n14120) );
  OAI22_X1 U16159 ( .A1(n14120), .A2(n14140), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14119), .ZN(n14122) );
  OAI22_X1 U16160 ( .A1(n14324), .A2(n14142), .B1(n14143), .B2(n14130), .ZN(
        n14121) );
  AOI211_X1 U16161 ( .C1(n14454), .C2(n14146), .A(n14122), .B(n14121), .ZN(
        n14123) );
  OAI21_X1 U16162 ( .B1(n14124), .B2(n14148), .A(n14123), .ZN(P2_U3205) );
  NAND2_X1 U16163 ( .A1(n14126), .A2(n14125), .ZN(n14127) );
  XOR2_X1 U16164 ( .A(n14128), .B(n14127), .Z(n14135) );
  OAI22_X1 U16165 ( .A1(n14130), .A2(n14325), .B1(n14129), .B2(n14323), .ZN(
        n14393) );
  AOI22_X1 U16166 ( .A1(n14393), .A2(n14131), .B1(P2_REG3_REG_18__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14132) );
  OAI21_X1 U16167 ( .B1(n14386), .B2(n14140), .A(n14132), .ZN(n14133) );
  AOI21_X1 U16168 ( .B1(n14390), .B2(n14146), .A(n14133), .ZN(n14134) );
  OAI21_X1 U16169 ( .B1(n14135), .B2(n14148), .A(n14134), .ZN(P2_U3210) );
  INV_X1 U16170 ( .A(n14247), .ZN(n14139) );
  OAI22_X1 U16171 ( .A1(n14140), .A2(n14139), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14138), .ZN(n14145) );
  OAI22_X1 U16172 ( .A1(n14286), .A2(n14143), .B1(n14142), .B2(n14141), .ZN(
        n14144) );
  AOI211_X1 U16173 ( .C1(n14420), .C2(n14146), .A(n14145), .B(n14144), .ZN(
        n14147) );
  OAI21_X1 U16174 ( .B1(n6775), .B2(n14148), .A(n14147), .ZN(P2_U3212) );
  INV_X2 U16175 ( .A(P2_U3947), .ZN(n14168) );
  MUX2_X1 U16176 ( .A(n14206), .B(P2_DATAO_REG_31__SCAN_IN), .S(n14168), .Z(
        P2_U3562) );
  MUX2_X1 U16177 ( .A(n14149), .B(P2_DATAO_REG_30__SCAN_IN), .S(n14168), .Z(
        P2_U3561) );
  MUX2_X1 U16178 ( .A(n14150), .B(P2_DATAO_REG_29__SCAN_IN), .S(n14168), .Z(
        P2_U3560) );
  MUX2_X1 U16179 ( .A(n14228), .B(P2_DATAO_REG_28__SCAN_IN), .S(n14168), .Z(
        P2_U3559) );
  MUX2_X1 U16180 ( .A(n14255), .B(P2_DATAO_REG_27__SCAN_IN), .S(n14168), .Z(
        P2_U3558) );
  MUX2_X1 U16181 ( .A(n14229), .B(P2_DATAO_REG_26__SCAN_IN), .S(n14168), .Z(
        P2_U3557) );
  MUX2_X1 U16182 ( .A(n14254), .B(P2_DATAO_REG_25__SCAN_IN), .S(n14168), .Z(
        P2_U3556) );
  MUX2_X1 U16183 ( .A(n14151), .B(P2_DATAO_REG_24__SCAN_IN), .S(n14168), .Z(
        P2_U3555) );
  MUX2_X1 U16184 ( .A(n14152), .B(P2_DATAO_REG_23__SCAN_IN), .S(n14168), .Z(
        P2_U3554) );
  MUX2_X1 U16185 ( .A(n14335), .B(P2_DATAO_REG_22__SCAN_IN), .S(n14168), .Z(
        P2_U3553) );
  MUX2_X1 U16186 ( .A(n14355), .B(P2_DATAO_REG_21__SCAN_IN), .S(n14168), .Z(
        P2_U3552) );
  MUX2_X1 U16187 ( .A(n14370), .B(P2_DATAO_REG_20__SCAN_IN), .S(n14168), .Z(
        P2_U3551) );
  MUX2_X1 U16188 ( .A(n14356), .B(P2_DATAO_REG_19__SCAN_IN), .S(n14168), .Z(
        P2_U3550) );
  MUX2_X1 U16189 ( .A(n14367), .B(P2_DATAO_REG_18__SCAN_IN), .S(n14168), .Z(
        P2_U3549) );
  MUX2_X1 U16190 ( .A(n14153), .B(P2_DATAO_REG_17__SCAN_IN), .S(n14168), .Z(
        P2_U3548) );
  MUX2_X1 U16191 ( .A(n14154), .B(P2_DATAO_REG_16__SCAN_IN), .S(n14168), .Z(
        P2_U3547) );
  MUX2_X1 U16192 ( .A(n14155), .B(P2_DATAO_REG_15__SCAN_IN), .S(n14168), .Z(
        P2_U3546) );
  MUX2_X1 U16193 ( .A(n14156), .B(P2_DATAO_REG_14__SCAN_IN), .S(n14168), .Z(
        P2_U3545) );
  MUX2_X1 U16194 ( .A(n14157), .B(P2_DATAO_REG_13__SCAN_IN), .S(n14168), .Z(
        P2_U3544) );
  MUX2_X1 U16195 ( .A(n14158), .B(P2_DATAO_REG_12__SCAN_IN), .S(n14168), .Z(
        P2_U3543) );
  MUX2_X1 U16196 ( .A(n14159), .B(P2_DATAO_REG_11__SCAN_IN), .S(n14168), .Z(
        P2_U3542) );
  MUX2_X1 U16197 ( .A(n14160), .B(P2_DATAO_REG_10__SCAN_IN), .S(n14168), .Z(
        P2_U3541) );
  MUX2_X1 U16198 ( .A(n14161), .B(P2_DATAO_REG_9__SCAN_IN), .S(n14168), .Z(
        P2_U3540) );
  MUX2_X1 U16199 ( .A(n14162), .B(P2_DATAO_REG_8__SCAN_IN), .S(n14168), .Z(
        P2_U3539) );
  MUX2_X1 U16200 ( .A(n14163), .B(P2_DATAO_REG_7__SCAN_IN), .S(n14168), .Z(
        P2_U3538) );
  MUX2_X1 U16201 ( .A(n14164), .B(P2_DATAO_REG_6__SCAN_IN), .S(n14168), .Z(
        P2_U3537) );
  MUX2_X1 U16202 ( .A(n14165), .B(P2_DATAO_REG_5__SCAN_IN), .S(n14168), .Z(
        P2_U3536) );
  MUX2_X1 U16203 ( .A(n14166), .B(P2_DATAO_REG_4__SCAN_IN), .S(n14168), .Z(
        P2_U3535) );
  MUX2_X1 U16204 ( .A(n14167), .B(P2_DATAO_REG_3__SCAN_IN), .S(n14168), .Z(
        P2_U3534) );
  MUX2_X1 U16205 ( .A(n14169), .B(P2_DATAO_REG_2__SCAN_IN), .S(n14168), .Z(
        P2_U3533) );
  MUX2_X1 U16206 ( .A(n14170), .B(P2_DATAO_REG_1__SCAN_IN), .S(n14168), .Z(
        P2_U3532) );
  AOI211_X1 U16207 ( .C1(n14173), .C2(n14172), .A(n14171), .B(n15461), .ZN(
        n14174) );
  INV_X1 U16208 ( .A(n14174), .ZN(n14182) );
  AOI22_X1 U16209 ( .A1(n15333), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n14181) );
  NAND2_X1 U16210 ( .A1(n7092), .A2(n14175), .ZN(n14180) );
  OAI211_X1 U16211 ( .C1(n14178), .C2(n14177), .A(n15484), .B(n14176), .ZN(
        n14179) );
  NAND4_X1 U16212 ( .A1(n14182), .A2(n14181), .A3(n14180), .A4(n14179), .ZN(
        P2_U3216) );
  AOI21_X1 U16213 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n14184), .A(n14183), 
        .ZN(n14185) );
  NOR2_X1 U16214 ( .A1(n14185), .A2(n15437), .ZN(n14186) );
  INV_X1 U16215 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n15441) );
  XNOR2_X1 U16216 ( .A(n15437), .B(n14185), .ZN(n15442) );
  NOR2_X1 U16217 ( .A1(n15441), .A2(n15442), .ZN(n15440) );
  NOR2_X1 U16218 ( .A1(n14186), .A2(n15440), .ZN(n15451) );
  XNOR2_X1 U16219 ( .A(n15457), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n15450) );
  NOR2_X1 U16220 ( .A1(n15451), .A2(n15450), .ZN(n15449) );
  AOI21_X1 U16221 ( .B1(n15457), .B2(P2_REG1_REG_16__SCAN_IN), .A(n15449), 
        .ZN(n15468) );
  XNOR2_X1 U16222 ( .A(n15471), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n15467) );
  NOR2_X1 U16223 ( .A1(n15468), .A2(n15467), .ZN(n15466) );
  AOI21_X1 U16224 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n15471), .A(n15466), 
        .ZN(n14187) );
  NOR2_X1 U16225 ( .A1(n14187), .A2(n15488), .ZN(n14188) );
  XNOR2_X1 U16226 ( .A(n15488), .B(n14187), .ZN(n15481) );
  NOR2_X1 U16227 ( .A1(n15480), .A2(n15481), .ZN(n15482) );
  NOR2_X1 U16228 ( .A1(n14188), .A2(n15482), .ZN(n14189) );
  XOR2_X1 U16229 ( .A(n14189), .B(n14461), .Z(n14200) );
  INV_X1 U16230 ( .A(n14200), .ZN(n14198) );
  NOR2_X1 U16231 ( .A1(n14192), .A2(n15437), .ZN(n14193) );
  NOR2_X1 U16232 ( .A1(n12372), .A2(n15439), .ZN(n15438) );
  NAND2_X1 U16233 ( .A1(n15457), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n14194) );
  OAI21_X1 U16234 ( .B1(n15457), .B2(P2_REG2_REG_16__SCAN_IN), .A(n14194), 
        .ZN(n15453) );
  XNOR2_X1 U16235 ( .A(n15471), .B(P2_REG2_REG_17__SCAN_IN), .ZN(n15463) );
  INV_X1 U16236 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n15476) );
  NAND2_X1 U16237 ( .A1(n15477), .A2(n15476), .ZN(n15475) );
  NAND2_X1 U16238 ( .A1(n14195), .A2(n15488), .ZN(n14196) );
  NAND2_X1 U16239 ( .A1(n15475), .A2(n14196), .ZN(n14197) );
  XNOR2_X1 U16240 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n14197), .ZN(n14199) );
  NAND2_X1 U16241 ( .A1(n14489), .A2(n14210), .ZN(n14209) );
  XNOR2_X1 U16242 ( .A(n14209), .B(n14484), .ZN(n14203) );
  INV_X1 U16243 ( .A(n14204), .ZN(n14205) );
  NAND2_X1 U16244 ( .A1(n14206), .A2(n14205), .ZN(n14409) );
  NOR2_X1 U16245 ( .A1(n6677), .A2(n14409), .ZN(n14212) );
  AOI21_X1 U16246 ( .B1(n6677), .B2(P2_REG2_REG_31__SCAN_IN), .A(n14212), .ZN(
        n14208) );
  NAND2_X1 U16247 ( .A1(n14484), .A2(n14389), .ZN(n14207) );
  OAI211_X1 U16248 ( .C1(n14405), .C2(n14214), .A(n14208), .B(n14207), .ZN(
        P2_U3234) );
  OAI211_X1 U16249 ( .C1(n14489), .C2(n14210), .A(n14398), .B(n14209), .ZN(
        n14410) );
  NOR2_X1 U16250 ( .A1(n14489), .A2(n15503), .ZN(n14211) );
  AOI211_X1 U16251 ( .C1(n6677), .C2(P2_REG2_REG_30__SCAN_IN), .A(n14212), .B(
        n14211), .ZN(n14213) );
  OAI21_X1 U16252 ( .B1(n14214), .B2(n14410), .A(n14213), .ZN(P2_U3235) );
  INV_X1 U16253 ( .A(n14215), .ZN(n14224) );
  NAND2_X1 U16254 ( .A1(n14216), .A2(n15498), .ZN(n14219) );
  AOI22_X1 U16255 ( .A1(n6677), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n14217), 
        .B2(n15499), .ZN(n14218) );
  OAI211_X1 U16256 ( .C1(n14220), .C2(n15503), .A(n14219), .B(n14218), .ZN(
        n14221) );
  AOI21_X1 U16257 ( .B1(n14222), .B2(n14397), .A(n14221), .ZN(n14223) );
  OAI21_X1 U16258 ( .B1(n14224), .B2(n14362), .A(n14223), .ZN(P2_U3236) );
  NAND3_X1 U16259 ( .A1(n14253), .A2(n7305), .A3(n14225), .ZN(n14226) );
  NAND2_X1 U16260 ( .A1(n14227), .A2(n14226), .ZN(n14230) );
  AOI222_X1 U16261 ( .A1(n14358), .A2(n14230), .B1(n14229), .B2(n14368), .C1(
        n14228), .C2(n14369), .ZN(n14417) );
  INV_X1 U16262 ( .A(n14231), .ZN(n14232) );
  AOI211_X1 U16263 ( .C1(n14415), .C2(n14244), .A(n12878), .B(n14232), .ZN(
        n14414) );
  AOI22_X1 U16264 ( .A1(n6677), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n14233), 
        .B2(n15499), .ZN(n14234) );
  OAI21_X1 U16265 ( .B1(n14235), .B2(n15503), .A(n14234), .ZN(n14236) );
  AOI21_X1 U16266 ( .B1(n14414), .B2(n15498), .A(n14236), .ZN(n14241) );
  NAND2_X1 U16267 ( .A1(n14239), .A2(n14238), .ZN(n14413) );
  NAND3_X1 U16268 ( .A1(n14237), .A2(n14413), .A3(n15496), .ZN(n14240) );
  OAI211_X1 U16269 ( .C1(n14417), .C2(n6677), .A(n14241), .B(n14240), .ZN(
        P2_U3238) );
  XNOR2_X1 U16270 ( .A(n14243), .B(n14242), .ZN(n14423) );
  INV_X1 U16271 ( .A(n14270), .ZN(n14246) );
  INV_X1 U16272 ( .A(n14244), .ZN(n14245) );
  AOI211_X1 U16273 ( .C1(n14420), .C2(n14246), .A(n12878), .B(n14245), .ZN(
        n14419) );
  AOI22_X1 U16274 ( .A1(n6677), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n14247), 
        .B2(n15499), .ZN(n14248) );
  OAI21_X1 U16275 ( .B1(n14249), .B2(n15503), .A(n14248), .ZN(n14258) );
  NAND3_X1 U16276 ( .A1(n14266), .A2(n14251), .A3(n14250), .ZN(n14252) );
  NAND2_X1 U16277 ( .A1(n14253), .A2(n14252), .ZN(n14256) );
  AOI222_X1 U16278 ( .A1(n14358), .A2(n14256), .B1(n14255), .B2(n14369), .C1(
        n14254), .C2(n14368), .ZN(n14422) );
  NOR2_X1 U16279 ( .A1(n14422), .A2(n6677), .ZN(n14257) );
  AOI211_X1 U16280 ( .C1(n14419), .C2(n15498), .A(n14258), .B(n14257), .ZN(
        n14259) );
  OAI21_X1 U16281 ( .B1(n14423), .B2(n14362), .A(n14259), .ZN(P2_U3239) );
  OAI21_X1 U16282 ( .B1(n6777), .B2(n14264), .A(n14260), .ZN(n14425) );
  INV_X1 U16283 ( .A(n14425), .ZN(n14277) );
  AND2_X1 U16284 ( .A1(n14262), .A2(n14261), .ZN(n14285) );
  NAND3_X1 U16285 ( .A1(n14285), .A2(n14264), .A3(n14263), .ZN(n14265) );
  AND2_X1 U16286 ( .A1(n14266), .A2(n14265), .ZN(n14267) );
  OAI222_X1 U16287 ( .A1(n14325), .A2(n14269), .B1(n14323), .B2(n14268), .C1(
        n14395), .C2(n14267), .ZN(n14424) );
  OAI21_X1 U16288 ( .B1(n14289), .B2(n14495), .A(n14398), .ZN(n14271) );
  NAND2_X1 U16289 ( .A1(n7603), .A2(n15498), .ZN(n14274) );
  AOI22_X1 U16290 ( .A1(n6677), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n14272), 
        .B2(n15499), .ZN(n14273) );
  OAI211_X1 U16291 ( .C1(n14495), .C2(n15503), .A(n14274), .B(n14273), .ZN(
        n14275) );
  AOI21_X1 U16292 ( .B1(n14424), .B2(n14397), .A(n14275), .ZN(n14276) );
  OAI21_X1 U16293 ( .B1(n14277), .B2(n14362), .A(n14276), .ZN(P2_U3240) );
  NAND2_X1 U16294 ( .A1(n14279), .A2(n14278), .ZN(n14280) );
  OR2_X1 U16295 ( .A1(n14300), .A2(n14299), .ZN(n14302) );
  NAND3_X1 U16296 ( .A1(n14302), .A2(n14283), .A3(n14282), .ZN(n14284) );
  AOI21_X1 U16297 ( .B1(n14285), .B2(n14284), .A(n14395), .ZN(n14288) );
  OAI22_X1 U16298 ( .A1(n14326), .A2(n14323), .B1(n14286), .B2(n14325), .ZN(
        n14287) );
  INV_X1 U16299 ( .A(n14430), .ZN(n14293) );
  AOI211_X1 U16300 ( .C1(n14430), .C2(n14307), .A(n12878), .B(n14289), .ZN(
        n14429) );
  NAND2_X1 U16301 ( .A1(n14429), .A2(n15498), .ZN(n14292) );
  AOI22_X1 U16302 ( .A1(n6677), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n14290), 
        .B2(n15499), .ZN(n14291) );
  OAI211_X1 U16303 ( .C1(n14293), .C2(n15503), .A(n14292), .B(n14291), .ZN(
        n14294) );
  AOI21_X1 U16304 ( .B1(n14428), .B2(n14295), .A(n14294), .ZN(n14296) );
  OAI21_X1 U16305 ( .B1(n14432), .B2(n6677), .A(n14296), .ZN(P2_U3241) );
  XNOR2_X1 U16306 ( .A(n14298), .B(n14297), .ZN(n14435) );
  INV_X1 U16307 ( .A(n14435), .ZN(n14314) );
  NAND2_X1 U16308 ( .A1(n14300), .A2(n14299), .ZN(n14301) );
  NAND2_X1 U16309 ( .A1(n14302), .A2(n14301), .ZN(n14303) );
  NAND2_X1 U16310 ( .A1(n14303), .A2(n14358), .ZN(n14305) );
  NAND2_X1 U16311 ( .A1(n14305), .A2(n14304), .ZN(n14437) );
  AOI21_X1 U16312 ( .B1(n14316), .B2(n14306), .A(n12878), .ZN(n14308) );
  AND2_X1 U16313 ( .A1(n14308), .A2(n14307), .ZN(n14436) );
  NAND2_X1 U16314 ( .A1(n14436), .A2(n15498), .ZN(n14311) );
  AOI22_X1 U16315 ( .A1(n14309), .A2(n15499), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(n6677), .ZN(n14310) );
  OAI211_X1 U16316 ( .C1(n7227), .C2(n15503), .A(n14311), .B(n14310), .ZN(
        n14312) );
  AOI21_X1 U16317 ( .B1(n14437), .B2(n14397), .A(n14312), .ZN(n14313) );
  OAI21_X1 U16318 ( .B1(n14314), .B2(n14362), .A(n14313), .ZN(P2_U3242) );
  OAI21_X1 U16319 ( .B1(n6739), .B2(n7228), .A(n14315), .ZN(n14446) );
  INV_X1 U16320 ( .A(n14316), .ZN(n14317) );
  AOI211_X1 U16321 ( .C1(n14443), .C2(n6990), .A(n12878), .B(n14317), .ZN(
        n14442) );
  INV_X1 U16322 ( .A(n14318), .ZN(n14319) );
  AOI22_X1 U16323 ( .A1(n14319), .A2(n15499), .B1(P2_REG2_REG_22__SCAN_IN), 
        .B2(n6677), .ZN(n14320) );
  OAI21_X1 U16324 ( .B1(n14321), .B2(n15503), .A(n14320), .ZN(n14331) );
  AOI21_X1 U16325 ( .B1(n14322), .B2(n7228), .A(n14395), .ZN(n14329) );
  OAI22_X1 U16326 ( .A1(n14326), .A2(n14325), .B1(n14324), .B2(n14323), .ZN(
        n14327) );
  AOI21_X1 U16327 ( .B1(n14329), .B2(n14328), .A(n14327), .ZN(n14445) );
  NOR2_X1 U16328 ( .A1(n14445), .A2(n6677), .ZN(n14330) );
  AOI211_X1 U16329 ( .C1(n14442), .C2(n15498), .A(n14331), .B(n14330), .ZN(
        n14332) );
  OAI21_X1 U16330 ( .B1(n14362), .B2(n14446), .A(n14332), .ZN(P2_U3243) );
  OAI21_X1 U16331 ( .B1(n14334), .B2(n14342), .A(n14333), .ZN(n14336) );
  AOI222_X1 U16332 ( .A1(n14358), .A2(n14336), .B1(n14370), .B2(n14368), .C1(
        n14335), .C2(n14369), .ZN(n14447) );
  AOI211_X1 U16333 ( .C1(n14338), .C2(n14348), .A(n12878), .B(n14337), .ZN(
        n14449) );
  INV_X1 U16334 ( .A(n14338), .ZN(n14504) );
  AOI22_X1 U16335 ( .A1(n14339), .A2(n15499), .B1(P2_REG2_REG_21__SCAN_IN), 
        .B2(n6677), .ZN(n14340) );
  OAI21_X1 U16336 ( .B1(n14504), .B2(n15503), .A(n14340), .ZN(n14341) );
  AOI21_X1 U16337 ( .B1(n14449), .B2(n15498), .A(n14341), .ZN(n14345) );
  XNOR2_X1 U16338 ( .A(n14343), .B(n14342), .ZN(n14450) );
  NAND2_X1 U16339 ( .A1(n14450), .A2(n15496), .ZN(n14344) );
  OAI211_X1 U16340 ( .C1(n14447), .C2(n6677), .A(n14345), .B(n14344), .ZN(
        P2_U3244) );
  XNOR2_X1 U16341 ( .A(n14346), .B(n14354), .ZN(n14457) );
  INV_X1 U16342 ( .A(n14348), .ZN(n14349) );
  AOI211_X1 U16343 ( .C1(n14454), .C2(n14374), .A(n12878), .B(n14349), .ZN(
        n14453) );
  AOI22_X1 U16344 ( .A1(n14350), .A2(n15499), .B1(n6677), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n14351) );
  OAI21_X1 U16345 ( .B1(n8712), .B2(n15503), .A(n14351), .ZN(n14360) );
  OAI21_X1 U16346 ( .B1(n14354), .B2(n14353), .A(n14352), .ZN(n14357) );
  AOI222_X1 U16347 ( .A1(n14358), .A2(n14357), .B1(n14356), .B2(n14368), .C1(
        n14355), .C2(n14369), .ZN(n14456) );
  NOR2_X1 U16348 ( .A1(n14456), .A2(n6677), .ZN(n14359) );
  AOI211_X1 U16349 ( .C1(n14453), .C2(n15498), .A(n14360), .B(n14359), .ZN(
        n14361) );
  OAI21_X1 U16350 ( .B1(n14457), .B2(n14362), .A(n14361), .ZN(P2_U3245) );
  XNOR2_X1 U16351 ( .A(n14363), .B(n14365), .ZN(n14460) );
  INV_X1 U16352 ( .A(n14460), .ZN(n14382) );
  AOI21_X1 U16353 ( .B1(n14365), .B2(n14364), .A(n6746), .ZN(n14373) );
  NAND2_X1 U16354 ( .A1(n14460), .A2(n14366), .ZN(n14372) );
  AOI22_X1 U16355 ( .A1(n14370), .A2(n14369), .B1(n14368), .B2(n14367), .ZN(
        n14371) );
  OAI211_X1 U16356 ( .C1(n14395), .C2(n14373), .A(n14372), .B(n14371), .ZN(
        n14458) );
  NAND2_X1 U16357 ( .A1(n14458), .A2(n14397), .ZN(n14380) );
  AOI211_X1 U16358 ( .C1(n14375), .C2(n14400), .A(n12878), .B(n14347), .ZN(
        n14459) );
  AOI22_X1 U16359 ( .A1(P2_REG2_REG_19__SCAN_IN), .A2(n6677), .B1(n14376), 
        .B2(n15499), .ZN(n14377) );
  OAI21_X1 U16360 ( .B1(n14509), .B2(n15503), .A(n14377), .ZN(n14378) );
  AOI21_X1 U16361 ( .B1(n14459), .B2(n15498), .A(n14378), .ZN(n14379) );
  OAI211_X1 U16362 ( .C1(n14382), .C2(n14381), .A(n14380), .B(n14379), .ZN(
        P2_U3246) );
  OAI21_X1 U16363 ( .B1(n14384), .B2(n14391), .A(n14383), .ZN(n14465) );
  NAND2_X1 U16364 ( .A1(n14465), .A2(n15496), .ZN(n14404) );
  NAND2_X1 U16365 ( .A1(n6677), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n14385) );
  OAI21_X1 U16366 ( .B1(n14387), .B2(n14386), .A(n14385), .ZN(n14388) );
  AOI21_X1 U16367 ( .B1(n14390), .B2(n14389), .A(n14388), .ZN(n14403) );
  XNOR2_X1 U16368 ( .A(n14392), .B(n14391), .ZN(n14396) );
  INV_X1 U16369 ( .A(n14393), .ZN(n14394) );
  OAI21_X1 U16370 ( .B1(n14396), .B2(n14395), .A(n14394), .ZN(n14463) );
  NAND2_X1 U16371 ( .A1(n14463), .A2(n14397), .ZN(n14402) );
  OR2_X1 U16372 ( .A1(n14513), .A2(n6800), .ZN(n14399) );
  AND3_X1 U16373 ( .A1(n14400), .A2(n14399), .A3(n14398), .ZN(n14464) );
  NAND2_X1 U16374 ( .A1(n14464), .A2(n15498), .ZN(n14401) );
  NAND4_X1 U16375 ( .A1(n14404), .A2(n14403), .A3(n14402), .A4(n14401), .ZN(
        P2_U3247) );
  NAND2_X1 U16376 ( .A1(n14405), .A2(n14409), .ZN(n14482) );
  MUX2_X1 U16377 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n14482), .S(n15550), .Z(
        n14406) );
  AOI21_X1 U16378 ( .B1(n14407), .B2(n14484), .A(n14406), .ZN(n14408) );
  INV_X1 U16379 ( .A(n14408), .ZN(P2_U3530) );
  INV_X1 U16380 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n14411) );
  AND2_X1 U16381 ( .A1(n14410), .A2(n14409), .ZN(n14486) );
  MUX2_X1 U16382 ( .A(n14411), .B(n14486), .S(n15550), .Z(n14412) );
  OAI21_X1 U16383 ( .B1(n14489), .B2(n14472), .A(n14412), .ZN(P2_U3529) );
  NAND3_X1 U16384 ( .A1(n14237), .A2(n15520), .A3(n14413), .ZN(n14418) );
  AOI21_X1 U16385 ( .B1(n15532), .B2(n14415), .A(n14414), .ZN(n14416) );
  NAND3_X1 U16386 ( .A1(n14418), .A2(n14417), .A3(n14416), .ZN(n14490) );
  MUX2_X1 U16387 ( .A(n14490), .B(P2_REG1_REG_27__SCAN_IN), .S(n15548), .Z(
        P2_U3526) );
  AOI21_X1 U16388 ( .B1(n15532), .B2(n14420), .A(n14419), .ZN(n14421) );
  OAI211_X1 U16389 ( .C1(n14423), .C2(n14478), .A(n14422), .B(n14421), .ZN(
        n14491) );
  MUX2_X1 U16390 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14491), .S(n15550), .Z(
        P2_U3525) );
  INV_X1 U16391 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n14426) );
  AOI211_X1 U16392 ( .C1(n15520), .C2(n14425), .A(n7603), .B(n14424), .ZN(
        n14492) );
  MUX2_X1 U16393 ( .A(n14426), .B(n14492), .S(n15550), .Z(n14427) );
  OAI21_X1 U16394 ( .B1(n14495), .B2(n14472), .A(n14427), .ZN(P2_U3524) );
  INV_X1 U16395 ( .A(n14428), .ZN(n14433) );
  AOI21_X1 U16396 ( .B1(n15532), .B2(n14430), .A(n14429), .ZN(n14431) );
  OAI211_X1 U16397 ( .C1(n14434), .C2(n14433), .A(n14432), .B(n14431), .ZN(
        n14496) );
  MUX2_X1 U16398 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14496), .S(n15550), .Z(
        P2_U3523) );
  INV_X1 U16399 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n14440) );
  NAND2_X1 U16400 ( .A1(n14435), .A2(n15520), .ZN(n14439) );
  NOR2_X1 U16401 ( .A1(n14437), .A2(n14436), .ZN(n14438) );
  MUX2_X1 U16402 ( .A(n14440), .B(n14497), .S(n15550), .Z(n14441) );
  OAI21_X1 U16403 ( .B1(n7227), .B2(n14472), .A(n14441), .ZN(P2_U3522) );
  AOI21_X1 U16404 ( .B1(n15532), .B2(n14443), .A(n14442), .ZN(n14444) );
  OAI211_X1 U16405 ( .C1(n14446), .C2(n14478), .A(n14445), .B(n14444), .ZN(
        n14500) );
  MUX2_X1 U16406 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n14500), .S(n15550), .Z(
        P2_U3521) );
  INV_X1 U16407 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n14451) );
  INV_X1 U16408 ( .A(n14447), .ZN(n14448) );
  AOI211_X1 U16409 ( .C1(n15520), .C2(n14450), .A(n14449), .B(n14448), .ZN(
        n14501) );
  MUX2_X1 U16410 ( .A(n14451), .B(n14501), .S(n15550), .Z(n14452) );
  OAI21_X1 U16411 ( .B1(n14504), .B2(n14472), .A(n14452), .ZN(P2_U3520) );
  AOI21_X1 U16412 ( .B1(n15532), .B2(n14454), .A(n14453), .ZN(n14455) );
  OAI211_X1 U16413 ( .C1(n14478), .C2(n14457), .A(n14456), .B(n14455), .ZN(
        n14505) );
  MUX2_X1 U16414 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14505), .S(n15550), .Z(
        P2_U3519) );
  AOI211_X1 U16415 ( .C1(n15537), .C2(n14460), .A(n14459), .B(n14458), .ZN(
        n14506) );
  MUX2_X1 U16416 ( .A(n14461), .B(n14506), .S(n15550), .Z(n14462) );
  OAI21_X1 U16417 ( .B1(n14509), .B2(n14472), .A(n14462), .ZN(P2_U3518) );
  AOI211_X1 U16418 ( .C1(n15520), .C2(n14465), .A(n14464), .B(n14463), .ZN(
        n14510) );
  MUX2_X1 U16419 ( .A(n15480), .B(n14510), .S(n15550), .Z(n14466) );
  OAI21_X1 U16420 ( .B1(n14513), .B2(n14472), .A(n14466), .ZN(P2_U3517) );
  AOI211_X1 U16421 ( .C1(n14469), .C2(n15520), .A(n14468), .B(n14467), .ZN(
        n14515) );
  MUX2_X1 U16422 ( .A(n14515), .B(n14470), .S(n15548), .Z(n14471) );
  OAI21_X1 U16423 ( .B1(n14518), .B2(n14472), .A(n14471), .ZN(P2_U3516) );
  AOI211_X1 U16424 ( .C1(n15532), .C2(n14475), .A(n14474), .B(n14473), .ZN(
        n14476) );
  OAI21_X1 U16425 ( .B1(n14478), .B2(n14477), .A(n14476), .ZN(n14519) );
  MUX2_X1 U16426 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14519), .S(n15550), .Z(
        P2_U3515) );
  OAI22_X1 U16427 ( .A1(n14479), .A2(n14478), .B1(n8711), .B2(n15525), .ZN(
        n14481) );
  OR2_X1 U16428 ( .A1(n14481), .A2(n14480), .ZN(n14520) );
  MUX2_X1 U16429 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n14520), .S(n15550), .Z(
        P2_U3514) );
  MUX2_X1 U16430 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n14482), .S(n15543), .Z(
        n14483) );
  AOI21_X1 U16431 ( .B1(n10162), .B2(n14484), .A(n14483), .ZN(n14485) );
  INV_X1 U16432 ( .A(n14485), .ZN(P2_U3498) );
  INV_X1 U16433 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n14487) );
  MUX2_X1 U16434 ( .A(n14487), .B(n14486), .S(n15543), .Z(n14488) );
  OAI21_X1 U16435 ( .B1(n14489), .B2(n14517), .A(n14488), .ZN(P2_U3497) );
  MUX2_X1 U16436 ( .A(n14490), .B(P2_REG0_REG_27__SCAN_IN), .S(n15541), .Z(
        P2_U3494) );
  MUX2_X1 U16437 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14491), .S(n15543), .Z(
        P2_U3493) );
  INV_X1 U16438 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n14493) );
  MUX2_X1 U16439 ( .A(n14493), .B(n14492), .S(n15543), .Z(n14494) );
  OAI21_X1 U16440 ( .B1(n14495), .B2(n14517), .A(n14494), .ZN(P2_U3492) );
  MUX2_X1 U16441 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14496), .S(n15543), .Z(
        P2_U3491) );
  INV_X1 U16442 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n14498) );
  MUX2_X1 U16443 ( .A(n14498), .B(n14497), .S(n15543), .Z(n14499) );
  OAI21_X1 U16444 ( .B1(n7227), .B2(n14517), .A(n14499), .ZN(P2_U3490) );
  MUX2_X1 U16445 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n14500), .S(n15543), .Z(
        P2_U3489) );
  INV_X1 U16446 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n14502) );
  MUX2_X1 U16447 ( .A(n14502), .B(n14501), .S(n15543), .Z(n14503) );
  OAI21_X1 U16448 ( .B1(n14504), .B2(n14517), .A(n14503), .ZN(P2_U3488) );
  MUX2_X1 U16449 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14505), .S(n15543), .Z(
        P2_U3487) );
  INV_X1 U16450 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n14507) );
  MUX2_X1 U16451 ( .A(n14507), .B(n14506), .S(n15543), .Z(n14508) );
  OAI21_X1 U16452 ( .B1(n14509), .B2(n14517), .A(n14508), .ZN(P2_U3486) );
  INV_X1 U16453 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n14511) );
  MUX2_X1 U16454 ( .A(n14511), .B(n14510), .S(n15543), .Z(n14512) );
  OAI21_X1 U16455 ( .B1(n14513), .B2(n14517), .A(n14512), .ZN(P2_U3484) );
  INV_X1 U16456 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n14514) );
  MUX2_X1 U16457 ( .A(n14515), .B(n14514), .S(n15541), .Z(n14516) );
  OAI21_X1 U16458 ( .B1(n14518), .B2(n14517), .A(n14516), .ZN(P2_U3481) );
  MUX2_X1 U16459 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n14519), .S(n15543), .Z(
        P2_U3478) );
  MUX2_X1 U16460 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n14520), .S(n15543), .Z(
        P2_U3475) );
  INV_X1 U16461 ( .A(n14521), .ZN(n14527) );
  NOR4_X1 U16462 ( .A1(n14523), .A2(P2_IR_REG_30__SCAN_IN), .A3(n14522), .A4(
        P2_U3088), .ZN(n14524) );
  AOI21_X1 U16463 ( .B1(n14525), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n14524), 
        .ZN(n14526) );
  OAI21_X1 U16464 ( .B1(n14527), .B2(n14531), .A(n14526), .ZN(P2_U3296) );
  OAI222_X1 U16465 ( .A1(n14531), .A2(n14530), .B1(P2_U3088), .B2(n14529), 
        .C1(n14528), .C2(n12959), .ZN(P2_U3298) );
  MUX2_X1 U16466 ( .A(n14532), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  AOI22_X1 U16467 ( .A1(n14587), .A2(n14643), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14535) );
  NAND2_X1 U16468 ( .A1(n14615), .A2(n14642), .ZN(n14534) );
  OAI211_X1 U16469 ( .C1(n15222), .C2(n14822), .A(n14535), .B(n14534), .ZN(
        n14536) );
  AOI21_X1 U16470 ( .B1(n14537), .B2(n15218), .A(n14536), .ZN(n14538) );
  XOR2_X1 U16471 ( .A(n14540), .B(n14539), .Z(n14545) );
  AND2_X1 U16472 ( .A1(n14898), .A2(n15224), .ZN(n15027) );
  AOI22_X1 U16473 ( .A1(n14587), .A2(n14888), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14542) );
  NAND2_X1 U16474 ( .A1(n14615), .A2(n14887), .ZN(n14541) );
  OAI211_X1 U16475 ( .C1(n15222), .C2(n14896), .A(n14542), .B(n14541), .ZN(
        n14543) );
  AOI21_X1 U16476 ( .B1(n15027), .B2(n14627), .A(n14543), .ZN(n14544) );
  OAI21_X1 U16477 ( .B1(n14545), .B2(n15212), .A(n14544), .ZN(P1_U3216) );
  AOI21_X1 U16478 ( .B1(n14546), .B2(n14547), .A(n15212), .ZN(n14549) );
  NAND2_X1 U16479 ( .A1(n14549), .A2(n14548), .ZN(n14554) );
  NAND2_X1 U16480 ( .A1(n14647), .A2(n14975), .ZN(n14551) );
  NAND2_X1 U16481 ( .A1(n14648), .A2(n14974), .ZN(n14550) );
  AND2_X1 U16482 ( .A1(n14551), .A2(n14550), .ZN(n15054) );
  NAND2_X1 U16483 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14767)
         );
  OAI21_X1 U16484 ( .B1(n15054), .B2(n14633), .A(n14767), .ZN(n14552) );
  AOI21_X1 U16485 ( .B1(n14961), .B2(n14636), .A(n14552), .ZN(n14553) );
  OAI211_X1 U16486 ( .C1(n7996), .C2(n15186), .A(n14554), .B(n14553), .ZN(
        P1_U3219) );
  INV_X1 U16487 ( .A(n14555), .ZN(n14556) );
  AOI21_X1 U16488 ( .B1(n14558), .B2(n14557), .A(n14556), .ZN(n14564) );
  NAND2_X1 U16489 ( .A1(n14647), .A2(n14974), .ZN(n14560) );
  NAND2_X1 U16490 ( .A1(n14888), .A2(n14975), .ZN(n14559) );
  NAND2_X1 U16491 ( .A1(n14560), .A2(n14559), .ZN(n14923) );
  AOI22_X1 U16492 ( .A1(n14923), .A2(n15183), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14561) );
  OAI21_X1 U16493 ( .B1(n14925), .B2(n15222), .A(n14561), .ZN(n14562) );
  AOI21_X1 U16494 ( .B1(n14928), .B2(n15218), .A(n14562), .ZN(n14563) );
  OAI21_X1 U16495 ( .B1(n14564), .B2(n15212), .A(n14563), .ZN(P1_U3223) );
  XOR2_X1 U16496 ( .A(n14566), .B(n14565), .Z(n14572) );
  NAND2_X1 U16497 ( .A1(n14887), .A2(n14974), .ZN(n14568) );
  NAND2_X1 U16498 ( .A1(n14643), .A2(n14975), .ZN(n14567) );
  NAND2_X1 U16499 ( .A1(n14568), .A2(n14567), .ZN(n15016) );
  AOI22_X1 U16500 ( .A1(n15183), .A2(n15016), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14569) );
  OAI21_X1 U16501 ( .B1(n14854), .B2(n15222), .A(n14569), .ZN(n14570) );
  AOI21_X1 U16502 ( .B1(n15017), .B2(n15218), .A(n14570), .ZN(n14571) );
  OAI21_X1 U16503 ( .B1(n14572), .B2(n15212), .A(n14571), .ZN(P1_U3225) );
  NAND2_X1 U16504 ( .A1(n14573), .A2(n15224), .ZN(n15064) );
  OAI21_X1 U16505 ( .B1(n14576), .B2(n14575), .A(n14574), .ZN(n14577) );
  NAND2_X1 U16506 ( .A1(n14577), .A2(n15179), .ZN(n14583) );
  AOI22_X1 U16507 ( .A1(n14615), .A2(n14648), .B1(P1_REG3_REG_17__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14578) );
  OAI21_X1 U16508 ( .B1(n14579), .B2(n15206), .A(n14578), .ZN(n14580) );
  AOI21_X1 U16509 ( .B1(n14581), .B2(n14636), .A(n14580), .ZN(n14582) );
  OAI211_X1 U16510 ( .C1(n14584), .C2(n15064), .A(n14583), .B(n14582), .ZN(
        P1_U3228) );
  XOR2_X1 U16511 ( .A(n14586), .B(n14585), .Z(n14592) );
  INV_X1 U16512 ( .A(n15224), .ZN(n15317) );
  NOR2_X1 U16513 ( .A1(n14880), .A2(n15317), .ZN(n15022) );
  AOI22_X1 U16514 ( .A1(n14587), .A2(n14645), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14589) );
  NAND2_X1 U16515 ( .A1(n14615), .A2(n14644), .ZN(n14588) );
  OAI211_X1 U16516 ( .C1(n15222), .C2(n14876), .A(n14589), .B(n14588), .ZN(
        n14590) );
  AOI21_X1 U16517 ( .B1(n15022), .B2(n14627), .A(n14590), .ZN(n14591) );
  OAI21_X1 U16518 ( .B1(n14592), .B2(n15212), .A(n14591), .ZN(P1_U3229) );
  OAI211_X1 U16519 ( .C1(n14595), .C2(n14594), .A(n14593), .B(n15179), .ZN(
        n14601) );
  OAI22_X1 U16520 ( .A1(n14597), .A2(n14869), .B1(n14596), .B2(n14871), .ZN(
        n14936) );
  AOI22_X1 U16521 ( .A1(n14936), .A2(n15183), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14598) );
  OAI21_X1 U16522 ( .B1(n14945), .B2(n15222), .A(n14598), .ZN(n14599) );
  AOI21_X1 U16523 ( .B1(n15048), .B2(n15218), .A(n14599), .ZN(n14600) );
  NAND2_X1 U16524 ( .A1(n14601), .A2(n14600), .ZN(P1_U3233) );
  OAI21_X1 U16525 ( .B1(n14604), .B2(n14603), .A(n14602), .ZN(n14605) );
  INV_X1 U16526 ( .A(n14605), .ZN(n14611) );
  NAND2_X1 U16527 ( .A1(n14646), .A2(n14974), .ZN(n14607) );
  NAND2_X1 U16528 ( .A1(n14645), .A2(n14975), .ZN(n14606) );
  NAND2_X1 U16529 ( .A1(n14607), .A2(n14606), .ZN(n15034) );
  AOI22_X1 U16530 ( .A1(n15183), .A2(n15034), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14608) );
  OAI21_X1 U16531 ( .B1(n14910), .B2(n15222), .A(n14608), .ZN(n14609) );
  AOI21_X1 U16532 ( .B1(n15035), .B2(n15218), .A(n14609), .ZN(n14610) );
  OAI21_X1 U16533 ( .B1(n14611), .B2(n15212), .A(n14610), .ZN(P1_U3235) );
  XOR2_X1 U16534 ( .A(n14613), .B(n14612), .Z(n14619) );
  NAND2_X1 U16535 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14738)
         );
  OAI21_X1 U16536 ( .B1(n15206), .B2(n15191), .A(n14738), .ZN(n14614) );
  AOI21_X1 U16537 ( .B1(n14615), .B2(n14976), .A(n14614), .ZN(n14616) );
  OAI21_X1 U16538 ( .B1(n14983), .B2(n15222), .A(n14616), .ZN(n14617) );
  AOI21_X1 U16539 ( .B1(n14991), .B2(n15218), .A(n14617), .ZN(n14618) );
  OAI21_X1 U16540 ( .B1(n14619), .B2(n15212), .A(n14618), .ZN(P1_U3238) );
  XOR2_X1 U16541 ( .A(n14621), .B(n14620), .Z(n14629) );
  AND2_X1 U16542 ( .A1(n14622), .A2(n15224), .ZN(n15010) );
  NAND2_X1 U16543 ( .A1(n14644), .A2(n14974), .ZN(n14624) );
  NAND2_X1 U16544 ( .A1(n14803), .A2(n14975), .ZN(n14623) );
  NAND2_X1 U16545 ( .A1(n14624), .A2(n14623), .ZN(n15009) );
  AOI22_X1 U16546 ( .A1(n15183), .A2(n15009), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14625) );
  OAI21_X1 U16547 ( .B1(n14837), .B2(n15222), .A(n14625), .ZN(n14626) );
  AOI21_X1 U16548 ( .B1(n15010), .B2(n14627), .A(n14626), .ZN(n14628) );
  OAI21_X1 U16549 ( .B1(n14629), .B2(n15212), .A(n14628), .ZN(P1_U3240) );
  OAI211_X1 U16550 ( .C1(n14632), .C2(n14631), .A(n14630), .B(n15179), .ZN(
        n14639) );
  NAND2_X1 U16551 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n15269)
         );
  OAI21_X1 U16552 ( .B1(n14634), .B2(n14633), .A(n15269), .ZN(n14635) );
  AOI21_X1 U16553 ( .B1(n14637), .B2(n14636), .A(n14635), .ZN(n14638) );
  OAI211_X1 U16554 ( .C1(n8211), .C2(n15186), .A(n14639), .B(n14638), .ZN(
        P1_U3241) );
  MUX2_X1 U16555 ( .A(n14773), .B(P1_DATAO_REG_31__SCAN_IN), .S(n14640), .Z(
        P1_U3591) );
  MUX2_X1 U16556 ( .A(n14641), .B(P1_DATAO_REG_30__SCAN_IN), .S(n14640), .Z(
        P1_U3590) );
  MUX2_X1 U16557 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14802), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16558 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14642), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16559 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14803), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16560 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14643), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16561 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14644), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16562 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14887), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16563 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14645), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16564 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14888), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16565 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14646), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16566 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14647), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16567 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14976), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U16568 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14648), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16569 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14973), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16570 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14649), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U16571 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14650), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16572 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14651), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16573 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14652), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U16574 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14653), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U16575 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14654), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U16576 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14655), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U16577 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14656), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U16578 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14657), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U16579 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14658), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U16580 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14659), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U16581 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14660), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U16582 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14661), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U16583 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14662), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U16584 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n14663), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U16585 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14664), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI22_X1 U16586 ( .A1(n15271), .A2(n9383), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14665), .ZN(n14666) );
  AOI21_X1 U16587 ( .B1(n14667), .B2(n15263), .A(n14666), .ZN(n14678) );
  AND2_X1 U16588 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n14669) );
  OAI211_X1 U16589 ( .C1(n14670), .C2(n14669), .A(n15260), .B(n14668), .ZN(
        n14677) );
  INV_X1 U16590 ( .A(n14671), .ZN(n14675) );
  MUX2_X1 U16591 ( .A(n14673), .B(P1_REG2_REG_1__SCAN_IN), .S(n14672), .Z(
        n14674) );
  OAI211_X1 U16592 ( .C1(n14675), .C2(n14674), .A(n14762), .B(n14685), .ZN(
        n14676) );
  NAND3_X1 U16593 ( .A1(n14678), .A2(n14677), .A3(n14676), .ZN(P1_U3244) );
  OAI22_X1 U16594 ( .A1(n15271), .A2(n9384), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14679), .ZN(n14680) );
  AOI21_X1 U16595 ( .B1(n14681), .B2(n15263), .A(n14680), .ZN(n14692) );
  INV_X1 U16596 ( .A(n14682), .ZN(n14687) );
  NAND3_X1 U16597 ( .A1(n14685), .A2(n14684), .A3(n14683), .ZN(n14686) );
  NAND3_X1 U16598 ( .A1(n14762), .A2(n14687), .A3(n14686), .ZN(n14691) );
  OAI211_X1 U16599 ( .C1(n14689), .C2(n14688), .A(n15260), .B(n7059), .ZN(
        n14690) );
  NAND4_X1 U16600 ( .A1(n14693), .A2(n14692), .A3(n14691), .A4(n14690), .ZN(
        P1_U3245) );
  NAND2_X1 U16601 ( .A1(n14707), .A2(n14696), .ZN(n14697) );
  NAND2_X1 U16602 ( .A1(n15259), .A2(n15258), .ZN(n15257) );
  NAND2_X1 U16603 ( .A1(n14697), .A2(n15257), .ZN(n14699) );
  XNOR2_X1 U16604 ( .A(n14716), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n14698) );
  NOR2_X1 U16605 ( .A1(n14699), .A2(n14698), .ZN(n14715) );
  AOI211_X1 U16606 ( .C1(n14699), .C2(n14698), .A(n14759), .B(n14715), .ZN(
        n14703) );
  NAND2_X1 U16607 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n15201)
         );
  INV_X1 U16608 ( .A(n15201), .ZN(n14700) );
  AOI21_X1 U16609 ( .B1(n14737), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n14700), 
        .ZN(n14701) );
  OAI21_X1 U16610 ( .B1(n14721), .B2(n14757), .A(n14701), .ZN(n14702) );
  NOR2_X1 U16611 ( .A1(n14703), .A2(n14702), .ZN(n14714) );
  OAI21_X1 U16612 ( .B1(n11763), .B2(n14705), .A(n14704), .ZN(n14706) );
  NOR2_X1 U16613 ( .A1(n15262), .A2(n14706), .ZN(n14708) );
  XOR2_X1 U16614 ( .A(n14707), .B(n14706), .Z(n15256) );
  NOR2_X1 U16615 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n15256), .ZN(n15255) );
  NOR2_X1 U16616 ( .A1(n14708), .A2(n15255), .ZN(n14712) );
  NAND2_X1 U16617 ( .A1(n14716), .A2(n14720), .ZN(n14709) );
  OAI21_X1 U16618 ( .B1(n14716), .B2(n14720), .A(n14709), .ZN(n14711) );
  NAND2_X1 U16619 ( .A1(n14721), .A2(n14720), .ZN(n14710) );
  OAI211_X1 U16620 ( .C1(n14721), .C2(n14720), .A(n14712), .B(n14710), .ZN(
        n14719) );
  OAI211_X1 U16621 ( .C1(n14712), .C2(n14711), .A(n14719), .B(n14762), .ZN(
        n14713) );
  NAND2_X1 U16622 ( .A1(n14714), .A2(n14713), .ZN(P1_U3259) );
  AOI21_X1 U16623 ( .B1(n14716), .B2(P1_REG1_REG_16__SCAN_IN), .A(n14715), 
        .ZN(n14718) );
  XNOR2_X1 U16624 ( .A(n14733), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n14717) );
  NOR2_X1 U16625 ( .A1(n14718), .A2(n14717), .ZN(n14732) );
  AOI211_X1 U16626 ( .C1(n14718), .C2(n14717), .A(n14759), .B(n14732), .ZN(
        n14731) );
  OAI21_X1 U16627 ( .B1(n14721), .B2(n14720), .A(n14719), .ZN(n14725) );
  NOR2_X1 U16628 ( .A1(n14736), .A2(n14722), .ZN(n14723) );
  AOI21_X1 U16629 ( .B1(n14722), .B2(n14736), .A(n14723), .ZN(n14724) );
  NAND2_X1 U16630 ( .A1(n14724), .A2(n14725), .ZN(n14735) );
  OAI211_X1 U16631 ( .C1(n14725), .C2(n14724), .A(n14735), .B(n14762), .ZN(
        n14729) );
  INV_X1 U16632 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n14726) );
  NOR2_X1 U16633 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14726), .ZN(n14727) );
  AOI21_X1 U16634 ( .B1(n14737), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n14727), 
        .ZN(n14728) );
  OAI211_X1 U16635 ( .C1(n14757), .C2(n14736), .A(n14729), .B(n14728), .ZN(
        n14730) );
  OR2_X1 U16636 ( .A1(n14731), .A2(n14730), .ZN(P1_U3260) );
  OAI21_X1 U16637 ( .B1(n14734), .B2(P1_REG1_REG_18__SCAN_IN), .A(n15260), 
        .ZN(n14744) );
  OAI21_X1 U16638 ( .B1(n14736), .B2(n14722), .A(n14735), .ZN(n14752) );
  XNOR2_X1 U16639 ( .A(n14752), .B(n14751), .ZN(n14749) );
  XNOR2_X1 U16640 ( .A(n14749), .B(P1_REG2_REG_18__SCAN_IN), .ZN(n14742) );
  NAND2_X1 U16641 ( .A1(n14737), .A2(P1_ADDR_REG_18__SCAN_IN), .ZN(n14739) );
  OAI211_X1 U16642 ( .C1(n14757), .C2(n14740), .A(n14739), .B(n14738), .ZN(
        n14741) );
  AOI21_X1 U16643 ( .B1(n14762), .B2(n14742), .A(n14741), .ZN(n14743) );
  OAI21_X1 U16644 ( .B1(n14744), .B2(n14746), .A(n14743), .ZN(P1_U3261) );
  NOR2_X1 U16645 ( .A1(n14746), .A2(n14745), .ZN(n14748) );
  INV_X1 U16646 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14747) );
  XOR2_X1 U16647 ( .A(n14748), .B(n14747), .Z(n14763) );
  INV_X1 U16648 ( .A(n14749), .ZN(n14750) );
  NAND2_X1 U16649 ( .A1(n14750), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n14754) );
  NAND2_X1 U16650 ( .A1(n14752), .A2(n14751), .ZN(n14753) );
  NAND2_X1 U16651 ( .A1(n14754), .A2(n14753), .ZN(n14755) );
  NAND2_X1 U16652 ( .A1(n14756), .A2(n14762), .ZN(n14758) );
  OAI211_X1 U16653 ( .C1(n14763), .C2(n14759), .A(n14758), .B(n14757), .ZN(
        n14760) );
  INV_X1 U16654 ( .A(n14760), .ZN(n14766) );
  AOI22_X1 U16655 ( .A1(n14763), .A2(n15260), .B1(n14762), .B2(n14761), .ZN(
        n14765) );
  OAI211_X1 U16656 ( .C1(n14769), .C2(n15271), .A(n14768), .B(n14767), .ZN(
        P1_U3262) );
  XNOR2_X1 U16657 ( .A(n14774), .B(n14777), .ZN(n14770) );
  INV_X1 U16658 ( .A(n14771), .ZN(n14772) );
  NAND2_X1 U16659 ( .A1(n14773), .A2(n14772), .ZN(n14999) );
  NOR2_X1 U16660 ( .A1(n14962), .A2(n14999), .ZN(n14780) );
  NOR2_X1 U16661 ( .A1(n15075), .A2(n14949), .ZN(n14775) );
  AOI211_X1 U16662 ( .C1(n14962), .C2(P1_REG2_REG_31__SCAN_IN), .A(n14780), 
        .B(n14775), .ZN(n14776) );
  OAI21_X1 U16663 ( .B1(n14988), .B2(n14994), .A(n14776), .ZN(P1_U3263) );
  OAI211_X1 U16664 ( .C1(n15079), .C2(n14778), .A(n15049), .B(n14777), .ZN(
        n15000) );
  NOR2_X1 U16665 ( .A1(n14913), .A2(n14779), .ZN(n14781) );
  AOI211_X1 U16666 ( .C1(n7145), .C2(n14992), .A(n14781), .B(n14780), .ZN(
        n14782) );
  OAI21_X1 U16667 ( .B1(n15000), .B2(n14988), .A(n14782), .ZN(P1_U3264) );
  NAND2_X1 U16668 ( .A1(n14783), .A2(n15279), .ZN(n14797) );
  INV_X1 U16669 ( .A(n14784), .ZN(n14787) );
  INV_X1 U16670 ( .A(n14785), .ZN(n14786) );
  AOI22_X1 U16671 ( .A1(n14788), .A2(n14787), .B1(n14786), .B2(n15277), .ZN(
        n14793) );
  NOR2_X1 U16672 ( .A1(n14913), .A2(n14789), .ZN(n14790) );
  AOI21_X1 U16673 ( .B1(n14791), .B2(n14913), .A(n14790), .ZN(n14792) );
  OAI211_X1 U16674 ( .C1(n7144), .C2(n14949), .A(n14793), .B(n14792), .ZN(
        n14794) );
  AOI21_X1 U16675 ( .B1(n14795), .B2(n14944), .A(n14794), .ZN(n14796) );
  OAI211_X1 U16676 ( .C1(n14798), .C2(n14969), .A(n14797), .B(n14796), .ZN(
        P1_U3356) );
  NAND2_X1 U16677 ( .A1(n14802), .A2(n14975), .ZN(n14805) );
  OAI21_X1 U16678 ( .B1(n6737), .B2(n14809), .A(n14808), .ZN(n15007) );
  INV_X1 U16679 ( .A(n15007), .ZN(n14819) );
  AOI21_X1 U16680 ( .B1(n14810), .B2(n15004), .A(n14958), .ZN(n14812) );
  NAND2_X1 U16681 ( .A1(n15003), .A2(n14944), .ZN(n14816) );
  INV_X1 U16682 ( .A(n14813), .ZN(n14814) );
  AOI22_X1 U16683 ( .A1(n14962), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n14814), 
        .B2(n15277), .ZN(n14815) );
  OAI211_X1 U16684 ( .C1(n14817), .C2(n14949), .A(n14816), .B(n14815), .ZN(
        n14818) );
  AOI21_X1 U16685 ( .B1(n14819), .B2(n15279), .A(n14818), .ZN(n14820) );
  OAI21_X1 U16686 ( .B1(n15006), .B2(n14962), .A(n14820), .ZN(P1_U3265) );
  NAND2_X1 U16687 ( .A1(n14821), .A2(n14944), .ZN(n14825) );
  INV_X1 U16688 ( .A(n14822), .ZN(n14823) );
  AOI22_X1 U16689 ( .A1(n14962), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n14823), 
        .B2(n15277), .ZN(n14824) );
  OAI211_X1 U16690 ( .C1(n14826), .C2(n14949), .A(n14825), .B(n14824), .ZN(
        n14827) );
  AOI21_X1 U16691 ( .B1(n14828), .B2(n14913), .A(n14827), .ZN(n14829) );
  INV_X1 U16692 ( .A(n14829), .ZN(P1_U3266) );
  XNOR2_X1 U16693 ( .A(n14830), .B(n14831), .ZN(n15008) );
  INV_X1 U16694 ( .A(n15008), .ZN(n14846) );
  OR2_X1 U16695 ( .A1(n14832), .A2(n14831), .ZN(n14833) );
  NAND2_X1 U16696 ( .A1(n14834), .A2(n14833), .ZN(n14835) );
  NAND2_X1 U16697 ( .A1(n14835), .A2(n6966), .ZN(n15012) );
  INV_X1 U16698 ( .A(n15009), .ZN(n14836) );
  OAI211_X1 U16699 ( .C1(n14837), .C2(n14982), .A(n15012), .B(n14836), .ZN(
        n14844) );
  OAI21_X1 U16700 ( .B1(n14853), .B2(n14841), .A(n15049), .ZN(n14838) );
  NOR2_X1 U16701 ( .A1(n15011), .A2(n14988), .ZN(n14843) );
  OAI22_X1 U16702 ( .A1(n14841), .A2(n14949), .B1(n14840), .B2(n14913), .ZN(
        n14842) );
  AOI211_X1 U16703 ( .C1(n14844), .C2(n14913), .A(n14843), .B(n14842), .ZN(
        n14845) );
  OAI21_X1 U16704 ( .B1(n14846), .B2(n14862), .A(n14845), .ZN(P1_U3267) );
  OAI21_X1 U16705 ( .B1(n14848), .B2(n8102), .A(n14847), .ZN(n15021) );
  OAI21_X1 U16706 ( .B1(n14851), .B2(n14850), .A(n14849), .ZN(n15018) );
  INV_X1 U16707 ( .A(n14852), .ZN(n14878) );
  AOI211_X1 U16708 ( .C1(n15017), .C2(n14878), .A(n14958), .B(n14853), .ZN(
        n15015) );
  NAND2_X1 U16709 ( .A1(n15015), .A2(n14944), .ZN(n14858) );
  OAI22_X1 U16710 ( .A1(n14913), .A2(n14855), .B1(n14854), .B2(n14982), .ZN(
        n14856) );
  AOI21_X1 U16711 ( .B1(n15016), .B2(n14913), .A(n14856), .ZN(n14857) );
  OAI211_X1 U16712 ( .C1(n14859), .C2(n14949), .A(n14858), .B(n14857), .ZN(
        n14860) );
  AOI21_X1 U16713 ( .B1(n15018), .B2(n15280), .A(n14860), .ZN(n14861) );
  OAI21_X1 U16714 ( .B1(n15021), .B2(n14862), .A(n14861), .ZN(P1_U3268) );
  OAI21_X1 U16715 ( .B1(n14866), .B2(n14864), .A(n14863), .ZN(n14875) );
  NAND3_X1 U16716 ( .A1(n14885), .A2(n14866), .A3(n14865), .ZN(n14867) );
  AOI21_X1 U16717 ( .B1(n14868), .B2(n14867), .A(n15286), .ZN(n14874) );
  OAI22_X1 U16718 ( .A1(n14872), .A2(n14871), .B1(n14870), .B2(n14869), .ZN(
        n14873) );
  AOI211_X1 U16719 ( .C1(n14875), .C2(n14980), .A(n14874), .B(n14873), .ZN(
        n15025) );
  OAI22_X1 U16720 ( .A1(n14913), .A2(n14877), .B1(n14876), .B2(n14982), .ZN(
        n14882) );
  INV_X1 U16721 ( .A(n14894), .ZN(n14879) );
  OAI211_X1 U16722 ( .C1(n14880), .C2(n14879), .A(n14878), .B(n15049), .ZN(
        n15023) );
  NOR2_X1 U16723 ( .A1(n15023), .A2(n14988), .ZN(n14881) );
  AOI211_X1 U16724 ( .C1(n14992), .C2(n14883), .A(n14882), .B(n14881), .ZN(
        n14884) );
  OAI21_X1 U16725 ( .B1(n15025), .B2(n14962), .A(n14884), .ZN(P1_U3269) );
  OAI21_X1 U16726 ( .B1(n14892), .B2(n14886), .A(n14885), .ZN(n14889) );
  AOI222_X1 U16727 ( .A1(n6966), .A2(n14889), .B1(n14888), .B2(n14974), .C1(
        n14887), .C2(n14975), .ZN(n15030) );
  AOI21_X1 U16728 ( .B1(n14892), .B2(n14891), .A(n14890), .ZN(n15026) );
  AOI21_X1 U16729 ( .B1(n14909), .B2(n14898), .A(n14958), .ZN(n14895) );
  NAND2_X1 U16730 ( .A1(n14895), .A2(n14894), .ZN(n15028) );
  INV_X1 U16731 ( .A(n14896), .ZN(n14897) );
  AOI22_X1 U16732 ( .A1(n14962), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n14897), 
        .B2(n15277), .ZN(n14900) );
  NAND2_X1 U16733 ( .A1(n14898), .A2(n14992), .ZN(n14899) );
  OAI211_X1 U16734 ( .C1(n15028), .C2(n14988), .A(n14900), .B(n14899), .ZN(
        n14901) );
  AOI21_X1 U16735 ( .B1(n15026), .B2(n15279), .A(n14901), .ZN(n14902) );
  OAI21_X1 U16736 ( .B1(n14962), .B2(n15030), .A(n14902), .ZN(P1_U3270) );
  INV_X1 U16737 ( .A(n14903), .ZN(n14904) );
  AOI21_X1 U16738 ( .B1(n14907), .B2(n14905), .A(n14904), .ZN(n15038) );
  OAI21_X1 U16739 ( .B1(n14908), .B2(n14907), .A(n14906), .ZN(n15032) );
  NAND2_X1 U16740 ( .A1(n15032), .A2(n15279), .ZN(n14918) );
  AOI211_X1 U16741 ( .C1(n15035), .C2(n14924), .A(n14958), .B(n14893), .ZN(
        n15033) );
  OAI22_X1 U16742 ( .A1(n14913), .A2(n14911), .B1(n14910), .B2(n14982), .ZN(
        n14912) );
  AOI21_X1 U16743 ( .B1(n14913), .B2(n15034), .A(n14912), .ZN(n14914) );
  OAI21_X1 U16744 ( .B1(n14915), .B2(n14949), .A(n14914), .ZN(n14916) );
  AOI21_X1 U16745 ( .B1(n15033), .B2(n14944), .A(n14916), .ZN(n14917) );
  OAI211_X1 U16746 ( .C1(n15038), .C2(n14969), .A(n14918), .B(n14917), .ZN(
        P1_U3271) );
  XNOR2_X1 U16747 ( .A(n14919), .B(n14920), .ZN(n15043) );
  XNOR2_X1 U16748 ( .A(n14921), .B(n14920), .ZN(n14922) );
  NAND2_X1 U16749 ( .A1(n14922), .A2(n6966), .ZN(n15041) );
  INV_X1 U16750 ( .A(n14923), .ZN(n15040) );
  AOI21_X1 U16751 ( .B1(n15041), .B2(n15040), .A(n14962), .ZN(n14931) );
  OAI211_X1 U16752 ( .C1(n14943), .C2(n15090), .A(n14924), .B(n15049), .ZN(
        n15039) );
  OAI22_X1 U16753 ( .A1(n14913), .A2(n14926), .B1(n14925), .B2(n14982), .ZN(
        n14927) );
  AOI21_X1 U16754 ( .B1(n14928), .B2(n14992), .A(n14927), .ZN(n14929) );
  OAI21_X1 U16755 ( .B1(n15039), .B2(n14988), .A(n14929), .ZN(n14930) );
  AOI211_X1 U16756 ( .C1(n15043), .C2(n15279), .A(n14931), .B(n14930), .ZN(
        n14932) );
  INV_X1 U16757 ( .A(n14932), .ZN(P1_U3272) );
  INV_X1 U16758 ( .A(n14933), .ZN(n14935) );
  AOI21_X1 U16759 ( .B1(n14935), .B2(n14934), .A(n15286), .ZN(n14938) );
  AOI21_X1 U16760 ( .B1(n14938), .B2(n14937), .A(n14936), .ZN(n15052) );
  AOI21_X1 U16761 ( .B1(n14941), .B2(n14940), .A(n14939), .ZN(n15047) );
  INV_X1 U16762 ( .A(n15048), .ZN(n14950) );
  AND2_X1 U16763 ( .A1(n14959), .A2(n15048), .ZN(n14942) );
  NOR2_X1 U16764 ( .A1(n14943), .A2(n14942), .ZN(n15050) );
  NAND3_X1 U16765 ( .A1(n15050), .A2(n15049), .A3(n14944), .ZN(n14948) );
  INV_X1 U16766 ( .A(n14945), .ZN(n14946) );
  AOI22_X1 U16767 ( .A1(n14962), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n14946), 
        .B2(n15277), .ZN(n14947) );
  OAI211_X1 U16768 ( .C1(n14950), .C2(n14949), .A(n14948), .B(n14947), .ZN(
        n14951) );
  AOI21_X1 U16769 ( .B1(n15047), .B2(n15279), .A(n14951), .ZN(n14952) );
  OAI21_X1 U16770 ( .B1(n14962), .B2(n15052), .A(n14952), .ZN(P1_U3273) );
  XNOR2_X1 U16771 ( .A(n14954), .B(n14953), .ZN(n15059) );
  OAI21_X1 U16772 ( .B1(n14957), .B2(n14956), .A(n14955), .ZN(n15057) );
  AOI21_X1 U16773 ( .B1(n14986), .B2(n14965), .A(n14958), .ZN(n14960) );
  NAND2_X1 U16774 ( .A1(n14960), .A2(n14959), .ZN(n15055) );
  AOI22_X1 U16775 ( .A1(n14962), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n14961), 
        .B2(n15277), .ZN(n14963) );
  OAI21_X1 U16776 ( .B1(n15054), .B2(n14962), .A(n14963), .ZN(n14964) );
  AOI21_X1 U16777 ( .B1(n14965), .B2(n14992), .A(n14964), .ZN(n14966) );
  OAI21_X1 U16778 ( .B1(n15055), .B2(n14988), .A(n14966), .ZN(n14967) );
  AOI21_X1 U16779 ( .B1(n15057), .B2(n15279), .A(n14967), .ZN(n14968) );
  OAI21_X1 U16780 ( .B1(n15059), .B2(n14969), .A(n14968), .ZN(P1_U3274) );
  XNOR2_X1 U16781 ( .A(n14970), .B(n14972), .ZN(n14981) );
  XNOR2_X1 U16782 ( .A(n14971), .B(n14972), .ZN(n14978) );
  AOI22_X1 U16783 ( .A1(n14976), .A2(n14975), .B1(n14974), .B2(n14973), .ZN(
        n14977) );
  OAI21_X1 U16784 ( .B1(n14978), .B2(n15286), .A(n14977), .ZN(n14979) );
  AOI21_X1 U16785 ( .B1(n14981), .B2(n14980), .A(n14979), .ZN(n15061) );
  INV_X1 U16786 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14984) );
  OAI22_X1 U16787 ( .A1(n14913), .A2(n14984), .B1(n14983), .B2(n14982), .ZN(
        n14990) );
  INV_X1 U16788 ( .A(n14985), .ZN(n14987) );
  OAI211_X1 U16789 ( .C1(n7137), .C2(n14987), .A(n14986), .B(n15049), .ZN(
        n15060) );
  NOR2_X1 U16790 ( .A1(n15060), .A2(n14988), .ZN(n14989) );
  AOI211_X1 U16791 ( .C1(n14992), .C2(n14991), .A(n14990), .B(n14989), .ZN(
        n14993) );
  OAI21_X1 U16792 ( .B1(n15061), .B2(n14962), .A(n14993), .ZN(P1_U3275) );
  OR2_X1 U16793 ( .A1(n15073), .A2(n15330), .ZN(n14997) );
  INV_X1 U16794 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n14995) );
  NAND2_X1 U16795 ( .A1(n15330), .A2(n14995), .ZN(n14996) );
  NAND2_X1 U16796 ( .A1(n14997), .A2(n14996), .ZN(n14998) );
  OAI21_X1 U16797 ( .B1(n15075), .B2(n15046), .A(n14998), .ZN(P1_U3559) );
  AND2_X1 U16798 ( .A1(n15000), .A2(n14999), .ZN(n15076) );
  MUX2_X1 U16799 ( .A(n15001), .B(n15076), .S(n15332), .Z(n15002) );
  OAI21_X1 U16800 ( .B1(n15079), .B2(n15046), .A(n15002), .ZN(P1_U3558) );
  INV_X1 U16801 ( .A(n15321), .ZN(n15287) );
  AOI21_X1 U16802 ( .B1(n15224), .B2(n15004), .A(n15003), .ZN(n15005) );
  OAI211_X1 U16803 ( .C1(n15007), .C2(n15287), .A(n15006), .B(n15005), .ZN(
        n15080) );
  MUX2_X1 U16804 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n15080), .S(n15332), .Z(
        P1_U3556) );
  NAND2_X1 U16805 ( .A1(n15008), .A2(n15321), .ZN(n15014) );
  NOR2_X1 U16806 ( .A1(n15010), .A2(n15009), .ZN(n15013) );
  NAND4_X1 U16807 ( .A1(n15014), .A2(n15013), .A3(n15012), .A4(n15011), .ZN(
        n15081) );
  MUX2_X1 U16808 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15081), .S(n15332), .Z(
        P1_U3554) );
  AOI211_X1 U16809 ( .C1(n15224), .C2(n15017), .A(n15016), .B(n15015), .ZN(
        n15020) );
  NAND2_X1 U16810 ( .A1(n15018), .A2(n6966), .ZN(n15019) );
  OAI211_X1 U16811 ( .C1(n15021), .C2(n15287), .A(n15020), .B(n15019), .ZN(
        n15082) );
  MUX2_X1 U16812 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n15082), .S(n15332), .Z(
        P1_U3553) );
  INV_X1 U16813 ( .A(n15022), .ZN(n15024) );
  NAND3_X1 U16814 ( .A1(n15025), .A2(n15024), .A3(n15023), .ZN(n15083) );
  MUX2_X1 U16815 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n15083), .S(n15332), .Z(
        P1_U3552) );
  NAND2_X1 U16816 ( .A1(n15026), .A2(n15321), .ZN(n15031) );
  INV_X1 U16817 ( .A(n15027), .ZN(n15029) );
  NAND4_X1 U16818 ( .A1(n15031), .A2(n15030), .A3(n15029), .A4(n15028), .ZN(
        n15084) );
  MUX2_X1 U16819 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15084), .S(n15332), .Z(
        P1_U3551) );
  NAND2_X1 U16820 ( .A1(n15032), .A2(n15321), .ZN(n15037) );
  AOI211_X1 U16821 ( .C1(n15224), .C2(n15035), .A(n15034), .B(n15033), .ZN(
        n15036) );
  OAI211_X1 U16822 ( .C1(n15286), .C2(n15038), .A(n15037), .B(n15036), .ZN(
        n15085) );
  MUX2_X1 U16823 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15085), .S(n15332), .Z(
        P1_U3550) );
  INV_X1 U16824 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n15044) );
  NAND3_X1 U16825 ( .A1(n15041), .A2(n15040), .A3(n15039), .ZN(n15042) );
  AOI21_X1 U16826 ( .B1(n15043), .B2(n15321), .A(n15042), .ZN(n15086) );
  MUX2_X1 U16827 ( .A(n15044), .B(n15086), .S(n15332), .Z(n15045) );
  OAI21_X1 U16828 ( .B1(n15090), .B2(n15046), .A(n15045), .ZN(P1_U3549) );
  INV_X1 U16829 ( .A(n15047), .ZN(n15053) );
  AOI22_X1 U16830 ( .A1(n15050), .A2(n15049), .B1(n15224), .B2(n15048), .ZN(
        n15051) );
  OAI211_X1 U16831 ( .C1(n15053), .C2(n15287), .A(n15052), .B(n15051), .ZN(
        n15091) );
  MUX2_X1 U16832 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n15091), .S(n15332), .Z(
        P1_U3548) );
  OAI211_X1 U16833 ( .C1(n7996), .C2(n15317), .A(n15055), .B(n15054), .ZN(
        n15056) );
  AOI21_X1 U16834 ( .B1(n15057), .B2(n15321), .A(n15056), .ZN(n15058) );
  OAI21_X1 U16835 ( .B1(n15286), .B2(n15059), .A(n15058), .ZN(n15092) );
  MUX2_X1 U16836 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15092), .S(n15332), .Z(
        P1_U3547) );
  OAI211_X1 U16837 ( .C1(n7137), .C2(n15317), .A(n15061), .B(n15060), .ZN(
        n15093) );
  MUX2_X1 U16838 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15093), .S(n15332), .Z(
        P1_U3546) );
  NAND2_X1 U16839 ( .A1(n15062), .A2(n15321), .ZN(n15066) );
  NAND4_X1 U16840 ( .A1(n15066), .A2(n15065), .A3(n15064), .A4(n15063), .ZN(
        n15094) );
  MUX2_X1 U16841 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15094), .S(n15332), .Z(
        P1_U3545) );
  NAND2_X1 U16842 ( .A1(n15067), .A2(n15321), .ZN(n15071) );
  AOI211_X1 U16843 ( .C1(n15224), .C2(n15200), .A(n15069), .B(n15068), .ZN(
        n15070) );
  OAI211_X1 U16844 ( .C1(n15286), .C2(n15072), .A(n15071), .B(n15070), .ZN(
        n15095) );
  MUX2_X1 U16845 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15095), .S(n15332), .Z(
        P1_U3544) );
  OAI21_X1 U16846 ( .B1(n15075), .B2(n15089), .A(n15074), .ZN(P1_U3527) );
  MUX2_X1 U16847 ( .A(n15077), .B(n15076), .S(n15324), .Z(n15078) );
  OAI21_X1 U16848 ( .B1(n15079), .B2(n15089), .A(n15078), .ZN(P1_U3526) );
  MUX2_X1 U16849 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n15080), .S(n15324), .Z(
        P1_U3524) );
  MUX2_X1 U16850 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15081), .S(n15324), .Z(
        P1_U3522) );
  MUX2_X1 U16851 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n15082), .S(n15324), .Z(
        P1_U3521) );
  MUX2_X1 U16852 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n15083), .S(n15324), .Z(
        P1_U3520) );
  MUX2_X1 U16853 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15084), .S(n15324), .Z(
        P1_U3519) );
  MUX2_X1 U16854 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15085), .S(n15324), .Z(
        P1_U3518) );
  MUX2_X1 U16855 ( .A(n15087), .B(n15086), .S(n15324), .Z(n15088) );
  OAI21_X1 U16856 ( .B1(n15090), .B2(n15089), .A(n15088), .ZN(P1_U3517) );
  MUX2_X1 U16857 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n15091), .S(n15324), .Z(
        P1_U3516) );
  MUX2_X1 U16858 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15092), .S(n15324), .Z(
        P1_U3515) );
  MUX2_X1 U16859 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15093), .S(n15324), .Z(
        P1_U3513) );
  MUX2_X1 U16860 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15094), .S(n15324), .Z(
        P1_U3510) );
  MUX2_X1 U16861 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15095), .S(n15324), .Z(
        P1_U3507) );
  MUX2_X1 U16862 ( .A(n15097), .B(n15096), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U16863 ( .A(n15098), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16864 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n15494) );
  AOI21_X1 U16865 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n15101) );
  OAI21_X1 U16866 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n15101), 
        .ZN(U28) );
  AOI21_X1 U16867 ( .B1(n15104), .B2(n15103), .A(n15102), .ZN(n15105) );
  XOR2_X1 U16868 ( .A(n15105), .B(P2_ADDR_REG_2__SCAN_IN), .Z(SUB_1596_U61) );
  OAI21_X1 U16869 ( .B1(n15107), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n15106), .ZN(
        n15108) );
  XOR2_X1 U16870 ( .A(n15109), .B(n15108), .Z(SUB_1596_U57) );
  INV_X1 U16871 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n15423) );
  XOR2_X1 U16872 ( .A(n15423), .B(n15110), .Z(SUB_1596_U55) );
  XOR2_X1 U16873 ( .A(n15111), .B(P2_ADDR_REG_9__SCAN_IN), .Z(SUB_1596_U54) );
  AOI21_X1 U16874 ( .B1(n15114), .B2(n15113), .A(n15112), .ZN(n15115) );
  XOR2_X1 U16875 ( .A(n15115), .B(P2_ADDR_REG_10__SCAN_IN), .Z(SUB_1596_U70)
         );
  OAI21_X1 U16876 ( .B1(n15117), .B2(n15317), .A(n15116), .ZN(n15119) );
  NOR2_X1 U16877 ( .A1(n15119), .A2(n15118), .ZN(n15121) );
  INV_X1 U16878 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n15120) );
  AOI22_X1 U16879 ( .A1(n15324), .A2(n15121), .B1(n15120), .B2(n10226), .ZN(
        P1_U3495) );
  AOI22_X1 U16880 ( .A1(n15332), .A2(n15121), .B1(n11713), .B2(n15330), .ZN(
        P1_U3540) );
  INV_X1 U16881 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n15474) );
  NOR2_X1 U16882 ( .A1(n15123), .A2(n15122), .ZN(n15124) );
  XNOR2_X1 U16883 ( .A(n15474), .B(n15124), .ZN(SUB_1596_U63) );
  AOI21_X1 U16884 ( .B1(n15127), .B2(n15126), .A(n15125), .ZN(n15141) );
  OAI21_X1 U16885 ( .B1(n15129), .B2(P3_REG1_REG_17__SCAN_IN), .A(n15128), 
        .ZN(n15139) );
  NAND2_X1 U16886 ( .A1(n15600), .A2(n15130), .ZN(n15132) );
  OAI211_X1 U16887 ( .C1(n15133), .C2(n15591), .A(n15132), .B(n15131), .ZN(
        n15138) );
  AOI211_X1 U16888 ( .C1(n15136), .C2(n15135), .A(n15595), .B(n15134), .ZN(
        n15137) );
  AOI211_X1 U16889 ( .C1(n15677), .C2(n15139), .A(n15138), .B(n15137), .ZN(
        n15140) );
  OAI21_X1 U16890 ( .B1(n15141), .B2(n15681), .A(n15140), .ZN(P3_U3199) );
  OAI22_X1 U16891 ( .A1(n15143), .A2(n15726), .B1(n15142), .B2(n15719), .ZN(
        n15144) );
  NOR2_X1 U16892 ( .A1(n15145), .A2(n15144), .ZN(n15155) );
  AOI22_X1 U16893 ( .A1(n15741), .A2(n15155), .B1(n9016), .B2(n15739), .ZN(
        P3_U3472) );
  NOR2_X1 U16894 ( .A1(n15146), .A2(n15719), .ZN(n15148) );
  AOI211_X1 U16895 ( .C1(n15724), .C2(n15149), .A(n15148), .B(n15147), .ZN(
        n15157) );
  AOI22_X1 U16896 ( .A1(n15741), .A2(n15157), .B1(n8989), .B2(n15739), .ZN(
        P3_U3471) );
  OAI22_X1 U16897 ( .A1(n15151), .A2(n15726), .B1(n15150), .B2(n15719), .ZN(
        n15152) );
  NOR2_X1 U16898 ( .A1(n15153), .A2(n15152), .ZN(n15159) );
  AOI22_X1 U16899 ( .A1(n15741), .A2(n15159), .B1(n8972), .B2(n15739), .ZN(
        P3_U3470) );
  INV_X1 U16900 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n15154) );
  AOI22_X1 U16901 ( .A1(n15734), .A2(n15155), .B1(n15154), .B2(n15732), .ZN(
        P3_U3429) );
  INV_X1 U16902 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n15156) );
  AOI22_X1 U16903 ( .A1(n15734), .A2(n15157), .B1(n15156), .B2(n15732), .ZN(
        P3_U3426) );
  INV_X1 U16904 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n15158) );
  AOI22_X1 U16905 ( .A1(n15734), .A2(n15159), .B1(n15158), .B2(n15732), .ZN(
        P3_U3423) );
  OAI21_X1 U16906 ( .B1(n15161), .B2(n15525), .A(n15160), .ZN(n15163) );
  AOI211_X1 U16907 ( .C1(n15537), .C2(n15164), .A(n15163), .B(n15162), .ZN(
        n15167) );
  AOI22_X1 U16908 ( .A1(n15550), .A2(n15167), .B1(n15165), .B2(n15548), .ZN(
        P2_U3511) );
  INV_X1 U16909 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n15166) );
  AOI22_X1 U16910 ( .A1(n15543), .A2(n15167), .B1(n15166), .B2(n15541), .ZN(
        P2_U3466) );
  OAI22_X1 U16911 ( .A1(n15168), .A2(n15206), .B1(n15205), .B2(n15192), .ZN(
        n15175) );
  INV_X1 U16912 ( .A(n13005), .ZN(n15171) );
  OAI21_X1 U16913 ( .B1(n15171), .B2(n15170), .A(n15169), .ZN(n15173) );
  AOI21_X1 U16914 ( .B1(n15173), .B2(n15172), .A(n15212), .ZN(n15174) );
  AOI211_X1 U16915 ( .C1(n15218), .C2(n15225), .A(n15175), .B(n15174), .ZN(
        n15177) );
  OAI211_X1 U16916 ( .C1(n15222), .C2(n15178), .A(n15177), .B(n15176), .ZN(
        P1_U3215) );
  OAI211_X1 U16917 ( .C1(n15181), .C2(n15180), .A(n15210), .B(n15179), .ZN(
        n15185) );
  AOI22_X1 U16918 ( .A1(n15183), .A2(n15182), .B1(P1_REG3_REG_10__SCAN_IN), 
        .B2(P1_U3086), .ZN(n15184) );
  OAI211_X1 U16919 ( .C1(n15187), .C2(n15186), .A(n15185), .B(n15184), .ZN(
        n15188) );
  INV_X1 U16920 ( .A(n15188), .ZN(n15189) );
  OAI21_X1 U16921 ( .B1(n15190), .B2(n15222), .A(n15189), .ZN(P1_U3217) );
  OAI22_X1 U16922 ( .A1(n15192), .A2(n15206), .B1(n15205), .B2(n15191), .ZN(
        n15199) );
  INV_X1 U16923 ( .A(n14630), .ZN(n15195) );
  OAI21_X1 U16924 ( .B1(n15195), .B2(n15194), .A(n15193), .ZN(n15197) );
  AOI21_X1 U16925 ( .B1(n15197), .B2(n15196), .A(n15212), .ZN(n15198) );
  AOI211_X1 U16926 ( .C1(n15218), .C2(n15200), .A(n15199), .B(n15198), .ZN(
        n15202) );
  OAI211_X1 U16927 ( .C1(n15222), .C2(n15203), .A(n15202), .B(n15201), .ZN(
        P1_U3226) );
  OAI22_X1 U16928 ( .A1(n15207), .A2(n15206), .B1(n15205), .B2(n15204), .ZN(
        n15216) );
  AOI21_X1 U16929 ( .B1(n15210), .B2(n15209), .A(n15208), .ZN(n15211) );
  INV_X1 U16930 ( .A(n15211), .ZN(n15214) );
  AOI21_X1 U16931 ( .B1(n15214), .B2(n15213), .A(n15212), .ZN(n15215) );
  AOI211_X1 U16932 ( .C1(n15218), .C2(n15217), .A(n15216), .B(n15215), .ZN(
        n15220) );
  OAI211_X1 U16933 ( .C1(n15222), .C2(n15221), .A(n15220), .B(n15219), .ZN(
        P1_U3236) );
  AOI21_X1 U16934 ( .B1(n15225), .B2(n15224), .A(n15223), .ZN(n15227) );
  OAI211_X1 U16935 ( .C1(n15228), .C2(n15287), .A(n15227), .B(n15226), .ZN(
        n15229) );
  AOI21_X1 U16936 ( .B1(n6966), .B2(n15230), .A(n15229), .ZN(n15232) );
  AOI22_X1 U16937 ( .A1(n15332), .A2(n15232), .B1(n7914), .B2(n15330), .ZN(
        P1_U3542) );
  INV_X1 U16938 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n15231) );
  AOI22_X1 U16939 ( .A1(n15324), .A2(n15232), .B1(n15231), .B2(n10226), .ZN(
        P1_U3501) );
  NOR2_X1 U16940 ( .A1(n15234), .A2(n15233), .ZN(n15235) );
  XOR2_X1 U16941 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n15235), .Z(SUB_1596_U69)
         );
  AOI21_X1 U16942 ( .B1(n15238), .B2(n15237), .A(n15236), .ZN(n15239) );
  XOR2_X1 U16943 ( .A(n15239), .B(P2_ADDR_REG_12__SCAN_IN), .Z(SUB_1596_U68)
         );
  NOR2_X1 U16944 ( .A1(n15241), .A2(n15240), .ZN(n15242) );
  XOR2_X1 U16945 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(n15242), .Z(SUB_1596_U67)
         );
  AOI21_X1 U16946 ( .B1(n15245), .B2(n15244), .A(n15243), .ZN(n15246) );
  XOR2_X1 U16947 ( .A(n15246), .B(P2_ADDR_REG_14__SCAN_IN), .Z(SUB_1596_U66)
         );
  OAI21_X1 U16948 ( .B1(n15249), .B2(n15248), .A(n15247), .ZN(n15250) );
  XOR2_X1 U16949 ( .A(n15250), .B(n15448), .Z(SUB_1596_U65) );
  OAI21_X1 U16950 ( .B1(n15253), .B2(n15252), .A(n15251), .ZN(n15254) );
  XOR2_X1 U16951 ( .A(n15254), .B(n15460), .Z(SUB_1596_U64) );
  AOI21_X1 U16952 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n15256), .A(n15255), 
        .ZN(n15267) );
  OAI21_X1 U16953 ( .B1(n15259), .B2(n15258), .A(n15257), .ZN(n15261) );
  NAND2_X1 U16954 ( .A1(n15261), .A2(n15260), .ZN(n15265) );
  NAND2_X1 U16955 ( .A1(n15263), .A2(n15262), .ZN(n15264) );
  OAI211_X1 U16956 ( .C1(n15267), .C2(n15266), .A(n15265), .B(n15264), .ZN(
        n15268) );
  INV_X1 U16957 ( .A(n15268), .ZN(n15270) );
  OAI211_X1 U16958 ( .C1(n15272), .C2(n15271), .A(n15270), .B(n15269), .ZN(
        P1_U3258) );
  NOR2_X1 U16959 ( .A1(n15274), .A2(n15273), .ZN(n15288) );
  NAND2_X1 U16960 ( .A1(n8213), .A2(n15275), .ZN(n15276) );
  AOI21_X1 U16961 ( .B1(n15288), .B2(n15276), .A(n15289), .ZN(n15283) );
  AOI22_X1 U16962 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n15277), .B1(
        P1_REG2_REG_0__SCAN_IN), .B2(n14962), .ZN(n15282) );
  INV_X1 U16963 ( .A(n15285), .ZN(n15278) );
  OAI21_X1 U16964 ( .B1(n15280), .B2(n15279), .A(n15278), .ZN(n15281) );
  OAI211_X1 U16965 ( .C1(n14962), .C2(n15283), .A(n15282), .B(n15281), .ZN(
        P1_U3293) );
  AND2_X1 U16966 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15284), .ZN(P1_U3294) );
  AND2_X1 U16967 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15284), .ZN(P1_U3295) );
  AND2_X1 U16968 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15284), .ZN(P1_U3296) );
  AND2_X1 U16969 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15284), .ZN(P1_U3297) );
  AND2_X1 U16970 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15284), .ZN(P1_U3298) );
  AND2_X1 U16971 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15284), .ZN(P1_U3299) );
  AND2_X1 U16972 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15284), .ZN(P1_U3300) );
  AND2_X1 U16973 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15284), .ZN(P1_U3301) );
  AND2_X1 U16974 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15284), .ZN(P1_U3302) );
  AND2_X1 U16975 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15284), .ZN(P1_U3303) );
  AND2_X1 U16976 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15284), .ZN(P1_U3304) );
  AND2_X1 U16977 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15284), .ZN(P1_U3305) );
  AND2_X1 U16978 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15284), .ZN(P1_U3306) );
  AND2_X1 U16979 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15284), .ZN(P1_U3307) );
  AND2_X1 U16980 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15284), .ZN(P1_U3308) );
  AND2_X1 U16981 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15284), .ZN(P1_U3309) );
  AND2_X1 U16982 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15284), .ZN(P1_U3310) );
  AND2_X1 U16983 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15284), .ZN(P1_U3311) );
  AND2_X1 U16984 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15284), .ZN(P1_U3312) );
  AND2_X1 U16985 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15284), .ZN(P1_U3313) );
  AND2_X1 U16986 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15284), .ZN(P1_U3314) );
  AND2_X1 U16987 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15284), .ZN(P1_U3315) );
  AND2_X1 U16988 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15284), .ZN(P1_U3316) );
  AND2_X1 U16989 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15284), .ZN(P1_U3317) );
  AND2_X1 U16990 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15284), .ZN(P1_U3318) );
  AND2_X1 U16991 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15284), .ZN(P1_U3319) );
  AND2_X1 U16992 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15284), .ZN(P1_U3320) );
  AND2_X1 U16993 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15284), .ZN(P1_U3321) );
  AND2_X1 U16994 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15284), .ZN(P1_U3322) );
  AND2_X1 U16995 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15284), .ZN(P1_U3323) );
  AOI21_X1 U16996 ( .B1(n15287), .B2(n15286), .A(n15285), .ZN(n15290) );
  NOR3_X1 U16997 ( .A1(n15290), .A2(n15289), .A3(n15288), .ZN(n15325) );
  INV_X1 U16998 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n15291) );
  AOI22_X1 U16999 ( .A1(n15324), .A2(n15325), .B1(n15291), .B2(n10226), .ZN(
        P1_U3459) );
  INV_X1 U17000 ( .A(n15292), .ZN(n15293) );
  OAI211_X1 U17001 ( .C1(n15295), .C2(n15317), .A(n15294), .B(n15293), .ZN(
        n15297) );
  AOI211_X1 U17002 ( .C1(n15321), .C2(n15298), .A(n15297), .B(n15296), .ZN(
        n15326) );
  INV_X1 U17003 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n15299) );
  AOI22_X1 U17004 ( .A1(n15324), .A2(n15326), .B1(n15299), .B2(n10226), .ZN(
        P1_U3462) );
  OAI21_X1 U17005 ( .B1(n15301), .B2(n15317), .A(n15300), .ZN(n15303) );
  AOI211_X1 U17006 ( .C1(n15321), .C2(n15304), .A(n15303), .B(n15302), .ZN(
        n15327) );
  INV_X1 U17007 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n15305) );
  AOI22_X1 U17008 ( .A1(n15324), .A2(n15327), .B1(n15305), .B2(n10226), .ZN(
        P1_U3465) );
  NAND3_X1 U17009 ( .A1(n15308), .A2(n15307), .A3(n15306), .ZN(n15309) );
  AOI211_X1 U17010 ( .C1(n15311), .C2(n15321), .A(n15310), .B(n15309), .ZN(
        n15328) );
  AOI22_X1 U17011 ( .A1(n15324), .A2(n15328), .B1(n7795), .B2(n10226), .ZN(
        P1_U3477) );
  NAND2_X1 U17012 ( .A1(n15313), .A2(n15312), .ZN(n15315) );
  NOR2_X1 U17013 ( .A1(n15315), .A2(n15314), .ZN(n15329) );
  AOI22_X1 U17014 ( .A1(n15324), .A2(n15329), .B1(n7807), .B2(n10226), .ZN(
        P1_U3480) );
  OAI21_X1 U17015 ( .B1(n15318), .B2(n15317), .A(n15316), .ZN(n15319) );
  AOI211_X1 U17016 ( .C1(n15322), .C2(n15321), .A(n15320), .B(n15319), .ZN(
        n15331) );
  INV_X1 U17017 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n15323) );
  AOI22_X1 U17018 ( .A1(n15324), .A2(n15331), .B1(n15323), .B2(n10226), .ZN(
        P1_U3483) );
  AOI22_X1 U17019 ( .A1(n15332), .A2(n15325), .B1(n10504), .B2(n15330), .ZN(
        P1_U3528) );
  AOI22_X1 U17020 ( .A1(n15332), .A2(n15326), .B1(n10353), .B2(n15330), .ZN(
        P1_U3529) );
  AOI22_X1 U17021 ( .A1(n15332), .A2(n15327), .B1(n7731), .B2(n15330), .ZN(
        P1_U3530) );
  AOI22_X1 U17022 ( .A1(n15332), .A2(n15328), .B1(n10473), .B2(n15330), .ZN(
        P1_U3534) );
  AOI22_X1 U17023 ( .A1(n15332), .A2(n15329), .B1(n10520), .B2(n15330), .ZN(
        P1_U3535) );
  AOI22_X1 U17024 ( .A1(n15332), .A2(n15331), .B1(n10643), .B2(n15330), .ZN(
        P1_U3536) );
  NOR2_X1 U17025 ( .A1(n15333), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U17026 ( .A1(n15333), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n15346) );
  OAI211_X1 U17027 ( .C1(n15336), .C2(n15335), .A(n15484), .B(n15334), .ZN(
        n15337) );
  INV_X1 U17028 ( .A(n15337), .ZN(n15343) );
  NAND2_X1 U17029 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n15341) );
  INV_X1 U17030 ( .A(n15338), .ZN(n15340) );
  AOI211_X1 U17031 ( .C1(n15341), .C2(n15340), .A(n15339), .B(n15461), .ZN(
        n15342) );
  AOI211_X1 U17032 ( .C1(n7092), .C2(n15344), .A(n15343), .B(n15342), .ZN(
        n15345) );
  NAND2_X1 U17033 ( .A1(n15346), .A2(n15345), .ZN(P2_U3215) );
  OAI211_X1 U17034 ( .C1(n15349), .C2(n15348), .A(n15484), .B(n15347), .ZN(
        n15350) );
  INV_X1 U17035 ( .A(n15350), .ZN(n15355) );
  AOI211_X1 U17036 ( .C1(n15353), .C2(n15352), .A(n15351), .B(n15461), .ZN(
        n15354) );
  AOI211_X1 U17037 ( .C1(n7092), .C2(n15356), .A(n15355), .B(n15354), .ZN(
        n15358) );
  NAND2_X1 U17038 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3088), .ZN(n15357) );
  OAI211_X1 U17039 ( .C1(n15493), .C2(n15359), .A(n15358), .B(n15357), .ZN(
        P2_U3217) );
  OAI211_X1 U17040 ( .C1(n15362), .C2(n15361), .A(n15484), .B(n15360), .ZN(
        n15363) );
  INV_X1 U17041 ( .A(n15363), .ZN(n15368) );
  AOI211_X1 U17042 ( .C1(n15366), .C2(n15365), .A(n15461), .B(n15364), .ZN(
        n15367) );
  AOI211_X1 U17043 ( .C1(n7092), .C2(n15369), .A(n15368), .B(n15367), .ZN(
        n15371) );
  NAND2_X1 U17044 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n15370) );
  OAI211_X1 U17045 ( .C1(n15493), .C2(n15372), .A(n15371), .B(n15370), .ZN(
        P2_U3218) );
  INV_X1 U17046 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15745) );
  OAI211_X1 U17047 ( .C1(n15375), .C2(n15374), .A(n15484), .B(n15373), .ZN(
        n15376) );
  INV_X1 U17048 ( .A(n15376), .ZN(n15381) );
  AOI211_X1 U17049 ( .C1(n15379), .C2(n15378), .A(n15461), .B(n15377), .ZN(
        n15380) );
  AOI211_X1 U17050 ( .C1(n7092), .C2(n15382), .A(n15381), .B(n15380), .ZN(
        n15384) );
  NAND2_X1 U17051 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n15383) );
  OAI211_X1 U17052 ( .C1(n15493), .C2(n15745), .A(n15384), .B(n15383), .ZN(
        P2_U3219) );
  INV_X1 U17053 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n15397) );
  OAI211_X1 U17054 ( .C1(n15387), .C2(n15386), .A(n15484), .B(n15385), .ZN(
        n15388) );
  INV_X1 U17055 ( .A(n15388), .ZN(n15393) );
  AOI211_X1 U17056 ( .C1(n15391), .C2(n15390), .A(n15461), .B(n15389), .ZN(
        n15392) );
  AOI211_X1 U17057 ( .C1(n7092), .C2(n15394), .A(n15393), .B(n15392), .ZN(
        n15396) );
  NAND2_X1 U17058 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n15395) );
  OAI211_X1 U17059 ( .C1(n15493), .C2(n15397), .A(n15396), .B(n15395), .ZN(
        P2_U3220) );
  OAI211_X1 U17060 ( .C1(n15400), .C2(n15399), .A(n15484), .B(n15398), .ZN(
        n15401) );
  INV_X1 U17061 ( .A(n15401), .ZN(n15406) );
  AOI211_X1 U17062 ( .C1(n15404), .C2(n15403), .A(n15461), .B(n15402), .ZN(
        n15405) );
  AOI211_X1 U17063 ( .C1(n7092), .C2(n15407), .A(n15406), .B(n15405), .ZN(
        n15409) );
  NAND2_X1 U17064 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n15408) );
  OAI211_X1 U17065 ( .C1(n15410), .C2(n15493), .A(n15409), .B(n15408), .ZN(
        P2_U3221) );
  AOI211_X1 U17066 ( .C1(n15413), .C2(n15412), .A(n15461), .B(n15411), .ZN(
        n15420) );
  OAI211_X1 U17067 ( .C1(n15416), .C2(n15415), .A(n15484), .B(n15414), .ZN(
        n15417) );
  OAI21_X1 U17068 ( .B1(n15489), .B2(n15418), .A(n15417), .ZN(n15419) );
  NOR2_X1 U17069 ( .A1(n15420), .A2(n15419), .ZN(n15422) );
  OAI211_X1 U17070 ( .C1(n15423), .C2(n15493), .A(n15422), .B(n15421), .ZN(
        P2_U3222) );
  INV_X1 U17071 ( .A(n15424), .ZN(n15425) );
  AOI211_X1 U17072 ( .C1(n15427), .C2(n15426), .A(n15465), .B(n15425), .ZN(
        n15432) );
  AOI211_X1 U17073 ( .C1(n15430), .C2(n15429), .A(n15461), .B(n15428), .ZN(
        n15431) );
  AOI211_X1 U17074 ( .C1(n7092), .C2(n15433), .A(n15432), .B(n15431), .ZN(
        n15435) );
  OAI211_X1 U17075 ( .C1(n15436), .C2(n15493), .A(n15435), .B(n15434), .ZN(
        P2_U3224) );
  INV_X1 U17076 ( .A(n15437), .ZN(n15445) );
  AOI211_X1 U17077 ( .C1(n15439), .C2(n12372), .A(n15438), .B(n15461), .ZN(
        n15444) );
  AOI211_X1 U17078 ( .C1(n15442), .C2(n15441), .A(n15440), .B(n15465), .ZN(
        n15443) );
  AOI211_X1 U17079 ( .C1(n7092), .C2(n15445), .A(n15444), .B(n15443), .ZN(
        n15447) );
  NAND2_X1 U17080 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3088), .ZN(n15446)
         );
  OAI211_X1 U17081 ( .C1(n15448), .C2(n15493), .A(n15447), .B(n15446), .ZN(
        P2_U3229) );
  AOI211_X1 U17082 ( .C1(n15451), .C2(n15450), .A(n15449), .B(n15465), .ZN(
        n15456) );
  AOI211_X1 U17083 ( .C1(n15454), .C2(n15453), .A(n15452), .B(n15461), .ZN(
        n15455) );
  AOI211_X1 U17084 ( .C1(n7092), .C2(n15457), .A(n15456), .B(n15455), .ZN(
        n15459) );
  OAI211_X1 U17085 ( .C1(n15460), .C2(n15493), .A(n15459), .B(n15458), .ZN(
        P2_U3230) );
  AOI211_X1 U17086 ( .C1(n15464), .C2(n15463), .A(n15462), .B(n15461), .ZN(
        n15470) );
  AOI211_X1 U17087 ( .C1(n15468), .C2(n15467), .A(n15466), .B(n15465), .ZN(
        n15469) );
  AOI211_X1 U17088 ( .C1(n7092), .C2(n15471), .A(n15470), .B(n15469), .ZN(
        n15473) );
  OAI211_X1 U17089 ( .C1(n15474), .C2(n15493), .A(n15473), .B(n15472), .ZN(
        P2_U3231) );
  OAI21_X1 U17090 ( .B1(n15477), .B2(n15476), .A(n15475), .ZN(n15479) );
  NAND2_X1 U17091 ( .A1(n15479), .A2(n15478), .ZN(n15487) );
  NAND2_X1 U17092 ( .A1(n15481), .A2(n15480), .ZN(n15485) );
  INV_X1 U17093 ( .A(n15482), .ZN(n15483) );
  NAND3_X1 U17094 ( .A1(n15485), .A2(n15484), .A3(n15483), .ZN(n15486) );
  OAI211_X1 U17095 ( .C1(n15489), .C2(n15488), .A(n15487), .B(n15486), .ZN(
        n15490) );
  INV_X1 U17096 ( .A(n15490), .ZN(n15492) );
  NAND2_X1 U17097 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3088), .ZN(n15491)
         );
  OAI211_X1 U17098 ( .C1(n15494), .C2(n15493), .A(n15492), .B(n15491), .ZN(
        P2_U3232) );
  AND2_X1 U17099 ( .A1(n15496), .A2(n15495), .ZN(n15505) );
  NAND2_X1 U17100 ( .A1(n15498), .A2(n15497), .ZN(n15501) );
  AOI22_X1 U17101 ( .A1(n6677), .A2(P2_REG2_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(n15499), .ZN(n15500) );
  OAI211_X1 U17102 ( .C1(n15503), .C2(n15502), .A(n15501), .B(n15500), .ZN(
        n15504) );
  NOR2_X1 U17103 ( .A1(n15505), .A2(n15504), .ZN(n15506) );
  OAI21_X1 U17104 ( .B1(n6677), .B2(n15507), .A(n15506), .ZN(P2_U3264) );
  AND2_X1 U17105 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15509), .ZN(P2_U3266) );
  AND2_X1 U17106 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15509), .ZN(P2_U3267) );
  AND2_X1 U17107 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15509), .ZN(P2_U3268) );
  AND2_X1 U17108 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15509), .ZN(P2_U3269) );
  AND2_X1 U17109 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15509), .ZN(P2_U3270) );
  AND2_X1 U17110 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15509), .ZN(P2_U3271) );
  AND2_X1 U17111 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15509), .ZN(P2_U3272) );
  AND2_X1 U17112 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15509), .ZN(P2_U3273) );
  AND2_X1 U17113 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15509), .ZN(P2_U3274) );
  AND2_X1 U17114 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15509), .ZN(P2_U3275) );
  AND2_X1 U17115 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15509), .ZN(P2_U3276) );
  AND2_X1 U17116 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15509), .ZN(P2_U3277) );
  AND2_X1 U17117 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15509), .ZN(P2_U3278) );
  AND2_X1 U17118 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15509), .ZN(P2_U3279) );
  AND2_X1 U17119 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15509), .ZN(P2_U3280) );
  AND2_X1 U17120 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15509), .ZN(P2_U3281) );
  AND2_X1 U17121 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15509), .ZN(P2_U3282) );
  AND2_X1 U17122 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15509), .ZN(P2_U3283) );
  AND2_X1 U17123 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15509), .ZN(P2_U3284) );
  AND2_X1 U17124 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15509), .ZN(P2_U3285) );
  AND2_X1 U17125 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15509), .ZN(P2_U3286) );
  AND2_X1 U17126 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15509), .ZN(P2_U3287) );
  AND2_X1 U17127 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15509), .ZN(P2_U3288) );
  AND2_X1 U17128 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15509), .ZN(P2_U3289) );
  AND2_X1 U17129 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15509), .ZN(P2_U3290) );
  AND2_X1 U17130 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15509), .ZN(P2_U3291) );
  AND2_X1 U17131 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15509), .ZN(P2_U3292) );
  AND2_X1 U17132 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15509), .ZN(P2_U3293) );
  AND2_X1 U17133 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15509), .ZN(P2_U3294) );
  AND2_X1 U17134 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15509), .ZN(P2_U3295) );
  AOI22_X1 U17135 ( .A1(n15512), .A2(n15511), .B1(n15510), .B2(n15514), .ZN(
        P2_U3416) );
  AOI21_X1 U17136 ( .B1(n15515), .B2(n15514), .A(n15513), .ZN(P2_U3417) );
  OAI211_X1 U17137 ( .C1(n15518), .C2(n15525), .A(n15517), .B(n15516), .ZN(
        n15519) );
  AOI21_X1 U17138 ( .B1(n15521), .B2(n15520), .A(n15519), .ZN(n15545) );
  INV_X1 U17139 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n15522) );
  AOI22_X1 U17140 ( .A1(n15543), .A2(n15545), .B1(n15522), .B2(n15541), .ZN(
        P2_U3451) );
  INV_X1 U17141 ( .A(n15523), .ZN(n15526) );
  OAI21_X1 U17142 ( .B1(n15526), .B2(n15525), .A(n15524), .ZN(n15527) );
  AOI21_X1 U17143 ( .B1(n15528), .B2(n15537), .A(n15527), .ZN(n15529) );
  AND2_X1 U17144 ( .A1(n15530), .A2(n15529), .ZN(n15547) );
  INV_X1 U17145 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n15531) );
  AOI22_X1 U17146 ( .A1(n15543), .A2(n15547), .B1(n15531), .B2(n15541), .ZN(
        P2_U3454) );
  NAND2_X1 U17147 ( .A1(n15533), .A2(n15532), .ZN(n15534) );
  NAND2_X1 U17148 ( .A1(n15535), .A2(n15534), .ZN(n15536) );
  AOI21_X1 U17149 ( .B1(n15538), .B2(n15537), .A(n15536), .ZN(n15539) );
  AND2_X1 U17150 ( .A1(n15540), .A2(n15539), .ZN(n15549) );
  INV_X1 U17151 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n15542) );
  AOI22_X1 U17152 ( .A1(n15543), .A2(n15549), .B1(n15542), .B2(n15541), .ZN(
        P2_U3460) );
  AOI22_X1 U17153 ( .A1(n15550), .A2(n15545), .B1(n15544), .B2(n15548), .ZN(
        P2_U3506) );
  AOI22_X1 U17154 ( .A1(n15550), .A2(n15547), .B1(n15546), .B2(n15548), .ZN(
        P2_U3507) );
  AOI22_X1 U17155 ( .A1(n15550), .A2(n15549), .B1(n11298), .B2(n15548), .ZN(
        P2_U3509) );
  NOR2_X1 U17156 ( .A1(P3_U3897), .A2(n15674), .ZN(P3_U3150) );
  AOI21_X1 U17157 ( .B1(n11852), .B2(n15552), .A(n15551), .ZN(n15566) );
  INV_X1 U17158 ( .A(n15553), .ZN(n15554) );
  OAI21_X1 U17159 ( .B1(n15591), .B2(n9796), .A(n15554), .ZN(n15560) );
  OR3_X1 U17160 ( .A1(n15557), .A2(n15556), .A3(n15555), .ZN(n15558) );
  AOI21_X1 U17161 ( .B1(n15573), .B2(n15558), .A(n15595), .ZN(n15559) );
  AOI211_X1 U17162 ( .C1(n15600), .C2(n15561), .A(n15560), .B(n15559), .ZN(
        n15565) );
  XNOR2_X1 U17163 ( .A(n15562), .B(P3_REG1_REG_3__SCAN_IN), .ZN(n15563) );
  NAND2_X1 U17164 ( .A1(n15677), .A2(n15563), .ZN(n15564) );
  OAI211_X1 U17165 ( .C1(n15566), .C2(n15681), .A(n15565), .B(n15564), .ZN(
        P3_U3185) );
  AOI21_X1 U17166 ( .B1(n15568), .B2(n15567), .A(n6820), .ZN(n15586) );
  INV_X1 U17167 ( .A(n15569), .ZN(n15570) );
  OAI21_X1 U17168 ( .B1(n15591), .B2(n9389), .A(n15570), .ZN(n15577) );
  INV_X1 U17169 ( .A(n15594), .ZN(n15575) );
  NAND3_X1 U17170 ( .A1(n15573), .A2(n15572), .A3(n15571), .ZN(n15574) );
  AOI21_X1 U17171 ( .B1(n15575), .B2(n15574), .A(n15595), .ZN(n15576) );
  AOI211_X1 U17172 ( .C1(n15600), .C2(n15578), .A(n15577), .B(n15576), .ZN(
        n15585) );
  AOI21_X1 U17173 ( .B1(n15581), .B2(n15580), .A(n15579), .ZN(n15582) );
  OR2_X1 U17174 ( .A1(n15583), .A2(n15582), .ZN(n15584) );
  OAI211_X1 U17175 ( .C1(n15586), .C2(n15681), .A(n15585), .B(n15584), .ZN(
        P3_U3186) );
  AOI21_X1 U17176 ( .B1(n11862), .B2(n15588), .A(n15587), .ZN(n15606) );
  INV_X1 U17177 ( .A(n15589), .ZN(n15590) );
  OAI21_X1 U17178 ( .B1(n15591), .B2(n9393), .A(n15590), .ZN(n15598) );
  OR3_X1 U17179 ( .A1(n15594), .A2(n15593), .A3(n15592), .ZN(n15596) );
  AOI21_X1 U17180 ( .B1(n15612), .B2(n15596), .A(n15595), .ZN(n15597) );
  AOI211_X1 U17181 ( .C1(n15600), .C2(n15599), .A(n15598), .B(n15597), .ZN(
        n15605) );
  XNOR2_X1 U17182 ( .A(n15602), .B(n15601), .ZN(n15603) );
  NAND2_X1 U17183 ( .A1(n15677), .A2(n15603), .ZN(n15604) );
  OAI211_X1 U17184 ( .C1(n15606), .C2(n15681), .A(n15605), .B(n15604), .ZN(
        P3_U3187) );
  AOI21_X1 U17185 ( .B1(n15609), .B2(n15608), .A(n15607), .ZN(n15624) );
  AND3_X1 U17186 ( .A1(n15612), .A2(n15611), .A3(n15610), .ZN(n15613) );
  OAI21_X1 U17187 ( .B1(n15629), .B2(n15613), .A(n15666), .ZN(n15614) );
  OAI21_X1 U17188 ( .B1(n15671), .B2(n15615), .A(n15614), .ZN(n15616) );
  AOI211_X1 U17189 ( .C1(P3_ADDR_REG_6__SCAN_IN), .C2(n15674), .A(n15617), .B(
        n15616), .ZN(n15623) );
  OAI21_X1 U17190 ( .B1(n15620), .B2(n15619), .A(n15618), .ZN(n15621) );
  NAND2_X1 U17191 ( .A1(n15677), .A2(n15621), .ZN(n15622) );
  OAI211_X1 U17192 ( .C1(n15624), .C2(n15681), .A(n15623), .B(n15622), .ZN(
        P3_U3188) );
  AOI21_X1 U17193 ( .B1(n11874), .B2(n15626), .A(n15625), .ZN(n15641) );
  INV_X1 U17194 ( .A(n15646), .ZN(n15631) );
  NOR3_X1 U17195 ( .A1(n15629), .A2(n15628), .A3(n15627), .ZN(n15630) );
  OAI21_X1 U17196 ( .B1(n15631), .B2(n15630), .A(n15666), .ZN(n15632) );
  OAI21_X1 U17197 ( .B1(n15671), .B2(n15633), .A(n15632), .ZN(n15634) );
  AOI211_X1 U17198 ( .C1(P3_ADDR_REG_7__SCAN_IN), .C2(n15674), .A(n15635), .B(
        n15634), .ZN(n15640) );
  OAI21_X1 U17199 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n15637), .A(n15636), .ZN(
        n15638) );
  NAND2_X1 U17200 ( .A1(n15638), .A2(n15677), .ZN(n15639) );
  OAI211_X1 U17201 ( .C1(n15641), .C2(n15681), .A(n15640), .B(n15639), .ZN(
        P3_U3189) );
  AOI21_X1 U17202 ( .B1(n6817), .B2(n15643), .A(n15642), .ZN(n15658) );
  AND3_X1 U17203 ( .A1(n15646), .A2(n15645), .A3(n15644), .ZN(n15647) );
  OAI21_X1 U17204 ( .B1(n15665), .B2(n15647), .A(n15666), .ZN(n15648) );
  OAI21_X1 U17205 ( .B1(n15671), .B2(n15649), .A(n15648), .ZN(n15650) );
  AOI211_X1 U17206 ( .C1(P3_ADDR_REG_8__SCAN_IN), .C2(n15674), .A(n15651), .B(
        n15650), .ZN(n15657) );
  OAI21_X1 U17207 ( .B1(n15654), .B2(n15653), .A(n15652), .ZN(n15655) );
  NAND2_X1 U17208 ( .A1(n15655), .A2(n15677), .ZN(n15656) );
  OAI211_X1 U17209 ( .C1(n15658), .C2(n15681), .A(n15657), .B(n15656), .ZN(
        P3_U3190) );
  AOI21_X1 U17210 ( .B1(n15661), .B2(n15660), .A(n15659), .ZN(n15682) );
  INV_X1 U17211 ( .A(n15662), .ZN(n15668) );
  NOR3_X1 U17212 ( .A1(n15665), .A2(n15664), .A3(n15663), .ZN(n15667) );
  OAI21_X1 U17213 ( .B1(n15668), .B2(n15667), .A(n15666), .ZN(n15669) );
  OAI21_X1 U17214 ( .B1(n15671), .B2(n15670), .A(n15669), .ZN(n15672) );
  AOI211_X1 U17215 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n15674), .A(n15673), .B(
        n15672), .ZN(n15680) );
  OAI21_X1 U17216 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n15676), .A(n15675), .ZN(
        n15678) );
  NAND2_X1 U17217 ( .A1(n15678), .A2(n15677), .ZN(n15679) );
  OAI211_X1 U17218 ( .C1(n15682), .C2(n15681), .A(n15680), .B(n15679), .ZN(
        P3_U3191) );
  NAND2_X1 U17219 ( .A1(n15683), .A2(n15684), .ZN(n15685) );
  XNOR2_X1 U17220 ( .A(n15685), .B(n15687), .ZN(n15695) );
  OAI21_X1 U17221 ( .B1(n15688), .B2(n15687), .A(n15686), .ZN(n15711) );
  OAI22_X1 U17222 ( .A1(n15691), .A2(n15690), .B1(n8839), .B2(n15689), .ZN(
        n15692) );
  AOI21_X1 U17223 ( .B1(n15711), .B2(n15693), .A(n15692), .ZN(n15694) );
  OAI21_X1 U17224 ( .B1(n15696), .B2(n15695), .A(n15694), .ZN(n15709) );
  NOR2_X1 U17225 ( .A1(n15697), .A2(n15719), .ZN(n15710) );
  AOI22_X1 U17226 ( .A1(n15711), .A2(n15699), .B1(n15710), .B2(n15698), .ZN(
        n15700) );
  INV_X1 U17227 ( .A(n15700), .ZN(n15701) );
  AOI211_X1 U17228 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n15702), .A(n15709), .B(
        n15701), .ZN(n15704) );
  AOI22_X1 U17229 ( .A1(n13921), .A2(n10951), .B1(n15704), .B2(n15703), .ZN(
        P3_U3231) );
  AOI211_X1 U17230 ( .C1(n15724), .C2(n15707), .A(n15706), .B(n15705), .ZN(
        n15735) );
  INV_X1 U17231 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15708) );
  AOI22_X1 U17232 ( .A1(n15734), .A2(n15735), .B1(n15708), .B2(n15732), .ZN(
        P3_U3393) );
  AOI211_X1 U17233 ( .C1(n15716), .C2(n15711), .A(n15710), .B(n15709), .ZN(
        n15736) );
  INV_X1 U17234 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15712) );
  AOI22_X1 U17235 ( .A1(n15734), .A2(n15736), .B1(n15712), .B2(n15732), .ZN(
        P3_U3396) );
  NOR2_X1 U17236 ( .A1(n15713), .A2(n15719), .ZN(n15715) );
  AOI211_X1 U17237 ( .C1(n15717), .C2(n15716), .A(n15715), .B(n15714), .ZN(
        n15737) );
  INV_X1 U17238 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15718) );
  AOI22_X1 U17239 ( .A1(n15734), .A2(n15737), .B1(n15718), .B2(n15732), .ZN(
        P3_U3399) );
  NOR2_X1 U17240 ( .A1(n15720), .A2(n15719), .ZN(n15722) );
  AOI211_X1 U17241 ( .C1(n15724), .C2(n15723), .A(n15722), .B(n15721), .ZN(
        n15738) );
  INV_X1 U17242 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15725) );
  AOI22_X1 U17243 ( .A1(n15734), .A2(n15738), .B1(n15725), .B2(n15732), .ZN(
        P3_U3408) );
  NOR2_X1 U17244 ( .A1(n15727), .A2(n15726), .ZN(n15729) );
  AOI211_X1 U17245 ( .C1(n15731), .C2(n15730), .A(n15729), .B(n15728), .ZN(
        n15740) );
  INV_X1 U17246 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15733) );
  AOI22_X1 U17247 ( .A1(n15734), .A2(n15740), .B1(n15733), .B2(n15732), .ZN(
        P3_U3420) );
  AOI22_X1 U17248 ( .A1(n15741), .A2(n15735), .B1(n10871), .B2(n15739), .ZN(
        P3_U3460) );
  AOI22_X1 U17249 ( .A1(n15741), .A2(n15736), .B1(n11899), .B2(n15739), .ZN(
        P3_U3461) );
  AOI22_X1 U17250 ( .A1(n15741), .A2(n15737), .B1(n11851), .B2(n15739), .ZN(
        P3_U3462) );
  AOI22_X1 U17251 ( .A1(n15741), .A2(n15738), .B1(n11867), .B2(n15739), .ZN(
        P3_U3465) );
  AOI22_X1 U17252 ( .A1(n15741), .A2(n15740), .B1(n11888), .B2(n15739), .ZN(
        P3_U3469) );
  XOR2_X1 U17253 ( .A(n15743), .B(n15742), .Z(SUB_1596_U59) );
  XOR2_X1 U17254 ( .A(n15745), .B(n15744), .Z(SUB_1596_U58) );
  AOI21_X1 U17255 ( .B1(n15747), .B2(n15746), .A(n15755), .ZN(SUB_1596_U53) );
  XOR2_X1 U17256 ( .A(n15749), .B(n15748), .Z(SUB_1596_U56) );
  AOI21_X1 U17257 ( .B1(n15752), .B2(n15751), .A(n15750), .ZN(n15753) );
  XOR2_X1 U17258 ( .A(n15753), .B(P2_ADDR_REG_3__SCAN_IN), .Z(SUB_1596_U60) );
  XOR2_X1 U17259 ( .A(n15755), .B(n15754), .Z(SUB_1596_U5) );
  CLKBUF_X1 U7427 ( .A(n12579), .Z(n6683) );
  NAND2_X1 U7429 ( .A1(n11159), .A2(n13679), .ZN(n11163) );
  OR2_X1 U7430 ( .A1(n14343), .A2(n7221), .ZN(n7218) );
  INV_X1 U7432 ( .A(n12970), .ZN(n11573) );
  INV_X2 U7444 ( .A(n12970), .ZN(n13364) );
  CLKBUF_X3 U7453 ( .A(n10697), .Z(n13112) );
  CLKBUF_X1 U7469 ( .A(n7779), .Z(n10200) );
  CLKBUF_X3 U7639 ( .A(n7770), .Z(n12751) );
  CLKBUF_X1 U9372 ( .A(n13667), .Z(n13629) );
  NAND4_X1 U14424 ( .A1(n7767), .A2(n7766), .A3(n7765), .A4(n7764), .ZN(n14660) );
endmodule

