

module b22_C_AntiSAT_k_256_10 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, SUB_1596_U4, SUB_1596_U62, 
        SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, 
        SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, 
        SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, 
        SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, 
        P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, 
        P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, 
        P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, 
        P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, 
        P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, 
        P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, 
        P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, 
        P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, 
        P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, 
        P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, 
        P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, 
        P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, 
        P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, 
        P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, 
        P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, 
        P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, 
        P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, 
        P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, 
        P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, 
        P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, 
        P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, 
        P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, 
        P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, 
        P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, 
        P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, 
        P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, 
        P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, 
        P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, 
        P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, 
        P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, 
        P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, 
        P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, 
        P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, 
        P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, 
        P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, 
        P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, 
        P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, 
        P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, 
        P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, 
        P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, 
        P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, 
        P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, 
        P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, 
        P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, 
        P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, 
        P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, 
        P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, 
        P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, 
        P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, 
        P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, 
        P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, 
        P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, 
        P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, 
        P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, 
        P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, 
        P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, 
        P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, 
        P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, 
        P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, 
        P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, 
        P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, 
        P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, 
        P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, 
        P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, 
        P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, 
        P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, 
        P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, 
        P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, 
        P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, 
        P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, 
        P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, 
        P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, 
        P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, 
        P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, 
        P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, 
        P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, 
        P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, 
        P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, 
        P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, 
        P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, 
        P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, 
        P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, 
        P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, 
        P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, 
        P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, 
        P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, 
        P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, 
        P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, 
        P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, 
        P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, 
        P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127,
         keyinput128, keyinput129, keyinput130, keyinput131, keyinput132,
         keyinput133, keyinput134, keyinput135, keyinput136, keyinput137,
         keyinput138, keyinput139, keyinput140, keyinput141, keyinput142,
         keyinput143, keyinput144, keyinput145, keyinput146, keyinput147,
         keyinput148, keyinput149, keyinput150, keyinput151, keyinput152,
         keyinput153, keyinput154, keyinput155, keyinput156, keyinput157,
         keyinput158, keyinput159, keyinput160, keyinput161, keyinput162,
         keyinput163, keyinput164, keyinput165, keyinput166, keyinput167,
         keyinput168, keyinput169, keyinput170, keyinput171, keyinput172,
         keyinput173, keyinput174, keyinput175, keyinput176, keyinput177,
         keyinput178, keyinput179, keyinput180, keyinput181, keyinput182,
         keyinput183, keyinput184, keyinput185, keyinput186, keyinput187,
         keyinput188, keyinput189, keyinput190, keyinput191, keyinput192,
         keyinput193, keyinput194, keyinput195, keyinput196, keyinput197,
         keyinput198, keyinput199, keyinput200, keyinput201, keyinput202,
         keyinput203, keyinput204, keyinput205, keyinput206, keyinput207,
         keyinput208, keyinput209, keyinput210, keyinput211, keyinput212,
         keyinput213, keyinput214, keyinput215, keyinput216, keyinput217,
         keyinput218, keyinput219, keyinput220, keyinput221, keyinput222,
         keyinput223, keyinput224, keyinput225, keyinput226, keyinput227,
         keyinput228, keyinput229, keyinput230, keyinput231, keyinput232,
         keyinput233, keyinput234, keyinput235, keyinput236, keyinput237,
         keyinput238, keyinput239, keyinput240, keyinput241, keyinput242,
         keyinput243, keyinput244, keyinput245, keyinput246, keyinput247,
         keyinput248, keyinput249, keyinput250, keyinput251, keyinput252,
         keyinput253, keyinput254, keyinput255;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
         n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
         n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
         n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
         n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
         n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
         n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
         n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
         n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
         n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
         n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
         n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
         n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,
         n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
         n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
         n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
         n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,
         n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
         n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
         n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,
         n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,
         n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
         n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
         n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
         n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
         n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118,
         n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,
         n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
         n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
         n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
         n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230,
         n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
         n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
         n15247, n15248, n15249, n15250, n15251, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564;

  NOR2_X1 U7384 ( .A1(n7211), .A2(n14406), .ZN(n14365) );
  OAI21_X1 U7385 ( .B1(n7441), .B2(n12584), .A(n6978), .ZN(n12612) );
  INV_X1 U7386 ( .A(n12712), .ZN(n12684) );
  OR2_X1 U7387 ( .A1(n11320), .A2(n11260), .ZN(n7361) );
  CLKBUF_X1 U7388 ( .A(n7853), .Z(n7929) );
  INV_X2 U7390 ( .A(n11957), .ZN(n11966) );
  CLKBUF_X2 U7391 ( .A(n12329), .Z(n6640) );
  NAND2_X2 U7392 ( .A1(n9611), .A2(n10184), .ZN(n11968) );
  BUF_X4 U7393 ( .A(n11048), .Z(n6638) );
  BUF_X2 U7394 ( .A(n9270), .Z(n12338) );
  NAND2_X1 U7395 ( .A1(n10529), .A2(n14038), .ZN(n9270) );
  INV_X2 U7396 ( .A(n14044), .ZN(n14198) );
  NAND2_X1 U7397 ( .A1(n14030), .A2(n7550), .ZN(n14044) );
  OR2_X1 U7398 ( .A1(n9151), .A2(n13840), .ZN(n8426) );
  AND2_X2 U7399 ( .A1(n11908), .A2(n8443), .ZN(n8497) );
  NOR2_X2 U7400 ( .A1(n14195), .A2(n14010), .ZN(n14038) );
  AND2_X1 U7401 ( .A1(n11909), .A2(n9258), .ZN(n9954) );
  AND3_X1 U7402 ( .A1(n9207), .A2(n9206), .A3(n9209), .ZN(n6668) );
  INV_X1 U7403 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n7536) );
  INV_X1 U7404 ( .A(n14038), .ZN(n9831) );
  NAND2_X1 U7405 ( .A1(n14699), .A2(n14352), .ZN(n14008) );
  OR2_X1 U7406 ( .A1(n10416), .A2(n7445), .ZN(n7443) );
  INV_X1 U7407 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9679) );
  OR2_X1 U7408 ( .A1(n11311), .A2(n11269), .ZN(n6985) );
  AND2_X1 U7409 ( .A1(n10945), .A2(n7885), .ZN(n11215) );
  NAND2_X1 U7410 ( .A1(n12051), .A2(n12050), .ZN(n10025) );
  NOR2_X1 U7411 ( .A1(n10145), .A2(n8069), .ZN(n7430) );
  INV_X1 U7412 ( .A(n6838), .ZN(n11961) );
  BUF_X1 U7413 ( .A(n11759), .Z(n6648) );
  OR2_X1 U7414 ( .A1(n14739), .A2(n14738), .ZN(n14740) );
  AND2_X1 U7415 ( .A1(n7635), .A2(n9235), .ZN(n7637) );
  INV_X1 U7416 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n7537) );
  INV_X1 U7417 ( .A(n6823), .ZN(n12390) );
  INV_X1 U7418 ( .A(n12743), .ZN(n12476) );
  OR2_X1 U7419 ( .A1(n15414), .A2(n7437), .ZN(n7436) );
  XNOR2_X1 U7420 ( .A(n11902), .B(n12633), .ZN(n12622) );
  NOR2_X1 U7422 ( .A1(n15059), .A2(n15060), .ZN(n15058) );
  NOR2_X1 U7423 ( .A1(n14406), .A2(n14608), .ZN(n14391) );
  NAND2_X1 U7424 ( .A1(n9108), .A2(n9075), .ZN(n9078) );
  INV_X1 U7425 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9484) );
  INV_X1 U7426 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9233) );
  NAND2_X1 U7427 ( .A1(n8263), .A2(n8246), .ZN(n9388) );
  INV_X1 U7428 ( .A(n14071), .ZN(n13978) );
  OAI21_X1 U7429 ( .B1(n9748), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9745), .ZN(
        n9878) );
  INV_X2 U7430 ( .A(n14352), .ZN(n14579) );
  AOI211_X1 U7431 ( .C1(n14603), .C2(n15191), .A(n14602), .B(n14601), .ZN(
        n14604) );
  XNOR2_X1 U7432 ( .A(n8807), .B(n8806), .ZN(n11670) );
  INV_X1 U7433 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9353) );
  AOI211_X1 U7434 ( .C1(n12652), .C2(n12651), .A(n12650), .B(n12649), .ZN(
        n12653) );
  BUF_X1 U7435 ( .A(n10317), .Z(n6641) );
  AND2_X1 U7436 ( .A1(n9614), .A2(n8463), .ZN(n6636) );
  NAND2_X2 U7437 ( .A1(n10127), .A2(n6832), .ZN(n11999) );
  INV_X1 U7438 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8069) );
  INV_X1 U7440 ( .A(n9270), .ZN(n11048) );
  INV_X1 U7441 ( .A(n12340), .ZN(n12329) );
  NOR2_X1 U7442 ( .A1(n10118), .A2(n7638), .ZN(n9236) );
  OR2_X1 U7443 ( .A1(n9288), .A2(n9233), .ZN(n9290) );
  NOR2_X2 U7444 ( .A1(n12201), .A2(n15463), .ZN(n15460) );
  NAND4_X2 U7445 ( .A1(n7790), .A2(n7792), .A3(n7791), .A4(n7789), .ZN(n15463)
         );
  NAND2_X2 U7446 ( .A1(n14985), .A2(n14987), .ZN(n8379) );
  XNOR2_X2 U7447 ( .A(n8245), .B(P3_IR_REG_26__SCAN_IN), .ZN(n8263) );
  NAND4_X2 U7448 ( .A1(n9851), .A2(n9850), .A3(n9849), .A4(n9848), .ZN(n14280)
         );
  AND2_X2 U7449 ( .A1(n9214), .A2(n7566), .ZN(n9240) );
  NOR2_X2 U7450 ( .A1(n10859), .A2(n14075), .ZN(n7202) );
  AOI21_X2 U7451 ( .B1(n11072), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10049), .ZN(
        n15004) );
  NOR2_X2 U7452 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n8412) );
  NAND2_X2 U7453 ( .A1(n8211), .A2(n12085), .ZN(n11146) );
  NOR2_X2 U7454 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n8431) );
  INV_X1 U7455 ( .A(n14062), .ZN(n11060) );
  OAI211_X2 U7456 ( .C1(n6845), .C2(n10324), .A(n10323), .B(n10322), .ZN(
        n14062) );
  NAND2_X2 U7457 ( .A1(n8654), .A2(n8653), .ZN(n8694) );
  XNOR2_X2 U7458 ( .A(n9078), .B(n9077), .ZN(n14692) );
  NAND2_X2 U7459 ( .A1(n15409), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n15406) );
  NAND4_X2 U7460 ( .A1(n8175), .A2(n8174), .A3(n8173), .A4(n8172), .ZN(n12699)
         );
  XNOR2_X2 U7461 ( .A(n8385), .B(n8384), .ZN(n14994) );
  NAND2_X1 U7462 ( .A1(n10520), .A2(n10519), .ZN(n10544) );
  XNOR2_X2 U7463 ( .A(n14644), .B(n14506), .ZN(n14495) );
  XNOR2_X1 U7464 ( .A(n8428), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8460) );
  NAND2_X2 U7465 ( .A1(n14989), .A2(n8381), .ZN(n8385) );
  INV_X4 U7466 ( .A(n14016), .ZN(n11774) );
  INV_X2 U7467 ( .A(n9954), .ZN(n14016) );
  OAI21_X2 U7468 ( .B1(n11032), .B2(n7138), .A(n7135), .ZN(n13973) );
  OAI21_X2 U7469 ( .B1(n8244), .B2(P3_IR_REG_25__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8245) );
  AOI21_X4 U7470 ( .B1(n13887), .B2(n12291), .A(n7677), .ZN(n13950) );
  NAND2_X2 U7471 ( .A1(n7144), .A2(n6770), .ZN(n13887) );
  INV_X1 U7472 ( .A(n15442), .ZN(n9995) );
  XNOR2_X2 U7473 ( .A(n8390), .B(n8389), .ZN(n14997) );
  NOR2_X1 U7474 ( .A1(n14048), .A2(n14047), .ZN(n14051) );
  XNOR2_X2 U7475 ( .A(n8426), .B(n8425), .ZN(n9571) );
  NAND2_X2 U7476 ( .A1(n14992), .A2(n8387), .ZN(n8390) );
  OAI222_X1 U7477 ( .A1(P2_U3088), .A2(n13538), .B1(n13854), .B2(n9336), .C1(
        n9337), .C2(n13852), .ZN(P2_U3325) );
  OR2_X1 U7478 ( .A1(n14025), .A2(n9336), .ZN(n9938) );
  XNOR2_X2 U7479 ( .A(n8364), .B(n7277), .ZN(n14711) );
  NAND2_X2 U7480 ( .A1(n15551), .A2(n8361), .ZN(n8364) );
  AOI22_X2 U7481 ( .A1(n10304), .A2(n10305), .B1(n10317), .B2(n10135), .ZN(
        n10430) );
  NOR2_X1 U7482 ( .A1(n15562), .A2(n8353), .ZN(n14707) );
  INV_X2 U7483 ( .A(n14044), .ZN(n6639) );
  INV_X4 U7484 ( .A(n14198), .ZN(n14187) );
  NOR2_X2 U7485 ( .A1(n12612), .A2(n11900), .ZN(n11902) );
  XNOR2_X2 U7486 ( .A(n8299), .B(n7272), .ZN(n8346) );
  NAND2_X2 U7487 ( .A1(n7275), .A2(n7273), .ZN(n8299) );
  XNOR2_X2 U7488 ( .A(n9286), .B(n7013), .ZN(n9802) );
  OAI21_X1 U7489 ( .B1(n6879), .B2(n6678), .A(n7559), .ZN(n14189) );
  AOI21_X1 U7490 ( .B1(n13858), .B2(n13859), .A(n6717), .ZN(n12346) );
  XNOR2_X1 U7491 ( .A(n12396), .B(n12699), .ZN(n12681) );
  NAND2_X1 U7492 ( .A1(n12406), .A2(n12373), .ZN(n12489) );
  OR2_X1 U7493 ( .A1(n14999), .A2(n15000), .ZN(n6856) );
  NAND2_X1 U7494 ( .A1(n7108), .A2(n11643), .ZN(n14608) );
  NAND2_X1 U7495 ( .A1(n12819), .A2(n12128), .ZN(n12831) );
  OAI21_X1 U7496 ( .B1(n7438), .B2(n12570), .A(n6976), .ZN(n6979) );
  OR2_X1 U7497 ( .A1(n12560), .A2(n11868), .ZN(n7438) );
  AOI21_X1 U7498 ( .B1(n11275), .B2(n11274), .A(n11273), .ZN(n15433) );
  NAND2_X1 U7499 ( .A1(n9837), .A2(n9838), .ZN(n10068) );
  INV_X2 U7500 ( .A(n12379), .ZN(n12416) );
  NAND2_X1 U7501 ( .A1(n9997), .A2(n7796), .ZN(n12051) );
  XNOR2_X1 U7502 ( .A(n11060), .B(n6897), .ZN(n10562) );
  INV_X1 U7503 ( .A(n14277), .ZN(n6897) );
  CLKBUF_X3 U7504 ( .A(n8186), .Z(n8170) );
  INV_X1 U7505 ( .A(n9935), .ZN(n10626) );
  CLKBUF_X3 U7507 ( .A(n7799), .Z(n12001) );
  INV_X1 U7508 ( .A(n11999), .ZN(n6820) );
  AND2_X1 U7509 ( .A1(n7702), .A2(n13027), .ZN(n7800) );
  INV_X8 U7510 ( .A(n9143), .ZN(n9113) );
  INV_X2 U7511 ( .A(n9121), .ZN(n9143) );
  NAND2_X1 U7512 ( .A1(n7330), .A2(n8474), .ZN(n9645) );
  BUF_X2 U7513 ( .A(n9115), .Z(n6860) );
  BUF_X2 U7514 ( .A(n9096), .Z(n6652) );
  AND2_X1 U7515 ( .A1(n9258), .A2(n9259), .ZN(n9942) );
  AOI21_X1 U7516 ( .B1(n9735), .B2(P1_REG1_REG_4__SCAN_IN), .A(n9726), .ZN(
        n9747) );
  CLKBUF_X3 U7517 ( .A(n8497), .Z(n6651) );
  CLKBUF_X2 U7518 ( .A(n8502), .Z(n9110) );
  AND2_X1 U7519 ( .A1(n8443), .A2(n8441), .ZN(n9096) );
  NAND2_X1 U7520 ( .A1(n7581), .A2(n8488), .ZN(n8527) );
  NAND2_X1 U7521 ( .A1(n9255), .A2(n14689), .ZN(n11621) );
  INV_X4 U7522 ( .A(n12187), .ZN(n6642) );
  INV_X2 U7523 ( .A(n8533), .ZN(n6643) );
  NAND2_X1 U7524 ( .A1(n9216), .A2(n6810), .ZN(n9248) );
  XNOR2_X1 U7525 ( .A(n9234), .B(n9235), .ZN(n9265) );
  NAND2_X1 U7526 ( .A1(n9240), .A2(n9215), .ZN(n9246) );
  NAND2_X1 U7527 ( .A1(n9823), .A2(n6672), .ZN(n14352) );
  CLKBUF_X1 U7529 ( .A(n8722), .Z(n8723) );
  AND2_X1 U7530 ( .A1(n8722), .A2(n8414), .ZN(n8421) );
  AND3_X1 U7531 ( .A1(n7686), .A2(n7479), .A3(n7196), .ZN(n7195) );
  NOR2_X1 U7532 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n9288) );
  INV_X1 U7533 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9284) );
  AOI21_X1 U7534 ( .B1(n6671), .B2(n6871), .A(n6825), .ZN(n12193) );
  MUX2_X1 U7535 ( .A(n12896), .B(n12964), .S(n15547), .Z(n12897) );
  NOR2_X1 U7536 ( .A1(n12894), .A2(n6687), .ZN(n12964) );
  OR2_X1 U7537 ( .A1(n12203), .A2(n14790), .ZN(n8236) );
  OR2_X1 U7538 ( .A1(n12203), .A2(n12888), .ZN(n6822) );
  AOI21_X1 U7539 ( .B1(n11831), .B2(n14841), .A(n11830), .ZN(n13764) );
  AOI22_X1 U7540 ( .A1(n13491), .A2(n13490), .B1(n7516), .B2(n7513), .ZN(
        n13504) );
  NAND2_X1 U7541 ( .A1(n7618), .A2(n14420), .ZN(n14419) );
  CLKBUF_X1 U7542 ( .A(n12396), .Z(n6864) );
  CLKBUF_X1 U7543 ( .A(n13679), .Z(n6911) );
  NAND2_X1 U7544 ( .A1(n13453), .A2(n11953), .ZN(n13420) );
  NAND2_X1 U7545 ( .A1(n12737), .A2(n12740), .ZN(n12739) );
  NAND2_X1 U7546 ( .A1(n13962), .A2(n13963), .ZN(n7144) );
  NAND2_X1 U7547 ( .A1(n8131), .A2(n8130), .ZN(n12483) );
  NAND2_X1 U7548 ( .A1(n13664), .A2(n13663), .ZN(n13662) );
  NAND2_X1 U7549 ( .A1(n13914), .A2(n12260), .ZN(n13962) );
  NAND2_X1 U7550 ( .A1(n8153), .A2(n8152), .ZN(n12898) );
  NAND2_X1 U7551 ( .A1(n13915), .A2(n13916), .ZN(n13914) );
  NAND2_X1 U7552 ( .A1(n11946), .A2(n11945), .ZN(n13449) );
  NAND2_X1 U7553 ( .A1(n11949), .A2(n13395), .ZN(n7532) );
  OAI21_X1 U7554 ( .B1(n7548), .B2(n7547), .A(n7546), .ZN(n14164) );
  NAND2_X1 U7555 ( .A1(n8142), .A2(n8141), .ZN(n12454) );
  NAND2_X1 U7556 ( .A1(n12489), .A2(n12488), .ZN(n12487) );
  NAND2_X1 U7557 ( .A1(n6922), .A2(n6956), .ZN(n14466) );
  OR2_X1 U7558 ( .A1(n13699), .A2(n13700), .ZN(n13697) );
  NAND2_X1 U7559 ( .A1(n13996), .A2(n13995), .ZN(n13993) );
  NAND2_X1 U7560 ( .A1(n8119), .A2(n8118), .ZN(n12749) );
  OAI21_X1 U7561 ( .B1(n13712), .B2(n11819), .A(n11820), .ZN(n13699) );
  XNOR2_X1 U7562 ( .A(n12248), .B(n12249), .ZN(n13996) );
  NAND2_X1 U7563 ( .A1(n6803), .A2(n8108), .ZN(n12985) );
  NAND2_X1 U7564 ( .A1(n8097), .A2(n8096), .ZN(n12989) );
  NAND2_X1 U7565 ( .A1(n13438), .A2(n11927), .ZN(n13483) );
  NAND2_X1 U7566 ( .A1(n13743), .A2(n13751), .ZN(n13742) );
  NAND2_X1 U7567 ( .A1(n13439), .A2(n13440), .ZN(n13438) );
  NAND2_X1 U7568 ( .A1(n14823), .A2(n11582), .ZN(n13743) );
  NAND2_X1 U7569 ( .A1(n13429), .A2(n11922), .ZN(n13439) );
  XNOR2_X1 U7570 ( .A(n9091), .B(n9090), .ZN(n11772) );
  NAND2_X1 U7571 ( .A1(n11444), .A2(n12095), .ZN(n14769) );
  AND2_X1 U7572 ( .A1(n12042), .A2(n12837), .ZN(n12852) );
  NAND2_X1 U7573 ( .A1(n11659), .A2(n11658), .ZN(n14431) );
  INV_X1 U7574 ( .A(n12831), .ZN(n6644) );
  NAND2_X1 U7575 ( .A1(n8909), .A2(n8908), .ZN(n13804) );
  OR2_X1 U7576 ( .A1(n11009), .A2(n11008), .ZN(n11011) );
  AND2_X1 U7577 ( .A1(n8025), .A2(n8024), .ZN(n12856) );
  OAI21_X1 U7578 ( .B1(n11146), .B2(n12092), .A(n12090), .ZN(n11328) );
  XNOR2_X1 U7579 ( .A(n8985), .B(SI_24_), .ZN(n8983) );
  AND2_X1 U7580 ( .A1(n14698), .A2(n6845), .ZN(n14639) );
  NAND2_X1 U7581 ( .A1(n11104), .A2(n14229), .ZN(n11416) );
  NAND2_X1 U7582 ( .A1(n6828), .A2(n6827), .ZN(n11278) );
  NAND2_X1 U7583 ( .A1(n7366), .A2(n7367), .ZN(n11104) );
  NAND2_X1 U7584 ( .A1(n7076), .A2(n7074), .ZN(n11213) );
  NAND3_X1 U7585 ( .A1(n7191), .A2(n7190), .A3(n6674), .ZN(n10910) );
  NAND2_X1 U7586 ( .A1(n11537), .A2(n11536), .ZN(n14956) );
  NAND2_X1 U7587 ( .A1(n11672), .A2(n11671), .ZN(n14921) );
  AND2_X1 U7588 ( .A1(n6901), .A2(n7739), .ZN(n7969) );
  NAND2_X1 U7589 ( .A1(n6965), .A2(n6662), .ZN(n7124) );
  OR2_X1 U7590 ( .A1(n7285), .A2(n8719), .ZN(n6901) );
  NAND2_X1 U7591 ( .A1(n8677), .A2(n8676), .ZN(n11170) );
  INV_X2 U7592 ( .A(n15477), .ZN(n12871) );
  NAND2_X1 U7593 ( .A1(n8748), .A2(n8747), .ZN(n8768) );
  AND2_X1 U7594 ( .A1(n12071), .A2(n12070), .ZN(n12025) );
  AND2_X1 U7595 ( .A1(n12058), .A2(n12043), .ZN(n12019) );
  INV_X1 U7596 ( .A(n10947), .ZN(n12547) );
  NAND2_X1 U7597 ( .A1(n9274), .A2(n9836), .ZN(n9835) );
  INV_X1 U7598 ( .A(n10114), .ZN(n12201) );
  NAND2_X1 U7599 ( .A1(n7803), .A2(n6694), .ZN(n15462) );
  NAND4_X1 U7600 ( .A1(n8501), .A2(n8500), .A3(n8499), .A4(n8498), .ZN(n13531)
         );
  NAND2_X1 U7601 ( .A1(n9249), .A2(n6647), .ZN(n12337) );
  AOI21_X1 U7602 ( .B1(n6969), .B2(n6972), .A(n6968), .ZN(n6967) );
  CLKBUF_X1 U7603 ( .A(n9821), .Z(n15120) );
  INV_X1 U7604 ( .A(n12340), .ZN(n9249) );
  AOI22_X1 U7605 ( .A1(n8862), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n6643), .B2(
        n9496), .ZN(n8511) );
  OAI21_X1 U7606 ( .B1(SI_2_), .B2(n8527), .A(n8508), .ZN(n8507) );
  NAND2_X1 U7607 ( .A1(n8240), .A2(n8244), .ZN(n11110) );
  XNOR2_X1 U7608 ( .A(n8242), .B(n8241), .ZN(n11254) );
  INV_X2 U7609 ( .A(n11800), .ZN(n14011) );
  AND2_X1 U7610 ( .A1(n8441), .A2(n13844), .ZN(n9115) );
  NAND2_X1 U7611 ( .A1(n8244), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8242) );
  NAND2_X1 U7612 ( .A1(n13022), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7698) );
  AND2_X2 U7613 ( .A1(n9477), .A2(n10827), .ZN(n14852) );
  INV_X1 U7614 ( .A(n13844), .ZN(n8443) );
  XNOR2_X1 U7615 ( .A(n8194), .B(n8193), .ZN(n12049) );
  XNOR2_X1 U7616 ( .A(n8192), .B(n8191), .ZN(n14725) );
  CLKBUF_X1 U7617 ( .A(n14832), .Z(n6843) );
  NAND2_X1 U7618 ( .A1(n7406), .A2(n7641), .ZN(n13844) );
  XNOR2_X1 U7619 ( .A(n7925), .B(n7924), .ZN(n15417) );
  BUF_X1 U7620 ( .A(n8442), .Z(n11908) );
  XNOR2_X1 U7621 ( .A(n9257), .B(P1_IR_REG_30__SCAN_IN), .ZN(n9259) );
  NAND2_X1 U7622 ( .A1(n9242), .A2(n9246), .ZN(n14195) );
  MUX2_X1 U7623 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7772), .S(
        P3_IR_REG_28__SCAN_IN), .Z(n7774) );
  AND3_X2 U7624 ( .A1(n6809), .A2(n9248), .A3(n6808), .ZN(n14699) );
  OAI21_X2 U7625 ( .B1(n9248), .B2(P1_IR_REG_23__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9219) );
  NAND2_X2 U7626 ( .A1(n9192), .A2(n9469), .ZN(n8533) );
  INV_X2 U7627 ( .A(n14691), .ZN(n11910) );
  NOR2_X1 U7628 ( .A1(n8523), .A2(n8524), .ZN(n8525) );
  CLKBUF_X1 U7629 ( .A(n9256), .Z(n14689) );
  AOI21_X1 U7630 ( .B1(n8811), .B2(n8411), .A(n6736), .ZN(n14832) );
  NAND2_X1 U7631 ( .A1(n8427), .A2(n8424), .ZN(n10827) );
  NAND2_X1 U7632 ( .A1(n9256), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9257) );
  OR2_X1 U7633 ( .A1(n9247), .A2(n6810), .ZN(n6809) );
  XNOR2_X1 U7634 ( .A(n7640), .B(n8440), .ZN(n8442) );
  AOI21_X1 U7635 ( .B1(n8459), .B2(n6707), .A(n7407), .ZN(n7406) );
  NAND2_X1 U7636 ( .A1(n7641), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7640) );
  OR2_X1 U7637 ( .A1(n7930), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7944) );
  NAND2_X1 U7638 ( .A1(n7775), .A2(n7776), .ZN(n7771) );
  NAND2_X1 U7639 ( .A1(n9231), .A2(n9230), .ZN(n14696) );
  INV_X1 U7640 ( .A(n9246), .ZN(n9216) );
  AND2_X1 U7641 ( .A1(n9245), .A2(n9244), .ZN(n14010) );
  XNOR2_X1 U7642 ( .A(n7894), .B(n7893), .ZN(n10928) );
  MUX2_X1 U7643 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8457), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n8458) );
  NAND2_X1 U7644 ( .A1(n9250), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9238) );
  OR2_X1 U7645 ( .A1(n9236), .A2(n9233), .ZN(n9234) );
  NAND2_X1 U7646 ( .A1(n8439), .A2(n6713), .ZN(n7641) );
  NAND2_X1 U7647 ( .A1(n7223), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8455) );
  NAND2_X1 U7648 ( .A1(n8421), .A2(n8429), .ZN(n8427) );
  NAND2_X1 U7649 ( .A1(n8297), .A2(n6833), .ZN(n8348) );
  AND2_X1 U7650 ( .A1(n6934), .A2(n7153), .ZN(n9214) );
  NOR2_X1 U7651 ( .A1(n8720), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n8722) );
  NAND2_X1 U7652 ( .A1(n7573), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n7109) );
  NAND2_X1 U7653 ( .A1(n7571), .A2(n7779), .ZN(n7110) );
  AND2_X2 U7654 ( .A1(n9485), .A2(n9212), .ZN(n7612) );
  AND2_X1 U7655 ( .A1(n9211), .A2(n9776), .ZN(n9212) );
  AND2_X2 U7656 ( .A1(n9288), .A2(n9289), .ZN(n9210) );
  NAND2_X1 U7657 ( .A1(n8351), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n8350) );
  AND3_X1 U7658 ( .A1(n9222), .A2(n9221), .A3(n9220), .ZN(n9226) );
  INV_X4 U7659 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7660 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n7987) );
  NOR2_X1 U7661 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n7216) );
  INV_X1 U7662 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n7953) );
  INV_X1 U7663 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9776) );
  INV_X1 U7664 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n7922) );
  NOR2_X1 U7665 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n8405) );
  NOR2_X1 U7666 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n8406) );
  NOR2_X1 U7667 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n9221) );
  INV_X1 U7668 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8425) );
  INV_X4 U7669 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7670 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8429) );
  NOR2_X1 U7671 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n8413) );
  XNOR2_X1 U7672 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n8349) );
  INV_X1 U7673 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n8351) );
  NOR2_X2 U7674 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n10145) );
  OAI21_X1 U7675 ( .B1(n10672), .B2(n10673), .A(n10603), .ZN(n10605) );
  NAND2_X2 U7676 ( .A1(n10127), .A2(n9800), .ZN(n8095) );
  NAND2_X2 U7677 ( .A1(n11737), .A2(n9800), .ZN(n14025) );
  OAI21_X2 U7678 ( .B1(n11329), .B2(n7449), .A(n7447), .ZN(n12876) );
  NAND2_X2 U7679 ( .A1(n15555), .A2(n8369), .ZN(n14714) );
  AOI21_X2 U7680 ( .B1(n13679), .B2(n6741), .A(n7416), .ZN(n13646) );
  BUF_X1 U7681 ( .A(n12337), .Z(n6645) );
  BUF_X4 U7682 ( .A(n12337), .Z(n6646) );
  AOI21_X2 U7683 ( .B1(n13646), .B2(n13645), .A(n6908), .ZN(n13627) );
  NOR2_X2 U7684 ( .A1(n13790), .A2(n13656), .ZN(n13641) );
  XNOR2_X2 U7685 ( .A(n8304), .B(n7282), .ZN(n8344) );
  NAND2_X2 U7686 ( .A1(n7283), .A2(n8303), .ZN(n8304) );
  INV_X1 U7687 ( .A(n9821), .ZN(n6647) );
  INV_X1 U7688 ( .A(n9821), .ZN(n15161) );
  NOR2_X1 U7689 ( .A1(n10059), .A2(n14010), .ZN(n9821) );
  NAND2_X1 U7690 ( .A1(n11737), .A2(n6832), .ZN(n11759) );
  AOI21_X2 U7691 ( .B1(n9883), .B2(P1_REG1_REG_6__SCAN_IN), .A(n9877), .ZN(
        n9892) );
  NAND2_X2 U7692 ( .A1(n9265), .A2(n9266), .ZN(n11737) );
  OAI21_X2 U7693 ( .B1(n8128), .B2(n7456), .A(n7454), .ZN(n12696) );
  AND2_X2 U7694 ( .A1(n6853), .A2(n6852), .ZN(n14727) );
  NOR2_X2 U7695 ( .A1(n10544), .A2(n10545), .ZN(n10543) );
  AOI21_X2 U7696 ( .B1(n15067), .B2(P1_REG1_REG_16__SCAN_IN), .A(n15058), .ZN(
        n15077) );
  AOI21_X2 U7697 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n14343), .A(n15076), .ZN(
        n14344) );
  NOR2_X2 U7698 ( .A1(n15077), .A2(n15078), .ZN(n15076) );
  OAI211_X1 U7699 ( .C1(n6845), .C2(n11619), .A(n9939), .B(n9938), .ZN(n15118)
         );
  NAND2_X1 U7700 ( .A1(n6686), .A2(n7107), .ZN(n7106) );
  NOR2_X1 U7701 ( .A1(n7693), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n7107) );
  BUF_X1 U7702 ( .A(n8070), .Z(n6916) );
  NAND2_X1 U7703 ( .A1(n7009), .A2(n7008), .ZN(n7338) );
  INV_X1 U7704 ( .A(n12602), .ZN(n7008) );
  INV_X1 U7705 ( .A(n6997), .ZN(n12638) );
  NAND2_X1 U7706 ( .A1(n11788), .A2(n11787), .ZN(n14372) );
  OAI21_X1 U7707 ( .B1(n7399), .B2(n6956), .A(n11744), .ZN(n6955) );
  AND3_X1 U7708 ( .A1(n14469), .A2(n14514), .A3(n7401), .ZN(n6954) );
  OR2_X1 U7709 ( .A1(n8542), .A2(n8541), .ZN(n7670) );
  NAND2_X1 U7710 ( .A1(n6797), .A2(n6795), .ZN(n7058) );
  INV_X1 U7711 ( .A(n6796), .ZN(n6795) );
  NAND2_X1 U7712 ( .A1(n7646), .A2(n7645), .ZN(n7644) );
  INV_X1 U7713 ( .A(n8921), .ZN(n7645) );
  INV_X1 U7714 ( .A(n8922), .ZN(n7646) );
  INV_X1 U7715 ( .A(n14190), .ZN(n7120) );
  NAND2_X1 U7716 ( .A1(n14185), .A2(n7560), .ZN(n7559) );
  INV_X1 U7717 ( .A(n7088), .ZN(n7087) );
  AOI21_X1 U7718 ( .B1(n13569), .B2(n9102), .A(n9120), .ZN(n9140) );
  NAND2_X1 U7719 ( .A1(n9131), .A2(n9029), .ZN(n9126) );
  AND2_X1 U7720 ( .A1(n9036), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n9018) );
  XNOR2_X1 U7721 ( .A(n10089), .B(n9998), .ZN(n9996) );
  INV_X1 U7722 ( .A(n7800), .ZN(n7932) );
  INV_X1 U7723 ( .A(n13027), .ZN(n7705) );
  NOR2_X1 U7724 ( .A1(n10310), .A2(n7341), .ZN(n10164) );
  NOR2_X1 U7725 ( .A1(n6641), .A2(n10162), .ZN(n7341) );
  AOI21_X1 U7726 ( .B1(n6985), .B2(n6984), .A(n6983), .ZN(n11893) );
  NOR2_X1 U7727 ( .A1(n11282), .A2(n14784), .ZN(n6983) );
  INV_X1 U7728 ( .A(n11890), .ZN(n6984) );
  OR2_X1 U7729 ( .A1(n12205), .A2(n12536), .ZN(n12176) );
  NOR2_X1 U7730 ( .A1(n8138), .A2(n7462), .ZN(n7461) );
  INV_X1 U7731 ( .A(n8127), .ZN(n7462) );
  OR2_X1 U7732 ( .A1(n12483), .A2(n12743), .ZN(n7460) );
  NOR2_X1 U7733 ( .A1(n12725), .A2(n12154), .ZN(n7094) );
  AND2_X1 U7734 ( .A1(n12759), .A2(n12758), .ZN(n12768) );
  OR2_X1 U7735 ( .A1(n12997), .A2(n12784), .ZN(n12137) );
  XNOR2_X1 U7736 ( .A(n15462), .B(n15442), .ZN(n8206) );
  INV_X1 U7737 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n7694) );
  INV_X1 U7738 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8005) );
  NAND2_X1 U7739 ( .A1(n11944), .A2(n11943), .ZN(n11948) );
  NAND2_X1 U7740 ( .A1(n7237), .A2(n13507), .ZN(n7236) );
  INV_X1 U7741 ( .A(n13767), .ZN(n7237) );
  NOR2_X1 U7742 ( .A1(n13645), .A2(n7264), .ZN(n7263) );
  INV_X1 U7743 ( .A(n7265), .ZN(n7264) );
  OR2_X1 U7744 ( .A1(n14830), .A2(n14849), .ZN(n7328) );
  NAND2_X1 U7745 ( .A1(n8533), .A2(n9800), .ZN(n8502) );
  INV_X1 U7746 ( .A(n7321), .ZN(n13584) );
  NAND2_X1 U7747 ( .A1(n7269), .A2(n13513), .ZN(n7268) );
  AND2_X1 U7748 ( .A1(n8555), .A2(n8437), .ZN(n7409) );
  NAND2_X1 U7749 ( .A1(n11036), .A2(n11035), .ZN(n7143) );
  NAND2_X1 U7750 ( .A1(n9831), .A2(n14008), .ZN(n10525) );
  NOR2_X1 U7751 ( .A1(n11036), .A2(n11035), .ZN(n7142) );
  OR2_X1 U7752 ( .A1(n14384), .A2(n14608), .ZN(n7213) );
  NAND2_X1 U7753 ( .A1(n14448), .A2(n12305), .ZN(n7379) );
  OR2_X1 U7754 ( .A1(n14667), .A2(n14530), .ZN(n14147) );
  OR2_X1 U7755 ( .A1(n14938), .A2(n12218), .ZN(n7605) );
  OR2_X1 U7756 ( .A1(n11381), .A2(n7611), .ZN(n7606) );
  OAI21_X1 U7757 ( .B1(n10807), .B2(n10806), .A(n10808), .ZN(n10870) );
  NAND2_X1 U7758 ( .A1(n7594), .A2(n7610), .ZN(n7593) );
  INV_X1 U7759 ( .A(n7601), .ZN(n7594) );
  AOI21_X1 U7760 ( .B1(n7603), .B2(n7602), .A(n14730), .ZN(n7601) );
  INV_X1 U7761 ( .A(n7607), .ZN(n7602) );
  NAND2_X1 U7762 ( .A1(n8992), .A2(n7039), .ZN(n9015) );
  OAI21_X1 U7763 ( .B1(n9032), .B2(n11304), .A(n9030), .ZN(n7039) );
  OAI21_X1 U7764 ( .B1(n9051), .B2(n9050), .A(n8990), .ZN(n9032) );
  AND2_X1 U7765 ( .A1(n8881), .A2(n8861), .ZN(n8879) );
  OAI21_X1 U7766 ( .B1(n7038), .B2(n6773), .A(n8858), .ZN(n8880) );
  INV_X1 U7767 ( .A(n7124), .ZN(n7038) );
  AND2_X2 U7768 ( .A1(n9208), .A2(n9213), .ZN(n7151) );
  INV_X1 U7769 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9211) );
  OAI211_X1 U7770 ( .C1(n8769), .C2(n6738), .A(n8809), .B(n7029), .ZN(n8834)
         );
  AOI21_X1 U7771 ( .B1(n6971), .B2(n6970), .A(n6731), .ZN(n6969) );
  INV_X1 U7772 ( .A(n6975), .ZN(n6970) );
  NAND2_X1 U7773 ( .A1(n8671), .A2(n8655), .ZN(n8672) );
  OR2_X1 U7774 ( .A1(n8694), .A2(n8689), .ZN(n8655) );
  NAND2_X1 U7775 ( .A1(n7037), .A2(n6705), .ZN(n8606) );
  NAND2_X1 U7776 ( .A1(n8565), .A2(n7117), .ZN(n7037) );
  NAND2_X1 U7777 ( .A1(n7117), .A2(n7118), .ZN(n7115) );
  NAND2_X1 U7778 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n7274), .ZN(n7273) );
  NOR2_X1 U7779 ( .A1(n12392), .A2(n12712), .ZN(n7169) );
  NAND2_X1 U7780 ( .A1(n7162), .A2(n7160), .ZN(n7159) );
  NAND2_X1 U7781 ( .A1(n7163), .A2(n7168), .ZN(n7162) );
  NAND2_X1 U7782 ( .A1(n7161), .A2(n7164), .ZN(n7160) );
  NAND2_X1 U7783 ( .A1(n7164), .A2(n7170), .ZN(n7163) );
  INV_X1 U7784 ( .A(n10844), .ZN(n7190) );
  NOR2_X1 U7785 ( .A1(n12656), .A2(n7307), .ZN(n7306) );
  NOR2_X1 U7786 ( .A1(n10930), .A2(n11301), .ZN(n11256) );
  NAND2_X1 U7787 ( .A1(n7363), .A2(n7362), .ZN(n7012) );
  INV_X1 U7788 ( .A(n15423), .ZN(n7362) );
  NOR2_X1 U7789 ( .A1(n11321), .A2(n14806), .ZN(n11320) );
  NAND2_X1 U7790 ( .A1(n7334), .A2(n7333), .ZN(n7332) );
  INV_X1 U7791 ( .A(n12568), .ZN(n7333) );
  XNOR2_X1 U7792 ( .A(n11858), .B(n11896), .ZN(n12587) );
  NOR2_X1 U7793 ( .A1(n12587), .A2(n12955), .ZN(n12586) );
  NAND2_X1 U7794 ( .A1(n8213), .A2(n12096), .ZN(n11445) );
  NOR2_X1 U7795 ( .A1(n12088), .A2(n7473), .ZN(n7472) );
  INV_X1 U7796 ( .A(n7899), .ZN(n7473) );
  INV_X1 U7797 ( .A(n15448), .ZN(n15461) );
  INV_X1 U7798 ( .A(n8095), .ZN(n11998) );
  INV_X1 U7799 ( .A(n10127), .ZN(n8072) );
  INV_X1 U7800 ( .A(n7763), .ZN(n6800) );
  XNOR2_X1 U7801 ( .A(n8071), .B(P3_IR_REG_19__SCAN_IN), .ZN(n12014) );
  NAND2_X1 U7802 ( .A1(n7749), .A2(n7748), .ZN(n8049) );
  AND2_X1 U7803 ( .A1(n7745), .A2(n7744), .ZN(n8019) );
  NOR2_X1 U7804 ( .A1(n8003), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n8006) );
  AND2_X1 U7805 ( .A1(n8006), .A2(n8005), .ZN(n8036) );
  AND2_X1 U7806 ( .A1(n7514), .A2(n7510), .ZN(n7508) );
  AND2_X1 U7807 ( .A1(n13790), .A2(n13511), .ZN(n6908) );
  XNOR2_X1 U7808 ( .A(n13790), .B(n13398), .ZN(n13645) );
  AOI21_X1 U7809 ( .B1(n7421), .B2(n13686), .A(n7423), .ZN(n7419) );
  AND2_X1 U7810 ( .A1(n13800), .A2(n13513), .ZN(n7423) );
  NAND2_X1 U7811 ( .A1(n6911), .A2(n6850), .ZN(n7422) );
  AND2_X1 U7812 ( .A1(n13804), .A2(n11822), .ZN(n6849) );
  AOI21_X1 U7813 ( .B1(n7249), .B2(n7247), .A(n6696), .ZN(n7246) );
  INV_X1 U7814 ( .A(n11814), .ZN(n7247) );
  AOI21_X1 U7815 ( .B1(n7257), .B2(n11574), .A(n6690), .ZN(n7255) );
  AND2_X2 U7816 ( .A1(n11909), .A2(n11621), .ZN(n11715) );
  XNOR2_X1 U7817 ( .A(n14614), .B(n13910), .ZN(n14410) );
  NAND2_X1 U7818 ( .A1(n7379), .A2(n7375), .ZN(n7374) );
  INV_X1 U7819 ( .A(n11757), .ZN(n7375) );
  NAND2_X1 U7820 ( .A1(n7373), .A2(n7379), .ZN(n7372) );
  INV_X1 U7821 ( .A(n7376), .ZN(n7373) );
  NOR2_X1 U7822 ( .A1(n7391), .A2(n14524), .ZN(n7389) );
  NAND2_X1 U7823 ( .A1(n14534), .A2(n7208), .ZN(n7207) );
  OAI21_X1 U7824 ( .B1(n11540), .B2(n11539), .A(n14118), .ZN(n11541) );
  INV_X1 U7825 ( .A(n6648), .ZN(n11700) );
  INV_X1 U7826 ( .A(n6845), .ZN(n11699) );
  NAND2_X1 U7827 ( .A1(n11416), .A2(n7387), .ZN(n7385) );
  INV_X1 U7828 ( .A(n7388), .ZN(n7387) );
  OAI21_X1 U7829 ( .B1(n14938), .B2(n14270), .A(n11415), .ZN(n7388) );
  BUF_X1 U7830 ( .A(n11737), .Z(n6845) );
  INV_X1 U7831 ( .A(n14025), .ZN(n14017) );
  NAND2_X1 U7832 ( .A1(n11792), .A2(n11791), .ZN(n14597) );
  OAI22_X1 U7833 ( .A1(n14372), .A2(n11789), .B1(n12339), .B2(n14384), .ZN(
        n11790) );
  XNOR2_X1 U7834 ( .A(n9069), .B(n9068), .ZN(n11809) );
  OAI21_X1 U7835 ( .B1(n9015), .B2(n8993), .A(n8994), .ZN(n9069) );
  XNOR2_X1 U7836 ( .A(n8949), .B(SI_22_), .ZN(n11735) );
  NAND2_X1 U7837 ( .A1(n7124), .A2(n7125), .ZN(n8856) );
  INV_X1 U7838 ( .A(n8490), .ZN(n6945) );
  AND2_X1 U7839 ( .A1(n7361), .A2(n7360), .ZN(n11854) );
  INV_X1 U7840 ( .A(n11261), .ZN(n7360) );
  NOR2_X1 U7841 ( .A1(n12552), .A2(n14798), .ZN(n12551) );
  OR2_X1 U7842 ( .A1(n12620), .A2(n11862), .ZN(n6997) );
  INV_X1 U7843 ( .A(n7336), .ZN(n11861) );
  XNOR2_X1 U7844 ( .A(n6961), .B(n6960), .ZN(n14598) );
  NAND2_X1 U7845 ( .A1(n6963), .A2(n6962), .ZN(n6961) );
  NAND2_X1 U7846 ( .A1(n14384), .A2(n14262), .ZN(n6962) );
  NAND2_X1 U7847 ( .A1(n6931), .A2(n6856), .ZN(n6930) );
  NAND2_X1 U7848 ( .A1(n8392), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n6931) );
  INV_X1 U7849 ( .A(n8561), .ZN(n7051) );
  NAND2_X1 U7850 ( .A1(n8583), .A2(n6793), .ZN(n7660) );
  INV_X1 U7851 ( .A(n14102), .ZN(n6888) );
  AOI21_X1 U7852 ( .B1(n6655), .B2(n7066), .A(n6737), .ZN(n7064) );
  INV_X1 U7853 ( .A(n14125), .ZN(n7543) );
  AOI21_X1 U7854 ( .B1(n15460), .B2(n12049), .A(n12048), .ZN(n12055) );
  NAND2_X1 U7855 ( .A1(n6728), .A2(n7652), .ZN(n7651) );
  NOR2_X1 U7856 ( .A1(n6722), .A2(n7060), .ZN(n7059) );
  NAND2_X1 U7857 ( .A1(n6730), .A2(n8786), .ZN(n7661) );
  NAND2_X1 U7858 ( .A1(n14157), .A2(n14159), .ZN(n7546) );
  AOI21_X1 U7859 ( .B1(n12171), .B2(n12124), .A(n12123), .ZN(n12129) );
  AND2_X1 U7860 ( .A1(n8921), .A2(n8922), .ZN(n7647) );
  OAI211_X1 U7861 ( .C1(n8878), .C2(n7668), .A(n7665), .B(n8900), .ZN(n8901)
         );
  NOR2_X1 U7862 ( .A1(n12151), .A2(n12152), .ZN(n6920) );
  NAND2_X1 U7863 ( .A1(n12749), .A2(n6918), .ZN(n6917) );
  NOR2_X1 U7864 ( .A1(n12728), .A2(n12161), .ZN(n6918) );
  NAND2_X1 U7865 ( .A1(n12155), .A2(n12154), .ZN(n6869) );
  AOI21_X1 U7866 ( .B1(n12978), .B2(n12743), .A(n12171), .ZN(n6868) );
  AOI21_X1 U7867 ( .B1(n8923), .B2(n7644), .A(n7642), .ZN(n7057) );
  NAND2_X1 U7868 ( .A1(n7643), .A2(n8946), .ZN(n7642) );
  NAND2_X1 U7869 ( .A1(n7647), .A2(n7644), .ZN(n7643) );
  NAND2_X1 U7870 ( .A1(n7644), .A2(n8947), .ZN(n7055) );
  INV_X1 U7871 ( .A(n8962), .ZN(n7655) );
  INV_X1 U7872 ( .A(n8961), .ZN(n7654) );
  INV_X1 U7873 ( .A(n14183), .ZN(n6816) );
  NOR2_X1 U7874 ( .A1(n8950), .A2(n8964), .ZN(n7032) );
  OR2_X1 U7875 ( .A1(n12985), .A2(n12442), .ZN(n12148) );
  NOR2_X1 U7876 ( .A1(n7470), .A2(n8018), .ZN(n7469) );
  INV_X1 U7877 ( .A(n7997), .ZN(n7470) );
  INV_X1 U7878 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8452) );
  NAND2_X1 U7879 ( .A1(n14192), .A2(n7535), .ZN(n7534) );
  OAI21_X1 U7880 ( .B1(n14189), .B2(n14188), .A(n6735), .ZN(n7121) );
  INV_X1 U7881 ( .A(n8994), .ZN(n7587) );
  OAI21_X1 U7882 ( .B1(n11734), .B2(n6913), .A(n6912), .ZN(n8554) );
  NAND2_X1 U7883 ( .A1(n11734), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n6912) );
  INV_X1 U7884 ( .A(n7168), .ZN(n7161) );
  INV_X1 U7885 ( .A(n10157), .ZN(n7446) );
  OR2_X1 U7886 ( .A1(n10460), .A2(n10459), .ZN(n10461) );
  NOR2_X1 U7887 ( .A1(n7354), .A2(n11864), .ZN(n7350) );
  AOI21_X1 U7888 ( .B1(n12637), .B2(n7350), .A(n7348), .ZN(n7347) );
  NOR2_X1 U7889 ( .A1(n7349), .A2(n7352), .ZN(n7348) );
  INV_X1 U7890 ( .A(n7354), .ZN(n7349) );
  INV_X1 U7891 ( .A(n7461), .ZN(n7455) );
  NAND2_X1 U7892 ( .A1(n12741), .A2(n12152), .ZN(n8128) );
  OR2_X1 U7894 ( .A1(n12788), .A2(n12799), .ZN(n12134) );
  INV_X1 U7895 ( .A(n7469), .ZN(n7464) );
  INV_X1 U7896 ( .A(n8017), .ZN(n7467) );
  OR2_X1 U7897 ( .A1(n11999), .A2(n9322), .ZN(n7788) );
  INV_X1 U7898 ( .A(n6915), .ZN(n6914) );
  OAI22_X1 U7899 ( .A1(n8095), .A2(n9323), .B1(n10127), .B2(n10253), .ZN(n6915) );
  NAND2_X1 U7900 ( .A1(n8166), .A2(n8165), .ZN(n12396) );
  OR2_X2 U7901 ( .A1(n14725), .A2(n12049), .ZN(n12161) );
  INV_X1 U7902 ( .A(n7758), .ZN(n7300) );
  AND2_X1 U7903 ( .A1(n6916), .A2(n7200), .ZN(n8265) );
  AND2_X1 U7904 ( .A1(n6658), .A2(n6749), .ZN(n7200) );
  INV_X1 U7905 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n13256) );
  NAND2_X1 U7906 ( .A1(n7288), .A2(n7286), .ZN(n7754) );
  AOI21_X1 U7907 ( .B1(n7289), .B2(n7291), .A(n7287), .ZN(n7286) );
  INV_X1 U7908 ( .A(n7753), .ZN(n7287) );
  INV_X1 U7909 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n7688) );
  INV_X1 U7910 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7695) );
  OR2_X1 U7911 ( .A1(n7528), .A2(n11914), .ZN(n7527) );
  AND2_X1 U7912 ( .A1(n11916), .A2(n11915), .ZN(n7528) );
  AND2_X1 U7913 ( .A1(n6745), .A2(n7482), .ZN(n7481) );
  NAND2_X1 U7914 ( .A1(n7483), .A2(n7486), .ZN(n7482) );
  INV_X1 U7915 ( .A(n13463), .ZN(n7491) );
  AOI21_X1 U7916 ( .B1(n13482), .B2(n7494), .A(n6781), .ZN(n7487) );
  NAND2_X1 U7917 ( .A1(n6729), .A2(n9138), .ZN(n7589) );
  AND2_X1 U7918 ( .A1(n9001), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n9036) );
  NOR2_X1 U7919 ( .A1(n7248), .A2(n7245), .ZN(n7244) );
  INV_X1 U7920 ( .A(n11584), .ZN(n7245) );
  INV_X1 U7921 ( .A(n7249), .ZN(n7248) );
  NOR2_X1 U7922 ( .A1(n11580), .A2(n7258), .ZN(n7257) );
  INV_X1 U7923 ( .A(n11578), .ZN(n7258) );
  OAI21_X1 U7924 ( .B1(n10727), .B2(n7415), .A(n10995), .ZN(n7414) );
  INV_X1 U7925 ( .A(n10764), .ZN(n7415) );
  AND2_X1 U7926 ( .A1(n10289), .A2(n10236), .ZN(n7238) );
  INV_X1 U7927 ( .A(n10240), .ZN(n7241) );
  AND2_X1 U7928 ( .A1(n9571), .A2(n10899), .ZN(n9477) );
  INV_X1 U7929 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8438) );
  NAND2_X1 U7930 ( .A1(n8453), .A2(n8452), .ZN(n7225) );
  INV_X1 U7931 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8430) );
  INV_X1 U7932 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n8404) );
  INV_X1 U7933 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8403) );
  NAND2_X1 U7934 ( .A1(n7212), .A2(n14593), .ZN(n7211) );
  INV_X1 U7935 ( .A(n7213), .ZN(n7212) );
  NOR2_X1 U7936 ( .A1(n14667), .A2(n14565), .ZN(n7208) );
  INV_X1 U7937 ( .A(n14237), .ZN(n7633) );
  INV_X1 U7938 ( .A(n7624), .ZN(n7623) );
  NAND2_X1 U7939 ( .A1(n14091), .A2(n7625), .ZN(n7624) );
  INV_X1 U7940 ( .A(n11085), .ZN(n7625) );
  NAND2_X1 U7941 ( .A1(n14050), .A2(n14049), .ZN(n14047) );
  NAND2_X1 U7942 ( .A1(n14570), .A2(n14123), .ZN(n7634) );
  NAND2_X1 U7943 ( .A1(n15106), .A2(n15108), .ZN(n9941) );
  OAI21_X1 U7944 ( .B1(n8983), .B2(n7122), .A(n8986), .ZN(n9051) );
  INV_X1 U7945 ( .A(n8984), .ZN(n7122) );
  OAI21_X1 U7946 ( .B1(n8880), .B2(n6657), .A(n7111), .ZN(n8949) );
  INV_X1 U7947 ( .A(n7112), .ZN(n7111) );
  OAI21_X1 U7948 ( .B1(n6657), .B2(n8879), .A(n8929), .ZN(n7112) );
  NOR2_X1 U7949 ( .A1(n7568), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n7566) );
  NAND2_X1 U7950 ( .A1(n7570), .A2(n7569), .ZN(n7568) );
  NOR2_X1 U7951 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n7569) );
  NOR2_X1 U7952 ( .A1(n7579), .A2(n8766), .ZN(n7578) );
  OAI21_X1 U7953 ( .B1(n7579), .B2(n7577), .A(n8790), .ZN(n7576) );
  NAND2_X1 U7954 ( .A1(n8767), .A2(n9377), .ZN(n7577) );
  INV_X1 U7955 ( .A(n8787), .ZN(n7579) );
  NAND2_X1 U7956 ( .A1(n8693), .A2(n7574), .ZN(n6974) );
  NOR2_X1 U7957 ( .A1(n8696), .A2(n6719), .ZN(n6975) );
  INV_X1 U7958 ( .A(n8566), .ZN(n7118) );
  AND3_X1 U7959 ( .A1(n6949), .A2(n6951), .A3(n6947), .ZN(n8565) );
  NAND2_X1 U7960 ( .A1(n8530), .A2(n8553), .ZN(n6951) );
  OAI21_X1 U7961 ( .B1(n11734), .B2(n7036), .A(n7035), .ZN(n7034) );
  NAND2_X1 U7962 ( .A1(n11734), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7035) );
  OAI21_X1 U7963 ( .B1(n7034), .B2(SI_3_), .A(n8528), .ZN(n8524) );
  INV_X1 U7964 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n7284) );
  INV_X1 U7965 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n7282) );
  INV_X1 U7966 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n13266) );
  OAI21_X1 U7967 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n11280), .A(n8320), .ZN(
        n8378) );
  OAI21_X1 U7968 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n8324), .A(n8323), .ZN(
        n8336) );
  AND2_X1 U7970 ( .A1(n8167), .A2(n12393), .ZN(n8169) );
  NOR2_X1 U7971 ( .A1(n7179), .A2(n7175), .ZN(n7174) );
  INV_X1 U7972 ( .A(n12467), .ZN(n7175) );
  INV_X1 U7973 ( .A(n12505), .ZN(n7179) );
  NAND2_X1 U7974 ( .A1(n12505), .A2(n7178), .ZN(n7177) );
  INV_X1 U7975 ( .A(n12368), .ZN(n7178) );
  INV_X1 U7976 ( .A(n12441), .ZN(n7188) );
  NAND2_X1 U7977 ( .A1(n10833), .A2(n7193), .ZN(n7192) );
  INV_X1 U7978 ( .A(n10472), .ZN(n7193) );
  NAND2_X1 U7979 ( .A1(n12015), .A2(n12013), .ZN(n7096) );
  NAND2_X1 U7980 ( .A1(n6862), .A2(n15444), .ZN(n6861) );
  NAND2_X1 U7981 ( .A1(n6863), .A2(n7097), .ZN(n6862) );
  NAND2_X1 U7982 ( .A1(n12181), .A2(n12180), .ZN(n6863) );
  NOR2_X1 U7983 ( .A1(n12179), .A2(n6804), .ZN(n12040) );
  NAND2_X1 U7984 ( .A1(n8264), .A2(n8263), .ZN(n9984) );
  XNOR2_X1 U7985 ( .A(n10164), .B(n10150), .ZN(n10436) );
  NAND2_X1 U7986 ( .A1(n10165), .A2(n10431), .ZN(n7339) );
  OAI22_X1 U7987 ( .A1(n10436), .A2(n7006), .B1(n7339), .B2(n10400), .ZN(
        n10399) );
  OR2_X1 U7988 ( .A1(n10400), .A2(n15532), .ZN(n7006) );
  XNOR2_X1 U7989 ( .A(n10169), .B(n10168), .ZN(n10420) );
  NAND2_X1 U7990 ( .A1(n7446), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7445) );
  NAND2_X1 U7991 ( .A1(n10155), .A2(n7446), .ZN(n7444) );
  NOR2_X1 U7992 ( .A1(n10416), .A2(n10417), .ZN(n10415) );
  OR2_X1 U7993 ( .A1(n10461), .A2(n10502), .ZN(n7358) );
  NAND2_X1 U7994 ( .A1(n7004), .A2(n10497), .ZN(n7003) );
  NAND2_X1 U7995 ( .A1(n7358), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n7004) );
  OR2_X1 U7996 ( .A1(n11256), .A2(n11257), .ZN(n7363) );
  AND2_X1 U7997 ( .A1(n15417), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7437) );
  AND4_X1 U7998 ( .A1(n7709), .A2(n7708), .A3(n7707), .A4(n7706), .ZN(n12683)
         );
  NAND2_X1 U7999 ( .A1(n8162), .A2(n8161), .ZN(n12679) );
  NOR2_X1 U8000 ( .A1(n12708), .A2(n7458), .ZN(n7457) );
  INV_X1 U8001 ( .A(n7460), .ZN(n7458) );
  NAND2_X1 U8002 ( .A1(n6846), .A2(n7461), .ZN(n7459) );
  OAI21_X1 U8003 ( .B1(n12790), .B2(n7102), .A(n7100), .ZN(n12737) );
  INV_X1 U8004 ( .A(n7101), .ZN(n7100) );
  OAI21_X1 U8005 ( .B1(n7102), .B2(n12134), .A(n8225), .ZN(n7101) );
  NAND2_X1 U8006 ( .A1(n8223), .A2(n7103), .ZN(n7102) );
  OR2_X1 U8007 ( .A1(n12989), .A2(n12755), .ZN(n12759) );
  AND2_X1 U8008 ( .A1(n8104), .A2(n8090), .ZN(n7477) );
  NOR2_X1 U8009 ( .A1(n8220), .A2(n7089), .ZN(n7088) );
  INV_X1 U8010 ( .A(n12125), .ZN(n7089) );
  AND2_X1 U8011 ( .A1(n12811), .A2(n8064), .ZN(n12798) );
  AND2_X1 U8012 ( .A1(n12041), .A2(n12120), .ZN(n12863) );
  AOI21_X1 U8013 ( .B1(n7450), .B2(n7448), .A(n6718), .ZN(n7447) );
  INV_X1 U8014 ( .A(n7450), .ZN(n7449) );
  INV_X1 U8015 ( .A(n7962), .ZN(n7448) );
  AND2_X1 U8016 ( .A1(n7975), .A2(n7974), .ZN(n14764) );
  AND4_X1 U8017 ( .A1(n7919), .A2(n7918), .A3(n7917), .A4(n7916), .ZN(n11443)
         );
  AOI21_X1 U8018 ( .B1(n6682), .B2(n7079), .A(n7075), .ZN(n7074) );
  INV_X1 U8019 ( .A(n12080), .ZN(n7075) );
  AND4_X1 U8020 ( .A1(n7859), .A2(n7858), .A3(n7857), .A4(n7856), .ZN(n10947)
         );
  AND4_X1 U8021 ( .A1(n7892), .A2(n7891), .A3(n7890), .A4(n7889), .ZN(n11142)
         );
  NAND2_X1 U8022 ( .A1(n12080), .A2(n12081), .ZN(n12022) );
  NAND2_X1 U8023 ( .A1(n10957), .A2(n12018), .ZN(n10959) );
  NAND2_X1 U8024 ( .A1(n10376), .A2(n12061), .ZN(n10379) );
  NAND2_X1 U8025 ( .A1(n10017), .A2(n12171), .ZN(n15450) );
  AND2_X1 U8026 ( .A1(n8235), .A2(n8270), .ZN(n15470) );
  NAND2_X1 U8027 ( .A1(n7308), .A2(n12000), .ZN(n12013) );
  NAND2_X1 U8028 ( .A1(n7781), .A2(n7780), .ZN(n12671) );
  NAND2_X1 U8029 ( .A1(n14725), .A2(n12049), .ZN(n15521) );
  OAI21_X1 U8030 ( .B1(n9388), .B2(P3_D_REG_0__SCAN_IN), .A(n8247), .ZN(n7154)
         );
  AND2_X1 U8031 ( .A1(n10125), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9387) );
  NOR2_X2 U8032 ( .A1(n7771), .A2(P3_IR_REG_28__SCAN_IN), .ZN(n7699) );
  OR2_X1 U8033 ( .A1(n11987), .A2(n11986), .ZN(n11995) );
  AOI21_X1 U8034 ( .B1(n7304), .B2(n7767), .A(n6791), .ZN(n7303) );
  NAND2_X1 U8035 ( .A1(n7762), .A2(n7761), .ZN(n7763) );
  OR2_X1 U8036 ( .A1(n7754), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7755) );
  NAND2_X1 U8037 ( .A1(n8081), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7756) );
  AND2_X1 U8038 ( .A1(n8197), .A2(n8237), .ZN(n8283) );
  NAND2_X1 U8039 ( .A1(n6916), .A2(n7694), .ZN(n8195) );
  XNOR2_X1 U8040 ( .A(n7754), .B(n10829), .ZN(n8081) );
  AND2_X1 U8041 ( .A1(n7753), .A2(n7752), .ZN(n8065) );
  INV_X1 U8042 ( .A(n7290), .ZN(n7289) );
  OAI21_X1 U8043 ( .B1(n8048), .B2(n7291), .A(n8065), .ZN(n7290) );
  INV_X1 U8044 ( .A(n7751), .ZN(n7291) );
  NAND2_X1 U8045 ( .A1(n8049), .A2(n8048), .ZN(n8051) );
  INV_X1 U8046 ( .A(n7296), .ZN(n7295) );
  OAI21_X1 U8047 ( .B1(n7999), .B2(n7297), .A(n8019), .ZN(n7296) );
  NAND2_X1 U8048 ( .A1(n8000), .A2(n7999), .ZN(n8002) );
  OR2_X1 U8049 ( .A1(n7986), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n8003) );
  NAND2_X1 U8050 ( .A1(n7731), .A2(n7730), .ZN(n7921) );
  OAI21_X1 U8051 ( .B1(n7864), .B2(n7721), .A(n7722), .ZN(n7876) );
  AND2_X1 U8052 ( .A1(n9350), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n7721) );
  INV_X1 U8054 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7686) );
  INV_X1 U8055 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n7479) );
  INV_X1 U8056 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7196) );
  XNOR2_X1 U8057 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n7845) );
  XNOR2_X1 U8058 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n7815) );
  NAND2_X1 U8059 ( .A1(n11928), .A2(n7495), .ZN(n7494) );
  INV_X1 U8060 ( .A(n11929), .ZN(n7495) );
  INV_X1 U8061 ( .A(n13385), .ZN(n7510) );
  AOI21_X1 U8062 ( .B1(n7513), .B2(n13419), .A(n7512), .ZN(n7511) );
  INV_X1 U8063 ( .A(n11960), .ZN(n7512) );
  OR2_X1 U8064 ( .A1(n6740), .A2(n7501), .ZN(n7497) );
  NAND2_X1 U8065 ( .A1(n7531), .A2(n13449), .ZN(n13448) );
  INV_X1 U8066 ( .A(n7532), .ZN(n7531) );
  NAND2_X1 U8067 ( .A1(n7530), .A2(n13450), .ZN(n13453) );
  INV_X1 U8068 ( .A(n11956), .ZN(n7515) );
  NAND2_X1 U8070 ( .A1(n9081), .A2(n9080), .ZN(n13566) );
  OAI21_X1 U8071 ( .B1(n14026), .B2(n9109), .A(n9111), .ZN(n13569) );
  AND2_X1 U8072 ( .A1(n7234), .A2(n11846), .ZN(n7227) );
  NAND2_X1 U8073 ( .A1(n7233), .A2(n7236), .ZN(n7232) );
  INV_X1 U8074 ( .A(n11846), .ZN(n7233) );
  INV_X1 U8075 ( .A(n7229), .ZN(n7228) );
  OAI21_X1 U8076 ( .B1(n7234), .B2(n7232), .A(n7230), .ZN(n7229) );
  NAND2_X1 U8077 ( .A1(n7231), .A2(n11846), .ZN(n7230) );
  INV_X1 U8078 ( .A(n7236), .ZN(n7231) );
  OR2_X1 U8079 ( .A1(n13785), .A2(n13510), .ZN(n7408) );
  NOR2_X1 U8080 ( .A1(n6691), .A2(n7266), .ZN(n7265) );
  INV_X1 U8081 ( .A(n7268), .ZN(n7266) );
  INV_X1 U8082 ( .A(n7421), .ZN(n7420) );
  NOR2_X1 U8083 ( .A1(n13663), .A2(n11840), .ZN(n7421) );
  AND2_X1 U8084 ( .A1(n7422), .A2(n7424), .ZN(n13673) );
  NOR2_X1 U8085 ( .A1(n6851), .A2(n6850), .ZN(n13689) );
  NOR2_X1 U8086 ( .A1(n7327), .A2(n11923), .ZN(n7325) );
  OAI21_X1 U8087 ( .B1(n14834), .B2(n7427), .A(n7425), .ZN(n11833) );
  INV_X1 U8088 ( .A(n7426), .ZN(n7425) );
  OAI21_X1 U8089 ( .B1(n7428), .B2(n7427), .A(n11585), .ZN(n7426) );
  INV_X1 U8090 ( .A(n11572), .ZN(n7427) );
  NAND2_X1 U8091 ( .A1(n13742), .A2(n11584), .ZN(n11815) );
  AND2_X1 U8092 ( .A1(n11571), .A2(n11570), .ZN(n7428) );
  NOR2_X1 U8093 ( .A1(n14850), .A2(n14849), .ZN(n14851) );
  NAND2_X1 U8094 ( .A1(n11011), .A2(n10990), .ZN(n11576) );
  NAND2_X1 U8095 ( .A1(n10757), .A2(n10756), .ZN(n10759) );
  NAND2_X1 U8096 ( .A1(n10728), .A2(n10727), .ZN(n10765) );
  NAND2_X1 U8097 ( .A1(n10237), .A2(n10236), .ZN(n7242) );
  NAND2_X1 U8098 ( .A1(n9565), .A2(n9564), .ZN(n14841) );
  NAND2_X1 U8099 ( .A1(n8968), .A2(n8967), .ZN(n13790) );
  NAND2_X1 U8100 ( .A1(n8702), .A2(n8701), .ZN(n11238) );
  AND2_X1 U8101 ( .A1(n15342), .A2(n15372), .ZN(n15350) );
  AND2_X1 U8102 ( .A1(n9477), .A2(n9476), .ZN(n15368) );
  OAI21_X1 U8103 ( .B1(n9152), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9154) );
  AND2_X1 U8104 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n8411) );
  NOR2_X1 U8105 ( .A1(n8419), .A2(n8418), .ZN(n8420) );
  INV_X1 U8106 ( .A(n11205), .ZN(n6925) );
  NAND2_X1 U8107 ( .A1(n11032), .A2(n7143), .ZN(n7140) );
  INV_X1 U8108 ( .A(n7142), .ZN(n7141) );
  NAND2_X1 U8109 ( .A1(n14917), .A2(n12254), .ZN(n13915) );
  NAND2_X1 U8110 ( .A1(n12229), .A2(n12230), .ZN(n7150) );
  NOR2_X1 U8111 ( .A1(n7149), .A2(n13898), .ZN(n7148) );
  INV_X1 U8112 ( .A(n12227), .ZN(n7149) );
  INV_X1 U8113 ( .A(n13941), .ZN(n6935) );
  INV_X1 U8114 ( .A(n14281), .ZN(n10072) );
  INV_X1 U8115 ( .A(n7139), .ZN(n7138) );
  AOI21_X1 U8116 ( .B1(n7139), .B2(n7137), .A(n7136), .ZN(n7135) );
  NOR2_X1 U8117 ( .A1(n7142), .A2(n11061), .ZN(n7139) );
  AND2_X1 U8118 ( .A1(n7133), .A2(n13907), .ZN(n7132) );
  OR2_X1 U8119 ( .A1(n13923), .A2(n7134), .ZN(n7133) );
  INV_X1 U8120 ( .A(n12313), .ZN(n7134) );
  NAND2_X1 U8121 ( .A1(n11775), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9945) );
  NOR2_X1 U8122 ( .A1(n10040), .A2(n7021), .ZN(n15008) );
  AND2_X1 U8123 ( .A1(n11072), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7021) );
  NOR2_X1 U8124 ( .A1(n15008), .A2(n15007), .ZN(n15006) );
  NOR2_X1 U8125 ( .A1(n15028), .A2(n15029), .ZN(n15027) );
  OR2_X1 U8126 ( .A1(n15062), .A2(n6786), .ZN(n7016) );
  AND2_X1 U8127 ( .A1(n7016), .A2(n7015), .ZN(n15072) );
  INV_X1 U8128 ( .A(n15074), .ZN(n7015) );
  NAND2_X1 U8129 ( .A1(n14019), .A2(n14018), .ZN(n14361) );
  AND2_X1 U8130 ( .A1(n14029), .A2(n14028), .ZN(n14366) );
  NOR2_X1 U8131 ( .A1(n14375), .A2(n14376), .ZN(n14374) );
  OAI21_X1 U8132 ( .B1(n14418), .B2(n7616), .A(n7613), .ZN(n14389) );
  AOI21_X1 U8133 ( .B1(n7615), .B2(n7614), .A(n6695), .ZN(n7613) );
  INV_X1 U8134 ( .A(n11785), .ZN(n7614) );
  XNOR2_X1 U8135 ( .A(n14608), .B(n13985), .ZN(n14398) );
  AND2_X1 U8136 ( .A1(n14416), .A2(n7370), .ZN(n7369) );
  NAND2_X1 U8137 ( .A1(n14452), .A2(n7372), .ZN(n7371) );
  NAND2_X1 U8138 ( .A1(n7372), .A2(n7374), .ZN(n7370) );
  NOR2_X1 U8139 ( .A1(n14440), .A2(n7377), .ZN(n7376) );
  INV_X1 U8140 ( .A(n11756), .ZN(n7377) );
  OR2_X1 U8141 ( .A1(n14452), .A2(n11757), .ZN(n7378) );
  NAND2_X1 U8142 ( .A1(n7630), .A2(n7629), .ZN(n14438) );
  AND2_X1 U8143 ( .A1(n14440), .A2(n11784), .ZN(n7629) );
  NAND2_X1 U8144 ( .A1(n14456), .A2(n14455), .ZN(n7630) );
  NAND2_X1 U8145 ( .A1(n14466), .A2(n7675), .ZN(n14456) );
  OR2_X1 U8146 ( .A1(n14497), .A2(n13961), .ZN(n7675) );
  OR2_X1 U8147 ( .A1(n14644), .A2(n13954), .ZN(n11783) );
  AOI21_X1 U8148 ( .B1(n7401), .B2(n14515), .A(n6721), .ZN(n7399) );
  AOI21_X1 U8149 ( .B1(n6656), .B2(n14528), .A(n6715), .ZN(n7627) );
  INV_X1 U8150 ( .A(n11684), .ZN(n7396) );
  NAND2_X1 U8151 ( .A1(n14558), .A2(n11782), .ZN(n14544) );
  OAI21_X1 U8152 ( .B1(n14965), .B2(n7404), .A(n7402), .ZN(n11674) );
  INV_X1 U8153 ( .A(n7403), .ZN(n7402) );
  NAND2_X1 U8154 ( .A1(n14965), .A2(n6676), .ZN(n11669) );
  NAND2_X1 U8155 ( .A1(n7591), .A2(n7592), .ZN(n11540) );
  AOI21_X1 U8156 ( .B1(n7597), .B2(n6654), .A(n6664), .ZN(n7592) );
  AND2_X1 U8157 ( .A1(n14119), .A2(n14118), .ZN(n14234) );
  NOR2_X1 U8158 ( .A1(n11515), .A2(n12218), .ZN(n7386) );
  NAND2_X1 U8159 ( .A1(n11074), .A2(n11073), .ZN(n14097) );
  AOI21_X1 U8160 ( .B1(n14231), .B2(n14076), .A(n6720), .ZN(n7367) );
  NAND2_X1 U8161 ( .A1(n10857), .A2(n7365), .ZN(n7366) );
  NAND2_X1 U8162 ( .A1(n7619), .A2(n10564), .ZN(n10807) );
  NAND2_X1 U8163 ( .A1(n10563), .A2(n10562), .ZN(n7619) );
  NAND2_X1 U8164 ( .A1(n10652), .A2(n14047), .ZN(n9952) );
  INV_X1 U8165 ( .A(n14533), .ZN(n14573) );
  INV_X1 U8166 ( .A(n14384), .ZN(n14600) );
  INV_X1 U8167 ( .A(n14391), .ZN(n14390) );
  NAND2_X1 U8168 ( .A1(n11748), .A2(n11747), .ZN(n14633) );
  AND2_X1 U8169 ( .A1(n9840), .A2(n10573), .ZN(n15187) );
  OR2_X1 U8170 ( .A1(n11811), .A2(P1_B_REG_SCAN_IN), .ZN(n9584) );
  AND2_X1 U8171 ( .A1(n10529), .A2(n9278), .ZN(n9846) );
  NAND2_X1 U8172 ( .A1(n9073), .A2(n9072), .ZN(n9106) );
  OR2_X1 U8173 ( .A1(n9106), .A2(n9105), .ZN(n9108) );
  NOR2_X1 U8174 ( .A1(n10118), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n6877) );
  XNOR2_X1 U8175 ( .A(n9015), .B(n9014), .ZN(n11642) );
  XNOR2_X1 U8176 ( .A(n8907), .B(n8906), .ZN(n11723) );
  AND2_X1 U8177 ( .A1(n6758), .A2(n9210), .ZN(n7152) );
  XNOR2_X1 U8178 ( .A(n8672), .B(SI_10_), .ZN(n11071) );
  NAND2_X1 U8179 ( .A1(n7034), .A2(SI_3_), .ZN(n8528) );
  NAND2_X1 U8180 ( .A1(n8526), .A2(n8525), .ZN(n6953) );
  NAND2_X1 U8181 ( .A1(n11734), .A2(n6941), .ZN(n6940) );
  NAND2_X1 U8182 ( .A1(n6946), .A2(n9322), .ZN(n8473) );
  XNOR2_X1 U8183 ( .A(n8349), .B(n8350), .ZN(n8352) );
  INV_X1 U8184 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7272) );
  INV_X1 U8185 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14310) );
  XNOR2_X1 U8186 ( .A(n8344), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n8359) );
  NOR2_X1 U8187 ( .A1(n14710), .A2(n8365), .ZN(n8367) );
  OAI21_X1 U8188 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n8312), .A(n8311), .ZN(
        n8341) );
  AND2_X1 U8189 ( .A1(n7184), .A2(n11526), .ZN(n7183) );
  NOR2_X1 U8190 ( .A1(n6663), .A2(n12520), .ZN(n7156) );
  NAND2_X1 U8191 ( .A1(n7159), .A2(n7165), .ZN(n7158) );
  NAND2_X1 U8192 ( .A1(n7166), .A2(n12417), .ZN(n7165) );
  INV_X1 U8193 ( .A(n7170), .ZN(n7166) );
  AND3_X1 U8194 ( .A1(n7912), .A2(n7911), .A3(n7910), .ZN(n10846) );
  AND4_X1 U8195 ( .A1(n7949), .A2(n7948), .A3(n7947), .A4(n7946), .ZN(n14762)
         );
  XNOR2_X1 U8196 ( .A(n12382), .B(n12380), .ZN(n12496) );
  NAND2_X1 U8197 ( .A1(n10016), .A2(n15443), .ZN(n12517) );
  INV_X1 U8198 ( .A(n12539), .ZN(n14763) );
  INV_X1 U8199 ( .A(n7010), .ZN(n11259) );
  INV_X1 U8200 ( .A(n6985), .ZN(n11891) );
  OR2_X1 U8201 ( .A1(n12551), .A2(n11856), .ZN(n7334) );
  AND2_X1 U8202 ( .A1(n7438), .A2(n6675), .ZN(n12571) );
  INV_X1 U8203 ( .A(n7332), .ZN(n12567) );
  XNOR2_X1 U8204 ( .A(n6979), .B(n11896), .ZN(n12584) );
  OR2_X1 U8205 ( .A1(n12586), .A2(n11859), .ZN(n7009) );
  INV_X1 U8206 ( .A(n7338), .ZN(n12601) );
  NOR2_X1 U8207 ( .A1(n12621), .A2(n12945), .ZN(n12620) );
  XNOR2_X1 U8208 ( .A(n6830), .B(n6829), .ZN(n11907) );
  INV_X1 U8209 ( .A(n11889), .ZN(n6829) );
  NAND2_X1 U8210 ( .A1(n12639), .A2(n11888), .ZN(n6830) );
  NOR2_X1 U8211 ( .A1(n12550), .A2(n10128), .ZN(n12652) );
  OAI211_X1 U8212 ( .C1(n12638), .C2(n7344), .A(n7342), .B(n6995), .ZN(n6994)
         );
  NOR2_X1 U8213 ( .A1(n11906), .A2(n6784), .ZN(n6995) );
  NAND2_X1 U8214 ( .A1(n7346), .A2(n7353), .ZN(n7344) );
  XNOR2_X1 U8215 ( .A(n7433), .B(n11905), .ZN(n7432) );
  NOR2_X1 U8216 ( .A1(n12646), .A2(n7434), .ZN(n7433) );
  NOR2_X1 U8217 ( .A1(n11887), .A2(n7435), .ZN(n7434) );
  NAND2_X1 U8218 ( .A1(n12667), .A2(n12666), .ZN(n12892) );
  OR2_X1 U8219 ( .A1(n12664), .A2(n12663), .ZN(n12667) );
  NAND2_X1 U8220 ( .A1(n9867), .A2(n15443), .ZN(n15477) );
  NAND2_X1 U8221 ( .A1(n8184), .A2(n8183), .ZN(n12205) );
  NAND2_X1 U8222 ( .A1(n12206), .A2(n8236), .ZN(n8293) );
  INV_X1 U8223 ( .A(n12671), .ZN(n12963) );
  NAND2_X1 U8224 ( .A1(n8074), .A2(n8073), .ZN(n12997) );
  OR2_X1 U8225 ( .A1(n15526), .A2(n15521), .ZN(n13014) );
  OR2_X1 U8226 ( .A1(n9388), .A2(P3_D_REG_1__SCAN_IN), .ZN(n8249) );
  XNOR2_X1 U8227 ( .A(n8022), .B(n8035), .ZN(n11899) );
  AOI21_X1 U8228 ( .B1(n13465), .B2(n13463), .A(n13462), .ZN(n13413) );
  NAND2_X1 U8229 ( .A1(n8726), .A2(n8725), .ZN(n14885) );
  NAND2_X1 U8230 ( .A1(n8931), .A2(n8930), .ZN(n13800) );
  NAND2_X1 U8231 ( .A1(n8839), .A2(n8838), .ZN(n13822) );
  INV_X1 U8232 ( .A(n13494), .ZN(n13510) );
  NAND2_X1 U8233 ( .A1(n7235), .A2(n6681), .ZN(n13580) );
  NAND2_X1 U8234 ( .A1(n9000), .A2(n8999), .ZN(n13767) );
  NAND2_X1 U8235 ( .A1(n12328), .A2(n12327), .ZN(n13858) );
  NAND2_X1 U8236 ( .A1(n11369), .A2(n11368), .ZN(n14909) );
  OR2_X1 U8237 ( .A1(n10518), .A2(n10517), .ZN(n10519) );
  NAND2_X1 U8238 ( .A1(n11667), .A2(n11666), .ZN(n14626) );
  INV_X1 U8239 ( .A(n14639), .ZN(n13961) );
  NOR2_X1 U8240 ( .A1(n15064), .A2(n15063), .ZN(n15062) );
  AND2_X1 U8241 ( .A1(n9385), .A2(n14254), .ZN(n15091) );
  NAND2_X1 U8242 ( .A1(n14419), .A2(n11785), .ZN(n14403) );
  NAND2_X1 U8243 ( .A1(n14654), .A2(n7401), .ZN(n14488) );
  NAND2_X1 U8244 ( .A1(n14654), .A2(n11722), .ZN(n14486) );
  NAND2_X1 U8245 ( .A1(n11702), .A2(n11701), .ZN(n14662) );
  NAND2_X1 U8246 ( .A1(n11384), .A2(n11383), .ZN(n14738) );
  NAND2_X1 U8247 ( .A1(n7600), .A2(n7603), .ZN(n14732) );
  INV_X1 U8248 ( .A(n6896), .ZN(n6895) );
  OAI21_X1 U8249 ( .B1(n14598), .B2(n14670), .A(n14596), .ZN(n6896) );
  XNOR2_X1 U8250 ( .A(n8352), .B(n6836), .ZN(n15563) );
  NOR2_X1 U8251 ( .A1(n14711), .A2(n14712), .ZN(n14710) );
  NAND2_X1 U8252 ( .A1(n14997), .A2(n14996), .ZN(n14995) );
  NAND2_X1 U8253 ( .A1(n6929), .A2(n7278), .ZN(n7280) );
  OR2_X1 U8254 ( .A1(n14756), .A2(n7281), .ZN(n7278) );
  NAND2_X1 U8255 ( .A1(n6930), .A2(n6714), .ZN(n6929) );
  INV_X1 U8256 ( .A(n14703), .ZN(n7279) );
  INV_X1 U8257 ( .A(n14049), .ZN(n7556) );
  OAI21_X1 U8258 ( .B1(n9121), .B2(n9161), .A(n9572), .ZN(n8462) );
  OR2_X1 U8259 ( .A1(n7553), .A2(n14073), .ZN(n7551) );
  NAND2_X1 U8260 ( .A1(n7659), .A2(n8582), .ZN(n7658) );
  INV_X1 U8261 ( .A(n8583), .ZN(n7659) );
  NAND2_X1 U8262 ( .A1(n6844), .A2(n8626), .ZN(n7669) );
  NAND2_X1 U8263 ( .A1(n6677), .A2(n7067), .ZN(n7065) );
  NOR2_X1 U8264 ( .A1(n6677), .A2(n7067), .ZN(n7066) );
  MUX2_X1 U8265 ( .A(n14266), .B(n14921), .S(n14187), .Z(n14142) );
  OAI21_X1 U8266 ( .B1(n8652), .B2(n8651), .A(n6732), .ZN(n6796) );
  INV_X1 U8267 ( .A(n8670), .ZN(n7061) );
  OAI21_X1 U8268 ( .B1(n6679), .B2(n6859), .A(n7557), .ZN(n14115) );
  NAND2_X1 U8269 ( .A1(n14110), .A2(n7558), .ZN(n7557) );
  INV_X1 U8270 ( .A(n8688), .ZN(n7652) );
  AND2_X1 U8271 ( .A1(n8670), .A2(n6743), .ZN(n7060) );
  NOR2_X1 U8272 ( .A1(n7542), .A2(n6882), .ZN(n6881) );
  INV_X1 U8273 ( .A(n14234), .ZN(n6882) );
  OR2_X1 U8274 ( .A1(n14146), .A2(n7543), .ZN(n7542) );
  OR2_X1 U8275 ( .A1(n14146), .A2(n6760), .ZN(n7539) );
  AND2_X1 U8276 ( .A1(n14524), .A2(n14149), .ZN(n7544) );
  NOR3_X1 U8277 ( .A1(n12069), .A2(n12068), .A3(n12067), .ZN(n12079) );
  OR2_X1 U8278 ( .A1(n8716), .A2(n8715), .ZN(n8741) );
  OAI21_X1 U8279 ( .B1(n14156), .B2(n14155), .A(n14154), .ZN(n14161) );
  NAND2_X1 U8280 ( .A1(n7661), .A2(n7070), .ZN(n7069) );
  NAND2_X1 U8281 ( .A1(n8805), .A2(n8804), .ZN(n7070) );
  NAND2_X1 U8282 ( .A1(n7565), .A2(n14170), .ZN(n7564) );
  AND2_X1 U8283 ( .A1(n8899), .A2(n7664), .ZN(n7663) );
  NAND2_X1 U8284 ( .A1(n7668), .A2(n7665), .ZN(n7664) );
  NAND2_X1 U8285 ( .A1(n7667), .A2(n7666), .ZN(n7665) );
  INV_X1 U8286 ( .A(n8876), .ZN(n7666) );
  INV_X1 U8287 ( .A(n8877), .ZN(n7667) );
  AND2_X1 U8288 ( .A1(n8876), .A2(n8877), .ZN(n7668) );
  NAND2_X1 U8289 ( .A1(n7563), .A2(n14178), .ZN(n7562) );
  NAND2_X1 U8290 ( .A1(n7127), .A2(n14186), .ZN(n7126) );
  INV_X1 U8291 ( .A(n14186), .ZN(n7560) );
  NAND2_X1 U8292 ( .A1(n12155), .A2(n12171), .ZN(n6867) );
  OAI21_X1 U8293 ( .B1(n8963), .B2(n7656), .A(n7653), .ZN(n8982) );
  AND2_X1 U8294 ( .A1(n8961), .A2(n8962), .ZN(n7656) );
  NAND2_X1 U8295 ( .A1(n7655), .A2(n7654), .ZN(n7653) );
  INV_X1 U8296 ( .A(n14193), .ZN(n7535) );
  AND2_X1 U8297 ( .A1(n14008), .A2(n14195), .ZN(n7549) );
  AND2_X1 U8298 ( .A1(n10928), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7005) );
  NOR2_X1 U8299 ( .A1(n11887), .A2(n12941), .ZN(n7354) );
  INV_X1 U8300 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7692) );
  NOR2_X1 U8301 ( .A1(P3_IR_REG_11__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n7689) );
  INV_X1 U8302 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8416) );
  OR2_X1 U8303 ( .A1(n8698), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n8609) );
  OAI21_X1 U8304 ( .B1(n11735), .B2(n6774), .A(n7033), .ZN(n8985) );
  INV_X1 U8305 ( .A(n8881), .ZN(n7113) );
  NAND2_X1 U8306 ( .A1(n6775), .A2(n6661), .ZN(n7590) );
  NAND2_X1 U8307 ( .A1(n8859), .A2(n9774), .ZN(n8881) );
  INV_X1 U8308 ( .A(n7125), .ZN(n7123) );
  INV_X1 U8309 ( .A(n7028), .ZN(n7027) );
  OAI21_X1 U8310 ( .B1(n7576), .B2(n7578), .A(n8806), .ZN(n7028) );
  INV_X1 U8311 ( .A(n8744), .ZN(n6968) );
  INV_X1 U8312 ( .A(n8689), .ZN(n8692) );
  INV_X1 U8313 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7572) );
  INV_X1 U8314 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7025) );
  INV_X1 U8315 ( .A(n12000), .ZN(n7307) );
  OR3_X1 U8316 ( .A1(n12725), .A2(n12152), .A3(n12035), .ZN(n12036) );
  OR4_X1 U8317 ( .A1(n8104), .A2(n12761), .A3(n12789), .A4(n12034), .ZN(n12035) );
  NOR2_X1 U8318 ( .A1(n12178), .A2(n6806), .ZN(n6805) );
  NAND2_X1 U8319 ( .A1(n6685), .A2(n6807), .ZN(n6806) );
  INV_X1 U8320 ( .A(n12038), .ZN(n6807) );
  NOR2_X1 U8321 ( .A1(n10306), .A2(n10149), .ZN(n10151) );
  AOI21_X1 U8322 ( .B1(P3_REG1_REG_4__SCAN_IN), .B2(n10167), .A(n10399), .ZN(
        n10169) );
  AND2_X1 U8323 ( .A1(n7000), .A2(n6999), .ZN(n11255) );
  NAND2_X1 U8324 ( .A1(n7358), .A2(n6998), .ZN(n7000) );
  AOI21_X1 U8325 ( .B1(n7001), .B2(n7002), .A(n7005), .ZN(n6999) );
  NOR2_X1 U8326 ( .A1(n10499), .A2(n15540), .ZN(n6998) );
  OR2_X1 U8327 ( .A1(n12671), .A2(n12683), .ZN(n8229) );
  OR2_X1 U8328 ( .A1(n12898), .A2(n12684), .ZN(n12162) );
  NAND2_X1 U8329 ( .A1(n12789), .A2(n12134), .ZN(n7103) );
  OR2_X1 U8330 ( .A1(n12150), .A2(n12759), .ZN(n8224) );
  AND2_X1 U8331 ( .A1(n12148), .A2(n12016), .ZN(n12146) );
  NAND2_X1 U8332 ( .A1(n7998), .A2(n7469), .ZN(n7468) );
  NAND2_X1 U8333 ( .A1(n12856), .A2(n12833), .ZN(n12042) );
  NOR2_X1 U8334 ( .A1(n7453), .A2(n7451), .ZN(n7450) );
  NAND2_X1 U8335 ( .A1(n7078), .A2(n12074), .ZN(n7077) );
  INV_X1 U8336 ( .A(n12074), .ZN(n7079) );
  OR2_X1 U8337 ( .A1(n9388), .A2(n8260), .ZN(n8280) );
  NAND2_X1 U8338 ( .A1(n8222), .A2(n12137), .ZN(n12790) );
  NOR2_X1 U8339 ( .A1(n7087), .A2(n7091), .ZN(n7086) );
  INV_X1 U8340 ( .A(n12130), .ZN(n7091) );
  INV_X1 U8341 ( .A(n7768), .ZN(n7305) );
  INV_X1 U8342 ( .A(n7743), .ZN(n7297) );
  NOR2_X1 U8343 ( .A1(n7297), .A2(n7294), .ZN(n7293) );
  INV_X1 U8344 ( .A(n7741), .ZN(n7294) );
  NAND2_X1 U8345 ( .A1(n7959), .A2(n7738), .ZN(n7285) );
  NAND2_X1 U8346 ( .A1(n7285), .A2(n8719), .ZN(n7739) );
  NOR2_X1 U8347 ( .A1(n7950), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n7954) );
  INV_X1 U8348 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n7733) );
  INV_X1 U8349 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7724) );
  AND2_X1 U8350 ( .A1(n7429), .A2(n7818), .ZN(n7478) );
  INV_X1 U8351 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n13315) );
  NAND2_X1 U8352 ( .A1(n7502), .A2(n6708), .ZN(n7501) );
  NAND2_X1 U8353 ( .A1(n10585), .A2(n6653), .ZN(n7502) );
  NOR2_X1 U8354 ( .A1(n7501), .A2(n7499), .ZN(n7498) );
  INV_X1 U8355 ( .A(n9923), .ZN(n7499) );
  OR2_X1 U8356 ( .A1(n7073), .A2(n9136), .ZN(n7072) );
  NAND2_X1 U8357 ( .A1(n6683), .A2(n9142), .ZN(n7073) );
  NOR2_X1 U8358 ( .A1(n9126), .A2(n9049), .ZN(n9087) );
  NOR2_X1 U8359 ( .A1(n9088), .A2(n9089), .ZN(n7040) );
  INV_X1 U8360 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8409) );
  NOR2_X1 U8361 ( .A1(n13767), .A2(n13596), .ZN(n7321) );
  NOR2_X1 U8362 ( .A1(n13628), .A2(n13779), .ZN(n7323) );
  NOR2_X1 U8363 ( .A1(n13800), .A2(n13681), .ZN(n7317) );
  AND2_X1 U8364 ( .A1(n8865), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8884) );
  NOR2_X1 U8365 ( .A1(n8840), .A2(n11185), .ZN(n8865) );
  NOR2_X1 U8366 ( .A1(n11818), .A2(n7250), .ZN(n7249) );
  INV_X1 U8367 ( .A(n11816), .ZN(n7250) );
  OR2_X1 U8368 ( .A1(n13750), .A2(n7328), .ZN(n7327) );
  NOR2_X1 U8369 ( .A1(n7256), .A2(n7254), .ZN(n7253) );
  INV_X1 U8370 ( .A(n10990), .ZN(n7254) );
  INV_X1 U8371 ( .A(n7257), .ZN(n7256) );
  INV_X1 U8372 ( .A(n10758), .ZN(n7221) );
  NOR2_X1 U8373 ( .A1(n10225), .A2(n10239), .ZN(n7315) );
  AND2_X1 U8374 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8543) );
  NAND2_X1 U8375 ( .A1(n7330), .A2(n7329), .ZN(n9641) );
  AND2_X1 U8376 ( .A1(n15307), .A2(n8474), .ZN(n7329) );
  INV_X1 U8377 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n7224) );
  INV_X1 U8378 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8451) );
  INV_X1 U8379 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8410) );
  OR2_X1 U8380 ( .A1(n8656), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n8674) );
  OR2_X1 U8381 ( .A1(n8636), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n8656) );
  INV_X1 U8382 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n7648) );
  INV_X1 U8383 ( .A(n7143), .ZN(n7137) );
  INV_X1 U8384 ( .A(n11062), .ZN(n7136) );
  OAI21_X1 U8385 ( .B1(n14204), .B2(n14203), .A(n14202), .ZN(n14209) );
  NAND2_X1 U8386 ( .A1(n14416), .A2(n11785), .ZN(n7617) );
  INV_X1 U8387 ( .A(n14263), .ZN(n13985) );
  INV_X1 U8388 ( .A(n14264), .ZN(n13986) );
  AND2_X1 U8389 ( .A1(n7392), .A2(n7394), .ZN(n7391) );
  INV_X1 U8390 ( .A(n11668), .ZN(n7404) );
  OAI21_X1 U8391 ( .B1(n6676), .B2(n7404), .A(n14238), .ZN(n7403) );
  AND2_X1 U8392 ( .A1(n7593), .A2(n14232), .ZN(n6654) );
  INV_X1 U8393 ( .A(n15108), .ZN(n14043) );
  AND2_X1 U8394 ( .A1(n11432), .A2(n14968), .ZN(n11552) );
  NOR2_X2 U8395 ( .A1(n14740), .A2(n14112), .ZN(n11432) );
  NAND2_X1 U8396 ( .A1(n7583), .A2(n7584), .ZN(n9091) );
  AOI21_X1 U8397 ( .B1(n7586), .B2(n8993), .A(n7585), .ZN(n7584) );
  INV_X1 U8398 ( .A(n9070), .ZN(n7585) );
  INV_X1 U8399 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9235) );
  NAND2_X1 U8400 ( .A1(n7114), .A2(n8881), .ZN(n8925) );
  NAND2_X1 U8401 ( .A1(n8880), .A2(n8879), .ZN(n7114) );
  INV_X1 U8402 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n7570) );
  NAND2_X1 U8403 ( .A1(n8833), .A2(SI_17_), .ZN(n7125) );
  INV_X1 U8404 ( .A(n8834), .ZN(n6965) );
  AND2_X1 U8405 ( .A1(n7612), .A2(n6668), .ZN(n6934) );
  AND3_X2 U8406 ( .A1(n13315), .A2(n7537), .A3(n7536), .ZN(n9485) );
  AND4_X2 U8407 ( .A1(n9284), .A2(n9353), .A3(n9679), .A4(n9484), .ZN(n9208)
         );
  NAND2_X1 U8408 ( .A1(n8345), .A2(n9300), .ZN(n7283) );
  OAI21_X1 U8409 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(n13266), .A(n8307), .ZN(
        n8308) );
  OAI21_X1 U8410 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n8314), .A(n8313), .ZN(
        n8315) );
  OAI21_X1 U8411 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n8319), .A(n8318), .ZN(
        n8338) );
  OAI21_X1 U8412 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(n8322), .A(n8321), .ZN(
        n8383) );
  OAI21_X1 U8413 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n12590), .A(n8325), .ZN(
        n8326) );
  NOR2_X1 U8414 ( .A1(n7186), .A2(n7182), .ZN(n7181) );
  INV_X1 U8415 ( .A(n11521), .ZN(n7182) );
  INV_X1 U8416 ( .A(n11524), .ZN(n7186) );
  NAND2_X1 U8417 ( .A1(n11524), .A2(n7185), .ZN(n7184) );
  INV_X1 U8418 ( .A(n11523), .ZN(n7185) );
  INV_X1 U8419 ( .A(n12417), .ZN(n7164) );
  AOI21_X1 U8420 ( .B1(n12415), .B2(n7169), .A(n6702), .ZN(n7168) );
  NAND2_X1 U8421 ( .A1(n12415), .A2(n7171), .ZN(n7170) );
  INV_X1 U8422 ( .A(n12512), .ZN(n7171) );
  AND2_X1 U8423 ( .A1(n10003), .A2(n9999), .ZN(n10028) );
  NAND2_X1 U8424 ( .A1(n8132), .A2(n12480), .ZN(n8143) );
  INV_X1 U8425 ( .A(n14764), .ZN(n11609) );
  OR2_X1 U8426 ( .A1(n7914), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7930) );
  NAND2_X1 U8427 ( .A1(n10471), .A2(n10472), .ZN(n10834) );
  AND4_X1 U8428 ( .A1(n12006), .A2(n8189), .A3(n8188), .A4(n8187), .ZN(n12536)
         );
  AND4_X1 U8429 ( .A1(n7874), .A2(n7873), .A3(n7872), .A4(n7871), .ZN(n12431)
         );
  NOR2_X1 U8430 ( .A1(n10258), .A2(n15529), .ZN(n10257) );
  NOR2_X1 U8431 ( .A1(n10255), .A2(n15476), .ZN(n10254) );
  INV_X1 U8432 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7429) );
  NAND2_X1 U8433 ( .A1(n7007), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7340) );
  INV_X1 U8434 ( .A(n10436), .ZN(n7007) );
  NOR2_X1 U8435 ( .A1(n10432), .A2(n10152), .ZN(n10398) );
  NOR2_X1 U8436 ( .A1(n10151), .A2(n10150), .ZN(n10152) );
  NOR2_X1 U8437 ( .A1(n10420), .A2(n15536), .ZN(n10419) );
  OAI21_X1 U8438 ( .B1(n10420), .B2(n7356), .A(n7355), .ZN(n10460) );
  NAND2_X1 U8439 ( .A1(n7357), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7356) );
  NAND2_X1 U8440 ( .A1(n10170), .A2(n7357), .ZN(n7355) );
  INV_X1 U8441 ( .A(n10172), .ZN(n7357) );
  INV_X1 U8442 ( .A(n10496), .ZN(n7440) );
  XNOR2_X1 U8443 ( .A(n11255), .B(n7439), .ZN(n10930) );
  OAI21_X1 U8444 ( .B1(n10919), .B2(n10928), .A(n10918), .ZN(n11275) );
  NOR2_X1 U8445 ( .A1(n10916), .A2(n6767), .ZN(n11263) );
  XNOR2_X1 U8446 ( .A(n7010), .B(n11268), .ZN(n11321) );
  INV_X1 U8447 ( .A(n11316), .ZN(n6827) );
  NAND2_X1 U8448 ( .A1(n7012), .A2(n7011), .ZN(n7010) );
  NAND2_X1 U8449 ( .A1(n15417), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7011) );
  INV_X1 U8450 ( .A(n7436), .ZN(n11267) );
  NOR2_X1 U8451 ( .A1(n11854), .A2(n7359), .ZN(n11855) );
  NOR2_X1 U8452 ( .A1(n11282), .A2(n14802), .ZN(n7359) );
  INV_X1 U8453 ( .A(n6977), .ZN(n6976) );
  OAI21_X1 U8454 ( .B1(n6675), .B2(n12570), .A(n11895), .ZN(n6977) );
  NAND2_X1 U8455 ( .A1(n7332), .A2(n11874), .ZN(n11858) );
  NAND2_X1 U8456 ( .A1(n7442), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7441) );
  NAND2_X1 U8457 ( .A1(n11897), .A2(n7442), .ZN(n6978) );
  INV_X1 U8458 ( .A(n12613), .ZN(n7442) );
  NAND2_X1 U8459 ( .A1(n7338), .A2(n7337), .ZN(n7336) );
  NAND2_X1 U8460 ( .A1(n11899), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n7337) );
  NOR2_X1 U8461 ( .A1(n6782), .A2(n15425), .ZN(n7343) );
  INV_X1 U8462 ( .A(n7350), .ZN(n7345) );
  NAND2_X1 U8463 ( .A1(n7351), .A2(n7347), .ZN(n7346) );
  OR2_X1 U8464 ( .A1(n12637), .A2(n7352), .ZN(n7351) );
  INV_X1 U8465 ( .A(n12409), .ZN(n7431) );
  OAI21_X1 U8466 ( .B1(n12622), .B2(n6981), .A(n6980), .ZN(n12646) );
  NAND2_X1 U8467 ( .A1(n6982), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n6981) );
  NAND2_X1 U8468 ( .A1(n11903), .A2(n6982), .ZN(n6980) );
  INV_X1 U8469 ( .A(n12647), .ZN(n6982) );
  AND2_X1 U8470 ( .A1(n8229), .A2(n8228), .ZN(n12669) );
  NOR2_X1 U8471 ( .A1(n12661), .A2(n12669), .ZN(n12664) );
  INV_X1 U8472 ( .A(n7457), .ZN(n7456) );
  AOI21_X1 U8473 ( .B1(n7457), .B2(n7455), .A(n6704), .ZN(n7454) );
  NAND2_X1 U8474 ( .A1(n6846), .A2(n8127), .ZN(n12724) );
  NAND2_X1 U8475 ( .A1(n12739), .A2(n12153), .ZN(n12723) );
  AND4_X1 U8476 ( .A1(n8103), .A2(n8102), .A3(n8101), .A4(n8100), .ZN(n12755)
         );
  INV_X1 U8477 ( .A(n12768), .ZN(n8104) );
  NAND2_X1 U8478 ( .A1(n12928), .A2(n12134), .ZN(n12776) );
  NAND2_X1 U8479 ( .A1(n12782), .A2(n8090), .ZN(n12769) );
  OR2_X1 U8480 ( .A1(n8098), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8109) );
  NAND2_X1 U8481 ( .A1(n12797), .A2(n8080), .ZN(n12783) );
  AND4_X1 U8482 ( .A1(n8089), .A2(n8088), .A3(n8087), .A4(n8086), .ZN(n12799)
         );
  NOR2_X1 U8483 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(n7674), .ZN(n8084) );
  OAI211_X1 U8484 ( .C1(n7998), .C2(n7465), .A(n7463), .B(n8063), .ZN(n12811)
         );
  INV_X1 U8485 ( .A(n7466), .ZN(n7465) );
  AND2_X1 U8486 ( .A1(n12125), .A2(n12136), .ZN(n12814) );
  INV_X1 U8487 ( .A(n12814), .ZN(n12821) );
  NAND2_X1 U8488 ( .A1(n7468), .A2(n7466), .ZN(n12829) );
  NAND2_X1 U8489 ( .A1(n7468), .A2(n8017), .ZN(n12845) );
  NOR2_X1 U8490 ( .A1(n8010), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8027) );
  AND2_X1 U8491 ( .A1(n8027), .A2(n8026), .ZN(n8041) );
  NOR2_X1 U8492 ( .A1(n8215), .A2(n7093), .ZN(n7092) );
  INV_X1 U8493 ( .A(n12111), .ZN(n7093) );
  INV_X1 U8494 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n11607) );
  NOR2_X1 U8495 ( .A1(n7944), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7976) );
  INV_X1 U8496 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n13326) );
  AND2_X1 U8497 ( .A1(n7887), .A2(n7886), .ZN(n7900) );
  OR2_X1 U8498 ( .A1(n7854), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7869) );
  NAND2_X1 U8499 ( .A1(n8209), .A2(n8208), .ZN(n10974) );
  NAND2_X1 U8500 ( .A1(n10379), .A2(n7474), .ZN(n10977) );
  AND2_X1 U8501 ( .A1(n12067), .A2(n7838), .ZN(n7474) );
  NAND2_X1 U8502 ( .A1(n10379), .A2(n7838), .ZN(n10975) );
  INV_X1 U8503 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n10418) );
  NAND2_X1 U8504 ( .A1(n15440), .A2(n12056), .ZN(n10480) );
  INV_X1 U8505 ( .A(n12019), .ZN(n7824) );
  NAND2_X1 U8506 ( .A1(n9863), .A2(n9862), .ZN(n9867) );
  AND4_X1 U8507 ( .A1(n12006), .A2(n12005), .A3(n12004), .A4(n12003), .ZN(
        n12656) );
  NAND2_X1 U8508 ( .A1(n7105), .A2(n7104), .ZN(n12928) );
  INV_X1 U8509 ( .A(n12789), .ZN(n7104) );
  INV_X1 U8510 ( .A(n12790), .ZN(n7105) );
  NOR2_X1 U8511 ( .A1(n8288), .A2(n8287), .ZN(n10013) );
  NOR2_X1 U8512 ( .A1(n8281), .A2(n8287), .ZN(n10015) );
  AND4_X2 U8513 ( .A1(n7785), .A2(n7784), .A3(n7783), .A4(n7782), .ZN(n15451)
         );
  NOR2_X1 U8514 ( .A1(n6706), .A2(n7476), .ZN(n7475) );
  NAND2_X1 U8515 ( .A1(n7694), .A2(n7201), .ZN(n7476) );
  INV_X1 U8516 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7776) );
  NAND2_X1 U8517 ( .A1(n7766), .A2(n7765), .ZN(n8151) );
  OAI21_X1 U8518 ( .B1(n7763), .B2(n7311), .A(n7310), .ZN(n8140) );
  NAND2_X1 U8519 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n11813), .ZN(n7310) );
  AND2_X1 U8520 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n11351), .ZN(n7311) );
  NOR2_X1 U8521 ( .A1(n8106), .A2(n7300), .ZN(n7299) );
  XNOR2_X1 U8522 ( .A(n8267), .B(n13256), .ZN(n10125) );
  INV_X1 U8523 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8191) );
  INV_X1 U8524 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8193) );
  NAND2_X1 U8525 ( .A1(n6916), .A2(n6658), .ZN(n8237) );
  AND2_X1 U8526 ( .A1(n7751), .A2(n7750), .ZN(n8048) );
  NAND2_X1 U8527 ( .A1(n8021), .A2(n7745), .ZN(n8034) );
  AND2_X1 U8528 ( .A1(n7741), .A2(n7740), .ZN(n7982) );
  OR2_X1 U8529 ( .A1(n7957), .A2(n7956), .ZN(n7959) );
  OR2_X1 U8530 ( .A1(n7937), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n7950) );
  NAND2_X1 U8531 ( .A1(n6802), .A2(n7728), .ZN(n7907) );
  INV_X1 U8532 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n7727) );
  XNOR2_X1 U8533 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n7895) );
  INV_X1 U8534 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n7198) );
  INV_X1 U8535 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n7687) );
  XNOR2_X1 U8536 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n7834) );
  XNOR2_X1 U8537 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n7805) );
  NAND2_X1 U8538 ( .A1(n8448), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7794) );
  INV_X1 U8539 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8448) );
  AND2_X1 U8540 ( .A1(n7504), .A2(n10099), .ZN(n7503) );
  INV_X1 U8541 ( .A(n10367), .ZN(n7504) );
  XNOR2_X1 U8542 ( .A(n11968), .B(n9568), .ZN(n9613) );
  AOI21_X1 U8543 ( .B1(n7521), .B2(n11160), .A(n7519), .ZN(n7518) );
  INV_X1 U8544 ( .A(n11241), .ZN(n7519) );
  AND2_X1 U8545 ( .A1(n7526), .A2(n7525), .ZN(n13430) );
  NAND2_X1 U8546 ( .A1(n11917), .A2(n11918), .ZN(n7525) );
  OR2_X1 U8547 ( .A1(n11913), .A2(n7527), .ZN(n7526) );
  NAND2_X1 U8548 ( .A1(n13430), .A2(n13431), .ZN(n13429) );
  NAND2_X1 U8549 ( .A1(n9921), .A2(n9920), .ZN(n9922) );
  NAND2_X1 U8550 ( .A1(n9791), .A2(n9790), .ZN(n9921) );
  OR2_X1 U8551 ( .A1(n8641), .A2(n8640), .ZN(n8661) );
  NOR2_X1 U8552 ( .A1(n8932), .A2(n13477), .ZN(n8953) );
  OR2_X1 U8553 ( .A1(n7489), .A2(n11939), .ZN(n7488) );
  OAI21_X1 U8554 ( .B1(n13483), .B2(n7484), .A(n7481), .ZN(n7490) );
  AND2_X1 U8555 ( .A1(n13412), .A2(n7492), .ZN(n7489) );
  NOR2_X1 U8556 ( .A1(n11164), .A2(n7522), .ZN(n7521) );
  INV_X1 U8557 ( .A(n7524), .ZN(n7522) );
  NAND2_X1 U8558 ( .A1(n11158), .A2(n11159), .ZN(n7524) );
  OR2_X1 U8559 ( .A1(n11161), .A2(n11160), .ZN(n7523) );
  NAND2_X1 U8560 ( .A1(n9478), .A2(n9469), .ZN(n13492) );
  AND2_X1 U8561 ( .A1(n9197), .A2(n6637), .ZN(n9478) );
  AND4_X1 U8562 ( .A1(n9100), .A2(n9099), .A3(n9098), .A4(n9097), .ZN(n11972)
         );
  AND4_X1 U8563 ( .A1(n9025), .A2(n9024), .A3(n9023), .A4(n9022), .ZN(n13493)
         );
  AND4_X1 U8564 ( .A1(n9061), .A2(n9060), .A3(n9059), .A4(n9058), .ZN(n13494)
         );
  INV_X1 U8565 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8408) );
  NAND2_X1 U8566 ( .A1(n7321), .A2(n7320), .ZN(n13570) );
  NOR2_X1 U8567 ( .A1(n13570), .A2(n13569), .ZN(n13571) );
  AND2_X1 U8568 ( .A1(n11844), .A2(n6681), .ZN(n7234) );
  AND2_X1 U8569 ( .A1(n9095), .A2(n9004), .ZN(n13586) );
  NAND2_X1 U8570 ( .A1(n7323), .A2(n7322), .ZN(n13596) );
  INV_X1 U8571 ( .A(n7323), .ZN(n13612) );
  AND2_X1 U8572 ( .A1(n9021), .A2(n9020), .ZN(n13598) );
  NOR2_X1 U8573 ( .A1(n13779), .A2(n13509), .ZN(n6898) );
  AND2_X1 U8574 ( .A1(n9039), .A2(n9038), .ZN(n13614) );
  INV_X1 U8575 ( .A(n7261), .ZN(n7260) );
  OAI22_X1 U8576 ( .A1(n13645), .A2(n7267), .B1(n13511), .B2(n13644), .ZN(
        n7261) );
  NAND2_X1 U8577 ( .A1(n7418), .A2(n11841), .ZN(n7416) );
  NAND2_X1 U8578 ( .A1(n7317), .A2(n7316), .ZN(n13656) );
  INV_X1 U8579 ( .A(n7317), .ZN(n13667) );
  NAND2_X1 U8580 ( .A1(n7319), .A2(n7318), .ZN(n13681) );
  INV_X1 U8581 ( .A(n13804), .ZN(n7318) );
  INV_X1 U8582 ( .A(n7319), .ZN(n13703) );
  INV_X1 U8583 ( .A(n13737), .ZN(n6893) );
  OR2_X1 U8584 ( .A1(n8817), .A2(n8816), .ZN(n8840) );
  NAND2_X1 U8585 ( .A1(n6848), .A2(n6847), .ZN(n14823) );
  NOR2_X1 U8586 ( .A1(n14850), .A2(n7328), .ZN(n14817) );
  OR2_X1 U8587 ( .A1(n8754), .A2(n13189), .ZN(n8775) );
  AOI21_X1 U8588 ( .B1(n7413), .B2(n7415), .A(n6711), .ZN(n7412) );
  AND2_X1 U8589 ( .A1(n10767), .A2(n15381), .ZN(n11013) );
  NAND2_X1 U8590 ( .A1(n10680), .A2(n15355), .ZN(n10679) );
  NOR2_X1 U8591 ( .A1(n10298), .A2(n15347), .ZN(n10680) );
  AOI21_X1 U8592 ( .B1(n10289), .B2(n7241), .A(n6710), .ZN(n7240) );
  NAND2_X1 U8593 ( .A1(n7315), .A2(n7314), .ZN(n10298) );
  INV_X1 U8594 ( .A(n7315), .ZN(n10246) );
  INV_X1 U8595 ( .A(n14841), .ZN(n14819) );
  INV_X1 U8596 ( .A(n10348), .ZN(n10346) );
  OR2_X1 U8597 ( .A1(n9336), .A2(n9109), .ZN(n8492) );
  NAND2_X1 U8598 ( .A1(n6643), .A2(n6858), .ZN(n6857) );
  CLKBUF_X1 U8599 ( .A(n9644), .Z(n6890) );
  NAND2_X1 U8600 ( .A1(n13662), .A2(n7268), .ZN(n13650) );
  NAND2_X1 U8601 ( .A1(n8639), .A2(n8638), .ZN(n15361) );
  CLKBUF_X1 U8602 ( .A(n9611), .Z(n15342) );
  INV_X1 U8603 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7639) );
  XNOR2_X1 U8604 ( .A(n9185), .B(P2_IR_REG_26__SCAN_IN), .ZN(n9462) );
  AND2_X1 U8605 ( .A1(n7533), .A2(n8434), .ZN(n8450) );
  CLKBUF_X1 U8606 ( .A(n9187), .Z(n9188) );
  INV_X1 U8607 ( .A(n8434), .ZN(n8697) );
  INV_X1 U8608 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8486) );
  INV_X1 U8609 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6941) );
  INV_X1 U8610 ( .A(n14262), .ZN(n12339) );
  AND2_X1 U8611 ( .A1(n11738), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n11749) );
  OR2_X1 U8612 ( .A1(n11356), .A2(n11357), .ZN(n7128) );
  AOI21_X1 U8613 ( .B1(n12333), .B2(n9935), .A(n9269), .ZN(n9274) );
  NAND2_X1 U8614 ( .A1(n14905), .A2(n6772), .ZN(n12248) );
  OR2_X1 U8615 ( .A1(n11397), .A2(n11370), .ZN(n11404) );
  NOR2_X1 U8616 ( .A1(n6886), .A2(n6885), .ZN(n6884) );
  INV_X1 U8617 ( .A(n14216), .ZN(n6886) );
  NOR2_X1 U8618 ( .A1(n14361), .A2(n14218), .ZN(n6885) );
  NAND2_X1 U8619 ( .A1(n9829), .A2(n9830), .ZN(n14281) );
  AND3_X1 U8620 ( .A1(n9828), .A2(n9827), .A3(n9826), .ZN(n9830) );
  OR2_X1 U8621 ( .A1(n9754), .A2(n9753), .ZN(n7023) );
  NOR2_X1 U8622 ( .A1(n15006), .A2(n6766), .ZN(n10042) );
  NAND2_X1 U8623 ( .A1(n10042), .A2(n10043), .ZN(n14326) );
  AOI21_X1 U8624 ( .B1(n15023), .B2(P1_REG1_REG_13__SCAN_IN), .A(n15018), .ZN(
        n15032) );
  NOR2_X1 U8625 ( .A1(n15015), .A2(n7020), .ZN(n15028) );
  AND2_X1 U8626 ( .A1(n15023), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7020) );
  INV_X1 U8627 ( .A(n14327), .ZN(n14328) );
  XNOR2_X1 U8628 ( .A(n15052), .B(n14340), .ZN(n15048) );
  NOR2_X1 U8629 ( .A1(n15027), .A2(n7019), .ZN(n14327) );
  AND2_X1 U8630 ( .A1(n14338), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7019) );
  NOR2_X1 U8631 ( .A1(n15072), .A2(n7014), .ZN(n14331) );
  AND2_X1 U8632 ( .A1(n14343), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7014) );
  INV_X1 U8633 ( .A(n7211), .ZN(n7209) );
  NAND2_X1 U8634 ( .A1(n7205), .A2(n14448), .ZN(n14443) );
  NAND2_X1 U8635 ( .A1(n7204), .A2(n14620), .ZN(n14421) );
  INV_X1 U8636 ( .A(n14443), .ZN(n7204) );
  OR2_X1 U8637 ( .A1(n11703), .A2(n13880), .ZN(n11714) );
  NOR2_X1 U8638 ( .A1(n14576), .A2(n7206), .ZN(n14548) );
  INV_X1 U8639 ( .A(n7208), .ZN(n7206) );
  OR2_X1 U8640 ( .A1(n14527), .A2(n14528), .ZN(n7628) );
  NAND2_X1 U8641 ( .A1(n14544), .A2(n7545), .ZN(n14543) );
  OAI21_X1 U8642 ( .B1(n11541), .B2(n7632), .A(n7631), .ZN(n7678) );
  NAND2_X1 U8643 ( .A1(n7634), .A2(n7676), .ZN(n7631) );
  NAND2_X1 U8644 ( .A1(n7676), .A2(n7633), .ZN(n7632) );
  NAND2_X1 U8645 ( .A1(n7678), .A2(n11781), .ZN(n14558) );
  NOR2_X1 U8646 ( .A1(n11404), .A2(n11403), .ZN(n11542) );
  AND2_X1 U8647 ( .A1(n11542), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n11678) );
  NAND2_X1 U8648 ( .A1(n11376), .A2(n7607), .ZN(n7600) );
  OR3_X1 U8649 ( .A1(n11091), .A2(n11090), .A3(n11089), .ZN(n11386) );
  NOR2_X1 U8650 ( .A1(n11122), .A2(n14097), .ZN(n11482) );
  INV_X1 U8651 ( .A(n7621), .ZN(n7620) );
  OAI21_X1 U8652 ( .B1(n7624), .B2(n14226), .A(n6688), .ZN(n7621) );
  NAND2_X1 U8653 ( .A1(n7202), .A2(n14079), .ZN(n11122) );
  OR2_X1 U8654 ( .A1(n11086), .A2(n7624), .ZN(n11124) );
  NOR2_X1 U8655 ( .A1(n11086), .A2(n11085), .ZN(n11125) );
  NAND2_X1 U8656 ( .A1(n11118), .A2(n14231), .ZN(n11120) );
  NAND2_X1 U8657 ( .A1(n11103), .A2(n11102), .ZN(n11118) );
  NAND2_X1 U8658 ( .A1(n10857), .A2(n10871), .ZN(n11103) );
  NOR2_X1 U8659 ( .A1(n10872), .A2(n10871), .ZN(n11086) );
  INV_X1 U8660 ( .A(n14225), .ZN(n10565) );
  NOR2_X1 U8661 ( .A1(n6697), .A2(n7381), .ZN(n7380) );
  INV_X1 U8662 ( .A(n9951), .ZN(n7381) );
  INV_X1 U8663 ( .A(n10562), .ZN(n14224) );
  NAND2_X1 U8664 ( .A1(n7203), .A2(n10536), .ZN(n10340) );
  INV_X1 U8665 ( .A(n10649), .ZN(n7203) );
  INV_X1 U8666 ( .A(n14047), .ZN(n14221) );
  NAND2_X1 U8667 ( .A1(n15122), .A2(n15179), .ZN(n10649) );
  NAND2_X1 U8668 ( .A1(n10561), .A2(n10560), .ZN(n11803) );
  NAND2_X1 U8669 ( .A1(n7628), .A2(n6656), .ZN(n14649) );
  INV_X1 U8670 ( .A(n14921), .ZN(n14951) );
  OR2_X1 U8671 ( .A1(n14960), .A2(n7634), .ZN(n14569) );
  NAND2_X1 U8672 ( .A1(n7595), .A2(n7593), .ZN(n11427) );
  NAND2_X1 U8673 ( .A1(n7596), .A2(n7598), .ZN(n7595) );
  INV_X1 U8674 ( .A(n14074), .ZN(n14087) );
  INV_X1 U8675 ( .A(n15187), .ZN(n14955) );
  XNOR2_X1 U8676 ( .A(n9218), .B(n9217), .ZN(n9587) );
  INV_X1 U8677 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9217) );
  OAI21_X1 U8678 ( .B1(n8769), .B2(n7579), .A(n7031), .ZN(n8807) );
  AOI21_X1 U8679 ( .B1(n8768), .B2(n7578), .A(n7576), .ZN(n7031) );
  OAI21_X1 U8680 ( .B1(n8768), .B2(n9377), .A(n8767), .ZN(n7580) );
  OR2_X1 U8681 ( .A1(n9608), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n9609) );
  OAI21_X1 U8682 ( .B1(n8694), .B2(n6972), .A(n6969), .ZN(n8745) );
  NAND2_X1 U8683 ( .A1(n8694), .A2(n6975), .ZN(n6973) );
  OAI21_X1 U8684 ( .B1(n8672), .B2(n9340), .A(n8671), .ZN(n8673) );
  OAI21_X1 U8685 ( .B1(n8606), .B2(n6939), .A(n6910), .ZN(n6909) );
  INV_X1 U8686 ( .A(n8607), .ZN(n6939) );
  AND2_X1 U8687 ( .A1(n6937), .A2(n8628), .ZN(n6910) );
  OAI21_X1 U8688 ( .B1(n9368), .B2(P1_IR_REG_8__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9550) );
  OR2_X1 U8689 ( .A1(n9363), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9368) );
  NAND2_X1 U8690 ( .A1(n6938), .A2(n8607), .ZN(n8629) );
  NAND2_X1 U8691 ( .A1(n8606), .A2(n8605), .ZN(n6938) );
  OR2_X1 U8692 ( .A1(n9356), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n9363) );
  INV_X1 U8693 ( .A(n7116), .ZN(n8585) );
  AOI21_X1 U8694 ( .B1(n8565), .B2(n8564), .A(n7118), .ZN(n7116) );
  INV_X1 U8695 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9351) );
  OAI21_X1 U8696 ( .B1(n8507), .B2(n8521), .A(n8508), .ZN(n8509) );
  NAND2_X1 U8697 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n6834), .ZN(n6833) );
  AND2_X1 U8698 ( .A1(n7270), .A2(n14981), .ZN(n8376) );
  OAI21_X1 U8699 ( .B1(n14983), .B2(n14982), .A(n7271), .ZN(n7270) );
  INV_X1 U8700 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7271) );
  INV_X1 U8701 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n7281) );
  AND3_X1 U8702 ( .A1(n7884), .A2(n7883), .A3(n7882), .ZN(n10778) );
  OR2_X1 U8703 ( .A1(n8169), .A2(n8168), .ZN(n12688) );
  INV_X1 U8704 ( .A(n7169), .ZN(n7167) );
  INV_X1 U8705 ( .A(n12415), .ZN(n6927) );
  AND4_X1 U8706 ( .A1(n7936), .A2(n7935), .A3(n7934), .A4(n7933), .ZN(n14777)
         );
  NAND2_X1 U8707 ( .A1(n10910), .A2(n10909), .ZN(n11226) );
  AND2_X1 U8708 ( .A1(n7177), .A2(n12371), .ZN(n7176) );
  NAND2_X1 U8709 ( .A1(n12487), .A2(n12376), .ZN(n12440) );
  AND3_X1 U8710 ( .A1(n7851), .A2(n7850), .A3(n7849), .ZN(n10476) );
  NAND2_X1 U8711 ( .A1(n12468), .A2(n12467), .ZN(n12466) );
  NAND2_X1 U8712 ( .A1(n7191), .A2(n6674), .ZN(n10843) );
  NAND2_X1 U8713 ( .A1(n8083), .A2(n8082), .ZN(n12788) );
  NAND2_X1 U8714 ( .A1(n7187), .A2(n11523), .ZN(n11614) );
  NAND2_X1 U8715 ( .A1(n11522), .A2(n11521), .ZN(n7187) );
  AND4_X2 U8716 ( .A1(n7814), .A2(n7813), .A3(n7812), .A4(n7811), .ZN(n15449)
         );
  NAND2_X1 U8717 ( .A1(n8170), .A2(n10488), .ZN(n7812) );
  AND4_X1 U8718 ( .A1(n8046), .A2(n8045), .A3(n8044), .A4(n8043), .ZN(n12816)
         );
  NAND2_X1 U8719 ( .A1(n12506), .A2(n12505), .ZN(n12504) );
  NAND2_X1 U8720 ( .A1(n12466), .A2(n12368), .ZN(n12506) );
  AND2_X1 U8721 ( .A1(n12524), .A2(n12358), .ZN(n7199) );
  AND2_X1 U8722 ( .A1(n12359), .A2(n12358), .ZN(n12525) );
  NOR2_X1 U8723 ( .A1(n12011), .A2(n12178), .ZN(n7098) );
  NAND2_X1 U8724 ( .A1(n6799), .A2(n6798), .ZN(n6825) );
  NAND2_X1 U8725 ( .A1(n12185), .A2(n12184), .ZN(n6799) );
  INV_X1 U8726 ( .A(n12183), .ZN(n6798) );
  INV_X1 U8727 ( .A(n12186), .ZN(n6871) );
  INV_X1 U8728 ( .A(n12800), .ZN(n12834) );
  INV_X1 U8729 ( .A(n12816), .ZN(n12849) );
  INV_X1 U8730 ( .A(n14777), .ZN(n12542) );
  INV_X1 U8731 ( .A(n11443), .ZN(n12543) );
  NAND2_X1 U8732 ( .A1(n7799), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7803) );
  OR2_X1 U8733 ( .A1(n9984), .A2(n13017), .ZN(n12550) );
  NOR2_X1 U8734 ( .A1(n12197), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n15402) );
  INV_X1 U8735 ( .A(n7340), .ZN(n10435) );
  AND2_X1 U8736 ( .A1(n7340), .A2(n7339), .ZN(n10401) );
  OAI22_X1 U8737 ( .A1(n10430), .A2(n10137), .B1(n10136), .B2(n10431), .ZN(
        n10395) );
  NAND2_X1 U8738 ( .A1(n7444), .A2(n7443), .ZN(n10445) );
  NAND2_X1 U8739 ( .A1(n6991), .A2(n6990), .ZN(n6989) );
  NAND2_X1 U8740 ( .A1(n7358), .A2(n10497), .ZN(n10462) );
  AND3_X1 U8741 ( .A1(n6989), .A2(n10492), .A3(P3_REG2_REG_7__SCAN_IN), .ZN(
        n10493) );
  INV_X1 U8742 ( .A(n10493), .ZN(n6988) );
  INV_X1 U8743 ( .A(n7003), .ZN(n10500) );
  AND2_X1 U8744 ( .A1(n7003), .A2(n7002), .ZN(n10927) );
  XNOR2_X1 U8745 ( .A(n11263), .B(n7439), .ZN(n10917) );
  INV_X1 U8746 ( .A(n7363), .ZN(n15424) );
  INV_X1 U8747 ( .A(n7012), .ZN(n15422) );
  NOR2_X1 U8748 ( .A1(n15416), .A2(n15415), .ZN(n15414) );
  XNOR2_X1 U8749 ( .A(n7436), .B(n11268), .ZN(n11312) );
  NOR2_X1 U8750 ( .A1(n11312), .A2(n11313), .ZN(n11311) );
  XNOR2_X1 U8751 ( .A(n11855), .B(n12564), .ZN(n12552) );
  INV_X1 U8752 ( .A(n7438), .ZN(n12559) );
  NOR2_X1 U8753 ( .A1(n12584), .A2(n12585), .ZN(n12583) );
  NOR2_X1 U8754 ( .A1(n12622), .A2(n11901), .ZN(n12624) );
  XNOR2_X1 U8755 ( .A(n7336), .B(n7335), .ZN(n12621) );
  NAND2_X1 U8756 ( .A1(n12686), .A2(n7084), .ZN(n12894) );
  OR2_X1 U8757 ( .A1(n12687), .A2(n15456), .ZN(n7084) );
  NAND2_X1 U8758 ( .A1(n7459), .A2(n7457), .ZN(n12710) );
  NAND2_X1 U8759 ( .A1(n7085), .A2(n7088), .ZN(n12805) );
  NAND2_X1 U8760 ( .A1(n7998), .A2(n7997), .ZN(n12859) );
  AND2_X1 U8761 ( .A1(n7452), .A2(n7683), .ZN(n14760) );
  NAND2_X1 U8762 ( .A1(n11329), .A2(n7962), .ZN(n7452) );
  NAND2_X1 U8763 ( .A1(n8214), .A2(n12111), .ZN(n14758) );
  AND3_X1 U8764 ( .A1(n7928), .A2(n7927), .A3(n7926), .ZN(n11336) );
  INV_X1 U8765 ( .A(n12885), .ZN(n12867) );
  NAND2_X1 U8766 ( .A1(n11214), .A2(n7899), .ZN(n11141) );
  INV_X1 U8767 ( .A(n12888), .ZN(n12869) );
  NAND2_X1 U8768 ( .A1(n10959), .A2(n12074), .ZN(n10944) );
  AND3_X1 U8769 ( .A1(n7822), .A2(n7821), .A3(n7820), .ZN(n15487) );
  NAND2_X1 U8770 ( .A1(n10124), .A2(n9864), .ZN(n15443) );
  AND2_X1 U8771 ( .A1(n15477), .A2(n15458), .ZN(n15474) );
  NAND2_X1 U8772 ( .A1(n7795), .A2(n6818), .ZN(n10114) );
  OR2_X1 U8773 ( .A1(n8095), .A2(n9334), .ZN(n7795) );
  AOI21_X1 U8774 ( .B1(n6820), .B2(SI_0_), .A(n6819), .ZN(n6818) );
  NOR2_X1 U8775 ( .A1(n10127), .A2(n9335), .ZN(n6819) );
  INV_X1 U8776 ( .A(n15443), .ZN(n15473) );
  AND2_X1 U8777 ( .A1(n15547), .A2(n15488), .ZN(n12951) );
  OR2_X1 U8778 ( .A1(n12656), .A2(n12655), .ZN(n14786) );
  INV_X1 U8779 ( .A(n6864), .ZN(n12966) );
  INV_X1 U8780 ( .A(n12454), .ZN(n12974) );
  INV_X1 U8781 ( .A(n12856), .ZN(n13008) );
  INV_X1 U8782 ( .A(n12360), .ZN(n13015) );
  INV_X1 U8783 ( .A(n7154), .ZN(n13018) );
  INV_X1 U8784 ( .A(n9387), .ZN(n13017) );
  XNOR2_X1 U8785 ( .A(n11997), .B(n11996), .ZN(n13024) );
  INV_X1 U8786 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13019) );
  INV_X1 U8787 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7697) );
  NAND2_X1 U8788 ( .A1(n11995), .A2(n11988), .ZN(n11990) );
  INV_X1 U8789 ( .A(SI_26_), .ZN(n11304) );
  INV_X1 U8790 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8241) );
  NAND2_X1 U8791 ( .A1(n7763), .A2(n11351), .ZN(n7312) );
  NAND2_X1 U8792 ( .A1(n6800), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n7313) );
  NAND2_X1 U8793 ( .A1(n7755), .A2(n7756), .ZN(n8092) );
  INV_X1 U8794 ( .A(n8283), .ZN(n10109) );
  INV_X1 U8795 ( .A(SI_19_), .ZN(n9774) );
  INV_X1 U8796 ( .A(n12014), .ZN(n12039) );
  OAI21_X1 U8797 ( .B1(n8049), .B2(n7291), .A(n7289), .ZN(n8068) );
  NAND2_X1 U8798 ( .A1(n8051), .A2(n7751), .ZN(n8066) );
  INV_X1 U8799 ( .A(SI_16_), .ZN(n9607) );
  NAND2_X1 U8800 ( .A1(n8002), .A2(n7743), .ZN(n8020) );
  INV_X1 U8801 ( .A(SI_15_), .ZN(n9547) );
  OR2_X1 U8802 ( .A1(n8007), .A2(n8036), .ZN(n11896) );
  INV_X1 U8803 ( .A(SI_14_), .ZN(n9377) );
  INV_X1 U8804 ( .A(SI_12_), .ZN(n9367) );
  INV_X1 U8805 ( .A(SI_10_), .ZN(n9340) );
  XNOR2_X1 U8806 ( .A(n7848), .B(P3_IR_REG_5__SCAN_IN), .ZN(n10168) );
  AND2_X1 U8807 ( .A1(n7195), .A2(n10145), .ZN(n7847) );
  AND2_X1 U8808 ( .A1(n8991), .A2(P3_U3151), .ZN(n13380) );
  AND2_X1 U8809 ( .A1(n9394), .A2(n9205), .ZN(n9395) );
  INV_X1 U8810 ( .A(n7500), .ZN(n10586) );
  AOI21_X1 U8811 ( .B1(n10100), .B2(n7503), .A(n6653), .ZN(n7500) );
  NAND2_X1 U8812 ( .A1(n7505), .A2(n7511), .ZN(n13386) );
  AND2_X1 U8813 ( .A1(n13449), .A2(n11949), .ZN(n13396) );
  OAI21_X1 U8814 ( .B1(n13483), .B2(n13482), .A(n7494), .ZN(n13406) );
  NAND2_X1 U8815 ( .A1(n8864), .A2(n8863), .ZN(n13818) );
  AOI21_X1 U8816 ( .B1(n7508), .B2(n7511), .A(n7507), .ZN(n7506) );
  NAND2_X1 U8817 ( .A1(n7511), .A2(n7510), .ZN(n7509) );
  NOR2_X1 U8818 ( .A1(n11965), .A2(n11964), .ZN(n7507) );
  NAND2_X1 U8819 ( .A1(n6839), .A2(n6837), .ZN(n9615) );
  NAND2_X1 U8820 ( .A1(n9669), .A2(n6636), .ZN(n6839) );
  NAND2_X1 U8821 ( .A1(n6838), .A2(n15307), .ZN(n6837) );
  INV_X1 U8822 ( .A(n11968), .ZN(n6838) );
  NAND2_X1 U8823 ( .A1(n9053), .A2(n9052), .ZN(n13785) );
  NAND2_X1 U8824 ( .A1(n7480), .A2(n7483), .ZN(n13465) );
  NAND2_X1 U8825 ( .A1(n13483), .A2(n7485), .ZN(n7480) );
  NAND2_X1 U8826 ( .A1(n8883), .A2(n8882), .ZN(n13813) );
  XNOR2_X1 U8827 ( .A(n11942), .B(n11940), .ZN(n13473) );
  NAND2_X1 U8828 ( .A1(n7523), .A2(n7524), .ZN(n11165) );
  OR2_X1 U8829 ( .A1(n9479), .A2(n9476), .ZN(n13476) );
  NAND2_X1 U8830 ( .A1(n10100), .A2(n10099), .ZN(n10368) );
  NAND2_X1 U8831 ( .A1(n6875), .A2(n7517), .ZN(n7516) );
  INV_X1 U8832 ( .A(n13420), .ZN(n6875) );
  NAND2_X1 U8833 ( .A1(n7516), .A2(n11956), .ZN(n13491) );
  CLKBUF_X1 U8834 ( .A(P2_DATAO_REG_1__SCAN_IN), .Z(n6866) );
  INV_X1 U8835 ( .A(n9646), .ZN(n13533) );
  INV_X1 U8836 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7778) );
  INV_X1 U8837 ( .A(n13569), .ZN(n13760) );
  NAND2_X1 U8838 ( .A1(n11829), .A2(n11828), .ZN(n11830) );
  AND2_X1 U8839 ( .A1(n9057), .A2(n9056), .ZN(n13631) );
  AOI21_X1 U8840 ( .B1(n13662), .B2(n7265), .A(n11824), .ZN(n13637) );
  OR2_X1 U8841 ( .A1(n6911), .A2(n7420), .ZN(n7417) );
  AND2_X1 U8842 ( .A1(n7422), .A2(n7421), .ZN(n13675) );
  AND2_X1 U8843 ( .A1(n13666), .A2(n13665), .ZN(n13802) );
  NAND2_X1 U8844 ( .A1(n7251), .A2(n11816), .ZN(n13724) );
  NAND2_X1 U8845 ( .A1(n11815), .A2(n11814), .ZN(n7251) );
  NAND2_X1 U8846 ( .A1(n14865), .A2(n11572), .ZN(n11573) );
  NAND2_X1 U8847 ( .A1(n8815), .A2(n8814), .ZN(n11923) );
  NAND2_X1 U8848 ( .A1(n14834), .A2(n7428), .ZN(n14865) );
  NAND2_X1 U8849 ( .A1(n14834), .A2(n11570), .ZN(n13752) );
  NAND2_X1 U8850 ( .A1(n7259), .A2(n11578), .ZN(n14839) );
  NAND2_X1 U8851 ( .A1(n11576), .A2(n11575), .ZN(n7259) );
  NAND2_X1 U8852 ( .A1(n8753), .A2(n8752), .ZN(n14849) );
  NAND2_X1 U8853 ( .A1(n10765), .A2(n10764), .ZN(n10996) );
  NAND2_X1 U8854 ( .A1(n10759), .A2(n10758), .ZN(n7222) );
  NAND2_X2 U8855 ( .A1(n8659), .A2(n8658), .ZN(n15369) );
  NAND2_X1 U8856 ( .A1(n7242), .A2(n10240), .ZN(n10290) );
  NAND2_X1 U8857 ( .A1(n9470), .A2(n15305), .ZN(n14827) );
  INV_X1 U8858 ( .A(n10200), .ZN(n15281) );
  OR2_X1 U8859 ( .A1(n15292), .A2(n14825), .ZN(n15282) );
  INV_X1 U8860 ( .A(n15282), .ZN(n14844) );
  INV_X2 U8861 ( .A(n15399), .ZN(n15401) );
  INV_X1 U8862 ( .A(n6900), .ZN(n6899) );
  AND2_X1 U8863 ( .A1(n9466), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15305) );
  INV_X1 U8864 ( .A(n15301), .ZN(n15298) );
  NOR2_X1 U8865 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n7407) );
  CLKBUF_X1 U8866 ( .A(n9192), .Z(n9193) );
  INV_X1 U8867 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n10829) );
  INV_X1 U8868 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10623) );
  INV_X1 U8869 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n9915) );
  INV_X1 U8870 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n9781) );
  INV_X1 U8871 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n13278) );
  INV_X1 U8872 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9444) );
  INV_X1 U8873 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9555) );
  INV_X1 U8874 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9373) );
  INV_X1 U8875 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9350) );
  INV_X1 U8876 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9342) );
  INV_X1 U8877 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9327) );
  INV_X1 U8878 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9337) );
  AND2_X1 U8879 ( .A1(n9587), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9278) );
  NAND2_X1 U8880 ( .A1(n11045), .A2(n6924), .ZN(n6923) );
  INV_X1 U8881 ( .A(n11046), .ZN(n6924) );
  NAND2_X1 U8882 ( .A1(n11642), .A2(n14017), .ZN(n7108) );
  AND4_X1 U8883 ( .A1(n11695), .A2(n11694), .A3(n11693), .A4(n11692), .ZN(
        n14530) );
  NAND2_X1 U8884 ( .A1(n7144), .A2(n12267), .ZN(n13878) );
  NOR2_X1 U8885 ( .A1(n6933), .A2(n10066), .ZN(n9838) );
  AND2_X1 U8886 ( .A1(n9834), .A2(n9833), .ZN(n6933) );
  NAND2_X1 U8887 ( .A1(n11723), .A2(n14017), .ZN(n6964) );
  NAND2_X1 U8888 ( .A1(n14933), .A2(n12227), .ZN(n13897) );
  NAND2_X1 U8889 ( .A1(n7131), .A2(n12313), .ZN(n13906) );
  NAND2_X1 U8890 ( .A1(n13922), .A2(n13923), .ZN(n7131) );
  NAND2_X1 U8891 ( .A1(n6680), .A2(n13993), .ZN(n14917) );
  NAND2_X1 U8892 ( .A1(n7140), .A2(n7141), .ZN(n11065) );
  AND2_X1 U8893 ( .A1(n10521), .A2(n10522), .ZN(n6874) );
  AND2_X1 U8894 ( .A1(n11713), .A2(n11712), .ZN(n14518) );
  NAND2_X1 U8895 ( .A1(n7147), .A2(n7150), .ZN(n7146) );
  INV_X1 U8896 ( .A(n7148), .ZN(n7147) );
  NAND2_X1 U8897 ( .A1(n14930), .A2(n12223), .ZN(n14933) );
  INV_X1 U8898 ( .A(n14271), .ZN(n14924) );
  NAND2_X1 U8899 ( .A1(n9842), .A2(n9841), .ZN(n14932) );
  AOI21_X1 U8900 ( .B1(n7132), .B2(n7134), .A(n6733), .ZN(n7129) );
  NAND2_X1 U8901 ( .A1(n11761), .A2(n11760), .ZN(n14614) );
  INV_X1 U8902 ( .A(n14956), .ZN(n14006) );
  AND4_X1 U8903 ( .A1(n11375), .A2(n11374), .A3(n11373), .A4(n11372), .ZN(
        n13999) );
  INV_X1 U8904 ( .A(n14941), .ZN(n14001) );
  BUF_X1 U8905 ( .A(n14281), .Z(n6932) );
  NAND2_X1 U8906 ( .A1(n14291), .A2(n14290), .ZN(n14289) );
  AND2_X1 U8907 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n14290) );
  AND2_X1 U8908 ( .A1(n9734), .A2(n7024), .ZN(n9754) );
  NAND2_X1 U8909 ( .A1(n9735), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7024) );
  INV_X1 U8910 ( .A(n7023), .ZN(n9752) );
  AND2_X1 U8911 ( .A1(n7023), .A2(n7022), .ZN(n9882) );
  NAND2_X1 U8912 ( .A1(n9748), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n7022) );
  NOR2_X1 U8913 ( .A1(n9740), .A2(n9739), .ZN(n9765) );
  NOR2_X1 U8914 ( .A1(n9893), .A2(n7018), .ZN(n9740) );
  AND2_X1 U8915 ( .A1(n10800), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7018) );
  NOR2_X1 U8916 ( .A1(n9765), .A2(n7017), .ZN(n9769) );
  AND2_X1 U8917 ( .A1(n10853), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7017) );
  NOR2_X1 U8918 ( .A1(n9769), .A2(n9768), .ZN(n9901) );
  INV_X1 U8919 ( .A(n7016), .ZN(n15073) );
  AND2_X1 U8920 ( .A1(n14349), .A2(n6902), .ZN(n14354) );
  INV_X1 U8921 ( .A(n6903), .ZN(n6902) );
  OAI21_X1 U8922 ( .B1(n14351), .B2(n15061), .A(n15100), .ZN(n6903) );
  INV_X1 U8923 ( .A(n14366), .ZN(n14587) );
  NAND2_X1 U8924 ( .A1(n11634), .A2(n11633), .ZN(n14384) );
  NAND2_X1 U8925 ( .A1(n7368), .A2(n7372), .ZN(n14417) );
  OR2_X1 U8926 ( .A1(n14452), .A2(n7374), .ZN(n7368) );
  NAND2_X1 U8927 ( .A1(n7378), .A2(n11756), .ZN(n14441) );
  NAND2_X1 U8928 ( .A1(n7630), .A2(n11784), .ZN(n14436) );
  NAND2_X1 U8929 ( .A1(n6734), .A2(n7399), .ZN(n14465) );
  NAND2_X1 U8930 ( .A1(n11721), .A2(n11720), .ZN(n14654) );
  INV_X1 U8931 ( .A(n14518), .ZN(n14652) );
  NAND2_X1 U8932 ( .A1(n7390), .A2(n7392), .ZN(n14525) );
  NAND2_X1 U8933 ( .A1(n14556), .A2(n7395), .ZN(n7390) );
  NAND2_X1 U8934 ( .A1(n11688), .A2(n11687), .ZN(n14667) );
  NAND2_X1 U8935 ( .A1(n7397), .A2(n11684), .ZN(n14542) );
  NAND2_X1 U8936 ( .A1(n7398), .A2(n6670), .ZN(n7397) );
  INV_X1 U8937 ( .A(n14556), .ZN(n7398) );
  NAND2_X1 U8938 ( .A1(n11677), .A2(n11676), .ZN(n14565) );
  NAND2_X1 U8939 ( .A1(n11669), .A2(n11668), .ZN(n14568) );
  NOR2_X1 U8940 ( .A1(n11541), .A2(n14237), .ZN(n14960) );
  AND2_X1 U8941 ( .A1(n14965), .A2(n11533), .ZN(n11538) );
  AND2_X1 U8942 ( .A1(n9846), .A2(n9824), .ZN(n15114) );
  NOR2_X1 U8943 ( .A1(n7382), .A2(n7386), .ZN(n14731) );
  INV_X1 U8944 ( .A(n7385), .ZN(n7382) );
  NAND2_X1 U8945 ( .A1(n11416), .A2(n11415), .ZN(n11481) );
  OR2_X1 U8946 ( .A1(n15129), .A2(n10573), .ZN(n15116) );
  OR2_X1 U8947 ( .A1(n15129), .A2(n10634), .ZN(n14584) );
  NAND2_X1 U8948 ( .A1(n9952), .A2(n9951), .ZN(n10320) );
  INV_X1 U8949 ( .A(n15114), .ZN(n14578) );
  INV_X1 U8950 ( .A(n14519), .ZN(n15125) );
  INV_X1 U8951 ( .A(n14584), .ZN(n14516) );
  INV_X1 U8952 ( .A(n15116), .ZN(n14737) );
  OAI21_X1 U8953 ( .B1(n9935), .B2(n10667), .A(n10635), .ZN(n14219) );
  NAND2_X1 U8954 ( .A1(n9108), .A2(n9107), .ZN(n14026) );
  MUX2_X1 U8955 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9252), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n9255) );
  CLKBUF_X1 U8956 ( .A(n9265), .Z(n14254) );
  NAND2_X1 U8957 ( .A1(n9228), .A2(n6669), .ZN(n11468) );
  OAI21_X1 U8958 ( .B1(n11735), .B2(n7575), .A(n8950), .ZN(n8965) );
  NAND2_X1 U8959 ( .A1(n6810), .A2(n9233), .ZN(n6808) );
  INV_X1 U8960 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n13291) );
  OAI21_X1 U8961 ( .B1(n10118), .B2(P1_IR_REG_18__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9822) );
  INV_X1 U8962 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n9876) );
  INV_X1 U8963 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n9779) );
  INV_X1 U8964 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n9703) );
  INV_X1 U8965 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9488) );
  INV_X1 U8966 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9552) );
  INV_X1 U8967 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n13149) );
  INV_X1 U8968 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10552) );
  NAND2_X1 U8969 ( .A1(n8525), .A2(n8527), .ZN(n6952) );
  NAND2_X1 U8970 ( .A1(n7364), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9292) );
  INV_X1 U8971 ( .A(n9210), .ZN(n7364) );
  NAND2_X1 U8972 ( .A1(n8473), .A2(n8488), .ZN(n8489) );
  NAND2_X1 U8973 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n7013) );
  AOI21_X1 U8974 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n8355), .A(n15558), .ZN(
        n15550) );
  XNOR2_X1 U8975 ( .A(n8360), .B(n6835), .ZN(n15553) );
  INV_X1 U8976 ( .A(n8359), .ZN(n6835) );
  NOR2_X1 U8977 ( .A1(n14727), .A2(n14728), .ZN(n14726) );
  XNOR2_X1 U8978 ( .A(n8379), .B(n7276), .ZN(n14991) );
  INV_X1 U8979 ( .A(n8380), .ZN(n7276) );
  NAND2_X1 U8980 ( .A1(n14991), .A2(n14990), .ZN(n14989) );
  INV_X1 U8981 ( .A(n8386), .ZN(n8384) );
  INV_X1 U8982 ( .A(n7280), .ZN(n14702) );
  AND2_X1 U8983 ( .A1(n12422), .A2(n12421), .ZN(n7172) );
  NAND2_X1 U8984 ( .A1(n7158), .A2(n12522), .ZN(n7157) );
  INV_X1 U8985 ( .A(n7361), .ZN(n11262) );
  INV_X1 U8986 ( .A(n7334), .ZN(n12569) );
  INV_X1 U8987 ( .A(n7009), .ZN(n12603) );
  XNOR2_X1 U8988 ( .A(n6997), .B(n12637), .ZN(n12654) );
  NAND2_X1 U8989 ( .A1(n7432), .A2(n15404), .ZN(n6992) );
  INV_X1 U8990 ( .A(n6994), .ZN(n6993) );
  AOI21_X1 U8991 ( .B1(n12205), .B2(n12885), .A(n12204), .ZN(n6821) );
  NAND2_X1 U8992 ( .A1(n7471), .A2(n6771), .ZN(P3_U3488) );
  NAND2_X1 U8993 ( .A1(n8293), .A2(n15547), .ZN(n7471) );
  INV_X1 U8994 ( .A(n6905), .ZN(n6904) );
  OAI22_X1 U8995 ( .A1(n12963), .A2(n12957), .B1(n15547), .B2(n12893), .ZN(
        n6905) );
  OAI21_X1 U8996 ( .B1(n8293), .B2(n15526), .A(n8292), .ZN(n8295) );
  INV_X1 U8997 ( .A(n6907), .ZN(n6906) );
  OAI22_X1 U8998 ( .A1(n12963), .A2(n13014), .B1(n15528), .B2(n12962), .ZN(
        n6907) );
  NAND2_X1 U8999 ( .A1(n7082), .A2(n7080), .ZN(P3_U3454) );
  INV_X1 U9000 ( .A(n7081), .ZN(n7080) );
  OR2_X1 U9001 ( .A1(n12964), .A2(n7083), .ZN(n7082) );
  OAI22_X1 U9002 ( .A1(n12966), .A2(n13014), .B1(n15528), .B2(n12965), .ZN(
        n7081) );
  NOR2_X1 U9003 ( .A1(n9200), .A2(n7679), .ZN(n9201) );
  OR2_X1 U9004 ( .A1(n15202), .A2(n6958), .ZN(n6957) );
  NAND2_X1 U9005 ( .A1(n14674), .A2(n15202), .ZN(n6959) );
  INV_X1 U9006 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6958) );
  INV_X1 U9007 ( .A(n6856), .ZN(n14998) );
  NOR2_X1 U9008 ( .A1(n14755), .A2(n14756), .ZN(n14754) );
  INV_X1 U9009 ( .A(n6930), .ZN(n14755) );
  NAND2_X1 U9010 ( .A1(n6855), .A2(n6716), .ZN(n6854) );
  AND2_X1 U9011 ( .A1(n10365), .A2(n10366), .ZN(n6653) );
  INV_X1 U9012 ( .A(n10431), .ZN(n10150) );
  INV_X1 U9013 ( .A(n9121), .ZN(n8574) );
  AND2_X1 U9014 ( .A1(n7669), .A2(n7065), .ZN(n6655) );
  AND2_X1 U9015 ( .A1(n14515), .A2(n6667), .ZN(n6656) );
  INV_X1 U9016 ( .A(n10132), .ZN(n12187) );
  OR2_X1 U9017 ( .A1(n7590), .A2(n7113), .ZN(n6657) );
  AND4_X2 U9018 ( .A1(n9947), .A2(n9946), .A3(n9945), .A4(n9944), .ZN(n10515)
         );
  AND2_X1 U9019 ( .A1(n7694), .A2(n7201), .ZN(n6658) );
  NAND2_X1 U9020 ( .A1(n11394), .A2(n11393), .ZN(n14112) );
  INV_X1 U9021 ( .A(n14112), .ZN(n7609) );
  AND2_X2 U9022 ( .A1(n14845), .A2(n11569), .ZN(n6659) );
  INV_X1 U9023 ( .A(n14515), .ZN(n11720) );
  OAI21_X1 U9024 ( .B1(n12305), .B2(n14626), .A(n14438), .ZN(n14418) );
  INV_X1 U9025 ( .A(n14418), .ZN(n7618) );
  AND2_X1 U9026 ( .A1(n8553), .A2(n8528), .ZN(n6660) );
  NAND2_X1 U9027 ( .A1(n9034), .A2(n9033), .ZN(n13779) );
  OR2_X1 U9028 ( .A1(n8927), .A2(SI_21_), .ZN(n6661) );
  OR2_X1 U9029 ( .A1(n8833), .A2(SI_17_), .ZN(n6662) );
  AND2_X1 U9030 ( .A1(n7159), .A2(n6723), .ZN(n6663) );
  AND2_X1 U9031 ( .A1(n7609), .A2(n14268), .ZN(n6664) );
  NAND2_X1 U9032 ( .A1(n7085), .A2(n8219), .ZN(n6665) );
  INV_X1 U9033 ( .A(n7401), .ZN(n7400) );
  INV_X1 U9034 ( .A(n13686), .ZN(n6850) );
  AND2_X1 U9035 ( .A1(n13795), .A2(n11823), .ZN(n11824) );
  INV_X1 U9036 ( .A(n10499), .ZN(n7002) );
  AND2_X1 U9037 ( .A1(n7440), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n6666) );
  INV_X1 U9038 ( .A(n14730), .ZN(n7384) );
  NOR2_X1 U9039 ( .A1(n7604), .A2(n7599), .ZN(n7598) );
  OR2_X1 U9040 ( .A1(n14534), .A2(n14545), .ZN(n6667) );
  BUF_X1 U9041 ( .A(n11715), .Z(n11775) );
  OR2_X1 U9042 ( .A1(n10118), .A2(n9227), .ZN(n6669) );
  INV_X1 U9043 ( .A(n10089), .ZN(n12379) );
  OAI211_X1 U9044 ( .C1(n6845), .C2(n9963), .A(n9962), .B(n9961), .ZN(n14053)
         );
  NAND2_X1 U9045 ( .A1(n9209), .A2(n9210), .ZN(n9283) );
  OR2_X1 U9046 ( .A1(n14565), .A2(n14574), .ZN(n6670) );
  XOR2_X1 U9047 ( .A(n6824), .B(n12014), .Z(n6671) );
  NAND4_X1 U9048 ( .A1(n7612), .A2(n7152), .A3(n7151), .A4(n6668), .ZN(n6672)
         );
  INV_X1 U9049 ( .A(n14245), .ZN(n6960) );
  OR2_X1 U9050 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6673) );
  AND2_X1 U9051 ( .A1(n10841), .A2(n7192), .ZN(n6674) );
  CLKBUF_X3 U9052 ( .A(n8991), .Z(n6832) );
  INV_X1 U9053 ( .A(n6972), .ZN(n6971) );
  NAND2_X1 U9054 ( .A1(n6974), .A2(n8717), .ZN(n6972) );
  OR2_X1 U9055 ( .A1(n12564), .A2(n11893), .ZN(n6675) );
  AND2_X1 U9056 ( .A1(n14237), .A2(n11533), .ZN(n6676) );
  AND2_X1 U9057 ( .A1(n8601), .A2(n8600), .ZN(n6677) );
  AND2_X1 U9058 ( .A1(n14181), .A2(n14180), .ZN(n6678) );
  AND2_X1 U9059 ( .A1(n14104), .A2(n14103), .ZN(n6679) );
  AND2_X1 U9060 ( .A1(n14915), .A2(n14914), .ZN(n6680) );
  INV_X1 U9061 ( .A(n8625), .ZN(n6844) );
  NAND2_X1 U9062 ( .A1(n13773), .A2(n13493), .ZN(n6681) );
  OR2_X1 U9063 ( .A1(n13490), .A2(n7515), .ZN(n7514) );
  AND2_X1 U9064 ( .A1(n12077), .A2(n7077), .ZN(n6682) );
  XOR2_X1 U9065 ( .A(n13566), .B(n9112), .Z(n6683) );
  INV_X1 U9066 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n8298) );
  NAND2_X1 U9067 ( .A1(n9017), .A2(n9016), .ZN(n13773) );
  INV_X1 U9068 ( .A(n13773), .ZN(n7322) );
  AND2_X1 U9069 ( .A1(n7417), .A2(n7419), .ZN(n6684) );
  INV_X1 U9070 ( .A(n14835), .ZN(n6847) );
  INV_X1 U9071 ( .A(n14495), .ZN(n14241) );
  INV_X1 U9072 ( .A(n14759), .ZN(n7451) );
  NAND2_X1 U9073 ( .A1(n8952), .A2(n8951), .ZN(n13795) );
  INV_X1 U9074 ( .A(n13795), .ZN(n7316) );
  AND3_X1 U9075 ( .A1(n12669), .A2(n12681), .A3(n12708), .ZN(n6685) );
  AND4_X1 U9076 ( .A1(n7690), .A2(n7689), .A3(n8005), .A4(n7987), .ZN(n6686)
         );
  AND2_X1 U9077 ( .A1(n12895), .A2(n15517), .ZN(n6687) );
  NAND2_X1 U9078 ( .A1(n8773), .A2(n8772), .ZN(n14830) );
  OR2_X1 U9079 ( .A1(n14079), .A2(n14272), .ZN(n6688) );
  OR2_X1 U9080 ( .A1(n6845), .A2(n14308), .ZN(n6689) );
  INV_X1 U9081 ( .A(n14111), .ZN(n7558) );
  AND2_X1 U9082 ( .A1(n14849), .A2(n11579), .ZN(n6690) );
  AND2_X1 U9083 ( .A1(n7316), .A2(n13512), .ZN(n6691) );
  INV_X1 U9084 ( .A(n8806), .ZN(n7030) );
  AND2_X1 U9085 ( .A1(n7378), .A2(n7376), .ZN(n6692) );
  OR2_X1 U9086 ( .A1(n11737), .A2(n9802), .ZN(n6693) );
  AOI21_X1 U9087 ( .B1(n11772), .B2(n14017), .A(n11771), .ZN(n14593) );
  AND3_X1 U9088 ( .A1(n7802), .A2(n7801), .A3(n7804), .ZN(n6694) );
  AND2_X1 U9089 ( .A1(n14614), .A2(n13910), .ZN(n6695) );
  AND2_X1 U9090 ( .A1(n13822), .A2(n11817), .ZN(n6696) );
  NOR2_X1 U9091 ( .A1(n14278), .A2(n14053), .ZN(n6697) );
  INV_X1 U9092 ( .A(n15307), .ZN(n9614) );
  AND3_X1 U9093 ( .A1(n7540), .A2(n7545), .A3(n7539), .ZN(n6698) );
  OR2_X1 U9094 ( .A1(n12749), .A2(n12754), .ZN(n12153) );
  NOR2_X1 U9095 ( .A1(n12583), .A2(n11897), .ZN(n6699) );
  NOR2_X1 U9096 ( .A1(n12624), .A2(n11903), .ZN(n6700) );
  OR2_X1 U9097 ( .A1(n14614), .A2(n14421), .ZN(n14406) );
  OR2_X1 U9098 ( .A1(n11468), .A2(n14696), .ZN(n6701) );
  AND2_X1 U9099 ( .A1(n12414), .A2(n12514), .ZN(n6702) );
  INV_X1 U9100 ( .A(n13404), .ZN(n7493) );
  AOI21_X1 U9101 ( .B1(n8563), .B2(n8566), .A(n8584), .ZN(n7117) );
  AND2_X1 U9102 ( .A1(n12223), .A2(n7150), .ZN(n6703) );
  AND2_X1 U9103 ( .A1(n11785), .A2(n11758), .ZN(n14420) );
  AND2_X1 U9104 ( .A1(n12454), .A2(n12727), .ZN(n6704) );
  AND2_X1 U9105 ( .A1(n7115), .A2(n8586), .ZN(n6705) );
  NAND4_X1 U9106 ( .A1(n6749), .A2(n7696), .A3(n13256), .A4(n7695), .ZN(n6706)
         );
  INV_X1 U9107 ( .A(n14171), .ZN(n7565) );
  INV_X1 U9108 ( .A(n14179), .ZN(n7563) );
  AND2_X1 U9109 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n6707) );
  NAND2_X1 U9110 ( .A1(n10583), .A2(n10584), .ZN(n6708) );
  INV_X1 U9111 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6836) );
  OR2_X1 U9112 ( .A1(n8852), .A2(n8851), .ZN(n6709) );
  AND2_X1 U9113 ( .A1(n10292), .A2(n10291), .ZN(n6710) );
  AND2_X1 U9114 ( .A1(n11170), .A2(n13523), .ZN(n6711) );
  INV_X1 U9115 ( .A(n7610), .ZN(n7599) );
  NAND2_X1 U9116 ( .A1(n14746), .A2(n14269), .ZN(n7610) );
  AND2_X1 U9117 ( .A1(n8491), .A2(n6857), .ZN(n6712) );
  OR2_X1 U9118 ( .A1(n14956), .A2(n14912), .ZN(n14123) );
  AND2_X1 U9119 ( .A1(n8438), .A2(n7639), .ZN(n6713) );
  INV_X1 U9120 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7201) );
  INV_X1 U9121 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6810) );
  NAND2_X1 U9122 ( .A1(n14756), .A2(n7281), .ZN(n6714) );
  AND2_X1 U9123 ( .A1(n14518), .A2(n14498), .ZN(n6715) );
  OR2_X1 U9124 ( .A1(n7280), .A2(n7279), .ZN(n6716) );
  AND2_X1 U9125 ( .A1(n12336), .A2(n12335), .ZN(n6717) );
  AND2_X1 U9126 ( .A1(n11609), .A2(n12540), .ZN(n6718) );
  AND2_X1 U9127 ( .A1(n8692), .A2(n9340), .ZN(n6719) );
  NOR2_X1 U9128 ( .A1(n14078), .A2(n14272), .ZN(n6720) );
  NOR2_X1 U9129 ( .A1(n14644), .A2(n14506), .ZN(n6721) );
  NOR2_X1 U9130 ( .A1(n7652), .A2(n6728), .ZN(n6722) );
  NAND2_X1 U9131 ( .A1(n14480), .A2(n14461), .ZN(n14453) );
  INV_X1 U9132 ( .A(n14453), .ZN(n7205) );
  INV_X1 U9133 ( .A(n7486), .ZN(n7485) );
  NAND2_X1 U9134 ( .A1(n7493), .A2(n7494), .ZN(n7486) );
  NAND2_X1 U9135 ( .A1(n7168), .A2(n7164), .ZN(n6723) );
  INV_X1 U9136 ( .A(n8696), .ZN(n7574) );
  AND2_X1 U9137 ( .A1(n6919), .A2(n6917), .ZN(n6724) );
  AND2_X1 U9138 ( .A1(n7459), .A2(n7460), .ZN(n6725) );
  OR2_X1 U9139 ( .A1(n8518), .A2(n8517), .ZN(n6726) );
  AND3_X1 U9140 ( .A1(n9260), .A2(n9262), .A3(n9263), .ZN(n6727) );
  AND2_X1 U9141 ( .A1(n8687), .A2(n8686), .ZN(n6728) );
  INV_X1 U9142 ( .A(n7484), .ZN(n7483) );
  NOR2_X1 U9143 ( .A1(n7487), .A2(n13404), .ZN(n7484) );
  INV_X1 U9144 ( .A(n11824), .ZN(n7267) );
  AND2_X1 U9145 ( .A1(n9104), .A2(n9103), .ZN(n6729) );
  INV_X1 U9146 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9237) );
  AND2_X1 U9147 ( .A1(n8783), .A2(n8782), .ZN(n6730) );
  AND2_X1 U9148 ( .A1(n8718), .A2(n9367), .ZN(n6731) );
  INV_X1 U9149 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9213) );
  NAND2_X1 U9150 ( .A1(n7062), .A2(n7061), .ZN(n6732) );
  AND2_X1 U9151 ( .A1(n12074), .A2(n12075), .ZN(n12018) );
  INV_X1 U9152 ( .A(n12018), .ZN(n7078) );
  AND2_X1 U9153 ( .A1(n12320), .A2(n12319), .ZN(n6733) );
  INV_X1 U9154 ( .A(n7616), .ZN(n7615) );
  NAND2_X1 U9155 ( .A1(n14402), .A2(n7617), .ZN(n7616) );
  OR2_X1 U9156 ( .A1(n7400), .A2(n11721), .ZN(n6734) );
  OR2_X1 U9157 ( .A1(n7535), .A2(n14192), .ZN(n6735) );
  OR2_X1 U9158 ( .A1(n8421), .A2(n8420), .ZN(n6736) );
  NOR2_X1 U9159 ( .A1(n6844), .A2(n8626), .ZN(n6737) );
  OR2_X1 U9160 ( .A1(n7030), .A2(n7579), .ZN(n6738) );
  INV_X1 U9161 ( .A(n7598), .ZN(n7597) );
  NOR3_X1 U9162 ( .A1(n14135), .A2(n14134), .A3(n14141), .ZN(n6739) );
  INV_X1 U9163 ( .A(n14185), .ZN(n7127) );
  AND2_X1 U9164 ( .A1(n7503), .A2(n10585), .ZN(n6740) );
  AND2_X1 U9165 ( .A1(n7419), .A2(n11842), .ZN(n6741) );
  NAND2_X1 U9166 ( .A1(n8795), .A2(n8794), .ZN(n13750) );
  AND2_X1 U9167 ( .A1(n6973), .A2(n6974), .ZN(n6742) );
  AND2_X1 U9168 ( .A1(n8668), .A2(n8667), .ZN(n6743) );
  NOR2_X1 U9169 ( .A1(n14902), .A2(n14903), .ZN(n6744) );
  INV_X1 U9170 ( .A(n14226), .ZN(n10871) );
  NOR2_X1 U9171 ( .A1(n11939), .A2(n7491), .ZN(n6745) );
  NOR2_X1 U9172 ( .A1(n14960), .A2(n11780), .ZN(n6746) );
  NAND2_X1 U9173 ( .A1(n12838), .A2(n12818), .ZN(n6747) );
  OR2_X1 U9174 ( .A1(n7322), .A2(n13493), .ZN(n6748) );
  AND2_X1 U9175 ( .A1(n8193), .A2(n8191), .ZN(n6749) );
  AND2_X1 U9176 ( .A1(n8176), .A2(n8161), .ZN(n6750) );
  AND2_X1 U9177 ( .A1(n6822), .A2(n6821), .ZN(n6751) );
  AND2_X1 U9178 ( .A1(n12145), .A2(n12146), .ZN(n6752) );
  OR2_X1 U9179 ( .A1(n8786), .A2(n6730), .ZN(n6753) );
  AND2_X1 U9180 ( .A1(n7188), .A2(n12376), .ZN(n6754) );
  OR2_X1 U9181 ( .A1(n7558), .A2(n14110), .ZN(n6755) );
  INV_X1 U9182 ( .A(n7393), .ZN(n7392) );
  OAI21_X1 U9183 ( .B1(n7394), .B2(n6670), .A(n11697), .ZN(n7393) );
  OR2_X1 U9184 ( .A1(n7565), .A2(n14170), .ZN(n6756) );
  OR2_X1 U9185 ( .A1(n7563), .A2(n14178), .ZN(n6757) );
  INV_X1 U9186 ( .A(n7611), .ZN(n7608) );
  NAND2_X1 U9187 ( .A1(n15188), .A2(n14271), .ZN(n7611) );
  AND2_X1 U9188 ( .A1(n7570), .A2(n7567), .ZN(n6758) );
  AND2_X1 U9189 ( .A1(n8452), .A2(n7224), .ZN(n6759) );
  INV_X1 U9190 ( .A(n7514), .ZN(n7513) );
  OR2_X1 U9191 ( .A1(n14122), .A2(n7543), .ZN(n6760) );
  NAND2_X1 U9192 ( .A1(n9087), .A2(n7040), .ZN(n6761) );
  AND2_X1 U9193 ( .A1(n14278), .A2(n14053), .ZN(n6762) );
  NAND2_X1 U9194 ( .A1(n7553), .A2(n14073), .ZN(n6763) );
  INV_X1 U9195 ( .A(n8526), .ZN(n7582) );
  AND2_X1 U9196 ( .A1(n7628), .A2(n6667), .ZN(n6764) );
  INV_X1 U9197 ( .A(n10525), .ZN(n12242) );
  INV_X1 U9198 ( .A(n12431), .ZN(n12546) );
  INV_X1 U9199 ( .A(n10929), .ZN(n7439) );
  INV_X1 U9200 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6942) );
  INV_X1 U9201 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7649) );
  OR2_X1 U9202 ( .A1(n14576), .A2(n14565), .ZN(n6765) );
  INV_X1 U9203 ( .A(n6866), .ZN(n6944) );
  AND2_X1 U9204 ( .A1(n14241), .A2(n11722), .ZN(n7401) );
  INV_X1 U9205 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n7036) );
  INV_X1 U9206 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6913) );
  AND2_X1 U9207 ( .A1(n11378), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6766) );
  AND2_X1 U9208 ( .A1(n10928), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n6767) );
  AND4_X1 U9209 ( .A1(n9208), .A2(n9210), .A3(n6668), .A4(n9485), .ZN(n6768)
         );
  INV_X1 U9210 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9751) );
  NAND2_X1 U9211 ( .A1(n9094), .A2(n9093), .ZN(n13762) );
  INV_X1 U9212 ( .A(n13762), .ZN(n7320) );
  AND4_X1 U9213 ( .A1(n9008), .A2(n9007), .A3(n9006), .A4(n9005), .ZN(n13387)
         );
  AND2_X1 U9214 ( .A1(n14933), .A2(n7148), .ZN(n6769) );
  AND2_X1 U9215 ( .A1(n12272), .A2(n12267), .ZN(n6770) );
  INV_X1 U9216 ( .A(n7395), .ZN(n7394) );
  NOR2_X1 U9217 ( .A1(n11696), .A2(n7396), .ZN(n7395) );
  AND4_X1 U9218 ( .A1(n9045), .A2(n9044), .A3(n9043), .A4(n9042), .ZN(n13421)
         );
  INV_X1 U9219 ( .A(n13421), .ZN(n13509) );
  AND2_X1 U9220 ( .A1(n8279), .A2(n8278), .ZN(n6771) );
  OR2_X1 U9221 ( .A1(n12239), .A2(n12238), .ZN(n6772) );
  OR2_X1 U9222 ( .A1(n8855), .A2(n7123), .ZN(n6773) );
  INV_X1 U9223 ( .A(n7326), .ZN(n13746) );
  NOR2_X1 U9224 ( .A1(n14850), .A2(n7327), .ZN(n7326) );
  NOR2_X1 U9225 ( .A1(n8770), .A2(P2_IR_REG_15__SCAN_IN), .ZN(n8791) );
  OR2_X1 U9226 ( .A1(n7575), .A2(n8964), .ZN(n6774) );
  INV_X1 U9227 ( .A(n13462), .ZN(n7492) );
  OR2_X1 U9228 ( .A1(n8924), .A2(SI_20_), .ZN(n6775) );
  AND2_X1 U9229 ( .A1(n12397), .A2(n12398), .ZN(n6776) );
  AND2_X1 U9230 ( .A1(n8966), .A2(SI_23_), .ZN(n6777) );
  AND2_X1 U9231 ( .A1(n8945), .A2(n8944), .ZN(n6778) );
  NAND2_X1 U9232 ( .A1(n10458), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n6779) );
  NAND2_X1 U9233 ( .A1(n9922), .A2(n9923), .ZN(n10100) );
  INV_X1 U9234 ( .A(n12520), .ZN(n12522) );
  INV_X1 U9235 ( .A(n15528), .ZN(n7083) );
  NOR2_X1 U9236 ( .A1(n8427), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n9151) );
  AND2_X1 U9237 ( .A1(n15405), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n6780) );
  INV_X1 U9238 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n7567) );
  AND2_X1 U9239 ( .A1(n11931), .A2(n11930), .ZN(n6781) );
  AND2_X1 U9240 ( .A1(n7347), .A2(n7345), .ZN(n6782) );
  INV_X1 U9241 ( .A(n11282), .ZN(n11892) );
  AND2_X1 U9242 ( .A1(n7955), .A2(n7986), .ZN(n11282) );
  INV_X1 U9243 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7277) );
  AND2_X1 U9244 ( .A1(n7523), .A2(n7521), .ZN(n6783) );
  NOR2_X1 U9245 ( .A1(n9068), .A2(n7587), .ZN(n7586) );
  INV_X1 U9246 ( .A(n7202), .ZN(n11121) );
  OR2_X1 U9247 ( .A1(n6780), .A2(n7431), .ZN(n6784) );
  NAND2_X1 U9248 ( .A1(n8450), .A2(n8555), .ZN(n6785) );
  INV_X1 U9249 ( .A(n7683), .ZN(n7453) );
  INV_X1 U9250 ( .A(n15425), .ZN(n7353) );
  INV_X1 U9251 ( .A(n12633), .ZN(n7335) );
  NAND2_X1 U9252 ( .A1(n8573), .A2(n8572), .ZN(n10292) );
  INV_X1 U9253 ( .A(n10292), .ZN(n7314) );
  INV_X1 U9254 ( .A(n10359), .ZN(n6842) );
  INV_X1 U9255 ( .A(n11864), .ZN(n7352) );
  AND2_X2 U9256 ( .A1(n9863), .A2(n8277), .ZN(n15547) );
  INV_X1 U9257 ( .A(n11887), .ZN(n12644) );
  AND2_X1 U9258 ( .A1(n15067), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6786) );
  NOR2_X1 U9259 ( .A1(n10415), .A2(n10155), .ZN(n6787) );
  NOR2_X1 U9260 ( .A1(n10419), .A2(n10170), .ZN(n6788) );
  AND2_X1 U9261 ( .A1(n10497), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n6789) );
  NAND2_X1 U9262 ( .A1(n10461), .A2(n10502), .ZN(n10497) );
  INV_X1 U9263 ( .A(n10497), .ZN(n7001) );
  AND2_X1 U9264 ( .A1(n7358), .A2(n6789), .ZN(n6790) );
  AND2_X1 U9265 ( .A1(n11911), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6791) );
  NOR2_X1 U9266 ( .A1(n7769), .A2(n7305), .ZN(n7304) );
  AND2_X1 U9267 ( .A1(n6988), .A2(n10492), .ZN(n6792) );
  INV_X1 U9268 ( .A(n13538), .ZN(n6858) );
  INV_X1 U9269 ( .A(n10502), .ZN(n6990) );
  INV_X1 U9270 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6834) );
  INV_X1 U9271 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7274) );
  INV_X1 U9272 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n7435) );
  INV_X1 U9273 ( .A(n15109), .ZN(n11791) );
  INV_X1 U9274 ( .A(n8948), .ZN(n7575) );
  INV_X1 U9275 ( .A(n14971), .ZN(n15109) );
  NOR2_X2 U9276 ( .A1(n10194), .A2(n6843), .ZN(n15285) );
  NAND2_X1 U9277 ( .A1(n12853), .A2(n12852), .ZN(n12838) );
  AOI21_X2 U9278 ( .B1(n12694), .B2(n8227), .A(n8226), .ZN(n12682) );
  NAND2_X1 U9279 ( .A1(n12721), .A2(n12155), .ZN(n12709) );
  NAND2_X1 U9280 ( .A1(n12873), .A2(n8218), .ZN(n12864) );
  OR2_X2 U9281 ( .A1(n7775), .A2(n8069), .ZN(n7777) );
  AND2_X2 U9282 ( .A1(n8070), .A2(n7475), .ZN(n7775) );
  NAND2_X1 U9283 ( .A1(n11202), .A2(n11201), .ZN(n11204) );
  NAND2_X1 U9284 ( .A1(n10069), .A2(n10070), .ZN(n10520) );
  NAND2_X1 U9285 ( .A1(n6926), .A2(n6925), .ZN(n11355) );
  NOR2_X2 U9286 ( .A1(n10543), .A2(n6874), .ZN(n11032) );
  NAND2_X1 U9287 ( .A1(n11050), .A2(n11049), .ZN(n11202) );
  OAI22_X1 U9288 ( .A1(n10072), .A2(n9270), .B1(n12340), .B2(n9972), .ZN(n9832) );
  NAND2_X1 U9289 ( .A1(n11497), .A2(n11496), .ZN(n11502) );
  NAND2_X1 U9290 ( .A1(n6936), .A2(n6935), .ZN(n13940) );
  NAND2_X1 U9291 ( .A1(n7145), .A2(n7146), .ZN(n13942) );
  AOI211_X2 U9292 ( .C1(n14608), .C2(n14955), .A(n14607), .B(n14606), .ZN(
        n14611) );
  NAND2_X2 U9293 ( .A1(n14577), .A2(n14951), .ZN(n14576) );
  AND2_X2 U9294 ( .A1(n10575), .A2(n13978), .ZN(n10805) );
  NAND2_X1 U9295 ( .A1(n11482), .A2(n11515), .ZN(n14739) );
  NAND2_X1 U9296 ( .A1(n14518), .A2(n14535), .ZN(n14517) );
  INV_X1 U9297 ( .A(n8650), .ZN(n6797) );
  OAI22_X1 U9298 ( .A1(n7068), .A2(n7069), .B1(n8804), .B2(n8805), .ZN(n8827)
         );
  INV_X1 U9299 ( .A(n8582), .ZN(n6793) );
  AOI21_X1 U9300 ( .B1(n6761), .B2(n7071), .A(n9149), .ZN(n9181) );
  NAND3_X1 U9301 ( .A1(n8434), .A2(n8555), .A3(n8408), .ZN(n8720) );
  AND4_X2 U9302 ( .A1(n8407), .A2(n8405), .A3(n8406), .A4(n8404), .ZN(n8434)
         );
  NAND3_X1 U9303 ( .A1(n7672), .A2(n6726), .A3(n7673), .ZN(n7671) );
  INV_X1 U9304 ( .A(n8421), .ZN(n8422) );
  AND2_X2 U9305 ( .A1(n6794), .A2(n9571), .ZN(n9570) );
  AND2_X1 U9306 ( .A1(n14832), .A2(n10827), .ZN(n6794) );
  NOR2_X1 U9307 ( .A1(n8923), .A2(n7647), .ZN(n7056) );
  NAND2_X1 U9308 ( .A1(n7650), .A2(n7651), .ZN(n7682) );
  NAND2_X1 U9309 ( .A1(n8831), .A2(n8830), .ZN(n8852) );
  NAND2_X1 U9310 ( .A1(n8743), .A2(n8742), .ZN(n8764) );
  NAND2_X1 U9311 ( .A1(n6801), .A2(n6867), .ZN(n12156) );
  NAND2_X1 U9312 ( .A1(n6868), .A2(n6869), .ZN(n6801) );
  NAND2_X1 U9313 ( .A1(n7896), .A2(n7895), .ZN(n6802) );
  NAND2_X1 U9314 ( .A1(n14723), .A2(n11998), .ZN(n6803) );
  NAND3_X1 U9315 ( .A1(n6805), .A2(n12175), .A3(n12037), .ZN(n6804) );
  XNOR2_X1 U9316 ( .A(n8129), .B(n11813), .ZN(n11107) );
  NAND2_X1 U9317 ( .A1(n7983), .A2(n7982), .ZN(n7985) );
  NAND2_X1 U9318 ( .A1(n7054), .A2(n6709), .ZN(n8878) );
  INV_X1 U9319 ( .A(n7331), .ZN(n7330) );
  NAND2_X1 U9320 ( .A1(n7760), .A2(n7759), .ZN(n8117) );
  NAND2_X1 U9321 ( .A1(n7044), .A2(n7041), .ZN(n8518) );
  NAND2_X1 U9322 ( .A1(n8094), .A2(n7758), .ZN(n8107) );
  OAI21_X1 U9323 ( .B1(n8480), .B2(n8479), .A(n8478), .ZN(n7049) );
  OAI21_X1 U9324 ( .B1(n7941), .B2(n7735), .A(n7736), .ZN(n7957) );
  AOI21_X1 U9325 ( .B1(n14051), .B2(n14052), .A(n7554), .ZN(n14056) );
  INV_X1 U9326 ( .A(n9950), .ZN(n15179) );
  INV_X1 U9327 ( .A(n14096), .ZN(n6812) );
  NAND2_X1 U9328 ( .A1(n14153), .A2(n14152), .ZN(n14156) );
  NAND2_X1 U9329 ( .A1(n6812), .A2(n6811), .ZN(n14101) );
  NAND2_X1 U9330 ( .A1(n6727), .A2(n9261), .ZN(n9935) );
  INV_X1 U9331 ( .A(n14095), .ZN(n6811) );
  NAND2_X1 U9332 ( .A1(n14101), .A2(n14102), .ZN(n14099) );
  NAND2_X1 U9333 ( .A1(n6817), .A2(n6816), .ZN(n14184) );
  INV_X1 U9334 ( .A(n14182), .ZN(n6817) );
  NAND3_X1 U9335 ( .A1(n6814), .A2(n6813), .A3(n6757), .ZN(n7561) );
  NAND2_X1 U9336 ( .A1(n14177), .A2(n14176), .ZN(n6813) );
  NAND2_X1 U9337 ( .A1(n14173), .A2(n14172), .ZN(n6814) );
  NAND2_X1 U9338 ( .A1(n6815), .A2(n7564), .ZN(n14174) );
  NAND3_X1 U9339 ( .A1(n14169), .A2(n14168), .A3(n6756), .ZN(n6815) );
  OAI21_X1 U9340 ( .B1(n14115), .B2(n14114), .A(n14113), .ZN(n14117) );
  MUX2_X1 U9341 ( .A(n7556), .B(n7555), .S(n6639), .Z(n7554) );
  NAND2_X2 U9342 ( .A1(n11230), .A2(n14777), .ZN(n11342) );
  OR2_X1 U9343 ( .A1(n10277), .A2(n10276), .ZN(n10470) );
  NAND2_X1 U9344 ( .A1(n12359), .A2(n7199), .ZN(n12523) );
  NAND2_X1 U9345 ( .A1(n12460), .A2(n12459), .ZN(n12458) );
  OAI21_X1 U9346 ( .B1(n12511), .B2(n12512), .A(n7167), .ZN(n6928) );
  INV_X1 U9347 ( .A(n7699), .ZN(n7773) );
  NAND2_X1 U9348 ( .A1(n12523), .A2(n12363), .ZN(n12460) );
  AOI21_X2 U9349 ( .B1(n12496), .B2(n12442), .A(n12383), .ZN(n12474) );
  AND4_X1 U9350 ( .A1(n10835), .A2(n12423), .A3(n10832), .A4(n10831), .ZN(
        n10833) );
  NAND2_X1 U9351 ( .A1(n7180), .A2(n7183), .ZN(n12355) );
  NAND2_X1 U9352 ( .A1(n12862), .A2(n12120), .ZN(n12853) );
  NAND2_X1 U9353 ( .A1(n6820), .A2(n9329), .ZN(n7807) );
  AOI21_X2 U9354 ( .B1(n12680), .B2(n12167), .A(n12166), .ZN(n12012) );
  NAND2_X1 U9355 ( .A1(n7302), .A2(n7303), .ZN(n8178) );
  NAND2_X1 U9356 ( .A1(n7720), .A2(n7719), .ZN(n7864) );
  INV_X1 U9357 ( .A(n12008), .ZN(n14787) );
  OAI22_X1 U9358 ( .A1(n11983), .A2(n11982), .B1(P2_DATAO_REG_29__SCAN_IN), 
        .B2(n13846), .ZN(n11987) );
  NAND2_X1 U9359 ( .A1(n10470), .A2(n10469), .ZN(n10471) );
  NAND2_X1 U9360 ( .A1(n10004), .A2(n10005), .ZN(n10092) );
  NAND2_X1 U9361 ( .A1(n12487), .A2(n6754), .ZN(n12438) );
  OAI21_X1 U9362 ( .B1(n6862), .B2(n8282), .A(n6861), .ZN(n12183) );
  NAND2_X1 U9363 ( .A1(n8094), .A2(n7299), .ZN(n7760) );
  AOI21_X1 U9364 ( .B1(n12165), .B2(n12164), .A(n8176), .ZN(n12172) );
  NAND2_X1 U9365 ( .A1(n7194), .A2(n7195), .ZN(n7860) );
  NAND2_X1 U9366 ( .A1(n6826), .A2(n12112), .ZN(n12875) );
  AOI21_X2 U9367 ( .B1(n7099), .B2(n7098), .A(n7095), .ZN(n6824) );
  NAND2_X1 U9368 ( .A1(n8217), .A2(n8216), .ZN(n12873) );
  NAND2_X1 U9369 ( .A1(n7090), .A2(n7086), .ZN(n8222) );
  NAND2_X1 U9370 ( .A1(n8210), .A2(n12071), .ZN(n10957) );
  NAND2_X1 U9371 ( .A1(n8214), .A2(n7092), .ZN(n6826) );
  NAND2_X1 U9372 ( .A1(n8207), .A2(n12058), .ZN(n10375) );
  INV_X1 U9373 ( .A(n8206), .ZN(n15446) );
  NOR2_X2 U9374 ( .A1(n7880), .A2(n7106), .ZN(n8070) );
  INV_X1 U9375 ( .A(n11328), .ZN(n8212) );
  NAND2_X1 U9376 ( .A1(n12682), .A2(n12681), .ZN(n12680) );
  NAND2_X1 U9377 ( .A1(n7877), .A2(n7688), .ZN(n7880) );
  NAND2_X1 U9378 ( .A1(n12012), .A2(n12176), .ZN(n7099) );
  INV_X1 U9379 ( .A(n11278), .ZN(n11314) );
  INV_X1 U9380 ( .A(n11315), .ZN(n6828) );
  NAND2_X1 U9381 ( .A1(n6831), .A2(n11872), .ZN(n12554) );
  OR2_X2 U9382 ( .A1(n11870), .A2(n11871), .ZN(n6831) );
  OR2_X2 U9383 ( .A1(n11877), .A2(n11878), .ZN(n12592) );
  NOR2_X2 U9384 ( .A1(n12628), .A2(n11884), .ZN(n11886) );
  NOR2_X2 U9385 ( .A1(n7860), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n7877) );
  NAND2_X1 U9386 ( .A1(n6739), .A2(n7541), .ZN(n7540) );
  NAND2_X1 U9387 ( .A1(n8348), .A2(n8347), .ZN(n7275) );
  INV_X1 U9388 ( .A(n14717), .ZN(n6853) );
  NAND2_X1 U9389 ( .A1(n14988), .A2(n15251), .ZN(n14985) );
  OAI21_X1 U9390 ( .B1(n12399), .B2(n12520), .A(n6776), .ZN(P3_U3154) );
  NAND2_X2 U9391 ( .A1(n14995), .A2(n8391), .ZN(n14999) );
  NAND2_X1 U9392 ( .A1(n15553), .A2(n15552), .ZN(n15551) );
  INV_X1 U9393 ( .A(n10835), .ZN(n12425) );
  NAND2_X1 U9394 ( .A1(n10891), .A2(n10890), .ZN(n11161) );
  AOI21_X1 U9395 ( .B1(n7682), .B2(n8714), .A(n8713), .ZN(n8716) );
  OAI21_X2 U9396 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(n8354), .A(n14706), .ZN(
        n15559) );
  NAND2_X1 U9397 ( .A1(n8371), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n6852) );
  NAND2_X1 U9398 ( .A1(n7490), .A2(n7488), .ZN(n11942) );
  NAND2_X1 U9399 ( .A1(n8902), .A2(n8901), .ZN(n8923) );
  NAND2_X1 U9400 ( .A1(n7520), .A2(n7518), .ZN(n11242) );
  NAND2_X1 U9401 ( .A1(n7496), .A2(n7497), .ZN(n10590) );
  NOR2_X1 U9402 ( .A1(n11459), .A2(n11460), .ZN(n11913) );
  NOR2_X1 U9403 ( .A1(n9673), .A2(n9672), .ZN(n9693) );
  AOI22_X1 U9404 ( .A1(n9787), .A2(n9786), .B1(n9785), .B2(n9784), .ZN(n9791)
         );
  INV_X1 U9405 ( .A(n14820), .ZN(n6848) );
  INV_X1 U9406 ( .A(n13687), .ZN(n6851) );
  AOI22_X1 U9407 ( .A1(n13622), .A2(n13621), .B1(n13494), .B2(n13785), .ZN(
        n13607) );
  OAI22_X1 U9408 ( .A1(n10609), .A2(n10608), .B1(n10607), .B2(n15347), .ZN(
        n10674) );
  NOR2_X1 U9409 ( .A1(n13689), .A2(n6849), .ZN(n13664) );
  NAND2_X1 U9410 ( .A1(n11242), .A2(n11243), .ZN(n11291) );
  NAND2_X2 U9411 ( .A1(n14852), .A2(n13587), .ZN(n9669) );
  INV_X1 U9412 ( .A(n9251), .ZN(n9254) );
  NAND2_X1 U9413 ( .A1(n6877), .A2(n7637), .ZN(n9251) );
  XNOR2_X2 U9414 ( .A(n14280), .B(n6840), .ZN(n15108) );
  INV_X2 U9415 ( .A(n15118), .ZN(n6840) );
  NAND2_X1 U9416 ( .A1(n14597), .A2(n6895), .ZN(n14674) );
  NAND2_X1 U9417 ( .A1(n10726), .A2(n10725), .ZN(n10728) );
  NAND2_X1 U9418 ( .A1(n13577), .A2(n11845), .ZN(n6841) );
  NAND2_X1 U9419 ( .A1(n11833), .A2(n11832), .ZN(n13736) );
  NAND2_X1 U9420 ( .A1(n6865), .A2(n11008), .ZN(n11004) );
  NAND2_X1 U9421 ( .A1(n10347), .A2(n10348), .ZN(n10190) );
  AOI21_X1 U9422 ( .B1(n13611), .B2(n11843), .A(n6898), .ZN(n13603) );
  XNOR2_X2 U9423 ( .A(n6841), .B(n11846), .ZN(n13765) );
  XNOR2_X2 U9424 ( .A(n13531), .B(n6842), .ZN(n10348) );
  NAND2_X1 U9425 ( .A1(n13734), .A2(n11834), .ZN(n13711) );
  OAI21_X1 U9426 ( .B1(n8764), .B2(n8763), .A(n6753), .ZN(n6873) );
  NOR2_X1 U9427 ( .A1(n9616), .A2(n9615), .ZN(n9668) );
  OAI22_X1 U9428 ( .A1(n11458), .A2(n11457), .B1(n11456), .B2(n11455), .ZN(
        n11459) );
  OAI22_X1 U9429 ( .A1(n6646), .A2(n10072), .B1(n9972), .B2(n9270), .ZN(n9833)
         );
  INV_X1 U9430 ( .A(n10632), .ZN(n9972) );
  NAND2_X1 U9431 ( .A1(n7214), .A2(n6693), .ZN(n10632) );
  OR2_X4 U9432 ( .A1(n6701), .A2(n11811), .ZN(n10529) );
  XNOR2_X2 U9433 ( .A(n9238), .B(n9237), .ZN(n9266) );
  INV_X1 U9434 ( .A(n7414), .ZN(n7413) );
  NAND2_X1 U9435 ( .A1(n6948), .A2(n6660), .ZN(n6947) );
  NAND2_X1 U9436 ( .A1(n7405), .A2(n10235), .ZN(n10286) );
  XNOR2_X2 U9437 ( .A(n8455), .B(n8454), .ZN(n9192) );
  INV_X1 U9438 ( .A(n12179), .ZN(n7097) );
  NAND2_X1 U9439 ( .A1(n7097), .A2(n7096), .ZN(n7095) );
  NAND2_X1 U9440 ( .A1(n7756), .A2(n7301), .ZN(n8094) );
  NAND2_X1 U9441 ( .A1(n7985), .A2(n7741), .ZN(n8000) );
  OAI21_X1 U9442 ( .B1(n8020), .B2(n8019), .A(n8021), .ZN(n9606) );
  NAND2_X1 U9443 ( .A1(n10210), .A2(n10209), .ZN(n10237) );
  NOR2_X1 U9444 ( .A1(n7588), .A2(n7072), .ZN(n7071) );
  NAND2_X1 U9445 ( .A1(n11355), .A2(n7128), .ZN(n11358) );
  XNOR2_X2 U9446 ( .A(n8302), .B(n7284), .ZN(n8345) );
  NAND2_X2 U9447 ( .A1(n8300), .A2(n8301), .ZN(n8302) );
  NOR2_X1 U9448 ( .A1(n14714), .A2(n14715), .ZN(n14713) );
  XNOR2_X1 U9449 ( .A(n6854), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  INV_X1 U9450 ( .A(n14701), .ZN(n6855) );
  NAND2_X1 U9451 ( .A1(n11004), .A2(n10997), .ZN(n11566) );
  NAND2_X1 U9452 ( .A1(n6892), .A2(n11568), .ZN(n14847) );
  NAND2_X1 U9453 ( .A1(n8527), .A2(SI_2_), .ZN(n8508) );
  NAND2_X2 U9454 ( .A1(n8492), .A2(n6712), .ZN(n10200) );
  NAND2_X1 U9455 ( .A1(n14109), .A2(n6755), .ZN(n6859) );
  OAI22_X1 U9456 ( .A1(n6944), .A2(n11759), .B1(n14025), .B2(n9801), .ZN(n7215) );
  NAND2_X1 U9457 ( .A1(n7636), .A2(n7637), .ZN(n9250) );
  OAI211_X1 U9458 ( .C1(n9948), .C2(n14025), .A(n9949), .B(n6689), .ZN(n9950)
         );
  XNOR2_X2 U9459 ( .A(n9219), .B(n9220), .ZN(n11811) );
  OAI21_X1 U9460 ( .B1(n11734), .B2(n6944), .A(n6943), .ZN(n8472) );
  INV_X1 U9461 ( .A(n9646), .ZN(n7218) );
  NAND2_X1 U9462 ( .A1(n10734), .A2(n10733), .ZN(n10757) );
  INV_X1 U9463 ( .A(n11006), .ZN(n6865) );
  NAND2_X1 U9464 ( .A1(n6872), .A2(n14838), .ZN(n14845) );
  NAND2_X1 U9465 ( .A1(n7969), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7972) );
  NAND2_X1 U9466 ( .A1(n8034), .A2(n7747), .ZN(n7749) );
  NAND3_X1 U9467 ( .A1(n6870), .A2(n12174), .A3(n12173), .ZN(n12177) );
  INV_X1 U9468 ( .A(n14847), .ZN(n6872) );
  NAND2_X2 U9469 ( .A1(n6659), .A2(n14835), .ZN(n14834) );
  OAI21_X1 U9470 ( .B1(n12170), .B2(n12169), .A(n12168), .ZN(n6870) );
  NAND2_X1 U9471 ( .A1(n7313), .A2(n7312), .ZN(n8129) );
  OR2_X2 U9472 ( .A1(n12852), .A2(n6644), .ZN(n8047) );
  NAND2_X1 U9473 ( .A1(n13771), .A2(n6748), .ZN(n13578) );
  NAND2_X1 U9474 ( .A1(n6894), .A2(n6893), .ZN(n13734) );
  NAND2_X1 U9475 ( .A1(n7411), .A2(n7412), .ZN(n11006) );
  NAND2_X1 U9476 ( .A1(n8542), .A2(n8541), .ZN(n7673) );
  NAND2_X1 U9477 ( .A1(n7063), .A2(n7064), .ZN(n8652) );
  OAI22_X1 U9478 ( .A1(n7057), .A2(n6778), .B1(n7056), .B2(n7055), .ZN(n8963)
         );
  INV_X1 U9479 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7779) );
  INV_X1 U9480 ( .A(n14832), .ZN(n13587) );
  INV_X1 U9481 ( .A(n8853), .ZN(n7054) );
  NAND2_X1 U9482 ( .A1(n13603), .A2(n13602), .ZN(n13771) );
  XNOR2_X2 U9483 ( .A(n10200), .B(n13532), .ZN(n10198) );
  NOR2_X1 U9484 ( .A1(n8765), .A2(n6873), .ZN(n7068) );
  NAND2_X1 U9485 ( .A1(n8473), .A2(n6945), .ZN(n7581) );
  NAND2_X1 U9486 ( .A1(n10602), .A2(n10601), .ZN(n10672) );
  NAND2_X1 U9487 ( .A1(n13625), .A2(n7408), .ZN(n13611) );
  NAND2_X1 U9488 ( .A1(n10192), .A2(n10191), .ZN(n10234) );
  NAND2_X1 U9489 ( .A1(n10605), .A2(n10604), .ZN(n10726) );
  NAND2_X1 U9490 ( .A1(n10288), .A2(n10287), .ZN(n10600) );
  NAND2_X1 U9491 ( .A1(n7043), .A2(n7042), .ZN(n7041) );
  NAND2_X1 U9492 ( .A1(n7049), .A2(n7048), .ZN(n7047) );
  OAI21_X1 U9493 ( .B1(n9067), .B2(n9066), .A(n7681), .ZN(n9150) );
  NAND2_X1 U9494 ( .A1(n9150), .A2(n7589), .ZN(n7588) );
  OAI211_X2 U9495 ( .C1(n12474), .C2(n12388), .A(n12387), .B(n12386), .ZN(
        n12449) );
  NAND2_X4 U9496 ( .A1(n10529), .A2(n9831), .ZN(n12340) );
  NAND2_X1 U9497 ( .A1(n7173), .A2(n7176), .ZN(n12408) );
  INV_X1 U9498 ( .A(n10833), .ZN(n7189) );
  XNOR2_X1 U9499 ( .A(n6928), .B(n6927), .ZN(n12399) );
  INV_X2 U9500 ( .A(n6645), .ZN(n12333) );
  NOR2_X1 U9501 ( .A1(n9693), .A2(n9692), .ZN(n9787) );
  NOR2_X1 U9502 ( .A1(n9668), .A2(n9667), .ZN(n9673) );
  NAND2_X1 U9503 ( .A1(n6876), .A2(n14042), .ZN(n6878) );
  NAND2_X1 U9504 ( .A1(n14039), .A2(n14040), .ZN(n6876) );
  NAND2_X1 U9505 ( .A1(n14217), .A2(n6884), .ZN(n6883) );
  INV_X1 U9506 ( .A(n14161), .ZN(n7548) );
  NAND2_X1 U9507 ( .A1(n6880), .A2(n6698), .ZN(n7538) );
  NAND2_X1 U9508 ( .A1(n14105), .A2(n14106), .ZN(n14104) );
  NAND2_X1 U9509 ( .A1(n6878), .A2(n14043), .ZN(n14052) );
  NAND2_X1 U9510 ( .A1(n14184), .A2(n7126), .ZN(n6879) );
  NAND3_X1 U9511 ( .A1(n14117), .A2(n14116), .A3(n6881), .ZN(n6880) );
  XNOR2_X1 U9512 ( .A(n8509), .B(n8524), .ZN(n9344) );
  NAND2_X1 U9513 ( .A1(n14100), .A2(n6887), .ZN(n14105) );
  NAND2_X1 U9514 ( .A1(n14061), .A2(n14060), .ZN(n14065) );
  NAND2_X1 U9515 ( .A1(n7552), .A2(n7551), .ZN(n14094) );
  INV_X1 U9516 ( .A(n14050), .ZN(n7555) );
  OAI21_X1 U9517 ( .B1(n7121), .B2(n7119), .A(n7534), .ZN(n14201) );
  OAI22_X1 U9518 ( .A1(n14252), .A2(n6883), .B1(n14251), .B2(n14250), .ZN(
        n14253) );
  NAND2_X1 U9519 ( .A1(n6889), .A2(n6888), .ZN(n6887) );
  INV_X1 U9520 ( .A(n14101), .ZN(n6889) );
  AOI21_X1 U9521 ( .B1(n14189), .B2(n14188), .A(n7120), .ZN(n7119) );
  OAI21_X1 U9522 ( .B1(n14157), .B2(n14159), .A(n14160), .ZN(n7547) );
  NAND2_X1 U9523 ( .A1(n10190), .A2(n10189), .ZN(n10217) );
  NAND2_X1 U9524 ( .A1(n6891), .A2(n11839), .ZN(n13679) );
  INV_X1 U9525 ( .A(n13736), .ZN(n6894) );
  NAND2_X2 U9526 ( .A1(n8458), .A2(n8459), .ZN(n9469) );
  NAND2_X1 U9527 ( .A1(n13696), .A2(n11838), .ZN(n6891) );
  NAND2_X1 U9528 ( .A1(n11566), .A2(n11565), .ZN(n6892) );
  NAND2_X1 U9529 ( .A1(n13769), .A2(n6899), .ZN(n13829) );
  OAI21_X1 U9530 ( .B1(n13770), .B2(n15350), .A(n13768), .ZN(n6900) );
  NOR2_X2 U9531 ( .A1(n12592), .A2(n12593), .ZN(n12591) );
  NAND2_X1 U9532 ( .A1(n11907), .A2(n12652), .ZN(n6996) );
  OAI22_X1 U9533 ( .A1(n10870), .A2(n10869), .B1(n14087), .B2(n14274), .ZN(
        n10872) );
  INV_X1 U9534 ( .A(n8525), .ZN(n6948) );
  INV_X1 U9535 ( .A(n14468), .ZN(n6922) );
  NAND2_X1 U9536 ( .A1(n6959), .A2(n6957), .ZN(P1_U3557) );
  NAND2_X1 U9537 ( .A1(n7622), .A2(n7620), .ZN(n11087) );
  NAND4_X2 U9538 ( .A1(n8485), .A2(n8484), .A3(n8483), .A4(n8482), .ZN(n13532)
         );
  NAND2_X1 U9539 ( .A1(n7262), .A2(n7260), .ZN(n13622) );
  NAND2_X1 U9540 ( .A1(n7235), .A2(n7234), .ZN(n13582) );
  NAND2_X1 U9541 ( .A1(n12677), .A2(n8177), .ZN(n12661) );
  NAND2_X1 U9542 ( .A1(n12771), .A2(n8105), .ZN(n12753) );
  NAND2_X1 U9543 ( .A1(n7309), .A2(n7734), .ZN(n7941) );
  NAND2_X1 U9544 ( .A1(n7726), .A2(n7725), .ZN(n7896) );
  NAND2_X1 U9545 ( .A1(n7466), .A2(n7464), .ZN(n7463) );
  XNOR2_X1 U9546 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n7787) );
  XNOR2_X2 U9547 ( .A(n9290), .B(n9289), .ZN(n11619) );
  OAI21_X1 U9548 ( .B1(n12961), .B2(n15544), .A(n6904), .ZN(P3_U3487) );
  OAI21_X1 U9549 ( .B1(n12961), .B2(n7083), .A(n6906), .ZN(P3_U3455) );
  NAND2_X1 U9550 ( .A1(n14983), .A2(n14982), .ZN(n14981) );
  NOR2_X1 U9551 ( .A1(n14719), .A2(n14718), .ZN(n14717) );
  NAND2_X1 U9552 ( .A1(n6909), .A2(n8630), .ZN(n8634) );
  NAND2_X1 U9553 ( .A1(n7371), .A2(n7369), .ZN(n14415) );
  AOI22_X1 U9554 ( .A1(n14411), .A2(n14410), .B1(n14614), .B2(n14424), .ZN(
        n14399) );
  AOI21_X1 U9555 ( .B1(n7380), .B2(n9952), .A(n6762), .ZN(n10325) );
  INV_X1 U9556 ( .A(n8472), .ZN(n6946) );
  INV_X1 U9557 ( .A(n14374), .ZN(n6963) );
  NAND2_X1 U9558 ( .A1(n7921), .A2(n7732), .ZN(n7309) );
  NAND2_X1 U9559 ( .A1(n7876), .A2(n7723), .ZN(n7726) );
  NAND2_X1 U9560 ( .A1(n7292), .A2(n7295), .ZN(n8021) );
  NAND2_X1 U9561 ( .A1(n7788), .A2(n6914), .ZN(n9998) );
  NAND2_X1 U9562 ( .A1(n6921), .A2(n6920), .ZN(n6919) );
  NAND2_X1 U9563 ( .A1(n12147), .A2(n6752), .ZN(n6921) );
  NAND2_X1 U9564 ( .A1(n11358), .A2(n11359), .ZN(n11497) );
  NAND2_X1 U9565 ( .A1(n13940), .A2(n6744), .ZN(n14905) );
  NAND2_X1 U9566 ( .A1(n13971), .A2(n6923), .ZN(n11050) );
  NAND2_X1 U9567 ( .A1(n13973), .A2(n13972), .ZN(n13971) );
  INV_X1 U9568 ( .A(n11204), .ZN(n6926) );
  XNOR2_X1 U9569 ( .A(n8367), .B(P2_ADDR_REG_7__SCAN_IN), .ZN(n15557) );
  NAND2_X1 U9570 ( .A1(n8346), .A2(n14310), .ZN(n8300) );
  AOI21_X2 U9571 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(n8372), .A(n14726), .ZN(
        n14983) );
  NAND2_X1 U9572 ( .A1(n7606), .A2(n7605), .ZN(n7604) );
  INV_X4 U9573 ( .A(n9800), .ZN(n8991) );
  INV_X1 U9574 ( .A(n11811), .ZN(n9588) );
  INV_X1 U9575 ( .A(n11502), .ZN(n11505) );
  NAND2_X2 U9576 ( .A1(n12458), .A2(n12365), .ZN(n12468) );
  AOI21_X2 U9577 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n8393), .A(n14701), .ZN(
        n8402) );
  NAND2_X1 U9578 ( .A1(n8450), .A2(n7409), .ZN(n8456) );
  OAI21_X2 U9579 ( .B1(n9644), .B2(n6636), .A(n9640), .ZN(n10186) );
  INV_X1 U9580 ( .A(n13942), .ZN(n6936) );
  NAND2_X1 U9581 ( .A1(n7130), .A2(n7129), .ZN(n13983) );
  INV_X1 U9582 ( .A(n7215), .ZN(n7214) );
  NAND4_X4 U9583 ( .A1(n7151), .A2(n7612), .A3(n9210), .A4(n6668), .ZN(n10118)
         );
  NAND2_X1 U9584 ( .A1(n8604), .A2(n8607), .ZN(n6937) );
  NAND2_X1 U9585 ( .A1(n11734), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6943) );
  OAI211_X1 U9586 ( .C1(n11734), .C2(P2_DATAO_REG_0__SCAN_IN), .A(n6940), .B(
        SI_0_), .ZN(n8490) );
  INV_X1 U9587 ( .A(n8527), .ZN(n6950) );
  NAND3_X1 U9588 ( .A1(n7582), .A2(n6660), .A3(n6950), .ZN(n6949) );
  NAND3_X1 U9589 ( .A1(n6953), .A2(n6952), .A3(n8528), .ZN(n8552) );
  INV_X1 U9590 ( .A(n14469), .ZN(n6956) );
  OR2_X2 U9591 ( .A1(n6955), .A2(n6954), .ZN(n14452) );
  NAND2_X2 U9592 ( .A1(n6964), .A2(n11725), .ZN(n14644) );
  NAND2_X1 U9593 ( .A1(n8694), .A2(n6969), .ZN(n6966) );
  NAND2_X1 U9594 ( .A1(n6967), .A2(n6966), .ZN(n8748) );
  INV_X2 U9595 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7197) );
  AND2_X1 U9596 ( .A1(n6979), .A2(n11896), .ZN(n11897) );
  NAND2_X1 U9597 ( .A1(n10494), .A2(n7440), .ZN(n6987) );
  NAND2_X1 U9598 ( .A1(n6987), .A2(n6986), .ZN(n10916) );
  NAND3_X1 U9599 ( .A1(n6989), .A2(n6666), .A3(n10492), .ZN(n6986) );
  NAND2_X1 U9600 ( .A1(n6989), .A2(n10492), .ZN(n10447) );
  INV_X1 U9601 ( .A(n10446), .ZN(n6991) );
  NAND3_X1 U9602 ( .A1(n6996), .A2(n6993), .A3(n6992), .ZN(P3_U3201) );
  MUX2_X1 U9603 ( .A(n10629), .B(P1_REG2_REG_1__SCAN_IN), .S(n9802), .Z(n14291) );
  INV_X1 U9604 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7026) );
  NAND3_X1 U9605 ( .A1(n7026), .A2(n7025), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n7573) );
  OAI21_X1 U9606 ( .B1(n8768), .B2(n7576), .A(n7027), .ZN(n7029) );
  NOR2_X1 U9607 ( .A1(n7032), .A2(n6777), .ZN(n7033) );
  INV_X1 U9608 ( .A(n8496), .ZN(n7042) );
  INV_X1 U9609 ( .A(n7047), .ZN(n7043) );
  NAND2_X1 U9610 ( .A1(n7046), .A2(n7045), .ZN(n7044) );
  INV_X1 U9611 ( .A(n8495), .ZN(n7045) );
  NAND2_X1 U9612 ( .A1(n7047), .A2(n8496), .ZN(n7046) );
  NAND2_X1 U9613 ( .A1(n8479), .A2(n8480), .ZN(n7048) );
  OAI211_X1 U9614 ( .C1(n8562), .C2(n7053), .A(n7050), .B(n7660), .ZN(n7657)
         );
  NAND2_X1 U9615 ( .A1(n7052), .A2(n7051), .ZN(n7050) );
  NAND2_X1 U9616 ( .A1(n7053), .A2(n8562), .ZN(n7052) );
  NAND2_X1 U9617 ( .A1(n7671), .A2(n7670), .ZN(n7053) );
  NAND2_X1 U9618 ( .A1(n7058), .A2(n7059), .ZN(n7650) );
  INV_X1 U9619 ( .A(n6743), .ZN(n7062) );
  NAND2_X1 U9620 ( .A1(n8603), .A2(n6655), .ZN(n7063) );
  INV_X1 U9621 ( .A(n8602), .ZN(n7067) );
  NAND2_X1 U9622 ( .A1(n10957), .A2(n6682), .ZN(n7076) );
  NAND2_X1 U9623 ( .A1(n12838), .A2(n8221), .ZN(n7090) );
  CLKBUF_X1 U9624 ( .A(n7090), .Z(n7085) );
  INV_X1 U9625 ( .A(n12875), .ZN(n8217) );
  NAND2_X1 U9626 ( .A1(n12739), .A2(n7094), .ZN(n12721) );
  NAND2_X4 U9627 ( .A1(n7110), .A2(n7109), .ZN(n11734) );
  NAND2_X1 U9628 ( .A1(n13922), .A2(n7132), .ZN(n7130) );
  NAND2_X1 U9629 ( .A1(n14930), .A2(n6703), .ZN(n7145) );
  AND2_X1 U9630 ( .A1(n9210), .A2(n9208), .ZN(n7153) );
  INV_X1 U9631 ( .A(n9214), .ZN(n9873) );
  OAI21_X2 U9632 ( .B1(n7154), .B2(n9992), .A(n9994), .ZN(n10089) );
  NAND2_X1 U9633 ( .A1(n12511), .A2(n7156), .ZN(n7155) );
  OAI211_X1 U9634 ( .C1(n12511), .C2(n7157), .A(n7155), .B(n7172), .ZN(
        P3_U3160) );
  NAND2_X1 U9635 ( .A1(n12468), .A2(n7174), .ZN(n7173) );
  NAND2_X1 U9636 ( .A1(n11522), .A2(n7181), .ZN(n7180) );
  NAND2_X1 U9637 ( .A1(n12438), .A2(n12378), .ZN(n12382) );
  OR2_X2 U9638 ( .A1(n10471), .A2(n7189), .ZN(n7191) );
  AND3_X2 U9639 ( .A1(n7198), .A2(n7197), .A3(n7687), .ZN(n7194) );
  NOR2_X2 U9640 ( .A1(n10340), .A2(n14062), .ZN(n10575) );
  NOR2_X1 U9641 ( .A1(n15119), .A2(n15118), .ZN(n15122) );
  NOR2_X2 U9642 ( .A1(n14489), .A2(n14639), .ZN(n14480) );
  NOR2_X2 U9643 ( .A1(n14576), .A2(n7207), .ZN(n14535) );
  NOR2_X1 U9644 ( .A1(n14406), .A2(n7213), .ZN(n14379) );
  INV_X1 U9645 ( .A(n14406), .ZN(n7210) );
  NAND3_X1 U9646 ( .A1(n7210), .A2(n7209), .A3(n14366), .ZN(n14364) );
  NAND3_X1 U9647 ( .A1(n7217), .A2(n8403), .A3(n7649), .ZN(n8505) );
  AND3_X2 U9648 ( .A1(n7217), .A2(n8403), .A3(n7216), .ZN(n8555) );
  NOR2_X2 U9649 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n7217) );
  XNOR2_X1 U9650 ( .A(n9645), .B(n7218), .ZN(n9644) );
  NAND2_X1 U9651 ( .A1(n7219), .A2(n10987), .ZN(n11009) );
  NAND2_X1 U9652 ( .A1(n10759), .A2(n7220), .ZN(n7219) );
  NOR2_X1 U9653 ( .A1(n10988), .A2(n7221), .ZN(n7220) );
  XNOR2_X1 U9654 ( .A(n7222), .B(n10988), .ZN(n10760) );
  NAND2_X1 U9655 ( .A1(n8453), .A2(n6759), .ZN(n7223) );
  NAND2_X1 U9656 ( .A1(n7225), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9185) );
  AND2_X1 U9657 ( .A1(n9191), .A2(n7225), .ZN(n9445) );
  NAND2_X1 U9658 ( .A1(n13593), .A2(n13592), .ZN(n7235) );
  NAND2_X1 U9659 ( .A1(n7235), .A2(n7227), .ZN(n7226) );
  OAI211_X1 U9660 ( .C1(n7235), .C2(n7232), .A(n7228), .B(n7226), .ZN(n11831)
         );
  NAND2_X1 U9661 ( .A1(n10237), .A2(n7238), .ZN(n7239) );
  NAND2_X1 U9662 ( .A1(n7239), .A2(n7240), .ZN(n10609) );
  NAND2_X1 U9663 ( .A1(n13742), .A2(n7244), .ZN(n7243) );
  NAND2_X1 U9664 ( .A1(n7243), .A2(n7246), .ZN(n13712) );
  NAND2_X1 U9665 ( .A1(n11011), .A2(n7253), .ZN(n7252) );
  NAND2_X1 U9666 ( .A1(n7252), .A2(n7255), .ZN(n14820) );
  NAND2_X1 U9667 ( .A1(n13662), .A2(n7263), .ZN(n7262) );
  INV_X1 U9668 ( .A(n13800), .ZN(n7269) );
  NOR2_X2 U9669 ( .A1(n8376), .A2(n8375), .ZN(n14986) );
  AND2_X2 U9670 ( .A1(n7280), .A2(n7279), .ZN(n14701) );
  NAND2_X1 U9671 ( .A1(n8049), .A2(n7289), .ZN(n7288) );
  NAND2_X1 U9672 ( .A1(n7985), .A2(n7293), .ZN(n7292) );
  INV_X1 U9673 ( .A(n7755), .ZN(n7298) );
  NOR2_X1 U9674 ( .A1(n7298), .A2(n8091), .ZN(n7301) );
  NAND2_X1 U9675 ( .A1(n8151), .A2(n7304), .ZN(n7302) );
  OAI21_X1 U9676 ( .B1(n8151), .B2(n7767), .A(n7768), .ZN(n8164) );
  NAND2_X1 U9677 ( .A1(n13024), .A2(n11998), .ZN(n7308) );
  NAND2_X1 U9678 ( .A1(n7308), .A2(n7306), .ZN(n12010) );
  NOR2_X2 U9679 ( .A1(n13717), .A2(n13813), .ZN(n7319) );
  INV_X1 U9680 ( .A(n14850), .ZN(n7324) );
  NAND2_X1 U9681 ( .A1(n7324), .A2(n7325), .ZN(n13729) );
  OAI22_X1 U9682 ( .A1(n9109), .A2(n9801), .B1(n8533), .B2(n15203), .ZN(n7331)
         );
  INV_X1 U9683 ( .A(n9645), .ZN(n9568) );
  NAND2_X1 U9684 ( .A1(n12638), .A2(n7343), .ZN(n7342) );
  NOR2_X1 U9685 ( .A1(n14091), .A2(n14226), .ZN(n7365) );
  NAND2_X1 U9686 ( .A1(n10325), .A2(n14224), .ZN(n10550) );
  NAND2_X1 U9687 ( .A1(n7385), .A2(n7383), .ZN(n11418) );
  NOR2_X1 U9688 ( .A1(n7386), .A2(n7384), .ZN(n7383) );
  OAI21_X1 U9689 ( .B1(n14556), .B2(n7393), .A(n7389), .ZN(n11710) );
  XNOR2_X1 U9690 ( .A(n6932), .B(n9972), .ZN(n14222) );
  NAND2_X1 U9691 ( .A1(n10286), .A2(n10285), .ZN(n10288) );
  NAND2_X1 U9692 ( .A1(n10234), .A2(n10233), .ZN(n7405) );
  NOR2_X2 U9693 ( .A1(n8433), .A2(n7410), .ZN(n7533) );
  NAND4_X1 U9694 ( .A1(n8432), .A2(n8431), .A3(n8430), .A4(n8429), .ZN(n7410)
         );
  NAND4_X1 U9695 ( .A1(n8413), .A2(n8412), .A3(n8416), .A4(n8409), .ZN(n8433)
         );
  NAND2_X1 U9696 ( .A1(n10728), .A2(n7413), .ZN(n7411) );
  NAND3_X1 U9697 ( .A1(n7419), .A2(n7420), .A3(n11842), .ZN(n7418) );
  INV_X1 U9698 ( .A(n11840), .ZN(n7424) );
  XNOR2_X2 U9699 ( .A(n7430), .B(n7429), .ZN(n10317) );
  NAND3_X1 U9700 ( .A1(n7444), .A2(n7443), .A3(n6779), .ZN(n10446) );
  NOR2_X2 U9701 ( .A1(n8047), .A2(n7467), .ZN(n7466) );
  NAND2_X1 U9702 ( .A1(n8162), .A2(n6750), .ZN(n12677) );
  NAND2_X1 U9703 ( .A1(n11214), .A2(n7472), .ZN(n11144) );
  NAND2_X2 U9704 ( .A1(n11215), .A2(n12021), .ZN(n11214) );
  NAND2_X1 U9705 ( .A1(n12782), .A2(n7477), .ZN(n12771) );
  NAND2_X1 U9706 ( .A1(n10145), .A2(n7429), .ZN(n7817) );
  NAND2_X1 U9707 ( .A1(n7478), .A2(n10145), .ZN(n7831) );
  NAND2_X1 U9708 ( .A1(n9922), .A2(n7498), .ZN(n7496) );
  NAND2_X1 U9709 ( .A1(n13420), .A2(n7513), .ZN(n7505) );
  OAI21_X1 U9710 ( .B1(n13420), .B2(n7509), .A(n7506), .ZN(n11971) );
  INV_X1 U9711 ( .A(n13419), .ZN(n7517) );
  NAND2_X1 U9712 ( .A1(n11161), .A2(n7521), .ZN(n7520) );
  NAND2_X2 U9713 ( .A1(n8533), .A2(n6832), .ZN(n9109) );
  NAND2_X1 U9714 ( .A1(n9568), .A2(n9646), .ZN(n9640) );
  OAI22_X1 U9715 ( .A1(n13461), .A2(n9568), .B1(n9617), .B2(n13476), .ZN(n9618) );
  NAND3_X1 U9716 ( .A1(n10388), .A2(n10387), .A3(n7529), .ZN(n10389) );
  OR2_X1 U9717 ( .A1(n15282), .A2(n9568), .ZN(n7529) );
  NAND2_X1 U9718 ( .A1(n13449), .A2(n7532), .ZN(n7530) );
  NAND4_X1 U9719 ( .A1(n8434), .A2(n8555), .A3(n7533), .A4(n8451), .ZN(n9187)
         );
  INV_X1 U9720 ( .A(n8433), .ZN(n8414) );
  INV_X1 U9721 ( .A(n14201), .ZN(n14203) );
  INV_X1 U9722 ( .A(n14146), .ZN(n7541) );
  NAND2_X1 U9723 ( .A1(n7544), .A2(n7538), .ZN(n14153) );
  INV_X1 U9724 ( .A(n14541), .ZN(n7545) );
  AOI21_X1 U9725 ( .B1(n7549), .B2(n14009), .A(n14038), .ZN(n14030) );
  NAND2_X1 U9726 ( .A1(n14009), .A2(n14008), .ZN(n14194) );
  NAND2_X1 U9727 ( .A1(n14194), .A2(n14010), .ZN(n7550) );
  NAND3_X1 U9728 ( .A1(n14070), .A2(n14069), .A3(n6763), .ZN(n7552) );
  INV_X1 U9729 ( .A(n14072), .ZN(n7553) );
  NAND2_X1 U9730 ( .A1(n7561), .A2(n7562), .ZN(n14182) );
  NAND3_X1 U9731 ( .A1(n7778), .A2(P3_ADDR_REG_19__SCAN_IN), .A3(n7572), .ZN(
        n7571) );
  NAND2_X1 U9732 ( .A1(n7580), .A2(n8769), .ZN(n8788) );
  NAND2_X1 U9733 ( .A1(n9015), .A2(n7586), .ZN(n7583) );
  NAND2_X1 U9734 ( .A1(n6654), .A2(n11376), .ZN(n7591) );
  INV_X1 U9735 ( .A(n11376), .ZN(n7596) );
  NOR2_X1 U9736 ( .A1(n11376), .A2(n7608), .ZN(n11486) );
  INV_X1 U9737 ( .A(n7604), .ZN(n7603) );
  INV_X1 U9738 ( .A(n11381), .ZN(n7607) );
  NAND2_X1 U9739 ( .A1(n10872), .A2(n7623), .ZN(n7622) );
  NAND2_X1 U9740 ( .A1(n14527), .A2(n6656), .ZN(n7626) );
  NAND2_X1 U9741 ( .A1(n7626), .A2(n7627), .ZN(n14496) );
  INV_X1 U9742 ( .A(n7628), .ZN(n14526) );
  INV_X1 U9743 ( .A(n10118), .ZN(n7636) );
  INV_X1 U9744 ( .A(n7635), .ZN(n7638) );
  NOR2_X2 U9745 ( .A1(n9227), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n7635) );
  NAND2_X1 U9746 ( .A1(n8439), .A2(n8438), .ZN(n8459) );
  NAND3_X1 U9747 ( .A1(n7649), .A2(n8486), .A3(n7648), .ZN(n8503) );
  NOR2_X1 U9748 ( .A1(n7682), .A2(n8714), .ZN(n8715) );
  NOR2_X1 U9749 ( .A1(n8982), .A2(n8981), .ZN(n9066) );
  NAND2_X1 U9750 ( .A1(n7657), .A2(n7658), .ZN(n8603) );
  NAND2_X1 U9751 ( .A1(n7662), .A2(n7663), .ZN(n8898) );
  NAND2_X1 U9752 ( .A1(n8878), .A2(n7665), .ZN(n7662) );
  NAND2_X1 U9753 ( .A1(n8516), .A2(n8515), .ZN(n7672) );
  NAND2_X1 U9754 ( .A1(n8266), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8267) );
  XNOR2_X1 U9755 ( .A(n10151), .B(n10150), .ZN(n10433) );
  AND2_X2 U9756 ( .A1(n7703), .A2(n7705), .ZN(n8186) );
  NAND2_X2 U9757 ( .A1(n8510), .A2(n8511), .ZN(n10359) );
  NOR2_X2 U9758 ( .A1(n10741), .A2(n15369), .ZN(n10767) );
  AOI22_X2 U9759 ( .A1(n12449), .A2(n12450), .B1(n12513), .B2(n12389), .ZN(
        n12511) );
  NAND2_X1 U9760 ( .A1(n11330), .A2(n12093), .ZN(n11329) );
  NAND2_X1 U9761 ( .A1(n11144), .A2(n7913), .ZN(n11330) );
  NAND2_X1 U9762 ( .A1(n12051), .A2(n15460), .ZN(n10001) );
  NAND2_X1 U9763 ( .A1(n7701), .A2(n13022), .ZN(n13027) );
  NAND2_X1 U9764 ( .A1(n7699), .A2(n7697), .ZN(n13022) );
  INV_X1 U9765 ( .A(n9187), .ZN(n8453) );
  NAND2_X1 U9767 ( .A1(n9998), .A2(n15451), .ZN(n12050) );
  INV_X1 U9768 ( .A(n15451), .ZN(n9997) );
  INV_X1 U9769 ( .A(n7877), .ZN(n7878) );
  INV_X2 U9770 ( .A(n14699), .ZN(n14007) );
  NAND2_X1 U9771 ( .A1(n9271), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n9267) );
  MUX2_X2 U9772 ( .A(P1_IR_REG_0__SCAN_IN), .B(n14700), .S(n11737), .Z(n10667)
         );
  CLKBUF_X3 U9773 ( .A(n9942), .Z(n11751) );
  NAND2_X1 U9774 ( .A1(n14167), .A2(n14166), .ZN(n14168) );
  OR2_X1 U9775 ( .A1(n11803), .A2(n14579), .ZN(n14519) );
  NAND2_X1 U9776 ( .A1(n9821), .A2(n14579), .ZN(n9929) );
  NAND2_X1 U9777 ( .A1(n14852), .A2(n6843), .ZN(n9579) );
  NAND2_X1 U9778 ( .A1(n9254), .A2(n9253), .ZN(n9256) );
  NAND2_X1 U9779 ( .A1(n14543), .A2(n14147), .ZN(n14527) );
  AND2_X1 U9780 ( .A1(n8476), .A2(n8475), .ZN(n8479) );
  INV_X1 U9781 ( .A(n11621), .ZN(n9258) );
  NAND2_X1 U9782 ( .A1(n9259), .A2(n11621), .ZN(n11800) );
  INV_X1 U9783 ( .A(n9240), .ZN(n9244) );
  AOI211_X1 U9784 ( .C1(n14210), .C2(n14361), .A(n14205), .B(n14209), .ZN(
        n14252) );
  INV_X1 U9785 ( .A(n8442), .ZN(n8441) );
  OR2_X1 U9786 ( .A1(n8056), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n7674) );
  INV_X2 U9787 ( .A(n15526), .ZN(n15528) );
  AND2_X1 U9788 ( .A1(n8290), .A2(n8289), .ZN(n15526) );
  OR2_X1 U9789 ( .A1(n14951), .A2(n14266), .ZN(n7676) );
  NOR2_X1 U9790 ( .A1(n12290), .A2(n13946), .ZN(n7677) );
  INV_X1 U9791 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9209) );
  NOR4_X1 U9792 ( .A1(n9199), .A2(n6637), .A3(n6843), .A4(n11137), .ZN(n7679)
         );
  INV_X1 U9793 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n8719) );
  INV_X1 U9794 ( .A(n13854), .ZN(n11136) );
  CLKBUF_X2 U9795 ( .A(P1_U4016), .Z(n14282) );
  INV_X1 U9796 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8774) );
  INV_X1 U9797 ( .A(SI_17_), .ZN(n9687) );
  CLKBUF_X3 U9798 ( .A(n8574), .Z(n9102) );
  AND2_X1 U9799 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7680) );
  AND2_X1 U9800 ( .A1(n9087), .A2(n9065), .ZN(n7681) );
  AND2_X1 U9801 ( .A1(n7968), .A2(n7967), .ZN(n7683) );
  NOR2_X1 U9802 ( .A1(n12303), .A2(n13869), .ZN(n7684) );
  OR2_X1 U9803 ( .A1(n10184), .A2(n13587), .ZN(n7685) );
  NAND2_X1 U9804 ( .A1(n11625), .A2(n10284), .ZN(n15288) );
  AND2_X2 U9805 ( .A1(n10194), .A2(n14827), .ZN(n15292) );
  NAND2_X1 U9806 ( .A1(n10035), .A2(n10034), .ZN(n15192) );
  INV_X2 U9807 ( .A(n15192), .ZN(n15194) );
  OR2_X1 U9808 ( .A1(n15281), .A2(n9121), .ZN(n8493) );
  INV_X1 U9809 ( .A(n8514), .ZN(n8515) );
  MUX2_X1 U9810 ( .A(n14046), .B(n14045), .S(n14280), .Z(n14048) );
  NAND2_X1 U9811 ( .A1(n14068), .A2(n14067), .ZN(n14069) );
  INV_X1 U9812 ( .A(n8899), .ZN(n8900) );
  INV_X1 U9813 ( .A(n8946), .ZN(n8947) );
  INV_X1 U9814 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n7691) );
  INV_X1 U9815 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10148) );
  AND2_X1 U9816 ( .A1(n8436), .A2(n8435), .ZN(n8437) );
  NOR2_X1 U9817 ( .A1(n6641), .A2(n10148), .ZN(n10149) );
  INV_X1 U9818 ( .A(n12681), .ZN(n8176) );
  AND2_X1 U9819 ( .A1(n9018), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n9002) );
  NOR2_X1 U9820 ( .A1(n14075), .A2(n11084), .ZN(n11085) );
  INV_X1 U9821 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10162) );
  AND2_X1 U9822 ( .A1(n11899), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n11900) );
  INV_X1 U9823 ( .A(n8219), .ZN(n8220) );
  AND2_X1 U9824 ( .A1(n9552), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n7735) );
  NOR2_X1 U9825 ( .A1(n8661), .A2(n8660), .ZN(n8678) );
  INV_X1 U9826 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n11185) );
  NOR2_X1 U9827 ( .A1(n8775), .A2(n8774), .ZN(n8796) );
  OR2_X1 U9828 ( .A1(n14565), .A2(n14913), .ZN(n11782) );
  INV_X1 U9829 ( .A(n14557), .ZN(n11781) );
  INV_X1 U9830 ( .A(n8854), .ZN(n8857) );
  OR2_X1 U9831 ( .A1(n7991), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8010) );
  NOR2_X1 U9832 ( .A1(n10433), .A2(n10434), .ZN(n10432) );
  INV_X1 U9833 ( .A(n12877), .ZN(n8216) );
  INV_X1 U9834 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n7886) );
  NAND2_X1 U9835 ( .A1(n8212), .A2(n12101), .ZN(n8213) );
  INV_X1 U9836 ( .A(n8280), .ZN(n8287) );
  NAND2_X1 U9837 ( .A1(n8140), .A2(n7764), .ZN(n7766) );
  AND2_X1 U9838 ( .A1(n7743), .A2(n7742), .ZN(n7999) );
  INV_X1 U9839 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8640) );
  AND2_X1 U9840 ( .A1(n8678), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8703) );
  OR2_X1 U9841 ( .A1(n8911), .A2(n8910), .ZN(n8932) );
  NAND2_X1 U9842 ( .A1(n8884), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8911) );
  INV_X1 U9843 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8998) );
  INV_X1 U9844 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8454) );
  AND3_X1 U9845 ( .A1(n8416), .A2(n8415), .A3(P2_IR_REG_19__SCAN_IN), .ZN(
        n8419) );
  OR2_X1 U9846 ( .A1(n12226), .A2(n12225), .ZN(n12227) );
  AND2_X1 U9847 ( .A1(n14928), .A2(n14929), .ZN(n12223) );
  INV_X2 U9848 ( .A(n12242), .ZN(n12341) );
  INV_X1 U9849 ( .A(n11739), .ZN(n11727) );
  INV_X1 U9850 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n11385) );
  OR2_X1 U9851 ( .A1(n9816), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9815) );
  INV_X1 U9852 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9253) );
  INV_X1 U9853 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n8314) );
  INV_X1 U9854 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n11280) );
  AND2_X1 U9855 ( .A1(n8120), .A2(n12400), .ZN(n8132) );
  INV_X1 U9856 ( .A(n12772), .ZN(n12442) );
  OR2_X1 U9857 ( .A1(n8143), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8154) );
  NAND2_X1 U9858 ( .A1(n8041), .A2(n8040), .ZN(n8056) );
  NAND2_X1 U9859 ( .A1(n7900), .A2(n13326), .ZN(n7914) );
  NOR2_X1 U9860 ( .A1(n8109), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8120) );
  NOR2_X1 U9861 ( .A1(n8154), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8167) );
  AND4_X1 U9862 ( .A1(n8061), .A2(n8060), .A3(n8059), .A4(n8058), .ZN(n12800)
         );
  AND2_X1 U9863 ( .A1(n8262), .A2(n8261), .ZN(n8264) );
  OR2_X1 U9864 ( .A1(n10124), .A2(n10123), .ZN(n10175) );
  INV_X1 U9865 ( .A(n12152), .ZN(n12740) );
  INV_X1 U9866 ( .A(n12146), .ZN(n12761) );
  INV_X1 U9867 ( .A(n12833), .ZN(n12861) );
  NOR2_X1 U9868 ( .A1(n7869), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7887) );
  AND2_X1 U9869 ( .A1(n10109), .A2(n12014), .ZN(n15444) );
  INV_X1 U9870 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n8291) );
  INV_X1 U9871 ( .A(n12848), .ZN(n12879) );
  INV_X1 U9872 ( .A(n12540), .ZN(n14778) );
  AND2_X1 U9873 ( .A1(n15470), .A2(n15522), .ZN(n14790) );
  INV_X1 U9874 ( .A(n15466), .ZN(n15456) );
  NAND2_X1 U9875 ( .A1(n10014), .A2(n12171), .ZN(n15448) );
  NAND2_X1 U9876 ( .A1(n7972), .A2(n7739), .ZN(n7983) );
  INV_X1 U9877 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9153) );
  OR2_X1 U9878 ( .A1(n8727), .A2(n9712), .ZN(n8754) );
  NAND2_X1 U9879 ( .A1(n9694), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13498) );
  AND4_X1 U9880 ( .A1(n8733), .A2(n8732), .A3(n8731), .A4(n8730), .ZN(n11577)
         );
  OR2_X1 U9881 ( .A1(n9517), .A2(n9516), .ZN(n15236) );
  INV_X1 U9882 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9712) );
  INV_X1 U9883 ( .A(n11571), .ZN(n13751) );
  INV_X1 U9884 ( .A(n14852), .ZN(n13728) );
  INV_X1 U9885 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8440) );
  OR2_X1 U9886 ( .A1(n6648), .A2(n11911), .ZN(n11643) );
  INV_X1 U9887 ( .A(n11503), .ZN(n11504) );
  AND2_X1 U9888 ( .A1(n12348), .A2(n12347), .ZN(n14599) );
  INV_X1 U9889 ( .A(n14424), .ZN(n13910) );
  NOR2_X1 U9890 ( .A1(n13275), .A2(n11714), .ZN(n11726) );
  INV_X1 U9891 ( .A(n11750), .ZN(n11738) );
  OR2_X1 U9892 ( .A1(n11690), .A2(n11689), .ZN(n11703) );
  AND3_X1 U9893 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n10331) );
  NAND2_X1 U9894 ( .A1(n14699), .A2(n9977), .ZN(n14022) );
  AND2_X1 U9895 ( .A1(n11773), .A2(n11645), .ZN(n14392) );
  INV_X1 U9896 ( .A(n9385), .ZN(n9301) );
  INV_X1 U9897 ( .A(n14410), .ZN(n14402) );
  INV_X1 U9898 ( .A(n14633), .ZN(n14461) );
  NOR2_X1 U9899 ( .A1(n11386), .A2(n11385), .ZN(n11395) );
  NAND2_X1 U9900 ( .A1(n10851), .A2(n10850), .ZN(n10857) );
  AND2_X1 U9901 ( .A1(n9933), .A2(n12341), .ZN(n10633) );
  INV_X1 U9902 ( .A(n14938), .ZN(n11515) );
  OR2_X1 U9903 ( .A1(n14255), .A2(n9852), .ZN(n10557) );
  AND2_X1 U9904 ( .A1(n9984), .A2(n9387), .ZN(n10124) );
  NAND2_X1 U9905 ( .A1(n9991), .A2(n9990), .ZN(n12530) );
  AND4_X1 U9906 ( .A1(n8125), .A2(n8124), .A3(n8123), .A4(n8122), .ZN(n12754)
         );
  INV_X1 U9907 ( .A(n11268), .ZN(n11325) );
  INV_X1 U9908 ( .A(n12645), .ZN(n15430) );
  OAI21_X1 U9909 ( .B1(n12682), .B2(n12681), .A(n12680), .ZN(n12895) );
  NAND2_X1 U9910 ( .A1(n8284), .A2(n12186), .ZN(n15466) );
  NOR2_X1 U9911 ( .A1(n12794), .A2(n15521), .ZN(n12885) );
  AND3_X1 U9912 ( .A1(n8281), .A2(n8269), .A3(n8288), .ZN(n9863) );
  INV_X1 U9913 ( .A(n14790), .ZN(n15497) );
  INV_X1 U9914 ( .A(n15522), .ZN(n15517) );
  OR2_X1 U9915 ( .A1(n8036), .A2(n8069), .ZN(n8022) );
  XNOR2_X1 U9916 ( .A(n9154), .B(n9153), .ZN(n9394) );
  INV_X1 U9917 ( .A(n13503), .ZN(n13454) );
  NAND2_X1 U9918 ( .A1(n9471), .A2(n14827), .ZN(n13501) );
  INV_X1 U9919 ( .A(n6652), .ZN(n8935) );
  INV_X1 U9920 ( .A(n6860), .ZN(n9041) );
  INV_X1 U9921 ( .A(n15225), .ZN(n15264) );
  AND2_X1 U9922 ( .A1(n9419), .A2(n9418), .ZN(n15271) );
  INV_X1 U9923 ( .A(n14827), .ZN(n15279) );
  INV_X1 U9924 ( .A(n15292), .ZN(n13748) );
  INV_X1 U9925 ( .A(n15368), .ZN(n15380) );
  INV_X1 U9926 ( .A(n15350), .ZN(n15377) );
  AND2_X1 U9927 ( .A1(n9394), .A2(n9204), .ZN(n9466) );
  AND2_X1 U9928 ( .A1(n8571), .A2(n8588), .ZN(n9594) );
  INV_X1 U9929 ( .A(n14005), .ZN(n14937) );
  INV_X1 U9930 ( .A(n14932), .ZN(n13994) );
  AND4_X1 U9931 ( .A1(n11719), .A2(n11718), .A3(n11717), .A4(n11716), .ZN(
        n14532) );
  AND4_X1 U9932 ( .A1(n11409), .A2(n11408), .A3(n11407), .A4(n11406), .ZN(
        n14912) );
  OR2_X1 U9933 ( .A1(n9301), .A2(n9853), .ZN(n15100) );
  INV_X1 U9934 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9886) );
  INV_X1 U9935 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9911) );
  INV_X1 U9936 ( .A(n15061), .ZN(n15096) );
  INV_X1 U9937 ( .A(n15100), .ZN(n15068) );
  INV_X1 U9938 ( .A(n14420), .ZN(n14416) );
  INV_X1 U9939 ( .A(n14531), .ZN(n14571) );
  NOR2_X1 U9940 ( .A1(n10557), .A2(n10558), .ZN(n9931) );
  AND2_X1 U9941 ( .A1(n11129), .A2(n15175), .ZN(n14670) );
  AND2_X1 U9942 ( .A1(n9930), .A2(n9929), .ZN(n10034) );
  INV_X1 U9943 ( .A(n14670), .ZN(n15191) );
  NAND3_X1 U9944 ( .A1(n9584), .A2(n9583), .A3(n9585), .ZN(n9816) );
  INV_X1 U9945 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9220) );
  AND2_X1 U9946 ( .A1(n9369), .A2(n9378), .ZN(n11080) );
  INV_X1 U9947 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9289) );
  INV_X1 U9948 ( .A(n8388), .ZN(n8389) );
  INV_X1 U9949 ( .A(n15421), .ZN(n15405) );
  INV_X1 U9950 ( .A(n12530), .ZN(n11236) );
  NAND2_X1 U9951 ( .A1(n10010), .A2(n10124), .ZN(n12520) );
  INV_X1 U9952 ( .A(n12799), .ZN(n12538) );
  INV_X1 U9953 ( .A(n12652), .ZN(n15434) );
  NAND2_X1 U9954 ( .A1(n10159), .A2(n10144), .ZN(n15438) );
  NAND2_X1 U9955 ( .A1(n10159), .A2(n6642), .ZN(n15425) );
  AND2_X1 U9956 ( .A1(n12803), .A2(n12802), .ZN(n12936) );
  AND2_X1 U9957 ( .A1(n12851), .A2(n12850), .ZN(n12949) );
  INV_X1 U9958 ( .A(n15474), .ZN(n12752) );
  INV_X1 U9959 ( .A(n15547), .ZN(n15544) );
  INV_X1 U9960 ( .A(n12013), .ZN(n12960) );
  INV_X1 U9961 ( .A(n10846), .ZN(n11310) );
  NAND2_X1 U9962 ( .A1(n9388), .A2(n9387), .ZN(n9391) );
  AND2_X1 U9963 ( .A1(n8249), .A2(n8248), .ZN(n13016) );
  INV_X1 U9964 ( .A(SI_18_), .ZN(n9690) );
  INV_X1 U9965 ( .A(SI_13_), .ZN(n9375) );
  INV_X1 U9966 ( .A(n13750), .ZN(n14868) );
  INV_X1 U9967 ( .A(n13501), .ZN(n13461) );
  OR3_X1 U9968 ( .A1(n9479), .A2(n9478), .A3(n15368), .ZN(n13503) );
  INV_X1 U9969 ( .A(n13387), .ZN(n13507) );
  OR2_X1 U9970 ( .A1(n15204), .A2(P2_U3088), .ZN(n15278) );
  AND2_X1 U9971 ( .A1(n11625), .A2(n10284), .ZN(n13738) );
  OR3_X1 U9972 ( .A1(n11021), .A2(n11020), .A3(n9581), .ZN(n15399) );
  OR3_X1 U9973 ( .A1(n11021), .A2(n11020), .A3(n11019), .ZN(n15385) );
  INV_X2 U9974 ( .A(n15385), .ZN(n15387) );
  INV_X1 U9975 ( .A(n15305), .ZN(n15302) );
  INV_X1 U9976 ( .A(n8460), .ZN(n10899) );
  INV_X1 U9977 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9638) );
  INV_X1 U9978 ( .A(n14662), .ZN(n14534) );
  AND2_X1 U9979 ( .A1(n10533), .A2(n14258), .ZN(n14941) );
  AOI21_X2 U9980 ( .B1(n9842), .B2(n9825), .A(n15114), .ZN(n14005) );
  INV_X1 U9981 ( .A(n14532), .ZN(n14498) );
  INV_X1 U9982 ( .A(n14530), .ZN(n14265) );
  NOR2_X1 U9983 ( .A1(n9232), .A2(n10529), .ZN(P1_U4016) );
  NAND2_X1 U9984 ( .A1(n9299), .A2(n9298), .ZN(n15104) );
  OAI21_X1 U9985 ( .B1(n11794), .B2(n11793), .A(n14552), .ZN(n11808) );
  AND2_X1 U9986 ( .A1(n14488), .A2(n14487), .ZN(n14648) );
  AND2_X2 U9987 ( .A1(n11803), .A2(n14578), .ZN(n15129) );
  INV_X1 U9988 ( .A(n15202), .ZN(n15200) );
  AND2_X2 U9989 ( .A1(n9931), .A2(n10034), .ZN(n15202) );
  AND2_X2 U9990 ( .A1(n9846), .A2(n9816), .ZN(n15160) );
  INV_X1 U9991 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10385) );
  INV_X1 U9992 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9683) );
  INV_X2 U9993 ( .A(n12550), .ZN(P3_U3897) );
  NAND2_X1 U9994 ( .A1(n8295), .A2(n8294), .ZN(P3_U3456) );
  AND2_X1 U9995 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9395), .ZN(P2_U3947) );
  XNOR2_X1 U9996 ( .A(n8402), .B(n8401), .ZN(SUB_1596_U4) );
  NOR2_X1 U9997 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_16__SCAN_IN), .ZN(
        n7690) );
  NAND4_X1 U9998 ( .A1(n7692), .A2(n7953), .A3(n7922), .A4(n7691), .ZN(n7693)
         );
  NOR2_X1 U9999 ( .A1(P3_IR_REG_25__SCAN_IN), .A2(P3_IR_REG_24__SCAN_IN), .ZN(
        n7696) );
  XNOR2_X2 U10000 ( .A(n7698), .B(n13019), .ZN(n7702) );
  INV_X1 U10001 ( .A(n7702), .ZN(n7703) );
  NAND2_X1 U10002 ( .A1(n7773), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7700) );
  MUX2_X1 U10003 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7700), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n7701) );
  AND2_X2 U10004 ( .A1(n7703), .A2(n13027), .ZN(n7799) );
  NAND2_X1 U10005 ( .A1(n12001), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n7709) );
  INV_X2 U10006 ( .A(n7932), .ZN(n12002) );
  NAND2_X1 U10007 ( .A1(n12002), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n7708) );
  NOR2_X1 U10008 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n7839) );
  NAND2_X1 U10009 ( .A1(n7839), .A2(n10418), .ZN(n7854) );
  NAND2_X1 U10010 ( .A1(n7976), .A2(n11607), .ZN(n7991) );
  INV_X1 U10011 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n8026) );
  INV_X1 U10012 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n8040) );
  INV_X1 U10013 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n12490) );
  NAND2_X1 U10014 ( .A1(n8084), .A2(n12490), .ZN(n8098) );
  INV_X1 U10015 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n12400) );
  INV_X1 U10016 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n12480) );
  INV_X1 U10017 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n12393) );
  INV_X1 U10018 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n12418) );
  NAND2_X1 U10019 ( .A1(n8169), .A2(n12418), .ZN(n12657) );
  OR2_X1 U10020 ( .A1(n8169), .A2(n12418), .ZN(n7704) );
  NAND2_X1 U10021 ( .A1(n12657), .A2(n7704), .ZN(n12672) );
  NAND2_X1 U10022 ( .A1(n8186), .A2(n12672), .ZN(n7707) );
  AND2_X2 U10023 ( .A1(n7702), .A2(n7705), .ZN(n7853) );
  NAND2_X1 U10024 ( .A1(n7929), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n7706) );
  INV_X1 U10025 ( .A(n12683), .ZN(n12537) );
  INV_X1 U10026 ( .A(n7794), .ZN(n7710) );
  NAND2_X1 U10027 ( .A1(n7787), .A2(n7710), .ZN(n7712) );
  INV_X1 U10028 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9349) );
  NAND2_X1 U10029 ( .A1(n9349), .A2(n6866), .ZN(n7711) );
  NAND2_X1 U10030 ( .A1(n7712), .A2(n7711), .ZN(n7806) );
  NAND2_X1 U10031 ( .A1(n7806), .A2(n7805), .ZN(n7714) );
  NAND2_X1 U10032 ( .A1(n9337), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7713) );
  NAND2_X1 U10033 ( .A1(n7714), .A2(n7713), .ZN(n7816) );
  NAND2_X1 U10034 ( .A1(n7816), .A2(n7815), .ZN(n7716) );
  INV_X1 U10035 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9345) );
  NAND2_X1 U10036 ( .A1(n9345), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7715) );
  NAND2_X1 U10037 ( .A1(n7716), .A2(n7715), .ZN(n7835) );
  NAND2_X1 U10038 ( .A1(n7835), .A2(n7834), .ZN(n7718) );
  NAND2_X1 U10039 ( .A1(n9327), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7717) );
  NAND2_X1 U10040 ( .A1(n7718), .A2(n7717), .ZN(n7846) );
  NAND2_X1 U10041 ( .A1(n7846), .A2(n7845), .ZN(n7720) );
  NAND2_X1 U10042 ( .A1(n9342), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n7719) );
  NAND2_X1 U10043 ( .A1(n10552), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7722) );
  XNOR2_X1 U10044 ( .A(n7724), .B(P1_DATAO_REG_7__SCAN_IN), .ZN(n7875) );
  INV_X1 U10045 ( .A(n7875), .ZN(n7723) );
  NAND2_X1 U10046 ( .A1(n7724), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7725) );
  NAND2_X1 U10047 ( .A1(n7727), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7728) );
  XNOR2_X1 U10048 ( .A(n9373), .B(P2_DATAO_REG_9__SCAN_IN), .ZN(n7906) );
  INV_X1 U10049 ( .A(n7906), .ZN(n7729) );
  NAND2_X1 U10050 ( .A1(n7907), .A2(n7729), .ZN(n7731) );
  NAND2_X1 U10051 ( .A1(n13149), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n7730) );
  XNOR2_X1 U10052 ( .A(n7733), .B(P1_DATAO_REG_10__SCAN_IN), .ZN(n7920) );
  INV_X1 U10053 ( .A(n7920), .ZN(n7732) );
  NAND2_X1 U10054 ( .A1(n7733), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n7734) );
  NAND2_X1 U10055 ( .A1(n9555), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n7736) );
  NAND2_X1 U10056 ( .A1(n9488), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n7738) );
  NAND2_X1 U10057 ( .A1(n9444), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n7737) );
  NAND2_X1 U10058 ( .A1(n7738), .A2(n7737), .ZN(n7956) );
  NAND2_X1 U10059 ( .A1(n9683), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n7741) );
  INV_X1 U10060 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n9684) );
  NAND2_X1 U10061 ( .A1(n9684), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n7740) );
  NAND2_X1 U10062 ( .A1(n9703), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n7743) );
  NAND2_X1 U10063 ( .A1(n13278), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n7742) );
  NAND2_X1 U10064 ( .A1(n9779), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n7745) );
  NAND2_X1 U10065 ( .A1(n9781), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n7744) );
  NAND2_X1 U10066 ( .A1(n9876), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n7748) );
  NAND2_X1 U10067 ( .A1(n9915), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n7746) );
  NAND2_X1 U10068 ( .A1(n7748), .A2(n7746), .ZN(n8033) );
  INV_X1 U10069 ( .A(n8033), .ZN(n7747) );
  INV_X1 U10070 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10120) );
  NAND2_X1 U10071 ( .A1(n10120), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n7751) );
  INV_X1 U10072 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10122) );
  NAND2_X1 U10073 ( .A1(n10122), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n7750) );
  NAND2_X1 U10074 ( .A1(n10385), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n7753) );
  NAND2_X1 U10075 ( .A1(n10623), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n7752) );
  INV_X1 U10076 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11724) );
  NAND2_X1 U10077 ( .A1(n11724), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n7758) );
  INV_X1 U10078 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n10900) );
  NAND2_X1 U10079 ( .A1(n10900), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n7757) );
  NAND2_X1 U10080 ( .A1(n7758), .A2(n7757), .ZN(n8091) );
  INV_X1 U10081 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11027) );
  XNOR2_X1 U10082 ( .A(n11027), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n8106) );
  NAND2_X1 U10083 ( .A1(n11027), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n7759) );
  XNOR2_X1 U10084 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n8116) );
  NAND2_X1 U10085 ( .A1(n8117), .A2(n8116), .ZN(n7762) );
  INV_X1 U10086 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11139) );
  NAND2_X1 U10087 ( .A1(n11139), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7761) );
  INV_X1 U10088 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11351) );
  INV_X1 U10089 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n11471) );
  NAND2_X1 U10090 ( .A1(n11471), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n7764) );
  INV_X1 U10091 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n11657) );
  NAND2_X1 U10092 ( .A1(n11657), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n7765) );
  INV_X1 U10093 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13853) );
  NOR2_X1 U10094 ( .A1(n13853), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n7767) );
  NAND2_X1 U10095 ( .A1(n13853), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n7768) );
  INV_X1 U10096 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n11632) );
  AND2_X1 U10097 ( .A1(n11632), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n7769) );
  INV_X1 U10098 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n11911) );
  XNOR2_X1 U10099 ( .A(n8998), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n7770) );
  XNOR2_X1 U10100 ( .A(n8178), .B(n7770), .ZN(n11978) );
  NAND2_X1 U10101 ( .A1(n7771), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7772) );
  NAND2_X2 U10102 ( .A1(n7774), .A2(n7773), .ZN(n8201) );
  XNOR2_X2 U10103 ( .A(n7777), .B(n7776), .ZN(n10132) );
  NAND2_X4 U10104 ( .A1(n8201), .A2(n10132), .ZN(n10127) );
  INV_X2 U10105 ( .A(n11734), .ZN(n9800) );
  NAND2_X1 U10106 ( .A1(n11978), .A2(n11998), .ZN(n7781) );
  NAND2_X1 U10107 ( .A1(n6650), .A2(SI_28_), .ZN(n7780) );
  NAND2_X1 U10108 ( .A1(n7853), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7785) );
  NAND2_X1 U10109 ( .A1(n7799), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n7784) );
  NAND2_X1 U10110 ( .A1(n8186), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n7783) );
  NAND2_X1 U10111 ( .A1(n7800), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n7782) );
  NAND2_X1 U10112 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n7786) );
  XNOR2_X2 U10113 ( .A(n7197), .B(n7786), .ZN(n10253) );
  INV_X1 U10114 ( .A(SI_1_), .ZN(n9322) );
  XNOR2_X1 U10115 ( .A(n7787), .B(n7794), .ZN(n9323) );
  INV_X1 U10116 ( .A(n9998), .ZN(n7796) );
  NAND2_X1 U10117 ( .A1(n7853), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n7792) );
  NAND2_X1 U10118 ( .A1(n7799), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7791) );
  NAND2_X1 U10119 ( .A1(n8186), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n7790) );
  NAND2_X1 U10120 ( .A1(n7800), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n7789) );
  INV_X1 U10121 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n9335) );
  INV_X1 U10122 ( .A(SI_0_), .ZN(n9333) );
  NAND2_X1 U10123 ( .A1(n6942), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7793) );
  AND2_X1 U10124 ( .A1(n7794), .A2(n7793), .ZN(n9334) );
  NAND2_X1 U10125 ( .A1(n15463), .A2(n10114), .ZN(n15465) );
  NAND2_X1 U10126 ( .A1(n10025), .A2(n15465), .ZN(n7798) );
  NAND2_X1 U10127 ( .A1(n15451), .A2(n7796), .ZN(n7797) );
  NAND2_X1 U10128 ( .A1(n7798), .A2(n7797), .ZN(n15447) );
  NAND2_X1 U10129 ( .A1(n7853), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7804) );
  NAND2_X1 U10130 ( .A1(n8186), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n7802) );
  NAND2_X1 U10131 ( .A1(n7800), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n7801) );
  XNOR2_X1 U10132 ( .A(n7806), .B(n7805), .ZN(n9328) );
  OR2_X1 U10133 ( .A1(n8095), .A2(n9328), .ZN(n7808) );
  OAI211_X1 U10134 ( .C1(n10317), .C2(n10127), .A(n7808), .B(n7807), .ZN(
        n15442) );
  NAND2_X1 U10135 ( .A1(n15447), .A2(n8206), .ZN(n7810) );
  INV_X1 U10136 ( .A(n15462), .ZN(n10482) );
  NAND2_X1 U10137 ( .A1(n10482), .A2(n15442), .ZN(n7809) );
  NAND2_X1 U10138 ( .A1(n7810), .A2(n7809), .ZN(n10485) );
  INV_X1 U10139 ( .A(n10485), .ZN(n7825) );
  NAND2_X1 U10140 ( .A1(n7853), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7814) );
  NAND2_X1 U10141 ( .A1(n12001), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7813) );
  INV_X1 U10142 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n10488) );
  NAND2_X1 U10143 ( .A1(n12002), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n7811) );
  OR2_X1 U10144 ( .A1(n11999), .A2(SI_3_), .ZN(n7822) );
  XNOR2_X1 U10145 ( .A(n7816), .B(n7815), .ZN(n13382) );
  OR2_X1 U10146 ( .A1(n8095), .A2(n13382), .ZN(n7821) );
  NAND2_X1 U10147 ( .A1(n7817), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7819) );
  INV_X1 U10148 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n7818) );
  XNOR2_X1 U10149 ( .A(n7819), .B(n7818), .ZN(n10431) );
  NAND2_X1 U10150 ( .A1(n8072), .A2(n10431), .ZN(n7820) );
  NAND2_X1 U10151 ( .A1(n15449), .A2(n15487), .ZN(n12058) );
  INV_X2 U10152 ( .A(n15449), .ZN(n12549) );
  INV_X1 U10153 ( .A(n15487), .ZN(n7823) );
  NAND2_X1 U10154 ( .A1(n12549), .A2(n7823), .ZN(n12043) );
  NAND2_X1 U10155 ( .A1(n7825), .A2(n7824), .ZN(n10483) );
  NAND2_X1 U10156 ( .A1(n12549), .A2(n15487), .ZN(n7826) );
  NAND2_X1 U10157 ( .A1(n10483), .A2(n7826), .ZN(n10376) );
  NAND2_X1 U10158 ( .A1(n7853), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7830) );
  NAND2_X1 U10159 ( .A1(n7799), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7829) );
  OR2_X1 U10160 ( .A1(n7680), .A2(n7839), .ZN(n10382) );
  NAND2_X1 U10161 ( .A1(n8186), .A2(n10382), .ZN(n7828) );
  NAND2_X1 U10162 ( .A1(n12002), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n7827) );
  NAND4_X1 U10163 ( .A1(n7830), .A2(n7829), .A3(n7828), .A4(n7827), .ZN(n12548) );
  NAND2_X1 U10164 ( .A1(n7831), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7833) );
  INV_X1 U10165 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7832) );
  XNOR2_X1 U10166 ( .A(n7833), .B(n7832), .ZN(n10167) );
  INV_X1 U10167 ( .A(n10167), .ZN(n10405) );
  XNOR2_X1 U10168 ( .A(n7835), .B(n7834), .ZN(n9315) );
  OR2_X1 U10169 ( .A1(n8095), .A2(n9315), .ZN(n7837) );
  OR2_X1 U10170 ( .A1(n11999), .A2(SI_4_), .ZN(n7836) );
  OAI211_X1 U10171 ( .C1(n10405), .C2(n10127), .A(n7837), .B(n7836), .ZN(
        n12064) );
  XNOR2_X1 U10172 ( .A(n12548), .B(n12064), .ZN(n12061) );
  INV_X1 U10173 ( .A(n12064), .ZN(n10280) );
  NAND2_X1 U10174 ( .A1(n12548), .A2(n10280), .ZN(n7838) );
  NAND2_X1 U10175 ( .A1(n7853), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7844) );
  NAND2_X1 U10176 ( .A1(n12001), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7843) );
  OR2_X1 U10177 ( .A1(n7839), .A2(n10418), .ZN(n7840) );
  NAND2_X1 U10178 ( .A1(n7854), .A2(n7840), .ZN(n10983) );
  NAND2_X1 U10179 ( .A1(n8170), .A2(n10983), .ZN(n7842) );
  NAND2_X1 U10180 ( .A1(n8171), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n7841) );
  AND4_X2 U10181 ( .A1(n7844), .A2(n7843), .A3(n7842), .A4(n7841), .ZN(n10963)
         );
  OR2_X1 U10182 ( .A1(n11999), .A2(SI_5_), .ZN(n7851) );
  XNOR2_X1 U10183 ( .A(n7846), .B(n7845), .ZN(n9313) );
  OR2_X1 U10184 ( .A1(n8095), .A2(n9313), .ZN(n7850) );
  OR2_X1 U10185 ( .A1(n7847), .A2(n8069), .ZN(n7848) );
  INV_X1 U10186 ( .A(n10168), .ZN(n10428) );
  NAND2_X1 U10187 ( .A1(n8072), .A2(n10428), .ZN(n7849) );
  NAND2_X1 U10188 ( .A1(n10963), .A2(n10476), .ZN(n12071) );
  INV_X1 U10189 ( .A(n10963), .ZN(n10468) );
  INV_X1 U10190 ( .A(n10476), .ZN(n10982) );
  NAND2_X1 U10191 ( .A1(n10468), .A2(n10982), .ZN(n12070) );
  NAND2_X1 U10192 ( .A1(n10963), .A2(n10982), .ZN(n7852) );
  NAND2_X1 U10193 ( .A1(n10977), .A2(n7852), .ZN(n10960) );
  INV_X1 U10194 ( .A(n10960), .ZN(n7867) );
  NAND2_X1 U10195 ( .A1(n7853), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n7859) );
  NAND2_X1 U10196 ( .A1(n12001), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7858) );
  NAND2_X1 U10197 ( .A1(n7854), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7855) );
  NAND2_X1 U10198 ( .A1(n7869), .A2(n7855), .ZN(n10970) );
  NAND2_X1 U10199 ( .A1(n8170), .A2(n10970), .ZN(n7857) );
  NAND2_X1 U10200 ( .A1(n8171), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n7856) );
  NAND2_X1 U10201 ( .A1(n7860), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7862) );
  INV_X1 U10202 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n7861) );
  XNOR2_X1 U10203 ( .A(n7862), .B(n7861), .ZN(n10458) );
  INV_X1 U10204 ( .A(SI_6_), .ZN(n9331) );
  OR2_X1 U10205 ( .A1(n11999), .A2(n9331), .ZN(n7866) );
  XNOR2_X1 U10206 ( .A(n9350), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n7863) );
  XNOR2_X1 U10207 ( .A(n7864), .B(n7863), .ZN(n9332) );
  OR2_X1 U10208 ( .A1(n8095), .A2(n9332), .ZN(n7865) );
  OAI211_X1 U10209 ( .C1(n10127), .C2(n10458), .A(n7866), .B(n7865), .ZN(
        n10660) );
  NAND2_X1 U10210 ( .A1(n10947), .A2(n10660), .ZN(n12074) );
  INV_X1 U10211 ( .A(n10660), .ZN(n10969) );
  NAND2_X1 U10212 ( .A1(n12547), .A2(n10969), .ZN(n12075) );
  NAND2_X1 U10213 ( .A1(n7867), .A2(n7078), .ZN(n10962) );
  NAND2_X1 U10214 ( .A1(n12547), .A2(n10660), .ZN(n7868) );
  NAND2_X1 U10215 ( .A1(n10962), .A2(n7868), .ZN(n10946) );
  NAND2_X1 U10216 ( .A1(n7853), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n7874) );
  NAND2_X1 U10217 ( .A1(n7799), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7873) );
  AND2_X1 U10218 ( .A1(n7869), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7870) );
  OR2_X1 U10219 ( .A1(n7870), .A2(n7887), .ZN(n10951) );
  NAND2_X1 U10220 ( .A1(n8186), .A2(n10951), .ZN(n7872) );
  NAND2_X1 U10221 ( .A1(n7800), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n7871) );
  OR2_X1 U10222 ( .A1(n11999), .A2(SI_7_), .ZN(n7884) );
  XNOR2_X1 U10223 ( .A(n7876), .B(n7875), .ZN(n9317) );
  OR2_X1 U10224 ( .A1(n8095), .A2(n9317), .ZN(n7883) );
  NAND2_X1 U10225 ( .A1(n7878), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7879) );
  MUX2_X1 U10226 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7879), .S(
        P3_IR_REG_7__SCAN_IN), .Z(n7881) );
  NAND2_X1 U10227 ( .A1(n7881), .A2(n7908), .ZN(n10502) );
  NAND2_X1 U10228 ( .A1(n8072), .A2(n10502), .ZN(n7882) );
  NAND2_X1 U10229 ( .A1(n12431), .A2(n10778), .ZN(n12080) );
  INV_X1 U10230 ( .A(n10778), .ZN(n15509) );
  NAND2_X1 U10231 ( .A1(n12546), .A2(n15509), .ZN(n12081) );
  NAND2_X1 U10232 ( .A1(n10946), .A2(n12022), .ZN(n10945) );
  NAND2_X1 U10233 ( .A1(n12546), .A2(n10778), .ZN(n7885) );
  NAND2_X1 U10234 ( .A1(n7853), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7892) );
  NAND2_X1 U10235 ( .A1(n7799), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7891) );
  NOR2_X1 U10236 ( .A1(n7887), .A2(n7886), .ZN(n7888) );
  OR2_X1 U10237 ( .A1(n7900), .A2(n7888), .ZN(n12433) );
  NAND2_X1 U10238 ( .A1(n8170), .A2(n12433), .ZN(n7890) );
  NAND2_X1 U10239 ( .A1(n8171), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n7889) );
  NAND2_X1 U10240 ( .A1(n7908), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7894) );
  INV_X1 U10241 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n7893) );
  INV_X1 U10242 ( .A(SI_8_), .ZN(n9320) );
  OR2_X1 U10243 ( .A1(n11999), .A2(n9320), .ZN(n7898) );
  XNOR2_X1 U10244 ( .A(n7896), .B(n7895), .ZN(n9321) );
  OR2_X1 U10245 ( .A1(n8095), .A2(n9321), .ZN(n7897) );
  OAI211_X1 U10246 ( .C1(n10127), .C2(n10928), .A(n7898), .B(n7897), .ZN(
        n12429) );
  NAND2_X1 U10247 ( .A1(n11142), .A2(n12429), .ZN(n12085) );
  INV_X1 U10248 ( .A(n11142), .ZN(n12545) );
  INV_X1 U10249 ( .A(n12429), .ZN(n11220) );
  NAND2_X1 U10250 ( .A1(n12545), .A2(n11220), .ZN(n12086) );
  NAND2_X1 U10251 ( .A1(n12085), .A2(n12086), .ZN(n12021) );
  NAND2_X1 U10252 ( .A1(n11142), .A2(n11220), .ZN(n7899) );
  NAND2_X1 U10253 ( .A1(n7929), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n7905) );
  NAND2_X1 U10254 ( .A1(n7799), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7904) );
  OR2_X1 U10255 ( .A1(n7900), .A2(n13326), .ZN(n7901) );
  NAND2_X1 U10256 ( .A1(n7914), .A2(n7901), .ZN(n11147) );
  NAND2_X1 U10257 ( .A1(n8170), .A2(n11147), .ZN(n7903) );
  NAND2_X1 U10258 ( .A1(n12002), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n7902) );
  NAND4_X1 U10259 ( .A1(n7905), .A2(n7904), .A3(n7903), .A4(n7902), .ZN(n12544) );
  XNOR2_X1 U10260 ( .A(n7907), .B(n7906), .ZN(n9324) );
  OR2_X1 U10261 ( .A1(n8095), .A2(n9324), .ZN(n7912) );
  OR2_X1 U10262 ( .A1(n11999), .A2(SI_9_), .ZN(n7911) );
  NOR2_X1 U10263 ( .A1(n7908), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n7923) );
  OR2_X1 U10264 ( .A1(n7923), .A2(n8069), .ZN(n7909) );
  XNOR2_X1 U10265 ( .A(n7909), .B(n7922), .ZN(n10929) );
  NAND2_X1 U10266 ( .A1(n8072), .A2(n10929), .ZN(n7910) );
  XNOR2_X1 U10267 ( .A(n12544), .B(n10846), .ZN(n12088) );
  NAND2_X1 U10268 ( .A1(n12544), .A2(n10846), .ZN(n7913) );
  NAND2_X1 U10269 ( .A1(n7853), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7919) );
  NAND2_X1 U10270 ( .A1(n7799), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7918) );
  NAND2_X1 U10271 ( .A1(n7914), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7915) );
  NAND2_X1 U10272 ( .A1(n7930), .A2(n7915), .ZN(n10905) );
  NAND2_X1 U10273 ( .A1(n8170), .A2(n10905), .ZN(n7917) );
  NAND2_X1 U10274 ( .A1(n8171), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n7916) );
  XNOR2_X1 U10275 ( .A(n7921), .B(n7920), .ZN(n9338) );
  OR2_X1 U10276 ( .A1(n8095), .A2(n9338), .ZN(n7928) );
  OR2_X1 U10277 ( .A1(n11999), .A2(SI_10_), .ZN(n7927) );
  NAND2_X1 U10278 ( .A1(n7923), .A2(n7922), .ZN(n7937) );
  NAND2_X1 U10279 ( .A1(n7937), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7925) );
  INV_X1 U10280 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n7924) );
  NAND2_X1 U10281 ( .A1(n8072), .A2(n15417), .ZN(n7926) );
  NAND2_X1 U10282 ( .A1(n11443), .A2(n11336), .ZN(n12096) );
  INV_X1 U10283 ( .A(n11336), .ZN(n15520) );
  NAND2_X1 U10284 ( .A1(n12543), .A2(n15520), .ZN(n12101) );
  NAND2_X1 U10285 ( .A1(n12096), .A2(n12101), .ZN(n12093) );
  NAND2_X1 U10286 ( .A1(n12543), .A2(n11336), .ZN(n11441) );
  NAND2_X1 U10287 ( .A1(n7929), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n7936) );
  NAND2_X1 U10288 ( .A1(n7799), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n7935) );
  NAND2_X1 U10289 ( .A1(n7930), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7931) );
  NAND2_X1 U10290 ( .A1(n7944), .A2(n7931), .ZN(n11447) );
  NAND2_X1 U10291 ( .A1(n8170), .A2(n11447), .ZN(n7934) );
  INV_X2 U10292 ( .A(n7932), .ZN(n8171) );
  NAND2_X1 U10293 ( .A1(n8171), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n7933) );
  NAND2_X1 U10294 ( .A1(n7950), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7939) );
  INV_X1 U10295 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n7938) );
  XNOR2_X1 U10296 ( .A(n7939), .B(n7938), .ZN(n11268) );
  OR2_X1 U10297 ( .A1(n11999), .A2(SI_11_), .ZN(n7943) );
  XNOR2_X1 U10298 ( .A(n9555), .B(P2_DATAO_REG_11__SCAN_IN), .ZN(n7940) );
  XNOR2_X1 U10299 ( .A(n7941), .B(n7940), .ZN(n9346) );
  OR2_X1 U10300 ( .A1(n8095), .A2(n9346), .ZN(n7942) );
  OAI211_X1 U10301 ( .C1(n11325), .C2(n10127), .A(n7943), .B(n7942), .ZN(
        n11446) );
  INV_X1 U10302 ( .A(n11446), .ZN(n12103) );
  NAND2_X1 U10303 ( .A1(n12542), .A2(n12103), .ZN(n14772) );
  NAND2_X1 U10304 ( .A1(n7799), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7949) );
  NAND2_X1 U10305 ( .A1(n12002), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n7948) );
  AND2_X1 U10306 ( .A1(n7944), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7945) );
  OR2_X1 U10307 ( .A1(n7945), .A2(n7976), .ZN(n14781) );
  NAND2_X1 U10308 ( .A1(n8170), .A2(n14781), .ZN(n7947) );
  NAND2_X1 U10309 ( .A1(n7929), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n7946) );
  INV_X1 U10310 ( .A(n14762), .ZN(n12541) );
  NOR2_X1 U10311 ( .A1(n7954), .A2(n8069), .ZN(n7951) );
  MUX2_X1 U10312 ( .A(n8069), .B(n7951), .S(P3_IR_REG_12__SCAN_IN), .Z(n7952)
         );
  INV_X1 U10313 ( .A(n7952), .ZN(n7955) );
  NAND2_X1 U10314 ( .A1(n7954), .A2(n7953), .ZN(n7986) );
  NAND2_X1 U10315 ( .A1(n7957), .A2(n7956), .ZN(n7958) );
  NAND2_X1 U10316 ( .A1(n7959), .A2(n7958), .ZN(n9366) );
  OR2_X1 U10317 ( .A1(n8095), .A2(n9366), .ZN(n7961) );
  OR2_X1 U10318 ( .A1(n11999), .A2(n9367), .ZN(n7960) );
  OAI211_X1 U10319 ( .C1(n10127), .C2(n11892), .A(n7961), .B(n7960), .ZN(
        n11346) );
  NAND2_X1 U10320 ( .A1(n12541), .A2(n11346), .ZN(n7963) );
  AND2_X1 U10321 ( .A1(n14772), .A2(n7963), .ZN(n7965) );
  AND2_X1 U10322 ( .A1(n11441), .A2(n7965), .ZN(n7962) );
  INV_X1 U10323 ( .A(n7963), .ZN(n7964) );
  NAND2_X1 U10324 ( .A1(n14762), .A2(n11346), .ZN(n12111) );
  INV_X1 U10325 ( .A(n11346), .ZN(n14780) );
  NAND2_X1 U10326 ( .A1(n12541), .A2(n14780), .ZN(n12102) );
  NAND2_X1 U10327 ( .A1(n12111), .A2(n12102), .ZN(n14774) );
  OR2_X1 U10328 ( .A1(n7964), .A2(n14774), .ZN(n7968) );
  INV_X1 U10329 ( .A(n7965), .ZN(n7966) );
  NAND2_X1 U10330 ( .A1(n14777), .A2(n11446), .ZN(n14770) );
  OR2_X1 U10331 ( .A1(n7966), .A2(n14770), .ZN(n7967) );
  INV_X1 U10332 ( .A(n7969), .ZN(n7970) );
  NAND2_X1 U10333 ( .A1(n7970), .A2(n9638), .ZN(n7971) );
  NAND2_X1 U10334 ( .A1(n7972), .A2(n7971), .ZN(n9374) );
  OR2_X1 U10335 ( .A1(n9374), .A2(n8095), .ZN(n7975) );
  NAND2_X1 U10336 ( .A1(n7986), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7973) );
  XNOR2_X1 U10337 ( .A(n7973), .B(P3_IR_REG_13__SCAN_IN), .ZN(n12564) );
  AOI22_X1 U10338 ( .A1(n6650), .A2(SI_13_), .B1(n8072), .B2(n12564), .ZN(
        n7974) );
  NAND2_X1 U10339 ( .A1(n7929), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n7981) );
  NAND2_X1 U10340 ( .A1(n7799), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n7980) );
  OR2_X1 U10341 ( .A1(n7976), .A2(n11607), .ZN(n7977) );
  NAND2_X1 U10342 ( .A1(n7991), .A2(n7977), .ZN(n14765) );
  NAND2_X1 U10343 ( .A1(n8170), .A2(n14765), .ZN(n7979) );
  NAND2_X1 U10344 ( .A1(n8171), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n7978) );
  NAND4_X1 U10345 ( .A1(n7981), .A2(n7980), .A3(n7979), .A4(n7978), .ZN(n12540) );
  NAND2_X1 U10346 ( .A1(n14764), .A2(n12540), .ZN(n12112) );
  NAND2_X1 U10347 ( .A1(n11609), .A2(n14778), .ZN(n12113) );
  NAND2_X1 U10348 ( .A1(n12112), .A2(n12113), .ZN(n14759) );
  OR2_X1 U10349 ( .A1(n7983), .A2(n7982), .ZN(n7984) );
  NAND2_X1 U10350 ( .A1(n7985), .A2(n7984), .ZN(n9376) );
  NAND2_X1 U10351 ( .A1(n9376), .A2(n11998), .ZN(n7990) );
  NAND2_X1 U10352 ( .A1(n8003), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7988) );
  XNOR2_X1 U10353 ( .A(n7988), .B(n7987), .ZN(n12578) );
  AOI22_X1 U10354 ( .A1(n6650), .A2(n9377), .B1(n8072), .B2(n12578), .ZN(n7989) );
  NAND2_X1 U10355 ( .A1(n7990), .A2(n7989), .ZN(n14789) );
  NAND2_X1 U10356 ( .A1(n12001), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n7996) );
  NAND2_X1 U10357 ( .A1(n7929), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n7995) );
  NAND2_X1 U10358 ( .A1(n7991), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7992) );
  NAND2_X1 U10359 ( .A1(n8010), .A2(n7992), .ZN(n12880) );
  NAND2_X1 U10360 ( .A1(n8170), .A2(n12880), .ZN(n7994) );
  NAND2_X1 U10361 ( .A1(n8171), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n7993) );
  NAND4_X1 U10362 ( .A1(n7996), .A2(n7995), .A3(n7994), .A4(n7993), .ZN(n12539) );
  XNOR2_X1 U10363 ( .A(n14789), .B(n12539), .ZN(n12877) );
  NAND2_X1 U10364 ( .A1(n12876), .A2(n12877), .ZN(n7998) );
  INV_X1 U10365 ( .A(n14789), .ZN(n12884) );
  NAND2_X1 U10366 ( .A1(n12884), .A2(n12539), .ZN(n7997) );
  OR2_X1 U10367 ( .A1(n8000), .A2(n7999), .ZN(n8001) );
  AND2_X1 U10368 ( .A1(n8002), .A2(n8001), .ZN(n9545) );
  NAND2_X1 U10369 ( .A1(n9545), .A2(n11998), .ZN(n8009) );
  NOR2_X1 U10370 ( .A1(n8006), .A2(n8069), .ZN(n8004) );
  MUX2_X1 U10371 ( .A(n8069), .B(n8004), .S(P3_IR_REG_15__SCAN_IN), .Z(n8007)
         );
  INV_X1 U10372 ( .A(n11896), .ZN(n12597) );
  AOI22_X1 U10373 ( .A1(n12597), .A2(n8072), .B1(n6650), .B2(SI_15_), .ZN(
        n8008) );
  NAND2_X1 U10374 ( .A1(n8009), .A2(n8008), .ZN(n12360) );
  NAND2_X1 U10375 ( .A1(n7929), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8016) );
  NAND2_X1 U10376 ( .A1(n12001), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8015) );
  INV_X1 U10377 ( .A(n8027), .ZN(n8012) );
  NAND2_X1 U10378 ( .A1(n8010), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8011) );
  NAND2_X1 U10379 ( .A1(n8012), .A2(n8011), .ZN(n12865) );
  NAND2_X1 U10380 ( .A1(n8170), .A2(n12865), .ZN(n8014) );
  NAND2_X1 U10381 ( .A1(n8171), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8013) );
  NAND4_X1 U10382 ( .A1(n8016), .A2(n8015), .A3(n8014), .A4(n8013), .ZN(n12848) );
  AND2_X1 U10383 ( .A1(n12360), .A2(n12848), .ZN(n8018) );
  NAND2_X1 U10384 ( .A1(n13015), .A2(n12879), .ZN(n8017) );
  OR2_X1 U10385 ( .A1(n9606), .A2(n8095), .ZN(n8025) );
  INV_X1 U10386 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8035) );
  OAI22_X1 U10387 ( .A1(n11899), .A2(n10127), .B1(n11999), .B2(n9607), .ZN(
        n8023) );
  INV_X1 U10388 ( .A(n8023), .ZN(n8024) );
  NAND2_X1 U10389 ( .A1(n7929), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8032) );
  NAND2_X1 U10390 ( .A1(n12001), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8031) );
  NOR2_X1 U10391 ( .A1(n8027), .A2(n8026), .ZN(n8028) );
  OR2_X1 U10392 ( .A1(n8041), .A2(n8028), .ZN(n12854) );
  NAND2_X1 U10393 ( .A1(n8170), .A2(n12854), .ZN(n8030) );
  NAND2_X1 U10394 ( .A1(n8171), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8029) );
  NAND4_X1 U10395 ( .A1(n8032), .A2(n8031), .A3(n8030), .A4(n8029), .ZN(n12833) );
  NAND2_X1 U10396 ( .A1(n13008), .A2(n12861), .ZN(n12837) );
  XNOR2_X1 U10397 ( .A(n8034), .B(n8033), .ZN(n9686) );
  NAND2_X1 U10398 ( .A1(n9686), .A2(n11998), .ZN(n8039) );
  NAND2_X1 U10399 ( .A1(n8036), .A2(n8035), .ZN(n8052) );
  NAND2_X1 U10400 ( .A1(n8052), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8037) );
  XNOR2_X1 U10401 ( .A(n8037), .B(P3_IR_REG_17__SCAN_IN), .ZN(n12633) );
  AOI22_X1 U10402 ( .A1(n12633), .A2(n8072), .B1(SI_17_), .B2(n6650), .ZN(
        n8038) );
  NAND2_X1 U10403 ( .A1(n8039), .A2(n8038), .ZN(n12465) );
  NAND2_X1 U10404 ( .A1(n7929), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8046) );
  NAND2_X1 U10405 ( .A1(n12001), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8045) );
  OR2_X1 U10406 ( .A1(n8041), .A2(n8040), .ZN(n8042) );
  NAND2_X1 U10407 ( .A1(n8056), .A2(n8042), .ZN(n12840) );
  NAND2_X1 U10408 ( .A1(n8170), .A2(n12840), .ZN(n8044) );
  NAND2_X1 U10409 ( .A1(n8171), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8043) );
  OR2_X1 U10410 ( .A1(n12465), .A2(n12816), .ZN(n12819) );
  NAND2_X1 U10411 ( .A1(n12465), .A2(n12816), .ZN(n12128) );
  OR2_X1 U10412 ( .A1(n8049), .A2(n8048), .ZN(n8050) );
  NAND2_X1 U10413 ( .A1(n8051), .A2(n8050), .ZN(n9689) );
  OR2_X1 U10414 ( .A1(n9689), .A2(n8095), .ZN(n8055) );
  OAI21_X1 U10415 ( .B1(n8052), .B2(P3_IR_REG_17__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8053) );
  XNOR2_X1 U10416 ( .A(n8053), .B(P3_IR_REG_18__SCAN_IN), .ZN(n11887) );
  AOI22_X1 U10417 ( .A1(n11887), .A2(n8072), .B1(SI_18_), .B2(n6650), .ZN(
        n8054) );
  NAND2_X1 U10418 ( .A1(n8055), .A2(n8054), .ZN(n12503) );
  NAND2_X1 U10419 ( .A1(n7929), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8061) );
  NAND2_X1 U10420 ( .A1(n12001), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8060) );
  NAND2_X1 U10421 ( .A1(n8056), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8057) );
  NAND2_X1 U10422 ( .A1(n8057), .A2(n7674), .ZN(n12822) );
  NAND2_X1 U10423 ( .A1(n8170), .A2(n12822), .ZN(n8059) );
  NAND2_X1 U10424 ( .A1(n8171), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8058) );
  OR2_X1 U10425 ( .A1(n12503), .A2(n12800), .ZN(n12125) );
  NAND2_X1 U10426 ( .A1(n12503), .A2(n12800), .ZN(n12136) );
  NAND2_X1 U10427 ( .A1(n12465), .A2(n12849), .ZN(n8062) );
  NAND2_X1 U10428 ( .A1(n13008), .A2(n12833), .ZN(n12827) );
  OR2_X1 U10429 ( .A1(n6644), .A2(n12827), .ZN(n12828) );
  AND2_X1 U10430 ( .A1(n8062), .A2(n12828), .ZN(n12810) );
  AND2_X1 U10431 ( .A1(n12821), .A2(n12810), .ZN(n8063) );
  OR2_X1 U10432 ( .A1(n12503), .A2(n12834), .ZN(n8064) );
  OR2_X1 U10433 ( .A1(n8066), .A2(n8065), .ZN(n8067) );
  NAND2_X1 U10434 ( .A1(n8068), .A2(n8067), .ZN(n9775) );
  NAND2_X1 U10435 ( .A1(n9775), .A2(n11998), .ZN(n8074) );
  OR2_X1 U10436 ( .A1(n6916), .A2(n8069), .ZN(n8071) );
  AOI22_X1 U10437 ( .A1(n6650), .A2(n9774), .B1(n8072), .B2(n12039), .ZN(n8073) );
  NAND2_X1 U10438 ( .A1(n7929), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8079) );
  NAND2_X1 U10439 ( .A1(n12001), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n8078) );
  AND2_X1 U10440 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(n7674), .ZN(n8075) );
  OR2_X1 U10441 ( .A1(n8075), .A2(n8084), .ZN(n12806) );
  NAND2_X1 U10442 ( .A1(n8170), .A2(n12806), .ZN(n8077) );
  NAND2_X1 U10443 ( .A1(n8171), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8076) );
  NAND4_X1 U10444 ( .A1(n8079), .A2(n8078), .A3(n8077), .A4(n8076), .ZN(n12784) );
  NAND2_X1 U10445 ( .A1(n12997), .A2(n12784), .ZN(n12130) );
  NAND2_X1 U10446 ( .A1(n12137), .A2(n12130), .ZN(n12804) );
  NAND2_X1 U10447 ( .A1(n12798), .A2(n12804), .ZN(n12797) );
  INV_X1 U10448 ( .A(n12784), .ZN(n12817) );
  OR2_X1 U10449 ( .A1(n12997), .A2(n12817), .ZN(n8080) );
  XNOR2_X1 U10450 ( .A(n8081), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n10108) );
  NAND2_X1 U10451 ( .A1(n10108), .A2(n11998), .ZN(n8083) );
  INV_X1 U10452 ( .A(SI_20_), .ZN(n10110) );
  OR2_X1 U10453 ( .A1(n11999), .A2(n10110), .ZN(n8082) );
  NAND2_X1 U10454 ( .A1(n7929), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n8089) );
  NAND2_X1 U10455 ( .A1(n12001), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n8088) );
  OR2_X1 U10456 ( .A1(n8084), .A2(n12490), .ZN(n8085) );
  NAND2_X1 U10457 ( .A1(n8098), .A2(n8085), .ZN(n12791) );
  NAND2_X1 U10458 ( .A1(n8170), .A2(n12791), .ZN(n8087) );
  NAND2_X1 U10459 ( .A1(n8171), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8086) );
  NAND2_X1 U10460 ( .A1(n12788), .A2(n12799), .ZN(n12135) );
  NAND2_X1 U10461 ( .A1(n12134), .A2(n12135), .ZN(n12789) );
  NAND2_X1 U10462 ( .A1(n12783), .A2(n12789), .ZN(n12782) );
  NAND2_X1 U10463 ( .A1(n12788), .A2(n12538), .ZN(n8090) );
  NAND2_X1 U10464 ( .A1(n8092), .A2(n8091), .ZN(n8093) );
  NAND2_X1 U10465 ( .A1(n8094), .A2(n8093), .ZN(n10267) );
  OR2_X1 U10466 ( .A1(n10267), .A2(n8095), .ZN(n8097) );
  NAND2_X1 U10467 ( .A1(n6650), .A2(SI_21_), .ZN(n8096) );
  NAND2_X1 U10468 ( .A1(n7929), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8103) );
  NAND2_X1 U10469 ( .A1(n12001), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n8102) );
  NAND2_X1 U10470 ( .A1(n8098), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8099) );
  NAND2_X1 U10471 ( .A1(n8109), .A2(n8099), .ZN(n12777) );
  NAND2_X1 U10472 ( .A1(n8170), .A2(n12777), .ZN(n8101) );
  NAND2_X1 U10473 ( .A1(n12002), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8100) );
  NAND2_X1 U10474 ( .A1(n12989), .A2(n12755), .ZN(n12758) );
  INV_X1 U10475 ( .A(n12755), .ZN(n12785) );
  OR2_X1 U10476 ( .A1(n12989), .A2(n12785), .ZN(n8105) );
  XNOR2_X1 U10477 ( .A(n8107), .B(n8106), .ZN(n14723) );
  NAND2_X1 U10478 ( .A1(n6650), .A2(SI_22_), .ZN(n8108) );
  NAND2_X1 U10479 ( .A1(n12001), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8114) );
  NAND2_X1 U10480 ( .A1(n7929), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8113) );
  AND2_X1 U10481 ( .A1(n8109), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8110) );
  OR2_X1 U10482 ( .A1(n8110), .A2(n8120), .ZN(n12763) );
  NAND2_X1 U10483 ( .A1(n8170), .A2(n12763), .ZN(n8112) );
  NAND2_X1 U10484 ( .A1(n12002), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8111) );
  NAND4_X1 U10485 ( .A1(n8114), .A2(n8113), .A3(n8112), .A4(n8111), .ZN(n12772) );
  NOR2_X1 U10486 ( .A1(n12985), .A2(n12772), .ZN(n8115) );
  INV_X1 U10487 ( .A(n12985), .ZN(n12765) );
  OAI22_X2 U10488 ( .A1(n12753), .A2(n8115), .B1(n12442), .B2(n12765), .ZN(
        n12741) );
  XNOR2_X1 U10489 ( .A(n8117), .B(n8116), .ZN(n10688) );
  NAND2_X1 U10490 ( .A1(n10688), .A2(n11998), .ZN(n8119) );
  NAND2_X1 U10491 ( .A1(n6650), .A2(SI_23_), .ZN(n8118) );
  NAND2_X1 U10492 ( .A1(n12001), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8125) );
  NAND2_X1 U10493 ( .A1(n7929), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8124) );
  NOR2_X1 U10494 ( .A1(n8120), .A2(n12400), .ZN(n8121) );
  OR2_X1 U10495 ( .A1(n8132), .A2(n8121), .ZN(n12746) );
  NAND2_X1 U10496 ( .A1(n8170), .A2(n12746), .ZN(n8123) );
  NAND2_X1 U10497 ( .A1(n12002), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8122) );
  NAND2_X1 U10498 ( .A1(n12749), .A2(n12754), .ZN(n8126) );
  NAND2_X1 U10499 ( .A1(n12153), .A2(n8126), .ZN(n12152) );
  INV_X1 U10500 ( .A(n12754), .ZN(n12728) );
  NAND2_X1 U10501 ( .A1(n12749), .A2(n12728), .ZN(n8127) );
  INV_X1 U10502 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11813) );
  NAND2_X1 U10503 ( .A1(n11107), .A2(n11998), .ZN(n8131) );
  NAND2_X1 U10504 ( .A1(n6650), .A2(SI_24_), .ZN(n8130) );
  NAND2_X1 U10505 ( .A1(n12001), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8137) );
  NAND2_X1 U10506 ( .A1(n8171), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8136) );
  OR2_X1 U10507 ( .A1(n8132), .A2(n12480), .ZN(n8133) );
  NAND2_X1 U10508 ( .A1(n8143), .A2(n8133), .ZN(n12732) );
  NAND2_X1 U10509 ( .A1(n8170), .A2(n12732), .ZN(n8135) );
  NAND2_X1 U10510 ( .A1(n7929), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8134) );
  NAND4_X1 U10511 ( .A1(n8137), .A2(n8136), .A3(n8135), .A4(n8134), .ZN(n12743) );
  AND2_X1 U10512 ( .A1(n12483), .A2(n12743), .ZN(n8138) );
  AOI22_X1 U10513 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(
        P1_DATAO_REG_25__SCAN_IN), .B1(n11471), .B2(n11657), .ZN(n8139) );
  XNOR2_X1 U10514 ( .A(n8140), .B(n8139), .ZN(n11251) );
  NAND2_X1 U10515 ( .A1(n11251), .A2(n11998), .ZN(n8142) );
  NAND2_X1 U10516 ( .A1(n6650), .A2(SI_25_), .ZN(n8141) );
  NAND2_X1 U10517 ( .A1(n7929), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8148) );
  NAND2_X1 U10518 ( .A1(n12001), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8147) );
  NAND2_X1 U10519 ( .A1(n8143), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8144) );
  NAND2_X1 U10520 ( .A1(n8154), .A2(n8144), .ZN(n12716) );
  NAND2_X1 U10521 ( .A1(n8170), .A2(n12716), .ZN(n8146) );
  NAND2_X1 U10522 ( .A1(n12002), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8145) );
  NAND4_X1 U10523 ( .A1(n8148), .A2(n8147), .A3(n8146), .A4(n8145), .ZN(n12727) );
  XNOR2_X1 U10524 ( .A(n12454), .B(n12727), .ZN(n12708) );
  INV_X1 U10525 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14695) );
  AOI22_X1 U10526 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n13853), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n14695), .ZN(n8149) );
  INV_X1 U10527 ( .A(n8149), .ZN(n8150) );
  XNOR2_X1 U10528 ( .A(n8151), .B(n8150), .ZN(n11303) );
  NAND2_X1 U10529 ( .A1(n11303), .A2(n11998), .ZN(n8153) );
  NAND2_X1 U10530 ( .A1(n6650), .A2(SI_26_), .ZN(n8152) );
  NAND2_X1 U10531 ( .A1(n12001), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8159) );
  NAND2_X1 U10532 ( .A1(n7929), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8158) );
  AND2_X1 U10533 ( .A1(n8154), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8155) );
  OR2_X1 U10534 ( .A1(n8155), .A2(n8167), .ZN(n12702) );
  NAND2_X1 U10535 ( .A1(n8186), .A2(n12702), .ZN(n8157) );
  NAND2_X1 U10536 ( .A1(n12002), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8156) );
  NAND4_X1 U10537 ( .A1(n8159), .A2(n8158), .A3(n8157), .A4(n8156), .ZN(n12712) );
  OR2_X1 U10538 ( .A1(n12898), .A2(n12712), .ZN(n8160) );
  NAND2_X1 U10539 ( .A1(n12696), .A2(n8160), .ZN(n8162) );
  NAND2_X1 U10540 ( .A1(n12898), .A2(n12712), .ZN(n8161) );
  XNOR2_X1 U10541 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n8163) );
  XNOR2_X1 U10542 ( .A(n8164), .B(n8163), .ZN(n11491) );
  NAND2_X1 U10543 ( .A1(n11491), .A2(n11998), .ZN(n8166) );
  NAND2_X1 U10544 ( .A1(n6650), .A2(SI_27_), .ZN(n8165) );
  NAND2_X1 U10545 ( .A1(n7929), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8175) );
  NAND2_X1 U10546 ( .A1(n12001), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8174) );
  NOR2_X1 U10547 ( .A1(n8167), .A2(n12393), .ZN(n8168) );
  NAND2_X1 U10548 ( .A1(n8170), .A2(n12688), .ZN(n8173) );
  NAND2_X1 U10549 ( .A1(n8171), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8172) );
  OR2_X1 U10550 ( .A1(n12699), .A2(n6864), .ZN(n8177) );
  NAND2_X1 U10551 ( .A1(n12671), .A2(n12683), .ZN(n8228) );
  AOI21_X1 U10552 ( .B1(n12537), .B2(n12671), .A(n12664), .ZN(n8190) );
  INV_X1 U10553 ( .A(n8178), .ZN(n8180) );
  INV_X1 U10554 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n11810) );
  NAND2_X1 U10555 ( .A1(n11810), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8179) );
  NAND2_X1 U10556 ( .A1(n8180), .A2(n8179), .ZN(n8182) );
  NAND2_X1 U10557 ( .A1(n8998), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8181) );
  NAND2_X1 U10558 ( .A1(n8182), .A2(n8181), .ZN(n11983) );
  XNOR2_X1 U10559 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n11981) );
  XNOR2_X1 U10560 ( .A(n11983), .B(n11981), .ZN(n13026) );
  NAND2_X1 U10561 ( .A1(n13026), .A2(n11998), .ZN(n8184) );
  NAND2_X1 U10562 ( .A1(n6650), .A2(SI_29_), .ZN(n8183) );
  INV_X1 U10563 ( .A(n12657), .ZN(n8185) );
  NAND2_X1 U10564 ( .A1(n8186), .A2(n8185), .ZN(n12006) );
  NAND2_X1 U10565 ( .A1(n12001), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8189) );
  NAND2_X1 U10566 ( .A1(n12002), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8188) );
  NAND2_X1 U10567 ( .A1(n7929), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8187) );
  NAND2_X1 U10568 ( .A1(n12205), .A2(n12536), .ZN(n12174) );
  NAND2_X1 U10569 ( .A1(n12176), .A2(n12174), .ZN(n12038) );
  XNOR2_X1 U10570 ( .A(n8190), .B(n12038), .ZN(n8205) );
  OAI21_X1 U10571 ( .B1(n8237), .B2(P3_IR_REG_21__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8192) );
  OR2_X1 U10572 ( .A1(n14725), .A2(n12039), .ZN(n8284) );
  NAND2_X1 U10573 ( .A1(n8237), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8194) );
  INV_X1 U10574 ( .A(n12049), .ZN(n12044) );
  NAND2_X1 U10575 ( .A1(n8195), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8196) );
  MUX2_X1 U10576 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8196), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n8197) );
  NAND2_X1 U10577 ( .A1(n12044), .A2(n8283), .ZN(n12186) );
  NAND2_X1 U10578 ( .A1(n7929), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8200) );
  NAND2_X1 U10579 ( .A1(n12001), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8199) );
  NAND2_X1 U10580 ( .A1(n12002), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8198) );
  AND4_X1 U10581 ( .A1(n12006), .A2(n8200), .A3(n8199), .A4(n8198), .ZN(n12007) );
  INV_X1 U10582 ( .A(n8201), .ZN(n10128) );
  NAND2_X1 U10583 ( .A1(n10128), .A2(n12187), .ZN(n10143) );
  NAND2_X1 U10584 ( .A1(n10143), .A2(n10127), .ZN(n10014) );
  INV_X1 U10585 ( .A(P3_B_REG_SCAN_IN), .ZN(n8202) );
  NOR2_X1 U10586 ( .A1(n8201), .A2(n8202), .ZN(n8203) );
  OR2_X1 U10587 ( .A1(n15448), .A2(n8203), .ZN(n12655) );
  INV_X1 U10588 ( .A(n10014), .ZN(n10017) );
  OAI22_X1 U10589 ( .A1(n12007), .A2(n12655), .B1(n12683), .B2(n15450), .ZN(
        n8204) );
  AOI21_X2 U10590 ( .B1(n8205), .B2(n15466), .A(n8204), .ZN(n12206) );
  NAND2_X1 U10591 ( .A1(n10001), .A2(n12050), .ZN(n15441) );
  NAND2_X1 U10592 ( .A1(n15441), .A2(n15446), .ZN(n15440) );
  NAND2_X1 U10593 ( .A1(n10482), .A2(n9995), .ZN(n12056) );
  NAND2_X1 U10594 ( .A1(n10480), .A2(n12019), .ZN(n8207) );
  INV_X1 U10595 ( .A(n12061), .ZN(n12020) );
  NAND2_X1 U10596 ( .A1(n10375), .A2(n12020), .ZN(n8209) );
  INV_X1 U10597 ( .A(n12548), .ZN(n12063) );
  NAND2_X1 U10598 ( .A1(n12063), .A2(n10280), .ZN(n8208) );
  NAND2_X1 U10599 ( .A1(n10974), .A2(n12025), .ZN(n8210) );
  INV_X1 U10600 ( .A(n12022), .ZN(n12077) );
  INV_X1 U10601 ( .A(n12021), .ZN(n12083) );
  NAND2_X1 U10602 ( .A1(n11213), .A2(n12083), .ZN(n8211) );
  NOR2_X1 U10603 ( .A1(n12544), .A2(n11310), .ZN(n12092) );
  NAND2_X1 U10604 ( .A1(n12544), .A2(n11310), .ZN(n12090) );
  XNOR2_X1 U10605 ( .A(n12542), .B(n12103), .ZN(n12106) );
  NAND2_X1 U10606 ( .A1(n11445), .A2(n12106), .ZN(n11444) );
  NAND2_X1 U10607 ( .A1(n14777), .A2(n12103), .ZN(n12095) );
  INV_X1 U10608 ( .A(n14774), .ZN(n14768) );
  NAND2_X1 U10609 ( .A1(n14769), .A2(n14768), .ZN(n8214) );
  INV_X1 U10610 ( .A(n12113), .ZN(n8215) );
  NAND2_X1 U10611 ( .A1(n12884), .A2(n14763), .ZN(n8218) );
  NAND2_X1 U10612 ( .A1(n13015), .A2(n12848), .ZN(n12041) );
  NAND2_X1 U10613 ( .A1(n12360), .A2(n12879), .ZN(n12120) );
  NAND2_X1 U10614 ( .A1(n12864), .A2(n12863), .ZN(n12862) );
  AND2_X1 U10615 ( .A1(n12837), .A2(n12128), .ZN(n12818) );
  AND2_X1 U10616 ( .A1(n12818), .A2(n12814), .ZN(n8221) );
  OR2_X1 U10617 ( .A1(n12821), .A2(n12819), .ZN(n8219) );
  NAND2_X1 U10618 ( .A1(n12985), .A2(n12442), .ZN(n12016) );
  AND2_X1 U10619 ( .A1(n12758), .A2(n12016), .ZN(n8223) );
  INV_X1 U10620 ( .A(n12016), .ZN(n12150) );
  AND2_X1 U10621 ( .A1(n8224), .A2(n12148), .ZN(n8225) );
  XNOR2_X1 U10622 ( .A(n12483), .B(n12476), .ZN(n12725) );
  NAND2_X1 U10623 ( .A1(n12483), .A2(n12476), .ZN(n12155) );
  NAND2_X1 U10624 ( .A1(n12709), .A2(n12708), .ZN(n12694) );
  INV_X1 U10625 ( .A(n12727), .ZN(n12513) );
  NAND2_X1 U10626 ( .A1(n12454), .A2(n12513), .ZN(n12693) );
  NAND2_X1 U10627 ( .A1(n12898), .A2(n12684), .ZN(n12163) );
  AND2_X1 U10628 ( .A1(n12693), .A2(n12163), .ZN(n8227) );
  INV_X1 U10629 ( .A(n12162), .ZN(n8226) );
  INV_X1 U10630 ( .A(n12699), .ZN(n12514) );
  NAND2_X1 U10631 ( .A1(n6864), .A2(n12514), .ZN(n12668) );
  AND2_X1 U10632 ( .A1(n8228), .A2(n12668), .ZN(n12167) );
  INV_X1 U10633 ( .A(n8229), .ZN(n12166) );
  XNOR2_X1 U10634 ( .A(n12012), .B(n12038), .ZN(n12203) );
  OAI21_X1 U10635 ( .B1(n14725), .B2(n8283), .A(n12014), .ZN(n8230) );
  NAND2_X1 U10636 ( .A1(n8230), .A2(n12049), .ZN(n8232) );
  OAI21_X1 U10637 ( .B1(n8283), .B2(n12044), .A(n14725), .ZN(n8231) );
  NAND2_X1 U10638 ( .A1(n8232), .A2(n8231), .ZN(n10006) );
  NAND2_X1 U10639 ( .A1(n10109), .A2(n12039), .ZN(n8282) );
  INV_X1 U10640 ( .A(n8282), .ZN(n12182) );
  AND2_X1 U10641 ( .A1(n15521), .A2(n12182), .ZN(n8233) );
  NAND2_X1 U10642 ( .A1(n10006), .A2(n8233), .ZN(n8235) );
  NAND2_X1 U10643 ( .A1(n8283), .A2(n12039), .ZN(n8234) );
  OR2_X1 U10644 ( .A1(n8234), .A2(n14725), .ZN(n8270) );
  NAND2_X1 U10645 ( .A1(n14725), .A2(n15444), .ZN(n15522) );
  NAND2_X1 U10646 ( .A1(n8265), .A2(n13256), .ZN(n8239) );
  NAND2_X1 U10647 ( .A1(n8239), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8238) );
  MUX2_X1 U10648 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8238), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8240) );
  OR2_X2 U10649 ( .A1(n8239), .A2(P3_IR_REG_24__SCAN_IN), .ZN(n8244) );
  XNOR2_X1 U10650 ( .A(n11110), .B(P3_B_REG_SCAN_IN), .ZN(n8243) );
  NAND2_X1 U10651 ( .A1(n8243), .A2(n11254), .ZN(n8246) );
  INV_X1 U10652 ( .A(n8263), .ZN(n11306) );
  NAND2_X1 U10653 ( .A1(n11306), .A2(n11110), .ZN(n8247) );
  NAND2_X1 U10654 ( .A1(n11306), .A2(n11254), .ZN(n8248) );
  NAND2_X1 U10655 ( .A1(n13018), .A2(n13016), .ZN(n8281) );
  NOR2_X1 U10656 ( .A1(P3_D_REG_25__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .ZN(
        n8253) );
  NOR4_X1 U10657 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_2__SCAN_IN), .A4(P3_D_REG_10__SCAN_IN), .ZN(n8252) );
  NOR4_X1 U10658 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n8251) );
  NOR4_X1 U10659 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_17__SCAN_IN), .A3(
        P3_D_REG_22__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n8250) );
  NAND4_X1 U10660 ( .A1(n8253), .A2(n8252), .A3(n8251), .A4(n8250), .ZN(n8259)
         );
  NOR4_X1 U10661 ( .A1(P3_D_REG_12__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n8257) );
  NOR4_X1 U10662 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_21__SCAN_IN), .ZN(n8256) );
  NOR4_X1 U10663 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8255) );
  NOR4_X1 U10664 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n8254) );
  NAND4_X1 U10665 ( .A1(n8257), .A2(n8256), .A3(n8255), .A4(n8254), .ZN(n8258)
         );
  NOR2_X1 U10666 ( .A1(n8259), .A2(n8258), .ZN(n8260) );
  INV_X1 U10667 ( .A(n11254), .ZN(n8262) );
  INV_X1 U10668 ( .A(n11110), .ZN(n8261) );
  INV_X1 U10669 ( .A(n8265), .ZN(n8266) );
  AND2_X1 U10670 ( .A1(n8280), .A2(n10124), .ZN(n8269) );
  INV_X1 U10671 ( .A(n13018), .ZN(n8268) );
  INV_X1 U10672 ( .A(n13016), .ZN(n8275) );
  NAND2_X1 U10673 ( .A1(n8268), .A2(n8275), .ZN(n8288) );
  NAND2_X1 U10674 ( .A1(n12171), .A2(n8282), .ZN(n9983) );
  NAND2_X1 U10675 ( .A1(n8270), .A2(n12161), .ZN(n9858) );
  AND2_X1 U10676 ( .A1(n9983), .A2(n9858), .ZN(n9860) );
  OAI22_X1 U10677 ( .A1(n15521), .A2(n8283), .B1(n12014), .B2(n14725), .ZN(
        n8271) );
  NAND2_X1 U10678 ( .A1(n8271), .A2(n8282), .ZN(n8272) );
  NAND2_X1 U10679 ( .A1(n8272), .A2(n12161), .ZN(n8273) );
  NAND2_X1 U10680 ( .A1(n8275), .A2(n8273), .ZN(n8274) );
  OAI21_X1 U10681 ( .B1(n8275), .B2(n9860), .A(n8274), .ZN(n8276) );
  INV_X1 U10682 ( .A(n8276), .ZN(n8277) );
  NAND2_X1 U10683 ( .A1(n15544), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8278) );
  INV_X1 U10684 ( .A(n15521), .ZN(n15488) );
  NAND2_X1 U10685 ( .A1(n12205), .A2(n12951), .ZN(n8279) );
  NOR2_X1 U10686 ( .A1(n12161), .A2(n8282), .ZN(n9865) );
  NAND2_X1 U10687 ( .A1(n10124), .A2(n9865), .ZN(n12188) );
  NAND2_X1 U10688 ( .A1(n12049), .A2(n8283), .ZN(n9992) );
  NOR2_X1 U10689 ( .A1(n8284), .A2(n9992), .ZN(n10007) );
  NAND2_X1 U10690 ( .A1(n10124), .A2(n10007), .ZN(n8285) );
  NAND2_X1 U10691 ( .A1(n12188), .A2(n8285), .ZN(n8286) );
  NAND2_X1 U10692 ( .A1(n10015), .A2(n8286), .ZN(n8290) );
  NAND3_X1 U10693 ( .A1(n10013), .A2(n10124), .A3(n10006), .ZN(n8289) );
  NAND2_X1 U10694 ( .A1(n15526), .A2(n8291), .ZN(n8292) );
  INV_X1 U10695 ( .A(n13014), .ZN(n13009) );
  NAND2_X1 U10696 ( .A1(n12205), .A2(n13009), .ZN(n8294) );
  INV_X1 U10697 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n15071) );
  INV_X1 U10698 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n12590) );
  INV_X1 U10699 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15056) );
  XOR2_X1 U10700 ( .A(n15056), .B(P3_ADDR_REG_15__SCAN_IN), .Z(n8335) );
  INV_X1 U10701 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n8324) );
  XOR2_X1 U10702 ( .A(n8324), .B(P1_ADDR_REG_14__SCAN_IN), .Z(n8382) );
  INV_X1 U10703 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n8322) );
  INV_X1 U10704 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n15026) );
  XOR2_X1 U10705 ( .A(n15026), .B(P3_ADDR_REG_13__SCAN_IN), .Z(n8377) );
  XOR2_X1 U10706 ( .A(n11280), .B(P1_ADDR_REG_12__SCAN_IN), .Z(n8337) );
  INV_X1 U10707 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n8319) );
  XOR2_X1 U10708 ( .A(n8319), .B(P1_ADDR_REG_11__SCAN_IN), .Z(n8373) );
  INV_X1 U10709 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9764) );
  XNOR2_X1 U10710 ( .A(n8314), .B(n9764), .ZN(n8340) );
  INV_X1 U10711 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n8312) );
  XOR2_X1 U10712 ( .A(n8312), .B(P1_ADDR_REG_8__SCAN_IN), .Z(n8342) );
  XNOR2_X1 U10713 ( .A(n9886), .B(n13266), .ZN(n8362) );
  XOR2_X1 U10714 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n8298), .Z(n8347) );
  INV_X1 U10715 ( .A(n8350), .ZN(n8296) );
  NAND2_X1 U10716 ( .A1(n8296), .A2(n8349), .ZN(n8297) );
  NAND2_X1 U10717 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n8299), .ZN(n8301) );
  NAND2_X1 U10718 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n8302), .ZN(n8303) );
  NAND2_X1 U10719 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n8304), .ZN(n8306) );
  NAND2_X1 U10720 ( .A1(n8344), .A2(n9751), .ZN(n8305) );
  NAND2_X1 U10721 ( .A1(n8306), .A2(n8305), .ZN(n8363) );
  NAND2_X1 U10722 ( .A1(n8362), .A2(n8363), .ZN(n8307) );
  NAND2_X1 U10723 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n8308), .ZN(n8310) );
  XOR2_X1 U10724 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n8308), .Z(n8368) );
  INV_X1 U10725 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9897) );
  NAND2_X1 U10726 ( .A1(n8368), .A2(n9897), .ZN(n8309) );
  NAND2_X1 U10727 ( .A1(n8310), .A2(n8309), .ZN(n8343) );
  NAND2_X1 U10728 ( .A1(n8342), .A2(n8343), .ZN(n8311) );
  NAND2_X1 U10729 ( .A1(n8340), .A2(n8341), .ZN(n8313) );
  NAND2_X1 U10730 ( .A1(n9911), .A2(n8315), .ZN(n8317) );
  XOR2_X1 U10731 ( .A(n9911), .B(n8315), .Z(n8339) );
  NAND2_X1 U10732 ( .A1(P3_ADDR_REG_10__SCAN_IN), .A2(n8339), .ZN(n8316) );
  NAND2_X1 U10733 ( .A1(n8317), .A2(n8316), .ZN(n8374) );
  NAND2_X1 U10734 ( .A1(n8373), .A2(n8374), .ZN(n8318) );
  NAND2_X1 U10735 ( .A1(n8337), .A2(n8338), .ZN(n8320) );
  NAND2_X1 U10736 ( .A1(n8377), .A2(n8378), .ZN(n8321) );
  NAND2_X1 U10737 ( .A1(n8382), .A2(n8383), .ZN(n8323) );
  NAND2_X1 U10738 ( .A1(n8335), .A2(n8336), .ZN(n8325) );
  NOR2_X1 U10739 ( .A1(n15071), .A2(n8326), .ZN(n8328) );
  XOR2_X1 U10740 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n8326), .Z(n8334) );
  NOR2_X1 U10741 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n8334), .ZN(n8327) );
  NOR2_X1 U10742 ( .A1(n8328), .A2(n8327), .ZN(n8329) );
  INV_X1 U10743 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n15086) );
  NAND2_X1 U10744 ( .A1(n8329), .A2(n15086), .ZN(n8331) );
  XNOR2_X1 U10745 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n8329), .ZN(n8333) );
  NAND2_X1 U10746 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n8333), .ZN(n8330) );
  NAND2_X1 U10747 ( .A1(n8331), .A2(n8330), .ZN(n8394) );
  INV_X1 U10748 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n8397) );
  NOR2_X1 U10749 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n8397), .ZN(n8332) );
  AOI21_X1 U10750 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n8397), .A(n8332), .ZN(
        n8395) );
  XOR2_X1 U10751 ( .A(n8394), .B(n8395), .Z(n14703) );
  XOR2_X1 U10752 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n8333), .Z(n14756) );
  INV_X1 U10753 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n13153) );
  XOR2_X1 U10754 ( .A(n13153), .B(n8334), .Z(n15000) );
  XOR2_X1 U10755 ( .A(n8336), .B(n8335), .Z(n8388) );
  XNOR2_X1 U10756 ( .A(n8338), .B(n8337), .ZN(n8375) );
  XOR2_X1 U10757 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(n8339), .Z(n14728) );
  XOR2_X1 U10758 ( .A(n8341), .B(n8340), .Z(n14719) );
  XOR2_X1 U10759 ( .A(n8343), .B(n8342), .Z(n14715) );
  XNOR2_X1 U10760 ( .A(n8345), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n8357) );
  INV_X1 U10761 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n8356) );
  NAND2_X1 U10762 ( .A1(n8357), .A2(n8356), .ZN(n8358) );
  XOR2_X1 U10763 ( .A(n8346), .B(n14310), .Z(n15560) );
  XOR2_X1 U10764 ( .A(n8348), .B(n8347), .Z(n14708) );
  NOR2_X1 U10765 ( .A1(n8352), .A2(n6836), .ZN(n8353) );
  OAI21_X1 U10766 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n8351), .A(n8350), .ZN(
        n15554) );
  NAND2_X1 U10767 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15554), .ZN(n15564) );
  NOR2_X1 U10768 ( .A1(n15564), .A2(n15563), .ZN(n15562) );
  NOR2_X1 U10769 ( .A1(n14708), .A2(n14707), .ZN(n8354) );
  NAND2_X1 U10770 ( .A1(n14708), .A2(n14707), .ZN(n14706) );
  NAND2_X1 U10771 ( .A1(n15560), .A2(n15559), .ZN(n8355) );
  NOR2_X1 U10772 ( .A1(n15560), .A2(n15559), .ZN(n15558) );
  XNOR2_X1 U10773 ( .A(n8357), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n15549) );
  NAND2_X1 U10774 ( .A1(n15550), .A2(n15549), .ZN(n15548) );
  NAND2_X1 U10775 ( .A1(n8358), .A2(n15548), .ZN(n8360) );
  NAND2_X1 U10776 ( .A1(n8359), .A2(n8360), .ZN(n8361) );
  INV_X1 U10777 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15552) );
  NOR2_X1 U10778 ( .A1(n8364), .A2(n7277), .ZN(n8365) );
  XOR2_X1 U10779 ( .A(n8363), .B(n8362), .Z(n14712) );
  INV_X1 U10780 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n8366) );
  NAND2_X1 U10781 ( .A1(n8367), .A2(n8366), .ZN(n8369) );
  XOR2_X1 U10782 ( .A(n8368), .B(n9897), .Z(n15556) );
  NAND2_X1 U10783 ( .A1(n15557), .A2(n15556), .ZN(n15555) );
  NAND2_X1 U10784 ( .A1(n14715), .A2(n14714), .ZN(n8370) );
  AOI21_X2 U10785 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(n8370), .A(n14713), .ZN(
        n14718) );
  NAND2_X1 U10786 ( .A1(n14719), .A2(n14718), .ZN(n8371) );
  NAND2_X1 U10787 ( .A1(n14728), .A2(n14727), .ZN(n8372) );
  XOR2_X1 U10788 ( .A(n8374), .B(n8373), .Z(n14982) );
  INV_X1 U10789 ( .A(n14986), .ZN(n14987) );
  INV_X1 U10790 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15251) );
  NAND2_X1 U10791 ( .A1(n8376), .A2(n8375), .ZN(n14988) );
  XOR2_X1 U10792 ( .A(n8378), .B(n8377), .Z(n8380) );
  INV_X1 U10793 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14990) );
  NAND2_X1 U10794 ( .A1(n8380), .A2(n8379), .ZN(n8381) );
  XOR2_X1 U10795 ( .A(n8383), .B(n8382), .Z(n8386) );
  INV_X1 U10796 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14993) );
  NAND2_X1 U10797 ( .A1(n14994), .A2(n14993), .ZN(n14992) );
  NAND2_X1 U10798 ( .A1(n8386), .A2(n8385), .ZN(n8387) );
  NAND2_X1 U10799 ( .A1(n8388), .A2(n8390), .ZN(n8391) );
  INV_X1 U10800 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n14996) );
  NAND2_X1 U10801 ( .A1(n15000), .A2(n14999), .ZN(n8392) );
  NAND2_X1 U10802 ( .A1(n14703), .A2(n14702), .ZN(n8393) );
  NAND2_X1 U10803 ( .A1(n8395), .A2(n8394), .ZN(n8396) );
  OAI21_X1 U10804 ( .B1(n8397), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n8396), .ZN(
        n8398) );
  XOR2_X1 U10805 ( .A(n8398), .B(P3_ADDR_REG_19__SCAN_IN), .Z(n8400) );
  XNOR2_X1 U10806 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n8399) );
  XNOR2_X1 U10807 ( .A(n8400), .B(n8399), .ZN(n8401) );
  NOR2_X1 U10808 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n8407) );
  NAND2_X1 U10809 ( .A1(n8723), .A2(n8409), .ZN(n8770) );
  NAND2_X1 U10810 ( .A1(n8791), .A2(n8410), .ZN(n8811) );
  INV_X1 U10811 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8415) );
  INV_X1 U10812 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8417) );
  XNOR2_X1 U10813 ( .A(n8417), .B(P2_IR_REG_31__SCAN_IN), .ZN(n8418) );
  NAND2_X1 U10814 ( .A1(n8422), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8423) );
  MUX2_X1 U10815 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8423), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n8424) );
  NAND2_X1 U10816 ( .A1(n8427), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8428) );
  NAND2_X4 U10817 ( .A1(n9570), .A2(n6637), .ZN(n9121) );
  NOR2_X1 U10818 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), 
        .ZN(n8432) );
  NOR2_X1 U10819 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), 
        .ZN(n8436) );
  NOR2_X1 U10820 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), 
        .ZN(n8435) );
  NAND2_X1 U10821 ( .A1(n9115), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8447) );
  NAND2_X1 U10822 ( .A1(n9096), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8446) );
  NAND2_X1 U10823 ( .A1(n8497), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8445) );
  AND2_X2 U10824 ( .A1(n11908), .A2(n13844), .ZN(n8481) );
  NAND2_X1 U10825 ( .A1(n8481), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8444) );
  NAND4_X1 U10826 ( .A1(n8447), .A2(n8446), .A3(n8445), .A4(n8444), .ZN(n8463)
         );
  NAND2_X1 U10827 ( .A1(n8991), .A2(SI_0_), .ZN(n8449) );
  XNOR2_X1 U10828 ( .A(n8449), .B(n6941), .ZN(n13856) );
  NAND2_X1 U10829 ( .A1(n8456), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8457) );
  MUX2_X2 U10830 ( .A(n7649), .B(n13856), .S(n8533), .Z(n15307) );
  AND2_X1 U10831 ( .A1(n8463), .A2(n15307), .ZN(n9161) );
  INV_X1 U10832 ( .A(n10184), .ZN(n9572) );
  NAND2_X1 U10833 ( .A1(n9121), .A2(n9614), .ZN(n8461) );
  NAND2_X1 U10834 ( .A1(n8462), .A2(n8461), .ZN(n8465) );
  OAI211_X1 U10835 ( .C1(n10184), .C2(n15307), .A(n9121), .B(n8463), .ZN(n8464) );
  NAND2_X1 U10836 ( .A1(n8465), .A2(n8464), .ZN(n8480) );
  NAND2_X1 U10837 ( .A1(n8481), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8469) );
  NAND2_X1 U10838 ( .A1(n9096), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n8468) );
  NAND2_X1 U10839 ( .A1(n9115), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8467) );
  NAND2_X1 U10840 ( .A1(n8497), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8466) );
  NAND2_X1 U10842 ( .A1(n8574), .A2(n13533), .ZN(n8476) );
  NAND2_X1 U10843 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8470) );
  MUX2_X1 U10844 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8470), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n8471) );
  NAND2_X1 U10845 ( .A1(n8471), .A2(n6673), .ZN(n15203) );
  OR2_X1 U10846 ( .A1(n8502), .A2(n9349), .ZN(n8474) );
  NAND2_X1 U10847 ( .A1(n8472), .A2(SI_1_), .ZN(n8488) );
  XNOR2_X1 U10848 ( .A(n8489), .B(n8490), .ZN(n9801) );
  NAND2_X1 U10849 ( .A1(n9121), .A2(n9645), .ZN(n8475) );
  NAND2_X1 U10850 ( .A1(n9121), .A2(n13533), .ZN(n8477) );
  OAI21_X1 U10851 ( .B1(n9121), .B2(n9568), .A(n8477), .ZN(n8478) );
  NAND2_X1 U10852 ( .A1(n9096), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n8485) );
  NAND2_X1 U10853 ( .A1(n9115), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8484) );
  NAND2_X1 U10854 ( .A1(n8497), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8483) );
  NAND2_X1 U10855 ( .A1(n8481), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8482) );
  NAND2_X1 U10856 ( .A1(n9121), .A2(n13532), .ZN(n8494) );
  NAND2_X1 U10857 ( .A1(n6673), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8487) );
  XNOR2_X1 U10858 ( .A(n8487), .B(n8486), .ZN(n13538) );
  INV_X1 U10859 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n11620) );
  MUX2_X1 U10860 ( .A(n11620), .B(n9337), .S(n11734), .Z(n8521) );
  XNOR2_X1 U10861 ( .A(n8521), .B(n8507), .ZN(n9336) );
  OR2_X1 U10862 ( .A1(n8502), .A2(n9337), .ZN(n8491) );
  NAND2_X1 U10863 ( .A1(n8494), .A2(n8493), .ZN(n8496) );
  AOI22_X1 U10864 ( .A1(n9143), .A2(n13532), .B1(n9121), .B2(n10200), .ZN(
        n8495) );
  INV_X1 U10865 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10352) );
  NAND2_X1 U10866 ( .A1(n9096), .A2(n10352), .ZN(n8501) );
  NAND2_X1 U10867 ( .A1(n9115), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n8500) );
  NAND2_X1 U10868 ( .A1(n8497), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8499) );
  NAND2_X1 U10869 ( .A1(n8481), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8498) );
  INV_X1 U10870 ( .A(n13531), .ZN(n10204) );
  OR2_X1 U10871 ( .A1(n9121), .A2(n10204), .ZN(n8513) );
  INV_X2 U10872 ( .A(n8502), .ZN(n8862) );
  NAND2_X1 U10873 ( .A1(n8503), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8504) );
  MUX2_X1 U10874 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8504), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n8506) );
  AND2_X1 U10875 ( .A1(n8506), .A2(n8505), .ZN(n9496) );
  INV_X4 U10876 ( .A(n9109), .ZN(n9092) );
  NAND2_X1 U10877 ( .A1(n9344), .A2(n9092), .ZN(n8510) );
  NAND2_X1 U10878 ( .A1(n9113), .A2(n10359), .ZN(n8512) );
  NAND2_X1 U10879 ( .A1(n8513), .A2(n8512), .ZN(n8517) );
  NAND2_X1 U10880 ( .A1(n8518), .A2(n8517), .ZN(n8516) );
  AOI22_X1 U10881 ( .A1(n9102), .A2(n10359), .B1(n9113), .B2(n13531), .ZN(
        n8514) );
  NAND2_X1 U10882 ( .A1(n8505), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8520) );
  INV_X1 U10883 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8519) );
  XNOR2_X1 U10884 ( .A(n8520), .B(n8519), .ZN(n9434) );
  INV_X1 U10885 ( .A(SI_2_), .ZN(n9329) );
  NOR2_X1 U10886 ( .A1(n8521), .A2(n9329), .ZN(n8526) );
  INV_X1 U10887 ( .A(n8521), .ZN(n8522) );
  NOR2_X1 U10888 ( .A1(n8522), .A2(SI_2_), .ZN(n8523) );
  MUX2_X1 U10889 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n11734), .Z(n8529) );
  NAND2_X1 U10890 ( .A1(n8529), .A2(SI_4_), .ZN(n8553) );
  OAI21_X1 U10891 ( .B1(n8529), .B2(SI_4_), .A(n8553), .ZN(n8530) );
  INV_X1 U10892 ( .A(n8530), .ZN(n8551) );
  XNOR2_X1 U10893 ( .A(n8552), .B(n8551), .ZN(n9959) );
  OR2_X1 U10894 ( .A1(n9959), .A2(n9109), .ZN(n8532) );
  OR2_X1 U10895 ( .A1(n9110), .A2(n9327), .ZN(n8531) );
  OAI211_X1 U10896 ( .C1(n8533), .C2(n9434), .A(n8532), .B(n8531), .ZN(n15324)
         );
  INV_X1 U10897 ( .A(n15324), .ZN(n10229) );
  OR2_X1 U10898 ( .A1(n9121), .A2(n10229), .ZN(n8540) );
  NAND2_X1 U10899 ( .A1(n8481), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8538) );
  NAND2_X1 U10900 ( .A1(n9115), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n8537) );
  INV_X1 U10901 ( .A(n8543), .ZN(n8545) );
  OAI21_X1 U10902 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n8545), .ZN(n10228) );
  INV_X1 U10903 ( .A(n10228), .ZN(n8534) );
  NAND2_X1 U10904 ( .A1(n9096), .A2(n8534), .ZN(n8536) );
  NAND2_X1 U10905 ( .A1(n8497), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8535) );
  NAND4_X1 U10906 ( .A1(n8538), .A2(n8537), .A3(n8536), .A4(n8535), .ZN(n13530) );
  NAND2_X1 U10907 ( .A1(n9113), .A2(n13530), .ZN(n8539) );
  NAND2_X1 U10908 ( .A1(n8540), .A2(n8539), .ZN(n8542) );
  AOI22_X1 U10909 ( .A1(n9143), .A2(n13530), .B1(n9113), .B2(n15324), .ZN(
        n8541) );
  NAND2_X1 U10910 ( .A1(n9035), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8550) );
  NAND2_X1 U10911 ( .A1(n6860), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8549) );
  NAND2_X1 U10912 ( .A1(n8543), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8594) );
  INV_X1 U10913 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8544) );
  NAND2_X1 U10914 ( .A1(n8545), .A2(n8544), .ZN(n8546) );
  AND2_X1 U10915 ( .A1(n8594), .A2(n8546), .ZN(n10195) );
  NAND2_X1 U10916 ( .A1(n6652), .A2(n10195), .ZN(n8548) );
  NAND2_X1 U10917 ( .A1(n6651), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8547) );
  NAND4_X1 U10918 ( .A1(n8550), .A2(n8549), .A3(n8548), .A4(n8547), .ZN(n13529) );
  INV_X1 U10919 ( .A(n13529), .ZN(n10238) );
  OR2_X1 U10920 ( .A1(n9121), .A2(n10238), .ZN(n8560) );
  NAND2_X1 U10921 ( .A1(n8554), .A2(SI_5_), .ZN(n8566) );
  OAI21_X1 U10922 ( .B1(n8554), .B2(SI_5_), .A(n8566), .ZN(n8563) );
  XNOR2_X1 U10923 ( .A(n8565), .B(n8563), .ZN(n9341) );
  NAND2_X1 U10924 ( .A1(n9341), .A2(n9092), .ZN(n8558) );
  INV_X1 U10925 ( .A(n8555), .ZN(n8698) );
  NAND2_X1 U10926 ( .A1(n8698), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8556) );
  XNOR2_X1 U10927 ( .A(n8556), .B(P2_IR_REG_5__SCAN_IN), .ZN(n9519) );
  AOI22_X1 U10928 ( .A1(n8862), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6643), .B2(
        n9519), .ZN(n8557) );
  NAND2_X1 U10929 ( .A1(n8558), .A2(n8557), .ZN(n10239) );
  NAND2_X1 U10930 ( .A1(n9113), .A2(n10239), .ZN(n8559) );
  NAND2_X1 U10931 ( .A1(n8560), .A2(n8559), .ZN(n8562) );
  AOI22_X1 U10932 ( .A1(n9102), .A2(n10239), .B1(n9113), .B2(n13529), .ZN(
        n8561) );
  INV_X1 U10933 ( .A(n8563), .ZN(n8564) );
  MUX2_X1 U10934 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n11734), .Z(n8567) );
  NAND2_X1 U10935 ( .A1(n8567), .A2(SI_6_), .ZN(n8586) );
  OAI21_X1 U10936 ( .B1(n8567), .B2(SI_6_), .A(n8586), .ZN(n8584) );
  XNOR2_X1 U10937 ( .A(n8585), .B(n8584), .ZN(n10551) );
  NAND2_X1 U10938 ( .A1(n10551), .A2(n9092), .ZN(n8573) );
  AND2_X1 U10939 ( .A1(n8609), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8568) );
  NAND2_X1 U10940 ( .A1(n8568), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n8571) );
  INV_X1 U10941 ( .A(n8568), .ZN(n8570) );
  INV_X1 U10942 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8569) );
  NAND2_X1 U10943 ( .A1(n8570), .A2(n8569), .ZN(n8588) );
  AOI22_X1 U10944 ( .A1(n8862), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6643), .B2(
        n9594), .ZN(n8572) );
  NAND2_X1 U10945 ( .A1(n10292), .A2(n9102), .ZN(n8580) );
  NAND2_X1 U10946 ( .A1(n6651), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8578) );
  NAND2_X1 U10947 ( .A1(n9035), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8577) );
  XNOR2_X1 U10948 ( .A(n8594), .B(P2_REG3_REG_6__SCAN_IN), .ZN(n10247) );
  NAND2_X1 U10949 ( .A1(n6652), .A2(n10247), .ZN(n8576) );
  NAND2_X1 U10950 ( .A1(n6860), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8575) );
  NAND4_X1 U10951 ( .A1(n8578), .A2(n8577), .A3(n8576), .A4(n8575), .ZN(n13528) );
  NAND2_X1 U10952 ( .A1(n9113), .A2(n13528), .ZN(n8579) );
  NAND2_X1 U10953 ( .A1(n8580), .A2(n8579), .ZN(n8583) );
  INV_X1 U10954 ( .A(n13528), .ZN(n10291) );
  NAND2_X1 U10955 ( .A1(n10292), .A2(n9113), .ZN(n8581) );
  OAI21_X1 U10956 ( .B1(n10291), .B2(n9121), .A(n8581), .ZN(n8582) );
  MUX2_X1 U10957 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n8991), .Z(n8587) );
  NAND2_X1 U10958 ( .A1(n8587), .A2(SI_7_), .ZN(n8607) );
  OAI21_X1 U10959 ( .B1(n8587), .B2(SI_7_), .A(n8607), .ZN(n8604) );
  XNOR2_X1 U10960 ( .A(n8606), .B(n8604), .ZN(n10799) );
  NAND2_X1 U10961 ( .A1(n10799), .A2(n9092), .ZN(n8591) );
  NAND2_X1 U10962 ( .A1(n8588), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8589) );
  XNOR2_X1 U10963 ( .A(n8589), .B(P2_IR_REG_7__SCAN_IN), .ZN(n13554) );
  AOI22_X1 U10964 ( .A1(n8862), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6643), .B2(
        n13554), .ZN(n8590) );
  NAND2_X1 U10965 ( .A1(n8591), .A2(n8590), .ZN(n15347) );
  NAND2_X1 U10966 ( .A1(n15347), .A2(n9113), .ZN(n8601) );
  NAND2_X1 U10967 ( .A1(n6651), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8599) );
  NAND2_X1 U10968 ( .A1(n9035), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8598) );
  NAND2_X1 U10969 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_REG3_REG_7__SCAN_IN), 
        .ZN(n8592) );
  NOR2_X1 U10970 ( .A1(n8594), .A2(n8592), .ZN(n8615) );
  INV_X1 U10971 ( .A(n8615), .ZN(n8616) );
  INV_X1 U10972 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8593) );
  INV_X1 U10973 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n13547) );
  OAI21_X1 U10974 ( .B1(n8594), .B2(n8593), .A(n13547), .ZN(n8595) );
  AND2_X1 U10975 ( .A1(n8616), .A2(n8595), .ZN(n10371) );
  NAND2_X1 U10976 ( .A1(n6652), .A2(n10371), .ZN(n8597) );
  NAND2_X1 U10977 ( .A1(n6860), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8596) );
  NAND4_X1 U10978 ( .A1(n8599), .A2(n8598), .A3(n8597), .A4(n8596), .ZN(n13527) );
  INV_X1 U10979 ( .A(n13527), .ZN(n10607) );
  OR2_X1 U10980 ( .A1(n9121), .A2(n10607), .ZN(n8600) );
  AOI22_X1 U10981 ( .A1(n15347), .A2(n9102), .B1(n9113), .B2(n13527), .ZN(
        n8602) );
  INV_X1 U10982 ( .A(n8604), .ZN(n8605) );
  MUX2_X1 U10983 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n8991), .Z(n8608) );
  NAND2_X1 U10984 ( .A1(n8608), .A2(SI_8_), .ZN(n8630) );
  OAI21_X1 U10985 ( .B1(n8608), .B2(SI_8_), .A(n8630), .ZN(n8627) );
  XNOR2_X1 U10986 ( .A(n8629), .B(n8627), .ZN(n10852) );
  NAND2_X1 U10987 ( .A1(n10852), .A2(n9092), .ZN(n8614) );
  INV_X1 U10988 ( .A(n8609), .ZN(n8611) );
  NOR2_X1 U10989 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n8610) );
  NAND2_X1 U10990 ( .A1(n8611), .A2(n8610), .ZN(n8636) );
  NAND2_X1 U10991 ( .A1(n8636), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8612) );
  XNOR2_X1 U10992 ( .A(n8612), .B(P2_IR_REG_8__SCAN_IN), .ZN(n9528) );
  AOI22_X1 U10993 ( .A1(n8862), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6643), .B2(
        n9528), .ZN(n8613) );
  NAND2_X1 U10994 ( .A1(n8614), .A2(n8613), .ZN(n10682) );
  NAND2_X1 U10995 ( .A1(n10682), .A2(n9102), .ZN(n8623) );
  NAND2_X1 U10996 ( .A1(n9035), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8621) );
  NAND2_X1 U10997 ( .A1(n6860), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8620) );
  NAND2_X1 U10998 ( .A1(n8615), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8641) );
  INV_X1 U10999 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n13257) );
  NAND2_X1 U11000 ( .A1(n8616), .A2(n13257), .ZN(n8617) );
  AND2_X1 U11001 ( .A1(n8641), .A2(n8617), .ZN(n10681) );
  NAND2_X1 U11002 ( .A1(n6652), .A2(n10681), .ZN(n8619) );
  NAND2_X1 U11003 ( .A1(n6651), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8618) );
  NAND4_X1 U11004 ( .A1(n8621), .A2(n8620), .A3(n8619), .A4(n8618), .ZN(n13526) );
  NAND2_X1 U11005 ( .A1(n9113), .A2(n13526), .ZN(n8622) );
  NAND2_X1 U11006 ( .A1(n8623), .A2(n8622), .ZN(n8626) );
  INV_X1 U11007 ( .A(n13526), .ZN(n10610) );
  NAND2_X1 U11008 ( .A1(n10682), .A2(n9113), .ZN(n8624) );
  OAI21_X1 U11009 ( .B1(n10610), .B2(n9121), .A(n8624), .ZN(n8625) );
  INV_X1 U11010 ( .A(n8627), .ZN(n8628) );
  MUX2_X1 U11011 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n6832), .Z(n8631) );
  NAND2_X1 U11012 ( .A1(n8631), .A2(SI_9_), .ZN(n8653) );
  OAI21_X1 U11013 ( .B1(n8631), .B2(SI_9_), .A(n8653), .ZN(n8632) );
  INV_X1 U11014 ( .A(n8632), .ZN(n8633) );
  NAND2_X1 U11015 ( .A1(n8634), .A2(n8633), .ZN(n8654) );
  OR2_X1 U11016 ( .A1(n8634), .A2(n8633), .ZN(n8635) );
  NAND2_X1 U11017 ( .A1(n8654), .A2(n8635), .ZN(n11079) );
  OR2_X1 U11018 ( .A1(n11079), .A2(n9109), .ZN(n8639) );
  NAND2_X1 U11019 ( .A1(n8656), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8637) );
  XNOR2_X1 U11020 ( .A(n8637), .B(P2_IR_REG_9__SCAN_IN), .ZN(n9629) );
  AOI22_X1 U11021 ( .A1(n8862), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6643), .B2(
        n9629), .ZN(n8638) );
  NAND2_X1 U11022 ( .A1(n15361), .A2(n9113), .ZN(n8648) );
  NAND2_X1 U11023 ( .A1(n6651), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8646) );
  NAND2_X1 U11024 ( .A1(n9035), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8645) );
  NAND2_X1 U11025 ( .A1(n8641), .A2(n8640), .ZN(n8642) );
  AND2_X1 U11026 ( .A1(n8661), .A2(n8642), .ZN(n10793) );
  NAND2_X1 U11027 ( .A1(n6652), .A2(n10793), .ZN(n8644) );
  NAND2_X1 U11028 ( .A1(n6860), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8643) );
  NAND4_X1 U11029 ( .A1(n8646), .A2(n8645), .A3(n8644), .A4(n8643), .ZN(n13525) );
  INV_X1 U11030 ( .A(n13525), .ZN(n10732) );
  OR2_X1 U11031 ( .A1(n9121), .A2(n10732), .ZN(n8647) );
  NAND2_X1 U11032 ( .A1(n8648), .A2(n8647), .ZN(n8651) );
  AOI22_X1 U11033 ( .A1(n15361), .A2(n9102), .B1(n9113), .B2(n13525), .ZN(
        n8649) );
  AOI21_X1 U11034 ( .B1(n8652), .B2(n8651), .A(n8649), .ZN(n8650) );
  MUX2_X1 U11035 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n8991), .Z(n8689) );
  NAND2_X1 U11036 ( .A1(n8694), .A2(n8689), .ZN(n8671) );
  NAND2_X1 U11037 ( .A1(n11071), .A2(n9092), .ZN(n8659) );
  NAND2_X1 U11038 ( .A1(n8674), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8657) );
  XNOR2_X1 U11039 ( .A(n8657), .B(P2_IR_REG_10__SCAN_IN), .ZN(n9533) );
  AOI22_X1 U11040 ( .A1(n8862), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6643), 
        .B2(n9533), .ZN(n8658) );
  NAND2_X1 U11041 ( .A1(n15369), .A2(n9102), .ZN(n8668) );
  NAND2_X1 U11042 ( .A1(n9035), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8666) );
  NAND2_X1 U11043 ( .A1(n6860), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n8665) );
  INV_X1 U11044 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8660) );
  INV_X1 U11045 ( .A(n8678), .ZN(n8680) );
  NAND2_X1 U11046 ( .A1(n8661), .A2(n8660), .ZN(n8662) );
  AND2_X1 U11047 ( .A1(n8680), .A2(n8662), .ZN(n10893) );
  NAND2_X1 U11048 ( .A1(n6652), .A2(n10893), .ZN(n8664) );
  NAND2_X1 U11049 ( .A1(n6651), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8663) );
  NAND4_X1 U11050 ( .A1(n8666), .A2(n8665), .A3(n8664), .A4(n8663), .ZN(n13524) );
  NAND2_X1 U11051 ( .A1(n9113), .A2(n13524), .ZN(n8667) );
  INV_X1 U11052 ( .A(n13524), .ZN(n10892) );
  NAND2_X1 U11053 ( .A1(n15369), .A2(n9113), .ZN(n8669) );
  OAI21_X1 U11054 ( .B1(n10892), .B2(n9121), .A(n8669), .ZN(n8670) );
  MUX2_X1 U11055 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n8991), .Z(n8695) );
  XNOR2_X1 U11056 ( .A(n8695), .B(SI_11_), .ZN(n8690) );
  XNOR2_X1 U11057 ( .A(n8690), .B(n8673), .ZN(n11377) );
  NAND2_X1 U11058 ( .A1(n11377), .A2(n9092), .ZN(n8677) );
  OAI21_X1 U11059 ( .B1(n8674), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8675) );
  XNOR2_X1 U11060 ( .A(n8675), .B(P2_IR_REG_11__SCAN_IN), .ZN(n9714) );
  AOI22_X1 U11061 ( .A1(n8862), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6643), 
        .B2(n9714), .ZN(n8676) );
  NAND2_X1 U11062 ( .A1(n11170), .A2(n9113), .ZN(n8687) );
  NAND2_X1 U11063 ( .A1(n6651), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8685) );
  NAND2_X1 U11064 ( .A1(n9035), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n8684) );
  INV_X1 U11065 ( .A(n8703), .ZN(n8705) );
  INV_X1 U11066 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8679) );
  NAND2_X1 U11067 ( .A1(n8680), .A2(n8679), .ZN(n8681) );
  AND2_X1 U11068 ( .A1(n8705), .A2(n8681), .ZN(n11169) );
  NAND2_X1 U11069 ( .A1(n6652), .A2(n11169), .ZN(n8683) );
  NAND2_X1 U11070 ( .A1(n6860), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8682) );
  NAND4_X1 U11071 ( .A1(n8685), .A2(n8684), .A3(n8683), .A4(n8682), .ZN(n13523) );
  INV_X1 U11072 ( .A(n13523), .ZN(n10986) );
  OR2_X1 U11073 ( .A1(n9121), .A2(n10986), .ZN(n8686) );
  AOI22_X1 U11074 ( .A1(n11170), .A2(n9102), .B1(n9113), .B2(n13523), .ZN(
        n8688) );
  INV_X1 U11075 ( .A(n8690), .ZN(n8691) );
  OAI21_X1 U11076 ( .B1(n8692), .B2(n9340), .A(n8691), .ZN(n8693) );
  NOR2_X1 U11077 ( .A1(n8695), .A2(SI_11_), .ZN(n8696) );
  MUX2_X1 U11078 ( .A(n9488), .B(n9444), .S(n8991), .Z(n8718) );
  XNOR2_X1 U11079 ( .A(n8718), .B(SI_12_), .ZN(n8717) );
  XNOR2_X1 U11080 ( .A(n6742), .B(n8717), .ZN(n11382) );
  NAND2_X1 U11081 ( .A1(n11382), .A2(n9092), .ZN(n8702) );
  OR2_X1 U11082 ( .A1(n8698), .A2(n8697), .ZN(n8699) );
  NAND2_X1 U11083 ( .A1(n8699), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8700) );
  XNOR2_X1 U11084 ( .A(n8700), .B(P2_IR_REG_12__SCAN_IN), .ZN(n9717) );
  AOI22_X1 U11085 ( .A1(n8862), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6643), 
        .B2(n9717), .ZN(n8701) );
  NAND2_X1 U11086 ( .A1(n11238), .A2(n9102), .ZN(n8712) );
  NAND2_X1 U11087 ( .A1(n6651), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8710) );
  NAND2_X1 U11088 ( .A1(n9035), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8709) );
  NAND2_X1 U11089 ( .A1(n8703), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8727) );
  INV_X1 U11090 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8704) );
  NAND2_X1 U11091 ( .A1(n8705), .A2(n8704), .ZN(n8706) );
  AND2_X1 U11092 ( .A1(n8727), .A2(n8706), .ZN(n11247) );
  NAND2_X1 U11093 ( .A1(n6652), .A2(n11247), .ZN(n8708) );
  NAND2_X1 U11094 ( .A1(n6860), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n8707) );
  NAND4_X1 U11095 ( .A1(n8710), .A2(n8709), .A3(n8708), .A4(n8707), .ZN(n13522) );
  NAND2_X1 U11096 ( .A1(n9113), .A2(n13522), .ZN(n8711) );
  NAND2_X1 U11097 ( .A1(n8712), .A2(n8711), .ZN(n8714) );
  AOI22_X1 U11098 ( .A1(n11238), .A2(n9113), .B1(n9102), .B2(n13522), .ZN(
        n8713) );
  MUX2_X1 U11099 ( .A(n8719), .B(n9638), .S(n6832), .Z(n8746) );
  XNOR2_X1 U11100 ( .A(n8746), .B(SI_13_), .ZN(n8744) );
  XNOR2_X1 U11101 ( .A(n8745), .B(n8744), .ZN(n11392) );
  NAND2_X1 U11102 ( .A1(n11392), .A2(n9092), .ZN(n8726) );
  NAND2_X1 U11103 ( .A1(n8720), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8721) );
  MUX2_X1 U11104 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8721), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n8724) );
  INV_X1 U11105 ( .A(n8723), .ZN(n8750) );
  AND2_X1 U11106 ( .A1(n8724), .A2(n8750), .ZN(n10079) );
  AOI22_X1 U11107 ( .A1(n8862), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6643), 
        .B2(n10079), .ZN(n8725) );
  NAND2_X1 U11108 ( .A1(n14885), .A2(n9113), .ZN(n8735) );
  NAND2_X1 U11109 ( .A1(n6651), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8733) );
  NAND2_X1 U11110 ( .A1(n8727), .A2(n9712), .ZN(n8728) );
  AND2_X1 U11111 ( .A1(n8754), .A2(n8728), .ZN(n11294) );
  NAND2_X1 U11112 ( .A1(n6652), .A2(n11294), .ZN(n8732) );
  INV_X1 U11113 ( .A(n9035), .ZN(n9083) );
  INV_X1 U11114 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8729) );
  OR2_X1 U11115 ( .A1(n9083), .A2(n8729), .ZN(n8731) );
  OR2_X1 U11116 ( .A1(n9041), .A2(n9713), .ZN(n8730) );
  OR2_X1 U11117 ( .A1(n9121), .A2(n11577), .ZN(n8734) );
  NAND2_X1 U11118 ( .A1(n8735), .A2(n8734), .ZN(n8740) );
  NAND2_X1 U11119 ( .A1(n8741), .A2(n8740), .ZN(n8739) );
  NAND2_X1 U11120 ( .A1(n14885), .A2(n9102), .ZN(n8737) );
  INV_X1 U11121 ( .A(n11577), .ZN(n11567) );
  NAND2_X1 U11122 ( .A1(n9113), .A2(n11567), .ZN(n8736) );
  NAND2_X1 U11123 ( .A1(n8737), .A2(n8736), .ZN(n8738) );
  NAND2_X1 U11124 ( .A1(n8739), .A2(n8738), .ZN(n8743) );
  OR2_X1 U11125 ( .A1(n8741), .A2(n8740), .ZN(n8742) );
  NAND2_X1 U11126 ( .A1(n8746), .A2(n9375), .ZN(n8747) );
  MUX2_X1 U11127 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n6832), .Z(n8766) );
  XNOR2_X1 U11128 ( .A(n8766), .B(n9377), .ZN(n8749) );
  XNOR2_X1 U11129 ( .A(n8768), .B(n8749), .ZN(n11367) );
  NAND2_X1 U11130 ( .A1(n11367), .A2(n9092), .ZN(n8753) );
  NAND2_X1 U11131 ( .A1(n8750), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8751) );
  XNOR2_X1 U11132 ( .A(n8751), .B(P2_IR_REG_14__SCAN_IN), .ZN(n10704) );
  AOI22_X1 U11133 ( .A1(n8862), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6643), 
        .B2(n10704), .ZN(n8752) );
  NAND2_X1 U11134 ( .A1(n14849), .A2(n9102), .ZN(n8761) );
  INV_X1 U11135 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n13189) );
  NAND2_X1 U11136 ( .A1(n8754), .A2(n13189), .ZN(n8755) );
  AND2_X1 U11137 ( .A1(n8775), .A2(n8755), .ZN(n14843) );
  NAND2_X1 U11138 ( .A1(n14843), .A2(n6652), .ZN(n8759) );
  NAND2_X1 U11139 ( .A1(n9035), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n8758) );
  NAND2_X1 U11140 ( .A1(n6860), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8757) );
  NAND2_X1 U11141 ( .A1(n6651), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8756) );
  NAND4_X1 U11142 ( .A1(n8759), .A2(n8758), .A3(n8757), .A4(n8756), .ZN(n13521) );
  NAND2_X1 U11143 ( .A1(n9113), .A2(n13521), .ZN(n8760) );
  NAND2_X1 U11144 ( .A1(n8761), .A2(n8760), .ZN(n8763) );
  AOI22_X1 U11145 ( .A1(n14849), .A2(n9113), .B1(n9102), .B2(n13521), .ZN(
        n8762) );
  AOI21_X1 U11146 ( .B1(n8764), .B2(n8763), .A(n8762), .ZN(n8765) );
  INV_X1 U11147 ( .A(n8766), .ZN(n8767) );
  NAND2_X1 U11148 ( .A1(n8768), .A2(n9377), .ZN(n8769) );
  MUX2_X1 U11149 ( .A(n9703), .B(n13278), .S(n6832), .Z(n8789) );
  XNOR2_X1 U11150 ( .A(n8789), .B(SI_15_), .ZN(n8787) );
  XNOR2_X1 U11151 ( .A(n8788), .B(n8787), .ZN(n11534) );
  NAND2_X1 U11152 ( .A1(n11534), .A2(n9092), .ZN(n8773) );
  NAND2_X1 U11153 ( .A1(n8770), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8771) );
  XNOR2_X1 U11154 ( .A(n8771), .B(P2_IR_REG_15__SCAN_IN), .ZN(n15253) );
  AOI22_X1 U11155 ( .A1(n8862), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6643), 
        .B2(n15253), .ZN(n8772) );
  NAND2_X1 U11156 ( .A1(n14830), .A2(n9113), .ZN(n8783) );
  INV_X1 U11157 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8781) );
  INV_X1 U11158 ( .A(n8796), .ZN(n8798) );
  NAND2_X1 U11159 ( .A1(n8775), .A2(n8774), .ZN(n8776) );
  NAND2_X1 U11160 ( .A1(n8798), .A2(n8776), .ZN(n14826) );
  OR2_X1 U11161 ( .A1(n14826), .A2(n8935), .ZN(n8780) );
  NAND2_X1 U11162 ( .A1(n6651), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8778) );
  NAND2_X1 U11163 ( .A1(n9035), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n8777) );
  AND2_X1 U11164 ( .A1(n8778), .A2(n8777), .ZN(n8779) );
  OAI211_X1 U11165 ( .C1(n9041), .C2(n8781), .A(n8780), .B(n8779), .ZN(n13520)
         );
  NAND2_X1 U11166 ( .A1(n9102), .A2(n13520), .ZN(n8782) );
  NAND2_X1 U11167 ( .A1(n14830), .A2(n9102), .ZN(n8785) );
  NAND2_X1 U11168 ( .A1(n9113), .A2(n13520), .ZN(n8784) );
  NAND2_X1 U11169 ( .A1(n8785), .A2(n8784), .ZN(n8786) );
  NAND2_X1 U11170 ( .A1(n8789), .A2(n9547), .ZN(n8790) );
  MUX2_X1 U11171 ( .A(n9779), .B(n9781), .S(n6832), .Z(n8808) );
  XNOR2_X1 U11172 ( .A(n8808), .B(SI_16_), .ZN(n8806) );
  NAND2_X1 U11173 ( .A1(n11670), .A2(n9092), .ZN(n8795) );
  INV_X1 U11174 ( .A(n8791), .ZN(n8792) );
  NAND2_X1 U11175 ( .A1(n8792), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8793) );
  XNOR2_X1 U11176 ( .A(n8793), .B(P2_IR_REG_16__SCAN_IN), .ZN(n10702) );
  AOI22_X1 U11177 ( .A1(n8862), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n10702), 
        .B2(n6643), .ZN(n8794) );
  NAND2_X1 U11178 ( .A1(n13750), .A2(n9102), .ZN(n8803) );
  INV_X1 U11179 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n10697) );
  NAND2_X1 U11180 ( .A1(n8796), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8817) );
  INV_X1 U11181 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8797) );
  NAND2_X1 U11182 ( .A1(n8798), .A2(n8797), .ZN(n8799) );
  NAND2_X1 U11183 ( .A1(n8817), .A2(n8799), .ZN(n13747) );
  OR2_X1 U11184 ( .A1(n13747), .A2(n8935), .ZN(n8801) );
  AOI22_X1 U11185 ( .A1(n9035), .A2(P2_REG0_REG_16__SCAN_IN), .B1(n6651), .B2(
        P2_REG1_REG_16__SCAN_IN), .ZN(n8800) );
  OAI211_X1 U11186 ( .C1(n9041), .C2(n10697), .A(n8801), .B(n8800), .ZN(n13519) );
  NAND2_X1 U11187 ( .A1(n9113), .A2(n13519), .ZN(n8802) );
  NAND2_X1 U11188 ( .A1(n8803), .A2(n8802), .ZN(n8805) );
  AOI22_X1 U11189 ( .A1(n13750), .A2(n9113), .B1(n9102), .B2(n13519), .ZN(
        n8804) );
  NAND2_X1 U11190 ( .A1(n8808), .A2(n9607), .ZN(n8809) );
  MUX2_X1 U11191 ( .A(n9876), .B(n9915), .S(n6832), .Z(n8832) );
  XNOR2_X1 U11192 ( .A(n8832), .B(SI_17_), .ZN(n8810) );
  XNOR2_X1 U11193 ( .A(n8834), .B(n8810), .ZN(n11675) );
  NAND2_X1 U11194 ( .A1(n11675), .A2(n9092), .ZN(n8815) );
  NAND2_X1 U11195 ( .A1(n8811), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8812) );
  MUX2_X1 U11196 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8812), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n8813) );
  OR2_X1 U11197 ( .A1(n8811), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n8836) );
  AND2_X1 U11198 ( .A1(n8813), .A2(n8836), .ZN(n11180) );
  AOI22_X1 U11199 ( .A1(n11180), .A2(n6643), .B1(P1_DATAO_REG_17__SCAN_IN), 
        .B2(n8862), .ZN(n8814) );
  INV_X1 U11200 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8816) );
  NAND2_X1 U11201 ( .A1(n8817), .A2(n8816), .ZN(n8818) );
  NAND2_X1 U11202 ( .A1(n8840), .A2(n8818), .ZN(n13442) );
  AOI22_X1 U11203 ( .A1(n9035), .A2(P2_REG0_REG_17__SCAN_IN), .B1(n6651), .B2(
        P2_REG1_REG_17__SCAN_IN), .ZN(n8820) );
  NAND2_X1 U11204 ( .A1(n6860), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8819) );
  OAI211_X1 U11205 ( .C1(n13442), .C2(n8935), .A(n8820), .B(n8819), .ZN(n13518) );
  AND2_X1 U11206 ( .A1(n13518), .A2(n9102), .ZN(n8821) );
  AOI21_X1 U11207 ( .B1(n11923), .B2(n9113), .A(n8821), .ZN(n8828) );
  INV_X1 U11208 ( .A(n8828), .ZN(n8822) );
  NAND2_X1 U11209 ( .A1(n8827), .A2(n8822), .ZN(n8826) );
  NAND2_X1 U11210 ( .A1(n11923), .A2(n9102), .ZN(n8824) );
  NAND2_X1 U11211 ( .A1(n13518), .A2(n9113), .ZN(n8823) );
  NAND2_X1 U11212 ( .A1(n8824), .A2(n8823), .ZN(n8825) );
  NAND2_X1 U11213 ( .A1(n8826), .A2(n8825), .ZN(n8831) );
  INV_X1 U11214 ( .A(n8827), .ZN(n8829) );
  NAND2_X1 U11215 ( .A1(n8829), .A2(n8828), .ZN(n8830) );
  INV_X1 U11216 ( .A(n8832), .ZN(n8833) );
  MUX2_X1 U11217 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n6832), .Z(n8854) );
  XNOR2_X1 U11218 ( .A(n8854), .B(SI_18_), .ZN(n8835) );
  XNOR2_X1 U11219 ( .A(n8856), .B(n8835), .ZN(n11685) );
  NAND2_X1 U11220 ( .A1(n11685), .A2(n9092), .ZN(n8839) );
  NAND2_X1 U11221 ( .A1(n8836), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8837) );
  XNOR2_X1 U11222 ( .A(n8837), .B(P2_IR_REG_18__SCAN_IN), .ZN(n11596) );
  AOI22_X1 U11223 ( .A1(n11596), .A2(n6643), .B1(P1_DATAO_REG_18__SCAN_IN), 
        .B2(n8862), .ZN(n8838) );
  NAND2_X1 U11224 ( .A1(n13822), .A2(n9102), .ZN(n8849) );
  INV_X1 U11225 ( .A(n8865), .ZN(n8867) );
  NAND2_X1 U11226 ( .A1(n8840), .A2(n11185), .ZN(n8841) );
  NAND2_X1 U11227 ( .A1(n8867), .A2(n8841), .ZN(n13730) );
  OR2_X1 U11228 ( .A1(n13730), .A2(n8935), .ZN(n8847) );
  INV_X1 U11229 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8844) );
  NAND2_X1 U11230 ( .A1(n9035), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8843) );
  NAND2_X1 U11231 ( .A1(n6651), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8842) );
  OAI211_X1 U11232 ( .C1(n8844), .C2(n9041), .A(n8843), .B(n8842), .ZN(n8845)
         );
  INV_X1 U11233 ( .A(n8845), .ZN(n8846) );
  NAND2_X1 U11234 ( .A1(n8847), .A2(n8846), .ZN(n13517) );
  NAND2_X1 U11235 ( .A1(n13517), .A2(n9113), .ZN(n8848) );
  NAND2_X1 U11236 ( .A1(n8849), .A2(n8848), .ZN(n8851) );
  AOI22_X1 U11237 ( .A1(n13822), .A2(n9113), .B1(n9102), .B2(n13517), .ZN(
        n8850) );
  AOI21_X1 U11238 ( .B1(n8852), .B2(n8851), .A(n8850), .ZN(n8853) );
  NOR2_X1 U11239 ( .A1(n8857), .A2(n9690), .ZN(n8855) );
  NAND2_X1 U11240 ( .A1(n8857), .A2(n9690), .ZN(n8858) );
  MUX2_X1 U11241 ( .A(n10385), .B(n10623), .S(n6832), .Z(n8859) );
  INV_X1 U11242 ( .A(n8859), .ZN(n8860) );
  NAND2_X1 U11243 ( .A1(n8860), .A2(SI_19_), .ZN(n8861) );
  XNOR2_X1 U11244 ( .A(n8880), .B(n8879), .ZN(n11698) );
  NAND2_X1 U11245 ( .A1(n11698), .A2(n9092), .ZN(n8864) );
  AOI22_X1 U11246 ( .A1(n6843), .A2(n6643), .B1(n8862), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n8863) );
  NAND2_X1 U11247 ( .A1(n13818), .A2(n9113), .ZN(n8875) );
  INV_X1 U11248 ( .A(n8884), .ZN(n8886) );
  INV_X1 U11249 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8866) );
  NAND2_X1 U11250 ( .A1(n8867), .A2(n8866), .ZN(n8868) );
  AND2_X1 U11251 ( .A1(n8886), .A2(n8868), .ZN(n13718) );
  NAND2_X1 U11252 ( .A1(n13718), .A2(n6652), .ZN(n8873) );
  INV_X1 U11253 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n13237) );
  NAND2_X1 U11254 ( .A1(n6651), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n8870) );
  NAND2_X1 U11255 ( .A1(n6860), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8869) );
  OAI211_X1 U11256 ( .C1(n9083), .C2(n13237), .A(n8870), .B(n8869), .ZN(n8871)
         );
  INV_X1 U11257 ( .A(n8871), .ZN(n8872) );
  NAND2_X1 U11258 ( .A1(n8873), .A2(n8872), .ZN(n13516) );
  NAND2_X1 U11259 ( .A1(n13516), .A2(n9102), .ZN(n8874) );
  NAND2_X1 U11260 ( .A1(n8875), .A2(n8874), .ZN(n8877) );
  AOI22_X1 U11261 ( .A1(n13818), .A2(n9102), .B1(n9113), .B2(n13516), .ZN(
        n8876) );
  XNOR2_X1 U11262 ( .A(n8925), .B(SI_20_), .ZN(n8903) );
  MUX2_X1 U11263 ( .A(n13291), .B(n10829), .S(n6832), .Z(n8926) );
  XNOR2_X1 U11264 ( .A(n8903), .B(n8926), .ZN(n11711) );
  NAND2_X1 U11265 ( .A1(n11711), .A2(n9092), .ZN(n8883) );
  OR2_X1 U11266 ( .A1(n9110), .A2(n10829), .ZN(n8882) );
  NAND2_X1 U11267 ( .A1(n13813), .A2(n9102), .ZN(n8895) );
  INV_X1 U11268 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8885) );
  NAND2_X1 U11269 ( .A1(n8886), .A2(n8885), .ZN(n8887) );
  NAND2_X1 U11270 ( .A1(n8911), .A2(n8887), .ZN(n13466) );
  OR2_X1 U11271 ( .A1(n13466), .A2(n8935), .ZN(n8893) );
  INV_X1 U11272 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8890) );
  NAND2_X1 U11273 ( .A1(n9035), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8889) );
  NAND2_X1 U11274 ( .A1(n6651), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8888) );
  OAI211_X1 U11275 ( .C1(n9041), .C2(n8890), .A(n8889), .B(n8888), .ZN(n8891)
         );
  INV_X1 U11276 ( .A(n8891), .ZN(n8892) );
  NAND2_X1 U11277 ( .A1(n8893), .A2(n8892), .ZN(n13515) );
  NAND2_X1 U11278 ( .A1(n13515), .A2(n9113), .ZN(n8894) );
  NAND2_X1 U11279 ( .A1(n8895), .A2(n8894), .ZN(n8899) );
  INV_X1 U11280 ( .A(n13515), .ZN(n9158) );
  NAND2_X1 U11281 ( .A1(n13813), .A2(n9113), .ZN(n8896) );
  OAI21_X1 U11282 ( .B1(n9158), .B2(n9121), .A(n8896), .ZN(n8897) );
  NAND2_X1 U11283 ( .A1(n8898), .A2(n8897), .ZN(n8902) );
  INV_X1 U11284 ( .A(n8926), .ZN(n8924) );
  NAND2_X1 U11285 ( .A1(n8903), .A2(n8924), .ZN(n8905) );
  OR2_X1 U11286 ( .A1(n8925), .A2(n10110), .ZN(n8904) );
  NAND2_X1 U11287 ( .A1(n8905), .A2(n8904), .ZN(n8907) );
  MUX2_X1 U11288 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n6832), .Z(n8927) );
  XNOR2_X1 U11289 ( .A(n8927), .B(SI_21_), .ZN(n8906) );
  NAND2_X1 U11290 ( .A1(n11723), .A2(n9092), .ZN(n8909) );
  OR2_X1 U11291 ( .A1(n9110), .A2(n10900), .ZN(n8908) );
  NAND2_X1 U11292 ( .A1(n13804), .A2(n9113), .ZN(n8920) );
  INV_X1 U11293 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8910) );
  NAND2_X1 U11294 ( .A1(n8911), .A2(n8910), .ZN(n8912) );
  AND2_X1 U11295 ( .A1(n8932), .A2(n8912), .ZN(n13682) );
  NAND2_X1 U11296 ( .A1(n13682), .A2(n6652), .ZN(n8918) );
  INV_X1 U11297 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8915) );
  NAND2_X1 U11298 ( .A1(n6651), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8914) );
  NAND2_X1 U11299 ( .A1(n6860), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8913) );
  OAI211_X1 U11300 ( .C1(n9083), .C2(n8915), .A(n8914), .B(n8913), .ZN(n8916)
         );
  INV_X1 U11301 ( .A(n8916), .ZN(n8917) );
  NAND2_X1 U11302 ( .A1(n8918), .A2(n8917), .ZN(n13514) );
  NAND2_X1 U11303 ( .A1(n13514), .A2(n9102), .ZN(n8919) );
  NAND2_X1 U11304 ( .A1(n8920), .A2(n8919), .ZN(n8922) );
  AOI22_X1 U11305 ( .A1(n13804), .A2(n9102), .B1(n9113), .B2(n13514), .ZN(
        n8921) );
  NOR2_X1 U11306 ( .A1(n8926), .A2(n10110), .ZN(n8928) );
  AOI22_X1 U11307 ( .A1(n8928), .A2(n6661), .B1(n8927), .B2(SI_21_), .ZN(n8929) );
  MUX2_X1 U11308 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n6832), .Z(n8948) );
  XNOR2_X1 U11309 ( .A(n11735), .B(n8948), .ZN(n11025) );
  NAND2_X1 U11310 ( .A1(n11025), .A2(n9092), .ZN(n8931) );
  OR2_X1 U11311 ( .A1(n9110), .A2(n11027), .ZN(n8930) );
  NAND2_X1 U11312 ( .A1(n13800), .A2(n9102), .ZN(n8943) );
  INV_X1 U11313 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13477) );
  NAND2_X1 U11314 ( .A1(n8932), .A2(n13477), .ZN(n8934) );
  INV_X1 U11315 ( .A(n8953), .ZN(n8933) );
  NAND2_X1 U11316 ( .A1(n8934), .A2(n8933), .ZN(n13669) );
  OR2_X1 U11317 ( .A1(n13669), .A2(n8935), .ZN(n8941) );
  INV_X1 U11318 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8938) );
  NAND2_X1 U11319 ( .A1(n6651), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8937) );
  NAND2_X1 U11320 ( .A1(n6860), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8936) );
  OAI211_X1 U11321 ( .C1(n9083), .C2(n8938), .A(n8937), .B(n8936), .ZN(n8939)
         );
  INV_X1 U11322 ( .A(n8939), .ZN(n8940) );
  NAND2_X1 U11323 ( .A1(n8941), .A2(n8940), .ZN(n13513) );
  NAND2_X1 U11324 ( .A1(n13513), .A2(n9113), .ZN(n8942) );
  NAND2_X1 U11325 ( .A1(n8943), .A2(n8942), .ZN(n8946) );
  NAND2_X1 U11326 ( .A1(n13800), .A2(n9113), .ZN(n8945) );
  NAND2_X1 U11327 ( .A1(n13513), .A2(n9102), .ZN(n8944) );
  NAND2_X1 U11328 ( .A1(n8949), .A2(SI_22_), .ZN(n8950) );
  MUX2_X1 U11329 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n6832), .Z(n8966) );
  XNOR2_X1 U11330 ( .A(n8966), .B(SI_23_), .ZN(n8964) );
  XNOR2_X1 U11331 ( .A(n8965), .B(n8964), .ZN(n11745) );
  NAND2_X1 U11332 ( .A1(n11745), .A2(n9092), .ZN(n8952) );
  OR2_X1 U11333 ( .A1(n9110), .A2(n11139), .ZN(n8951) );
  NAND2_X1 U11334 ( .A1(n13795), .A2(n9113), .ZN(n8960) );
  NAND2_X1 U11335 ( .A1(n6651), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8958) );
  NAND2_X1 U11336 ( .A1(n9035), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8957) );
  NAND2_X1 U11337 ( .A1(n8953), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8969) );
  OAI21_X1 U11338 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(n8953), .A(n8969), .ZN(
        n13654) );
  INV_X1 U11339 ( .A(n13654), .ZN(n8954) );
  NAND2_X1 U11340 ( .A1(n6652), .A2(n8954), .ZN(n8956) );
  NAND2_X1 U11341 ( .A1(n6860), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8955) );
  NAND4_X1 U11342 ( .A1(n8958), .A2(n8957), .A3(n8956), .A4(n8955), .ZN(n13512) );
  INV_X1 U11343 ( .A(n13512), .ZN(n11823) );
  OR2_X1 U11344 ( .A1(n9121), .A2(n11823), .ZN(n8959) );
  NAND2_X1 U11345 ( .A1(n8960), .A2(n8959), .ZN(n8962) );
  AOI22_X1 U11346 ( .A1(n13795), .A2(n9102), .B1(n9113), .B2(n13512), .ZN(
        n8961) );
  MUX2_X1 U11347 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n8991), .Z(n8984) );
  XNOR2_X1 U11348 ( .A(n8983), .B(n8984), .ZN(n11665) );
  NAND2_X1 U11349 ( .A1(n11665), .A2(n9092), .ZN(n8968) );
  OR2_X1 U11350 ( .A1(n9110), .A2(n11351), .ZN(n8967) );
  NAND2_X1 U11351 ( .A1(n13790), .A2(n9102), .ZN(n8977) );
  NAND2_X1 U11352 ( .A1(n6651), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8975) );
  NAND2_X1 U11353 ( .A1(n9035), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8974) );
  INV_X1 U11354 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13457) );
  NAND2_X1 U11355 ( .A1(n13457), .A2(n8969), .ZN(n8971) );
  INV_X1 U11356 ( .A(n8969), .ZN(n8970) );
  NAND2_X1 U11357 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(n8970), .ZN(n9055) );
  AND2_X1 U11358 ( .A1(n8971), .A2(n9055), .ZN(n13642) );
  NAND2_X1 U11359 ( .A1(n6652), .A2(n13642), .ZN(n8973) );
  NAND2_X1 U11360 ( .A1(n6860), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8972) );
  NAND4_X1 U11361 ( .A1(n8975), .A2(n8974), .A3(n8973), .A4(n8972), .ZN(n13511) );
  NAND2_X1 U11362 ( .A1(n9113), .A2(n13511), .ZN(n8976) );
  NAND2_X1 U11363 ( .A1(n8977), .A2(n8976), .ZN(n8981) );
  INV_X1 U11364 ( .A(n13511), .ZN(n13398) );
  NAND2_X1 U11365 ( .A1(n13790), .A2(n9113), .ZN(n8978) );
  OAI21_X1 U11366 ( .B1(n13398), .B2(n9113), .A(n8978), .ZN(n8979) );
  INV_X1 U11367 ( .A(n8979), .ZN(n8980) );
  AOI21_X1 U11368 ( .B1(n8982), .B2(n8981), .A(n8980), .ZN(n9067) );
  NAND2_X1 U11369 ( .A1(n8985), .A2(SI_24_), .ZN(n8986) );
  MUX2_X1 U11370 ( .A(n11657), .B(n11471), .S(n8991), .Z(n8987) );
  INV_X1 U11371 ( .A(SI_25_), .ZN(n11253) );
  NAND2_X1 U11372 ( .A1(n8987), .A2(n11253), .ZN(n8990) );
  INV_X1 U11373 ( .A(n8987), .ZN(n8988) );
  NAND2_X1 U11374 ( .A1(n8988), .A2(SI_25_), .ZN(n8989) );
  NAND2_X1 U11375 ( .A1(n8990), .A2(n8989), .ZN(n9050) );
  MUX2_X1 U11376 ( .A(n14695), .B(n13853), .S(n6832), .Z(n9030) );
  NAND2_X1 U11377 ( .A1(n9032), .A2(n11304), .ZN(n8992) );
  MUX2_X1 U11378 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n8991), .Z(n9012) );
  NOR2_X1 U11379 ( .A1(n9012), .A2(SI_27_), .ZN(n8993) );
  NAND2_X1 U11380 ( .A1(n9012), .A2(SI_27_), .ZN(n8994) );
  MUX2_X1 U11381 ( .A(n11810), .B(n8998), .S(n8991), .Z(n8995) );
  INV_X1 U11382 ( .A(SI_28_), .ZN(n11979) );
  NAND2_X1 U11383 ( .A1(n8995), .A2(n11979), .ZN(n9070) );
  INV_X1 U11384 ( .A(n8995), .ZN(n8996) );
  NAND2_X1 U11385 ( .A1(n8996), .A2(SI_28_), .ZN(n8997) );
  NAND2_X1 U11386 ( .A1(n9070), .A2(n8997), .ZN(n9068) );
  NAND2_X1 U11387 ( .A1(n11809), .A2(n9092), .ZN(n9000) );
  OR2_X1 U11388 ( .A1(n9110), .A2(n8998), .ZN(n8999) );
  NAND2_X1 U11389 ( .A1(n9035), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n9008) );
  NAND2_X1 U11390 ( .A1(n6860), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n9007) );
  INV_X1 U11391 ( .A(n9055), .ZN(n9001) );
  NAND2_X1 U11392 ( .A1(n9002), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n9095) );
  INV_X1 U11393 ( .A(n9002), .ZN(n9021) );
  INV_X1 U11394 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9003) );
  NAND2_X1 U11395 ( .A1(n9021), .A2(n9003), .ZN(n9004) );
  NAND2_X1 U11396 ( .A1(n6652), .A2(n13586), .ZN(n9006) );
  NAND2_X1 U11397 ( .A1(n6651), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n9005) );
  NOR2_X1 U11398 ( .A1(n9121), .A2(n13387), .ZN(n9009) );
  AOI21_X1 U11399 ( .B1(n13767), .B2(n9113), .A(n9009), .ZN(n9135) );
  NAND2_X1 U11400 ( .A1(n13767), .A2(n9102), .ZN(n9011) );
  NAND2_X1 U11401 ( .A1(n9113), .A2(n13507), .ZN(n9010) );
  NAND2_X1 U11402 ( .A1(n9011), .A2(n9010), .ZN(n9134) );
  NAND2_X1 U11403 ( .A1(n9135), .A2(n9134), .ZN(n9131) );
  INV_X1 U11404 ( .A(n9012), .ZN(n9013) );
  XNOR2_X1 U11405 ( .A(n9013), .B(SI_27_), .ZN(n9014) );
  NAND2_X1 U11406 ( .A1(n11642), .A2(n9092), .ZN(n9017) );
  OR2_X1 U11407 ( .A1(n9110), .A2(n11632), .ZN(n9016) );
  NAND2_X1 U11408 ( .A1(n6651), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n9025) );
  NAND2_X1 U11409 ( .A1(n9035), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n9024) );
  INV_X1 U11410 ( .A(n9018), .ZN(n9039) );
  INV_X1 U11411 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9019) );
  NAND2_X1 U11412 ( .A1(n9039), .A2(n9019), .ZN(n9020) );
  NAND2_X1 U11413 ( .A1(n6652), .A2(n13598), .ZN(n9023) );
  NAND2_X1 U11414 ( .A1(n6860), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n9022) );
  NOR2_X1 U11415 ( .A1(n9121), .A2(n13493), .ZN(n9026) );
  AOI21_X1 U11416 ( .B1(n13773), .B2(n9113), .A(n9026), .ZN(n9128) );
  NAND2_X1 U11417 ( .A1(n13773), .A2(n9102), .ZN(n9028) );
  INV_X1 U11418 ( .A(n13493), .ZN(n13508) );
  NAND2_X1 U11419 ( .A1(n9113), .A2(n13508), .ZN(n9027) );
  NAND2_X1 U11420 ( .A1(n9028), .A2(n9027), .ZN(n9127) );
  NAND2_X1 U11421 ( .A1(n9128), .A2(n9127), .ZN(n9029) );
  XNOR2_X1 U11422 ( .A(n9030), .B(SI_26_), .ZN(n9031) );
  XNOR2_X1 U11423 ( .A(n9032), .B(n9031), .ZN(n13851) );
  NAND2_X1 U11424 ( .A1(n13851), .A2(n9092), .ZN(n9034) );
  OR2_X1 U11425 ( .A1(n9110), .A2(n13853), .ZN(n9033) );
  NAND2_X1 U11426 ( .A1(n9035), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n9045) );
  INV_X1 U11427 ( .A(n9036), .ZN(n9057) );
  INV_X1 U11428 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9037) );
  NAND2_X1 U11429 ( .A1(n9057), .A2(n9037), .ZN(n9038) );
  NAND2_X1 U11430 ( .A1(n6652), .A2(n13614), .ZN(n9044) );
  NAND2_X1 U11431 ( .A1(n6651), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n9043) );
  INV_X1 U11432 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n9040) );
  OR2_X1 U11433 ( .A1(n9041), .A2(n9040), .ZN(n9042) );
  NOR2_X1 U11434 ( .A1(n9121), .A2(n13421), .ZN(n9046) );
  AOI21_X1 U11435 ( .B1(n13779), .B2(n9113), .A(n9046), .ZN(n9125) );
  NAND2_X1 U11436 ( .A1(n13779), .A2(n9102), .ZN(n9048) );
  NAND2_X1 U11437 ( .A1(n9113), .A2(n13509), .ZN(n9047) );
  NAND2_X1 U11438 ( .A1(n9048), .A2(n9047), .ZN(n9124) );
  AND2_X1 U11439 ( .A1(n9125), .A2(n9124), .ZN(n9049) );
  XNOR2_X1 U11440 ( .A(n9051), .B(n9050), .ZN(n11656) );
  NAND2_X1 U11441 ( .A1(n11656), .A2(n9092), .ZN(n9053) );
  OR2_X1 U11442 ( .A1(n9110), .A2(n11471), .ZN(n9052) );
  NAND2_X1 U11443 ( .A1(n6651), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n9061) );
  NAND2_X1 U11444 ( .A1(n9035), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n9060) );
  INV_X1 U11445 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9054) );
  NAND2_X1 U11446 ( .A1(n9055), .A2(n9054), .ZN(n9056) );
  NAND2_X1 U11447 ( .A1(n6652), .A2(n13631), .ZN(n9059) );
  NAND2_X1 U11448 ( .A1(n6860), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n9058) );
  NOR2_X1 U11449 ( .A1(n9113), .A2(n13494), .ZN(n9062) );
  AOI21_X1 U11450 ( .B1(n13785), .B2(n9113), .A(n9062), .ZN(n9089) );
  NAND2_X1 U11451 ( .A1(n13785), .A2(n9102), .ZN(n9064) );
  NAND2_X1 U11452 ( .A1(n9113), .A2(n13510), .ZN(n9063) );
  NAND2_X1 U11453 ( .A1(n9064), .A2(n9063), .ZN(n9088) );
  NAND2_X1 U11454 ( .A1(n9089), .A2(n9088), .ZN(n9065) );
  INV_X1 U11455 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n11770) );
  INV_X1 U11456 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13846) );
  MUX2_X1 U11457 ( .A(n11770), .B(n13846), .S(n8991), .Z(n9071) );
  XNOR2_X1 U11458 ( .A(n9071), .B(SI_29_), .ZN(n9090) );
  NAND2_X1 U11459 ( .A1(n9091), .A2(n9090), .ZN(n9073) );
  INV_X1 U11460 ( .A(SI_29_), .ZN(n13030) );
  NAND2_X1 U11461 ( .A1(n9071), .A2(n13030), .ZN(n9072) );
  MUX2_X1 U11462 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n8991), .Z(n9074) );
  NAND2_X1 U11463 ( .A1(n9074), .A2(SI_30_), .ZN(n9075) );
  OAI21_X1 U11464 ( .B1(n9074), .B2(SI_30_), .A(n9075), .ZN(n9105) );
  MUX2_X1 U11465 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n8991), .Z(n9076) );
  XNOR2_X1 U11466 ( .A(n9076), .B(SI_31_), .ZN(n9077) );
  NAND2_X1 U11467 ( .A1(n14692), .A2(n9092), .ZN(n9081) );
  INV_X1 U11468 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9079) );
  OR2_X1 U11469 ( .A1(n9110), .A2(n9079), .ZN(n9080) );
  NAND2_X1 U11470 ( .A1(n6651), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n9086) );
  NAND2_X1 U11471 ( .A1(n6860), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9085) );
  INV_X1 U11472 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9082) );
  OR2_X1 U11473 ( .A1(n9083), .A2(n9082), .ZN(n9084) );
  AND3_X1 U11474 ( .A1(n9086), .A2(n9085), .A3(n9084), .ZN(n9112) );
  NAND2_X1 U11475 ( .A1(n11772), .A2(n9092), .ZN(n9094) );
  OR2_X1 U11476 ( .A1(n9110), .A2(n13846), .ZN(n9093) );
  NAND2_X1 U11477 ( .A1(n6651), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n9100) );
  NAND2_X1 U11478 ( .A1(n9035), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n9099) );
  INV_X1 U11479 ( .A(n9095), .ZN(n11848) );
  NAND2_X1 U11480 ( .A1(n6652), .A2(n11848), .ZN(n9098) );
  NAND2_X1 U11481 ( .A1(n6860), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n9097) );
  NOR2_X1 U11482 ( .A1(n9121), .A2(n11972), .ZN(n9101) );
  AOI21_X1 U11483 ( .B1(n13762), .B2(n9113), .A(n9101), .ZN(n9137) );
  NAND2_X1 U11484 ( .A1(n13762), .A2(n9102), .ZN(n9104) );
  INV_X1 U11485 ( .A(n11972), .ZN(n13506) );
  NAND2_X1 U11486 ( .A1(n9113), .A2(n13506), .ZN(n9103) );
  NAND2_X1 U11487 ( .A1(n9106), .A2(n9105), .ZN(n9107) );
  INV_X1 U11488 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n11984) );
  OR2_X1 U11489 ( .A1(n9110), .A2(n11984), .ZN(n9111) );
  INV_X1 U11490 ( .A(n9112), .ZN(n13564) );
  NAND2_X1 U11491 ( .A1(n9113), .A2(n13564), .ZN(n9144) );
  INV_X1 U11492 ( .A(n9571), .ZN(n9197) );
  AND2_X1 U11493 ( .A1(n9197), .A2(n6843), .ZN(n9562) );
  NAND2_X1 U11494 ( .A1(n13587), .A2(n10827), .ZN(n9476) );
  NAND2_X1 U11495 ( .A1(n9476), .A2(n6637), .ZN(n9114) );
  AOI21_X1 U11496 ( .B1(n9562), .B2(n10827), .A(n9114), .ZN(n9119) );
  NAND2_X1 U11497 ( .A1(n6651), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n9118) );
  NAND2_X1 U11498 ( .A1(n6860), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9117) );
  NAND2_X1 U11499 ( .A1(n9035), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9116) );
  AND3_X1 U11500 ( .A1(n9118), .A2(n9117), .A3(n9116), .ZN(n11827) );
  AOI21_X1 U11501 ( .B1(n9144), .B2(n9119), .A(n11827), .ZN(n9120) );
  NAND2_X1 U11502 ( .A1(n13569), .A2(n9113), .ZN(n9123) );
  OR2_X1 U11503 ( .A1(n9121), .A2(n11827), .ZN(n9122) );
  NAND2_X1 U11504 ( .A1(n9123), .A2(n9122), .ZN(n9139) );
  NAND2_X1 U11505 ( .A1(n9140), .A2(n9139), .ZN(n9142) );
  OR3_X1 U11506 ( .A1(n9126), .A2(n9125), .A3(n9124), .ZN(n9133) );
  INV_X1 U11507 ( .A(n9127), .ZN(n9130) );
  INV_X1 U11508 ( .A(n9128), .ZN(n9129) );
  NAND3_X1 U11509 ( .A1(n9131), .A2(n9130), .A3(n9129), .ZN(n9132) );
  OAI211_X1 U11510 ( .C1(n9135), .C2(n9134), .A(n9133), .B(n9132), .ZN(n9136)
         );
  INV_X1 U11511 ( .A(n9137), .ZN(n9138) );
  OAI22_X1 U11512 ( .A1(n9140), .A2(n9139), .B1(n6729), .B2(n9138), .ZN(n9141)
         );
  NAND3_X1 U11513 ( .A1(n6683), .A2(n9142), .A3(n9141), .ZN(n9148) );
  NAND2_X1 U11514 ( .A1(n9143), .A2(n13564), .ZN(n9146) );
  NAND2_X1 U11515 ( .A1(n9144), .A2(n9113), .ZN(n9145) );
  MUX2_X1 U11516 ( .A(n9146), .B(n9145), .S(n13566), .Z(n9147) );
  NAND2_X1 U11517 ( .A1(n9148), .A2(n9147), .ZN(n9149) );
  MUX2_X1 U11518 ( .A(n10899), .B(n9571), .S(n10827), .Z(n9156) );
  INV_X1 U11519 ( .A(n9151), .ZN(n9152) );
  INV_X1 U11520 ( .A(n9394), .ZN(n9155) );
  NAND2_X1 U11521 ( .A1(n9155), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11137) );
  NOR4_X2 U11522 ( .A1(n9181), .A2(n9156), .A3(n13587), .A4(n11137), .ZN(n9180) );
  XNOR2_X1 U11523 ( .A(n13569), .B(n11827), .ZN(n9176) );
  XNOR2_X1 U11524 ( .A(n13762), .B(n11972), .ZN(n11846) );
  XNOR2_X1 U11525 ( .A(n13773), .B(n13493), .ZN(n13602) );
  NAND2_X1 U11526 ( .A1(n13767), .A2(n13507), .ZN(n11845) );
  OR2_X1 U11527 ( .A1(n13767), .A2(n13507), .ZN(n9157) );
  NAND2_X1 U11528 ( .A1(n11845), .A2(n9157), .ZN(n11844) );
  OR2_X1 U11529 ( .A1(n13795), .A2(n13512), .ZN(n11841) );
  NAND2_X1 U11530 ( .A1(n13795), .A2(n13512), .ZN(n11842) );
  NAND2_X1 U11531 ( .A1(n11841), .A2(n11842), .ZN(n13651) );
  NAND2_X1 U11532 ( .A1(n13813), .A2(n9158), .ZN(n11821) );
  OR2_X1 U11533 ( .A1(n13813), .A2(n9158), .ZN(n9159) );
  NAND2_X1 U11534 ( .A1(n11821), .A2(n9159), .ZN(n13700) );
  OR2_X1 U11535 ( .A1(n13818), .A2(n13516), .ZN(n11836) );
  NAND2_X1 U11536 ( .A1(n13818), .A2(n13516), .ZN(n11835) );
  NAND2_X1 U11537 ( .A1(n11836), .A2(n11835), .ZN(n13713) );
  INV_X1 U11538 ( .A(n13518), .ZN(n13484) );
  XNOR2_X1 U11539 ( .A(n11923), .B(n13484), .ZN(n11585) );
  INV_X1 U11540 ( .A(n13519), .ZN(n11583) );
  XNOR2_X1 U11541 ( .A(n13750), .B(n11583), .ZN(n11571) );
  XNOR2_X1 U11542 ( .A(n14885), .B(n11577), .ZN(n11574) );
  XNOR2_X1 U11543 ( .A(n11170), .B(n10986), .ZN(n10988) );
  INV_X1 U11544 ( .A(n13522), .ZN(n10989) );
  XNOR2_X1 U11545 ( .A(n11238), .B(n10989), .ZN(n11008) );
  NAND2_X1 U11546 ( .A1(n15369), .A2(n13524), .ZN(n10764) );
  OR2_X1 U11547 ( .A1(n15369), .A2(n13524), .ZN(n9160) );
  NAND2_X1 U11548 ( .A1(n10764), .A2(n9160), .ZN(n10756) );
  XNOR2_X1 U11549 ( .A(n15347), .B(n10607), .ZN(n10599) );
  XNOR2_X1 U11550 ( .A(n10292), .B(n13528), .ZN(n10289) );
  INV_X1 U11551 ( .A(n8463), .ZN(n9473) );
  NAND2_X1 U11552 ( .A1(n9473), .A2(n9614), .ZN(n9475) );
  INV_X1 U11553 ( .A(n9161), .ZN(n9162) );
  AND2_X1 U11554 ( .A1(n9475), .A2(n9162), .ZN(n15308) );
  INV_X1 U11555 ( .A(n10827), .ZN(n9563) );
  NAND4_X1 U11556 ( .A1(n15308), .A2(n6890), .A3(n10198), .A4(n9563), .ZN(
        n9163) );
  INV_X1 U11557 ( .A(n13530), .ZN(n10208) );
  XNOR2_X1 U11558 ( .A(n15324), .B(n10208), .ZN(n10218) );
  NOR2_X1 U11559 ( .A1(n9163), .A2(n10218), .ZN(n9164) );
  XNOR2_X1 U11560 ( .A(n10239), .B(n13529), .ZN(n10236) );
  NAND4_X1 U11561 ( .A1(n10289), .A2(n9164), .A3(n10236), .A4(n10346), .ZN(
        n9165) );
  NOR2_X1 U11562 ( .A1(n10599), .A2(n9165), .ZN(n9166) );
  XNOR2_X1 U11563 ( .A(n10682), .B(n13526), .ZN(n10673) );
  XNOR2_X1 U11564 ( .A(n15361), .B(n13525), .ZN(n10730) );
  NAND4_X1 U11565 ( .A1(n10756), .A2(n9166), .A3(n10673), .A4(n10730), .ZN(
        n9167) );
  OR4_X1 U11566 ( .A1(n11574), .A2(n10988), .A3(n11008), .A4(n9167), .ZN(n9168) );
  INV_X1 U11567 ( .A(n13520), .ZN(n11581) );
  XNOR2_X1 U11568 ( .A(n14830), .B(n11581), .ZN(n14835) );
  INV_X1 U11569 ( .A(n13521), .ZN(n11579) );
  XNOR2_X1 U11570 ( .A(n14849), .B(n11579), .ZN(n14838) );
  OR4_X1 U11571 ( .A1(n11571), .A2(n9168), .A3(n14835), .A4(n14838), .ZN(n9169) );
  NOR2_X1 U11572 ( .A1(n11585), .A2(n9169), .ZN(n9170) );
  XNOR2_X1 U11573 ( .A(n13822), .B(n13517), .ZN(n13737) );
  NAND3_X1 U11574 ( .A1(n13713), .A2(n9170), .A3(n13737), .ZN(n9171) );
  NOR2_X1 U11575 ( .A1(n13700), .A2(n9171), .ZN(n9172) );
  XNOR2_X1 U11576 ( .A(n13804), .B(n13514), .ZN(n13686) );
  XNOR2_X1 U11577 ( .A(n13800), .B(n13513), .ZN(n13663) );
  NAND4_X1 U11578 ( .A1(n13651), .A2(n9172), .A3(n13686), .A4(n13663), .ZN(
        n9173) );
  NOR2_X1 U11579 ( .A1(n13645), .A2(n9173), .ZN(n9174) );
  XNOR2_X1 U11580 ( .A(n13779), .B(n13509), .ZN(n13610) );
  XNOR2_X1 U11581 ( .A(n13785), .B(n13510), .ZN(n13621) );
  NAND4_X1 U11582 ( .A1(n11844), .A2(n9174), .A3(n13610), .A4(n13621), .ZN(
        n9175) );
  NOR4_X1 U11583 ( .A1(n9176), .A2(n11846), .A3(n13602), .A4(n9175), .ZN(n9177) );
  NAND2_X1 U11584 ( .A1(n6683), .A2(n9177), .ZN(n9199) );
  INV_X1 U11585 ( .A(n11137), .ZN(n9184) );
  NAND4_X1 U11586 ( .A1(n9199), .A2(n6843), .A3(n9184), .A4(n10899), .ZN(n9178) );
  AOI21_X1 U11587 ( .B1(n9181), .B2(n10827), .A(n9178), .ZN(n9179) );
  NOR2_X1 U11588 ( .A1(n9180), .A2(n9179), .ZN(n9203) );
  NAND2_X1 U11589 ( .A1(n13587), .A2(n6637), .ZN(n9182) );
  OAI211_X1 U11590 ( .C1(n9197), .C2(n10184), .A(n9182), .B(n9476), .ZN(n9183)
         );
  NAND3_X1 U11591 ( .A1(n9181), .A2(n9184), .A3(n9183), .ZN(n9202) );
  NAND2_X1 U11592 ( .A1(n6785), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9186) );
  MUX2_X1 U11593 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9186), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n9189) );
  NAND2_X1 U11594 ( .A1(n9189), .A2(n9188), .ZN(n11350) );
  INV_X1 U11595 ( .A(n11350), .ZN(n9461) );
  NAND2_X1 U11596 ( .A1(n9188), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9190) );
  MUX2_X1 U11597 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9190), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n9191) );
  NAND3_X1 U11598 ( .A1(n9462), .A2(n9461), .A3(n9445), .ZN(n9204) );
  INV_X1 U11599 ( .A(n9193), .ZN(n9418) );
  INV_X1 U11600 ( .A(n9476), .ZN(n9195) );
  INV_X1 U11601 ( .A(n9469), .ZN(n9194) );
  AND2_X2 U11602 ( .A1(n9478), .A2(n9194), .ZN(n13475) );
  NAND4_X1 U11603 ( .A1(n15305), .A2(n9418), .A3(n9195), .A4(n13475), .ZN(
        n9196) );
  OAI211_X1 U11604 ( .C1(n9197), .C2(n11137), .A(n9196), .B(P2_B_REG_SCAN_IN), 
        .ZN(n9198) );
  INV_X1 U11605 ( .A(n9198), .ZN(n9200) );
  NAND3_X1 U11606 ( .A1(n9203), .A2(n9202), .A3(n9201), .ZN(P2_U3328) );
  INV_X1 U11607 ( .A(n9204), .ZN(n9205) );
  NOR2_X1 U11608 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n9207) );
  NOR2_X1 U11609 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n9206) );
  INV_X1 U11610 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9215) );
  NAND2_X1 U11611 ( .A1(n9248), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9218) );
  INV_X1 U11612 ( .A(n9278), .ZN(n9232) );
  NOR2_X1 U11613 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n9222) );
  INV_X1 U11614 ( .A(n9226), .ZN(n9223) );
  OAI21_X1 U11615 ( .B1(n6672), .B2(n9223), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9224) );
  MUX2_X1 U11616 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9224), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n9228) );
  NOR3_X1 U11617 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .A3(P1_IR_REG_25__SCAN_IN), .ZN(n9225) );
  NAND2_X1 U11618 ( .A1(n9226), .A2(n9225), .ZN(n9227) );
  NAND2_X1 U11619 ( .A1(n6669), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9229) );
  MUX2_X1 U11620 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9229), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n9231) );
  INV_X1 U11621 ( .A(n9236), .ZN(n9230) );
  INV_X2 U11622 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U11623 ( .A(n14254), .ZN(n11797) );
  INV_X1 U11624 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9239) );
  AOI21_X1 U11625 ( .B1(n11797), .B2(n9239), .A(n9266), .ZN(n9382) );
  NAND2_X1 U11626 ( .A1(n9244), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9241) );
  MUX2_X1 U11627 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9241), .S(
        P1_IR_REG_21__SCAN_IN), .Z(n9242) );
  NAND2_X1 U11628 ( .A1(n6672), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9243) );
  MUX2_X1 U11629 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9243), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n9245) );
  NAND2_X1 U11630 ( .A1(n9246), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9247) );
  NAND2_X1 U11631 ( .A1(n14007), .A2(n14195), .ZN(n10059) );
  NAND2_X1 U11632 ( .A1(n9251), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9252) );
  NAND2_X1 U11633 ( .A1(n9942), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n9263) );
  INV_X1 U11634 ( .A(n9259), .ZN(n11909) );
  NAND2_X1 U11635 ( .A1(n9954), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9262) );
  INV_X2 U11636 ( .A(n11800), .ZN(n11093) );
  NAND2_X1 U11637 ( .A1(n11093), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9261) );
  NAND2_X1 U11638 ( .A1(n11715), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9260) );
  NOR2_X1 U11639 ( .A1(n6832), .A2(n9333), .ZN(n9264) );
  XNOR2_X1 U11640 ( .A(n9264), .B(n6942), .ZN(n14700) );
  NAND2_X1 U11641 ( .A1(n11048), .A2(n10667), .ZN(n9268) );
  INV_X1 U11642 ( .A(n10529), .ZN(n9271) );
  NAND2_X1 U11643 ( .A1(n9268), .A2(n9267), .ZN(n9269) );
  OR2_X1 U11644 ( .A1(n10626), .A2(n12338), .ZN(n9273) );
  AOI22_X1 U11645 ( .A1(n12329), .A2(n10667), .B1(n9271), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n9272) );
  NAND2_X1 U11646 ( .A1(n9273), .A2(n9272), .ZN(n9836) );
  OAI21_X1 U11647 ( .B1(n9274), .B2(n9836), .A(n9835), .ZN(n9275) );
  INV_X1 U11648 ( .A(n9275), .ZN(n9872) );
  MUX2_X1 U11649 ( .A(n14290), .B(n9872), .S(n14254), .Z(n9276) );
  INV_X1 U11650 ( .A(n9266), .ZN(n9853) );
  NAND2_X1 U11651 ( .A1(n9276), .A2(n9853), .ZN(n9277) );
  OAI211_X1 U11652 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n9382), .A(n9277), .B(
        n14282), .ZN(n14307) );
  INV_X1 U11653 ( .A(n14307), .ZN(n9312) );
  INV_X1 U11654 ( .A(n9846), .ZN(n9820) );
  INV_X1 U11655 ( .A(n9587), .ZN(n9279) );
  NAND2_X1 U11656 ( .A1(n9279), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14258) );
  NAND2_X1 U11657 ( .A1(n9820), .A2(n14258), .ZN(n9299) );
  INV_X1 U11658 ( .A(n14195), .ZN(n9977) );
  INV_X1 U11659 ( .A(n14022), .ZN(n9854) );
  NAND2_X1 U11660 ( .A1(n9854), .A2(n9587), .ZN(n9280) );
  NAND2_X1 U11661 ( .A1(n9280), .A2(n6845), .ZN(n9298) );
  INV_X1 U11662 ( .A(n9298), .ZN(n9281) );
  AND2_X1 U11663 ( .A1(n9299), .A2(n9281), .ZN(n9385) );
  OR2_X1 U11664 ( .A1(n9266), .A2(n14254), .ZN(n9282) );
  OR2_X1 U11665 ( .A1(n9301), .A2(n9282), .ZN(n15061) );
  NAND2_X1 U11666 ( .A1(n9283), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9285) );
  XNOR2_X1 U11667 ( .A(n9285), .B(n9284), .ZN(n9963) );
  XNOR2_X1 U11668 ( .A(n9963), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n9296) );
  INV_X1 U11669 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10629) );
  INV_X1 U11670 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n9286) );
  INV_X1 U11671 ( .A(n9802), .ZN(n14285) );
  NAND2_X1 U11672 ( .A1(n14285), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9287) );
  NAND2_X1 U11673 ( .A1(n14289), .A2(n9287), .ZN(n14299) );
  INV_X1 U11674 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n15113) );
  MUX2_X1 U11675 ( .A(n15113), .B(P1_REG2_REG_2__SCAN_IN), .S(n11619), .Z(
        n14300) );
  NAND2_X1 U11676 ( .A1(n14299), .A2(n14300), .ZN(n14298) );
  INV_X1 U11677 ( .A(n11619), .ZN(n14297) );
  NAND2_X1 U11678 ( .A1(n14297), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9291) );
  NAND2_X1 U11679 ( .A1(n14298), .A2(n9291), .ZN(n14314) );
  XNOR2_X1 U11680 ( .A(n9292), .B(n9209), .ZN(n14308) );
  XNOR2_X1 U11681 ( .A(n14308), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n14315) );
  NAND2_X1 U11682 ( .A1(n14314), .A2(n14315), .ZN(n14313) );
  INV_X1 U11683 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n9293) );
  OR2_X1 U11684 ( .A1(n14308), .A2(n9293), .ZN(n9294) );
  NAND2_X1 U11685 ( .A1(n14313), .A2(n9294), .ZN(n9295) );
  NAND2_X1 U11686 ( .A1(n9295), .A2(n9296), .ZN(n9734) );
  OAI21_X1 U11687 ( .B1(n9296), .B2(n9295), .A(n9734), .ZN(n9297) );
  NOR2_X1 U11688 ( .A1(n15061), .A2(n9297), .ZN(n9311) );
  INV_X1 U11689 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9300) );
  NAND2_X1 U11690 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n10535) );
  OAI21_X1 U11691 ( .B1(n15104), .B2(n9300), .A(n10535), .ZN(n9310) );
  XNOR2_X1 U11692 ( .A(n9963), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n9307) );
  INV_X1 U11693 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n15195) );
  MUX2_X1 U11694 ( .A(n15195), .B(P1_REG1_REG_1__SCAN_IN), .S(n9802), .Z(
        n14288) );
  AND2_X1 U11695 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n14287) );
  NAND2_X1 U11696 ( .A1(n14288), .A2(n14287), .ZN(n14286) );
  NAND2_X1 U11697 ( .A1(n14285), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9302) );
  NAND2_X1 U11698 ( .A1(n14286), .A2(n9302), .ZN(n14302) );
  INV_X1 U11699 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n15197) );
  MUX2_X1 U11700 ( .A(n15197), .B(P1_REG1_REG_2__SCAN_IN), .S(n11619), .Z(
        n14303) );
  NAND2_X1 U11701 ( .A1(n14302), .A2(n14303), .ZN(n14301) );
  NAND2_X1 U11702 ( .A1(n14297), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9303) );
  NAND2_X1 U11703 ( .A1(n14301), .A2(n9303), .ZN(n14317) );
  XNOR2_X1 U11704 ( .A(n14308), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n14318) );
  NAND2_X1 U11705 ( .A1(n14317), .A2(n14318), .ZN(n14316) );
  INV_X1 U11706 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9304) );
  OR2_X1 U11707 ( .A1(n14308), .A2(n9304), .ZN(n9305) );
  NAND2_X1 U11708 ( .A1(n14316), .A2(n9305), .ZN(n9306) );
  NAND2_X1 U11709 ( .A1(n9306), .A2(n9307), .ZN(n9725) );
  OAI211_X1 U11710 ( .C1(n9307), .C2(n9306), .A(n15091), .B(n9725), .ZN(n9308)
         );
  OAI21_X1 U11711 ( .B1(n15100), .B2(n9963), .A(n9308), .ZN(n9309) );
  OR4_X1 U11712 ( .A1(n9312), .A2(n9311), .A3(n9310), .A4(n9309), .ZN(P1_U3247) );
  NOR2_X1 U11713 ( .A1(n6832), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13381) );
  AOI222_X1 U11714 ( .A1(n9313), .A2(n13381), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10168), .C1(SI_5_), .C2(n13380), .ZN(n9314) );
  INV_X1 U11715 ( .A(n9314), .ZN(P3_U3290) );
  AOI222_X1 U11716 ( .A1(n9315), .A2(n13381), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10405), .C1(SI_4_), .C2(n13380), .ZN(n9316) );
  INV_X1 U11717 ( .A(n9316), .ZN(P3_U3291) );
  INV_X2 U11718 ( .A(n13380), .ZN(n14721) );
  INV_X1 U11719 ( .A(SI_7_), .ZN(n9319) );
  INV_X2 U11720 ( .A(n13381), .ZN(n14722) );
  INV_X1 U11721 ( .A(n9317), .ZN(n9318) );
  OAI222_X1 U11722 ( .A1(P3_U3151), .A2(n10502), .B1(n14721), .B2(n9319), .C1(
        n14722), .C2(n9318), .ZN(P3_U3288) );
  OAI222_X1 U11723 ( .A1(n14722), .A2(n9321), .B1(n14721), .B2(n9320), .C1(
        P3_U3151), .C2(n10928), .ZN(P3_U3287) );
  OAI222_X1 U11724 ( .A1(n14722), .A2(n9323), .B1(n14721), .B2(n9322), .C1(
        P3_U3151), .C2(n10253), .ZN(P3_U3294) );
  INV_X1 U11725 ( .A(SI_9_), .ZN(n9326) );
  INV_X1 U11726 ( .A(n9324), .ZN(n9325) );
  OAI222_X1 U11727 ( .A1(P3_U3151), .A2(n10929), .B1(n14721), .B2(n9326), .C1(
        n14722), .C2(n9325), .ZN(P3_U3286) );
  NOR2_X1 U11728 ( .A1(n8991), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13848) );
  INV_X2 U11729 ( .A(n13848), .ZN(n13852) );
  NAND2_X2 U11730 ( .A1(n8991), .A2(P2_U3088), .ZN(n13854) );
  OAI222_X1 U11731 ( .A1(n13852), .A2(n9327), .B1(n13854), .B2(n9959), .C1(
        P2_U3088), .C2(n9434), .ZN(P2_U3323) );
  INV_X1 U11732 ( .A(n6641), .ZN(n10163) );
  INV_X1 U11733 ( .A(n9328), .ZN(n9330) );
  OAI222_X1 U11734 ( .A1(n10163), .A2(P3_U3151), .B1(n14722), .B2(n9330), .C1(
        n9329), .C2(n14721), .ZN(P3_U3293) );
  OAI222_X1 U11735 ( .A1(P3_U3151), .A2(n10458), .B1(n14722), .B2(n9332), .C1(
        n9331), .C2(n14721), .ZN(P3_U3289) );
  OAI222_X1 U11736 ( .A1(P3_U3151), .A2(n9335), .B1(n14722), .B2(n9334), .C1(
        n9333), .C2(n14721), .ZN(P3_U3295) );
  NAND2_X2 U11737 ( .A1(n6832), .A2(P1_U3086), .ZN(n14694) );
  INV_X1 U11738 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9960) );
  NOR2_X1 U11739 ( .A1(n6832), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14691) );
  OAI222_X1 U11740 ( .A1(n14694), .A2(n9960), .B1(n11910), .B2(n9959), .C1(
        P1_U3086), .C2(n9963), .ZN(P1_U3351) );
  INV_X1 U11741 ( .A(n9338), .ZN(n9339) );
  OAI222_X1 U11742 ( .A1(P3_U3151), .A2(n15417), .B1(n14721), .B2(n9340), .C1(
        n14722), .C2(n9339), .ZN(P3_U3285) );
  INV_X1 U11743 ( .A(n9341), .ZN(n10321) );
  INV_X1 U11744 ( .A(n9519), .ZN(n9443) );
  OAI222_X1 U11745 ( .A1(n13852), .A2(n9342), .B1(n13854), .B2(n10321), .C1(
        P2_U3088), .C2(n9443), .ZN(P2_U3322) );
  NOR2_X1 U11746 ( .A1(n9283), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n9352) );
  OR2_X1 U11747 ( .A1(n9352), .A2(n9233), .ZN(n9343) );
  XNOR2_X1 U11748 ( .A(n9343), .B(n9351), .ZN(n10324) );
  OAI222_X1 U11749 ( .A1(n14694), .A2(n6913), .B1(n11910), .B2(n10321), .C1(
        P1_U3086), .C2(n10324), .ZN(P1_U3350) );
  INV_X1 U11750 ( .A(n9344), .ZN(n9948) );
  OAI222_X1 U11751 ( .A1(n14694), .A2(n7036), .B1(n11910), .B2(n9948), .C1(
        P1_U3086), .C2(n14308), .ZN(P1_U3352) );
  INV_X1 U11752 ( .A(n9496), .ZN(n9503) );
  OAI222_X1 U11753 ( .A1(n13852), .A2(n9345), .B1(n13854), .B2(n9948), .C1(
        P2_U3088), .C2(n9503), .ZN(P2_U3324) );
  OAI222_X1 U11754 ( .A1(n11910), .A2(n9801), .B1(n9802), .B2(P1_U3086), .C1(
        n6944), .C2(n14694), .ZN(P1_U3354) );
  INV_X1 U11755 ( .A(SI_11_), .ZN(n9348) );
  INV_X1 U11756 ( .A(n9346), .ZN(n9347) );
  OAI222_X1 U11757 ( .A1(P3_U3151), .A2(n11268), .B1(n14721), .B2(n9348), .C1(
        n14722), .C2(n9347), .ZN(P3_U3284) );
  OAI222_X1 U11758 ( .A1(P2_U3088), .A2(n15203), .B1(n13854), .B2(n9801), .C1(
        n9349), .C2(n13852), .ZN(P2_U3326) );
  INV_X1 U11759 ( .A(n10551), .ZN(n9355) );
  INV_X1 U11760 ( .A(n9594), .ZN(n9605) );
  OAI222_X1 U11761 ( .A1(n13852), .A2(n9350), .B1(n13854), .B2(n9355), .C1(
        P2_U3088), .C2(n9605), .ZN(P2_U3321) );
  NAND2_X1 U11762 ( .A1(n9352), .A2(n9351), .ZN(n9356) );
  NAND2_X1 U11763 ( .A1(n9356), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9354) );
  XNOR2_X1 U11764 ( .A(n9354), .B(n9353), .ZN(n10555) );
  OAI222_X1 U11765 ( .A1(n14694), .A2(n10552), .B1(n11910), .B2(n9355), .C1(
        P1_U3086), .C2(n10555), .ZN(P1_U3349) );
  INV_X1 U11766 ( .A(n10799), .ZN(n9360) );
  NAND2_X1 U11767 ( .A1(n9363), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9357) );
  XNOR2_X1 U11768 ( .A(n9357), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10800) );
  INV_X1 U11769 ( .A(n14694), .ZN(n9380) );
  AOI22_X1 U11770 ( .A1(n10800), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n9380), .ZN(n9358) );
  OAI21_X1 U11771 ( .B1(n9360), .B2(n11910), .A(n9358), .ZN(P1_U3348) );
  INV_X1 U11772 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9361) );
  INV_X1 U11773 ( .A(n13554), .ZN(n9359) );
  OAI222_X1 U11774 ( .A1(n13852), .A2(n9361), .B1(n13854), .B2(n9360), .C1(
        P2_U3088), .C2(n9359), .ZN(P2_U3320) );
  NAND2_X1 U11775 ( .A1(n11567), .A2(P2_U3947), .ZN(n9362) );
  OAI21_X1 U11776 ( .B1(n8719), .B2(P2_U3947), .A(n9362), .ZN(P2_U3544) );
  INV_X1 U11777 ( .A(n10852), .ZN(n9371) );
  NAND2_X1 U11778 ( .A1(n9368), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9364) );
  XNOR2_X1 U11779 ( .A(n9364), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10853) );
  AOI22_X1 U11780 ( .A1(n10853), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9380), .ZN(n9365) );
  OAI21_X1 U11781 ( .B1(n9371), .B2(n11910), .A(n9365), .ZN(P1_U3347) );
  OAI222_X1 U11782 ( .A1(n14721), .A2(n9367), .B1(n14722), .B2(n9366), .C1(
        n11892), .C2(P3_U3151), .ZN(P3_U3283) );
  OR2_X1 U11783 ( .A1(n9550), .A2(n7537), .ZN(n9369) );
  NAND2_X1 U11784 ( .A1(n9550), .A2(n7537), .ZN(n9378) );
  INV_X1 U11785 ( .A(n11080), .ZN(n9370) );
  OAI222_X1 U11786 ( .A1(n11910), .A2(n11079), .B1(n9370), .B2(P1_U3086), .C1(
        n13149), .C2(n14694), .ZN(P1_U3346) );
  INV_X1 U11787 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9372) );
  INV_X1 U11788 ( .A(n9528), .ZN(n9665) );
  OAI222_X1 U11789 ( .A1(n13852), .A2(n9372), .B1(n13854), .B2(n9371), .C1(
        P2_U3088), .C2(n9665), .ZN(P2_U3319) );
  INV_X1 U11790 ( .A(n9629), .ZN(n9636) );
  OAI222_X1 U11791 ( .A1(P2_U3088), .A2(n9636), .B1(n13854), .B2(n11079), .C1(
        n9373), .C2(n13852), .ZN(P2_U3318) );
  INV_X1 U11792 ( .A(n12564), .ZN(n11894) );
  OAI222_X1 U11793 ( .A1(n14721), .A2(n9375), .B1(n14722), .B2(n9374), .C1(
        n11894), .C2(P3_U3151), .ZN(P3_U3282) );
  OAI222_X1 U11794 ( .A1(P3_U3151), .A2(n12578), .B1(n14721), .B2(n9377), .C1(
        n14722), .C2(n9376), .ZN(P3_U3281) );
  INV_X1 U11795 ( .A(n11071), .ZN(n9390) );
  NAND2_X1 U11796 ( .A1(n9378), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9379) );
  XNOR2_X1 U11797 ( .A(n9379), .B(P1_IR_REG_10__SCAN_IN), .ZN(n11072) );
  AOI22_X1 U11798 ( .A1(n11072), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9380), .ZN(n9381) );
  OAI21_X1 U11799 ( .B1(n9390), .B2(n11910), .A(n9381), .ZN(P1_U3345) );
  OAI21_X1 U11800 ( .B1(n11797), .B2(P1_REG1_REG_0__SCAN_IN), .A(n9382), .ZN(
        n9383) );
  XNOR2_X1 U11801 ( .A(n9383), .B(P1_IR_REG_0__SCAN_IN), .ZN(n9384) );
  AOI22_X1 U11802 ( .A1(n9385), .A2(n9384), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n9386) );
  OAI21_X1 U11803 ( .B1(n15104), .B2(n8351), .A(n9386), .ZN(P1_U3243) );
  AND2_X1 U11804 ( .A1(n9391), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U11805 ( .A1(n9391), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U11806 ( .A1(n9391), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U11807 ( .A1(n9391), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U11808 ( .A1(n9391), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U11809 ( .A1(n9391), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U11810 ( .A1(n9391), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U11811 ( .A1(n9391), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U11812 ( .A1(n9391), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U11813 ( .A1(n9391), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U11814 ( .A1(n9391), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U11815 ( .A1(n9391), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U11816 ( .A1(n9391), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U11817 ( .A1(n9391), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U11818 ( .A1(n9391), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U11819 ( .A1(n9391), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U11820 ( .A1(n9391), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U11821 ( .A1(n9391), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U11822 ( .A1(n9391), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U11823 ( .A1(n9391), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U11824 ( .A1(n9391), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U11825 ( .A1(n9391), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U11826 ( .A1(n9391), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U11827 ( .A1(n9391), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U11828 ( .A1(n9391), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  INV_X1 U11829 ( .A(n9533), .ZN(n15218) );
  INV_X1 U11830 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9389) );
  OAI222_X1 U11831 ( .A1(P2_U3088), .A2(n15218), .B1(n13854), .B2(n9390), .C1(
        n9389), .C2(n13852), .ZN(P2_U3317) );
  INV_X1 U11832 ( .A(n9391), .ZN(n9393) );
  INV_X1 U11833 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n13151) );
  NOR2_X1 U11834 ( .A1(n9393), .A2(n13151), .ZN(P3_U3263) );
  INV_X1 U11835 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n9392) );
  NOR2_X1 U11836 ( .A1(n9393), .A2(n9392), .ZN(P3_U3255) );
  INV_X1 U11837 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n13217) );
  NOR2_X1 U11838 ( .A1(n9393), .A2(n13217), .ZN(P3_U3240) );
  INV_X1 U11839 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n13292) );
  NOR2_X1 U11840 ( .A1(n9393), .A2(n13292), .ZN(P3_U3254) );
  INV_X1 U11841 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n13208) );
  NOR2_X1 U11842 ( .A1(n9393), .A2(n13208), .ZN(P3_U3262) );
  AOI21_X1 U11843 ( .B1(n9478), .B2(n9394), .A(n6643), .ZN(n9396) );
  OR2_X1 U11844 ( .A1(n9396), .A2(n9395), .ZN(n9408) );
  NAND2_X1 U11845 ( .A1(n9408), .A2(n9469), .ZN(n15204) );
  NOR2_X1 U11846 ( .A1(n9469), .A2(P2_U3088), .ZN(n13847) );
  NAND2_X1 U11847 ( .A1(n9408), .A2(n13847), .ZN(n9417) );
  OR2_X1 U11848 ( .A1(n9417), .A2(n9418), .ZN(n15225) );
  INV_X1 U11849 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9397) );
  MUX2_X1 U11850 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n9397), .S(n9496), .Z(n9402)
         );
  XNOR2_X1 U11851 ( .A(n15203), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n15211) );
  AND2_X1 U11852 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n15210) );
  NAND2_X1 U11853 ( .A1(n15211), .A2(n15210), .ZN(n15209) );
  INV_X1 U11854 ( .A(n15203), .ZN(n9410) );
  NAND2_X1 U11855 ( .A1(n9410), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9398) );
  NAND2_X1 U11856 ( .A1(n15209), .A2(n9398), .ZN(n13535) );
  XNOR2_X1 U11857 ( .A(n13538), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n13536) );
  NAND2_X1 U11858 ( .A1(n13535), .A2(n13536), .ZN(n9401) );
  INV_X1 U11859 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9399) );
  OR2_X1 U11860 ( .A1(n13538), .A2(n9399), .ZN(n9400) );
  NAND2_X1 U11861 ( .A1(n9401), .A2(n9400), .ZN(n9489) );
  NAND2_X1 U11862 ( .A1(n9402), .A2(n9489), .ZN(n9490) );
  NAND2_X1 U11863 ( .A1(n9496), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9406) );
  NAND2_X1 U11864 ( .A1(n9490), .A2(n9406), .ZN(n9404) );
  INV_X1 U11865 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9426) );
  MUX2_X1 U11866 ( .A(n9426), .B(P2_REG1_REG_4__SCAN_IN), .S(n9434), .Z(n9403)
         );
  NAND2_X1 U11867 ( .A1(n9404), .A2(n9403), .ZN(n9432) );
  MUX2_X1 U11868 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n9426), .S(n9434), .Z(n9405)
         );
  NAND3_X1 U11869 ( .A1(n9490), .A2(n9406), .A3(n9405), .ZN(n9407) );
  NAND3_X1 U11870 ( .A1(n15264), .A2(n9432), .A3(n9407), .ZN(n9425) );
  OR2_X1 U11871 ( .A1(n9408), .A2(P2_U3088), .ZN(n15250) );
  INV_X1 U11872 ( .A(n15250), .ZN(n15270) );
  NAND2_X1 U11873 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n9794) );
  INV_X1 U11874 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9409) );
  MUX2_X1 U11875 ( .A(n9409), .B(P2_REG2_REG_1__SCAN_IN), .S(n15203), .Z(
        n15207) );
  AND2_X1 U11876 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n15208) );
  NAND2_X1 U11877 ( .A1(n15207), .A2(n15208), .ZN(n15206) );
  NAND2_X1 U11878 ( .A1(n9410), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n13540) );
  NAND2_X1 U11879 ( .A1(n15206), .A2(n13540), .ZN(n9412) );
  INV_X1 U11880 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9413) );
  MUX2_X1 U11881 ( .A(n9413), .B(P2_REG2_REG_2__SCAN_IN), .S(n13538), .Z(n9411) );
  NAND2_X1 U11882 ( .A1(n9412), .A2(n9411), .ZN(n13542) );
  OR2_X1 U11883 ( .A1(n13538), .A2(n9413), .ZN(n9498) );
  NAND2_X1 U11884 ( .A1(n13542), .A2(n9498), .ZN(n9415) );
  INV_X1 U11885 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10354) );
  MUX2_X1 U11886 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10354), .S(n9496), .Z(n9414) );
  NAND2_X1 U11887 ( .A1(n9415), .A2(n9414), .ZN(n9500) );
  NAND2_X1 U11888 ( .A1(n9496), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9416) );
  NAND2_X1 U11889 ( .A1(n9500), .A2(n9416), .ZN(n9421) );
  INV_X1 U11890 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10224) );
  MUX2_X1 U11891 ( .A(n10224), .B(P2_REG2_REG_4__SCAN_IN), .S(n9434), .Z(n9420) );
  INV_X1 U11892 ( .A(n9417), .ZN(n9419) );
  NAND2_X1 U11893 ( .A1(n9421), .A2(n9420), .ZN(n9436) );
  OAI211_X1 U11894 ( .C1(n9421), .C2(n9420), .A(n15271), .B(n9436), .ZN(n9422)
         );
  NAND2_X1 U11895 ( .A1(n9794), .A2(n9422), .ZN(n9423) );
  AOI21_X1 U11896 ( .B1(n15270), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n9423), .ZN(
        n9424) );
  OAI211_X1 U11897 ( .C1(n15278), .C2(n9434), .A(n9425), .B(n9424), .ZN(
        P2_U3218) );
  OR2_X1 U11898 ( .A1(n9434), .A2(n9426), .ZN(n9431) );
  NAND2_X1 U11899 ( .A1(n9432), .A2(n9431), .ZN(n9429) );
  INV_X1 U11900 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9427) );
  MUX2_X1 U11901 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n9427), .S(n9519), .Z(n9428)
         );
  NAND2_X1 U11902 ( .A1(n9429), .A2(n9428), .ZN(n9521) );
  MUX2_X1 U11903 ( .A(n9427), .B(P2_REG1_REG_5__SCAN_IN), .S(n9519), .Z(n9430)
         );
  NAND3_X1 U11904 ( .A1(n9432), .A2(n9431), .A3(n9430), .ZN(n9433) );
  NAND3_X1 U11905 ( .A1(n15264), .A2(n9521), .A3(n9433), .ZN(n9442) );
  NAND2_X1 U11906 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n9925) );
  OR2_X1 U11907 ( .A1(n9434), .A2(n10224), .ZN(n9435) );
  NAND2_X1 U11908 ( .A1(n9436), .A2(n9435), .ZN(n9438) );
  INV_X1 U11909 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10214) );
  MUX2_X1 U11910 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10214), .S(n9519), .Z(n9437) );
  NAND2_X1 U11911 ( .A1(n9438), .A2(n9437), .ZN(n9597) );
  OAI211_X1 U11912 ( .C1(n9438), .C2(n9437), .A(n15271), .B(n9597), .ZN(n9439)
         );
  NAND2_X1 U11913 ( .A1(n9925), .A2(n9439), .ZN(n9440) );
  AOI21_X1 U11914 ( .B1(n15270), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n9440), .ZN(
        n9441) );
  OAI211_X1 U11915 ( .C1(n15278), .C2(n9443), .A(n9442), .B(n9441), .ZN(
        P2_U3219) );
  INV_X1 U11916 ( .A(n9717), .ZN(n15246) );
  INV_X1 U11917 ( .A(n11382), .ZN(n9487) );
  OAI222_X1 U11918 ( .A1(P2_U3088), .A2(n15246), .B1(n13854), .B2(n9487), .C1(
        n9444), .C2(n13852), .ZN(P2_U3315) );
  INV_X1 U11919 ( .A(n9445), .ZN(n11469) );
  XNOR2_X1 U11920 ( .A(n11350), .B(P2_B_REG_SCAN_IN), .ZN(n9446) );
  NAND2_X1 U11921 ( .A1(n11469), .A2(n9446), .ZN(n9447) );
  AND2_X1 U11922 ( .A1(n9447), .A2(n9462), .ZN(n15293) );
  INV_X1 U11923 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15303) );
  NAND2_X1 U11924 ( .A1(n15293), .A2(n15303), .ZN(n9449) );
  INV_X1 U11925 ( .A(n9462), .ZN(n13855) );
  NAND2_X1 U11926 ( .A1(n13855), .A2(n11469), .ZN(n9448) );
  NAND2_X1 U11927 ( .A1(n9449), .A2(n9448), .ZN(n15304) );
  NOR4_X1 U11928 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n9453) );
  NOR4_X1 U11929 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n9452) );
  NOR4_X1 U11930 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9451) );
  NOR4_X1 U11931 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n9450) );
  AND4_X1 U11932 ( .A1(n9453), .A2(n9452), .A3(n9451), .A4(n9450), .ZN(n9459)
         );
  NOR2_X1 U11933 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .ZN(
        n9457) );
  NOR4_X1 U11934 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n9456) );
  NOR4_X1 U11935 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n9455) );
  NOR4_X1 U11936 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n9454) );
  AND4_X1 U11937 ( .A1(n9457), .A2(n9456), .A3(n9455), .A4(n9454), .ZN(n9458)
         );
  NAND2_X1 U11938 ( .A1(n9459), .A2(n9458), .ZN(n9460) );
  AND2_X1 U11939 ( .A1(n15293), .A2(n9460), .ZN(n9576) );
  NOR2_X1 U11940 ( .A1(n15304), .A2(n9576), .ZN(n10182) );
  INV_X1 U11941 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15299) );
  NAND2_X1 U11942 ( .A1(n15293), .A2(n15299), .ZN(n9464) );
  NOR2_X1 U11943 ( .A1(n9462), .A2(n9461), .ZN(n15300) );
  INV_X1 U11944 ( .A(n15300), .ZN(n9463) );
  AND2_X1 U11945 ( .A1(n9464), .A2(n9463), .ZN(n11019) );
  NAND2_X1 U11946 ( .A1(n10182), .A2(n11019), .ZN(n9465) );
  NAND2_X1 U11947 ( .A1(n9579), .A2(n9465), .ZN(n9468) );
  NAND2_X1 U11948 ( .A1(n9478), .A2(n9476), .ZN(n9580) );
  AND2_X1 U11949 ( .A1(n9466), .A2(n9580), .ZN(n9467) );
  NAND2_X1 U11950 ( .A1(n9468), .A2(n9467), .ZN(n9694) );
  OR2_X1 U11951 ( .A1(n9694), .A2(P2_U3088), .ZN(n9676) );
  INV_X1 U11952 ( .A(n9676), .ZN(n9483) );
  INV_X1 U11953 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n11626) );
  NAND3_X1 U11954 ( .A1(n15305), .A2(n11019), .A3(n10182), .ZN(n9479) );
  INV_X1 U11955 ( .A(n13476), .ZN(n13496) );
  OR2_X1 U11956 ( .A1(n13492), .A2(n9646), .ZN(n11623) );
  INV_X1 U11957 ( .A(n11623), .ZN(n9472) );
  INV_X1 U11958 ( .A(n9477), .ZN(n15306) );
  OR2_X1 U11959 ( .A1(n15306), .A2(n10827), .ZN(n14825) );
  OR2_X1 U11960 ( .A1(n9479), .A2(n14825), .ZN(n9471) );
  INV_X1 U11961 ( .A(n9579), .ZN(n9470) );
  AOI22_X1 U11962 ( .A1(n13496), .A2(n9472), .B1(n13501), .B2(n9614), .ZN(
        n9482) );
  NOR2_X1 U11963 ( .A1(n11966), .A2(n9473), .ZN(n9474) );
  MUX2_X1 U11964 ( .A(n11966), .B(n9474), .S(n15307), .Z(n9480) );
  INV_X1 U11965 ( .A(n9475), .ZN(n9643) );
  OAI21_X1 U11966 ( .B1(n9480), .B2(n9643), .A(n13454), .ZN(n9481) );
  OAI211_X1 U11967 ( .C1(n9483), .C2(n11626), .A(n9482), .B(n9481), .ZN(
        P2_U3204) );
  OR2_X1 U11968 ( .A1(n9485), .A2(n9233), .ZN(n9486) );
  NAND2_X1 U11969 ( .A1(n9550), .A2(n9486), .ZN(n9608) );
  XNOR2_X1 U11970 ( .A(n9484), .B(n9608), .ZN(n14337) );
  INV_X1 U11971 ( .A(n14337), .ZN(n10048) );
  OAI222_X1 U11972 ( .A1(n14694), .A2(n9488), .B1(P1_U3086), .B2(n10048), .C1(
        n9487), .C2(n11910), .ZN(P1_U3343) );
  NAND2_X1 U11973 ( .A1(P2_U3088), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n9697) );
  INV_X1 U11974 ( .A(n9697), .ZN(n9495) );
  INV_X1 U11975 ( .A(n9489), .ZN(n9493) );
  MUX2_X1 U11976 ( .A(n9397), .B(P2_REG1_REG_3__SCAN_IN), .S(n9496), .Z(n9492)
         );
  INV_X1 U11977 ( .A(n9490), .ZN(n9491) );
  AOI211_X1 U11978 ( .C1(n9493), .C2(n9492), .A(n9491), .B(n15225), .ZN(n9494)
         );
  AOI211_X1 U11979 ( .C1(n15270), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n9495), .B(
        n9494), .ZN(n9502) );
  MUX2_X1 U11980 ( .A(n10354), .B(P2_REG2_REG_3__SCAN_IN), .S(n9496), .Z(n9497) );
  NAND3_X1 U11981 ( .A1(n13542), .A2(n9498), .A3(n9497), .ZN(n9499) );
  NAND3_X1 U11982 ( .A1(n15271), .A2(n9500), .A3(n9499), .ZN(n9501) );
  OAI211_X1 U11983 ( .C1(n15278), .C2(n9503), .A(n9502), .B(n9501), .ZN(
        P2_U3217) );
  NAND2_X1 U11984 ( .A1(n9519), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9596) );
  NAND2_X1 U11985 ( .A1(n9597), .A2(n9596), .ZN(n9505) );
  INV_X1 U11986 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10244) );
  MUX2_X1 U11987 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10244), .S(n9594), .Z(n9504) );
  NAND2_X1 U11988 ( .A1(n9505), .A2(n9504), .ZN(n13557) );
  NAND2_X1 U11989 ( .A1(n9594), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n13556) );
  NAND2_X1 U11990 ( .A1(n13557), .A2(n13556), .ZN(n9507) );
  INV_X1 U11991 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10297) );
  MUX2_X1 U11992 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10297), .S(n13554), .Z(
        n9506) );
  NAND2_X1 U11993 ( .A1(n9507), .A2(n9506), .ZN(n13559) );
  NAND2_X1 U11994 ( .A1(n13554), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9508) );
  NAND2_X1 U11995 ( .A1(n13559), .A2(n9508), .ZN(n9659) );
  INV_X1 U11996 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10678) );
  MUX2_X1 U11997 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10678), .S(n9528), .Z(n9658) );
  NAND2_X1 U11998 ( .A1(n9659), .A2(n9658), .ZN(n9657) );
  NAND2_X1 U11999 ( .A1(n9528), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9509) );
  NAND2_X1 U12000 ( .A1(n9657), .A2(n9509), .ZN(n9625) );
  INV_X1 U12001 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n9624) );
  MUX2_X1 U12002 ( .A(n9624), .B(P2_REG2_REG_9__SCAN_IN), .S(n9629), .Z(n9510)
         );
  OR2_X1 U12003 ( .A1(n9625), .A2(n9510), .ZN(n9627) );
  OR2_X1 U12004 ( .A1(n9629), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n9511) );
  NAND2_X1 U12005 ( .A1(n9627), .A2(n9511), .ZN(n15221) );
  INV_X1 U12006 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n9512) );
  MUX2_X1 U12007 ( .A(n9512), .B(P2_REG2_REG_10__SCAN_IN), .S(n9533), .Z(
        n15222) );
  OR2_X1 U12008 ( .A1(n15221), .A2(n15222), .ZN(n15223) );
  NAND2_X1 U12009 ( .A1(n9533), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n9513) );
  NAND2_X1 U12010 ( .A1(n15223), .A2(n9513), .ZN(n9517) );
  INV_X1 U12011 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n9514) );
  MUX2_X1 U12012 ( .A(n9514), .B(P2_REG2_REG_11__SCAN_IN), .S(n9714), .Z(n9516) );
  INV_X1 U12013 ( .A(n15236), .ZN(n9515) );
  AOI21_X1 U12014 ( .B1(n9517), .B2(n9516), .A(n9515), .ZN(n9542) );
  INV_X1 U12015 ( .A(n15271), .ZN(n15220) );
  AND2_X1 U12016 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n11168) );
  INV_X1 U12017 ( .A(n9714), .ZN(n9553) );
  NOR2_X1 U12018 ( .A1(n15278), .A2(n9553), .ZN(n9518) );
  AOI211_X1 U12019 ( .C1(n15270), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n11168), 
        .B(n9518), .ZN(n9541) );
  NAND2_X1 U12020 ( .A1(n9519), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9520) );
  NAND2_X1 U12021 ( .A1(n9521), .A2(n9520), .ZN(n9600) );
  INV_X1 U12022 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9522) );
  MUX2_X1 U12023 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n9522), .S(n9594), .Z(n9599)
         );
  NAND2_X1 U12024 ( .A1(n9600), .A2(n9599), .ZN(n13551) );
  NAND2_X1 U12025 ( .A1(n9594), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n13550) );
  NAND2_X1 U12026 ( .A1(n13551), .A2(n13550), .ZN(n9525) );
  INV_X1 U12027 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9523) );
  MUX2_X1 U12028 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n9523), .S(n13554), .Z(n9524) );
  NAND2_X1 U12029 ( .A1(n9525), .A2(n9524), .ZN(n13553) );
  NAND2_X1 U12030 ( .A1(n13554), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9526) );
  NAND2_X1 U12031 ( .A1(n13553), .A2(n9526), .ZN(n9656) );
  INV_X1 U12032 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9527) );
  MUX2_X1 U12033 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9527), .S(n9528), .Z(n9655)
         );
  NAND2_X1 U12034 ( .A1(n9656), .A2(n9655), .ZN(n9654) );
  NAND2_X1 U12035 ( .A1(n9528), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9529) );
  NAND2_X1 U12036 ( .A1(n9654), .A2(n9529), .ZN(n9621) );
  INV_X1 U12037 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9530) );
  MUX2_X1 U12038 ( .A(n9530), .B(P2_REG1_REG_9__SCAN_IN), .S(n9629), .Z(n9531)
         );
  OR2_X1 U12039 ( .A1(n9621), .A2(n9531), .ZN(n9631) );
  OR2_X1 U12040 ( .A1(n9629), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n9532) );
  NAND2_X1 U12041 ( .A1(n9631), .A2(n9532), .ZN(n15226) );
  INV_X1 U12042 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n15397) );
  MUX2_X1 U12043 ( .A(n15397), .B(P2_REG1_REG_10__SCAN_IN), .S(n9533), .Z(
        n15227) );
  OR2_X1 U12044 ( .A1(n15226), .A2(n15227), .ZN(n15228) );
  NAND2_X1 U12045 ( .A1(n9533), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n9538) );
  NAND2_X1 U12046 ( .A1(n15228), .A2(n9538), .ZN(n9536) );
  INV_X1 U12047 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n9534) );
  MUX2_X1 U12048 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n9534), .S(n9714), .Z(n9535) );
  NAND2_X1 U12049 ( .A1(n9536), .A2(n9535), .ZN(n9706) );
  MUX2_X1 U12050 ( .A(n9534), .B(P2_REG1_REG_11__SCAN_IN), .S(n9714), .Z(n9537) );
  NAND3_X1 U12051 ( .A1(n15228), .A2(n9538), .A3(n9537), .ZN(n9539) );
  NAND3_X1 U12052 ( .A1(n9706), .A2(n15264), .A3(n9539), .ZN(n9540) );
  OAI211_X1 U12053 ( .C1(n9542), .C2(n15220), .A(n9541), .B(n9540), .ZN(
        P2_U3225) );
  INV_X1 U12054 ( .A(P3_DATAO_REG_5__SCAN_IN), .ZN(n13297) );
  NAND2_X1 U12055 ( .A1(n10468), .A2(P3_U3897), .ZN(n9543) );
  OAI21_X1 U12056 ( .B1(P3_U3897), .B2(n13297), .A(n9543), .ZN(P3_U3496) );
  INV_X1 U12057 ( .A(P3_DATAO_REG_2__SCAN_IN), .ZN(n13247) );
  NAND2_X1 U12058 ( .A1(n15462), .A2(P3_U3897), .ZN(n9544) );
  OAI21_X1 U12059 ( .B1(P3_U3897), .B2(n13247), .A(n9544), .ZN(P3_U3493) );
  INV_X1 U12060 ( .A(n9545), .ZN(n9546) );
  OAI222_X1 U12061 ( .A1(n14721), .A2(n9547), .B1(n14722), .B2(n9546), .C1(
        n11896), .C2(P3_U3151), .ZN(P3_U3280) );
  INV_X1 U12062 ( .A(n11377), .ZN(n9554) );
  OR2_X1 U12063 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n9548) );
  NAND2_X1 U12064 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n9548), .ZN(n9549) );
  NAND2_X1 U12065 ( .A1(n9550), .A2(n9549), .ZN(n9551) );
  XNOR2_X1 U12066 ( .A(n9551), .B(n7536), .ZN(n11378) );
  INV_X1 U12067 ( .A(n11378), .ZN(n15005) );
  OAI222_X1 U12068 ( .A1(n14694), .A2(n9552), .B1(n11910), .B2(n9554), .C1(
        P1_U3086), .C2(n15005), .ZN(P1_U3344) );
  OAI222_X1 U12069 ( .A1(n13852), .A2(n9555), .B1(n13854), .B2(n9554), .C1(
        P2_U3088), .C2(n9553), .ZN(P2_U3316) );
  INV_X1 U12070 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n11627) );
  NAND2_X1 U12071 ( .A1(n15271), .A2(n11627), .ZN(n9556) );
  OAI211_X1 U12072 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n15225), .A(n9556), .B(
        n15278), .ZN(n9557) );
  INV_X1 U12073 ( .A(n9557), .ZN(n9559) );
  AOI22_X1 U12074 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(n15264), .B1(n15271), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n9558) );
  MUX2_X1 U12075 ( .A(n9559), .B(n9558), .S(n7649), .Z(n9561) );
  AOI22_X1 U12076 ( .A1(n15270), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n9560) );
  NAND2_X1 U12077 ( .A1(n9561), .A2(n9560), .ZN(P2_U3214) );
  XNOR2_X1 U12078 ( .A(n6890), .B(n9643), .ZN(n9567) );
  INV_X1 U12079 ( .A(n9562), .ZN(n9565) );
  NAND2_X1 U12080 ( .A1(n9563), .A2(n6637), .ZN(n9564) );
  INV_X1 U12081 ( .A(n13492), .ZN(n13474) );
  AOI22_X1 U12082 ( .A1(n13474), .A2(n13532), .B1(n13475), .B2(n8463), .ZN(
        n9617) );
  INV_X1 U12083 ( .A(n9617), .ZN(n9566) );
  AOI21_X1 U12084 ( .B1(n9567), .B2(n14841), .A(n9566), .ZN(n10392) );
  NAND2_X1 U12085 ( .A1(n9614), .A2(n9645), .ZN(n9569) );
  AND3_X1 U12086 ( .A1(n9641), .A2(n14852), .A3(n9569), .ZN(n10386) );
  AOI21_X1 U12087 ( .B1(n15368), .B2(n9645), .A(n10386), .ZN(n9575) );
  XNOR2_X1 U12088 ( .A(n9571), .B(n9572), .ZN(n9573) );
  NAND2_X1 U12089 ( .A1(n9573), .A2(n13587), .ZN(n9611) );
  INV_X1 U12090 ( .A(n15342), .ZN(n11622) );
  XNOR2_X1 U12091 ( .A(n6636), .B(n6890), .ZN(n10390) );
  OAI21_X1 U12092 ( .B1(n9570), .B2(n11622), .A(n10390), .ZN(n9574) );
  AND3_X1 U12093 ( .A1(n10392), .A2(n9575), .A3(n9574), .ZN(n15313) );
  INV_X1 U12094 ( .A(n9576), .ZN(n9577) );
  AND2_X1 U12095 ( .A1(n9577), .A2(n15304), .ZN(n9578) );
  NAND2_X1 U12096 ( .A1(n9579), .A2(n9578), .ZN(n11021) );
  NAND2_X1 U12097 ( .A1(n15305), .A2(n9580), .ZN(n11020) );
  INV_X1 U12098 ( .A(n11019), .ZN(n9581) );
  NAND2_X1 U12099 ( .A1(n15399), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9582) );
  OAI21_X1 U12100 ( .B1(n15313), .B2(n15399), .A(n9582), .ZN(P2_U3500) );
  NAND3_X1 U12101 ( .A1(n11811), .A2(P1_B_REG_SCAN_IN), .A3(n11468), .ZN(n9583) );
  INV_X1 U12102 ( .A(n14696), .ZN(n9585) );
  NOR2_X1 U12103 ( .A1(n9585), .A2(P1_U3086), .ZN(n9586) );
  NAND2_X1 U12104 ( .A1(n9587), .A2(n9586), .ZN(n9590) );
  OAI22_X1 U12105 ( .A1(n15160), .A2(P1_D_REG_0__SCAN_IN), .B1(n9588), .B2(
        n9590), .ZN(n9589) );
  INV_X1 U12106 ( .A(n9589), .ZN(P1_U3445) );
  INV_X1 U12107 ( .A(n11468), .ZN(n9591) );
  OAI22_X1 U12108 ( .A1(n15160), .A2(P1_D_REG_1__SCAN_IN), .B1(n9591), .B2(
        n9590), .ZN(n9592) );
  INV_X1 U12109 ( .A(n9592), .ZN(P1_U3446) );
  INV_X1 U12110 ( .A(P3_DATAO_REG_18__SCAN_IN), .ZN(n13268) );
  NAND2_X1 U12111 ( .A1(n12834), .A2(P3_U3897), .ZN(n9593) );
  OAI21_X1 U12112 ( .B1(P3_U3897), .B2(n13268), .A(n9593), .ZN(P3_U3509) );
  MUX2_X1 U12113 ( .A(n10244), .B(P2_REG2_REG_6__SCAN_IN), .S(n9594), .Z(n9595) );
  NAND3_X1 U12114 ( .A1(n9597), .A2(n9596), .A3(n9595), .ZN(n9598) );
  NAND3_X1 U12115 ( .A1(n15271), .A2(n13557), .A3(n9598), .ZN(n9604) );
  NAND2_X1 U12116 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n10103) );
  OAI211_X1 U12117 ( .C1(n9600), .C2(n9599), .A(n15264), .B(n13551), .ZN(n9601) );
  NAND2_X1 U12118 ( .A1(n10103), .A2(n9601), .ZN(n9602) );
  AOI21_X1 U12119 ( .B1(n15270), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n9602), .ZN(
        n9603) );
  OAI211_X1 U12120 ( .C1(n15278), .C2(n9605), .A(n9604), .B(n9603), .ZN(
        P2_U3220) );
  OAI222_X1 U12121 ( .A1(n14721), .A2(n9607), .B1(n14722), .B2(n9606), .C1(
        n11899), .C2(P3_U3151), .ZN(P3_U3279) );
  INV_X1 U12122 ( .A(n11392), .ZN(n9639) );
  NAND2_X1 U12123 ( .A1(n9609), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9680) );
  XNOR2_X1 U12124 ( .A(n9680), .B(P1_IR_REG_13__SCAN_IN), .ZN(n15023) );
  INV_X1 U12125 ( .A(n15023), .ZN(n9610) );
  OAI222_X1 U12126 ( .A1(n11910), .A2(n9639), .B1(n14694), .B2(n8719), .C1(
        P1_U3086), .C2(n9610), .ZN(P1_U3342) );
  NAND2_X1 U12127 ( .A1(n9669), .A2(n13533), .ZN(n9612) );
  NAND2_X1 U12128 ( .A1(n9613), .A2(n9612), .ZN(n9666) );
  OAI21_X1 U12129 ( .B1(n9613), .B2(n9612), .A(n9666), .ZN(n9616) );
  AOI21_X1 U12130 ( .B1(n9616), .B2(n9615), .A(n9668), .ZN(n9620) );
  AOI21_X1 U12131 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n9676), .A(n9618), .ZN(
        n9619) );
  OAI21_X1 U12132 ( .B1(n9620), .B2(n13503), .A(n9619), .ZN(P2_U3194) );
  NOR2_X1 U12133 ( .A1(n15220), .A2(n9624), .ZN(n9623) );
  INV_X1 U12134 ( .A(n15278), .ZN(n15254) );
  INV_X1 U12135 ( .A(n9621), .ZN(n9630) );
  NOR3_X1 U12136 ( .A1(n15225), .A2(n9530), .A3(n9630), .ZN(n9622) );
  AOI211_X1 U12137 ( .C1(n9623), .C2(n9625), .A(n15254), .B(n9622), .ZN(n9637)
         );
  AND2_X1 U12138 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n10792) );
  NAND3_X1 U12139 ( .A1(n9625), .A2(n9636), .A3(n9624), .ZN(n9626) );
  AOI21_X1 U12140 ( .B1(n9627), .B2(n9626), .A(n15220), .ZN(n9628) );
  AOI211_X1 U12141 ( .C1(n15270), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n10792), .B(
        n9628), .ZN(n9635) );
  NOR3_X1 U12142 ( .A1(n9630), .A2(n9629), .A3(P2_REG1_REG_9__SCAN_IN), .ZN(
        n9633) );
  INV_X1 U12143 ( .A(n9631), .ZN(n9632) );
  OAI21_X1 U12144 ( .B1(n9633), .B2(n9632), .A(n15264), .ZN(n9634) );
  OAI211_X1 U12145 ( .C1(n9637), .C2(n9636), .A(n9635), .B(n9634), .ZN(
        P2_U3223) );
  INV_X1 U12146 ( .A(n10079), .ZN(n9710) );
  OAI222_X1 U12147 ( .A1(P2_U3088), .A2(n9710), .B1(n13854), .B2(n9639), .C1(
        n9638), .C2(n13852), .ZN(P2_U3314) );
  INV_X1 U12148 ( .A(n10198), .ZN(n10185) );
  XNOR2_X1 U12149 ( .A(n10186), .B(n10185), .ZN(n15287) );
  INV_X1 U12150 ( .A(n9570), .ZN(n15372) );
  INV_X1 U12151 ( .A(n9641), .ZN(n9642) );
  OR2_X1 U12152 ( .A1(n9641), .A2(n10200), .ZN(n10355) );
  OAI211_X1 U12153 ( .C1(n9642), .C2(n15281), .A(n14852), .B(n10355), .ZN(
        n15284) );
  OAI21_X1 U12154 ( .B1(n15281), .B2(n15380), .A(n15284), .ZN(n9652) );
  NAND2_X1 U12155 ( .A1(n9644), .A2(n9643), .ZN(n9648) );
  NAND2_X1 U12156 ( .A1(n9646), .A2(n9645), .ZN(n9647) );
  NAND2_X1 U12157 ( .A1(n9648), .A2(n9647), .ZN(n10199) );
  XNOR2_X1 U12158 ( .A(n10199), .B(n10198), .ZN(n9650) );
  AOI22_X1 U12159 ( .A1(n13474), .A2(n13531), .B1(n13475), .B2(n13533), .ZN(
        n9674) );
  INV_X1 U12160 ( .A(n9674), .ZN(n9649) );
  AOI21_X1 U12161 ( .B1(n14841), .B2(n9650), .A(n9649), .ZN(n15291) );
  INV_X1 U12162 ( .A(n15291), .ZN(n9651) );
  AOI211_X1 U12163 ( .C1(n15287), .C2(n15377), .A(n9652), .B(n9651), .ZN(
        n15315) );
  NAND2_X1 U12164 ( .A1(n15399), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9653) );
  OAI21_X1 U12165 ( .B1(n15315), .B2(n15399), .A(n9653), .ZN(P2_U3501) );
  OAI211_X1 U12166 ( .C1(n9656), .C2(n9655), .A(n15264), .B(n9654), .ZN(n9661)
         );
  OAI211_X1 U12167 ( .C1(n9659), .C2(n9658), .A(n15271), .B(n9657), .ZN(n9660)
         );
  NAND2_X1 U12168 ( .A1(n9661), .A2(n9660), .ZN(n9663) );
  NAND2_X1 U12169 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n10594) );
  INV_X1 U12170 ( .A(n10594), .ZN(n9662) );
  AOI211_X1 U12171 ( .C1(n15270), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n9663), .B(
        n9662), .ZN(n9664) );
  OAI21_X1 U12172 ( .B1(n9665), .B2(n15278), .A(n9664), .ZN(P2_U3222) );
  INV_X1 U12173 ( .A(n9666), .ZN(n9667) );
  XNOR2_X1 U12174 ( .A(n11968), .B(n15281), .ZN(n9671) );
  NAND2_X1 U12175 ( .A1(n9669), .A2(n13532), .ZN(n9670) );
  NAND2_X1 U12176 ( .A1(n9671), .A2(n9670), .ZN(n9691) );
  OAI21_X1 U12177 ( .B1(n9671), .B2(n9670), .A(n9691), .ZN(n9672) );
  AOI21_X1 U12178 ( .B1(n9673), .B2(n9672), .A(n9693), .ZN(n9678) );
  OAI22_X1 U12179 ( .A1(n13461), .A2(n15281), .B1(n9674), .B2(n13476), .ZN(
        n9675) );
  AOI21_X1 U12180 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n9676), .A(n9675), .ZN(
        n9677) );
  OAI21_X1 U12181 ( .B1(n9678), .B2(n13503), .A(n9677), .ZN(P2_U3209) );
  INV_X1 U12182 ( .A(n11367), .ZN(n9685) );
  NAND2_X1 U12183 ( .A1(n9680), .A2(n9679), .ZN(n9681) );
  NAND2_X1 U12184 ( .A1(n9681), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9682) );
  XNOR2_X1 U12185 ( .A(n9682), .B(P1_IR_REG_14__SCAN_IN), .ZN(n14338) );
  INV_X1 U12186 ( .A(n14338), .ZN(n15037) );
  OAI222_X1 U12187 ( .A1(n11910), .A2(n9685), .B1(n15037), .B2(P1_U3086), .C1(
        n9683), .C2(n14694), .ZN(P1_U3341) );
  INV_X1 U12188 ( .A(n10704), .ZN(n10693) );
  OAI222_X1 U12189 ( .A1(P2_U3088), .A2(n10693), .B1(n13854), .B2(n9685), .C1(
        n9684), .C2(n13852), .ZN(P2_U3313) );
  INV_X1 U12190 ( .A(n9686), .ZN(n9688) );
  OAI222_X1 U12191 ( .A1(n7335), .A2(P3_U3151), .B1(n14722), .B2(n9688), .C1(
        n9687), .C2(n14721), .ZN(P3_U3278) );
  OAI222_X1 U12192 ( .A1(P3_U3151), .A2(n12644), .B1(n14721), .B2(n9690), .C1(
        n14722), .C2(n9689), .ZN(P3_U3277) );
  INV_X1 U12193 ( .A(n9691), .ZN(n9692) );
  XNOR2_X1 U12194 ( .A(n11968), .B(n10359), .ZN(n9784) );
  NAND2_X1 U12195 ( .A1(n9669), .A2(n13531), .ZN(n9783) );
  XNOR2_X1 U12196 ( .A(n9784), .B(n9783), .ZN(n9786) );
  XNOR2_X1 U12197 ( .A(n9787), .B(n9786), .ZN(n9701) );
  INV_X1 U12198 ( .A(n13498), .ZN(n13467) );
  NAND2_X1 U12199 ( .A1(n13475), .A2(n13532), .ZN(n9696) );
  OR2_X1 U12200 ( .A1(n13492), .A2(n10208), .ZN(n9695) );
  AND2_X1 U12201 ( .A1(n9696), .A2(n9695), .ZN(n15317) );
  OAI21_X1 U12202 ( .B1(n13476), .B2(n15317), .A(n9697), .ZN(n9699) );
  NOR2_X1 U12203 ( .A1(n13461), .A2(n6842), .ZN(n9698) );
  AOI211_X1 U12204 ( .C1(n13467), .C2(n10352), .A(n9699), .B(n9698), .ZN(n9700) );
  OAI21_X1 U12205 ( .B1(n9701), .B2(n13503), .A(n9700), .ZN(P2_U3190) );
  INV_X1 U12206 ( .A(n15104), .ZN(n10044) );
  NOR2_X1 U12207 ( .A1(n10044), .A2(n14282), .ZN(P1_U3085) );
  INV_X1 U12208 ( .A(n11534), .ZN(n9704) );
  OR2_X1 U12209 ( .A1(n6768), .A2(n9233), .ZN(n9702) );
  XNOR2_X1 U12210 ( .A(n9702), .B(n9776), .ZN(n15052) );
  OAI222_X1 U12211 ( .A1(n11910), .A2(n9704), .B1(n15052), .B2(P1_U3086), .C1(
        n9703), .C2(n14694), .ZN(P1_U3340) );
  INV_X1 U12212 ( .A(n15253), .ZN(n10707) );
  OAI222_X1 U12213 ( .A1(P2_U3088), .A2(n10707), .B1(n13854), .B2(n9704), .C1(
        n13278), .C2(n13852), .ZN(P2_U3312) );
  NOR2_X1 U12214 ( .A1(n10079), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n9707) );
  NAND2_X1 U12215 ( .A1(n9714), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n9705) );
  AND2_X1 U12216 ( .A1(n9706), .A2(n9705), .ZN(n15242) );
  INV_X1 U12217 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n13312) );
  MUX2_X1 U12218 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n13312), .S(n9717), .Z(
        n15241) );
  NAND2_X1 U12219 ( .A1(n15242), .A2(n15241), .ZN(n15240) );
  OAI21_X1 U12220 ( .B1(n9717), .B2(P2_REG1_REG_12__SCAN_IN), .A(n15240), .ZN(
        n9709) );
  AOI211_X1 U12221 ( .C1(P2_REG1_REG_13__SCAN_IN), .C2(n10079), .A(n9707), .B(
        n9709), .ZN(n10078) );
  NAND2_X1 U12222 ( .A1(n9710), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n9708) );
  OAI211_X1 U12223 ( .C1(P2_REG1_REG_13__SCAN_IN), .C2(n9710), .A(n9709), .B(
        n9708), .ZN(n9711) );
  NAND2_X1 U12224 ( .A1(n9711), .A2(n15264), .ZN(n9724) );
  OAI22_X1 U12225 ( .A1(n15250), .A2(n14990), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9712), .ZN(n9722) );
  INV_X1 U12226 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n9713) );
  MUX2_X1 U12227 ( .A(n9713), .B(P2_REG2_REG_13__SCAN_IN), .S(n10079), .Z(
        n9720) );
  OR2_X1 U12228 ( .A1(n9714), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n15234) );
  NAND2_X1 U12229 ( .A1(n15236), .A2(n15234), .ZN(n9716) );
  INV_X1 U12230 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n9715) );
  MUX2_X1 U12231 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n9715), .S(n9717), .Z(
        n15233) );
  NAND2_X1 U12232 ( .A1(n9716), .A2(n15233), .ZN(n15238) );
  OAI21_X1 U12233 ( .B1(n9717), .B2(P2_REG2_REG_12__SCAN_IN), .A(n15238), .ZN(
        n9719) );
  NOR2_X1 U12234 ( .A1(n10079), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n9718) );
  AOI211_X1 U12235 ( .C1(P2_REG2_REG_13__SCAN_IN), .C2(n10079), .A(n9718), .B(
        n9719), .ZN(n10076) );
  AOI211_X1 U12236 ( .C1(n9720), .C2(n9719), .A(n15220), .B(n10076), .ZN(n9721) );
  AOI211_X1 U12237 ( .C1(n15254), .C2(n10079), .A(n9722), .B(n9721), .ZN(n9723) );
  OAI21_X1 U12238 ( .B1(n10078), .B2(n9724), .A(n9723), .ZN(P2_U3227) );
  INV_X1 U12239 ( .A(n10555), .ZN(n9883) );
  INV_X1 U12240 ( .A(n10324), .ZN(n9748) );
  INV_X1 U12241 ( .A(n9963), .ZN(n9735) );
  INV_X1 U12242 ( .A(n9725), .ZN(n9726) );
  INV_X1 U12243 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9727) );
  MUX2_X1 U12244 ( .A(n9727), .B(P1_REG1_REG_5__SCAN_IN), .S(n10324), .Z(n9746) );
  NAND2_X1 U12245 ( .A1(n9747), .A2(n9746), .ZN(n9745) );
  XOR2_X1 U12246 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10555), .Z(n9879) );
  NOR2_X1 U12247 ( .A1(n9878), .A2(n9879), .ZN(n9877) );
  INV_X1 U12248 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9728) );
  MUX2_X1 U12249 ( .A(n9728), .B(P1_REG1_REG_7__SCAN_IN), .S(n10800), .Z(n9891) );
  NOR2_X1 U12250 ( .A1(n9892), .A2(n9891), .ZN(n9890) );
  AOI21_X1 U12251 ( .B1(n10800), .B2(P1_REG1_REG_7__SCAN_IN), .A(n9890), .ZN(
        n9731) );
  INV_X1 U12252 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9729) );
  MUX2_X1 U12253 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n9729), .S(n10853), .Z(n9730) );
  NAND2_X1 U12254 ( .A1(n9731), .A2(n9730), .ZN(n9760) );
  OAI21_X1 U12255 ( .B1(n9731), .B2(n9730), .A(n9760), .ZN(n9743) );
  INV_X1 U12256 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9733) );
  NAND2_X1 U12257 ( .A1(n15068), .A2(n10853), .ZN(n9732) );
  NAND2_X1 U12258 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n11208) );
  OAI211_X1 U12259 ( .C1(n15104), .C2(n9733), .A(n9732), .B(n11208), .ZN(n9742) );
  INV_X1 U12260 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9736) );
  MUX2_X1 U12261 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n9736), .S(n10324), .Z(n9753) );
  INV_X1 U12262 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10574) );
  XNOR2_X1 U12263 ( .A(n10555), .B(n10574), .ZN(n9881) );
  NOR2_X1 U12264 ( .A1(n9882), .A2(n9881), .ZN(n9880) );
  AOI21_X1 U12265 ( .B1(n9883), .B2(P1_REG2_REG_6__SCAN_IN), .A(n9880), .ZN(
        n9895) );
  INV_X1 U12266 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9737) );
  MUX2_X1 U12267 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n9737), .S(n10800), .Z(n9738) );
  INV_X1 U12268 ( .A(n9738), .ZN(n9894) );
  NOR2_X1 U12269 ( .A1(n9895), .A2(n9894), .ZN(n9893) );
  XNOR2_X1 U12270 ( .A(n10853), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n9739) );
  AOI211_X1 U12271 ( .C1(n9740), .C2(n9739), .A(n15061), .B(n9765), .ZN(n9741)
         );
  AOI211_X1 U12272 ( .C1(n15091), .C2(n9743), .A(n9742), .B(n9741), .ZN(n9744)
         );
  INV_X1 U12273 ( .A(n9744), .ZN(P1_U3251) );
  OAI21_X1 U12274 ( .B1(n9747), .B2(n9746), .A(n9745), .ZN(n9757) );
  NAND2_X1 U12275 ( .A1(n15068), .A2(n9748), .ZN(n9750) );
  NAND2_X1 U12276 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9749) );
  OAI211_X1 U12277 ( .C1(n9751), .C2(n15104), .A(n9750), .B(n9749), .ZN(n9756)
         );
  AOI211_X1 U12278 ( .C1(n9754), .C2(n9753), .A(n9752), .B(n15061), .ZN(n9755)
         );
  AOI211_X1 U12279 ( .C1(n15091), .C2(n9757), .A(n9756), .B(n9755), .ZN(n9758)
         );
  INV_X1 U12280 ( .A(n9758), .ZN(P1_U3248) );
  INV_X1 U12281 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9759) );
  MUX2_X1 U12282 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n9759), .S(n11080), .Z(n9762) );
  OAI21_X1 U12283 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n10853), .A(n9760), .ZN(
        n9761) );
  NAND2_X1 U12284 ( .A1(n9761), .A2(n9762), .ZN(n9907) );
  OAI21_X1 U12285 ( .B1(n9762), .B2(n9761), .A(n9907), .ZN(n9772) );
  NAND2_X1 U12286 ( .A1(n15068), .A2(n11080), .ZN(n9763) );
  NAND2_X1 U12287 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n11361) );
  OAI211_X1 U12288 ( .C1(n9764), .C2(n15104), .A(n9763), .B(n11361), .ZN(n9771) );
  INV_X1 U12289 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9766) );
  MUX2_X1 U12290 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n9766), .S(n11080), .Z(n9767) );
  INV_X1 U12291 ( .A(n9767), .ZN(n9768) );
  AOI211_X1 U12292 ( .C1(n9769), .C2(n9768), .A(n15061), .B(n9901), .ZN(n9770)
         );
  AOI211_X1 U12293 ( .C1(n15091), .C2(n9772), .A(n9771), .B(n9770), .ZN(n9773)
         );
  INV_X1 U12294 ( .A(n9773), .ZN(P1_U3252) );
  OAI222_X1 U12295 ( .A1(n14722), .A2(n9775), .B1(n14721), .B2(n9774), .C1(
        P3_U3151), .C2(n12039), .ZN(P3_U3276) );
  INV_X1 U12296 ( .A(n11670), .ZN(n9782) );
  AND2_X1 U12297 ( .A1(n6768), .A2(n9776), .ZN(n9777) );
  OR2_X1 U12298 ( .A1(n9777), .A2(n9233), .ZN(n9778) );
  XNOR2_X1 U12299 ( .A(n9778), .B(P1_IR_REG_16__SCAN_IN), .ZN(n15067) );
  INV_X1 U12300 ( .A(n15067), .ZN(n9780) );
  OAI222_X1 U12301 ( .A1(n11910), .A2(n9782), .B1(n9780), .B2(P1_U3086), .C1(
        n9779), .C2(n14694), .ZN(P1_U3339) );
  INV_X1 U12302 ( .A(n10702), .ZN(n11182) );
  OAI222_X1 U12303 ( .A1(P2_U3088), .A2(n11182), .B1(n13854), .B2(n9782), .C1(
        n9781), .C2(n13852), .ZN(P2_U3311) );
  INV_X1 U12304 ( .A(n9783), .ZN(n9785) );
  BUF_X2 U12305 ( .A(n9669), .Z(n11957) );
  AND2_X1 U12306 ( .A1(n11957), .A2(n13530), .ZN(n9789) );
  XNOR2_X1 U12307 ( .A(n11968), .B(n15324), .ZN(n9788) );
  NOR2_X1 U12308 ( .A1(n9788), .A2(n9789), .ZN(n9919) );
  AOI21_X1 U12309 ( .B1(n9789), .B2(n9788), .A(n9919), .ZN(n9790) );
  OAI21_X1 U12310 ( .B1(n9791), .B2(n9790), .A(n9921), .ZN(n9798) );
  NOR2_X1 U12311 ( .A1(n13498), .A2(n10228), .ZN(n9797) );
  NAND2_X1 U12312 ( .A1(n13475), .A2(n13531), .ZN(n9793) );
  OR2_X1 U12313 ( .A1(n13492), .A2(n10238), .ZN(n9792) );
  AND2_X1 U12314 ( .A1(n9793), .A2(n9792), .ZN(n10220) );
  NAND2_X1 U12315 ( .A1(n13501), .A2(n15324), .ZN(n9795) );
  OAI211_X1 U12316 ( .C1(n10220), .C2(n13476), .A(n9795), .B(n9794), .ZN(n9796) );
  AOI211_X1 U12317 ( .C1(n9798), .C2(n13454), .A(n9797), .B(n9796), .ZN(n9799)
         );
  INV_X1 U12318 ( .A(n9799), .ZN(P2_U3202) );
  NOR4_X1 U12319 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n9806) );
  NOR4_X1 U12320 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n9805) );
  NOR4_X1 U12321 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9804) );
  NOR4_X1 U12322 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n9803) );
  NAND4_X1 U12323 ( .A1(n9806), .A2(n9805), .A3(n9804), .A4(n9803), .ZN(n9812)
         );
  NOR2_X1 U12324 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .ZN(
        n9810) );
  NOR4_X1 U12325 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n9809) );
  NOR4_X1 U12326 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n9808) );
  NOR4_X1 U12327 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n9807) );
  NAND4_X1 U12328 ( .A1(n9810), .A2(n9809), .A3(n9808), .A4(n9807), .ZN(n9811)
         );
  NOR2_X1 U12329 ( .A1(n9812), .A2(n9811), .ZN(n9813) );
  NOR2_X1 U12330 ( .A1(n9816), .A2(n9813), .ZN(n9852) );
  INV_X1 U12331 ( .A(n9852), .ZN(n9819) );
  NAND2_X1 U12332 ( .A1(n11811), .A2(n14696), .ZN(n9814) );
  NAND2_X1 U12333 ( .A1(n9815), .A2(n9814), .ZN(n10558) );
  INV_X1 U12334 ( .A(n10558), .ZN(n10033) );
  OR2_X1 U12335 ( .A1(n9816), .A2(P1_D_REG_1__SCAN_IN), .ZN(n9818) );
  NAND2_X1 U12336 ( .A1(n11468), .A2(n14696), .ZN(n9817) );
  NAND2_X1 U12337 ( .A1(n9818), .A2(n9817), .ZN(n9930) );
  INV_X1 U12338 ( .A(n9930), .ZN(n10559) );
  NAND3_X1 U12339 ( .A1(n9819), .A2(n10033), .A3(n10559), .ZN(n9844) );
  NOR2_X1 U12340 ( .A1(n9844), .A2(n9820), .ZN(n9842) );
  AND2_X1 U12341 ( .A1(n14195), .A2(n14010), .ZN(n14249) );
  NAND2_X1 U12342 ( .A1(n14007), .A2(n14249), .ZN(n10573) );
  INV_X1 U12343 ( .A(n10573), .ZN(n9825) );
  MUX2_X1 U12344 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9822), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n9823) );
  INV_X1 U12345 ( .A(n9929), .ZN(n9824) );
  NAND2_X1 U12346 ( .A1(n11715), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n9828) );
  NAND2_X1 U12347 ( .A1(n9954), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9827) );
  NAND2_X1 U12348 ( .A1(n9942), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n9826) );
  NAND2_X1 U12349 ( .A1(n11093), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9829) );
  XNOR2_X1 U12350 ( .A(n9832), .B(n10525), .ZN(n9834) );
  NOR2_X1 U12351 ( .A1(n9834), .A2(n9833), .ZN(n10066) );
  OAI21_X1 U12352 ( .B1(n12242), .B2(n9836), .A(n9835), .ZN(n9837) );
  OAI21_X1 U12353 ( .B1(n9838), .B2(n9837), .A(n10068), .ZN(n9843) );
  INV_X1 U12354 ( .A(n10059), .ZN(n9839) );
  NAND2_X1 U12355 ( .A1(n9839), .A2(n14579), .ZN(n9840) );
  AND2_X1 U12356 ( .A1(n15187), .A2(n14022), .ZN(n9841) );
  NAND2_X1 U12357 ( .A1(n9843), .A2(n13994), .ZN(n9857) );
  NAND2_X1 U12358 ( .A1(n9844), .A2(n9929), .ZN(n10531) );
  INV_X1 U12359 ( .A(n14010), .ZN(n14020) );
  NAND2_X1 U12360 ( .A1(n14020), .A2(n14352), .ZN(n9845) );
  NAND2_X1 U12361 ( .A1(n9854), .A2(n9845), .ZN(n10530) );
  NAND2_X1 U12362 ( .A1(n9846), .A2(n10530), .ZN(n14255) );
  INV_X1 U12363 ( .A(n14255), .ZN(n9847) );
  NAND2_X1 U12364 ( .A1(n10531), .A2(n9847), .ZN(n10073) );
  NAND2_X1 U12365 ( .A1(n11775), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n9851) );
  NAND2_X1 U12366 ( .A1(n11093), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9850) );
  NAND2_X1 U12367 ( .A1(n9954), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9849) );
  NAND2_X1 U12368 ( .A1(n9942), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9848) );
  INV_X1 U12369 ( .A(n14280), .ZN(n10062) );
  NAND2_X1 U12370 ( .A1(n9931), .A2(n10559), .ZN(n13918) );
  NAND2_X1 U12371 ( .A1(n9854), .A2(n9266), .ZN(n14533) );
  OR2_X1 U12372 ( .A1(n13918), .A2(n14533), .ZN(n14926) );
  NAND2_X1 U12373 ( .A1(n9854), .A2(n9853), .ZN(n14531) );
  OR2_X1 U12374 ( .A1(n13918), .A2(n14531), .ZN(n14925) );
  OAI22_X1 U12375 ( .A1(n10062), .A2(n14926), .B1(n14925), .B2(n10626), .ZN(
        n9855) );
  AOI21_X1 U12376 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n10073), .A(n9855), .ZN(
        n9856) );
  OAI211_X1 U12377 ( .C1(n9972), .C2(n14005), .A(n9857), .B(n9856), .ZN(
        P1_U3222) );
  INV_X1 U12378 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10146) );
  NAND2_X1 U12379 ( .A1(n13016), .A2(n9858), .ZN(n9859) );
  OAI21_X1 U12380 ( .B1(n13016), .B2(n9860), .A(n9859), .ZN(n9861) );
  INV_X1 U12381 ( .A(n9861), .ZN(n9862) );
  INV_X1 U12382 ( .A(n15444), .ZN(n15471) );
  NOR2_X1 U12383 ( .A1(n15521), .A2(n15471), .ZN(n9864) );
  AND2_X1 U12384 ( .A1(n12201), .A2(n15463), .ZN(n12017) );
  NOR2_X1 U12385 ( .A1(n15460), .A2(n12017), .ZN(n10117) );
  OR3_X1 U12386 ( .A1(n10117), .A2(n15488), .A3(n9865), .ZN(n9866) );
  OAI21_X1 U12387 ( .B1(n15451), .B2(n15448), .A(n9866), .ZN(n12199) );
  AOI22_X1 U12388 ( .A1(n12199), .A2(n15477), .B1(P3_REG3_REG_0__SCAN_IN), 
        .B2(n15473), .ZN(n9869) );
  OR2_X1 U12389 ( .A1(n9867), .A2(n15444), .ZN(n12794) );
  NAND2_X1 U12390 ( .A1(n12885), .A2(n10114), .ZN(n9868) );
  OAI211_X1 U12391 ( .C1(n10146), .C2(n15477), .A(n9869), .B(n9868), .ZN(
        P3_U3233) );
  INV_X1 U12392 ( .A(n14926), .ZN(n13997) );
  AOI22_X1 U12393 ( .A1(n13997), .A2(n6932), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n10073), .ZN(n9871) );
  NAND2_X1 U12394 ( .A1(n14937), .A2(n10667), .ZN(n9870) );
  OAI211_X1 U12395 ( .C1(n9872), .C2(n14932), .A(n9871), .B(n9870), .ZN(
        P1_U3232) );
  INV_X1 U12396 ( .A(n11675), .ZN(n9916) );
  NAND2_X1 U12397 ( .A1(n9873), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9874) );
  MUX2_X1 U12398 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9874), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n9875) );
  AND2_X1 U12399 ( .A1(n9875), .A2(n10118), .ZN(n14343) );
  INV_X1 U12400 ( .A(n14343), .ZN(n15082) );
  OAI222_X1 U12401 ( .A1(n11910), .A2(n9916), .B1(n15082), .B2(P1_U3086), .C1(
        n9876), .C2(n14694), .ZN(P1_U3338) );
  INV_X1 U12402 ( .A(n15091), .ZN(n15057) );
  AOI211_X1 U12403 ( .C1(n9879), .C2(n9878), .A(n9877), .B(n15057), .ZN(n9889)
         );
  AOI211_X1 U12404 ( .C1(n9882), .C2(n9881), .A(n9880), .B(n15061), .ZN(n9888)
         );
  NAND2_X1 U12405 ( .A1(n15068), .A2(n9883), .ZN(n9885) );
  NAND2_X1 U12406 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n9884) );
  OAI211_X1 U12407 ( .C1(n9886), .C2(n15104), .A(n9885), .B(n9884), .ZN(n9887)
         );
  OR3_X1 U12408 ( .A1(n9889), .A2(n9888), .A3(n9887), .ZN(P1_U3249) );
  AOI211_X1 U12409 ( .C1(n9892), .C2(n9891), .A(n9890), .B(n15057), .ZN(n9900)
         );
  AOI211_X1 U12410 ( .C1(n9895), .C2(n9894), .A(n15061), .B(n9893), .ZN(n9899)
         );
  NAND2_X1 U12411 ( .A1(n15068), .A2(n10800), .ZN(n9896) );
  NAND2_X1 U12412 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n11053) );
  OAI211_X1 U12413 ( .C1(n9897), .C2(n15104), .A(n9896), .B(n11053), .ZN(n9898) );
  OR3_X1 U12414 ( .A1(n9900), .A2(n9899), .A3(n9898), .ZN(P1_U3250) );
  AOI21_X1 U12415 ( .B1(n11080), .B2(P1_REG2_REG_9__SCAN_IN), .A(n9901), .ZN(
        n9905) );
  INV_X1 U12416 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n9902) );
  MUX2_X1 U12417 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n9902), .S(n11072), .Z(
        n9903) );
  INV_X1 U12418 ( .A(n9903), .ZN(n9904) );
  NOR2_X1 U12419 ( .A1(n9905), .A2(n9904), .ZN(n10040) );
  AOI211_X1 U12420 ( .C1(n9905), .C2(n9904), .A(n15061), .B(n10040), .ZN(n9914) );
  INV_X1 U12421 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9906) );
  MUX2_X1 U12422 ( .A(n9906), .B(P1_REG1_REG_10__SCAN_IN), .S(n11072), .Z(
        n9909) );
  OAI21_X1 U12423 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n11080), .A(n9907), .ZN(
        n9908) );
  NOR2_X1 U12424 ( .A1(n9908), .A2(n9909), .ZN(n10049) );
  AOI211_X1 U12425 ( .C1(n9909), .C2(n9908), .A(n15057), .B(n10049), .ZN(n9913) );
  NAND2_X1 U12426 ( .A1(n15068), .A2(n11072), .ZN(n9910) );
  NAND2_X1 U12427 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n11507)
         );
  OAI211_X1 U12428 ( .C1(n9911), .C2(n15104), .A(n9910), .B(n11507), .ZN(n9912) );
  OR3_X1 U12429 ( .A1(n9914), .A2(n9913), .A3(n9912), .ZN(P1_U3253) );
  INV_X1 U12430 ( .A(n11180), .ZN(n15277) );
  OAI222_X1 U12431 ( .A1(P2_U3088), .A2(n15277), .B1(n13854), .B2(n9916), .C1(
        n9915), .C2(n13852), .ZN(P2_U3310) );
  INV_X1 U12432 ( .A(n10239), .ZN(n15333) );
  AND2_X1 U12433 ( .A1(n11957), .A2(n13529), .ZN(n9918) );
  XNOR2_X1 U12434 ( .A(n11968), .B(n10239), .ZN(n9917) );
  NOR2_X1 U12435 ( .A1(n9917), .A2(n9918), .ZN(n10098) );
  AOI21_X1 U12436 ( .B1(n9918), .B2(n9917), .A(n10098), .ZN(n9923) );
  INV_X1 U12437 ( .A(n9919), .ZN(n9920) );
  OAI21_X1 U12438 ( .B1(n9923), .B2(n9922), .A(n10100), .ZN(n9924) );
  NAND2_X1 U12439 ( .A1(n9924), .A2(n13454), .ZN(n9928) );
  AOI22_X1 U12440 ( .A1(n13474), .A2(n13528), .B1(n13475), .B2(n13530), .ZN(
        n10211) );
  OAI21_X1 U12441 ( .B1(n13476), .B2(n10211), .A(n9925), .ZN(n9926) );
  AOI21_X1 U12442 ( .B1(n10195), .B2(n13467), .A(n9926), .ZN(n9927) );
  OAI211_X1 U12443 ( .C1(n15333), .C2(n13461), .A(n9928), .B(n9927), .ZN(
        P2_U3199) );
  INV_X1 U12444 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9982) );
  INV_X1 U12445 ( .A(n14008), .ZN(n9932) );
  NAND2_X1 U12446 ( .A1(n9932), .A2(n14038), .ZN(n9933) );
  NAND2_X1 U12447 ( .A1(n10633), .A2(n14352), .ZN(n11129) );
  NOR2_X1 U12448 ( .A1(n14010), .A2(n14352), .ZN(n9934) );
  NAND2_X1 U12449 ( .A1(n14007), .A2(n9934), .ZN(n15175) );
  NAND2_X1 U12450 ( .A1(n9935), .A2(n10667), .ZN(n10635) );
  NAND2_X1 U12451 ( .A1(n14222), .A2(n10635), .ZN(n9937) );
  NAND2_X1 U12452 ( .A1(n10072), .A2(n9972), .ZN(n9936) );
  NAND2_X1 U12453 ( .A1(n9937), .A2(n9936), .ZN(n15106) );
  OR2_X1 U12454 ( .A1(n6649), .A2(n11620), .ZN(n9939) );
  NAND2_X1 U12455 ( .A1(n10062), .A2(n6840), .ZN(n9940) );
  NAND2_X1 U12456 ( .A1(n9941), .A2(n9940), .ZN(n10652) );
  INV_X1 U12457 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9943) );
  NAND2_X1 U12458 ( .A1(n11751), .A2(n9943), .ZN(n9947) );
  NAND2_X1 U12459 ( .A1(n9954), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9946) );
  NAND2_X1 U12460 ( .A1(n11093), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9944) );
  INV_X1 U12461 ( .A(n10515), .ZN(n14279) );
  OR2_X1 U12462 ( .A1(n6648), .A2(n7036), .ZN(n9949) );
  NAND2_X1 U12463 ( .A1(n14279), .A2(n15179), .ZN(n14050) );
  NAND2_X1 U12464 ( .A1(n10515), .A2(n9950), .ZN(n14049) );
  NAND2_X1 U12465 ( .A1(n10515), .A2(n15179), .ZN(n9951) );
  INV_X1 U12466 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n9953) );
  XNOR2_X1 U12467 ( .A(n9953), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n10716) );
  NAND2_X1 U12468 ( .A1(n11751), .A2(n10716), .ZN(n9958) );
  NAND2_X1 U12469 ( .A1(n11774), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9957) );
  NAND2_X1 U12470 ( .A1(n11093), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9956) );
  BUF_X2 U12471 ( .A(n11715), .Z(n14012) );
  NAND2_X1 U12472 ( .A1(n14012), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9955) );
  NAND4_X1 U12473 ( .A1(n9958), .A2(n9957), .A3(n9956), .A4(n9955), .ZN(n14278) );
  OR2_X1 U12474 ( .A1(n14025), .A2(n9959), .ZN(n9962) );
  OR2_X1 U12475 ( .A1(n6649), .A2(n9960), .ZN(n9961) );
  XNOR2_X1 U12476 ( .A(n14278), .B(n14053), .ZN(n14220) );
  XNOR2_X1 U12477 ( .A(n10320), .B(n14220), .ZN(n10724) );
  OR2_X1 U12478 ( .A1(n10515), .A2(n14531), .ZN(n9970) );
  AOI21_X1 U12479 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9964) );
  NOR2_X1 U12480 ( .A1(n9964), .A2(n10331), .ZN(n11069) );
  NAND2_X1 U12481 ( .A1(n11751), .A2(n11069), .ZN(n9968) );
  NAND2_X1 U12482 ( .A1(n11774), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9967) );
  NAND2_X1 U12483 ( .A1(n11775), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9966) );
  NAND2_X1 U12484 ( .A1(n14011), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9965) );
  NAND4_X1 U12485 ( .A1(n9968), .A2(n9967), .A3(n9966), .A4(n9965), .ZN(n14277) );
  NAND2_X1 U12486 ( .A1(n14277), .A2(n14573), .ZN(n9969) );
  NAND2_X1 U12487 ( .A1(n9970), .A2(n9969), .ZN(n10717) );
  OR2_X1 U12488 ( .A1(n10632), .A2(n10667), .ZN(n15119) );
  INV_X1 U12489 ( .A(n10340), .ZN(n9971) );
  AOI211_X1 U12490 ( .C1(n14053), .C2(n10649), .A(n15161), .B(n9971), .ZN(
        n10715) );
  AOI211_X1 U12491 ( .C1(n14053), .C2(n14955), .A(n10717), .B(n10715), .ZN(
        n9980) );
  NAND2_X1 U12492 ( .A1(n10626), .A2(n10667), .ZN(n14033) );
  NAND2_X1 U12493 ( .A1(n6932), .A2(n9972), .ZN(n14034) );
  INV_X1 U12494 ( .A(n14034), .ZN(n9973) );
  NAND2_X1 U12495 ( .A1(n10072), .A2(n10632), .ZN(n14041) );
  OAI21_X1 U12496 ( .B1(n14033), .B2(n9973), .A(n14041), .ZN(n15107) );
  NAND2_X1 U12497 ( .A1(n15107), .A2(n14043), .ZN(n9975) );
  NAND2_X1 U12498 ( .A1(n10062), .A2(n15118), .ZN(n9974) );
  NAND2_X1 U12499 ( .A1(n9975), .A2(n9974), .ZN(n10646) );
  NAND2_X1 U12500 ( .A1(n10646), .A2(n14221), .ZN(n9976) );
  NAND2_X1 U12501 ( .A1(n9976), .A2(n14049), .ZN(n10327) );
  XNOR2_X1 U12502 ( .A(n10327), .B(n14220), .ZN(n10722) );
  NAND2_X1 U12503 ( .A1(n9977), .A2(n14010), .ZN(n9978) );
  OAI21_X2 U12504 ( .B1(n14007), .B2(n14352), .A(n9978), .ZN(n14971) );
  NAND2_X1 U12505 ( .A1(n10722), .A2(n14971), .ZN(n9979) );
  OAI211_X1 U12506 ( .C1(n14670), .C2(n10724), .A(n9980), .B(n9979), .ZN(
        n10036) );
  NAND2_X1 U12507 ( .A1(n10036), .A2(n15202), .ZN(n9981) );
  OAI21_X1 U12508 ( .B1(n15202), .B2(n9982), .A(n9981), .ZN(P1_U3532) );
  INV_X1 U12509 ( .A(n10006), .ZN(n9988) );
  AND3_X1 U12510 ( .A1(n9984), .A2(n10125), .A3(n9983), .ZN(n9987) );
  INV_X1 U12511 ( .A(n10007), .ZN(n9985) );
  OR2_X1 U12512 ( .A1(n10013), .A2(n9985), .ZN(n9986) );
  OAI211_X1 U12513 ( .C1(n10015), .C2(n9988), .A(n9987), .B(n9986), .ZN(n9989)
         );
  NAND2_X1 U12514 ( .A1(n9989), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9991) );
  OR2_X1 U12515 ( .A1(n10013), .A2(n12188), .ZN(n9990) );
  NOR2_X1 U12516 ( .A1(n12530), .A2(P3_U3151), .ZN(n10112) );
  INV_X1 U12517 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n10022) );
  INV_X1 U12518 ( .A(n9992), .ZN(n12184) );
  NAND2_X1 U12519 ( .A1(n12049), .A2(n12014), .ZN(n9993) );
  NAND2_X1 U12520 ( .A1(n9993), .A2(n10109), .ZN(n9994) );
  XNOR2_X1 U12521 ( .A(n9995), .B(n10089), .ZN(n10088) );
  XNOR2_X1 U12522 ( .A(n10088), .B(n15462), .ZN(n10005) );
  NAND2_X1 U12523 ( .A1(n9996), .A2(n15451), .ZN(n10003) );
  NAND3_X1 U12524 ( .A1(n9997), .A2(n12379), .A3(n9998), .ZN(n9999) );
  NAND2_X1 U12525 ( .A1(n12379), .A2(n15465), .ZN(n10000) );
  NAND2_X1 U12526 ( .A1(n10001), .A2(n10000), .ZN(n10002) );
  NAND2_X1 U12527 ( .A1(n10028), .A2(n10002), .ZN(n10027) );
  NAND2_X1 U12528 ( .A1(n10027), .A2(n10003), .ZN(n10004) );
  OAI21_X1 U12529 ( .B1(n10005), .B2(n10004), .A(n10092), .ZN(n10011) );
  NAND3_X1 U12530 ( .A1(n10015), .A2(n10006), .A3(n15521), .ZN(n10009) );
  NAND2_X1 U12531 ( .A1(n10013), .A2(n10007), .ZN(n10008) );
  NAND2_X1 U12532 ( .A1(n10009), .A2(n10008), .ZN(n10010) );
  NAND2_X1 U12533 ( .A1(n10011), .A2(n12522), .ZN(n10021) );
  INV_X1 U12534 ( .A(n12188), .ZN(n10012) );
  NAND2_X1 U12535 ( .A1(n10013), .A2(n10012), .ZN(n10018) );
  OR2_X2 U12536 ( .A1(n10018), .A2(n10014), .ZN(n12527) );
  INV_X1 U12537 ( .A(n12527), .ZN(n10024) );
  NAND3_X1 U12538 ( .A1(n10015), .A2(n15488), .A3(n10124), .ZN(n10016) );
  INV_X1 U12539 ( .A(n12517), .ZN(n12533) );
  OR2_X2 U12540 ( .A1(n10018), .A2(n10017), .ZN(n12526) );
  OAI22_X1 U12541 ( .A1(n12533), .A2(n15442), .B1(n15449), .B2(n12526), .ZN(
        n10019) );
  AOI21_X1 U12542 ( .B1(n10024), .B2(n9997), .A(n10019), .ZN(n10020) );
  OAI211_X1 U12543 ( .C1(n10112), .C2(n10022), .A(n10021), .B(n10020), .ZN(
        P3_U3177) );
  INV_X1 U12544 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10032) );
  OAI22_X1 U12545 ( .A1(n12533), .A2(n7796), .B1(n10482), .B2(n12526), .ZN(
        n10023) );
  AOI21_X1 U12546 ( .B1(n10024), .B2(n15463), .A(n10023), .ZN(n10031) );
  INV_X1 U12547 ( .A(n15460), .ZN(n12023) );
  NAND3_X1 U12548 ( .A1(n12023), .A2(n10025), .A3(n12390), .ZN(n10026) );
  OAI211_X1 U12549 ( .C1(n10028), .C2(n15465), .A(n10027), .B(n10026), .ZN(
        n10029) );
  NAND2_X1 U12550 ( .A1(n10029), .A2(n12522), .ZN(n10030) );
  OAI211_X1 U12551 ( .C1(n10112), .C2(n10032), .A(n10031), .B(n10030), .ZN(
        P3_U3162) );
  NOR2_X1 U12552 ( .A1(n10557), .A2(n10033), .ZN(n10035) );
  INV_X1 U12553 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10038) );
  NAND2_X1 U12554 ( .A1(n10036), .A2(n15194), .ZN(n10037) );
  OAI21_X1 U12555 ( .B1(n15194), .B2(n10038), .A(n10037), .ZN(P1_U3471) );
  INV_X1 U12556 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10039) );
  AOI22_X1 U12557 ( .A1(n14337), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n10039), 
        .B2(n10048), .ZN(n10043) );
  NAND2_X1 U12558 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n11378), .ZN(n10041) );
  OAI21_X1 U12559 ( .B1(n11378), .B2(P1_REG2_REG_11__SCAN_IN), .A(n10041), 
        .ZN(n15007) );
  OAI21_X1 U12560 ( .B1(n10043), .B2(n10042), .A(n14326), .ZN(n10047) );
  NAND2_X1 U12561 ( .A1(n10044), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n10045) );
  NAND2_X1 U12562 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n13902)
         );
  OAI211_X1 U12563 ( .C1(n15100), .C2(n10048), .A(n10045), .B(n13902), .ZN(
        n10046) );
  AOI21_X1 U12564 ( .B1(n10047), .B2(n15096), .A(n10046), .ZN(n10055) );
  INV_X1 U12565 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n14752) );
  AOI22_X1 U12566 ( .A1(n14337), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n14752), 
        .B2(n10048), .ZN(n10052) );
  INV_X1 U12567 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10050) );
  MUX2_X1 U12568 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10050), .S(n11378), .Z(
        n15003) );
  NAND2_X1 U12569 ( .A1(n15004), .A2(n15003), .ZN(n15002) );
  OAI21_X1 U12570 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n11378), .A(n15002), 
        .ZN(n10051) );
  NAND2_X1 U12571 ( .A1(n10052), .A2(n10051), .ZN(n14336) );
  OAI21_X1 U12572 ( .B1(n10052), .B2(n10051), .A(n14336), .ZN(n10053) );
  NAND2_X1 U12573 ( .A1(n10053), .A2(n15091), .ZN(n10054) );
  NAND2_X1 U12574 ( .A1(n10055), .A2(n10054), .ZN(P1_U3255) );
  INV_X1 U12575 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10061) );
  INV_X1 U12576 ( .A(n10667), .ZN(n10058) );
  INV_X1 U12577 ( .A(n14219), .ZN(n10056) );
  OAI21_X1 U12578 ( .B1(n15191), .B2(n14971), .A(n10056), .ZN(n10057) );
  OR2_X1 U12579 ( .A1(n10072), .A2(n14533), .ZN(n10665) );
  OAI211_X1 U12580 ( .C1(n10059), .C2(n10058), .A(n10057), .B(n10665), .ZN(
        n14671) );
  NAND2_X1 U12581 ( .A1(n14671), .A2(n15194), .ZN(n10060) );
  OAI21_X1 U12582 ( .B1(n15194), .B2(n10061), .A(n10060), .ZN(P1_U3459) );
  OAI22_X1 U12583 ( .A1(n10062), .A2(n6646), .B1(n6840), .B2(n12338), .ZN(
        n10517) );
  NAND2_X1 U12584 ( .A1(n14280), .A2(n11048), .ZN(n10064) );
  NAND2_X1 U12585 ( .A1(n12329), .A2(n15118), .ZN(n10063) );
  NAND2_X1 U12586 ( .A1(n10064), .A2(n10063), .ZN(n10065) );
  XNOR2_X1 U12587 ( .A(n10065), .B(n10525), .ZN(n10518) );
  XOR2_X1 U12588 ( .A(n10517), .B(n10518), .Z(n10070) );
  INV_X1 U12589 ( .A(n10066), .ZN(n10067) );
  NAND2_X1 U12590 ( .A1(n10068), .A2(n10067), .ZN(n10069) );
  OAI21_X1 U12591 ( .B1(n10070), .B2(n10069), .A(n10520), .ZN(n10071) );
  NAND2_X1 U12592 ( .A1(n10071), .A2(n13994), .ZN(n10075) );
  INV_X1 U12593 ( .A(n13918), .ZN(n13987) );
  OAI22_X1 U12594 ( .A1(n10072), .A2(n14531), .B1(n10515), .B2(n14533), .ZN(
        n15112) );
  AOI22_X1 U12595 ( .A1(n13987), .A2(n15112), .B1(n10073), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n10074) );
  OAI211_X1 U12596 ( .C1(n6840), .C2(n14005), .A(n10075), .B(n10074), .ZN(
        P1_U3237) );
  AOI21_X1 U12597 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n10079), .A(n10076), 
        .ZN(n10694) );
  INV_X1 U12598 ( .A(n10694), .ZN(n10077) );
  XNOR2_X1 U12599 ( .A(n10077), .B(n10704), .ZN(n10692) );
  XOR2_X1 U12600 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n10692), .Z(n10087) );
  NAND2_X1 U12601 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n11462)
         );
  AOI21_X1 U12602 ( .B1(n10079), .B2(P2_REG1_REG_13__SCAN_IN), .A(n10078), 
        .ZN(n10081) );
  INV_X1 U12603 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n14883) );
  MUX2_X1 U12604 ( .A(n14883), .B(P2_REG1_REG_14__SCAN_IN), .S(n10704), .Z(
        n10080) );
  NOR2_X1 U12605 ( .A1(n10081), .A2(n10080), .ZN(n10703) );
  AOI211_X1 U12606 ( .C1(n10081), .C2(n10080), .A(n10703), .B(n15225), .ZN(
        n10082) );
  INV_X1 U12607 ( .A(n10082), .ZN(n10083) );
  NAND2_X1 U12608 ( .A1(n11462), .A2(n10083), .ZN(n10085) );
  NOR2_X1 U12609 ( .A1(n15278), .A2(n10693), .ZN(n10084) );
  AOI211_X1 U12610 ( .C1(n15270), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n10085), 
        .B(n10084), .ZN(n10086) );
  OAI21_X1 U12611 ( .B1(n10087), .B2(n15220), .A(n10086), .ZN(P2_U3228) );
  NAND2_X1 U12612 ( .A1(n10088), .A2(n10482), .ZN(n10090) );
  AND2_X1 U12613 ( .A1(n10092), .A2(n10090), .ZN(n10094) );
  XNOR2_X1 U12614 ( .A(n10089), .B(n15487), .ZN(n10268) );
  XNOR2_X1 U12615 ( .A(n10268), .B(n12549), .ZN(n10093) );
  AND2_X1 U12616 ( .A1(n10093), .A2(n10090), .ZN(n10091) );
  NAND2_X1 U12617 ( .A1(n10092), .A2(n10091), .ZN(n10271) );
  OAI211_X1 U12618 ( .C1(n10094), .C2(n10093), .A(n12522), .B(n10271), .ZN(
        n10097) );
  NOR2_X1 U12619 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10488), .ZN(n10439) );
  OAI22_X1 U12620 ( .A1(n10482), .A2(n12527), .B1(n12526), .B2(n12063), .ZN(
        n10095) );
  AOI211_X1 U12621 ( .C1(n15487), .C2(n12517), .A(n10439), .B(n10095), .ZN(
        n10096) );
  OAI211_X1 U12622 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n11236), .A(n10097), .B(
        n10096), .ZN(P3_U3158) );
  INV_X1 U12623 ( .A(n10098), .ZN(n10099) );
  XNOR2_X1 U12624 ( .A(n11968), .B(n10292), .ZN(n10365) );
  NOR2_X1 U12625 ( .A1(n11966), .A2(n10291), .ZN(n10366) );
  XNOR2_X1 U12626 ( .A(n10365), .B(n10366), .ZN(n10367) );
  XNOR2_X1 U12627 ( .A(n10368), .B(n10367), .ZN(n10107) );
  NAND2_X1 U12628 ( .A1(n13475), .A2(n13529), .ZN(n10102) );
  OR2_X1 U12629 ( .A1(n13492), .A2(n10607), .ZN(n10101) );
  AND2_X1 U12630 ( .A1(n10102), .A2(n10101), .ZN(n10241) );
  OAI21_X1 U12631 ( .B1(n13476), .B2(n10241), .A(n10103), .ZN(n10105) );
  NOR2_X1 U12632 ( .A1(n13461), .A2(n7314), .ZN(n10104) );
  AOI211_X1 U12633 ( .C1(n13467), .C2(n10247), .A(n10105), .B(n10104), .ZN(
        n10106) );
  OAI21_X1 U12634 ( .B1(n10107), .B2(n13503), .A(n10106), .ZN(P2_U3211) );
  INV_X1 U12635 ( .A(n10108), .ZN(n10111) );
  OAI222_X1 U12636 ( .A1(n14722), .A2(n10111), .B1(n14721), .B2(n10110), .C1(
        P3_U3151), .C2(n10109), .ZN(P3_U3275) );
  INV_X1 U12637 ( .A(n10112), .ZN(n10113) );
  NAND2_X1 U12638 ( .A1(n10113), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10116) );
  INV_X1 U12639 ( .A(n12526), .ZN(n11608) );
  AOI22_X1 U12640 ( .A1(n11608), .A2(n9997), .B1(n12517), .B2(n10114), .ZN(
        n10115) );
  OAI211_X1 U12641 ( .C1(n10117), .C2(n12520), .A(n10116), .B(n10115), .ZN(
        P3_U3172) );
  INV_X1 U12642 ( .A(n11685), .ZN(n10121) );
  NAND2_X1 U12643 ( .A1(n10118), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10119) );
  XNOR2_X1 U12644 ( .A(n10119), .B(n7567), .ZN(n15099) );
  OAI222_X1 U12645 ( .A1(n14694), .A2(n10120), .B1(n11910), .B2(n10121), .C1(
        P1_U3086), .C2(n15099), .ZN(P1_U3337) );
  INV_X1 U12646 ( .A(n11596), .ZN(n11189) );
  OAI222_X1 U12647 ( .A1(n13852), .A2(n10122), .B1(n13854), .B2(n10121), .C1(
        P2_U3088), .C2(n11189), .ZN(P2_U3309) );
  OR2_X1 U12648 ( .A1(n10125), .A2(P3_U3151), .ZN(n12192) );
  INV_X1 U12649 ( .A(n12192), .ZN(n10123) );
  NAND2_X1 U12650 ( .A1(n12171), .A2(n10125), .ZN(n10126) );
  AND2_X1 U12651 ( .A1(n10127), .A2(n10126), .ZN(n10173) );
  NAND2_X1 U12652 ( .A1(n10175), .A2(n10173), .ZN(n10142) );
  MUX2_X1 U12653 ( .A(n10142), .B(n12550), .S(n10128), .Z(n12645) );
  MUX2_X1 U12654 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n6642), .Z(n10448) );
  INV_X1 U12655 ( .A(n10458), .ZN(n10129) );
  XNOR2_X1 U12656 ( .A(n10448), .B(n10129), .ZN(n10141) );
  MUX2_X1 U12657 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n6642), .Z(n10130) );
  OR2_X1 U12658 ( .A1(n10130), .A2(n10428), .ZN(n10139) );
  XNOR2_X1 U12659 ( .A(n10130), .B(n10168), .ZN(n10414) );
  MUX2_X1 U12660 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n6642), .Z(n10131) );
  OR2_X1 U12661 ( .A1(n10131), .A2(n10167), .ZN(n10138) );
  XNOR2_X1 U12662 ( .A(n10131), .B(n10405), .ZN(n10394) );
  MUX2_X1 U12663 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n10132), .Z(n10133) );
  XNOR2_X1 U12664 ( .A(n10133), .B(n10253), .ZN(n10252) );
  INV_X1 U12665 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n12197) );
  MUX2_X1 U12666 ( .A(n10146), .B(n12197), .S(n6642), .Z(n15409) );
  OAI22_X1 U12667 ( .A1(n10252), .A2(n15406), .B1(n10133), .B2(n10253), .ZN(
        n10304) );
  MUX2_X1 U12668 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n6642), .Z(n10134) );
  XNOR2_X1 U12669 ( .A(n10134), .B(n6641), .ZN(n10305) );
  INV_X1 U12670 ( .A(n10134), .ZN(n10135) );
  MUX2_X1 U12671 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n6642), .Z(n10136) );
  XOR2_X1 U12672 ( .A(n10431), .B(n10136), .Z(n10429) );
  INV_X1 U12673 ( .A(n10429), .ZN(n10137) );
  NAND2_X1 U12674 ( .A1(n10394), .A2(n10395), .ZN(n10393) );
  NAND2_X1 U12675 ( .A1(n10138), .A2(n10393), .ZN(n10413) );
  NAND2_X1 U12676 ( .A1(n10414), .A2(n10413), .ZN(n10412) );
  NAND2_X1 U12677 ( .A1(n10139), .A2(n10412), .ZN(n10140) );
  NAND2_X1 U12678 ( .A1(n10141), .A2(n10140), .ZN(n10449) );
  OAI21_X1 U12679 ( .B1(n10141), .B2(n10140), .A(n10449), .ZN(n10180) );
  INV_X1 U12680 ( .A(n10142), .ZN(n10159) );
  INV_X1 U12681 ( .A(n10143), .ZN(n10144) );
  NOR2_X1 U12682 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n10146), .ZN(n15403) );
  NAND2_X1 U12683 ( .A1(n10145), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10147) );
  OAI21_X1 U12684 ( .B1(n10253), .B2(n15403), .A(n10147), .ZN(n10255) );
  INV_X1 U12685 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n15476) );
  AOI21_X1 U12686 ( .B1(n10145), .B2(P3_REG2_REG_0__SCAN_IN), .A(n10254), .ZN(
        n10307) );
  XNOR2_X1 U12687 ( .A(n10317), .B(n10148), .ZN(n10308) );
  NOR2_X1 U12688 ( .A1(n10307), .A2(n10308), .ZN(n10306) );
  INV_X1 U12689 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10434) );
  NAND2_X1 U12690 ( .A1(P3_REG2_REG_4__SCAN_IN), .A2(n10167), .ZN(n10153) );
  OAI21_X1 U12691 ( .B1(P3_REG2_REG_4__SCAN_IN), .B2(n10167), .A(n10153), .ZN(
        n10397) );
  NOR2_X1 U12692 ( .A1(n10398), .A2(n10397), .ZN(n10396) );
  AOI21_X1 U12693 ( .B1(P3_REG2_REG_4__SCAN_IN), .B2(n10167), .A(n10396), .ZN(
        n10154) );
  NOR2_X1 U12694 ( .A1(n10168), .A2(n10154), .ZN(n10155) );
  INV_X1 U12695 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n10417) );
  XNOR2_X1 U12696 ( .A(n10154), .B(n10168), .ZN(n10416) );
  NAND2_X1 U12697 ( .A1(P3_REG2_REG_6__SCAN_IN), .A2(n10458), .ZN(n10156) );
  OAI21_X1 U12698 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n10458), .A(n10156), .ZN(
        n10157) );
  AOI21_X1 U12699 ( .B1(n6787), .B2(n10157), .A(n10445), .ZN(n10158) );
  NOR2_X1 U12700 ( .A1(n15438), .A2(n10158), .ZN(n10179) );
  INV_X1 U12701 ( .A(n15402), .ZN(n10160) );
  AOI22_X1 U12702 ( .A1(n10253), .A2(n10160), .B1(P3_IR_REG_1__SCAN_IN), .B2(
        n15402), .ZN(n10258) );
  INV_X1 U12703 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n15529) );
  NOR2_X1 U12704 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10160), .ZN(n10161) );
  NOR2_X1 U12705 ( .A1(n10257), .A2(n10161), .ZN(n10311) );
  XNOR2_X1 U12706 ( .A(n10317), .B(n10162), .ZN(n10312) );
  NOR2_X1 U12707 ( .A1(n10311), .A2(n10312), .ZN(n10310) );
  INV_X1 U12708 ( .A(n10164), .ZN(n10165) );
  INV_X1 U12709 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15532) );
  NAND2_X1 U12710 ( .A1(P3_REG1_REG_4__SCAN_IN), .A2(n10167), .ZN(n10166) );
  OAI21_X1 U12711 ( .B1(P3_REG1_REG_4__SCAN_IN), .B2(n10167), .A(n10166), .ZN(
        n10400) );
  NOR2_X1 U12712 ( .A1(n10168), .A2(n10169), .ZN(n10170) );
  INV_X1 U12713 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15536) );
  NAND2_X1 U12714 ( .A1(P3_REG1_REG_6__SCAN_IN), .A2(n10458), .ZN(n10171) );
  OAI21_X1 U12715 ( .B1(P3_REG1_REG_6__SCAN_IN), .B2(n10458), .A(n10171), .ZN(
        n10172) );
  AOI21_X1 U12716 ( .B1(n6788), .B2(n10172), .A(n10460), .ZN(n10177) );
  INV_X1 U12717 ( .A(n10173), .ZN(n10174) );
  NAND2_X1 U12718 ( .A1(n10175), .A2(n10174), .ZN(n15421) );
  AND2_X1 U12719 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n10659) );
  AOI21_X1 U12720 ( .B1(n15405), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n10659), .ZN(
        n10176) );
  OAI21_X1 U12721 ( .B1(n15425), .B2(n10177), .A(n10176), .ZN(n10178) );
  AOI211_X1 U12722 ( .C1(n12652), .C2(n10180), .A(n10179), .B(n10178), .ZN(
        n10181) );
  OAI21_X1 U12723 ( .B1(n10458), .B2(n12645), .A(n10181), .ZN(P3_U3188) );
  INV_X1 U12724 ( .A(n10182), .ZN(n10183) );
  OR3_X1 U12725 ( .A1(n11020), .A2(n11019), .A3(n10183), .ZN(n10194) );
  OR2_X1 U12726 ( .A1(n15292), .A2(n7685), .ZN(n11625) );
  OR2_X1 U12727 ( .A1(n10194), .A2(n15342), .ZN(n10284) );
  NAND2_X1 U12728 ( .A1(n10186), .A2(n10185), .ZN(n10188) );
  INV_X1 U12729 ( .A(n13532), .ZN(n10201) );
  NAND2_X1 U12730 ( .A1(n15281), .A2(n10201), .ZN(n10187) );
  NAND2_X1 U12731 ( .A1(n10188), .A2(n10187), .ZN(n10347) );
  OR2_X1 U12732 ( .A1(n10359), .A2(n13531), .ZN(n10189) );
  NAND2_X1 U12733 ( .A1(n10217), .A2(n10218), .ZN(n10192) );
  NAND2_X1 U12734 ( .A1(n10229), .A2(n10208), .ZN(n10191) );
  XNOR2_X1 U12735 ( .A(n10234), .B(n10236), .ZN(n15334) );
  NOR2_X1 U12736 ( .A1(n10355), .A2(n10359), .ZN(n10358) );
  NAND2_X1 U12737 ( .A1(n10358), .A2(n10229), .ZN(n10225) );
  INV_X1 U12738 ( .A(n10246), .ZN(n10193) );
  AOI211_X1 U12739 ( .C1(n10239), .C2(n10225), .A(n13728), .B(n10193), .ZN(
        n15330) );
  INV_X1 U12740 ( .A(n10195), .ZN(n10196) );
  OAI22_X1 U12741 ( .A1(n15282), .A2(n15333), .B1(n14827), .B2(n10196), .ZN(
        n10197) );
  AOI21_X1 U12742 ( .B1(n15330), .B2(n15285), .A(n10197), .ZN(n10216) );
  NAND2_X1 U12743 ( .A1(n10199), .A2(n10198), .ZN(n10203) );
  NAND2_X1 U12744 ( .A1(n10201), .A2(n10200), .ZN(n10202) );
  NAND2_X1 U12745 ( .A1(n10203), .A2(n10202), .ZN(n10349) );
  NAND2_X1 U12746 ( .A1(n10349), .A2(n10346), .ZN(n10206) );
  NAND2_X1 U12747 ( .A1(n10359), .A2(n10204), .ZN(n10205) );
  NAND2_X1 U12748 ( .A1(n10206), .A2(n10205), .ZN(n10219) );
  INV_X1 U12749 ( .A(n10218), .ZN(n10207) );
  NAND2_X1 U12750 ( .A1(n10219), .A2(n10207), .ZN(n10210) );
  NAND2_X1 U12751 ( .A1(n15324), .A2(n10208), .ZN(n10209) );
  XNOR2_X1 U12752 ( .A(n10237), .B(n10236), .ZN(n10213) );
  INV_X1 U12753 ( .A(n10211), .ZN(n10212) );
  AOI21_X1 U12754 ( .B1(n10213), .B2(n14841), .A(n10212), .ZN(n15331) );
  MUX2_X1 U12755 ( .A(n10214), .B(n15331), .S(n13748), .Z(n10215) );
  OAI211_X1 U12756 ( .C1(n13738), .C2(n15334), .A(n10216), .B(n10215), .ZN(
        P2_U3260) );
  XNOR2_X1 U12757 ( .A(n10217), .B(n10218), .ZN(n10223) );
  INV_X1 U12758 ( .A(n10223), .ZN(n15327) );
  XNOR2_X1 U12759 ( .A(n10219), .B(n10218), .ZN(n10221) );
  OAI21_X1 U12760 ( .B1(n10221), .B2(n14819), .A(n10220), .ZN(n10222) );
  AOI21_X1 U12761 ( .B1(n11622), .B2(n10223), .A(n10222), .ZN(n15325) );
  MUX2_X1 U12762 ( .A(n10224), .B(n15325), .S(n13748), .Z(n10232) );
  INV_X1 U12763 ( .A(n10358), .ZN(n10227) );
  INV_X1 U12764 ( .A(n10225), .ZN(n10226) );
  AOI211_X1 U12765 ( .C1(n15324), .C2(n10227), .A(n13728), .B(n10226), .ZN(
        n15323) );
  OAI22_X1 U12766 ( .A1(n15282), .A2(n10229), .B1(n10228), .B2(n14827), .ZN(
        n10230) );
  AOI21_X1 U12767 ( .B1(n15323), .B2(n15285), .A(n10230), .ZN(n10231) );
  OAI211_X1 U12768 ( .C1(n15327), .C2(n11625), .A(n10232), .B(n10231), .ZN(
        P2_U3261) );
  INV_X1 U12769 ( .A(n10236), .ZN(n10233) );
  OR2_X1 U12770 ( .A1(n10239), .A2(n13529), .ZN(n10235) );
  XNOR2_X1 U12771 ( .A(n10286), .B(n10289), .ZN(n15341) );
  NAND2_X1 U12772 ( .A1(n10239), .A2(n10238), .ZN(n10240) );
  XNOR2_X1 U12773 ( .A(n10290), .B(n10289), .ZN(n10243) );
  INV_X1 U12774 ( .A(n10241), .ZN(n10242) );
  AOI21_X1 U12775 ( .B1(n10243), .B2(n14841), .A(n10242), .ZN(n15339) );
  MUX2_X1 U12776 ( .A(n10244), .B(n15339), .S(n13748), .Z(n10251) );
  INV_X1 U12777 ( .A(n10298), .ZN(n10245) );
  AOI211_X1 U12778 ( .C1(n10292), .C2(n10246), .A(n13728), .B(n10245), .ZN(
        n15338) );
  INV_X1 U12779 ( .A(n10247), .ZN(n10248) );
  OAI22_X1 U12780 ( .A1(n15282), .A2(n7314), .B1(n10248), .B2(n14827), .ZN(
        n10249) );
  AOI21_X1 U12781 ( .B1(n15338), .B2(n15285), .A(n10249), .ZN(n10250) );
  OAI211_X1 U12782 ( .C1(n13738), .C2(n15341), .A(n10251), .B(n10250), .ZN(
        P2_U3259) );
  XOR2_X1 U12783 ( .A(n15406), .B(n10252), .Z(n10265) );
  INV_X1 U12784 ( .A(n10253), .ZN(n10263) );
  AOI21_X1 U12785 ( .B1(n15476), .B2(n10255), .A(n10254), .ZN(n10256) );
  NOR2_X1 U12786 ( .A1(n15438), .A2(n10256), .ZN(n10262) );
  AOI21_X1 U12787 ( .B1(n10258), .B2(n15529), .A(n10257), .ZN(n10260) );
  AOI22_X1 U12788 ( .A1(n15405), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10259) );
  OAI21_X1 U12789 ( .B1(n10260), .B2(n15425), .A(n10259), .ZN(n10261) );
  AOI211_X1 U12790 ( .C1(n15430), .C2(n10263), .A(n10262), .B(n10261), .ZN(
        n10264) );
  OAI21_X1 U12791 ( .B1(n15434), .B2(n10265), .A(n10264), .ZN(P3_U3183) );
  INV_X1 U12792 ( .A(SI_21_), .ZN(n10266) );
  OAI222_X1 U12793 ( .A1(n14722), .A2(n10267), .B1(n14721), .B2(n10266), .C1(
        P3_U3151), .C2(n12049), .ZN(P3_U3274) );
  INV_X1 U12794 ( .A(n10268), .ZN(n10269) );
  NAND2_X1 U12795 ( .A1(n10269), .A2(n12549), .ZN(n10270) );
  NAND2_X1 U12796 ( .A1(n10271), .A2(n10270), .ZN(n10277) );
  XNOR2_X1 U12797 ( .A(n12416), .B(n10280), .ZN(n10272) );
  NAND2_X1 U12798 ( .A1(n10272), .A2(n12063), .ZN(n10469) );
  INV_X1 U12799 ( .A(n10272), .ZN(n10273) );
  NAND2_X1 U12800 ( .A1(n10273), .A2(n12548), .ZN(n10274) );
  NAND2_X1 U12801 ( .A1(n10469), .A2(n10274), .ZN(n10276) );
  INV_X1 U12802 ( .A(n10470), .ZN(n10275) );
  AOI21_X1 U12803 ( .B1(n10277), .B2(n10276), .A(n10275), .ZN(n10283) );
  INV_X1 U12804 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n10278) );
  NOR2_X1 U12805 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10278), .ZN(n10404) );
  OAI22_X1 U12806 ( .A1(n15449), .A2(n12527), .B1(n12526), .B2(n10963), .ZN(
        n10279) );
  AOI211_X1 U12807 ( .C1(n10280), .C2(n12517), .A(n10404), .B(n10279), .ZN(
        n10282) );
  NAND2_X1 U12808 ( .A1(n12530), .A2(n10382), .ZN(n10281) );
  OAI211_X1 U12809 ( .C1(n10283), .C2(n12520), .A(n10282), .B(n10281), .ZN(
        P3_U3170) );
  INV_X1 U12810 ( .A(n10289), .ZN(n10285) );
  OR2_X1 U12811 ( .A1(n10292), .A2(n13528), .ZN(n10287) );
  XOR2_X1 U12812 ( .A(n10600), .B(n10599), .Z(n15351) );
  XOR2_X1 U12813 ( .A(n10609), .B(n10599), .Z(n10296) );
  NAND2_X1 U12814 ( .A1(n13475), .A2(n13528), .ZN(n10294) );
  OR2_X1 U12815 ( .A1(n13492), .A2(n10610), .ZN(n10293) );
  AND2_X1 U12816 ( .A1(n10294), .A2(n10293), .ZN(n10369) );
  INV_X1 U12817 ( .A(n10369), .ZN(n10295) );
  AOI21_X1 U12818 ( .B1(n10296), .B2(n14841), .A(n10295), .ZN(n15348) );
  MUX2_X1 U12819 ( .A(n10297), .B(n15348), .S(n13748), .Z(n10303) );
  AOI211_X1 U12820 ( .C1(n15347), .C2(n10298), .A(n13728), .B(n10680), .ZN(
        n15346) );
  INV_X1 U12821 ( .A(n15347), .ZN(n10300) );
  INV_X1 U12822 ( .A(n10371), .ZN(n10299) );
  OAI22_X1 U12823 ( .A1(n15282), .A2(n10300), .B1(n14827), .B2(n10299), .ZN(
        n10301) );
  AOI21_X1 U12824 ( .B1(n15346), .B2(n15285), .A(n10301), .ZN(n10302) );
  OAI211_X1 U12825 ( .C1(n13738), .C2(n15351), .A(n10303), .B(n10302), .ZN(
        P2_U3258) );
  XOR2_X1 U12826 ( .A(n10305), .B(n10304), .Z(n10319) );
  AOI21_X1 U12827 ( .B1(n10308), .B2(n10307), .A(n10306), .ZN(n10309) );
  NOR2_X1 U12828 ( .A1(n15438), .A2(n10309), .ZN(n10316) );
  AOI21_X1 U12829 ( .B1(n10312), .B2(n10311), .A(n10310), .ZN(n10314) );
  AOI22_X1 U12830 ( .A1(n15405), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10313) );
  OAI21_X1 U12831 ( .B1(n10314), .B2(n15425), .A(n10313), .ZN(n10315) );
  AOI211_X1 U12832 ( .C1(n15430), .C2(n6641), .A(n10316), .B(n10315), .ZN(
        n10318) );
  OAI21_X1 U12833 ( .B1(n10319), .B2(n15434), .A(n10318), .ZN(P3_U3184) );
  OR2_X1 U12834 ( .A1(n14025), .A2(n10321), .ZN(n10323) );
  OR2_X1 U12835 ( .A1(n6649), .A2(n6913), .ZN(n10322) );
  OAI21_X1 U12836 ( .B1(n10325), .B2(n14224), .A(n10550), .ZN(n10642) );
  INV_X1 U12837 ( .A(n10642), .ZN(n10344) );
  INV_X1 U12838 ( .A(n14053), .ZN(n10536) );
  NAND2_X1 U12839 ( .A1(n14278), .A2(n10536), .ZN(n10326) );
  NAND2_X1 U12840 ( .A1(n10327), .A2(n10326), .ZN(n10330) );
  INV_X1 U12841 ( .A(n14278), .ZN(n10328) );
  NAND2_X1 U12842 ( .A1(n10328), .A2(n14053), .ZN(n10329) );
  NAND2_X1 U12843 ( .A1(n10330), .A2(n10329), .ZN(n10563) );
  XNOR2_X1 U12844 ( .A(n10563), .B(n10562), .ZN(n10339) );
  NAND2_X1 U12845 ( .A1(n14278), .A2(n14571), .ZN(n10338) );
  NAND2_X1 U12846 ( .A1(n11774), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10336) );
  NAND2_X1 U12847 ( .A1(n10331), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10812) );
  OAI21_X1 U12848 ( .B1(n10331), .B2(P1_REG3_REG_6__SCAN_IN), .A(n10812), .ZN(
        n13977) );
  INV_X1 U12849 ( .A(n13977), .ZN(n10332) );
  NAND2_X1 U12850 ( .A1(n11751), .A2(n10332), .ZN(n10335) );
  NAND2_X1 U12851 ( .A1(n11093), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10334) );
  NAND2_X1 U12852 ( .A1(n14012), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n10333) );
  NAND4_X1 U12853 ( .A1(n10336), .A2(n10335), .A3(n10334), .A4(n10333), .ZN(
        n14276) );
  NAND2_X1 U12854 ( .A1(n14276), .A2(n14573), .ZN(n10337) );
  NAND2_X1 U12855 ( .A1(n10338), .A2(n10337), .ZN(n11058) );
  AOI21_X1 U12856 ( .B1(n10339), .B2(n14971), .A(n11058), .ZN(n10645) );
  NAND2_X1 U12857 ( .A1(n10340), .A2(n14062), .ZN(n10341) );
  NAND2_X1 U12858 ( .A1(n10341), .A2(n15120), .ZN(n10342) );
  NOR2_X1 U12859 ( .A1(n10575), .A2(n10342), .ZN(n10641) );
  AOI21_X1 U12860 ( .B1(n14062), .B2(n14955), .A(n10641), .ZN(n10343) );
  OAI211_X1 U12861 ( .C1(n10344), .C2(n14670), .A(n10645), .B(n10343), .ZN(
        n10362) );
  NAND2_X1 U12862 ( .A1(n10362), .A2(n15202), .ZN(n10345) );
  OAI21_X1 U12863 ( .B1(n15202), .B2(n9727), .A(n10345), .ZN(P1_U3533) );
  XNOR2_X1 U12864 ( .A(n10347), .B(n10346), .ZN(n15316) );
  INV_X1 U12865 ( .A(n15317), .ZN(n10351) );
  XNOR2_X1 U12866 ( .A(n10348), .B(n10349), .ZN(n10350) );
  NOR2_X1 U12867 ( .A1(n10350), .A2(n14819), .ZN(n15320) );
  AOI211_X1 U12868 ( .C1(n15279), .C2(n10352), .A(n10351), .B(n15320), .ZN(
        n10353) );
  MUX2_X1 U12869 ( .A(n10354), .B(n10353), .S(n13748), .Z(n10361) );
  NAND2_X1 U12870 ( .A1(n10355), .A2(n10359), .ZN(n10356) );
  NAND2_X1 U12871 ( .A1(n10356), .A2(n14852), .ZN(n10357) );
  NOR2_X1 U12872 ( .A1(n10358), .A2(n10357), .ZN(n15319) );
  AOI22_X1 U12873 ( .A1(n14844), .A2(n10359), .B1(n15319), .B2(n15285), .ZN(
        n10360) );
  OAI211_X1 U12874 ( .C1(n13738), .C2(n15316), .A(n10361), .B(n10360), .ZN(
        P2_U3262) );
  INV_X1 U12875 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10364) );
  NAND2_X1 U12876 ( .A1(n10362), .A2(n15194), .ZN(n10363) );
  OAI21_X1 U12877 ( .B1(n15194), .B2(n10364), .A(n10363), .ZN(P1_U3474) );
  XNOR2_X1 U12878 ( .A(n15347), .B(n11968), .ZN(n10583) );
  NAND2_X1 U12879 ( .A1(n9669), .A2(n13527), .ZN(n10582) );
  XNOR2_X1 U12880 ( .A(n10583), .B(n10582), .ZN(n10585) );
  XNOR2_X1 U12881 ( .A(n10586), .B(n10585), .ZN(n10374) );
  OAI22_X1 U12882 ( .A1(n13476), .A2(n10369), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13547), .ZN(n10370) );
  AOI21_X1 U12883 ( .B1(n10371), .B2(n13467), .A(n10370), .ZN(n10373) );
  NAND2_X1 U12884 ( .A1(n13501), .A2(n15347), .ZN(n10372) );
  OAI211_X1 U12885 ( .C1(n10374), .C2(n13503), .A(n10373), .B(n10372), .ZN(
        P2_U3185) );
  NAND2_X1 U12886 ( .A1(n12044), .A2(n15444), .ZN(n10481) );
  NAND2_X1 U12887 ( .A1(n15470), .A2(n10481), .ZN(n14779) );
  NAND2_X1 U12888 ( .A1(n15477), .A2(n14779), .ZN(n12888) );
  XNOR2_X1 U12889 ( .A(n10375), .B(n12061), .ZN(n15493) );
  INV_X1 U12890 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10381) );
  INV_X1 U12891 ( .A(n10376), .ZN(n10377) );
  AOI21_X1 U12892 ( .B1(n10377), .B2(n12020), .A(n15456), .ZN(n10380) );
  OAI22_X1 U12893 ( .A1(n15449), .A2(n15450), .B1(n10963), .B2(n15448), .ZN(
        n10378) );
  AOI21_X1 U12894 ( .B1(n10380), .B2(n10379), .A(n10378), .ZN(n15494) );
  MUX2_X1 U12895 ( .A(n10381), .B(n15494), .S(n15477), .Z(n10384) );
  INV_X1 U12896 ( .A(n12794), .ZN(n14782) );
  NOR2_X1 U12897 ( .A1(n12064), .A2(n15521), .ZN(n15496) );
  AOI22_X1 U12898 ( .A1(n14782), .A2(n15496), .B1(n15473), .B2(n10382), .ZN(
        n10383) );
  OAI211_X1 U12899 ( .C1(n12888), .C2(n15493), .A(n10384), .B(n10383), .ZN(
        P3_U3229) );
  INV_X1 U12900 ( .A(n11698), .ZN(n10624) );
  OAI222_X1 U12901 ( .A1(n11910), .A2(n10624), .B1(P1_U3086), .B2(n14352), 
        .C1(n10385), .C2(n14694), .ZN(P1_U3336) );
  AOI22_X1 U12902 ( .A1(n15285), .A2(n10386), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n15279), .ZN(n10388) );
  NAND2_X1 U12903 ( .A1(n15292), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10387) );
  AOI21_X1 U12904 ( .B1(n10390), .B2(n15288), .A(n10389), .ZN(n10391) );
  OAI21_X1 U12905 ( .B1(n15292), .B2(n10392), .A(n10391), .ZN(P2_U3264) );
  OAI21_X1 U12906 ( .B1(n10395), .B2(n10394), .A(n10393), .ZN(n10410) );
  AOI21_X1 U12907 ( .B1(n10398), .B2(n10397), .A(n10396), .ZN(n10408) );
  AOI21_X1 U12908 ( .B1(n10401), .B2(n10400), .A(n10399), .ZN(n10402) );
  NOR2_X1 U12909 ( .A1(n15425), .A2(n10402), .ZN(n10403) );
  AOI211_X1 U12910 ( .C1(n15405), .C2(P3_ADDR_REG_4__SCAN_IN), .A(n10404), .B(
        n10403), .ZN(n10407) );
  NAND2_X1 U12911 ( .A1(n15430), .A2(n10405), .ZN(n10406) );
  OAI211_X1 U12912 ( .C1(n10408), .C2(n15438), .A(n10407), .B(n10406), .ZN(
        n10409) );
  AOI21_X1 U12913 ( .B1(n12652), .B2(n10410), .A(n10409), .ZN(n10411) );
  INV_X1 U12914 ( .A(n10411), .ZN(P3_U3186) );
  OAI21_X1 U12915 ( .B1(n10414), .B2(n10413), .A(n10412), .ZN(n10426) );
  AOI21_X1 U12916 ( .B1(n10417), .B2(n10416), .A(n10415), .ZN(n10424) );
  NOR2_X1 U12917 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10418), .ZN(n10475) );
  AOI21_X1 U12918 ( .B1(n15536), .B2(n10420), .A(n10419), .ZN(n10421) );
  NOR2_X1 U12919 ( .A1(n15425), .A2(n10421), .ZN(n10422) );
  AOI211_X1 U12920 ( .C1(n15405), .C2(P3_ADDR_REG_5__SCAN_IN), .A(n10475), .B(
        n10422), .ZN(n10423) );
  OAI21_X1 U12921 ( .B1(n10424), .B2(n15438), .A(n10423), .ZN(n10425) );
  AOI21_X1 U12922 ( .B1(n12652), .B2(n10426), .A(n10425), .ZN(n10427) );
  OAI21_X1 U12923 ( .B1(n10428), .B2(n12645), .A(n10427), .ZN(P3_U3187) );
  XNOR2_X1 U12924 ( .A(n10430), .B(n10429), .ZN(n10444) );
  AOI21_X1 U12925 ( .B1(n10434), .B2(n10433), .A(n10432), .ZN(n10441) );
  AOI21_X1 U12926 ( .B1(n15532), .B2(n10436), .A(n10435), .ZN(n10437) );
  NOR2_X1 U12927 ( .A1(n15425), .A2(n10437), .ZN(n10438) );
  AOI211_X1 U12928 ( .C1(n15405), .C2(P3_ADDR_REG_3__SCAN_IN), .A(n10439), .B(
        n10438), .ZN(n10440) );
  OAI21_X1 U12929 ( .B1(n10441), .B2(n15438), .A(n10440), .ZN(n10442) );
  AOI21_X1 U12930 ( .B1(n10150), .B2(n15430), .A(n10442), .ZN(n10443) );
  OAI21_X1 U12931 ( .B1(n10444), .B2(n15434), .A(n10443), .ZN(P3_U3185) );
  NAND2_X1 U12932 ( .A1(n10446), .A2(n10502), .ZN(n10492) );
  INV_X1 U12933 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n10952) );
  AOI21_X1 U12934 ( .B1(n10447), .B2(n10952), .A(n10493), .ZN(n10467) );
  INV_X1 U12935 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n10457) );
  MUX2_X1 U12936 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n6642), .Z(n10503) );
  XOR2_X1 U12937 ( .A(n10502), .B(n10503), .Z(n10452) );
  OR2_X1 U12938 ( .A1(n10448), .A2(n10458), .ZN(n10450) );
  NAND2_X1 U12939 ( .A1(n10450), .A2(n10449), .ZN(n10451) );
  NAND2_X1 U12940 ( .A1(n10452), .A2(n10451), .ZN(n10504) );
  OAI21_X1 U12941 ( .B1(n10452), .B2(n10451), .A(n10504), .ZN(n10453) );
  NAND2_X1 U12942 ( .A1(n10453), .A2(n12652), .ZN(n10456) );
  INV_X1 U12943 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n10454) );
  NOR2_X1 U12944 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10454), .ZN(n10777) );
  INV_X1 U12945 ( .A(n10777), .ZN(n10455) );
  OAI211_X1 U12946 ( .C1(n15421), .C2(n10457), .A(n10456), .B(n10455), .ZN(
        n10465) );
  AND2_X1 U12947 ( .A1(n10458), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n10459) );
  INV_X1 U12948 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15540) );
  AOI21_X1 U12949 ( .B1(n10462), .B2(n15540), .A(n6790), .ZN(n10463) );
  NOR2_X1 U12950 ( .A1(n10463), .A2(n15425), .ZN(n10464) );
  AOI211_X1 U12951 ( .C1(n15430), .C2(n6990), .A(n10465), .B(n10464), .ZN(
        n10466) );
  OAI21_X1 U12952 ( .B1(n10467), .B2(n15438), .A(n10466), .ZN(P3_U3189) );
  INV_X1 U12953 ( .A(n10983), .ZN(n10479) );
  XNOR2_X1 U12954 ( .A(n12416), .B(n10476), .ZN(n10655) );
  XNOR2_X1 U12955 ( .A(n10655), .B(n10468), .ZN(n10472) );
  OAI21_X1 U12956 ( .B1(n10472), .B2(n10471), .A(n10834), .ZN(n10473) );
  NAND2_X1 U12957 ( .A1(n10473), .A2(n12522), .ZN(n10478) );
  OAI22_X1 U12958 ( .A1(n12063), .A2(n12527), .B1(n12526), .B2(n10947), .ZN(
        n10474) );
  AOI211_X1 U12959 ( .C1(n10476), .C2(n12517), .A(n10475), .B(n10474), .ZN(
        n10477) );
  OAI211_X1 U12960 ( .C1(n10479), .C2(n11236), .A(n10478), .B(n10477), .ZN(
        P3_U3167) );
  XNOR2_X1 U12961 ( .A(n10480), .B(n12019), .ZN(n15489) );
  INV_X1 U12962 ( .A(n15489), .ZN(n10491) );
  INV_X1 U12963 ( .A(n10481), .ZN(n15458) );
  INV_X1 U12964 ( .A(n15470), .ZN(n15453) );
  OAI22_X1 U12965 ( .A1(n10482), .A2(n15450), .B1(n12063), .B2(n15448), .ZN(
        n10487) );
  INV_X1 U12966 ( .A(n10483), .ZN(n10484) );
  AOI211_X1 U12967 ( .C1(n12019), .C2(n10485), .A(n15456), .B(n10484), .ZN(
        n10486) );
  AOI211_X1 U12968 ( .C1(n15489), .C2(n15453), .A(n10487), .B(n10486), .ZN(
        n15491) );
  MUX2_X1 U12969 ( .A(n10434), .B(n15491), .S(n15477), .Z(n10490) );
  AOI22_X1 U12970 ( .A1(n12885), .A2(n15487), .B1(n15473), .B2(n10488), .ZN(
        n10489) );
  OAI211_X1 U12971 ( .C1(n10491), .C2(n12752), .A(n10490), .B(n10489), .ZN(
        P3_U3230) );
  INV_X1 U12972 ( .A(n10492), .ZN(n10494) );
  NAND2_X1 U12973 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n10928), .ZN(n10495) );
  OAI21_X1 U12974 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n10928), .A(n10495), .ZN(
        n10496) );
  AOI21_X1 U12975 ( .B1(n6792), .B2(n10496), .A(n10916), .ZN(n10514) );
  NAND2_X1 U12976 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n10928), .ZN(n10498) );
  OAI21_X1 U12977 ( .B1(P3_REG1_REG_8__SCAN_IN), .B2(n10928), .A(n10498), .ZN(
        n10499) );
  AOI21_X1 U12978 ( .B1(n10500), .B2(n10499), .A(n10927), .ZN(n10501) );
  NOR2_X1 U12979 ( .A1(n10501), .A2(n15425), .ZN(n10512) );
  AND2_X1 U12980 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n12428) );
  AOI21_X1 U12981 ( .B1(n15405), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n12428), .ZN(
        n10510) );
  MUX2_X1 U12982 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n6642), .Z(n10919) );
  XOR2_X1 U12983 ( .A(n10928), .B(n10919), .Z(n10507) );
  OR2_X1 U12984 ( .A1(n10503), .A2(n10502), .ZN(n10505) );
  NAND2_X1 U12985 ( .A1(n10505), .A2(n10504), .ZN(n10506) );
  NAND2_X1 U12986 ( .A1(n10507), .A2(n10506), .ZN(n10918) );
  OAI21_X1 U12987 ( .B1(n10507), .B2(n10506), .A(n10918), .ZN(n10508) );
  NAND2_X1 U12988 ( .A1(n10508), .A2(n12652), .ZN(n10509) );
  OAI211_X1 U12989 ( .C1(n12645), .C2(n10928), .A(n10510), .B(n10509), .ZN(
        n10511) );
  NOR2_X1 U12990 ( .A1(n10512), .A2(n10511), .ZN(n10513) );
  OAI21_X1 U12991 ( .B1(n10514), .B2(n15438), .A(n10513), .ZN(P3_U3190) );
  OAI22_X1 U12992 ( .A1(n10515), .A2(n6646), .B1(n15179), .B2(n12338), .ZN(
        n10522) );
  OAI22_X1 U12993 ( .A1(n10515), .A2(n12338), .B1(n15179), .B2(n12340), .ZN(
        n10516) );
  XNOR2_X1 U12994 ( .A(n10516), .B(n10525), .ZN(n10521) );
  XNOR2_X1 U12995 ( .A(n10521), .B(n10522), .ZN(n10545) );
  NAND2_X1 U12996 ( .A1(n14278), .A2(n6638), .ZN(n10524) );
  NAND2_X1 U12997 ( .A1(n6640), .A2(n14053), .ZN(n10523) );
  NAND2_X1 U12998 ( .A1(n10524), .A2(n10523), .ZN(n10526) );
  XNOR2_X1 U12999 ( .A(n10526), .B(n12242), .ZN(n11034) );
  NOR2_X1 U13000 ( .A1(n12338), .A2(n10536), .ZN(n10527) );
  AOI21_X1 U13001 ( .B1(n12333), .B2(n14278), .A(n10527), .ZN(n11033) );
  XNOR2_X1 U13002 ( .A(n11034), .B(n11033), .ZN(n10528) );
  XNOR2_X1 U13003 ( .A(n11032), .B(n10528), .ZN(n10539) );
  NAND3_X1 U13004 ( .A1(n10531), .A2(n10530), .A3(n10529), .ZN(n10532) );
  NAND2_X1 U13005 ( .A1(n10532), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10533) );
  NAND2_X1 U13006 ( .A1(n13987), .A2(n10717), .ZN(n10534) );
  OAI211_X1 U13007 ( .C1(n14005), .C2(n10536), .A(n10535), .B(n10534), .ZN(
        n10537) );
  AOI21_X1 U13008 ( .B1(n10716), .B2(n14001), .A(n10537), .ZN(n10538) );
  OAI21_X1 U13009 ( .B1(n10539), .B2(n14932), .A(n10538), .ZN(P1_U3230) );
  NAND2_X1 U13010 ( .A1(n14280), .A2(n14571), .ZN(n10541) );
  NAND2_X1 U13011 ( .A1(n14278), .A2(n14573), .ZN(n10540) );
  NAND2_X1 U13012 ( .A1(n10541), .A2(n10540), .ZN(n10647) );
  AOI22_X1 U13013 ( .A1(n13987), .A2(n10647), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10542) );
  OAI21_X1 U13014 ( .B1(n14005), .B2(n15179), .A(n10542), .ZN(n10547) );
  AOI211_X1 U13015 ( .C1(n10545), .C2(n10544), .A(n14932), .B(n10543), .ZN(
        n10546) );
  AOI211_X1 U13016 ( .C1(n9943), .C2(n14001), .A(n10547), .B(n10546), .ZN(
        n10548) );
  INV_X1 U13017 ( .A(n10548), .ZN(P1_U3218) );
  NAND2_X1 U13018 ( .A1(n6897), .A2(n11060), .ZN(n10549) );
  NAND2_X1 U13019 ( .A1(n10550), .A2(n10549), .ZN(n10556) );
  NAND2_X1 U13020 ( .A1(n10551), .A2(n14017), .ZN(n10554) );
  OR2_X1 U13021 ( .A1(n6649), .A2(n10552), .ZN(n10553) );
  OAI211_X1 U13022 ( .C1(n6845), .C2(n10555), .A(n10554), .B(n10553), .ZN(
        n14071) );
  XNOR2_X1 U13023 ( .A(n14276), .B(n14071), .ZN(n14225) );
  NAND2_X1 U13024 ( .A1(n10556), .A2(n10565), .ZN(n10798) );
  OAI21_X1 U13025 ( .B1(n10556), .B2(n10565), .A(n10798), .ZN(n10750) );
  INV_X1 U13026 ( .A(n10750), .ZN(n10581) );
  INV_X1 U13027 ( .A(n10557), .ZN(n10561) );
  AND2_X1 U13028 ( .A1(n10559), .A2(n10558), .ZN(n10560) );
  NAND2_X1 U13029 ( .A1(n14038), .A2(n14579), .ZN(n14023) );
  OR2_X1 U13030 ( .A1(n15129), .A2(n14023), .ZN(n10936) );
  NAND2_X1 U13031 ( .A1(n6897), .A2(n14062), .ZN(n10564) );
  XNOR2_X1 U13032 ( .A(n10807), .B(n10565), .ZN(n10572) );
  INV_X1 U13033 ( .A(n11129), .ZN(n15183) );
  NAND2_X1 U13034 ( .A1(n10750), .A2(n15183), .ZN(n10571) );
  XNOR2_X1 U13035 ( .A(n10812), .B(P1_REG3_REG_7__SCAN_IN), .ZN(n11028) );
  NAND2_X1 U13036 ( .A1(n11751), .A2(n11028), .ZN(n10569) );
  NAND2_X1 U13037 ( .A1(n11774), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10568) );
  NAND2_X1 U13038 ( .A1(n14012), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n10567) );
  NAND2_X1 U13039 ( .A1(n11093), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10566) );
  NAND4_X1 U13040 ( .A1(n10569), .A2(n10568), .A3(n10567), .A4(n10566), .ZN(
        n14274) );
  AOI22_X1 U13041 ( .A1(n14571), .A2(n14277), .B1(n14274), .B2(n14573), .ZN(
        n10570) );
  OAI211_X1 U13042 ( .C1(n15109), .C2(n10572), .A(n10571), .B(n10570), .ZN(
        n10748) );
  NAND2_X1 U13043 ( .A1(n10748), .A2(n14552), .ZN(n10580) );
  OAI22_X1 U13044 ( .A1(n14552), .A2(n10574), .B1(n13977), .B2(n14578), .ZN(
        n10578) );
  NOR2_X1 U13045 ( .A1(n14519), .A2(n15161), .ZN(n14503) );
  INV_X1 U13046 ( .A(n14503), .ZN(n14371) );
  NOR2_X1 U13047 ( .A1(n10575), .A2(n13978), .ZN(n10576) );
  OR2_X1 U13048 ( .A1(n10805), .A2(n10576), .ZN(n10747) );
  NOR2_X1 U13049 ( .A1(n14371), .A2(n10747), .ZN(n10577) );
  AOI211_X1 U13050 ( .C1(n14737), .C2(n14071), .A(n10578), .B(n10577), .ZN(
        n10579) );
  OAI211_X1 U13051 ( .C1(n10581), .C2(n10936), .A(n10580), .B(n10579), .ZN(
        P1_U3287) );
  INV_X1 U13052 ( .A(n10582), .ZN(n10584) );
  AND2_X1 U13053 ( .A1(n11957), .A2(n13526), .ZN(n10588) );
  XNOR2_X1 U13054 ( .A(n10682), .B(n11961), .ZN(n10587) );
  NOR2_X1 U13055 ( .A1(n10587), .A2(n10588), .ZN(n10784) );
  AOI21_X1 U13056 ( .B1(n10588), .B2(n10587), .A(n10784), .ZN(n10589) );
  NAND2_X1 U13057 ( .A1(n10590), .A2(n10589), .ZN(n10786) );
  OAI21_X1 U13058 ( .B1(n10590), .B2(n10589), .A(n10786), .ZN(n10591) );
  NAND2_X1 U13059 ( .A1(n10591), .A2(n13454), .ZN(n10598) );
  NAND2_X1 U13060 ( .A1(n13475), .A2(n13527), .ZN(n10593) );
  OR2_X1 U13061 ( .A1(n13492), .A2(n10732), .ZN(n10592) );
  AND2_X1 U13062 ( .A1(n10593), .A2(n10592), .ZN(n10675) );
  OAI21_X1 U13063 ( .B1(n13476), .B2(n10675), .A(n10594), .ZN(n10596) );
  INV_X1 U13064 ( .A(n10682), .ZN(n15355) );
  NOR2_X1 U13065 ( .A1(n15355), .A2(n13461), .ZN(n10595) );
  AOI211_X1 U13066 ( .C1(n13467), .C2(n10681), .A(n10596), .B(n10595), .ZN(
        n10597) );
  NAND2_X1 U13067 ( .A1(n10598), .A2(n10597), .ZN(P2_U3193) );
  NAND2_X1 U13068 ( .A1(n10600), .A2(n10599), .ZN(n10602) );
  OR2_X1 U13069 ( .A1(n15347), .A2(n13527), .ZN(n10601) );
  NAND2_X1 U13070 ( .A1(n10682), .A2(n13526), .ZN(n10603) );
  INV_X1 U13071 ( .A(n10730), .ZN(n10604) );
  OR2_X1 U13072 ( .A1(n10605), .A2(n10604), .ZN(n10606) );
  NAND2_X1 U13073 ( .A1(n10726), .A2(n10606), .ZN(n15364) );
  AND2_X1 U13074 ( .A1(n15347), .A2(n10607), .ZN(n10608) );
  NAND2_X1 U13075 ( .A1(n10674), .A2(n10673), .ZN(n10612) );
  OR2_X1 U13076 ( .A1(n10682), .A2(n10610), .ZN(n10611) );
  NAND2_X1 U13077 ( .A1(n10612), .A2(n10611), .ZN(n10731) );
  XNOR2_X1 U13078 ( .A(n10731), .B(n10730), .ZN(n10616) );
  NAND2_X1 U13079 ( .A1(n13475), .A2(n13526), .ZN(n10614) );
  OR2_X1 U13080 ( .A1(n13492), .A2(n10892), .ZN(n10613) );
  AND2_X1 U13081 ( .A1(n10614), .A2(n10613), .ZN(n10790) );
  OR2_X1 U13082 ( .A1(n15364), .A2(n15342), .ZN(n10615) );
  OAI211_X1 U13083 ( .C1(n10616), .C2(n14819), .A(n10790), .B(n10615), .ZN(
        n15366) );
  NAND2_X1 U13084 ( .A1(n15366), .A2(n13748), .ZN(n10622) );
  AOI21_X1 U13085 ( .B1(n10679), .B2(n15361), .A(n13728), .ZN(n10617) );
  OR2_X2 U13086 ( .A1(n10679), .A2(n15361), .ZN(n10741) );
  NAND2_X1 U13087 ( .A1(n10617), .A2(n10741), .ZN(n15363) );
  INV_X1 U13088 ( .A(n15363), .ZN(n10620) );
  INV_X1 U13089 ( .A(n15361), .ZN(n10796) );
  AOI22_X1 U13090 ( .A1(n15292), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n10793), 
        .B2(n15279), .ZN(n10618) );
  OAI21_X1 U13091 ( .B1(n10796), .B2(n15282), .A(n10618), .ZN(n10619) );
  AOI21_X1 U13092 ( .B1(n10620), .B2(n15285), .A(n10619), .ZN(n10621) );
  OAI211_X1 U13093 ( .C1(n15364), .C2(n11625), .A(n10622), .B(n10621), .ZN(
        P2_U3256) );
  OAI222_X1 U13094 ( .A1(P2_U3088), .A2(n13587), .B1(n13854), .B2(n10624), 
        .C1(n10623), .C2(n13852), .ZN(P2_U3308) );
  NAND2_X1 U13095 ( .A1(n10632), .A2(n10667), .ZN(n10625) );
  NAND2_X1 U13096 ( .A1(n15119), .A2(n10625), .ZN(n15162) );
  XNOR2_X1 U13097 ( .A(n6932), .B(n15162), .ZN(n10627) );
  MUX2_X1 U13098 ( .A(n14222), .B(n10627), .S(n10626), .Z(n10628) );
  AOI222_X1 U13099 ( .A1(n14971), .A2(n10628), .B1(n14280), .B2(n14573), .C1(
        n9935), .C2(n14571), .ZN(n15163) );
  INV_X1 U13100 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n14283) );
  OAI22_X1 U13101 ( .A1(n14552), .A2(n10629), .B1(n14283), .B2(n14578), .ZN(
        n10631) );
  NOR2_X1 U13102 ( .A1(n14371), .A2(n15162), .ZN(n10630) );
  AOI211_X1 U13103 ( .C1(n14737), .C2(n10632), .A(n10631), .B(n10630), .ZN(
        n10637) );
  INV_X1 U13104 ( .A(n10633), .ZN(n10634) );
  XNOR2_X1 U13105 ( .A(n14222), .B(n10635), .ZN(n15166) );
  NAND2_X1 U13106 ( .A1(n14516), .A2(n15166), .ZN(n10636) );
  OAI211_X1 U13107 ( .C1(n15129), .C2(n15163), .A(n10637), .B(n10636), .ZN(
        P1_U3292) );
  NOR2_X1 U13108 ( .A1(n15116), .A2(n11060), .ZN(n10640) );
  INV_X1 U13109 ( .A(n11069), .ZN(n10638) );
  OAI22_X1 U13110 ( .A1(n14552), .A2(n9736), .B1(n10638), .B2(n14578), .ZN(
        n10639) );
  AOI211_X1 U13111 ( .C1(n10641), .C2(n15125), .A(n10640), .B(n10639), .ZN(
        n10644) );
  NAND2_X1 U13112 ( .A1(n10642), .A2(n14516), .ZN(n10643) );
  OAI211_X1 U13113 ( .C1(n10645), .C2(n15129), .A(n10644), .B(n10643), .ZN(
        P1_U3288) );
  XNOR2_X1 U13114 ( .A(n10646), .B(n14221), .ZN(n10648) );
  AOI21_X1 U13115 ( .B1(n10648), .B2(n14971), .A(n10647), .ZN(n15178) );
  OAI211_X1 U13116 ( .C1(n15122), .C2(n15179), .A(n15120), .B(n10649), .ZN(
        n15177) );
  OAI22_X1 U13117 ( .A1(n14519), .A2(n15177), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14578), .ZN(n10651) );
  NOR2_X1 U13118 ( .A1(n15116), .A2(n15179), .ZN(n10650) );
  AOI211_X1 U13119 ( .C1(n15129), .C2(P1_REG2_REG_3__SCAN_IN), .A(n10651), .B(
        n10650), .ZN(n10654) );
  XNOR2_X1 U13120 ( .A(n10652), .B(n14221), .ZN(n15176) );
  INV_X1 U13121 ( .A(n15176), .ZN(n15182) );
  NAND2_X1 U13122 ( .A1(n15182), .A2(n14516), .ZN(n10653) );
  OAI211_X1 U13123 ( .C1(n15129), .C2(n15178), .A(n10654), .B(n10653), .ZN(
        P1_U3290) );
  INV_X1 U13124 ( .A(n10970), .ZN(n10663) );
  NAND2_X1 U13125 ( .A1(n10655), .A2(n10963), .ZN(n10831) );
  AND2_X1 U13126 ( .A1(n10834), .A2(n10831), .ZN(n10657) );
  XNOR2_X1 U13127 ( .A(n12416), .B(n10660), .ZN(n10830) );
  XNOR2_X1 U13128 ( .A(n10830), .B(n12547), .ZN(n10656) );
  NAND2_X1 U13129 ( .A1(n10657), .A2(n10656), .ZN(n10775) );
  OAI211_X1 U13130 ( .C1(n10657), .C2(n10656), .A(n10775), .B(n12522), .ZN(
        n10662) );
  OAI22_X1 U13131 ( .A1(n10963), .A2(n12527), .B1(n12526), .B2(n12431), .ZN(
        n10658) );
  AOI211_X1 U13132 ( .C1(n10660), .C2(n12517), .A(n10659), .B(n10658), .ZN(
        n10661) );
  OAI211_X1 U13133 ( .C1(n10663), .C2(n11236), .A(n10662), .B(n10661), .ZN(
        P3_U3179) );
  NAND2_X1 U13134 ( .A1(n14552), .A2(n14971), .ZN(n14483) );
  INV_X1 U13135 ( .A(n14483), .ZN(n14505) );
  NOR2_X1 U13136 ( .A1(n14505), .A2(n14516), .ZN(n10670) );
  INV_X1 U13137 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10664) );
  OAI22_X1 U13138 ( .A1(n15129), .A2(n10665), .B1(n10664), .B2(n14578), .ZN(
        n10666) );
  AOI21_X1 U13139 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n15129), .A(n10666), .ZN(
        n10669) );
  OAI21_X1 U13140 ( .B1(n14737), .B2(n14503), .A(n10667), .ZN(n10668) );
  OAI211_X1 U13141 ( .C1(n10670), .C2(n14219), .A(n10669), .B(n10668), .ZN(
        P1_U3293) );
  INV_X1 U13142 ( .A(n10673), .ZN(n10671) );
  XNOR2_X1 U13143 ( .A(n10672), .B(n10671), .ZN(n15359) );
  INV_X1 U13144 ( .A(n15359), .ZN(n10687) );
  XNOR2_X1 U13145 ( .A(n10674), .B(n10673), .ZN(n10676) );
  OAI21_X1 U13146 ( .B1(n10676), .B2(n14819), .A(n10675), .ZN(n10677) );
  AOI21_X1 U13147 ( .B1(n11622), .B2(n15359), .A(n10677), .ZN(n15356) );
  MUX2_X1 U13148 ( .A(n10678), .B(n15356), .S(n13748), .Z(n10686) );
  OAI211_X1 U13149 ( .C1(n10680), .C2(n15355), .A(n14852), .B(n10679), .ZN(
        n15354) );
  INV_X1 U13150 ( .A(n15285), .ZN(n13685) );
  AOI22_X1 U13151 ( .A1(n14844), .A2(n10682), .B1(n10681), .B2(n15279), .ZN(
        n10683) );
  OAI21_X1 U13152 ( .B1(n15354), .B2(n13685), .A(n10683), .ZN(n10684) );
  INV_X1 U13153 ( .A(n10684), .ZN(n10685) );
  OAI211_X1 U13154 ( .C1(n10687), .C2(n11625), .A(n10686), .B(n10685), .ZN(
        P2_U3257) );
  INV_X1 U13155 ( .A(SI_23_), .ZN(n10690) );
  NAND2_X1 U13156 ( .A1(n10688), .A2(n13381), .ZN(n10689) );
  OAI211_X1 U13157 ( .C1(n10690), .C2(n14721), .A(n10689), .B(n12192), .ZN(
        P3_U3272) );
  INV_X1 U13158 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n10691) );
  OAI22_X1 U13159 ( .A1(n10694), .A2(n10693), .B1(n10692), .B2(n10691), .ZN(
        n10695) );
  NAND2_X1 U13160 ( .A1(n15253), .A2(n10695), .ZN(n10696) );
  XOR2_X1 U13161 ( .A(n15253), .B(n10695), .Z(n15256) );
  NAND2_X1 U13162 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n15256), .ZN(n15255) );
  NAND2_X1 U13163 ( .A1(n10696), .A2(n15255), .ZN(n10700) );
  NOR2_X1 U13164 ( .A1(n11182), .A2(n10697), .ZN(n10698) );
  AOI21_X1 U13165 ( .B1(n10697), .B2(n11182), .A(n10698), .ZN(n10699) );
  NAND2_X1 U13166 ( .A1(n10699), .A2(n10700), .ZN(n11176) );
  OAI211_X1 U13167 ( .C1(n10700), .C2(n10699), .A(n15271), .B(n11176), .ZN(
        n10714) );
  NAND2_X1 U13168 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n13433)
         );
  NOR2_X1 U13169 ( .A1(n10702), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n10701) );
  AOI21_X1 U13170 ( .B1(n10702), .B2(P2_REG1_REG_16__SCAN_IN), .A(n10701), 
        .ZN(n10710) );
  AOI21_X1 U13171 ( .B1(n10704), .B2(P2_REG1_REG_14__SCAN_IN), .A(n10703), 
        .ZN(n10708) );
  INV_X1 U13172 ( .A(n10708), .ZN(n10705) );
  XNOR2_X1 U13173 ( .A(n10705), .B(n15253), .ZN(n15257) );
  INV_X1 U13174 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n10706) );
  OAI22_X1 U13175 ( .A1(n10708), .A2(n10707), .B1(n15257), .B2(n10706), .ZN(
        n10709) );
  NAND2_X1 U13176 ( .A1(n10710), .A2(n10709), .ZN(n11181) );
  OAI211_X1 U13177 ( .C1(n10710), .C2(n10709), .A(n15264), .B(n11181), .ZN(
        n10711) );
  NAND2_X1 U13178 ( .A1(n13433), .A2(n10711), .ZN(n10712) );
  AOI21_X1 U13179 ( .B1(n15270), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n10712), 
        .ZN(n10713) );
  OAI211_X1 U13180 ( .C1(n15278), .C2(n11182), .A(n10714), .B(n10713), .ZN(
        P2_U3230) );
  INV_X1 U13181 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10720) );
  AOI22_X1 U13182 ( .A1(n10715), .A2(n15125), .B1(n14737), .B2(n14053), .ZN(
        n10719) );
  AOI22_X1 U13183 ( .A1(n14552), .A2(n10717), .B1(n10716), .B2(n15114), .ZN(
        n10718) );
  OAI211_X1 U13184 ( .C1(n10720), .C2(n14552), .A(n10719), .B(n10718), .ZN(
        n10721) );
  AOI21_X1 U13185 ( .B1(n14505), .B2(n10722), .A(n10721), .ZN(n10723) );
  OAI21_X1 U13186 ( .B1(n14584), .B2(n10724), .A(n10723), .ZN(P1_U3289) );
  NAND2_X1 U13187 ( .A1(n15361), .A2(n13525), .ZN(n10725) );
  INV_X1 U13188 ( .A(n10756), .ZN(n10727) );
  OR2_X1 U13189 ( .A1(n10728), .A2(n10727), .ZN(n10729) );
  NAND2_X1 U13190 ( .A1(n10765), .A2(n10729), .ZN(n15373) );
  NAND2_X1 U13191 ( .A1(n10731), .A2(n10730), .ZN(n10734) );
  OR2_X1 U13192 ( .A1(n15361), .A2(n10732), .ZN(n10733) );
  XNOR2_X1 U13193 ( .A(n10756), .B(n10757), .ZN(n10738) );
  OR2_X1 U13194 ( .A1(n15373), .A2(n15342), .ZN(n10737) );
  NAND2_X1 U13195 ( .A1(n13475), .A2(n13525), .ZN(n10736) );
  OR2_X1 U13196 ( .A1(n13492), .A2(n10986), .ZN(n10735) );
  AND2_X1 U13197 ( .A1(n10736), .A2(n10735), .ZN(n10895) );
  OAI211_X1 U13198 ( .C1(n10738), .C2(n14819), .A(n10737), .B(n10895), .ZN(
        n15375) );
  NAND2_X1 U13199 ( .A1(n15375), .A2(n13748), .ZN(n10746) );
  INV_X1 U13200 ( .A(n10893), .ZN(n10739) );
  OAI22_X1 U13201 ( .A1(n13748), .A2(n9512), .B1(n10739), .B2(n14827), .ZN(
        n10744) );
  NAND2_X1 U13202 ( .A1(n10741), .A2(n15369), .ZN(n10740) );
  NAND2_X1 U13203 ( .A1(n10740), .A2(n14852), .ZN(n10742) );
  OR2_X1 U13204 ( .A1(n10742), .A2(n10767), .ZN(n15371) );
  NOR2_X1 U13205 ( .A1(n15371), .A2(n13685), .ZN(n10743) );
  AOI211_X1 U13206 ( .C1(n14844), .C2(n15369), .A(n10744), .B(n10743), .ZN(
        n10745) );
  OAI211_X1 U13207 ( .C1(n15373), .C2(n11625), .A(n10746), .B(n10745), .ZN(
        P2_U3255) );
  INV_X1 U13208 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10752) );
  INV_X1 U13209 ( .A(n15175), .ZN(n15173) );
  OAI22_X1 U13210 ( .A1(n10747), .A2(n15161), .B1(n13978), .B2(n15187), .ZN(
        n10749) );
  AOI211_X1 U13211 ( .C1(n15173), .C2(n10750), .A(n10749), .B(n10748), .ZN(
        n10753) );
  OR2_X1 U13212 ( .A1(n10753), .A2(n15200), .ZN(n10751) );
  OAI21_X1 U13213 ( .B1(n15202), .B2(n10752), .A(n10751), .ZN(P1_U3534) );
  INV_X1 U13214 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10755) );
  OR2_X1 U13215 ( .A1(n10753), .A2(n15192), .ZN(n10754) );
  OAI21_X1 U13216 ( .B1(n15194), .B2(n10755), .A(n10754), .ZN(P1_U3477) );
  INV_X1 U13217 ( .A(n11711), .ZN(n10828) );
  OAI222_X1 U13218 ( .A1(n11910), .A2(n10828), .B1(P1_U3086), .B2(n14020), 
        .C1(n13291), .C2(n14694), .ZN(P1_U3335) );
  OR2_X1 U13219 ( .A1(n15369), .A2(n10892), .ZN(n10758) );
  NAND2_X1 U13220 ( .A1(n10760), .A2(n14841), .ZN(n10763) );
  NAND2_X1 U13221 ( .A1(n13475), .A2(n13524), .ZN(n10762) );
  OR2_X1 U13222 ( .A1(n13492), .A2(n10989), .ZN(n10761) );
  AND2_X1 U13223 ( .A1(n10762), .A2(n10761), .ZN(n11166) );
  NAND2_X1 U13224 ( .A1(n10763), .A2(n11166), .ZN(n15383) );
  INV_X1 U13225 ( .A(n15383), .ZN(n10773) );
  INV_X1 U13226 ( .A(n10988), .ZN(n10766) );
  XNOR2_X1 U13227 ( .A(n10996), .B(n10766), .ZN(n15378) );
  INV_X1 U13228 ( .A(n11170), .ZN(n15381) );
  OAI21_X1 U13229 ( .B1(n10767), .B2(n15381), .A(n14852), .ZN(n10768) );
  OR2_X1 U13230 ( .A1(n11013), .A2(n10768), .ZN(n15379) );
  AOI22_X1 U13231 ( .A1(n15292), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n11169), 
        .B2(n15279), .ZN(n10770) );
  NAND2_X1 U13232 ( .A1(n11170), .A2(n14844), .ZN(n10769) );
  OAI211_X1 U13233 ( .C1(n15379), .C2(n13685), .A(n10770), .B(n10769), .ZN(
        n10771) );
  AOI21_X1 U13234 ( .B1(n15378), .B2(n15288), .A(n10771), .ZN(n10772) );
  OAI21_X1 U13235 ( .B1(n10773), .B2(n15292), .A(n10772), .ZN(P2_U3254) );
  INV_X1 U13236 ( .A(n10830), .ZN(n10774) );
  NAND2_X1 U13237 ( .A1(n10774), .A2(n12547), .ZN(n10836) );
  NAND2_X1 U13238 ( .A1(n10775), .A2(n10836), .ZN(n12424) );
  XNOR2_X1 U13239 ( .A(n12022), .B(n6823), .ZN(n12423) );
  XNOR2_X1 U13240 ( .A(n12424), .B(n12423), .ZN(n10781) );
  OAI22_X1 U13241 ( .A1(n10947), .A2(n12527), .B1(n12526), .B2(n11142), .ZN(
        n10776) );
  AOI211_X1 U13242 ( .C1(n10778), .C2(n12517), .A(n10777), .B(n10776), .ZN(
        n10780) );
  NAND2_X1 U13243 ( .A1(n12530), .A2(n10951), .ZN(n10779) );
  OAI211_X1 U13244 ( .C1(n10781), .C2(n12520), .A(n10780), .B(n10779), .ZN(
        P3_U3153) );
  AND2_X1 U13245 ( .A1(n9669), .A2(n13525), .ZN(n10783) );
  XNOR2_X1 U13246 ( .A(n15361), .B(n11968), .ZN(n10782) );
  NOR2_X1 U13247 ( .A1(n10782), .A2(n10783), .ZN(n10889) );
  AOI21_X1 U13248 ( .B1(n10783), .B2(n10782), .A(n10889), .ZN(n10788) );
  INV_X1 U13249 ( .A(n10784), .ZN(n10785) );
  NAND2_X1 U13250 ( .A1(n10786), .A2(n10785), .ZN(n10787) );
  NAND2_X1 U13251 ( .A1(n10787), .A2(n10788), .ZN(n10891) );
  OAI21_X1 U13252 ( .B1(n10788), .B2(n10787), .A(n10891), .ZN(n10789) );
  NAND2_X1 U13253 ( .A1(n10789), .A2(n13454), .ZN(n10795) );
  NOR2_X1 U13254 ( .A1(n13476), .A2(n10790), .ZN(n10791) );
  AOI211_X1 U13255 ( .C1(n13467), .C2(n10793), .A(n10792), .B(n10791), .ZN(
        n10794) );
  OAI211_X1 U13256 ( .C1(n10796), .C2(n13461), .A(n10795), .B(n10794), .ZN(
        P2_U3203) );
  INV_X1 U13257 ( .A(n14276), .ZN(n11030) );
  NAND2_X1 U13258 ( .A1(n11030), .A2(n13978), .ZN(n10797) );
  NAND2_X1 U13259 ( .A1(n10798), .A2(n10797), .ZN(n10803) );
  NAND2_X1 U13260 ( .A1(n10799), .A2(n14017), .ZN(n10802) );
  AOI22_X1 U13261 ( .A1(n11700), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n11699), 
        .B2(n10800), .ZN(n10801) );
  NAND2_X1 U13262 ( .A1(n10802), .A2(n10801), .ZN(n14074) );
  XNOR2_X1 U13263 ( .A(n14274), .B(n14074), .ZN(n14227) );
  INV_X1 U13264 ( .A(n14227), .ZN(n10809) );
  NAND2_X1 U13265 ( .A1(n10803), .A2(n10809), .ZN(n10851) );
  OR2_X1 U13266 ( .A1(n10803), .A2(n10809), .ZN(n10804) );
  NAND2_X1 U13267 ( .A1(n10851), .A2(n10804), .ZN(n10942) );
  NAND2_X1 U13268 ( .A1(n10805), .A2(n14087), .ZN(n10859) );
  OAI211_X1 U13269 ( .C1(n10805), .C2(n14087), .A(n15120), .B(n10859), .ZN(
        n10938) );
  OAI21_X1 U13270 ( .B1(n14087), .B2(n15187), .A(n10938), .ZN(n10825) );
  NAND2_X1 U13271 ( .A1(n10942), .A2(n15183), .ZN(n10824) );
  NOR2_X1 U13272 ( .A1(n14276), .A2(n13978), .ZN(n10806) );
  NAND2_X1 U13273 ( .A1(n14276), .A2(n13978), .ZN(n10808) );
  XNOR2_X1 U13274 ( .A(n10870), .B(n10809), .ZN(n10822) );
  NAND2_X1 U13275 ( .A1(n14276), .A2(n14571), .ZN(n10820) );
  INV_X1 U13276 ( .A(n10812), .ZN(n10810) );
  AOI21_X1 U13277 ( .B1(n10810), .B2(P1_REG3_REG_7__SCAN_IN), .A(
        P1_REG3_REG_8__SCAN_IN), .ZN(n10813) );
  NAND2_X1 U13278 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n10811) );
  NOR2_X1 U13279 ( .A1(n10812), .A2(n10811), .ZN(n10860) );
  OR2_X1 U13280 ( .A1(n10813), .A2(n10860), .ZN(n11209) );
  INV_X1 U13281 ( .A(n11209), .ZN(n10814) );
  NAND2_X1 U13282 ( .A1(n11751), .A2(n10814), .ZN(n10818) );
  NAND2_X1 U13283 ( .A1(n11774), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n10817) );
  NAND2_X1 U13284 ( .A1(n11715), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n10816) );
  NAND2_X1 U13285 ( .A1(n14011), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10815) );
  NAND4_X1 U13286 ( .A1(n10818), .A2(n10817), .A3(n10816), .A4(n10815), .ZN(
        n14273) );
  NAND2_X1 U13287 ( .A1(n14273), .A2(n14573), .ZN(n10819) );
  NAND2_X1 U13288 ( .A1(n10820), .A2(n10819), .ZN(n10821) );
  AOI21_X1 U13289 ( .B1(n10822), .B2(n14971), .A(n10821), .ZN(n10823) );
  NAND2_X1 U13290 ( .A1(n10824), .A2(n10823), .ZN(n10939) );
  AOI211_X1 U13291 ( .C1(n15173), .C2(n10942), .A(n10825), .B(n10939), .ZN(
        n10902) );
  NAND2_X1 U13292 ( .A1(n15200), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10826) );
  OAI21_X1 U13293 ( .B1(n10902), .B2(n15200), .A(n10826), .ZN(P1_U3535) );
  OAI222_X1 U13294 ( .A1(n13852), .A2(n10829), .B1(n13854), .B2(n10828), .C1(
        n10827), .C2(P2_U3088), .ZN(P2_U3307) );
  XNOR2_X1 U13295 ( .A(n12416), .B(n11310), .ZN(n10906) );
  XNOR2_X1 U13296 ( .A(n10906), .B(n12544), .ZN(n10844) );
  XNOR2_X1 U13297 ( .A(n12416), .B(n11220), .ZN(n10838) );
  XNOR2_X1 U13298 ( .A(n10838), .B(n11142), .ZN(n10835) );
  NAND2_X1 U13299 ( .A1(n10830), .A2(n10947), .ZN(n10832) );
  OAI21_X1 U13300 ( .B1(n12425), .B2(n10836), .A(n12423), .ZN(n10840) );
  INV_X1 U13301 ( .A(n12423), .ZN(n10837) );
  OAI21_X1 U13302 ( .B1(n12425), .B2(n12431), .A(n10837), .ZN(n10839) );
  AOI22_X1 U13303 ( .A1(n10840), .A2(n10839), .B1(n10838), .B2(n12545), .ZN(
        n10841) );
  INV_X1 U13304 ( .A(n10910), .ZN(n10842) );
  AOI21_X1 U13305 ( .B1(n10844), .B2(n10843), .A(n10842), .ZN(n10849) );
  NOR2_X1 U13306 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13326), .ZN(n10924) );
  OAI22_X1 U13307 ( .A1(n11142), .A2(n12527), .B1(n12526), .B2(n11443), .ZN(
        n10845) );
  AOI211_X1 U13308 ( .C1(n10846), .C2(n12517), .A(n10924), .B(n10845), .ZN(
        n10848) );
  NAND2_X1 U13309 ( .A1(n12530), .A2(n11147), .ZN(n10847) );
  OAI211_X1 U13310 ( .C1(n10849), .C2(n12520), .A(n10848), .B(n10847), .ZN(
        P3_U3171) );
  INV_X1 U13311 ( .A(n14274), .ZN(n14088) );
  NAND2_X1 U13312 ( .A1(n14088), .A2(n14087), .ZN(n10850) );
  NAND2_X1 U13313 ( .A1(n10852), .A2(n14017), .ZN(n10855) );
  AOI22_X1 U13314 ( .A1(n11700), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n11699), 
        .B2(n10853), .ZN(n10854) );
  NAND2_X1 U13315 ( .A1(n10855), .A2(n10854), .ZN(n14075) );
  NOR2_X1 U13316 ( .A1(n14075), .A2(n14273), .ZN(n14076) );
  INV_X1 U13317 ( .A(n14076), .ZN(n11102) );
  NAND2_X1 U13318 ( .A1(n14075), .A2(n14273), .ZN(n10856) );
  NAND2_X1 U13319 ( .A1(n11102), .A2(n10856), .ZN(n14226) );
  OAI21_X1 U13320 ( .B1(n10857), .B2(n10871), .A(n11103), .ZN(n10858) );
  INV_X1 U13321 ( .A(n10858), .ZN(n10885) );
  AOI21_X1 U13322 ( .B1(n14075), .B2(n10859), .A(n7202), .ZN(n10880) );
  INV_X1 U13323 ( .A(n14075), .ZN(n11083) );
  NOR2_X1 U13324 ( .A1(n11083), .A2(n15187), .ZN(n10868) );
  NAND2_X1 U13325 ( .A1(n14274), .A2(n14571), .ZN(n10867) );
  NAND2_X1 U13326 ( .A1(n10860), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n11091) );
  OR2_X1 U13327 ( .A1(n10860), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n10861) );
  AND2_X1 U13328 ( .A1(n11091), .A2(n10861), .ZN(n11364) );
  NAND2_X1 U13329 ( .A1(n11751), .A2(n11364), .ZN(n10865) );
  NAND2_X1 U13330 ( .A1(n11774), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n10864) );
  NAND2_X1 U13331 ( .A1(n14012), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n10863) );
  NAND2_X1 U13332 ( .A1(n14011), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10862) );
  NAND4_X1 U13333 ( .A1(n10865), .A2(n10864), .A3(n10863), .A4(n10862), .ZN(
        n14272) );
  NAND2_X1 U13334 ( .A1(n14272), .A2(n14573), .ZN(n10866) );
  NAND2_X1 U13335 ( .A1(n10867), .A2(n10866), .ZN(n11206) );
  AOI211_X1 U13336 ( .C1(n10880), .C2(n15120), .A(n10868), .B(n11206), .ZN(
        n10874) );
  NOR2_X1 U13337 ( .A1(n14088), .A2(n14074), .ZN(n10869) );
  INV_X1 U13338 ( .A(n11086), .ZN(n10882) );
  NAND2_X1 U13339 ( .A1(n10872), .A2(n10871), .ZN(n10881) );
  NAND3_X1 U13340 ( .A1(n10882), .A2(n14971), .A3(n10881), .ZN(n10873) );
  OAI211_X1 U13341 ( .C1(n10885), .C2(n14670), .A(n10874), .B(n10873), .ZN(
        n10886) );
  NAND2_X1 U13342 ( .A1(n10886), .A2(n15202), .ZN(n10875) );
  OAI21_X1 U13343 ( .B1(n15202), .B2(n9729), .A(n10875), .ZN(P1_U3536) );
  INV_X1 U13344 ( .A(n11206), .ZN(n10876) );
  OAI22_X1 U13345 ( .A1(n15129), .A2(n10876), .B1(n11209), .B2(n14578), .ZN(
        n10877) );
  AOI21_X1 U13346 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n15129), .A(n10877), .ZN(
        n10878) );
  OAI21_X1 U13347 ( .B1(n11083), .B2(n15116), .A(n10878), .ZN(n10879) );
  AOI21_X1 U13348 ( .B1(n10880), .B2(n14503), .A(n10879), .ZN(n10884) );
  NAND3_X1 U13349 ( .A1(n10882), .A2(n14505), .A3(n10881), .ZN(n10883) );
  OAI211_X1 U13350 ( .C1(n10885), .C2(n14584), .A(n10884), .B(n10883), .ZN(
        P1_U3285) );
  INV_X1 U13351 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10888) );
  NAND2_X1 U13352 ( .A1(n10886), .A2(n15194), .ZN(n10887) );
  OAI21_X1 U13353 ( .B1(n15194), .B2(n10888), .A(n10887), .ZN(P1_U3483) );
  INV_X1 U13354 ( .A(n10889), .ZN(n10890) );
  XNOR2_X1 U13355 ( .A(n15369), .B(n11961), .ZN(n11158) );
  NOR2_X1 U13356 ( .A1(n11966), .A2(n10892), .ZN(n11159) );
  XNOR2_X1 U13357 ( .A(n11158), .B(n11159), .ZN(n11160) );
  XNOR2_X1 U13358 ( .A(n11161), .B(n11160), .ZN(n10898) );
  NAND2_X1 U13359 ( .A1(n13467), .A2(n10893), .ZN(n10894) );
  NAND2_X1 U13360 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n15217)
         );
  OAI211_X1 U13361 ( .C1(n10895), .C2(n13476), .A(n10894), .B(n15217), .ZN(
        n10896) );
  AOI21_X1 U13362 ( .B1(n15369), .B2(n13501), .A(n10896), .ZN(n10897) );
  OAI21_X1 U13363 ( .B1(n10898), .B2(n13503), .A(n10897), .ZN(P2_U3189) );
  INV_X1 U13364 ( .A(n11723), .ZN(n10901) );
  OAI222_X1 U13365 ( .A1(n13852), .A2(n10900), .B1(n13854), .B2(n10901), .C1(
        P2_U3088), .C2(n10899), .ZN(P2_U3306) );
  OAI222_X1 U13366 ( .A1(n14694), .A2(n11724), .B1(n11910), .B2(n10901), .C1(
        n14195), .C2(P1_U3086), .ZN(P1_U3334) );
  INV_X1 U13367 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10904) );
  OR2_X1 U13368 ( .A1(n10902), .A2(n15192), .ZN(n10903) );
  OAI21_X1 U13369 ( .B1(n15194), .B2(n10904), .A(n10903), .ZN(P1_U3480) );
  INV_X1 U13370 ( .A(n10905), .ZN(n11333) );
  INV_X1 U13371 ( .A(n10906), .ZN(n10907) );
  INV_X1 U13372 ( .A(n12544), .ZN(n12430) );
  NAND2_X1 U13373 ( .A1(n10907), .A2(n12430), .ZN(n10908) );
  AND2_X1 U13374 ( .A1(n10910), .A2(n10908), .ZN(n10912) );
  XNOR2_X1 U13375 ( .A(n12390), .B(n11336), .ZN(n11223) );
  XNOR2_X1 U13376 ( .A(n11223), .B(n12543), .ZN(n10911) );
  AND2_X1 U13377 ( .A1(n10911), .A2(n10908), .ZN(n10909) );
  OAI211_X1 U13378 ( .C1(n10912), .C2(n10911), .A(n12522), .B(n11226), .ZN(
        n10915) );
  AND2_X1 U13379 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n15418) );
  OAI22_X1 U13380 ( .A1(n12430), .A2(n12527), .B1(n12526), .B2(n14777), .ZN(
        n10913) );
  AOI211_X1 U13381 ( .C1(n11336), .C2(n12517), .A(n15418), .B(n10913), .ZN(
        n10914) );
  OAI211_X1 U13382 ( .C1(n11333), .C2(n11236), .A(n10915), .B(n10914), .ZN(
        P3_U3157) );
  INV_X1 U13383 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n10920) );
  NOR2_X1 U13384 ( .A1(n10920), .A2(n10917), .ZN(n11264) );
  AOI21_X1 U13385 ( .B1(n10920), .B2(n10917), .A(n11264), .ZN(n10935) );
  INV_X1 U13386 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11301) );
  MUX2_X1 U13387 ( .A(n10920), .B(n11301), .S(n6642), .Z(n10921) );
  NAND2_X1 U13388 ( .A1(n10921), .A2(n7439), .ZN(n11272) );
  INV_X1 U13389 ( .A(n10921), .ZN(n10922) );
  NAND2_X1 U13390 ( .A1(n10922), .A2(n10929), .ZN(n11274) );
  NAND2_X1 U13391 ( .A1(n11272), .A2(n11274), .ZN(n10923) );
  XNOR2_X1 U13392 ( .A(n11275), .B(n10923), .ZN(n10926) );
  AOI21_X1 U13393 ( .B1(n15405), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n10924), .ZN(
        n10925) );
  OAI21_X1 U13394 ( .B1(n15434), .B2(n10926), .A(n10925), .ZN(n10933) );
  AOI21_X1 U13395 ( .B1(n11301), .B2(n10930), .A(n11256), .ZN(n10931) );
  NOR2_X1 U13396 ( .A1(n10931), .A2(n15425), .ZN(n10932) );
  AOI211_X1 U13397 ( .C1(n15430), .C2(n7439), .A(n10933), .B(n10932), .ZN(
        n10934) );
  OAI21_X1 U13398 ( .B1(n10935), .B2(n15438), .A(n10934), .ZN(P3_U3191) );
  INV_X1 U13399 ( .A(n10936), .ZN(n15126) );
  AOI22_X1 U13400 ( .A1(n14737), .A2(n14074), .B1(n11028), .B2(n15114), .ZN(
        n10937) );
  OAI21_X1 U13401 ( .B1(n14519), .B2(n10938), .A(n10937), .ZN(n10941) );
  MUX2_X1 U13402 ( .A(n10939), .B(P1_REG2_REG_7__SCAN_IN), .S(n15129), .Z(
        n10940) );
  AOI211_X1 U13403 ( .C1(n15126), .C2(n10942), .A(n10941), .B(n10940), .ZN(
        n10943) );
  INV_X1 U13404 ( .A(n10943), .ZN(P1_U3286) );
  XNOR2_X1 U13405 ( .A(n10944), .B(n12022), .ZN(n15510) );
  OAI211_X1 U13406 ( .C1(n10946), .C2(n12022), .A(n10945), .B(n15466), .ZN(
        n10950) );
  OAI22_X1 U13407 ( .A1(n10947), .A2(n15450), .B1(n11142), .B2(n15448), .ZN(
        n10948) );
  INV_X1 U13408 ( .A(n10948), .ZN(n10949) );
  OAI211_X1 U13409 ( .C1(n15510), .C2(n15470), .A(n10950), .B(n10949), .ZN(
        n15512) );
  AOI21_X1 U13410 ( .B1(n15473), .B2(n10951), .A(n15512), .ZN(n10956) );
  INV_X1 U13411 ( .A(n15510), .ZN(n10954) );
  OAI22_X1 U13412 ( .A1(n12867), .A2(n15509), .B1(n10952), .B2(n15477), .ZN(
        n10953) );
  AOI21_X1 U13413 ( .B1(n10954), .B2(n15474), .A(n10953), .ZN(n10955) );
  OAI21_X1 U13414 ( .B1(n10956), .B2(n12871), .A(n10955), .ZN(P3_U3226) );
  OR2_X1 U13415 ( .A1(n10957), .A2(n12018), .ZN(n10958) );
  NAND2_X1 U13416 ( .A1(n10959), .A2(n10958), .ZN(n15507) );
  INV_X1 U13417 ( .A(n15507), .ZN(n10973) );
  NAND2_X1 U13418 ( .A1(n10960), .A2(n12018), .ZN(n10961) );
  NAND3_X1 U13419 ( .A1(n10962), .A2(n15466), .A3(n10961), .ZN(n10967) );
  OAI22_X1 U13420 ( .A1(n10963), .A2(n15450), .B1(n12431), .B2(n15448), .ZN(
        n10964) );
  INV_X1 U13421 ( .A(n10964), .ZN(n10966) );
  NAND2_X1 U13422 ( .A1(n15507), .A2(n15453), .ZN(n10965) );
  NAND3_X1 U13423 ( .A1(n10967), .A2(n10966), .A3(n10965), .ZN(n15505) );
  MUX2_X1 U13424 ( .A(n15505), .B(P3_REG2_REG_6__SCAN_IN), .S(n12871), .Z(
        n10968) );
  INV_X1 U13425 ( .A(n10968), .ZN(n10972) );
  NOR2_X1 U13426 ( .A1(n10969), .A2(n15521), .ZN(n15506) );
  AOI22_X1 U13427 ( .A1(n14782), .A2(n15506), .B1(n15473), .B2(n10970), .ZN(
        n10971) );
  OAI211_X1 U13428 ( .C1(n10973), .C2(n12752), .A(n10972), .B(n10971), .ZN(
        P3_U3227) );
  INV_X1 U13429 ( .A(n12025), .ZN(n12067) );
  XNOR2_X1 U13430 ( .A(n10974), .B(n12067), .ZN(n15500) );
  NAND2_X1 U13431 ( .A1(n10975), .A2(n12025), .ZN(n10976) );
  NAND2_X1 U13432 ( .A1(n10977), .A2(n10976), .ZN(n10978) );
  NAND2_X1 U13433 ( .A1(n10978), .A2(n15466), .ZN(n10980) );
  INV_X1 U13434 ( .A(n15450), .ZN(n15464) );
  AOI22_X1 U13435 ( .A1(n12547), .A2(n15461), .B1(n15464), .B2(n12548), .ZN(
        n10979) );
  OAI211_X1 U13436 ( .C1(n15500), .C2(n15470), .A(n10980), .B(n10979), .ZN(
        n15501) );
  MUX2_X1 U13437 ( .A(n15501), .B(P3_REG2_REG_5__SCAN_IN), .S(n12871), .Z(
        n10981) );
  INV_X1 U13438 ( .A(n10981), .ZN(n10985) );
  NOR2_X1 U13439 ( .A1(n10982), .A2(n15521), .ZN(n15502) );
  AOI22_X1 U13440 ( .A1(n14782), .A2(n15502), .B1(n15473), .B2(n10983), .ZN(
        n10984) );
  OAI211_X1 U13441 ( .C1(n15500), .C2(n12752), .A(n10985), .B(n10984), .ZN(
        P3_U3228) );
  NAND2_X1 U13442 ( .A1(n11170), .A2(n10986), .ZN(n10987) );
  OR2_X1 U13443 ( .A1(n11238), .A2(n10989), .ZN(n10990) );
  XNOR2_X1 U13444 ( .A(n11576), .B(n11574), .ZN(n10991) );
  NAND2_X1 U13445 ( .A1(n10991), .A2(n14841), .ZN(n10994) );
  NAND2_X1 U13446 ( .A1(n13475), .A2(n13522), .ZN(n10993) );
  OR2_X1 U13447 ( .A1(n11579), .A2(n13492), .ZN(n10992) );
  AND2_X1 U13448 ( .A1(n10993), .A2(n10992), .ZN(n11292) );
  NAND2_X1 U13449 ( .A1(n10994), .A2(n11292), .ZN(n14889) );
  INV_X1 U13450 ( .A(n14889), .ZN(n11003) );
  OR2_X1 U13451 ( .A1(n11170), .A2(n13523), .ZN(n10995) );
  INV_X1 U13452 ( .A(n11008), .ZN(n11007) );
  OR2_X1 U13453 ( .A1(n11238), .A2(n13522), .ZN(n10997) );
  XNOR2_X1 U13454 ( .A(n11566), .B(n11574), .ZN(n14884) );
  INV_X1 U13455 ( .A(n11238), .ZN(n11250) );
  NAND2_X1 U13456 ( .A1(n11013), .A2(n11250), .ZN(n11014) );
  AOI21_X1 U13457 ( .B1(n11014), .B2(n14885), .A(n13728), .ZN(n10998) );
  OR2_X2 U13458 ( .A1(n11014), .A2(n14885), .ZN(n14850) );
  NAND2_X1 U13459 ( .A1(n10998), .A2(n14850), .ZN(n14887) );
  AOI22_X1 U13460 ( .A1(n15292), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n11294), 
        .B2(n15279), .ZN(n11000) );
  NAND2_X1 U13461 ( .A1(n14885), .A2(n14844), .ZN(n10999) );
  OAI211_X1 U13462 ( .C1(n14887), .C2(n13685), .A(n11000), .B(n10999), .ZN(
        n11001) );
  AOI21_X1 U13463 ( .B1(n14884), .B2(n15288), .A(n11001), .ZN(n11002) );
  OAI21_X1 U13464 ( .B1(n11003), .B2(n15292), .A(n11002), .ZN(P2_U3252) );
  INV_X1 U13465 ( .A(n11004), .ZN(n11005) );
  AOI21_X1 U13466 ( .B1(n11007), .B2(n11006), .A(n11005), .ZN(n11112) );
  AOI21_X1 U13467 ( .B1(n11009), .B2(n11008), .A(n14819), .ZN(n11012) );
  AOI22_X1 U13468 ( .A1(n13474), .A2(n11567), .B1(n13475), .B2(n13523), .ZN(
        n11245) );
  INV_X1 U13469 ( .A(n11245), .ZN(n11010) );
  AOI21_X1 U13470 ( .B1(n11012), .B2(n11011), .A(n11010), .ZN(n11117) );
  INV_X1 U13471 ( .A(n11013), .ZN(n11016) );
  INV_X1 U13472 ( .A(n11014), .ZN(n11015) );
  AOI211_X1 U13473 ( .C1(n11238), .C2(n11016), .A(n13728), .B(n11015), .ZN(
        n11115) );
  AOI21_X1 U13474 ( .B1(n15368), .B2(n11238), .A(n11115), .ZN(n11017) );
  OAI211_X1 U13475 ( .C1(n11112), .C2(n15350), .A(n11117), .B(n11017), .ZN(
        n11022) );
  NAND2_X1 U13476 ( .A1(n11022), .A2(n15401), .ZN(n11018) );
  OAI21_X1 U13477 ( .B1(n15401), .B2(n13312), .A(n11018), .ZN(P2_U3511) );
  INV_X1 U13478 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n11024) );
  NAND2_X1 U13479 ( .A1(n11022), .A2(n15387), .ZN(n11023) );
  OAI21_X1 U13480 ( .B1(n15387), .B2(n11024), .A(n11023), .ZN(P2_U3466) );
  INV_X1 U13481 ( .A(n11025), .ZN(n11026) );
  OAI222_X1 U13482 ( .A1(n13852), .A2(n11027), .B1(n13854), .B2(n11026), .C1(
        n9571), .C2(P2_U3088), .ZN(P2_U3305) );
  INV_X1 U13483 ( .A(n11028), .ZN(n11057) );
  NOR2_X1 U13484 ( .A1(n12338), .A2(n13978), .ZN(n11029) );
  AOI21_X1 U13485 ( .B1(n12333), .B2(n14276), .A(n11029), .ZN(n11046) );
  OAI22_X1 U13486 ( .A1(n11030), .A2(n12338), .B1(n13978), .B2(n12340), .ZN(
        n11031) );
  XNOR2_X1 U13487 ( .A(n11031), .B(n12341), .ZN(n11045) );
  INV_X1 U13488 ( .A(n11033), .ZN(n11036) );
  INV_X1 U13489 ( .A(n11034), .ZN(n11035) );
  NAND2_X1 U13490 ( .A1(n14277), .A2(n6638), .ZN(n11038) );
  NAND2_X1 U13491 ( .A1(n6640), .A2(n14062), .ZN(n11037) );
  NAND2_X1 U13492 ( .A1(n11038), .A2(n11037), .ZN(n11039) );
  XNOR2_X1 U13493 ( .A(n11039), .B(n12242), .ZN(n11041) );
  NOR2_X1 U13494 ( .A1(n12338), .A2(n11060), .ZN(n11040) );
  AOI21_X1 U13495 ( .B1(n12333), .B2(n14277), .A(n11040), .ZN(n11042) );
  AND2_X1 U13496 ( .A1(n11041), .A2(n11042), .ZN(n11061) );
  INV_X1 U13497 ( .A(n11041), .ZN(n11044) );
  INV_X1 U13498 ( .A(n11042), .ZN(n11043) );
  NAND2_X1 U13499 ( .A1(n11044), .A2(n11043), .ZN(n11062) );
  XNOR2_X1 U13500 ( .A(n11045), .B(n11046), .ZN(n13972) );
  OAI22_X1 U13501 ( .A1(n14088), .A2(n12338), .B1(n14087), .B2(n12340), .ZN(
        n11047) );
  XNOR2_X1 U13502 ( .A(n11047), .B(n12341), .ZN(n11199) );
  AOI22_X1 U13503 ( .A1(n12333), .A2(n14274), .B1(n6638), .B2(n14074), .ZN(
        n11198) );
  XNOR2_X1 U13504 ( .A(n11199), .B(n11198), .ZN(n11049) );
  OAI211_X1 U13505 ( .C1(n11050), .C2(n11049), .A(n11202), .B(n13994), .ZN(
        n11056) );
  OR2_X1 U13506 ( .A1(n14005), .A2(n14087), .ZN(n11054) );
  INV_X1 U13507 ( .A(n14925), .ZN(n13964) );
  NAND2_X1 U13508 ( .A1(n13964), .A2(n14276), .ZN(n11052) );
  NAND2_X1 U13509 ( .A1(n13997), .A2(n14273), .ZN(n11051) );
  AND4_X1 U13510 ( .A1(n11054), .A2(n11053), .A3(n11052), .A4(n11051), .ZN(
        n11055) );
  OAI211_X1 U13511 ( .C1(n14941), .C2(n11057), .A(n11056), .B(n11055), .ZN(
        P1_U3213) );
  AOI22_X1 U13512 ( .A1(n13987), .A2(n11058), .B1(P1_REG3_REG_5__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11059) );
  OAI21_X1 U13513 ( .B1(n14005), .B2(n11060), .A(n11059), .ZN(n11068) );
  INV_X1 U13514 ( .A(n11061), .ZN(n11063) );
  NAND2_X1 U13515 ( .A1(n11063), .A2(n11062), .ZN(n11064) );
  XNOR2_X1 U13516 ( .A(n11065), .B(n11064), .ZN(n11066) );
  NOR2_X1 U13517 ( .A1(n11066), .A2(n14932), .ZN(n11067) );
  AOI211_X1 U13518 ( .C1(n11069), .C2(n14001), .A(n11068), .B(n11067), .ZN(
        n11070) );
  INV_X1 U13519 ( .A(n11070), .ZN(P1_U3227) );
  NAND2_X1 U13520 ( .A1(n11071), .A2(n14017), .ZN(n11074) );
  AOI22_X1 U13521 ( .A1(n11700), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n11699), 
        .B2(n11072), .ZN(n11073) );
  XNOR2_X1 U13522 ( .A(n11091), .B(P1_REG3_REG_10__SCAN_IN), .ZN(n11510) );
  NAND2_X1 U13523 ( .A1(n11751), .A2(n11510), .ZN(n11078) );
  NAND2_X1 U13524 ( .A1(n11774), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n11077) );
  NAND2_X1 U13525 ( .A1(n11093), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n11076) );
  NAND2_X1 U13526 ( .A1(n11775), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n11075) );
  NAND4_X1 U13527 ( .A1(n11078), .A2(n11077), .A3(n11076), .A4(n11075), .ZN(
        n14271) );
  XNOR2_X1 U13528 ( .A(n14097), .B(n14924), .ZN(n14229) );
  OR2_X1 U13529 ( .A1(n11079), .A2(n14025), .ZN(n11082) );
  AOI22_X1 U13530 ( .A1(n11700), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n11699), 
        .B2(n11080), .ZN(n11081) );
  NAND2_X1 U13531 ( .A1(n11082), .A2(n11081), .ZN(n14078) );
  INV_X1 U13532 ( .A(n14078), .ZN(n14079) );
  INV_X1 U13533 ( .A(n14273), .ZN(n11084) );
  XNOR2_X1 U13534 ( .A(n14078), .B(n14272), .ZN(n14091) );
  NOR2_X1 U13535 ( .A1(n11087), .A2(n14229), .ZN(n11376) );
  AOI211_X1 U13536 ( .C1(n14229), .C2(n11087), .A(n15109), .B(n11376), .ZN(
        n11088) );
  AOI21_X1 U13537 ( .B1(n14571), .B2(n14272), .A(n11088), .ZN(n15186) );
  INV_X1 U13538 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n11089) );
  INV_X1 U13539 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n11090) );
  OAI21_X1 U13540 ( .B1(n11091), .B2(n11089), .A(n11090), .ZN(n11092) );
  NAND2_X1 U13541 ( .A1(n11092), .A2(n11386), .ZN(n14940) );
  INV_X1 U13542 ( .A(n14940), .ZN(n11483) );
  NAND2_X1 U13543 ( .A1(n11751), .A2(n11483), .ZN(n11097) );
  NAND2_X1 U13544 ( .A1(n11774), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n11096) );
  NAND2_X1 U13545 ( .A1(n14012), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n11095) );
  NAND2_X1 U13546 ( .A1(n11093), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n11094) );
  NAND4_X1 U13547 ( .A1(n11097), .A2(n11096), .A3(n11095), .A4(n11094), .ZN(
        n14270) );
  AOI211_X1 U13548 ( .C1(n14097), .C2(n11122), .A(n15161), .B(n11482), .ZN(
        n11098) );
  AOI21_X1 U13549 ( .B1(n14573), .B2(n14270), .A(n11098), .ZN(n15185) );
  INV_X1 U13550 ( .A(n15185), .ZN(n11101) );
  INV_X1 U13551 ( .A(n14097), .ZN(n15188) );
  AOI22_X1 U13552 ( .A1(n15129), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n11510), 
        .B2(n15114), .ZN(n11099) );
  OAI21_X1 U13553 ( .B1(n15116), .B2(n15188), .A(n11099), .ZN(n11100) );
  AOI21_X1 U13554 ( .B1(n11101), .B2(n15125), .A(n11100), .ZN(n11106) );
  INV_X1 U13555 ( .A(n14091), .ZN(n14231) );
  OAI21_X1 U13556 ( .B1(n11104), .B2(n14229), .A(n11416), .ZN(n15190) );
  NAND2_X1 U13557 ( .A1(n15190), .A2(n14516), .ZN(n11105) );
  OAI211_X1 U13558 ( .C1(n15186), .C2(n15129), .A(n11106), .B(n11105), .ZN(
        P1_U3283) );
  INV_X1 U13559 ( .A(n11107), .ZN(n11109) );
  INV_X1 U13560 ( .A(SI_24_), .ZN(n11108) );
  OAI222_X1 U13561 ( .A1(n11110), .A2(P3_U3151), .B1(n14722), .B2(n11109), 
        .C1(n11108), .C2(n14721), .ZN(P3_U3271) );
  AOI22_X1 U13562 ( .A1(n15292), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n11247), 
        .B2(n15279), .ZN(n11111) );
  OAI21_X1 U13563 ( .B1(n11250), .B2(n15282), .A(n11111), .ZN(n11114) );
  NOR2_X1 U13564 ( .A1(n11112), .A2(n13738), .ZN(n11113) );
  AOI211_X1 U13565 ( .C1(n11115), .C2(n15285), .A(n11114), .B(n11113), .ZN(
        n11116) );
  OAI21_X1 U13566 ( .B1(n15292), .B2(n11117), .A(n11116), .ZN(P2_U3253) );
  OR2_X1 U13567 ( .A1(n11118), .A2(n14231), .ZN(n11119) );
  AND2_X1 U13568 ( .A1(n11120), .A2(n11119), .ZN(n11130) );
  INV_X1 U13569 ( .A(n11130), .ZN(n11156) );
  AOI21_X1 U13570 ( .B1(n11121), .B2(n14078), .A(n15161), .ZN(n11123) );
  NAND2_X1 U13571 ( .A1(n11123), .A2(n11122), .ZN(n11152) );
  OAI21_X1 U13572 ( .B1(n14079), .B2(n15187), .A(n11152), .ZN(n11131) );
  OAI21_X1 U13573 ( .B1(n11125), .B2(n14091), .A(n11124), .ZN(n11126) );
  NAND2_X1 U13574 ( .A1(n11126), .A2(n14971), .ZN(n11128) );
  AOI22_X1 U13575 ( .A1(n14571), .A2(n14273), .B1(n14271), .B2(n14573), .ZN(
        n11127) );
  OAI211_X1 U13576 ( .C1(n11130), .C2(n11129), .A(n11128), .B(n11127), .ZN(
        n11153) );
  AOI211_X1 U13577 ( .C1(n15173), .C2(n11156), .A(n11131), .B(n11153), .ZN(
        n11133) );
  OR2_X1 U13578 ( .A1(n11133), .A2(n15200), .ZN(n11132) );
  OAI21_X1 U13579 ( .B1(n15202), .B2(n9759), .A(n11132), .ZN(P1_U3537) );
  INV_X1 U13580 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n11135) );
  OR2_X1 U13581 ( .A1(n11133), .A2(n15192), .ZN(n11134) );
  OAI21_X1 U13582 ( .B1(n15194), .B2(n11135), .A(n11134), .ZN(P1_U3486) );
  NAND2_X1 U13583 ( .A1(n11745), .A2(n11136), .ZN(n11138) );
  OAI211_X1 U13584 ( .C1(n11139), .C2(n13852), .A(n11138), .B(n11137), .ZN(
        P2_U3304) );
  INV_X1 U13585 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11746) );
  NAND2_X1 U13586 ( .A1(n11745), .A2(n14691), .ZN(n11140) );
  OAI211_X1 U13587 ( .C1(n11746), .C2(n14694), .A(n11140), .B(n14258), .ZN(
        P1_U3332) );
  AOI21_X1 U13588 ( .B1(n11141), .B2(n12088), .A(n15456), .ZN(n11145) );
  OAI22_X1 U13589 ( .A1(n11142), .A2(n15450), .B1(n11443), .B2(n15448), .ZN(
        n11143) );
  AOI21_X1 U13590 ( .B1(n11145), .B2(n11144), .A(n11143), .ZN(n11300) );
  XNOR2_X1 U13591 ( .A(n11146), .B(n12088), .ZN(n11298) );
  AOI22_X1 U13592 ( .A1(n12871), .A2(P3_REG2_REG_9__SCAN_IN), .B1(n15473), 
        .B2(n11147), .ZN(n11148) );
  OAI21_X1 U13593 ( .B1(n12867), .B2(n11310), .A(n11148), .ZN(n11149) );
  AOI21_X1 U13594 ( .B1(n11298), .B2(n12869), .A(n11149), .ZN(n11150) );
  OAI21_X1 U13595 ( .B1(n11300), .B2(n12871), .A(n11150), .ZN(P3_U3224) );
  AOI22_X1 U13596 ( .A1(n14737), .A2(n14078), .B1(n11364), .B2(n15114), .ZN(
        n11151) );
  OAI21_X1 U13597 ( .B1(n11152), .B2(n14519), .A(n11151), .ZN(n11155) );
  MUX2_X1 U13598 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n11153), .S(n14552), .Z(
        n11154) );
  AOI211_X1 U13599 ( .C1(n15126), .C2(n11156), .A(n11155), .B(n11154), .ZN(
        n11157) );
  INV_X1 U13600 ( .A(n11157), .ZN(P1_U3284) );
  XNOR2_X1 U13601 ( .A(n11170), .B(n6838), .ZN(n11163) );
  NAND2_X1 U13602 ( .A1(n11957), .A2(n13523), .ZN(n11162) );
  NAND2_X1 U13603 ( .A1(n11163), .A2(n11162), .ZN(n11241) );
  OAI21_X1 U13604 ( .B1(n11163), .B2(n11162), .A(n11241), .ZN(n11164) );
  AOI21_X1 U13605 ( .B1(n11165), .B2(n11164), .A(n6783), .ZN(n11173) );
  NOR2_X1 U13606 ( .A1(n13476), .A2(n11166), .ZN(n11167) );
  AOI211_X1 U13607 ( .C1(n13467), .C2(n11169), .A(n11168), .B(n11167), .ZN(
        n11172) );
  NAND2_X1 U13608 ( .A1(n11170), .A2(n13501), .ZN(n11171) );
  OAI211_X1 U13609 ( .C1(n11173), .C2(n13503), .A(n11172), .B(n11171), .ZN(
        P2_U3208) );
  NAND2_X1 U13610 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n11180), .ZN(n11177) );
  INV_X1 U13611 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n11175) );
  INV_X1 U13612 ( .A(n11177), .ZN(n11174) );
  AOI21_X1 U13613 ( .B1(n11175), .B2(n15277), .A(n11174), .ZN(n15274) );
  OAI21_X1 U13614 ( .B1(n11182), .B2(n10697), .A(n11176), .ZN(n15273) );
  NAND2_X1 U13615 ( .A1(n15274), .A2(n15273), .ZN(n15272) );
  NAND2_X1 U13616 ( .A1(n11177), .A2(n15272), .ZN(n11591) );
  XNOR2_X1 U13617 ( .A(n11596), .B(n11591), .ZN(n11178) );
  NOR2_X1 U13618 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n11178), .ZN(n11593) );
  AOI21_X1 U13619 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n11178), .A(n11593), 
        .ZN(n11192) );
  INV_X1 U13620 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n14863) );
  NOR2_X1 U13621 ( .A1(n11180), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n11179) );
  AOI21_X1 U13622 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n11180), .A(n11179), 
        .ZN(n15266) );
  INV_X1 U13623 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n14871) );
  OAI21_X1 U13624 ( .B1(n11182), .B2(n14871), .A(n11181), .ZN(n15265) );
  NAND2_X1 U13625 ( .A1(n15266), .A2(n15265), .ZN(n15263) );
  OAI21_X1 U13626 ( .B1(n15277), .B2(n14863), .A(n15263), .ZN(n11595) );
  INV_X1 U13627 ( .A(n11595), .ZN(n11183) );
  XNOR2_X1 U13628 ( .A(n11596), .B(n11183), .ZN(n11184) );
  NAND2_X1 U13629 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n11184), .ZN(n11598) );
  OAI211_X1 U13630 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n11184), .A(n15264), 
        .B(n11598), .ZN(n11188) );
  NOR2_X1 U13631 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11185), .ZN(n11186) );
  AOI21_X1 U13632 ( .B1(n15270), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n11186), 
        .ZN(n11187) );
  OAI211_X1 U13633 ( .C1(n15278), .C2(n11189), .A(n11188), .B(n11187), .ZN(
        n11190) );
  INV_X1 U13634 ( .A(n11190), .ZN(n11191) );
  OAI21_X1 U13635 ( .B1(n11192), .B2(n15220), .A(n11191), .ZN(P2_U3232) );
  NAND2_X1 U13636 ( .A1(n14075), .A2(n6640), .ZN(n11194) );
  NAND2_X1 U13637 ( .A1(n14273), .A2(n6638), .ZN(n11193) );
  NAND2_X1 U13638 ( .A1(n11194), .A2(n11193), .ZN(n11195) );
  XNOR2_X1 U13639 ( .A(n11195), .B(n12341), .ZN(n11356) );
  NAND2_X1 U13640 ( .A1(n12333), .A2(n14273), .ZN(n11197) );
  NAND2_X1 U13641 ( .A1(n14075), .A2(n6638), .ZN(n11196) );
  NAND2_X1 U13642 ( .A1(n11197), .A2(n11196), .ZN(n11357) );
  XNOR2_X1 U13643 ( .A(n11356), .B(n11357), .ZN(n11205) );
  INV_X1 U13644 ( .A(n11198), .ZN(n11200) );
  NAND2_X1 U13645 ( .A1(n11200), .A2(n11199), .ZN(n11201) );
  INV_X1 U13646 ( .A(n11355), .ZN(n11203) );
  AOI21_X1 U13647 ( .B1(n11205), .B2(n11204), .A(n11203), .ZN(n11212) );
  NAND2_X1 U13648 ( .A1(n13987), .A2(n11206), .ZN(n11207) );
  OAI211_X1 U13649 ( .C1(n14941), .C2(n11209), .A(n11208), .B(n11207), .ZN(
        n11210) );
  AOI21_X1 U13650 ( .B1(n14075), .B2(n14937), .A(n11210), .ZN(n11211) );
  OAI21_X1 U13651 ( .B1(n11212), .B2(n14932), .A(n11211), .ZN(P1_U3221) );
  XNOR2_X1 U13652 ( .A(n11213), .B(n12021), .ZN(n15514) );
  OAI21_X1 U13653 ( .B1(n11215), .B2(n12021), .A(n11214), .ZN(n11216) );
  NAND2_X1 U13654 ( .A1(n11216), .A2(n15466), .ZN(n11218) );
  AOI22_X1 U13655 ( .A1(n12546), .A2(n15464), .B1(n15461), .B2(n12544), .ZN(
        n11217) );
  OAI211_X1 U13656 ( .C1(n15470), .C2(n15514), .A(n11218), .B(n11217), .ZN(
        n15515) );
  MUX2_X1 U13657 ( .A(n15515), .B(P3_REG2_REG_8__SCAN_IN), .S(n12871), .Z(
        n11219) );
  INV_X1 U13658 ( .A(n11219), .ZN(n11222) );
  NOR2_X1 U13659 ( .A1(n11220), .A2(n15521), .ZN(n15516) );
  AOI22_X1 U13660 ( .A1(n14782), .A2(n15516), .B1(n15473), .B2(n12433), .ZN(
        n11221) );
  OAI211_X1 U13661 ( .C1(n15514), .C2(n12752), .A(n11222), .B(n11221), .ZN(
        P3_U3225) );
  INV_X1 U13662 ( .A(n11447), .ZN(n11237) );
  INV_X1 U13663 ( .A(n11223), .ZN(n11224) );
  NAND2_X1 U13664 ( .A1(n11224), .A2(n12543), .ZN(n11225) );
  NAND2_X1 U13665 ( .A1(n11226), .A2(n11225), .ZN(n11228) );
  XNOR2_X1 U13666 ( .A(n12416), .B(n11446), .ZN(n11227) );
  OR2_X2 U13667 ( .A1(n11228), .A2(n11227), .ZN(n11341) );
  NAND2_X1 U13668 ( .A1(n11228), .A2(n11227), .ZN(n11229) );
  AND2_X2 U13669 ( .A1(n11341), .A2(n11229), .ZN(n11230) );
  OAI21_X1 U13670 ( .B1(n14777), .B2(n11230), .A(n11342), .ZN(n11231) );
  NAND2_X1 U13671 ( .A1(n11231), .A2(n12522), .ZN(n11235) );
  INV_X1 U13672 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11232) );
  NOR2_X1 U13673 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11232), .ZN(n11317) );
  OAI22_X1 U13674 ( .A1(n11443), .A2(n12527), .B1(n12526), .B2(n14762), .ZN(
        n11233) );
  AOI211_X1 U13675 ( .C1(n12103), .C2(n12517), .A(n11317), .B(n11233), .ZN(
        n11234) );
  OAI211_X1 U13676 ( .C1(n11237), .C2(n11236), .A(n11235), .B(n11234), .ZN(
        P3_U3176) );
  AND2_X1 U13677 ( .A1(n11957), .A2(n13522), .ZN(n11240) );
  XNOR2_X1 U13678 ( .A(n11238), .B(n11961), .ZN(n11239) );
  NOR2_X1 U13679 ( .A1(n11239), .A2(n11240), .ZN(n11289) );
  AOI21_X1 U13680 ( .B1(n11240), .B2(n11239), .A(n11289), .ZN(n11243) );
  OAI21_X1 U13681 ( .B1(n11243), .B2(n11242), .A(n11291), .ZN(n11244) );
  NAND2_X1 U13682 ( .A1(n11244), .A2(n13454), .ZN(n11249) );
  NAND2_X1 U13683 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n15248)
         );
  OAI21_X1 U13684 ( .B1(n13476), .B2(n11245), .A(n15248), .ZN(n11246) );
  AOI21_X1 U13685 ( .B1(n11247), .B2(n13467), .A(n11246), .ZN(n11248) );
  OAI211_X1 U13686 ( .C1(n11250), .C2(n13461), .A(n11249), .B(n11248), .ZN(
        P2_U3196) );
  INV_X1 U13687 ( .A(n11251), .ZN(n11252) );
  OAI222_X1 U13688 ( .A1(P3_U3151), .A2(n11254), .B1(n14721), .B2(n11253), 
        .C1(n14722), .C2(n11252), .ZN(P3_U3270) );
  NOR2_X1 U13689 ( .A1(n7439), .A2(n11255), .ZN(n11257) );
  NAND2_X1 U13690 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n15417), .ZN(n11258) );
  OAI21_X1 U13691 ( .B1(P3_REG1_REG_10__SCAN_IN), .B2(n15417), .A(n11258), 
        .ZN(n15423) );
  NOR2_X1 U13692 ( .A1(n11325), .A2(n11259), .ZN(n11260) );
  INV_X1 U13693 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14806) );
  INV_X1 U13694 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14802) );
  AOI22_X1 U13695 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n11282), .B1(n11892), 
        .B2(n14802), .ZN(n11261) );
  AOI21_X1 U13696 ( .B1(n11262), .B2(n11261), .A(n11854), .ZN(n11288) );
  NOR2_X1 U13697 ( .A1(n7439), .A2(n11263), .ZN(n11265) );
  NOR2_X1 U13698 ( .A1(n11265), .A2(n11264), .ZN(n15416) );
  NAND2_X1 U13699 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n15417), .ZN(n11266) );
  OAI21_X1 U13700 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n15417), .A(n11266), 
        .ZN(n15415) );
  NOR2_X1 U13701 ( .A1(n11325), .A2(n11267), .ZN(n11269) );
  INV_X1 U13702 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11313) );
  INV_X1 U13703 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n14784) );
  AOI22_X1 U13704 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n11282), .B1(n11892), 
        .B2(n14784), .ZN(n11890) );
  XNOR2_X1 U13705 ( .A(n11891), .B(n11890), .ZN(n11286) );
  INV_X1 U13706 ( .A(n15438), .ZN(n15404) );
  MUX2_X1 U13707 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n6642), .Z(n11869) );
  XNOR2_X1 U13708 ( .A(n11869), .B(n11892), .ZN(n11871) );
  MUX2_X1 U13709 ( .A(n11313), .B(n14806), .S(n6642), .Z(n11277) );
  NAND2_X1 U13710 ( .A1(n11277), .A2(n11325), .ZN(n11279) );
  MUX2_X1 U13711 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n6642), .Z(n11270) );
  NOR2_X1 U13712 ( .A1(n11270), .A2(n15417), .ZN(n11276) );
  AOI21_X1 U13713 ( .B1(n11270), .B2(n15417), .A(n11276), .ZN(n11271) );
  INV_X1 U13714 ( .A(n11271), .ZN(n15432) );
  INV_X1 U13715 ( .A(n11272), .ZN(n11273) );
  NOR2_X1 U13716 ( .A1(n15432), .A2(n15433), .ZN(n15431) );
  NOR2_X1 U13717 ( .A1(n11276), .A2(n15431), .ZN(n11315) );
  OAI21_X1 U13718 ( .B1(n11277), .B2(n11325), .A(n11279), .ZN(n11316) );
  NAND2_X1 U13719 ( .A1(n11279), .A2(n11278), .ZN(n11870) );
  XNOR2_X1 U13720 ( .A(n11871), .B(n11870), .ZN(n11284) );
  INV_X1 U13721 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n13261) );
  NOR2_X1 U13722 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13261), .ZN(n11345) );
  NOR2_X1 U13723 ( .A1(n15421), .A2(n11280), .ZN(n11281) );
  AOI211_X1 U13724 ( .C1(n15430), .C2(n11282), .A(n11345), .B(n11281), .ZN(
        n11283) );
  OAI21_X1 U13725 ( .B1(n11284), .B2(n15434), .A(n11283), .ZN(n11285) );
  AOI21_X1 U13726 ( .B1(n11286), .B2(n15404), .A(n11285), .ZN(n11287) );
  OAI21_X1 U13727 ( .B1(n11288), .B2(n15425), .A(n11287), .ZN(P3_U3194) );
  INV_X1 U13728 ( .A(n11289), .ZN(n11290) );
  NAND2_X1 U13729 ( .A1(n11291), .A2(n11290), .ZN(n11458) );
  NAND2_X1 U13730 ( .A1(n11957), .A2(n11567), .ZN(n11455) );
  XNOR2_X1 U13731 ( .A(n14885), .B(n11961), .ZN(n11454) );
  XOR2_X1 U13732 ( .A(n11455), .B(n11454), .Z(n11457) );
  XNOR2_X1 U13733 ( .A(n11458), .B(n11457), .ZN(n11297) );
  OAI22_X1 U13734 ( .A1(n13476), .A2(n11292), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9712), .ZN(n11293) );
  AOI21_X1 U13735 ( .B1(n11294), .B2(n13467), .A(n11293), .ZN(n11296) );
  NAND2_X1 U13736 ( .A1(n14885), .A2(n13501), .ZN(n11295) );
  OAI211_X1 U13737 ( .C1(n11297), .C2(n13503), .A(n11296), .B(n11295), .ZN(
        P2_U3206) );
  INV_X1 U13738 ( .A(n12951), .ZN(n12957) );
  NAND2_X1 U13739 ( .A1(n11298), .A2(n15497), .ZN(n11299) );
  AND2_X1 U13740 ( .A1(n11300), .A2(n11299), .ZN(n11308) );
  MUX2_X1 U13741 ( .A(n11301), .B(n11308), .S(n15547), .Z(n11302) );
  OAI21_X1 U13742 ( .B1(n12957), .B2(n11310), .A(n11302), .ZN(P3_U3468) );
  INV_X1 U13743 ( .A(n11303), .ZN(n11305) );
  OAI222_X1 U13744 ( .A1(n11306), .A2(P3_U3151), .B1(n14722), .B2(n11305), 
        .C1(n11304), .C2(n14721), .ZN(P3_U3269) );
  INV_X1 U13745 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n11307) );
  MUX2_X1 U13746 ( .A(n11308), .B(n11307), .S(n15526), .Z(n11309) );
  OAI21_X1 U13747 ( .B1(n13014), .B2(n11310), .A(n11309), .ZN(P3_U3417) );
  AOI21_X1 U13748 ( .B1(n11313), .B2(n11312), .A(n11311), .ZN(n11327) );
  AOI21_X1 U13749 ( .B1(n11316), .B2(n11315), .A(n11314), .ZN(n11319) );
  AOI21_X1 U13750 ( .B1(n15405), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n11317), 
        .ZN(n11318) );
  OAI21_X1 U13751 ( .B1(n11319), .B2(n15434), .A(n11318), .ZN(n11324) );
  AOI21_X1 U13752 ( .B1(n14806), .B2(n11321), .A(n11320), .ZN(n11322) );
  NOR2_X1 U13753 ( .A1(n11322), .A2(n15425), .ZN(n11323) );
  AOI211_X1 U13754 ( .C1(n15430), .C2(n11325), .A(n11324), .B(n11323), .ZN(
        n11326) );
  OAI21_X1 U13755 ( .B1(n11327), .B2(n15438), .A(n11326), .ZN(P3_U3193) );
  INV_X1 U13756 ( .A(n12093), .ZN(n12024) );
  XNOR2_X1 U13757 ( .A(n11328), .B(n12024), .ZN(n15523) );
  OAI211_X1 U13758 ( .C1(n11330), .C2(n12093), .A(n11329), .B(n15466), .ZN(
        n11332) );
  AOI22_X1 U13759 ( .A1(n12542), .A2(n15461), .B1(n15464), .B2(n12544), .ZN(
        n11331) );
  OAI211_X1 U13760 ( .C1(n15470), .C2(n15523), .A(n11332), .B(n11331), .ZN(
        n15525) );
  NAND2_X1 U13761 ( .A1(n15525), .A2(n15477), .ZN(n11338) );
  INV_X1 U13762 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11334) );
  OAI22_X1 U13763 ( .A1(n15477), .A2(n11334), .B1(n11333), .B2(n15443), .ZN(
        n11335) );
  AOI21_X1 U13764 ( .B1(n12885), .B2(n11336), .A(n11335), .ZN(n11337) );
  OAI211_X1 U13765 ( .C1(n15523), .C2(n12752), .A(n11338), .B(n11337), .ZN(
        P3_U3223) );
  XNOR2_X1 U13766 ( .A(n12390), .B(n11346), .ZN(n11340) );
  INV_X1 U13767 ( .A(n11340), .ZN(n11339) );
  NAND2_X1 U13768 ( .A1(n11339), .A2(n12541), .ZN(n11523) );
  NAND2_X1 U13769 ( .A1(n11340), .A2(n14762), .ZN(n11521) );
  NAND2_X1 U13770 ( .A1(n11523), .A2(n11521), .ZN(n11343) );
  AND2_X2 U13771 ( .A1(n11342), .A2(n11341), .ZN(n11522) );
  XOR2_X1 U13772 ( .A(n11343), .B(n11522), .Z(n11349) );
  OAI22_X1 U13773 ( .A1(n14777), .A2(n12527), .B1(n12526), .B2(n14778), .ZN(
        n11344) );
  AOI211_X1 U13774 ( .C1(n11346), .C2(n12517), .A(n11345), .B(n11344), .ZN(
        n11348) );
  NAND2_X1 U13775 ( .A1(n12530), .A2(n14781), .ZN(n11347) );
  OAI211_X1 U13776 ( .C1(n11349), .C2(n12520), .A(n11348), .B(n11347), .ZN(
        P3_U3164) );
  INV_X1 U13777 ( .A(n11665), .ZN(n11812) );
  OAI222_X1 U13778 ( .A1(n13852), .A2(n11351), .B1(n13854), .B2(n11812), .C1(
        n11350), .C2(P2_U3088), .ZN(P2_U3303) );
  INV_X1 U13779 ( .A(n14272), .ZN(n14080) );
  OAI22_X1 U13780 ( .A1(n14079), .A2(n12338), .B1(n14080), .B2(n6646), .ZN(
        n11494) );
  NAND2_X1 U13781 ( .A1(n14078), .A2(n6640), .ZN(n11353) );
  NAND2_X1 U13782 ( .A1(n14272), .A2(n6638), .ZN(n11352) );
  NAND2_X1 U13783 ( .A1(n11353), .A2(n11352), .ZN(n11354) );
  XNOR2_X1 U13784 ( .A(n11354), .B(n12341), .ZN(n11495) );
  XOR2_X1 U13785 ( .A(n11494), .B(n11495), .Z(n11359) );
  OAI21_X1 U13786 ( .B1(n11359), .B2(n11358), .A(n11497), .ZN(n11360) );
  NAND2_X1 U13787 ( .A1(n11360), .A2(n13994), .ZN(n11366) );
  NAND2_X1 U13788 ( .A1(n13964), .A2(n14273), .ZN(n11362) );
  OAI211_X1 U13789 ( .C1(n14924), .C2(n14926), .A(n11362), .B(n11361), .ZN(
        n11363) );
  AOI21_X1 U13790 ( .B1(n11364), .B2(n14001), .A(n11363), .ZN(n11365) );
  OAI211_X1 U13791 ( .C1(n14079), .C2(n14005), .A(n11366), .B(n11365), .ZN(
        P1_U3231) );
  NAND2_X1 U13792 ( .A1(n11367), .A2(n14017), .ZN(n11369) );
  AOI22_X1 U13793 ( .A1(n11700), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n11699), 
        .B2(n14338), .ZN(n11368) );
  NAND2_X1 U13794 ( .A1(n11395), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n11397) );
  INV_X1 U13795 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n11370) );
  NAND2_X1 U13796 ( .A1(n11397), .A2(n11370), .ZN(n11371) );
  NAND2_X1 U13797 ( .A1(n11404), .A2(n11371), .ZN(n14911) );
  INV_X1 U13798 ( .A(n14911), .ZN(n11410) );
  NAND2_X1 U13799 ( .A1(n11751), .A2(n11410), .ZN(n11375) );
  NAND2_X1 U13800 ( .A1(n11774), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n11374) );
  NAND2_X1 U13801 ( .A1(n14011), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11373) );
  NAND2_X1 U13802 ( .A1(n14012), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n11372) );
  OR2_X1 U13803 ( .A1(n14909), .A2(n13999), .ZN(n14119) );
  NAND2_X1 U13804 ( .A1(n14909), .A2(n13999), .ZN(n14118) );
  NAND2_X1 U13805 ( .A1(n11377), .A2(n14017), .ZN(n11380) );
  AOI22_X1 U13806 ( .A1(n11700), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n11699), 
        .B2(n11378), .ZN(n11379) );
  NAND2_X2 U13807 ( .A1(n11380), .A2(n11379), .ZN(n14938) );
  NOR2_X1 U13808 ( .A1(n11515), .A2(n14270), .ZN(n11381) );
  INV_X1 U13809 ( .A(n14270), .ZN(n12218) );
  NAND2_X1 U13810 ( .A1(n11382), .A2(n14017), .ZN(n11384) );
  AOI22_X1 U13811 ( .A1(n11700), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n11699), 
        .B2(n14337), .ZN(n11383) );
  AND2_X1 U13812 ( .A1(n11386), .A2(n11385), .ZN(n11387) );
  NOR2_X1 U13813 ( .A1(n11395), .A2(n11387), .ZN(n14736) );
  NAND2_X1 U13814 ( .A1(n11751), .A2(n14736), .ZN(n11391) );
  NAND2_X1 U13815 ( .A1(n11774), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n11390) );
  NAND2_X1 U13816 ( .A1(n14012), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n11389) );
  NAND2_X1 U13817 ( .A1(n14011), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n11388) );
  NAND4_X1 U13818 ( .A1(n11391), .A2(n11390), .A3(n11389), .A4(n11388), .ZN(
        n14269) );
  INV_X1 U13819 ( .A(n14269), .ZN(n14927) );
  XNOR2_X1 U13820 ( .A(n14738), .B(n14927), .ZN(n14730) );
  INV_X1 U13821 ( .A(n14738), .ZN(n14746) );
  NAND2_X1 U13822 ( .A1(n11392), .A2(n14017), .ZN(n11394) );
  AOI22_X1 U13823 ( .A1(n11700), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n11699), 
        .B2(n15023), .ZN(n11393) );
  OR2_X1 U13824 ( .A1(n11395), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n11396) );
  AND2_X1 U13825 ( .A1(n11397), .A2(n11396), .ZN(n11429) );
  NAND2_X1 U13826 ( .A1(n11751), .A2(n11429), .ZN(n11401) );
  NAND2_X1 U13827 ( .A1(n11774), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n11400) );
  NAND2_X1 U13828 ( .A1(n11715), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n11399) );
  NAND2_X1 U13829 ( .A1(n14011), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11398) );
  NAND4_X1 U13830 ( .A1(n11401), .A2(n11400), .A3(n11399), .A4(n11398), .ZN(
        n14268) );
  XNOR2_X1 U13831 ( .A(n14112), .B(n14268), .ZN(n14232) );
  INV_X1 U13832 ( .A(n14232), .ZN(n11419) );
  INV_X1 U13833 ( .A(n14268), .ZN(n14901) );
  XOR2_X1 U13834 ( .A(n14234), .B(n11540), .Z(n14972) );
  INV_X1 U13835 ( .A(n14972), .ZN(n11425) );
  INV_X1 U13836 ( .A(n14909), .ZN(n14968) );
  INV_X1 U13837 ( .A(n11552), .ZN(n11402) );
  OAI211_X1 U13838 ( .C1(n14968), .C2(n11432), .A(n11402), .B(n15120), .ZN(
        n14967) );
  INV_X1 U13839 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n11403) );
  AND2_X1 U13840 ( .A1(n11404), .A2(n11403), .ZN(n11405) );
  NOR2_X1 U13841 ( .A1(n11542), .A2(n11405), .ZN(n14002) );
  NAND2_X1 U13842 ( .A1(n11751), .A2(n14002), .ZN(n11409) );
  NAND2_X1 U13843 ( .A1(n11774), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n11408) );
  NAND2_X1 U13844 ( .A1(n14012), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n11407) );
  NAND2_X1 U13845 ( .A1(n14011), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n11406) );
  INV_X1 U13846 ( .A(n14912), .ZN(n14572) );
  AOI22_X1 U13847 ( .A1(n14572), .A2(n14573), .B1(n14571), .B2(n14268), .ZN(
        n14966) );
  NAND2_X1 U13848 ( .A1(n15114), .A2(n11410), .ZN(n11411) );
  OAI211_X1 U13849 ( .C1(n14967), .C2(n14579), .A(n14966), .B(n11411), .ZN(
        n11414) );
  INV_X1 U13850 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11412) );
  INV_X1 U13851 ( .A(n15129), .ZN(n14552) );
  OAI22_X1 U13852 ( .A1(n14968), .A2(n15116), .B1(n11412), .B2(n14552), .ZN(
        n11413) );
  AOI21_X1 U13853 ( .B1(n11414), .B2(n14552), .A(n11413), .ZN(n11424) );
  OR2_X1 U13854 ( .A1(n14097), .A2(n14271), .ZN(n11415) );
  OR2_X1 U13855 ( .A1(n14738), .A2(n14269), .ZN(n11417) );
  NAND2_X1 U13856 ( .A1(n11418), .A2(n11417), .ZN(n11426) );
  NAND2_X1 U13857 ( .A1(n11426), .A2(n11419), .ZN(n11421) );
  OR2_X1 U13858 ( .A1(n14112), .A2(n14268), .ZN(n11420) );
  NAND2_X1 U13859 ( .A1(n11421), .A2(n11420), .ZN(n11422) );
  OR2_X2 U13860 ( .A1(n11422), .A2(n14234), .ZN(n14965) );
  NAND2_X1 U13861 ( .A1(n11422), .A2(n14234), .ZN(n14964) );
  NAND3_X1 U13862 ( .A1(n14965), .A2(n14964), .A3(n14516), .ZN(n11423) );
  OAI211_X1 U13863 ( .C1(n11425), .C2(n14483), .A(n11424), .B(n11423), .ZN(
        P1_U3279) );
  XNOR2_X1 U13864 ( .A(n11426), .B(n14232), .ZN(n11475) );
  XNOR2_X1 U13865 ( .A(n11427), .B(n14232), .ZN(n11428) );
  NAND2_X1 U13866 ( .A1(n11428), .A2(n14971), .ZN(n11474) );
  INV_X1 U13867 ( .A(n11474), .ZN(n11438) );
  INV_X1 U13868 ( .A(n11429), .ZN(n13939) );
  NAND2_X1 U13869 ( .A1(n14740), .A2(n14112), .ZN(n11430) );
  NAND2_X1 U13870 ( .A1(n11430), .A2(n15120), .ZN(n11431) );
  NOR2_X1 U13871 ( .A1(n11432), .A2(n11431), .ZN(n11472) );
  NAND2_X1 U13872 ( .A1(n11472), .A2(n14352), .ZN(n11436) );
  OR2_X1 U13873 ( .A1(n13999), .A2(n14533), .ZN(n11434) );
  NAND2_X1 U13874 ( .A1(n14269), .A2(n14571), .ZN(n11433) );
  NAND2_X1 U13875 ( .A1(n11434), .A2(n11433), .ZN(n13937) );
  INV_X1 U13876 ( .A(n13937), .ZN(n11435) );
  OAI211_X1 U13877 ( .C1(n14578), .C2(n13939), .A(n11436), .B(n11435), .ZN(
        n11437) );
  OAI21_X1 U13878 ( .B1(n11438), .B2(n11437), .A(n14552), .ZN(n11440) );
  AOI22_X1 U13879 ( .A1(n14112), .A2(n14737), .B1(P1_REG2_REG_13__SCAN_IN), 
        .B2(n15129), .ZN(n11439) );
  OAI211_X1 U13880 ( .C1(n11475), .C2(n14584), .A(n11440), .B(n11439), .ZN(
        P1_U3280) );
  NAND2_X1 U13881 ( .A1(n11329), .A2(n11441), .ZN(n14771) );
  INV_X1 U13882 ( .A(n12106), .ZN(n12097) );
  XNOR2_X1 U13883 ( .A(n14771), .B(n12097), .ZN(n11442) );
  OAI222_X1 U13884 ( .A1(n15448), .A2(n14762), .B1(n15450), .B2(n11443), .C1(
        n11442), .C2(n15456), .ZN(n14803) );
  INV_X1 U13885 ( .A(n14803), .ZN(n11451) );
  OAI21_X1 U13886 ( .B1(n11445), .B2(n12106), .A(n11444), .ZN(n14805) );
  NOR2_X1 U13887 ( .A1(n11446), .A2(n15521), .ZN(n14804) );
  AOI22_X1 U13888 ( .A1(n14782), .A2(n14804), .B1(n15473), .B2(n11447), .ZN(
        n11448) );
  OAI21_X1 U13889 ( .B1(n11313), .B2(n15477), .A(n11448), .ZN(n11449) );
  AOI21_X1 U13890 ( .B1(n14805), .B2(n12869), .A(n11449), .ZN(n11450) );
  OAI21_X1 U13891 ( .B1(n11451), .B2(n12871), .A(n11450), .ZN(P3_U3222) );
  XNOR2_X1 U13892 ( .A(n14849), .B(n6838), .ZN(n11453) );
  NAND2_X1 U13893 ( .A1(n11957), .A2(n13521), .ZN(n11452) );
  NAND2_X1 U13894 ( .A1(n11453), .A2(n11452), .ZN(n11558) );
  OAI21_X1 U13895 ( .B1(n11453), .B2(n11452), .A(n11558), .ZN(n11460) );
  INV_X1 U13896 ( .A(n11454), .ZN(n11456) );
  AOI21_X1 U13897 ( .B1(n11460), .B2(n11459), .A(n11913), .ZN(n11467) );
  INV_X1 U13898 ( .A(n14843), .ZN(n11464) );
  NAND2_X1 U13899 ( .A1(n13475), .A2(n11567), .ZN(n11461) );
  OAI21_X1 U13900 ( .B1(n13492), .B2(n11581), .A(n11461), .ZN(n14840) );
  NAND2_X1 U13901 ( .A1(n13496), .A2(n14840), .ZN(n11463) );
  OAI211_X1 U13902 ( .C1(n13498), .C2(n11464), .A(n11463), .B(n11462), .ZN(
        n11465) );
  AOI21_X1 U13903 ( .B1(n14849), .B2(n13501), .A(n11465), .ZN(n11466) );
  OAI21_X1 U13904 ( .B1(n11467), .B2(n13503), .A(n11466), .ZN(P2_U3187) );
  INV_X1 U13905 ( .A(n11656), .ZN(n11470) );
  OAI222_X1 U13906 ( .A1(n14694), .A2(n11657), .B1(n11910), .B2(n11470), .C1(
        n11468), .C2(P1_U3086), .ZN(P1_U3330) );
  OAI222_X1 U13907 ( .A1(n13852), .A2(n11471), .B1(n13854), .B2(n11470), .C1(
        n11469), .C2(P2_U3088), .ZN(P2_U3302) );
  INV_X1 U13908 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11477) );
  AOI211_X1 U13909 ( .C1(n14112), .C2(n14955), .A(n13937), .B(n11472), .ZN(
        n11473) );
  OAI211_X1 U13910 ( .C1(n14670), .C2(n11475), .A(n11474), .B(n11473), .ZN(
        n11478) );
  NAND2_X1 U13911 ( .A1(n11478), .A2(n15202), .ZN(n11476) );
  OAI21_X1 U13912 ( .B1(n15202), .B2(n11477), .A(n11476), .ZN(P1_U3541) );
  INV_X1 U13913 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n11480) );
  NAND2_X1 U13914 ( .A1(n11478), .A2(n15194), .ZN(n11479) );
  OAI21_X1 U13915 ( .B1(n15194), .B2(n11480), .A(n11479), .ZN(P1_U3498) );
  XNOR2_X1 U13916 ( .A(n14938), .B(n14270), .ZN(n14233) );
  XOR2_X1 U13917 ( .A(n14233), .B(n11481), .Z(n11517) );
  OAI211_X1 U13918 ( .C1(n11482), .C2(n11515), .A(n15120), .B(n14739), .ZN(
        n11513) );
  AOI22_X1 U13919 ( .A1(n15129), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n11483), 
        .B2(n15114), .ZN(n11485) );
  NAND2_X1 U13920 ( .A1(n14737), .A2(n14938), .ZN(n11484) );
  OAI211_X1 U13921 ( .C1(n11513), .C2(n14519), .A(n11485), .B(n11484), .ZN(
        n11489) );
  XNOR2_X1 U13922 ( .A(n11486), .B(n14233), .ZN(n11487) );
  AOI222_X1 U13923 ( .A1(n14271), .A2(n14571), .B1(n14269), .B2(n14573), .C1(
        n14971), .C2(n11487), .ZN(n11514) );
  NOR2_X1 U13924 ( .A1(n11514), .A2(n15129), .ZN(n11488) );
  AOI211_X1 U13925 ( .C1(n11517), .C2(n14516), .A(n11489), .B(n11488), .ZN(
        n11490) );
  INV_X1 U13926 ( .A(n11490), .ZN(P1_U3282) );
  INV_X1 U13927 ( .A(n11491), .ZN(n11493) );
  INV_X1 U13928 ( .A(SI_27_), .ZN(n11492) );
  OAI222_X1 U13929 ( .A1(P3_U3151), .A2(n10132), .B1(n14722), .B2(n11493), 
        .C1(n11492), .C2(n14721), .ZN(P3_U3268) );
  OR2_X1 U13930 ( .A1(n11495), .A2(n11494), .ZN(n11496) );
  NOR2_X1 U13931 ( .A1(n14924), .A2(n6646), .ZN(n11498) );
  AOI21_X1 U13932 ( .B1(n14097), .B2(n6638), .A(n11498), .ZN(n12220) );
  NAND2_X1 U13933 ( .A1(n14097), .A2(n6640), .ZN(n11500) );
  NAND2_X1 U13934 ( .A1(n14271), .A2(n6638), .ZN(n11499) );
  NAND2_X1 U13935 ( .A1(n11500), .A2(n11499), .ZN(n11501) );
  XNOR2_X1 U13936 ( .A(n11501), .B(n12341), .ZN(n12222) );
  XOR2_X1 U13937 ( .A(n12220), .B(n12222), .Z(n11503) );
  AOI21_X1 U13938 ( .B1(n11502), .B2(n11503), .A(n14932), .ZN(n11506) );
  NAND2_X2 U13939 ( .A1(n11505), .A2(n11504), .ZN(n14930) );
  NAND2_X1 U13940 ( .A1(n11506), .A2(n14930), .ZN(n11512) );
  NAND2_X1 U13941 ( .A1(n13997), .A2(n14270), .ZN(n11508) );
  OAI211_X1 U13942 ( .C1(n14080), .C2(n14925), .A(n11508), .B(n11507), .ZN(
        n11509) );
  AOI21_X1 U13943 ( .B1(n11510), .B2(n14001), .A(n11509), .ZN(n11511) );
  OAI211_X1 U13944 ( .C1(n15188), .C2(n14005), .A(n11512), .B(n11511), .ZN(
        P1_U3217) );
  OAI211_X1 U13945 ( .C1(n11515), .C2(n15187), .A(n11514), .B(n11513), .ZN(
        n11516) );
  AOI21_X1 U13946 ( .B1(n11517), .B2(n15191), .A(n11516), .ZN(n11520) );
  OR2_X1 U13947 ( .A1(n15202), .A2(n10050), .ZN(n11518) );
  OAI21_X1 U13948 ( .B1(n11520), .B2(n15200), .A(n11518), .ZN(P1_U3539) );
  NAND2_X1 U13949 ( .A1(n15192), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n11519) );
  OAI21_X1 U13950 ( .B1(n11520), .B2(n15192), .A(n11519), .ZN(P1_U3492) );
  XNOR2_X1 U13951 ( .A(n14764), .B(n6823), .ZN(n11612) );
  NAND2_X1 U13952 ( .A1(n11612), .A2(n14778), .ZN(n11524) );
  INV_X1 U13953 ( .A(n11612), .ZN(n11525) );
  NAND2_X1 U13954 ( .A1(n11525), .A2(n12540), .ZN(n11526) );
  XNOR2_X1 U13955 ( .A(n14789), .B(n12416), .ZN(n12356) );
  XNOR2_X1 U13956 ( .A(n12356), .B(n14763), .ZN(n11527) );
  XNOR2_X1 U13957 ( .A(n12355), .B(n11527), .ZN(n11532) );
  NAND2_X1 U13958 ( .A1(n12530), .A2(n12880), .ZN(n11529) );
  AND2_X1 U13959 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n12572) );
  AOI21_X1 U13960 ( .B1(n11608), .B2(n12848), .A(n12572), .ZN(n11528) );
  OAI211_X1 U13961 ( .C1(n14778), .C2(n12527), .A(n11529), .B(n11528), .ZN(
        n11530) );
  AOI21_X1 U13962 ( .B1(n12884), .B2(n12517), .A(n11530), .ZN(n11531) );
  OAI21_X1 U13963 ( .B1(n11532), .B2(n12520), .A(n11531), .ZN(P3_U3155) );
  INV_X1 U13964 ( .A(n13999), .ZN(n14267) );
  NAND2_X1 U13965 ( .A1(n14909), .A2(n14267), .ZN(n11533) );
  NAND2_X1 U13966 ( .A1(n11534), .A2(n14017), .ZN(n11537) );
  INV_X1 U13967 ( .A(n15052), .ZN(n11535) );
  AOI22_X1 U13968 ( .A1(n11700), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n11699), 
        .B2(n11535), .ZN(n11536) );
  NAND2_X1 U13969 ( .A1(n14956), .A2(n14912), .ZN(n14124) );
  NAND2_X1 U13970 ( .A1(n14123), .A2(n14124), .ZN(n14237) );
  OAI21_X1 U13971 ( .B1(n11538), .B2(n14237), .A(n11669), .ZN(n14963) );
  INV_X1 U13972 ( .A(n14963), .ZN(n11557) );
  INV_X1 U13973 ( .A(n14119), .ZN(n11539) );
  AND2_X1 U13974 ( .A1(n11541), .A2(n14237), .ZN(n14959) );
  OR3_X1 U13975 ( .A1(n14960), .A2(n14959), .A3(n14483), .ZN(n11556) );
  NOR2_X1 U13976 ( .A1(n11542), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n11543) );
  OR2_X1 U13977 ( .A1(n11678), .A2(n11543), .ZN(n14923) );
  INV_X1 U13978 ( .A(n14923), .ZN(n11544) );
  NAND2_X1 U13979 ( .A1(n11751), .A2(n11544), .ZN(n11548) );
  NAND2_X1 U13980 ( .A1(n11774), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n11547) );
  NAND2_X1 U13981 ( .A1(n14011), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n11546) );
  NAND2_X1 U13982 ( .A1(n14012), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n11545) );
  NAND4_X1 U13983 ( .A1(n11548), .A2(n11547), .A3(n11546), .A4(n11545), .ZN(
        n14266) );
  INV_X1 U13984 ( .A(n14266), .ZN(n14128) );
  OAI22_X1 U13985 ( .A1(n14128), .A2(n14533), .B1(n13999), .B2(n14531), .ZN(
        n14954) );
  AOI21_X1 U13986 ( .B1(n14002), .B2(n15114), .A(n14954), .ZN(n11550) );
  NAND2_X1 U13987 ( .A1(n15129), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n11549) );
  OAI21_X1 U13988 ( .B1(n11550), .B2(n15129), .A(n11549), .ZN(n11554) );
  AND2_X2 U13989 ( .A1(n11552), .A2(n14006), .ZN(n14577) );
  INV_X1 U13990 ( .A(n14577), .ZN(n11551) );
  OAI21_X1 U13991 ( .B1(n14006), .B2(n11552), .A(n11551), .ZN(n14958) );
  NOR2_X1 U13992 ( .A1(n14958), .A2(n14371), .ZN(n11553) );
  AOI211_X1 U13993 ( .C1(n14737), .C2(n14956), .A(n11554), .B(n11553), .ZN(
        n11555) );
  OAI211_X1 U13994 ( .C1(n11557), .C2(n14584), .A(n11556), .B(n11555), .ZN(
        P1_U3278) );
  INV_X1 U13995 ( .A(n11558), .ZN(n11914) );
  NOR2_X1 U13996 ( .A1(n11913), .A2(n11914), .ZN(n11560) );
  XNOR2_X1 U13997 ( .A(n14830), .B(n6838), .ZN(n11916) );
  NAND2_X1 U13998 ( .A1(n11957), .A2(n13520), .ZN(n11915) );
  INV_X1 U13999 ( .A(n11915), .ZN(n11918) );
  XNOR2_X1 U14000 ( .A(n11916), .B(n11918), .ZN(n11559) );
  XNOR2_X1 U14001 ( .A(n11560), .B(n11559), .ZN(n11564) );
  NOR2_X1 U14002 ( .A1(n13498), .A2(n14826), .ZN(n11562) );
  AOI22_X1 U14003 ( .A1(n13474), .A2(n13519), .B1(n13475), .B2(n13521), .ZN(
        n14821) );
  OAI22_X1 U14004 ( .A1(n13476), .A2(n14821), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8774), .ZN(n11561) );
  AOI211_X1 U14005 ( .C1(n14830), .C2(n13501), .A(n11562), .B(n11561), .ZN(
        n11563) );
  OAI21_X1 U14006 ( .B1(n11564), .B2(n13503), .A(n11563), .ZN(P2_U3213) );
  NAND2_X1 U14007 ( .A1(n14885), .A2(n11567), .ZN(n11565) );
  OR2_X1 U14008 ( .A1(n14885), .A2(n11567), .ZN(n11568) );
  INV_X1 U14009 ( .A(n14838), .ZN(n14848) );
  NAND2_X1 U14010 ( .A1(n14849), .A2(n13521), .ZN(n11569) );
  OR2_X1 U14011 ( .A1(n14830), .A2(n13520), .ZN(n11570) );
  NAND2_X1 U14012 ( .A1(n13750), .A2(n13519), .ZN(n11572) );
  OAI21_X1 U14013 ( .B1(n11573), .B2(n11585), .A(n11833), .ZN(n14857) );
  INV_X1 U14014 ( .A(n11574), .ZN(n11575) );
  OR2_X1 U14015 ( .A1(n14885), .A2(n11577), .ZN(n11578) );
  NOR2_X1 U14016 ( .A1(n14849), .A2(n11579), .ZN(n11580) );
  OR2_X1 U14017 ( .A1(n14830), .A2(n11581), .ZN(n11582) );
  OR2_X1 U14018 ( .A1(n13750), .A2(n11583), .ZN(n11584) );
  XOR2_X1 U14019 ( .A(n11815), .B(n11585), .Z(n11586) );
  AOI22_X1 U14020 ( .A1(n13517), .A2(n13474), .B1(n13475), .B2(n13519), .ZN(
        n13443) );
  OAI21_X1 U14021 ( .B1(n11586), .B2(n14819), .A(n13443), .ZN(n14860) );
  NAND2_X1 U14022 ( .A1(n14860), .A2(n13748), .ZN(n11590) );
  OAI22_X1 U14023 ( .A1(n13748), .A2(n11175), .B1(n13442), .B2(n14827), .ZN(
        n11588) );
  INV_X1 U14024 ( .A(n14830), .ZN(n14874) );
  INV_X1 U14025 ( .A(n11923), .ZN(n14859) );
  OAI211_X1 U14026 ( .C1(n7326), .C2(n14859), .A(n14852), .B(n13729), .ZN(
        n14858) );
  NOR2_X1 U14027 ( .A1(n14858), .A2(n13685), .ZN(n11587) );
  AOI211_X1 U14028 ( .C1(n14844), .C2(n11923), .A(n11588), .B(n11587), .ZN(
        n11589) );
  OAI211_X1 U14029 ( .C1(n13738), .C2(n14857), .A(n11590), .B(n11589), .ZN(
        P2_U3248) );
  NOR2_X1 U14030 ( .A1(n11596), .A2(n11591), .ZN(n11592) );
  NOR2_X1 U14031 ( .A1(n11593), .A2(n11592), .ZN(n11594) );
  XOR2_X1 U14032 ( .A(n11594), .B(P2_REG2_REG_19__SCAN_IN), .Z(n11603) );
  INV_X1 U14033 ( .A(n11603), .ZN(n11601) );
  NAND2_X1 U14034 ( .A1(n11596), .A2(n11595), .ZN(n11597) );
  NAND2_X1 U14035 ( .A1(n11598), .A2(n11597), .ZN(n11599) );
  XOR2_X1 U14036 ( .A(n11599), .B(P2_REG1_REG_19__SCAN_IN), .Z(n11602) );
  OAI21_X1 U14037 ( .B1(n11602), .B2(n15225), .A(n15278), .ZN(n11600) );
  AOI21_X1 U14038 ( .B1(n11601), .B2(n15271), .A(n11600), .ZN(n11605) );
  AOI22_X1 U14039 ( .A1(n11603), .A2(n15271), .B1(n15264), .B2(n11602), .ZN(
        n11604) );
  MUX2_X1 U14040 ( .A(n11605), .B(n11604), .S(n13587), .Z(n11606) );
  NAND2_X1 U14041 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13407)
         );
  OAI211_X1 U14042 ( .C1(n7778), .C2(n15250), .A(n11606), .B(n13407), .ZN(
        P2_U3233) );
  NOR2_X1 U14043 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11607), .ZN(n12556) );
  AOI21_X1 U14044 ( .B1(n11608), .B2(n12539), .A(n12556), .ZN(n11611) );
  NAND2_X1 U14045 ( .A1(n12517), .A2(n11609), .ZN(n11610) );
  OAI211_X1 U14046 ( .C1(n14762), .C2(n12527), .A(n11611), .B(n11610), .ZN(
        n11617) );
  XNOR2_X1 U14047 ( .A(n11612), .B(n12540), .ZN(n11613) );
  XNOR2_X1 U14048 ( .A(n11614), .B(n11613), .ZN(n11615) );
  NOR2_X1 U14049 ( .A1(n11615), .A2(n12520), .ZN(n11616) );
  AOI211_X1 U14050 ( .C1(n14765), .C2(n12530), .A(n11617), .B(n11616), .ZN(
        n11618) );
  INV_X1 U14051 ( .A(n11618), .ZN(P3_U3174) );
  OAI222_X1 U14052 ( .A1(n14694), .A2(n11620), .B1(n11619), .B2(P1_U3086), 
        .C1(n11910), .C2(n9336), .ZN(P1_U3353) );
  INV_X1 U14053 ( .A(n11772), .ZN(n13845) );
  OAI222_X1 U14054 ( .A1(n11910), .A2(n13845), .B1(n11621), .B2(P1_U3086), 
        .C1(n11770), .C2(n14694), .ZN(P1_U3326) );
  AOI21_X1 U14055 ( .B1(n11966), .B2(n13748), .A(n14844), .ZN(n11631) );
  NOR2_X1 U14056 ( .A1(n11622), .A2(n14841), .ZN(n11624) );
  OAI21_X1 U14057 ( .B1(n11624), .B2(n15308), .A(n11623), .ZN(n15310) );
  NOR2_X1 U14058 ( .A1(n11625), .A2(n15308), .ZN(n11629) );
  OAI22_X1 U14059 ( .A1(n13748), .A2(n11627), .B1(n11626), .B2(n14827), .ZN(
        n11628) );
  AOI211_X1 U14060 ( .C1(n13748), .C2(n15310), .A(n11629), .B(n11628), .ZN(
        n11630) );
  OAI21_X1 U14061 ( .B1(n11631), .B2(n15307), .A(n11630), .ZN(P2_U3265) );
  INV_X1 U14062 ( .A(n11642), .ZN(n11912) );
  OAI222_X1 U14063 ( .A1(P2_U3088), .A2(n9193), .B1(n13854), .B2(n11912), .C1(
        n11632), .C2(n13852), .ZN(P2_U3300) );
  NAND2_X1 U14064 ( .A1(n11809), .A2(n14017), .ZN(n11634) );
  OR2_X1 U14065 ( .A1(n6648), .A2(n11810), .ZN(n11633) );
  NAND2_X1 U14066 ( .A1(n11774), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n11641) );
  INV_X1 U14067 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13275) );
  NAND2_X1 U14068 ( .A1(n11678), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n11690) );
  INV_X1 U14069 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n11689) );
  INV_X1 U14070 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n13880) );
  NAND2_X1 U14071 ( .A1(n11726), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n11739) );
  NAND2_X1 U14072 ( .A1(n11727), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n11750) );
  NAND2_X1 U14073 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(n11749), .ZN(n11660) );
  INV_X1 U14074 ( .A(n11660), .ZN(n11635) );
  NAND2_X1 U14075 ( .A1(n11635), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n11763) );
  INV_X1 U14076 ( .A(n11763), .ZN(n11636) );
  NAND2_X1 U14077 ( .A1(n11636), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n11765) );
  INV_X1 U14078 ( .A(n11765), .ZN(n11637) );
  NAND2_X1 U14079 ( .A1(n11637), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n11773) );
  XNOR2_X1 U14080 ( .A(n11773), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n14380) );
  NAND2_X1 U14081 ( .A1(n11751), .A2(n14380), .ZN(n11640) );
  NAND2_X1 U14082 ( .A1(n14011), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n11639) );
  NAND2_X1 U14083 ( .A1(n11775), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n11638) );
  NAND4_X1 U14084 ( .A1(n11641), .A2(n11640), .A3(n11639), .A4(n11638), .ZN(
        n14262) );
  INV_X1 U14085 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n11644) );
  NAND2_X1 U14086 ( .A1(n11765), .A2(n11644), .ZN(n11645) );
  NAND2_X1 U14087 ( .A1(n11751), .A2(n14392), .ZN(n11649) );
  NAND2_X1 U14088 ( .A1(n11774), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n11648) );
  NAND2_X1 U14089 ( .A1(n11715), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n11647) );
  NAND2_X1 U14090 ( .A1(n14011), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n11646) );
  NAND4_X1 U14091 ( .A1(n11649), .A2(n11648), .A3(n11647), .A4(n11646), .ZN(
        n14263) );
  INV_X1 U14092 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n11650) );
  NAND2_X1 U14093 ( .A1(n11660), .A2(n11650), .ZN(n11651) );
  AND2_X1 U14094 ( .A1(n11763), .A2(n11651), .ZN(n14427) );
  NAND2_X1 U14095 ( .A1(n11751), .A2(n14427), .ZN(n11655) );
  NAND2_X1 U14096 ( .A1(n11774), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n11654) );
  NAND2_X1 U14097 ( .A1(n14012), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n11653) );
  NAND2_X1 U14098 ( .A1(n14011), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n11652) );
  NAND4_X1 U14099 ( .A1(n11655), .A2(n11654), .A3(n11653), .A4(n11652), .ZN(
        n14264) );
  NAND2_X1 U14100 ( .A1(n11656), .A2(n14017), .ZN(n11659) );
  OR2_X1 U14101 ( .A1(n6648), .A2(n11657), .ZN(n11658) );
  INV_X1 U14102 ( .A(n14431), .ZN(n14620) );
  OAI21_X1 U14103 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n11749), .A(n11660), 
        .ZN(n13927) );
  INV_X1 U14104 ( .A(n13927), .ZN(n14445) );
  NAND2_X1 U14105 ( .A1(n11751), .A2(n14445), .ZN(n11664) );
  NAND2_X1 U14106 ( .A1(n11774), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n11663) );
  NAND2_X1 U14107 ( .A1(n14012), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n11662) );
  NAND2_X1 U14108 ( .A1(n14011), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n11661) );
  NAND4_X1 U14109 ( .A1(n11664), .A2(n11663), .A3(n11662), .A4(n11661), .ZN(
        n14423) );
  INV_X1 U14110 ( .A(n14423), .ZN(n12305) );
  NAND2_X1 U14111 ( .A1(n11665), .A2(n14017), .ZN(n11667) );
  OR2_X1 U14112 ( .A1(n6648), .A2(n11813), .ZN(n11666) );
  INV_X1 U14113 ( .A(n14626), .ZN(n14448) );
  OR2_X1 U14114 ( .A1(n14956), .A2(n14572), .ZN(n11668) );
  NAND2_X1 U14115 ( .A1(n11670), .A2(n14017), .ZN(n11672) );
  AOI22_X1 U14116 ( .A1(n11700), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n11699), 
        .B2(n15067), .ZN(n11671) );
  XNOR2_X1 U14117 ( .A(n14921), .B(n14128), .ZN(n14238) );
  OR2_X1 U14118 ( .A1(n14921), .A2(n14266), .ZN(n11673) );
  NAND2_X1 U14119 ( .A1(n11674), .A2(n11673), .ZN(n14556) );
  NAND2_X1 U14120 ( .A1(n11675), .A2(n14017), .ZN(n11677) );
  AOI22_X1 U14121 ( .A1(n11700), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n11699), 
        .B2(n14343), .ZN(n11676) );
  OR2_X1 U14122 ( .A1(n11678), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n11679) );
  AND2_X1 U14123 ( .A1(n11690), .A2(n11679), .ZN(n14562) );
  NAND2_X1 U14124 ( .A1(n11751), .A2(n14562), .ZN(n11683) );
  NAND2_X1 U14125 ( .A1(n11774), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n11682) );
  NAND2_X1 U14126 ( .A1(n11775), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n11681) );
  NAND2_X1 U14127 ( .A1(n14011), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n11680) );
  NAND4_X1 U14128 ( .A1(n11683), .A2(n11682), .A3(n11681), .A4(n11680), .ZN(
        n14574) );
  NAND2_X1 U14129 ( .A1(n14565), .A2(n14574), .ZN(n11684) );
  NAND2_X1 U14130 ( .A1(n11685), .A2(n14017), .ZN(n11688) );
  INV_X1 U14131 ( .A(n15099), .ZN(n11686) );
  AOI22_X1 U14132 ( .A1(n11700), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n11699), 
        .B2(n11686), .ZN(n11687) );
  NAND2_X1 U14133 ( .A1(n11774), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n11695) );
  NAND2_X1 U14134 ( .A1(n11690), .A2(n11689), .ZN(n11691) );
  AND2_X1 U14135 ( .A1(n11703), .A2(n11691), .ZN(n14549) );
  NAND2_X1 U14136 ( .A1(n11751), .A2(n14549), .ZN(n11694) );
  NAND2_X1 U14137 ( .A1(n14011), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n11693) );
  NAND2_X1 U14138 ( .A1(n14012), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n11692) );
  AND2_X1 U14139 ( .A1(n14667), .A2(n14265), .ZN(n11696) );
  OR2_X1 U14140 ( .A1(n14667), .A2(n14265), .ZN(n11697) );
  NAND2_X1 U14141 ( .A1(n11698), .A2(n14017), .ZN(n11702) );
  AOI22_X1 U14142 ( .A1(n11700), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14579), 
        .B2(n11699), .ZN(n11701) );
  NAND2_X1 U14143 ( .A1(n11703), .A2(n13880), .ZN(n11704) );
  NAND2_X1 U14144 ( .A1(n11714), .A2(n11704), .ZN(n14537) );
  INV_X1 U14145 ( .A(n14537), .ZN(n13883) );
  NAND2_X1 U14146 ( .A1(n11751), .A2(n13883), .ZN(n11708) );
  NAND2_X1 U14147 ( .A1(n11774), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n11707) );
  NAND2_X1 U14148 ( .A1(n14012), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n11706) );
  NAND2_X1 U14149 ( .A1(n14011), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n11705) );
  NAND4_X1 U14150 ( .A1(n11708), .A2(n11707), .A3(n11706), .A4(n11705), .ZN(
        n14545) );
  XNOR2_X1 U14151 ( .A(n14662), .B(n14545), .ZN(n14524) );
  INV_X1 U14152 ( .A(n14524), .ZN(n14528) );
  OR2_X1 U14153 ( .A1(n14662), .A2(n14545), .ZN(n11709) );
  NAND2_X1 U14154 ( .A1(n11710), .A2(n11709), .ZN(n14514) );
  INV_X1 U14155 ( .A(n14514), .ZN(n11721) );
  NAND2_X1 U14156 ( .A1(n11711), .A2(n14017), .ZN(n11713) );
  OR2_X1 U14157 ( .A1(n6649), .A2(n13291), .ZN(n11712) );
  AOI21_X1 U14158 ( .B1(n11714), .B2(n13275), .A(n11726), .ZN(n14509) );
  NAND2_X1 U14159 ( .A1(n11751), .A2(n14509), .ZN(n11719) );
  NAND2_X1 U14160 ( .A1(n11774), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n11718) );
  NAND2_X1 U14161 ( .A1(n11715), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n11717) );
  NAND2_X1 U14162 ( .A1(n14011), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n11716) );
  XNOR2_X1 U14163 ( .A(n14652), .B(n14498), .ZN(n14515) );
  OR2_X1 U14164 ( .A1(n14518), .A2(n14532), .ZN(n11722) );
  OR2_X1 U14165 ( .A1(n6648), .A2(n11724), .ZN(n11725) );
  INV_X1 U14166 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n11729) );
  INV_X1 U14167 ( .A(n11726), .ZN(n11728) );
  AOI21_X1 U14168 ( .B1(n11729), .B2(n11728), .A(n11727), .ZN(n14491) );
  NAND2_X1 U14169 ( .A1(n11751), .A2(n14491), .ZN(n11733) );
  NAND2_X1 U14170 ( .A1(n11774), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n11732) );
  NAND2_X1 U14171 ( .A1(n14012), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n11731) );
  NAND2_X1 U14172 ( .A1(n14011), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n11730) );
  NAND4_X1 U14173 ( .A1(n11733), .A2(n11732), .A3(n11731), .A4(n11730), .ZN(
        n14506) );
  INV_X1 U14174 ( .A(n14506), .ZN(n13954) );
  OR2_X1 U14175 ( .A1(n11735), .A2(n6832), .ZN(n11736) );
  XNOR2_X1 U14176 ( .A(n11736), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14698) );
  INV_X1 U14177 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13955) );
  AOI21_X1 U14178 ( .B1(n13955), .B2(n11739), .A(n11738), .ZN(n14473) );
  NAND2_X1 U14179 ( .A1(n11751), .A2(n14473), .ZN(n11743) );
  NAND2_X1 U14180 ( .A1(n11774), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n11742) );
  NAND2_X1 U14181 ( .A1(n11775), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n11741) );
  NAND2_X1 U14182 ( .A1(n14011), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n11740) );
  NAND4_X1 U14183 ( .A1(n11743), .A2(n11742), .A3(n11741), .A4(n11740), .ZN(
        n14497) );
  XNOR2_X1 U14184 ( .A(n13961), .B(n14497), .ZN(n14469) );
  OR2_X1 U14185 ( .A1(n14639), .A2(n14497), .ZN(n11744) );
  NAND2_X1 U14186 ( .A1(n11745), .A2(n14017), .ZN(n11748) );
  OR2_X1 U14187 ( .A1(n6649), .A2(n11746), .ZN(n11747) );
  INV_X1 U14188 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n13872) );
  AOI21_X1 U14189 ( .B1(n13872), .B2(n11750), .A(n11749), .ZN(n14459) );
  NAND2_X1 U14190 ( .A1(n11751), .A2(n14459), .ZN(n11755) );
  NAND2_X1 U14191 ( .A1(n11774), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n11754) );
  NAND2_X1 U14192 ( .A1(n14012), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n11753) );
  NAND2_X1 U14193 ( .A1(n14011), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n11752) );
  NAND4_X1 U14194 ( .A1(n11755), .A2(n11754), .A3(n11753), .A4(n11752), .ZN(
        n14470) );
  NOR2_X1 U14195 ( .A1(n14633), .A2(n14470), .ZN(n11757) );
  NAND2_X1 U14196 ( .A1(n14633), .A2(n14470), .ZN(n11756) );
  XNOR2_X1 U14197 ( .A(n14626), .B(n14423), .ZN(n14440) );
  NAND2_X1 U14198 ( .A1(n14431), .A2(n13986), .ZN(n11785) );
  OR2_X1 U14199 ( .A1(n14431), .A2(n13986), .ZN(n11758) );
  OAI21_X1 U14200 ( .B1(n13986), .B2(n14620), .A(n14415), .ZN(n14411) );
  NAND2_X1 U14201 ( .A1(n13851), .A2(n14017), .ZN(n11761) );
  OR2_X1 U14202 ( .A1(n6649), .A2(n14695), .ZN(n11760) );
  INV_X1 U14203 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n11762) );
  NAND2_X1 U14204 ( .A1(n11763), .A2(n11762), .ZN(n11764) );
  AND2_X1 U14205 ( .A1(n11765), .A2(n11764), .ZN(n14407) );
  NAND2_X1 U14206 ( .A1(n11751), .A2(n14407), .ZN(n11769) );
  NAND2_X1 U14207 ( .A1(n11774), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n11768) );
  NAND2_X1 U14208 ( .A1(n14012), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n11767) );
  NAND2_X1 U14209 ( .A1(n14011), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n11766) );
  NAND4_X1 U14210 ( .A1(n11769), .A2(n11768), .A3(n11767), .A4(n11766), .ZN(
        n14424) );
  NAND2_X1 U14211 ( .A1(n14399), .A2(n14398), .ZN(n14397) );
  OAI21_X1 U14212 ( .B1(n14608), .B2(n14263), .A(n14397), .ZN(n14375) );
  XNOR2_X1 U14213 ( .A(n14384), .B(n12339), .ZN(n14373) );
  INV_X1 U14214 ( .A(n14373), .ZN(n14376) );
  NOR2_X1 U14215 ( .A1(n6649), .A2(n11770), .ZN(n11771) );
  INV_X1 U14216 ( .A(n14593), .ZN(n11796) );
  INV_X1 U14217 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n12349) );
  NOR2_X1 U14218 ( .A1(n11773), .A2(n12349), .ZN(n11801) );
  NAND2_X1 U14219 ( .A1(n11751), .A2(n11801), .ZN(n11779) );
  NAND2_X1 U14220 ( .A1(n11774), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n11778) );
  NAND2_X1 U14221 ( .A1(n11775), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n11777) );
  NAND2_X1 U14222 ( .A1(n14011), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n11776) );
  AND4_X1 U14223 ( .A1(n11779), .A2(n11778), .A3(n11777), .A4(n11776), .ZN(
        n14191) );
  INV_X1 U14224 ( .A(n14191), .ZN(n14261) );
  XNOR2_X1 U14225 ( .A(n11796), .B(n14261), .ZN(n14245) );
  INV_X1 U14226 ( .A(n14123), .ZN(n11780) );
  INV_X1 U14227 ( .A(n14238), .ZN(n14570) );
  XOR2_X1 U14228 ( .A(n14574), .B(n14565), .Z(n14557) );
  INV_X1 U14229 ( .A(n14574), .ZN(n14913) );
  NAND2_X1 U14230 ( .A1(n14667), .A2(n14530), .ZN(n14148) );
  NAND2_X1 U14231 ( .A1(n14147), .A2(n14148), .ZN(n14541) );
  NAND2_X1 U14232 ( .A1(n14496), .A2(n14495), .ZN(n14494) );
  NAND2_X1 U14233 ( .A1(n14494), .A2(n11783), .ZN(n14468) );
  XNOR2_X1 U14234 ( .A(n14633), .B(n14470), .ZN(n14455) );
  INV_X1 U14235 ( .A(n14470), .ZN(n13956) );
  NAND2_X1 U14236 ( .A1(n14633), .A2(n13956), .ZN(n11784) );
  INV_X1 U14237 ( .A(n14440), .ZN(n14435) );
  INV_X1 U14238 ( .A(n14398), .ZN(n11786) );
  NAND2_X1 U14239 ( .A1(n14389), .A2(n11786), .ZN(n11788) );
  NAND2_X1 U14240 ( .A1(n14608), .A2(n13985), .ZN(n11787) );
  NOR2_X1 U14241 ( .A1(n14600), .A2(n14262), .ZN(n11789) );
  XNOR2_X1 U14242 ( .A(n11790), .B(n6960), .ZN(n11792) );
  INV_X1 U14243 ( .A(n14597), .ZN(n11794) );
  NAND2_X1 U14244 ( .A1(n14262), .A2(n14571), .ZN(n14591) );
  INV_X1 U14245 ( .A(n14591), .ZN(n11793) );
  OR2_X2 U14246 ( .A1(n14517), .A2(n14644), .ZN(n14489) );
  INV_X1 U14247 ( .A(n14379), .ZN(n11795) );
  AOI21_X1 U14248 ( .B1(n11796), .B2(n11795), .A(n14365), .ZN(n14595) );
  AOI21_X1 U14249 ( .B1(n11797), .B2(P1_B_REG_SCAN_IN), .A(n14533), .ZN(n14360) );
  INV_X1 U14250 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n14367) );
  NAND2_X1 U14251 ( .A1(n11774), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n11799) );
  NAND2_X1 U14252 ( .A1(n14012), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n11798) );
  OAI211_X1 U14253 ( .C1(n11800), .C2(n14367), .A(n11799), .B(n11798), .ZN(
        n14260) );
  NAND2_X1 U14254 ( .A1(n14360), .A2(n14260), .ZN(n14592) );
  INV_X1 U14255 ( .A(n11801), .ZN(n11802) );
  OAI22_X1 U14256 ( .A1(n11803), .A2(n14592), .B1(n11802), .B2(n14578), .ZN(
        n11804) );
  AOI21_X1 U14257 ( .B1(P1_REG2_REG_29__SCAN_IN), .B2(n15129), .A(n11804), 
        .ZN(n11805) );
  OAI21_X1 U14258 ( .B1(n14593), .B2(n15116), .A(n11805), .ZN(n11806) );
  AOI21_X1 U14259 ( .B1(n14595), .B2(n14503), .A(n11806), .ZN(n11807) );
  OAI211_X1 U14260 ( .C1(n14598), .C2(n14584), .A(n11808), .B(n11807), .ZN(
        P1_U3356) );
  INV_X1 U14261 ( .A(n11809), .ZN(n13850) );
  OAI222_X1 U14262 ( .A1(n14694), .A2(n11810), .B1(n11910), .B2(n13850), .C1(
        P1_U3086), .C2(n9266), .ZN(P1_U3327) );
  OAI222_X1 U14263 ( .A1(n14694), .A2(n11813), .B1(n11910), .B2(n11812), .C1(
        n11811), .C2(P1_U3086), .ZN(P1_U3331) );
  INV_X1 U14264 ( .A(n13513), .ZN(n13399) );
  INV_X1 U14265 ( .A(n13514), .ZN(n11822) );
  NAND2_X1 U14266 ( .A1(n11923), .A2(n13484), .ZN(n11814) );
  OR2_X1 U14267 ( .A1(n11923), .A2(n13484), .ZN(n11816) );
  INV_X1 U14268 ( .A(n13517), .ZN(n11817) );
  NOR2_X1 U14269 ( .A1(n13822), .A2(n11817), .ZN(n11818) );
  INV_X1 U14270 ( .A(n13516), .ZN(n13485) );
  AND2_X1 U14271 ( .A1(n13818), .A2(n13485), .ZN(n11819) );
  OR2_X1 U14272 ( .A1(n13818), .A2(n13485), .ZN(n11820) );
  NAND2_X1 U14273 ( .A1(n13697), .A2(n11821), .ZN(n13687) );
  INV_X1 U14274 ( .A(n13790), .ZN(n13644) );
  INV_X1 U14275 ( .A(n13610), .ZN(n13606) );
  INV_X1 U14276 ( .A(n13779), .ZN(n13617) );
  OAI22_X1 U14277 ( .A1(n13607), .A2(n13606), .B1(n13617), .B2(n13509), .ZN(
        n13593) );
  INV_X1 U14278 ( .A(n13602), .ZN(n13592) );
  NAND2_X1 U14279 ( .A1(n13507), .A2(n13475), .ZN(n11829) );
  INV_X1 U14280 ( .A(P2_B_REG_SCAN_IN), .ZN(n11825) );
  NOR2_X1 U14281 ( .A1(n9193), .A2(n11825), .ZN(n11826) );
  NOR2_X1 U14282 ( .A1(n13492), .A2(n11826), .ZN(n13565) );
  INV_X1 U14283 ( .A(n11827), .ZN(n13505) );
  NAND2_X1 U14284 ( .A1(n13565), .A2(n13505), .ZN(n11828) );
  NAND2_X1 U14285 ( .A1(n11923), .A2(n13518), .ZN(n11832) );
  OR2_X1 U14286 ( .A1(n13822), .A2(n13517), .ZN(n11834) );
  NAND2_X1 U14287 ( .A1(n13711), .A2(n11835), .ZN(n11837) );
  NAND2_X1 U14288 ( .A1(n11837), .A2(n11836), .ZN(n13696) );
  NAND2_X1 U14289 ( .A1(n13813), .A2(n13515), .ZN(n11838) );
  OR2_X1 U14290 ( .A1(n13813), .A2(n13515), .ZN(n11839) );
  NOR2_X1 U14291 ( .A1(n13804), .A2(n13514), .ZN(n11840) );
  INV_X1 U14292 ( .A(n13663), .ZN(n13672) );
  INV_X1 U14293 ( .A(n13621), .ZN(n13626) );
  NAND2_X1 U14294 ( .A1(n13627), .A2(n13626), .ZN(n13625) );
  NAND2_X1 U14295 ( .A1(n13779), .A2(n13509), .ZN(n11843) );
  INV_X1 U14296 ( .A(n11844), .ZN(n13579) );
  NAND2_X1 U14297 ( .A1(n13578), .A2(n13579), .ZN(n13577) );
  INV_X1 U14298 ( .A(n13765), .ZN(n11852) );
  INV_X1 U14299 ( .A(n13785), .ZN(n13634) );
  INV_X1 U14300 ( .A(n13818), .ZN(n13721) );
  NOR2_X1 U14301 ( .A1(n13822), .A2(n13729), .ZN(n13727) );
  NAND2_X1 U14302 ( .A1(n13721), .A2(n13727), .ZN(n13717) );
  NAND2_X1 U14303 ( .A1(n13634), .A2(n13641), .ZN(n13628) );
  AOI21_X1 U14304 ( .B1(n13762), .B2(n13584), .A(n13728), .ZN(n11847) );
  AND2_X1 U14305 ( .A1(n11847), .A2(n13570), .ZN(n13761) );
  NAND2_X1 U14306 ( .A1(n13761), .A2(n15285), .ZN(n11850) );
  AOI22_X1 U14307 ( .A1(n15292), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n11848), 
        .B2(n15279), .ZN(n11849) );
  OAI211_X1 U14308 ( .C1(n7320), .C2(n15282), .A(n11850), .B(n11849), .ZN(
        n11851) );
  AOI21_X1 U14309 ( .B1(n11852), .B2(n15288), .A(n11851), .ZN(n11853) );
  OAI21_X1 U14310 ( .B1(n13764), .B2(n15292), .A(n11853), .ZN(P2_U3236) );
  NAND2_X1 U14311 ( .A1(n12578), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n11874) );
  NOR2_X1 U14312 ( .A1(n12564), .A2(n11855), .ZN(n11856) );
  INV_X1 U14313 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n14798) );
  OR2_X1 U14314 ( .A1(n12578), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n11857) );
  NAND2_X1 U14315 ( .A1(n11874), .A2(n11857), .ZN(n12568) );
  AND2_X1 U14316 ( .A1(n11896), .A2(n11858), .ZN(n11859) );
  INV_X1 U14317 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12955) );
  NAND2_X1 U14318 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n11899), .ZN(n11860) );
  OAI21_X1 U14319 ( .B1(P3_REG1_REG_16__SCAN_IN), .B2(n11899), .A(n11860), 
        .ZN(n12602) );
  NOR2_X1 U14320 ( .A1(n12633), .A2(n11861), .ZN(n11862) );
  INV_X1 U14321 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12945) );
  INV_X1 U14322 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12941) );
  AOI22_X1 U14323 ( .A1(P3_REG1_REG_18__SCAN_IN), .A2(n11887), .B1(n12644), 
        .B2(n12941), .ZN(n12637) );
  XNOR2_X1 U14324 ( .A(n12014), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n11864) );
  INV_X1 U14325 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n11863) );
  MUX2_X1 U14326 ( .A(P3_REG2_REG_19__SCAN_IN), .B(n11863), .S(n12014), .Z(
        n11905) );
  MUX2_X1 U14327 ( .A(n11905), .B(n7352), .S(n6642), .Z(n11889) );
  INV_X1 U14328 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n11901) );
  MUX2_X1 U14329 ( .A(n11901), .B(n12945), .S(n6642), .Z(n11882) );
  NOR2_X1 U14330 ( .A1(n12633), .A2(n11882), .ZN(n11884) );
  MUX2_X1 U14331 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n6642), .Z(n11865) );
  AND2_X1 U14332 ( .A1(n11899), .A2(n11865), .ZN(n12604) );
  NAND2_X1 U14333 ( .A1(n12578), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n11895) );
  OR2_X1 U14334 ( .A1(n12578), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n11866) );
  NAND2_X1 U14335 ( .A1(n11895), .A2(n11866), .ZN(n12570) );
  MUX2_X1 U14336 ( .A(n12568), .B(n12570), .S(n12187), .Z(n11867) );
  INV_X1 U14337 ( .A(n11867), .ZN(n12574) );
  INV_X1 U14338 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n11868) );
  MUX2_X1 U14339 ( .A(n11868), .B(n14798), .S(n6642), .Z(n11873) );
  XNOR2_X1 U14340 ( .A(n11873), .B(n12564), .ZN(n12555) );
  NAND2_X1 U14341 ( .A1(n11869), .A2(n11892), .ZN(n11872) );
  NOR2_X1 U14342 ( .A1(n12555), .A2(n12554), .ZN(n12553) );
  AOI21_X1 U14343 ( .B1(n11873), .B2(n12564), .A(n12553), .ZN(n12575) );
  NAND2_X1 U14344 ( .A1(n12574), .A2(n12575), .ZN(n12573) );
  MUX2_X1 U14345 ( .A(n11874), .B(n11895), .S(n12187), .Z(n11875) );
  NAND2_X1 U14346 ( .A1(n12573), .A2(n11875), .ZN(n11876) );
  NOR2_X1 U14347 ( .A1(n11876), .A2(n11896), .ZN(n11878) );
  AND2_X1 U14348 ( .A1(n11876), .A2(n11896), .ZN(n11877) );
  MUX2_X1 U14349 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n6642), .Z(n12593) );
  NOR2_X1 U14350 ( .A1(n11878), .A2(n12591), .ZN(n12608) );
  INV_X1 U14351 ( .A(n11899), .ZN(n12609) );
  INV_X1 U14352 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n11880) );
  INV_X1 U14353 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n11879) );
  MUX2_X1 U14354 ( .A(n11880), .B(n11879), .S(n6642), .Z(n11881) );
  NAND2_X1 U14355 ( .A1(n12609), .A2(n11881), .ZN(n12606) );
  OAI21_X1 U14356 ( .B1(n12604), .B2(n12608), .A(n12606), .ZN(n12630) );
  AOI21_X1 U14357 ( .B1(n12633), .B2(n11882), .A(n11884), .ZN(n11883) );
  INV_X1 U14358 ( .A(n11883), .ZN(n12629) );
  NOR2_X1 U14359 ( .A1(n12630), .A2(n12629), .ZN(n12628) );
  INV_X1 U14360 ( .A(n11886), .ZN(n11885) );
  XNOR2_X1 U14361 ( .A(n11887), .B(n11885), .ZN(n12641) );
  MUX2_X1 U14362 ( .A(n7435), .B(n12941), .S(n6642), .Z(n12640) );
  NAND2_X1 U14363 ( .A1(n12641), .A2(n12640), .ZN(n12639) );
  NAND2_X1 U14364 ( .A1(n11887), .A2(n11886), .ZN(n11888) );
  NOR2_X1 U14365 ( .A1(n12645), .A2(n12039), .ZN(n11906) );
  XOR2_X1 U14366 ( .A(n11894), .B(n11893), .Z(n12560) );
  INV_X1 U14367 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12585) );
  NAND2_X1 U14368 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n11899), .ZN(n11898) );
  OAI21_X1 U14369 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n11899), .A(n11898), 
        .ZN(n12613) );
  NOR2_X1 U14370 ( .A1(n12633), .A2(n11902), .ZN(n11903) );
  NAND2_X1 U14371 ( .A1(P3_REG2_REG_18__SCAN_IN), .A2(n12644), .ZN(n11904) );
  OAI21_X1 U14372 ( .B1(P3_REG2_REG_18__SCAN_IN), .B2(n12644), .A(n11904), 
        .ZN(n12647) );
  NAND2_X1 U14373 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12409)
         );
  OAI222_X1 U14374 ( .A1(n13852), .A2(n11984), .B1(n13854), .B2(n14026), .C1(
        n11908), .C2(P2_U3088), .ZN(P2_U3297) );
  INV_X1 U14375 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14027) );
  OAI222_X1 U14376 ( .A1(n11910), .A2(n14026), .B1(n11909), .B2(P1_U3086), 
        .C1(n14027), .C2(n14694), .ZN(P1_U3325) );
  OAI222_X1 U14377 ( .A1(n11910), .A2(n11912), .B1(n14254), .B2(P1_U3086), 
        .C1(n11911), .C2(n14694), .ZN(P1_U3328) );
  INV_X1 U14378 ( .A(n11916), .ZN(n11917) );
  AND2_X1 U14379 ( .A1(n11957), .A2(n13519), .ZN(n11920) );
  XNOR2_X1 U14380 ( .A(n13750), .B(n11961), .ZN(n11919) );
  NOR2_X1 U14381 ( .A1(n11919), .A2(n11920), .ZN(n11921) );
  AOI21_X1 U14382 ( .B1(n11920), .B2(n11919), .A(n11921), .ZN(n13431) );
  INV_X1 U14383 ( .A(n11921), .ZN(n11922) );
  AND2_X1 U14384 ( .A1(n11957), .A2(n13518), .ZN(n11925) );
  XNOR2_X1 U14385 ( .A(n11923), .B(n11961), .ZN(n11924) );
  NOR2_X1 U14386 ( .A1(n11924), .A2(n11925), .ZN(n11926) );
  AOI21_X1 U14387 ( .B1(n11925), .B2(n11924), .A(n11926), .ZN(n13440) );
  INV_X1 U14388 ( .A(n11926), .ZN(n11927) );
  NAND2_X1 U14389 ( .A1(n13517), .A2(n11957), .ZN(n11929) );
  XNOR2_X1 U14390 ( .A(n13822), .B(n11961), .ZN(n11928) );
  XOR2_X1 U14391 ( .A(n11929), .B(n11928), .Z(n13482) );
  XNOR2_X1 U14392 ( .A(n13818), .B(n6838), .ZN(n11931) );
  NAND2_X1 U14393 ( .A1(n13516), .A2(n11957), .ZN(n11930) );
  NOR2_X1 U14394 ( .A1(n11931), .A2(n11930), .ZN(n13404) );
  XNOR2_X1 U14395 ( .A(n13813), .B(n6838), .ZN(n11935) );
  INV_X1 U14396 ( .A(n11935), .ZN(n11933) );
  NAND2_X1 U14397 ( .A1(n13515), .A2(n11957), .ZN(n11934) );
  INV_X1 U14398 ( .A(n11934), .ZN(n11932) );
  NAND2_X1 U14399 ( .A1(n11933), .A2(n11932), .ZN(n13463) );
  AND2_X1 U14400 ( .A1(n11935), .A2(n11934), .ZN(n13462) );
  XNOR2_X1 U14401 ( .A(n13804), .B(n11961), .ZN(n11936) );
  NAND2_X1 U14402 ( .A1(n13514), .A2(n11957), .ZN(n11937) );
  XNOR2_X1 U14403 ( .A(n11936), .B(n11937), .ZN(n13412) );
  INV_X1 U14404 ( .A(n11936), .ZN(n11938) );
  NOR2_X1 U14405 ( .A1(n11938), .A2(n11937), .ZN(n11939) );
  XNOR2_X1 U14406 ( .A(n13800), .B(n11961), .ZN(n11940) );
  NOR2_X1 U14407 ( .A1(n13399), .A2(n11966), .ZN(n13472) );
  NAND2_X1 U14408 ( .A1(n13473), .A2(n13472), .ZN(n11944) );
  INV_X1 U14409 ( .A(n11940), .ZN(n11941) );
  OR2_X1 U14410 ( .A1(n11942), .A2(n11941), .ZN(n11943) );
  INV_X1 U14411 ( .A(n11948), .ZN(n11946) );
  XNOR2_X1 U14412 ( .A(n13795), .B(n11961), .ZN(n11947) );
  INV_X1 U14413 ( .A(n11947), .ZN(n11945) );
  NAND2_X1 U14414 ( .A1(n11948), .A2(n11947), .ZN(n11949) );
  NAND2_X1 U14415 ( .A1(n11957), .A2(n13512), .ZN(n13395) );
  XNOR2_X1 U14416 ( .A(n13790), .B(n11961), .ZN(n11950) );
  NAND2_X1 U14417 ( .A1(n9669), .A2(n13511), .ZN(n11951) );
  XNOR2_X1 U14418 ( .A(n11950), .B(n11951), .ZN(n13450) );
  INV_X1 U14419 ( .A(n11950), .ZN(n11952) );
  NAND2_X1 U14420 ( .A1(n11952), .A2(n11951), .ZN(n11953) );
  XNOR2_X1 U14421 ( .A(n13785), .B(n11961), .ZN(n11955) );
  NOR2_X1 U14422 ( .A1(n11966), .A2(n13494), .ZN(n11954) );
  XNOR2_X1 U14423 ( .A(n11955), .B(n11954), .ZN(n13419) );
  NAND2_X1 U14424 ( .A1(n11955), .A2(n11954), .ZN(n11956) );
  XNOR2_X1 U14425 ( .A(n13779), .B(n6838), .ZN(n11959) );
  NAND2_X1 U14426 ( .A1(n11957), .A2(n13509), .ZN(n11958) );
  NAND2_X1 U14427 ( .A1(n11959), .A2(n11958), .ZN(n11960) );
  OAI21_X1 U14428 ( .B1(n11959), .B2(n11958), .A(n11960), .ZN(n13490) );
  XNOR2_X1 U14429 ( .A(n13773), .B(n11961), .ZN(n11962) );
  NOR2_X1 U14430 ( .A1(n11966), .A2(n13493), .ZN(n11963) );
  XNOR2_X1 U14431 ( .A(n11962), .B(n11963), .ZN(n13385) );
  INV_X1 U14432 ( .A(n11962), .ZN(n11965) );
  INV_X1 U14433 ( .A(n11963), .ZN(n11964) );
  NOR2_X1 U14434 ( .A1(n11966), .A2(n13387), .ZN(n11967) );
  XOR2_X1 U14435 ( .A(n11968), .B(n11967), .Z(n11969) );
  XNOR2_X1 U14436 ( .A(n13767), .B(n11969), .ZN(n11970) );
  XNOR2_X1 U14437 ( .A(n11971), .B(n11970), .ZN(n11977) );
  INV_X1 U14438 ( .A(n13586), .ZN(n11974) );
  INV_X1 U14439 ( .A(n13475), .ZN(n13495) );
  OAI22_X1 U14440 ( .A1(n13495), .A2(n13493), .B1(n11972), .B2(n13492), .ZN(
        n13581) );
  AOI22_X1 U14441 ( .A1(n13496), .A2(n13581), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11973) );
  OAI21_X1 U14442 ( .B1(n11974), .B2(n13498), .A(n11973), .ZN(n11975) );
  AOI21_X1 U14443 ( .B1(n13767), .B2(n13501), .A(n11975), .ZN(n11976) );
  OAI21_X1 U14444 ( .B1(n11977), .B2(n13503), .A(n11976), .ZN(P2_U3192) );
  INV_X1 U14445 ( .A(n11978), .ZN(n11980) );
  OAI222_X1 U14446 ( .A1(n14722), .A2(n11980), .B1(n14721), .B2(n11979), .C1(
        P3_U3151), .C2(n8201), .ZN(P3_U3267) );
  INV_X1 U14447 ( .A(n11981), .ZN(n11982) );
  NAND2_X1 U14448 ( .A1(n11984), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n11994) );
  NAND2_X1 U14449 ( .A1(n14027), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n11985) );
  NAND2_X1 U14450 ( .A1(n11994), .A2(n11985), .ZN(n11986) );
  NAND2_X1 U14451 ( .A1(n11987), .A2(n11986), .ZN(n11988) );
  INV_X1 U14452 ( .A(n11990), .ZN(n11989) );
  INV_X1 U14453 ( .A(SI_30_), .ZN(n11991) );
  OAI222_X1 U14454 ( .A1(P3_U3151), .A2(n7702), .B1(n14722), .B2(n11989), .C1(
        n11991), .C2(n14721), .ZN(P3_U3265) );
  NAND2_X1 U14455 ( .A1(n11990), .A2(n11998), .ZN(n11993) );
  OR2_X1 U14456 ( .A1(n11999), .A2(n11991), .ZN(n11992) );
  NAND2_X1 U14457 ( .A1(n11993), .A2(n11992), .ZN(n12008) );
  INV_X1 U14458 ( .A(n12007), .ZN(n12535) );
  AND2_X1 U14459 ( .A1(n14787), .A2(n12535), .ZN(n12015) );
  NAND2_X1 U14460 ( .A1(n11995), .A2(n11994), .ZN(n11997) );
  XNOR2_X1 U14461 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n11996) );
  INV_X1 U14462 ( .A(SI_31_), .ZN(n13020) );
  OR2_X1 U14463 ( .A1(n11999), .A2(n13020), .ZN(n12000) );
  NAND2_X1 U14464 ( .A1(n7929), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12005) );
  NAND2_X1 U14465 ( .A1(n12001), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12004) );
  NAND2_X1 U14466 ( .A1(n12002), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12003) );
  INV_X1 U14467 ( .A(n12656), .ZN(n12534) );
  NOR2_X1 U14468 ( .A1(n12960), .A2(n12534), .ZN(n12179) );
  NAND2_X1 U14469 ( .A1(n12008), .A2(n12007), .ZN(n12009) );
  NAND2_X1 U14470 ( .A1(n12010), .A2(n12009), .ZN(n12178) );
  OAI21_X1 U14471 ( .B1(n14787), .B2(n12534), .A(n12174), .ZN(n12011) );
  INV_X1 U14472 ( .A(n12015), .ZN(n12175) );
  NAND2_X1 U14473 ( .A1(n12162), .A2(n12163), .ZN(n12697) );
  INV_X1 U14474 ( .A(n12804), .ZN(n12033) );
  NOR2_X1 U14475 ( .A1(n10025), .A2(n12017), .ZN(n12047) );
  NAND4_X1 U14476 ( .A1(n12047), .A2(n12020), .A3(n12019), .A4(n12018), .ZN(
        n12028) );
  NOR2_X1 U14477 ( .A1(n12022), .A2(n12021), .ZN(n12026) );
  NAND4_X1 U14478 ( .A1(n12026), .A2(n12025), .A3(n12024), .A4(n12023), .ZN(
        n12027) );
  OR2_X1 U14479 ( .A1(n12028), .A2(n12027), .ZN(n12030) );
  NAND3_X1 U14480 ( .A1(n14768), .A2(n15446), .A3(n12088), .ZN(n12029) );
  NOR4_X1 U14481 ( .A1(n12030), .A2(n12029), .A3(n12097), .A4(n14759), .ZN(
        n12031) );
  AND4_X1 U14482 ( .A1(n12852), .A2(n8216), .A3(n12863), .A4(n12031), .ZN(
        n12032) );
  NAND4_X1 U14483 ( .A1(n12033), .A2(n12814), .A3(n6644), .A4(n12032), .ZN(
        n12034) );
  NOR2_X1 U14484 ( .A1(n12697), .A2(n12036), .ZN(n12037) );
  XNOR2_X1 U14485 ( .A(n12040), .B(n12039), .ZN(n12185) );
  INV_X1 U14486 ( .A(n12749), .ZN(n12982) );
  INV_X1 U14487 ( .A(n12042), .ZN(n12124) );
  AND2_X1 U14488 ( .A1(n12042), .A2(n12041), .ZN(n12119) );
  INV_X1 U14489 ( .A(n12043), .ZN(n12062) );
  INV_X1 U14490 ( .A(n14725), .ZN(n12189) );
  NAND3_X1 U14491 ( .A1(n15463), .A2(n12201), .A3(n14725), .ZN(n12045) );
  NAND2_X1 U14492 ( .A1(n12045), .A2(n12044), .ZN(n12046) );
  AOI22_X1 U14493 ( .A1(n12047), .A2(n12189), .B1(n12050), .B2(n12046), .ZN(
        n12048) );
  MUX2_X1 U14494 ( .A(n12051), .B(n12050), .S(n12171), .Z(n12052) );
  NAND2_X1 U14495 ( .A1(n12052), .A2(n15446), .ZN(n12054) );
  AOI21_X1 U14496 ( .B1(n15462), .B2(n15442), .A(n12062), .ZN(n12053) );
  OAI22_X1 U14497 ( .A1(n12055), .A2(n12054), .B1(n12053), .B2(n12161), .ZN(
        n12059) );
  AOI21_X1 U14498 ( .B1(n12058), .B2(n12056), .A(n12171), .ZN(n12057) );
  AOI21_X1 U14499 ( .B1(n12059), .B2(n12058), .A(n12057), .ZN(n12060) );
  AOI211_X1 U14500 ( .C1(n12062), .C2(n12161), .A(n12061), .B(n12060), .ZN(
        n12069) );
  NOR2_X1 U14501 ( .A1(n12548), .A2(n12171), .ZN(n12066) );
  NOR2_X1 U14502 ( .A1(n12063), .A2(n12161), .ZN(n12065) );
  MUX2_X1 U14503 ( .A(n12066), .B(n12065), .S(n12064), .Z(n12068) );
  NAND2_X1 U14504 ( .A1(n12075), .A2(n12070), .ZN(n12073) );
  NAND2_X1 U14505 ( .A1(n12074), .A2(n12071), .ZN(n12072) );
  MUX2_X1 U14506 ( .A(n12073), .B(n12072), .S(n12171), .Z(n12078) );
  MUX2_X1 U14507 ( .A(n12075), .B(n12074), .S(n12161), .Z(n12076) );
  OAI211_X1 U14508 ( .C1(n12079), .C2(n12078), .A(n12077), .B(n12076), .ZN(
        n12084) );
  MUX2_X1 U14509 ( .A(n12081), .B(n12080), .S(n12171), .Z(n12082) );
  NAND3_X1 U14510 ( .A1(n12084), .A2(n12083), .A3(n12082), .ZN(n12089) );
  MUX2_X1 U14511 ( .A(n12086), .B(n12085), .S(n12161), .Z(n12087) );
  NAND3_X1 U14512 ( .A1(n12089), .A2(n12088), .A3(n12087), .ZN(n12100) );
  INV_X1 U14513 ( .A(n12090), .ZN(n12091) );
  MUX2_X1 U14514 ( .A(n12092), .B(n12091), .S(n12161), .Z(n12094) );
  NOR3_X1 U14515 ( .A1(n12094), .A2(n12097), .A3(n12093), .ZN(n12099) );
  OAI211_X1 U14516 ( .C1(n12097), .C2(n12096), .A(n12111), .B(n12095), .ZN(
        n12098) );
  AOI22_X1 U14517 ( .A1(n12100), .A2(n12099), .B1(n12161), .B2(n12098), .ZN(
        n12109) );
  INV_X1 U14518 ( .A(n12102), .ZN(n12108) );
  INV_X1 U14519 ( .A(n12101), .ZN(n12105) );
  OAI21_X1 U14520 ( .B1(n14777), .B2(n12103), .A(n12102), .ZN(n12104) );
  AOI21_X1 U14521 ( .B1(n12106), .B2(n12105), .A(n12104), .ZN(n12107) );
  OAI22_X1 U14522 ( .A1(n12109), .A2(n12108), .B1(n12107), .B2(n12161), .ZN(
        n12110) );
  OAI211_X1 U14523 ( .C1(n12111), .C2(n12161), .A(n12110), .B(n7451), .ZN(
        n12115) );
  MUX2_X1 U14524 ( .A(n12113), .B(n12112), .S(n12171), .Z(n12114) );
  NAND4_X1 U14525 ( .A1(n12115), .A2(n12863), .A3(n8216), .A4(n12114), .ZN(
        n12118) );
  MUX2_X1 U14526 ( .A(n14763), .B(n12161), .S(n14789), .Z(n12116) );
  OAI211_X1 U14527 ( .C1(n12171), .C2(n12539), .A(n12863), .B(n12116), .ZN(
        n12117) );
  OAI211_X1 U14528 ( .C1(n12171), .C2(n12119), .A(n12118), .B(n12117), .ZN(
        n12122) );
  AOI21_X1 U14529 ( .B1(n12837), .B2(n12120), .A(n12161), .ZN(n12121) );
  AOI21_X1 U14530 ( .B1(n12122), .B2(n12837), .A(n12121), .ZN(n12123) );
  NAND2_X1 U14531 ( .A1(n12125), .A2(n12819), .ZN(n12126) );
  AOI21_X1 U14532 ( .B1(n12126), .B2(n12136), .A(n12161), .ZN(n12127) );
  AND2_X1 U14533 ( .A1(n12127), .A2(n12130), .ZN(n12138) );
  OAI22_X1 U14534 ( .A1(n12129), .A2(n12831), .B1(n12138), .B2(n12128), .ZN(
        n12133) );
  MUX2_X1 U14535 ( .A(n12130), .B(n12137), .S(n12171), .Z(n12131) );
  INV_X1 U14536 ( .A(n12131), .ZN(n12132) );
  NOR2_X1 U14537 ( .A1(n12789), .A2(n12132), .ZN(n12141) );
  NAND3_X1 U14538 ( .A1(n12133), .A2(n12141), .A3(n12814), .ZN(n12144) );
  MUX2_X1 U14539 ( .A(n12135), .B(n12134), .S(n12171), .Z(n12143) );
  NAND3_X1 U14540 ( .A1(n12137), .A2(n12136), .A3(n12161), .ZN(n12140) );
  INV_X1 U14541 ( .A(n12138), .ZN(n12139) );
  NAND3_X1 U14542 ( .A1(n12141), .A2(n12140), .A3(n12139), .ZN(n12142) );
  NAND4_X1 U14543 ( .A1(n12144), .A2(n12768), .A3(n12143), .A4(n12142), .ZN(
        n12147) );
  MUX2_X1 U14544 ( .A(n12758), .B(n12759), .S(n12161), .Z(n12145) );
  INV_X1 U14545 ( .A(n12148), .ZN(n12149) );
  MUX2_X1 U14546 ( .A(n12150), .B(n12149), .S(n12171), .Z(n12151) );
  INV_X1 U14547 ( .A(n12153), .ZN(n12154) );
  INV_X1 U14548 ( .A(n12483), .ZN(n12978) );
  OAI211_X1 U14549 ( .C1(n6724), .C2(n12725), .A(n12156), .B(n12708), .ZN(
        n12160) );
  INV_X1 U14550 ( .A(n12697), .ZN(n12159) );
  NAND2_X1 U14551 ( .A1(n12974), .A2(n12727), .ZN(n12157) );
  MUX2_X1 U14552 ( .A(n12693), .B(n12157), .S(n12171), .Z(n12158) );
  NAND3_X1 U14553 ( .A1(n12160), .A2(n12159), .A3(n12158), .ZN(n12165) );
  MUX2_X1 U14554 ( .A(n12163), .B(n12162), .S(n12161), .Z(n12164) );
  AOI21_X1 U14555 ( .B1(n12966), .B2(n12699), .A(n12172), .ZN(n12170) );
  INV_X1 U14556 ( .A(n12669), .ZN(n12169) );
  AOI21_X1 U14557 ( .B1(n12167), .B2(n12171), .A(n12166), .ZN(n12168) );
  NAND3_X1 U14558 ( .A1(n12172), .A2(n12171), .A3(n12669), .ZN(n12173) );
  NAND3_X1 U14559 ( .A1(n12177), .A2(n12176), .A3(n12175), .ZN(n12181) );
  INV_X1 U14560 ( .A(n12178), .ZN(n12180) );
  NOR3_X1 U14561 ( .A1(n12188), .A2(n12187), .A3(n8201), .ZN(n12191) );
  OAI21_X1 U14562 ( .B1(n12192), .B2(n12189), .A(P3_B_REG_SCAN_IN), .ZN(n12190) );
  OAI22_X1 U14563 ( .A1(n12193), .A2(n12192), .B1(n12191), .B2(n12190), .ZN(
        P3_U3296) );
  INV_X1 U14564 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n12194) );
  NOR2_X1 U14565 ( .A1(n15528), .A2(n12194), .ZN(n12195) );
  AOI21_X1 U14566 ( .B1(n15528), .B2(n12199), .A(n12195), .ZN(n12196) );
  OAI21_X1 U14567 ( .B1(n12201), .B2(n13014), .A(n12196), .ZN(P3_U3390) );
  NOR2_X1 U14568 ( .A1(n15547), .A2(n12197), .ZN(n12198) );
  AOI21_X1 U14569 ( .B1(n12199), .B2(n15547), .A(n12198), .ZN(n12200) );
  OAI21_X1 U14570 ( .B1(n12201), .B2(n12957), .A(n12200), .ZN(P3_U3459) );
  INV_X1 U14571 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n12202) );
  OAI22_X1 U14572 ( .A1(n15477), .A2(n12202), .B1(n12657), .B2(n15443), .ZN(
        n12204) );
  OAI21_X1 U14573 ( .B1(n12206), .B2(n12871), .A(n6751), .ZN(P3_U3204) );
  NAND2_X1 U14574 ( .A1(n14909), .A2(n6640), .ZN(n12208) );
  NAND2_X1 U14575 ( .A1(n14267), .A2(n6638), .ZN(n12207) );
  NAND2_X1 U14576 ( .A1(n12208), .A2(n12207), .ZN(n12209) );
  XNOR2_X1 U14577 ( .A(n12209), .B(n12242), .ZN(n12234) );
  INV_X1 U14578 ( .A(n12234), .ZN(n12239) );
  NOR2_X1 U14579 ( .A1(n13999), .A2(n6646), .ZN(n12210) );
  AOI21_X1 U14580 ( .B1(n14909), .B2(n6638), .A(n12210), .ZN(n12233) );
  INV_X1 U14581 ( .A(n12233), .ZN(n12238) );
  NOR2_X1 U14582 ( .A1(n14927), .A2(n6646), .ZN(n12211) );
  AOI21_X1 U14583 ( .B1(n14738), .B2(n6638), .A(n12211), .ZN(n12228) );
  INV_X1 U14584 ( .A(n12228), .ZN(n12230) );
  NAND2_X1 U14585 ( .A1(n14738), .A2(n6640), .ZN(n12213) );
  NAND2_X1 U14586 ( .A1(n14269), .A2(n6638), .ZN(n12212) );
  NAND2_X1 U14587 ( .A1(n12213), .A2(n12212), .ZN(n12214) );
  XNOR2_X1 U14588 ( .A(n12214), .B(n12341), .ZN(n12229) );
  NAND2_X1 U14589 ( .A1(n14938), .A2(n6640), .ZN(n12216) );
  NAND2_X1 U14590 ( .A1(n14270), .A2(n6638), .ZN(n12215) );
  NAND2_X1 U14591 ( .A1(n12216), .A2(n12215), .ZN(n12217) );
  XNOR2_X1 U14592 ( .A(n12217), .B(n12341), .ZN(n12226) );
  NOR2_X1 U14593 ( .A1(n12218), .A2(n6646), .ZN(n12219) );
  AOI21_X1 U14594 ( .B1(n14938), .B2(n6638), .A(n12219), .ZN(n12224) );
  XNOR2_X1 U14595 ( .A(n12226), .B(n12224), .ZN(n14928) );
  INV_X1 U14596 ( .A(n12220), .ZN(n12221) );
  NAND2_X1 U14597 ( .A1(n12222), .A2(n12221), .ZN(n14929) );
  INV_X1 U14598 ( .A(n12224), .ZN(n12225) );
  XOR2_X1 U14599 ( .A(n12228), .B(n12229), .Z(n13898) );
  NOR2_X1 U14600 ( .A1(n14901), .A2(n6646), .ZN(n12231) );
  AOI21_X1 U14601 ( .B1(n14112), .B2(n6638), .A(n12231), .ZN(n12236) );
  OAI22_X1 U14602 ( .A1(n7609), .A2(n12340), .B1(n14901), .B2(n12338), .ZN(
        n12232) );
  XNOR2_X1 U14603 ( .A(n12232), .B(n12341), .ZN(n12235) );
  XOR2_X1 U14604 ( .A(n12236), .B(n12235), .Z(n13941) );
  XNOR2_X1 U14605 ( .A(n12234), .B(n12233), .ZN(n14902) );
  INV_X1 U14606 ( .A(n12235), .ZN(n12237) );
  NOR2_X1 U14607 ( .A1(n12237), .A2(n12236), .ZN(n14903) );
  NAND2_X1 U14608 ( .A1(n14956), .A2(n6640), .ZN(n12241) );
  NAND2_X1 U14609 ( .A1(n14572), .A2(n6638), .ZN(n12240) );
  NAND2_X1 U14610 ( .A1(n12241), .A2(n12240), .ZN(n12243) );
  XNOR2_X1 U14611 ( .A(n12243), .B(n12341), .ZN(n12249) );
  OAI22_X1 U14612 ( .A1(n14006), .A2(n12338), .B1(n14912), .B2(n6646), .ZN(
        n13995) );
  NAND2_X1 U14613 ( .A1(n14921), .A2(n6640), .ZN(n12245) );
  NAND2_X1 U14614 ( .A1(n14266), .A2(n6638), .ZN(n12244) );
  NAND2_X1 U14615 ( .A1(n12245), .A2(n12244), .ZN(n12246) );
  XNOR2_X1 U14616 ( .A(n12246), .B(n12341), .ZN(n12251) );
  NOR2_X1 U14617 ( .A1(n14128), .A2(n6646), .ZN(n12247) );
  AOI21_X1 U14618 ( .B1(n14921), .B2(n6638), .A(n12247), .ZN(n12252) );
  XNOR2_X1 U14619 ( .A(n12251), .B(n12252), .ZN(n14914) );
  INV_X1 U14620 ( .A(n12248), .ZN(n12250) );
  NAND2_X1 U14621 ( .A1(n12250), .A2(n12249), .ZN(n14915) );
  INV_X1 U14622 ( .A(n12251), .ZN(n12253) );
  NAND2_X1 U14623 ( .A1(n12253), .A2(n12252), .ZN(n12254) );
  INV_X1 U14624 ( .A(n14565), .ZN(n14944) );
  OAI22_X1 U14625 ( .A1(n14944), .A2(n12340), .B1(n14913), .B2(n12338), .ZN(
        n12255) );
  XNOR2_X1 U14626 ( .A(n12255), .B(n12341), .ZN(n12257) );
  NOR2_X1 U14627 ( .A1(n14913), .A2(n6646), .ZN(n12256) );
  AOI21_X1 U14628 ( .B1(n14565), .B2(n6638), .A(n12256), .ZN(n12258) );
  XNOR2_X1 U14629 ( .A(n12257), .B(n12258), .ZN(n13916) );
  INV_X1 U14630 ( .A(n12257), .ZN(n12259) );
  NAND2_X1 U14631 ( .A1(n12259), .A2(n12258), .ZN(n12260) );
  NAND2_X1 U14632 ( .A1(n14667), .A2(n6640), .ZN(n12262) );
  NAND2_X1 U14633 ( .A1(n14265), .A2(n6638), .ZN(n12261) );
  NAND2_X1 U14634 ( .A1(n12262), .A2(n12261), .ZN(n12263) );
  XNOR2_X1 U14635 ( .A(n12263), .B(n12341), .ZN(n12264) );
  AOI22_X1 U14636 ( .A1(n14667), .A2(n6638), .B1(n12333), .B2(n14265), .ZN(
        n12265) );
  XNOR2_X1 U14637 ( .A(n12264), .B(n12265), .ZN(n13963) );
  INV_X1 U14638 ( .A(n12264), .ZN(n12266) );
  NAND2_X1 U14639 ( .A1(n12266), .A2(n12265), .ZN(n12267) );
  INV_X1 U14640 ( .A(n14545), .ZN(n13966) );
  NOR2_X1 U14641 ( .A1(n13966), .A2(n6646), .ZN(n12268) );
  AOI21_X1 U14642 ( .B1(n14662), .B2(n6638), .A(n12268), .ZN(n12273) );
  NAND2_X1 U14643 ( .A1(n14662), .A2(n6640), .ZN(n12270) );
  NAND2_X1 U14644 ( .A1(n14545), .A2(n6638), .ZN(n12269) );
  NAND2_X1 U14645 ( .A1(n12270), .A2(n12269), .ZN(n12271) );
  XNOR2_X1 U14646 ( .A(n12271), .B(n12341), .ZN(n12275) );
  XOR2_X1 U14647 ( .A(n12273), .B(n12275), .Z(n13877) );
  INV_X1 U14648 ( .A(n13877), .ZN(n12272) );
  INV_X1 U14649 ( .A(n12273), .ZN(n12274) );
  NAND2_X1 U14650 ( .A1(n12275), .A2(n12274), .ZN(n13886) );
  NAND2_X1 U14651 ( .A1(n14639), .A2(n6640), .ZN(n12277) );
  NAND2_X1 U14652 ( .A1(n14497), .A2(n6638), .ZN(n12276) );
  NAND2_X1 U14653 ( .A1(n12277), .A2(n12276), .ZN(n12278) );
  XNOR2_X1 U14654 ( .A(n12278), .B(n12341), .ZN(n12292) );
  AOI22_X1 U14655 ( .A1(n14639), .A2(n6638), .B1(n12333), .B2(n14497), .ZN(
        n12293) );
  XNOR2_X1 U14656 ( .A(n12292), .B(n12293), .ZN(n13952) );
  AOI22_X1 U14657 ( .A1(n14644), .A2(n6640), .B1(n6638), .B2(n14506), .ZN(
        n12279) );
  XNOR2_X1 U14658 ( .A(n12279), .B(n12341), .ZN(n12281) );
  AOI22_X1 U14659 ( .A1(n14644), .A2(n6638), .B1(n12333), .B2(n14506), .ZN(
        n12280) );
  NAND2_X1 U14660 ( .A1(n12281), .A2(n12280), .ZN(n12289) );
  INV_X1 U14661 ( .A(n12289), .ZN(n12285) );
  XNOR2_X1 U14662 ( .A(n12281), .B(n12280), .ZN(n13891) );
  OAI22_X1 U14663 ( .A1(n14518), .A2(n12340), .B1(n14532), .B2(n12338), .ZN(
        n12282) );
  XNOR2_X1 U14664 ( .A(n12282), .B(n12341), .ZN(n12287) );
  OAI22_X1 U14665 ( .A1(n14518), .A2(n12338), .B1(n14532), .B2(n6646), .ZN(
        n12288) );
  NAND2_X1 U14666 ( .A1(n12287), .A2(n12288), .ZN(n13888) );
  INV_X1 U14667 ( .A(n13888), .ZN(n12283) );
  NOR2_X1 U14668 ( .A1(n13891), .A2(n12283), .ZN(n12284) );
  OR2_X1 U14669 ( .A1(n12285), .A2(n12284), .ZN(n13948) );
  AND2_X1 U14670 ( .A1(n13952), .A2(n13948), .ZN(n12286) );
  AND2_X1 U14671 ( .A1(n13886), .A2(n12286), .ZN(n12291) );
  INV_X1 U14672 ( .A(n12286), .ZN(n12290) );
  XOR2_X1 U14673 ( .A(n12288), .B(n12287), .Z(n13932) );
  AND2_X1 U14674 ( .A1(n13932), .A2(n12289), .ZN(n13946) );
  INV_X1 U14675 ( .A(n12292), .ZN(n12294) );
  NAND2_X1 U14676 ( .A1(n12294), .A2(n12293), .ZN(n13867) );
  NAND2_X1 U14677 ( .A1(n14633), .A2(n6640), .ZN(n12296) );
  NAND2_X1 U14678 ( .A1(n14470), .A2(n6638), .ZN(n12295) );
  NAND2_X1 U14679 ( .A1(n12296), .A2(n12295), .ZN(n12297) );
  XNOR2_X1 U14680 ( .A(n12297), .B(n12341), .ZN(n12301) );
  INV_X1 U14681 ( .A(n12301), .ZN(n12299) );
  OAI22_X1 U14682 ( .A1(n14461), .A2(n12338), .B1(n13956), .B2(n6646), .ZN(
        n12302) );
  INV_X1 U14683 ( .A(n12302), .ZN(n12298) );
  NAND2_X1 U14684 ( .A1(n12299), .A2(n12298), .ZN(n12300) );
  AND2_X1 U14685 ( .A1(n13867), .A2(n12300), .ZN(n12304) );
  INV_X1 U14686 ( .A(n12300), .ZN(n12303) );
  XOR2_X1 U14687 ( .A(n12302), .B(n12301), .Z(n13869) );
  AOI21_X2 U14688 ( .B1(n13950), .B2(n12304), .A(n7684), .ZN(n13922) );
  OAI22_X1 U14689 ( .A1(n14448), .A2(n12338), .B1(n12305), .B2(n6646), .ZN(
        n12310) );
  NAND2_X1 U14690 ( .A1(n14626), .A2(n6640), .ZN(n12307) );
  NAND2_X1 U14691 ( .A1(n14423), .A2(n6638), .ZN(n12306) );
  NAND2_X1 U14692 ( .A1(n12307), .A2(n12306), .ZN(n12308) );
  XNOR2_X1 U14693 ( .A(n12308), .B(n12341), .ZN(n12309) );
  XOR2_X1 U14694 ( .A(n12310), .B(n12309), .Z(n13923) );
  INV_X1 U14695 ( .A(n12309), .ZN(n12312) );
  INV_X1 U14696 ( .A(n12310), .ZN(n12311) );
  NAND2_X1 U14697 ( .A1(n12312), .A2(n12311), .ZN(n12313) );
  OAI22_X1 U14698 ( .A1(n14620), .A2(n12338), .B1(n13986), .B2(n6646), .ZN(
        n12318) );
  NAND2_X1 U14699 ( .A1(n14431), .A2(n6640), .ZN(n12315) );
  NAND2_X1 U14700 ( .A1(n14264), .A2(n6638), .ZN(n12314) );
  NAND2_X1 U14701 ( .A1(n12315), .A2(n12314), .ZN(n12316) );
  XNOR2_X1 U14702 ( .A(n12316), .B(n12341), .ZN(n12317) );
  XOR2_X1 U14703 ( .A(n12318), .B(n12317), .Z(n13907) );
  INV_X1 U14704 ( .A(n12317), .ZN(n12320) );
  INV_X1 U14705 ( .A(n12318), .ZN(n12319) );
  NAND2_X1 U14706 ( .A1(n14614), .A2(n6640), .ZN(n12322) );
  NAND2_X1 U14707 ( .A1(n14424), .A2(n6638), .ZN(n12321) );
  NAND2_X1 U14708 ( .A1(n12322), .A2(n12321), .ZN(n12323) );
  XNOR2_X1 U14709 ( .A(n12323), .B(n12341), .ZN(n12324) );
  AOI22_X1 U14710 ( .A1(n14614), .A2(n6638), .B1(n12333), .B2(n14424), .ZN(
        n12325) );
  XNOR2_X1 U14711 ( .A(n12324), .B(n12325), .ZN(n13984) );
  NAND2_X1 U14712 ( .A1(n13983), .A2(n13984), .ZN(n12328) );
  INV_X1 U14713 ( .A(n12324), .ZN(n12326) );
  NAND2_X1 U14714 ( .A1(n12326), .A2(n12325), .ZN(n12327) );
  NAND2_X1 U14715 ( .A1(n14608), .A2(n6640), .ZN(n12331) );
  NAND2_X1 U14716 ( .A1(n14263), .A2(n6638), .ZN(n12330) );
  NAND2_X1 U14717 ( .A1(n12331), .A2(n12330), .ZN(n12332) );
  XNOR2_X1 U14718 ( .A(n12332), .B(n12341), .ZN(n12334) );
  AOI22_X1 U14719 ( .A1(n14608), .A2(n6638), .B1(n12333), .B2(n14263), .ZN(
        n12335) );
  XNOR2_X1 U14720 ( .A(n12334), .B(n12335), .ZN(n13859) );
  INV_X1 U14721 ( .A(n12334), .ZN(n12336) );
  OAI22_X1 U14722 ( .A1(n14600), .A2(n12338), .B1(n12339), .B2(n6646), .ZN(
        n12344) );
  OAI22_X1 U14723 ( .A1(n14600), .A2(n12340), .B1(n12339), .B2(n12338), .ZN(
        n12342) );
  XNOR2_X1 U14724 ( .A(n12342), .B(n12341), .ZN(n12343) );
  XOR2_X1 U14725 ( .A(n12344), .B(n12343), .Z(n12345) );
  XNOR2_X1 U14726 ( .A(n12346), .B(n12345), .ZN(n12353) );
  OR2_X1 U14727 ( .A1(n14191), .A2(n14533), .ZN(n12348) );
  NAND2_X1 U14728 ( .A1(n14263), .A2(n14571), .ZN(n12347) );
  OAI22_X1 U14729 ( .A1(n13918), .A2(n14599), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12349), .ZN(n12351) );
  NOR2_X1 U14730 ( .A1(n14600), .A2(n14005), .ZN(n12350) );
  AOI211_X1 U14731 ( .C1(n14380), .C2(n14001), .A(n12351), .B(n12350), .ZN(
        n12352) );
  OAI21_X1 U14732 ( .B1(n12353), .B2(n14932), .A(n12352), .ZN(P1_U3220) );
  XNOR2_X1 U14733 ( .A(n6864), .B(n12390), .ZN(n12414) );
  XNOR2_X1 U14734 ( .A(n12414), .B(n12699), .ZN(n12415) );
  AND2_X1 U14735 ( .A1(n12356), .A2(n12539), .ZN(n12354) );
  OR2_X2 U14736 ( .A1(n12355), .A2(n12354), .ZN(n12359) );
  INV_X1 U14737 ( .A(n12356), .ZN(n12357) );
  NAND2_X1 U14738 ( .A1(n12357), .A2(n14763), .ZN(n12358) );
  XNOR2_X1 U14739 ( .A(n12360), .B(n12390), .ZN(n12361) );
  XNOR2_X1 U14740 ( .A(n12361), .B(n12848), .ZN(n12524) );
  INV_X1 U14741 ( .A(n12361), .ZN(n12362) );
  NAND2_X1 U14742 ( .A1(n12362), .A2(n12848), .ZN(n12363) );
  XNOR2_X1 U14743 ( .A(n12856), .B(n12390), .ZN(n12364) );
  XNOR2_X1 U14744 ( .A(n12364), .B(n12861), .ZN(n12459) );
  NAND2_X1 U14745 ( .A1(n12364), .A2(n12833), .ZN(n12365) );
  XNOR2_X1 U14746 ( .A(n12465), .B(n12416), .ZN(n12366) );
  XNOR2_X1 U14747 ( .A(n12366), .B(n12849), .ZN(n12467) );
  INV_X1 U14748 ( .A(n12366), .ZN(n12367) );
  NAND2_X1 U14749 ( .A1(n12367), .A2(n12849), .ZN(n12368) );
  XNOR2_X1 U14750 ( .A(n12503), .B(n12390), .ZN(n12369) );
  XNOR2_X1 U14751 ( .A(n12369), .B(n12834), .ZN(n12505) );
  INV_X1 U14752 ( .A(n12369), .ZN(n12370) );
  NAND2_X1 U14753 ( .A1(n12370), .A2(n12834), .ZN(n12371) );
  XNOR2_X1 U14754 ( .A(n12997), .B(n12390), .ZN(n12372) );
  XNOR2_X1 U14755 ( .A(n12372), .B(n12817), .ZN(n12407) );
  NAND2_X1 U14756 ( .A1(n12408), .A2(n12407), .ZN(n12406) );
  NAND2_X1 U14757 ( .A1(n12372), .A2(n12784), .ZN(n12373) );
  XNOR2_X1 U14758 ( .A(n12788), .B(n12416), .ZN(n12374) );
  XNOR2_X1 U14759 ( .A(n12374), .B(n12538), .ZN(n12488) );
  INV_X1 U14760 ( .A(n12374), .ZN(n12375) );
  NAND2_X1 U14761 ( .A1(n12375), .A2(n12538), .ZN(n12376) );
  XNOR2_X1 U14762 ( .A(n12989), .B(n12390), .ZN(n12377) );
  XNOR2_X1 U14763 ( .A(n12377), .B(n12755), .ZN(n12441) );
  NAND2_X1 U14764 ( .A1(n12377), .A2(n12755), .ZN(n12378) );
  XNOR2_X1 U14765 ( .A(n12985), .B(n6823), .ZN(n12380) );
  INV_X1 U14766 ( .A(n12380), .ZN(n12381) );
  AND2_X1 U14767 ( .A1(n12382), .A2(n12381), .ZN(n12383) );
  XNOR2_X1 U14768 ( .A(n12483), .B(n12416), .ZN(n12477) );
  XNOR2_X1 U14769 ( .A(n12749), .B(n12390), .ZN(n12385) );
  OAI22_X1 U14770 ( .A1(n12477), .A2(n12476), .B1(n12754), .B2(n12385), .ZN(
        n12388) );
  INV_X1 U14771 ( .A(n12385), .ZN(n12473) );
  OAI21_X1 U14772 ( .B1(n12473), .B2(n12728), .A(n12743), .ZN(n12384) );
  NAND2_X1 U14773 ( .A1(n12477), .A2(n12384), .ZN(n12387) );
  NAND3_X1 U14774 ( .A1(n12385), .A2(n12754), .A3(n12476), .ZN(n12386) );
  XNOR2_X1 U14775 ( .A(n12454), .B(n12390), .ZN(n12389) );
  XNOR2_X1 U14776 ( .A(n12389), .B(n12727), .ZN(n12450) );
  XNOR2_X1 U14777 ( .A(n12898), .B(n12390), .ZN(n12391) );
  XNOR2_X1 U14778 ( .A(n12391), .B(n12684), .ZN(n12512) );
  INV_X1 U14779 ( .A(n12391), .ZN(n12392) );
  NOR2_X1 U14780 ( .A1(n12526), .A2(n12683), .ZN(n12395) );
  OAI22_X1 U14781 ( .A1(n12527), .A2(n12684), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12393), .ZN(n12394) );
  AOI211_X1 U14782 ( .C1(n12688), .C2(n12530), .A(n12395), .B(n12394), .ZN(
        n12398) );
  NAND2_X1 U14783 ( .A1(n6864), .A2(n12517), .ZN(n12397) );
  XNOR2_X1 U14784 ( .A(n12474), .B(n12473), .ZN(n12475) );
  XNOR2_X1 U14785 ( .A(n12475), .B(n12754), .ZN(n12405) );
  NOR2_X1 U14786 ( .A1(n12527), .A2(n12442), .ZN(n12402) );
  OAI22_X1 U14787 ( .A1(n12526), .A2(n12476), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12400), .ZN(n12401) );
  AOI211_X1 U14788 ( .C1(n12746), .C2(n12530), .A(n12402), .B(n12401), .ZN(
        n12404) );
  NAND2_X1 U14789 ( .A1(n12749), .A2(n12517), .ZN(n12403) );
  OAI211_X1 U14790 ( .C1(n12405), .C2(n12520), .A(n12404), .B(n12403), .ZN(
        P3_U3156) );
  OAI211_X1 U14791 ( .C1(n12408), .C2(n12407), .A(n12406), .B(n12522), .ZN(
        n12413) );
  NOR2_X1 U14792 ( .A1(n12527), .A2(n12800), .ZN(n12411) );
  OAI21_X1 U14793 ( .B1(n12526), .B2(n12799), .A(n12409), .ZN(n12410) );
  AOI211_X1 U14794 ( .C1(n12806), .C2(n12530), .A(n12411), .B(n12410), .ZN(
        n12412) );
  OAI211_X1 U14795 ( .C1(n12533), .C2(n12997), .A(n12413), .B(n12412), .ZN(
        P3_U3159) );
  XNOR2_X1 U14796 ( .A(n12669), .B(n12416), .ZN(n12417) );
  NOR2_X1 U14797 ( .A1(n12526), .A2(n12536), .ZN(n12420) );
  OAI22_X1 U14798 ( .A1(n12527), .A2(n12514), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12418), .ZN(n12419) );
  AOI211_X1 U14799 ( .C1(n12672), .C2(n12530), .A(n12420), .B(n12419), .ZN(
        n12422) );
  NAND2_X1 U14800 ( .A1(n12671), .A2(n12517), .ZN(n12421) );
  MUX2_X1 U14801 ( .A(n12546), .B(n12424), .S(n12423), .Z(n12426) );
  XNOR2_X1 U14802 ( .A(n12426), .B(n12425), .ZN(n12427) );
  NAND2_X1 U14803 ( .A1(n12427), .A2(n12522), .ZN(n12437) );
  AOI21_X1 U14804 ( .B1(n12517), .B2(n12429), .A(n12428), .ZN(n12436) );
  OAI22_X1 U14805 ( .A1(n12431), .A2(n12527), .B1(n12526), .B2(n12430), .ZN(
        n12432) );
  INV_X1 U14806 ( .A(n12432), .ZN(n12435) );
  NAND2_X1 U14807 ( .A1(n12530), .A2(n12433), .ZN(n12434) );
  NAND4_X1 U14808 ( .A1(n12437), .A2(n12436), .A3(n12435), .A4(n12434), .ZN(
        P3_U3161) );
  INV_X1 U14809 ( .A(n12438), .ZN(n12439) );
  AOI21_X1 U14810 ( .B1(n12441), .B2(n12440), .A(n12439), .ZN(n12448) );
  NOR2_X1 U14811 ( .A1(n12526), .A2(n12442), .ZN(n12445) );
  INV_X1 U14812 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n12443) );
  OAI22_X1 U14813 ( .A1(n12527), .A2(n12799), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12443), .ZN(n12444) );
  AOI211_X1 U14814 ( .C1(n12777), .C2(n12530), .A(n12445), .B(n12444), .ZN(
        n12447) );
  NAND2_X1 U14815 ( .A1(n12989), .A2(n12517), .ZN(n12446) );
  OAI211_X1 U14816 ( .C1(n12448), .C2(n12520), .A(n12447), .B(n12446), .ZN(
        P3_U3163) );
  XOR2_X1 U14817 ( .A(n12450), .B(n12449), .Z(n12457) );
  NOR2_X1 U14818 ( .A1(n12527), .A2(n12476), .ZN(n12453) );
  INV_X1 U14819 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n12451) );
  OAI22_X1 U14820 ( .A1(n12526), .A2(n12684), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12451), .ZN(n12452) );
  AOI211_X1 U14821 ( .C1(n12716), .C2(n12530), .A(n12453), .B(n12452), .ZN(
        n12456) );
  NAND2_X1 U14822 ( .A1(n12454), .A2(n12517), .ZN(n12455) );
  OAI211_X1 U14823 ( .C1(n12457), .C2(n12520), .A(n12456), .B(n12455), .ZN(
        P3_U3165) );
  OAI211_X1 U14824 ( .C1(n12460), .C2(n12459), .A(n12458), .B(n12522), .ZN(
        n12464) );
  NOR2_X1 U14825 ( .A1(n12527), .A2(n12879), .ZN(n12462) );
  NAND2_X1 U14826 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12610)
         );
  OAI21_X1 U14827 ( .B1(n12526), .B2(n12816), .A(n12610), .ZN(n12461) );
  AOI211_X1 U14828 ( .C1(n12854), .C2(n12530), .A(n12462), .B(n12461), .ZN(
        n12463) );
  OAI211_X1 U14829 ( .C1(n12856), .C2(n12533), .A(n12464), .B(n12463), .ZN(
        P3_U3166) );
  INV_X1 U14830 ( .A(n12465), .ZN(n13005) );
  OAI211_X1 U14831 ( .C1(n12468), .C2(n12467), .A(n12466), .B(n12522), .ZN(
        n12472) );
  NOR2_X1 U14832 ( .A1(n12527), .A2(n12861), .ZN(n12470) );
  NAND2_X1 U14833 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12626)
         );
  OAI21_X1 U14834 ( .B1(n12526), .B2(n12800), .A(n12626), .ZN(n12469) );
  AOI211_X1 U14835 ( .C1(n12840), .C2(n12530), .A(n12470), .B(n12469), .ZN(
        n12471) );
  OAI211_X1 U14836 ( .C1(n13005), .C2(n12533), .A(n12472), .B(n12471), .ZN(
        P3_U3168) );
  OAI22_X1 U14837 ( .A1(n12475), .A2(n12728), .B1(n12474), .B2(n12473), .ZN(
        n12479) );
  XNOR2_X1 U14838 ( .A(n12477), .B(n12476), .ZN(n12478) );
  XNOR2_X1 U14839 ( .A(n12479), .B(n12478), .ZN(n12486) );
  NOR2_X1 U14840 ( .A1(n12527), .A2(n12754), .ZN(n12482) );
  OAI22_X1 U14841 ( .A1(n12526), .A2(n12513), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12480), .ZN(n12481) );
  AOI211_X1 U14842 ( .C1(n12732), .C2(n12530), .A(n12482), .B(n12481), .ZN(
        n12485) );
  NAND2_X1 U14843 ( .A1(n12483), .A2(n12517), .ZN(n12484) );
  OAI211_X1 U14844 ( .C1(n12486), .C2(n12520), .A(n12485), .B(n12484), .ZN(
        P3_U3169) );
  INV_X1 U14845 ( .A(n12788), .ZN(n12495) );
  OAI211_X1 U14846 ( .C1(n12489), .C2(n12488), .A(n12487), .B(n12522), .ZN(
        n12494) );
  NOR2_X1 U14847 ( .A1(n12527), .A2(n12817), .ZN(n12492) );
  OAI22_X1 U14848 ( .A1(n12526), .A2(n12755), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12490), .ZN(n12491) );
  AOI211_X1 U14849 ( .C1(n12791), .C2(n12530), .A(n12492), .B(n12491), .ZN(
        n12493) );
  OAI211_X1 U14850 ( .C1(n12495), .C2(n12533), .A(n12494), .B(n12493), .ZN(
        P3_U3173) );
  XNOR2_X1 U14851 ( .A(n12496), .B(n12772), .ZN(n12502) );
  NOR2_X1 U14852 ( .A1(n12526), .A2(n12754), .ZN(n12499) );
  INV_X1 U14853 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n12497) );
  OAI22_X1 U14854 ( .A1(n12527), .A2(n12755), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12497), .ZN(n12498) );
  AOI211_X1 U14855 ( .C1(n12763), .C2(n12530), .A(n12499), .B(n12498), .ZN(
        n12501) );
  NAND2_X1 U14856 ( .A1(n12985), .A2(n12517), .ZN(n12500) );
  OAI211_X1 U14857 ( .C1(n12502), .C2(n12520), .A(n12501), .B(n12500), .ZN(
        P3_U3175) );
  INV_X1 U14858 ( .A(n12503), .ZN(n13001) );
  OAI211_X1 U14859 ( .C1(n12506), .C2(n12505), .A(n12504), .B(n12522), .ZN(
        n12510) );
  NOR2_X1 U14860 ( .A1(n12527), .A2(n12816), .ZN(n12508) );
  NAND2_X1 U14861 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12643)
         );
  OAI21_X1 U14862 ( .B1(n12526), .B2(n12817), .A(n12643), .ZN(n12507) );
  AOI211_X1 U14863 ( .C1(n12822), .C2(n12530), .A(n12508), .B(n12507), .ZN(
        n12509) );
  OAI211_X1 U14864 ( .C1(n13001), .C2(n12533), .A(n12510), .B(n12509), .ZN(
        P3_U3178) );
  XOR2_X1 U14865 ( .A(n12512), .B(n12511), .Z(n12521) );
  NOR2_X1 U14866 ( .A1(n12527), .A2(n12513), .ZN(n12516) );
  INV_X1 U14867 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n13159) );
  OAI22_X1 U14868 ( .A1(n12526), .A2(n12514), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13159), .ZN(n12515) );
  AOI211_X1 U14869 ( .C1(n12702), .C2(n12530), .A(n12516), .B(n12515), .ZN(
        n12519) );
  NAND2_X1 U14870 ( .A1(n12898), .A2(n12517), .ZN(n12518) );
  OAI211_X1 U14871 ( .C1(n12521), .C2(n12520), .A(n12519), .B(n12518), .ZN(
        P3_U3180) );
  OAI211_X1 U14872 ( .C1(n12525), .C2(n12524), .A(n12523), .B(n12522), .ZN(
        n12532) );
  NOR2_X1 U14873 ( .A1(n12526), .A2(n12861), .ZN(n12529) );
  NAND2_X1 U14874 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12589)
         );
  OAI21_X1 U14875 ( .B1(n12527), .B2(n14763), .A(n12589), .ZN(n12528) );
  AOI211_X1 U14876 ( .C1(n12865), .C2(n12530), .A(n12529), .B(n12528), .ZN(
        n12531) );
  OAI211_X1 U14877 ( .C1(n13015), .C2(n12533), .A(n12532), .B(n12531), .ZN(
        P3_U3181) );
  MUX2_X1 U14878 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12534), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14879 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(n12535), .S(P3_U3897), .Z(
        P3_U3521) );
  INV_X1 U14880 ( .A(n12536), .ZN(n12665) );
  MUX2_X1 U14881 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(n12665), .S(P3_U3897), .Z(
        P3_U3520) );
  MUX2_X1 U14882 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12537), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14883 ( .A(n12699), .B(P3_DATAO_REG_27__SCAN_IN), .S(n12550), .Z(
        P3_U3518) );
  MUX2_X1 U14884 ( .A(n12712), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12550), .Z(
        P3_U3517) );
  MUX2_X1 U14885 ( .A(n12727), .B(P3_DATAO_REG_25__SCAN_IN), .S(n12550), .Z(
        P3_U3516) );
  MUX2_X1 U14886 ( .A(n12743), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12550), .Z(
        P3_U3515) );
  MUX2_X1 U14887 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n12728), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U14888 ( .A(n12772), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12550), .Z(
        P3_U3513) );
  MUX2_X1 U14889 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12785), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14890 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12538), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14891 ( .A(n12784), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12550), .Z(
        P3_U3510) );
  MUX2_X1 U14892 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12849), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14893 ( .A(n12833), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12550), .Z(
        P3_U3507) );
  MUX2_X1 U14894 ( .A(n12848), .B(P3_DATAO_REG_15__SCAN_IN), .S(n12550), .Z(
        P3_U3506) );
  MUX2_X1 U14895 ( .A(n12539), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12550), .Z(
        P3_U3505) );
  MUX2_X1 U14896 ( .A(n12540), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12550), .Z(
        P3_U3504) );
  MUX2_X1 U14897 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12541), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14898 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n12542), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U14899 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12543), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14900 ( .A(n12544), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12550), .Z(
        P3_U3500) );
  MUX2_X1 U14901 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12545), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14902 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12546), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14903 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12547), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14904 ( .A(n12548), .B(P3_DATAO_REG_4__SCAN_IN), .S(n12550), .Z(
        P3_U3495) );
  MUX2_X1 U14905 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12549), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14906 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n9997), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U14907 ( .A(n15463), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12550), .Z(
        P3_U3491) );
  AOI21_X1 U14908 ( .B1(n14798), .B2(n12552), .A(n12551), .ZN(n12566) );
  AOI21_X1 U14909 ( .B1(n12555), .B2(n12554), .A(n12553), .ZN(n12558) );
  AOI21_X1 U14910 ( .B1(n15405), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n12556), 
        .ZN(n12557) );
  OAI21_X1 U14911 ( .B1(n12558), .B2(n15434), .A(n12557), .ZN(n12563) );
  AOI21_X1 U14912 ( .B1(n11868), .B2(n12560), .A(n12559), .ZN(n12561) );
  NOR2_X1 U14913 ( .A1(n12561), .A2(n15438), .ZN(n12562) );
  AOI211_X1 U14914 ( .C1(n15430), .C2(n12564), .A(n12563), .B(n12562), .ZN(
        n12565) );
  OAI21_X1 U14915 ( .B1(n12566), .B2(n15425), .A(n12565), .ZN(P3_U3195) );
  AOI21_X1 U14916 ( .B1(n12569), .B2(n12568), .A(n12567), .ZN(n12582) );
  XNOR2_X1 U14917 ( .A(n12571), .B(n12570), .ZN(n12580) );
  AOI21_X1 U14918 ( .B1(n15405), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n12572), 
        .ZN(n12577) );
  OAI211_X1 U14919 ( .C1(n12575), .C2(n12574), .A(n12652), .B(n12573), .ZN(
        n12576) );
  OAI211_X1 U14920 ( .C1(n12645), .C2(n12578), .A(n12577), .B(n12576), .ZN(
        n12579) );
  AOI21_X1 U14921 ( .B1(n12580), .B2(n15404), .A(n12579), .ZN(n12581) );
  OAI21_X1 U14922 ( .B1(n12582), .B2(n15425), .A(n12581), .ZN(P3_U3196) );
  AOI21_X1 U14923 ( .B1(n12585), .B2(n12584), .A(n12583), .ZN(n12600) );
  AOI21_X1 U14924 ( .B1(n12955), .B2(n12587), .A(n12586), .ZN(n12588) );
  OR2_X1 U14925 ( .A1(n12588), .A2(n15425), .ZN(n12599) );
  OAI21_X1 U14926 ( .B1(n15421), .B2(n12590), .A(n12589), .ZN(n12596) );
  AOI21_X1 U14927 ( .B1(n12593), .B2(n12592), .A(n12591), .ZN(n12594) );
  NOR2_X1 U14928 ( .A1(n12594), .A2(n15434), .ZN(n12595) );
  AOI211_X1 U14929 ( .C1(n15430), .C2(n12597), .A(n12596), .B(n12595), .ZN(
        n12598) );
  OAI211_X1 U14930 ( .C1(n12600), .C2(n15438), .A(n12599), .B(n12598), .ZN(
        P3_U3197) );
  AOI21_X1 U14931 ( .B1(n12603), .B2(n12602), .A(n12601), .ZN(n12619) );
  INV_X1 U14932 ( .A(n12604), .ZN(n12605) );
  NAND2_X1 U14933 ( .A1(n12606), .A2(n12605), .ZN(n12607) );
  XNOR2_X1 U14934 ( .A(n12608), .B(n12607), .ZN(n12617) );
  NAND2_X1 U14935 ( .A1(n15430), .A2(n12609), .ZN(n12611) );
  OAI211_X1 U14936 ( .C1(n13153), .C2(n15421), .A(n12611), .B(n12610), .ZN(
        n12616) );
  AOI21_X1 U14937 ( .B1(n6699), .B2(n12613), .A(n12612), .ZN(n12614) );
  NOR2_X1 U14938 ( .A1(n12614), .A2(n15438), .ZN(n12615) );
  AOI211_X1 U14939 ( .C1(n12652), .C2(n12617), .A(n12616), .B(n12615), .ZN(
        n12618) );
  OAI21_X1 U14940 ( .B1(n12619), .B2(n15425), .A(n12618), .ZN(P3_U3198) );
  AOI21_X1 U14941 ( .B1(n12945), .B2(n12621), .A(n12620), .ZN(n12636) );
  INV_X1 U14942 ( .A(n12622), .ZN(n12623) );
  NOR2_X1 U14943 ( .A1(n12623), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n12625) );
  OAI21_X1 U14944 ( .B1(n12625), .B2(n12624), .A(n15404), .ZN(n12635) );
  INV_X1 U14945 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n12627) );
  OAI21_X1 U14946 ( .B1(n15421), .B2(n12627), .A(n12626), .ZN(n12632) );
  AOI211_X1 U14947 ( .C1(n12630), .C2(n12629), .A(n12628), .B(n15434), .ZN(
        n12631) );
  AOI211_X1 U14948 ( .C1(n15430), .C2(n12633), .A(n12632), .B(n12631), .ZN(
        n12634) );
  OAI211_X1 U14949 ( .C1(n12636), .C2(n15425), .A(n12635), .B(n12634), .ZN(
        P3_U3199) );
  OAI21_X1 U14950 ( .B1(n12641), .B2(n12640), .A(n12639), .ZN(n12651) );
  NAND2_X1 U14951 ( .A1(n15405), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n12642) );
  OAI211_X1 U14952 ( .C1(n12645), .C2(n12644), .A(n12643), .B(n12642), .ZN(
        n12650) );
  AOI21_X1 U14953 ( .B1(n6700), .B2(n12647), .A(n12646), .ZN(n12648) );
  NOR2_X1 U14954 ( .A1(n12648), .A2(n15438), .ZN(n12649) );
  OAI21_X1 U14955 ( .B1(n12654), .B2(n15425), .A(n12653), .ZN(P3_U3200) );
  OAI22_X1 U14956 ( .A1(n12871), .A2(n14786), .B1(n12657), .B2(n15443), .ZN(
        n12659) );
  AOI21_X1 U14957 ( .B1(n12871), .B2(P3_REG2_REG_31__SCAN_IN), .A(n12659), 
        .ZN(n12658) );
  OAI21_X1 U14958 ( .B1(n12960), .B2(n12867), .A(n12658), .ZN(P3_U3202) );
  AOI21_X1 U14959 ( .B1(n12871), .B2(P3_REG2_REG_30__SCAN_IN), .A(n12659), 
        .ZN(n12660) );
  OAI21_X1 U14960 ( .B1(n14787), .B2(n12867), .A(n12660), .ZN(P3_U3203) );
  NAND2_X1 U14961 ( .A1(n12661), .A2(n12669), .ZN(n12662) );
  NAND2_X1 U14962 ( .A1(n12662), .A2(n15466), .ZN(n12663) );
  AOI22_X1 U14963 ( .A1(n12665), .A2(n15461), .B1(n15464), .B2(n12699), .ZN(
        n12666) );
  INV_X1 U14964 ( .A(n12892), .ZN(n12676) );
  NAND2_X1 U14965 ( .A1(n12680), .A2(n12668), .ZN(n12670) );
  XNOR2_X1 U14966 ( .A(n12670), .B(n12669), .ZN(n12890) );
  AOI22_X1 U14967 ( .A1(n12871), .A2(P3_REG2_REG_28__SCAN_IN), .B1(n15473), 
        .B2(n12672), .ZN(n12673) );
  OAI21_X1 U14968 ( .B1(n12963), .B2(n12867), .A(n12673), .ZN(n12674) );
  AOI21_X1 U14969 ( .B1(n12890), .B2(n12869), .A(n12674), .ZN(n12675) );
  OAI21_X1 U14970 ( .B1(n12676), .B2(n12871), .A(n12675), .ZN(P3_U3205) );
  INV_X1 U14971 ( .A(n12677), .ZN(n12678) );
  AOI21_X1 U14972 ( .B1(n12681), .B2(n12679), .A(n12678), .ZN(n12687) );
  OAI22_X1 U14973 ( .A1(n12684), .A2(n15450), .B1(n12683), .B2(n15448), .ZN(
        n12685) );
  AOI21_X1 U14974 ( .B1(n12895), .B2(n15453), .A(n12685), .ZN(n12686) );
  INV_X1 U14975 ( .A(n12894), .ZN(n12692) );
  AOI22_X1 U14976 ( .A1(n12871), .A2(P3_REG2_REG_27__SCAN_IN), .B1(n15473), 
        .B2(n12688), .ZN(n12689) );
  OAI21_X1 U14977 ( .B1(n12966), .B2(n12867), .A(n12689), .ZN(n12690) );
  AOI21_X1 U14978 ( .B1(n12895), .B2(n15474), .A(n12690), .ZN(n12691) );
  OAI21_X1 U14979 ( .B1(n12692), .B2(n12871), .A(n12691), .ZN(P3_U3206) );
  NAND2_X1 U14980 ( .A1(n12694), .A2(n12693), .ZN(n12695) );
  XNOR2_X1 U14981 ( .A(n12695), .B(n12697), .ZN(n12899) );
  XOR2_X1 U14982 ( .A(n12696), .B(n12697), .Z(n12698) );
  NAND2_X1 U14983 ( .A1(n12698), .A2(n15466), .ZN(n12701) );
  AOI22_X1 U14984 ( .A1(n15461), .A2(n12699), .B1(n12727), .B2(n15464), .ZN(
        n12700) );
  OAI211_X1 U14985 ( .C1(n15470), .C2(n12899), .A(n12701), .B(n12700), .ZN(
        n12900) );
  NAND2_X1 U14986 ( .A1(n12900), .A2(n15477), .ZN(n12707) );
  INV_X1 U14987 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n12704) );
  INV_X1 U14988 ( .A(n12702), .ZN(n12703) );
  OAI22_X1 U14989 ( .A1(n15477), .A2(n12704), .B1(n12703), .B2(n15443), .ZN(
        n12705) );
  AOI21_X1 U14990 ( .B1(n12898), .B2(n12885), .A(n12705), .ZN(n12706) );
  OAI211_X1 U14991 ( .C1(n12752), .C2(n12899), .A(n12707), .B(n12706), .ZN(
        P3_U3207) );
  INV_X1 U14992 ( .A(n12708), .ZN(n12711) );
  XNOR2_X1 U14993 ( .A(n12709), .B(n12711), .ZN(n12715) );
  OAI211_X1 U14994 ( .C1(n6725), .C2(n12711), .A(n12710), .B(n15466), .ZN(
        n12714) );
  AOI22_X1 U14995 ( .A1(n15464), .A2(n12743), .B1(n12712), .B2(n15461), .ZN(
        n12713) );
  OAI211_X1 U14996 ( .C1(n15470), .C2(n12715), .A(n12714), .B(n12713), .ZN(
        n12904) );
  INV_X1 U14997 ( .A(n12904), .ZN(n12720) );
  INV_X1 U14998 ( .A(n12715), .ZN(n12905) );
  AOI22_X1 U14999 ( .A1(n12871), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n15473), 
        .B2(n12716), .ZN(n12717) );
  OAI21_X1 U15000 ( .B1(n12974), .B2(n12867), .A(n12717), .ZN(n12718) );
  AOI21_X1 U15001 ( .B1(n12905), .B2(n15474), .A(n12718), .ZN(n12719) );
  OAI21_X1 U15002 ( .B1(n12720), .B2(n12871), .A(n12719), .ZN(P3_U3208) );
  INV_X1 U15003 ( .A(n12721), .ZN(n12722) );
  AOI21_X1 U15004 ( .B1(n12725), .B2(n12723), .A(n12722), .ZN(n12731) );
  XOR2_X1 U15005 ( .A(n12725), .B(n12724), .Z(n12726) );
  NAND2_X1 U15006 ( .A1(n12726), .A2(n15466), .ZN(n12730) );
  AOI22_X1 U15007 ( .A1(n12728), .A2(n15464), .B1(n15461), .B2(n12727), .ZN(
        n12729) );
  OAI211_X1 U15008 ( .C1(n15470), .C2(n12731), .A(n12730), .B(n12729), .ZN(
        n12908) );
  INV_X1 U15009 ( .A(n12908), .ZN(n12736) );
  INV_X1 U15010 ( .A(n12731), .ZN(n12909) );
  AOI22_X1 U15011 ( .A1(n12871), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n15473), 
        .B2(n12732), .ZN(n12733) );
  OAI21_X1 U15012 ( .B1(n12978), .B2(n12867), .A(n12733), .ZN(n12734) );
  AOI21_X1 U15013 ( .B1(n12909), .B2(n15474), .A(n12734), .ZN(n12735) );
  OAI21_X1 U15014 ( .B1(n12736), .B2(n12871), .A(n12735), .ZN(P3_U3209) );
  OR2_X1 U15015 ( .A1(n12737), .A2(n12740), .ZN(n12738) );
  NAND2_X1 U15016 ( .A1(n12739), .A2(n12738), .ZN(n12912) );
  XNOR2_X1 U15017 ( .A(n12741), .B(n12740), .ZN(n12742) );
  NAND2_X1 U15018 ( .A1(n12742), .A2(n15466), .ZN(n12745) );
  AOI22_X1 U15019 ( .A1(n15464), .A2(n12772), .B1(n12743), .B2(n15461), .ZN(
        n12744) );
  OAI211_X1 U15020 ( .C1(n15470), .C2(n12912), .A(n12745), .B(n12744), .ZN(
        n12913) );
  NAND2_X1 U15021 ( .A1(n12913), .A2(n15477), .ZN(n12751) );
  INV_X1 U15022 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n13302) );
  INV_X1 U15023 ( .A(n12746), .ZN(n12747) );
  OAI22_X1 U15024 ( .A1(n15477), .A2(n13302), .B1(n12747), .B2(n15443), .ZN(
        n12748) );
  AOI21_X1 U15025 ( .B1(n12749), .B2(n12885), .A(n12748), .ZN(n12750) );
  OAI211_X1 U15026 ( .C1(n12912), .C2(n12752), .A(n12751), .B(n12750), .ZN(
        P3_U3210) );
  XNOR2_X1 U15027 ( .A(n12753), .B(n12761), .ZN(n12757) );
  OAI22_X1 U15028 ( .A1(n12755), .A2(n15450), .B1(n12754), .B2(n15448), .ZN(
        n12756) );
  AOI21_X1 U15029 ( .B1(n12757), .B2(n15466), .A(n12756), .ZN(n12919) );
  NAND2_X1 U15030 ( .A1(n12776), .A2(n12758), .ZN(n12760) );
  NAND2_X1 U15031 ( .A1(n12760), .A2(n12759), .ZN(n12762) );
  XNOR2_X1 U15032 ( .A(n12762), .B(n12761), .ZN(n12917) );
  AOI22_X1 U15033 ( .A1(n12871), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n15473), 
        .B2(n12763), .ZN(n12764) );
  OAI21_X1 U15034 ( .B1(n12765), .B2(n12867), .A(n12764), .ZN(n12766) );
  AOI21_X1 U15035 ( .B1(n12917), .B2(n12869), .A(n12766), .ZN(n12767) );
  OAI21_X1 U15036 ( .B1(n12919), .B2(n12871), .A(n12767), .ZN(P3_U3211) );
  NAND2_X1 U15037 ( .A1(n12769), .A2(n12768), .ZN(n12770) );
  NAND2_X1 U15038 ( .A1(n12771), .A2(n12770), .ZN(n12775) );
  NAND2_X1 U15039 ( .A1(n12772), .A2(n15461), .ZN(n12773) );
  OAI21_X1 U15040 ( .B1(n12799), .B2(n15450), .A(n12773), .ZN(n12774) );
  AOI21_X1 U15041 ( .B1(n12775), .B2(n15466), .A(n12774), .ZN(n12924) );
  XNOR2_X1 U15042 ( .A(n12776), .B(n8104), .ZN(n12922) );
  INV_X1 U15043 ( .A(n12989), .ZN(n12779) );
  AOI22_X1 U15044 ( .A1(n12871), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15473), 
        .B2(n12777), .ZN(n12778) );
  OAI21_X1 U15045 ( .B1(n12779), .B2(n12867), .A(n12778), .ZN(n12780) );
  AOI21_X1 U15046 ( .B1(n12922), .B2(n12869), .A(n12780), .ZN(n12781) );
  OAI21_X1 U15047 ( .B1(n12924), .B2(n12871), .A(n12781), .ZN(P3_U3212) );
  OAI211_X1 U15048 ( .C1(n12783), .C2(n12789), .A(n12782), .B(n15466), .ZN(
        n12787) );
  AOI22_X1 U15049 ( .A1(n12785), .A2(n15461), .B1(n15464), .B2(n12784), .ZN(
        n12786) );
  NAND2_X1 U15050 ( .A1(n12787), .A2(n12786), .ZN(n12932) );
  NAND2_X1 U15051 ( .A1(n12788), .A2(n15488), .ZN(n12929) );
  NAND2_X1 U15052 ( .A1(n12790), .A2(n12789), .ZN(n12927) );
  NAND3_X1 U15053 ( .A1(n12928), .A2(n12927), .A3(n12869), .ZN(n12793) );
  AOI22_X1 U15054 ( .A1(n12871), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15473), 
        .B2(n12791), .ZN(n12792) );
  OAI211_X1 U15055 ( .C1(n12929), .C2(n12794), .A(n12793), .B(n12792), .ZN(
        n12795) );
  AOI21_X1 U15056 ( .B1(n12932), .B2(n15477), .A(n12795), .ZN(n12796) );
  INV_X1 U15057 ( .A(n12796), .ZN(P3_U3213) );
  OAI211_X1 U15058 ( .C1(n12798), .C2(n12804), .A(n12797), .B(n15466), .ZN(
        n12803) );
  OAI22_X1 U15059 ( .A1(n12800), .A2(n15450), .B1(n12799), .B2(n15448), .ZN(
        n12801) );
  INV_X1 U15060 ( .A(n12801), .ZN(n12802) );
  XNOR2_X1 U15061 ( .A(n12805), .B(n12804), .ZN(n12934) );
  AOI22_X1 U15062 ( .A1(n12871), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15473), 
        .B2(n12806), .ZN(n12807) );
  OAI21_X1 U15063 ( .B1(n12997), .B2(n12867), .A(n12807), .ZN(n12808) );
  AOI21_X1 U15064 ( .B1(n12934), .B2(n12869), .A(n12808), .ZN(n12809) );
  OAI21_X1 U15065 ( .B1(n12936), .B2(n12871), .A(n12809), .ZN(P3_U3214) );
  NAND2_X1 U15066 ( .A1(n12829), .A2(n12810), .ZN(n12813) );
  INV_X1 U15067 ( .A(n12811), .ZN(n12812) );
  AOI21_X1 U15068 ( .B1(n12814), .B2(n12813), .A(n12812), .ZN(n12815) );
  OAI222_X1 U15069 ( .A1(n15448), .A2(n12817), .B1(n15450), .B2(n12816), .C1(
        n15456), .C2(n12815), .ZN(n12939) );
  INV_X1 U15070 ( .A(n12939), .ZN(n12826) );
  AND2_X1 U15071 ( .A1(n6747), .A2(n12819), .ZN(n12820) );
  AOI21_X1 U15072 ( .B1(n12821), .B2(n12820), .A(n6665), .ZN(n12940) );
  AOI22_X1 U15073 ( .A1(n12871), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n15473), 
        .B2(n12822), .ZN(n12823) );
  OAI21_X1 U15074 ( .B1(n13001), .B2(n12867), .A(n12823), .ZN(n12824) );
  AOI21_X1 U15075 ( .B1(n12940), .B2(n12869), .A(n12824), .ZN(n12825) );
  OAI21_X1 U15076 ( .B1(n12826), .B2(n12871), .A(n12825), .ZN(P3_U3215) );
  OR2_X1 U15077 ( .A1(n12845), .A2(n12852), .ZN(n12847) );
  NAND2_X1 U15078 ( .A1(n12847), .A2(n12827), .ZN(n12832) );
  AND2_X1 U15079 ( .A1(n12829), .A2(n12828), .ZN(n12830) );
  OAI211_X1 U15080 ( .C1(n12832), .C2(n12831), .A(n12830), .B(n15466), .ZN(
        n12836) );
  AOI22_X1 U15081 ( .A1(n12834), .A2(n15461), .B1(n15464), .B2(n12833), .ZN(
        n12835) );
  NAND2_X1 U15082 ( .A1(n12836), .A2(n12835), .ZN(n12943) );
  INV_X1 U15083 ( .A(n12943), .ZN(n12844) );
  NAND2_X1 U15084 ( .A1(n12838), .A2(n12837), .ZN(n12839) );
  XNOR2_X1 U15085 ( .A(n12839), .B(n6644), .ZN(n12944) );
  AOI22_X1 U15086 ( .A1(n12871), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15473), 
        .B2(n12840), .ZN(n12841) );
  OAI21_X1 U15087 ( .B1(n13005), .B2(n12867), .A(n12841), .ZN(n12842) );
  AOI21_X1 U15088 ( .B1(n12944), .B2(n12869), .A(n12842), .ZN(n12843) );
  OAI21_X1 U15089 ( .B1(n12844), .B2(n12871), .A(n12843), .ZN(P3_U3216) );
  NAND2_X1 U15090 ( .A1(n12845), .A2(n12852), .ZN(n12846) );
  NAND3_X1 U15091 ( .A1(n12847), .A2(n15466), .A3(n12846), .ZN(n12851) );
  AOI22_X1 U15092 ( .A1(n12849), .A2(n15461), .B1(n15464), .B2(n12848), .ZN(
        n12850) );
  XNOR2_X1 U15093 ( .A(n12853), .B(n12852), .ZN(n12947) );
  AOI22_X1 U15094 ( .A1(n12871), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15473), 
        .B2(n12854), .ZN(n12855) );
  OAI21_X1 U15095 ( .B1(n12867), .B2(n12856), .A(n12855), .ZN(n12857) );
  AOI21_X1 U15096 ( .B1(n12947), .B2(n12869), .A(n12857), .ZN(n12858) );
  OAI21_X1 U15097 ( .B1(n12949), .B2(n12871), .A(n12858), .ZN(P3_U3217) );
  XOR2_X1 U15098 ( .A(n12859), .B(n12863), .Z(n12860) );
  OAI222_X1 U15099 ( .A1(n15448), .A2(n12861), .B1(n15450), .B2(n14763), .C1(
        n12860), .C2(n15456), .ZN(n12953) );
  INV_X1 U15100 ( .A(n12953), .ZN(n12872) );
  OAI21_X1 U15101 ( .B1(n12864), .B2(n12863), .A(n12862), .ZN(n12954) );
  AOI22_X1 U15102 ( .A1(n12871), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15473), 
        .B2(n12865), .ZN(n12866) );
  OAI21_X1 U15103 ( .B1(n12867), .B2(n13015), .A(n12866), .ZN(n12868) );
  AOI21_X1 U15104 ( .B1(n12954), .B2(n12869), .A(n12868), .ZN(n12870) );
  OAI21_X1 U15105 ( .B1(n12872), .B2(n12871), .A(n12870), .ZN(P3_U3218) );
  INV_X1 U15106 ( .A(n12873), .ZN(n12874) );
  AOI21_X1 U15107 ( .B1(n12877), .B2(n12875), .A(n12874), .ZN(n14791) );
  XNOR2_X1 U15108 ( .A(n12876), .B(n12877), .ZN(n12878) );
  OAI222_X1 U15109 ( .A1(n15448), .A2(n12879), .B1(n15450), .B2(n14778), .C1(
        n12878), .C2(n15456), .ZN(n14793) );
  NAND2_X1 U15110 ( .A1(n14793), .A2(n15477), .ZN(n12887) );
  INV_X1 U15111 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n12882) );
  INV_X1 U15112 ( .A(n12880), .ZN(n12881) );
  OAI22_X1 U15113 ( .A1(n15477), .A2(n12882), .B1(n12881), .B2(n15443), .ZN(
        n12883) );
  AOI21_X1 U15114 ( .B1(n12885), .B2(n12884), .A(n12883), .ZN(n12886) );
  OAI211_X1 U15115 ( .C1(n14791), .C2(n12888), .A(n12887), .B(n12886), .ZN(
        P3_U3219) );
  INV_X1 U15116 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n13324) );
  MUX2_X1 U15117 ( .A(n13324), .B(n14786), .S(n15547), .Z(n12889) );
  OAI21_X1 U15118 ( .B1(n12960), .B2(n12957), .A(n12889), .ZN(P3_U3490) );
  INV_X1 U15119 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n12893) );
  AND2_X1 U15120 ( .A1(n12890), .A2(n15497), .ZN(n12891) );
  NOR2_X1 U15121 ( .A1(n12892), .A2(n12891), .ZN(n12961) );
  INV_X1 U15122 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n12896) );
  OAI21_X1 U15123 ( .B1(n12966), .B2(n12957), .A(n12897), .ZN(P3_U3486) );
  INV_X1 U15124 ( .A(n12898), .ZN(n12970) );
  INV_X1 U15125 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12902) );
  INV_X1 U15126 ( .A(n12899), .ZN(n12901) );
  AOI21_X1 U15127 ( .B1(n15517), .B2(n12901), .A(n12900), .ZN(n12967) );
  MUX2_X1 U15128 ( .A(n12902), .B(n12967), .S(n15547), .Z(n12903) );
  OAI21_X1 U15129 ( .B1(n12970), .B2(n12957), .A(n12903), .ZN(P3_U3485) );
  INV_X1 U15130 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n12906) );
  AOI21_X1 U15131 ( .B1(n15517), .B2(n12905), .A(n12904), .ZN(n12971) );
  MUX2_X1 U15132 ( .A(n12906), .B(n12971), .S(n15547), .Z(n12907) );
  OAI21_X1 U15133 ( .B1(n12974), .B2(n12957), .A(n12907), .ZN(P3_U3484) );
  INV_X1 U15134 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12910) );
  AOI21_X1 U15135 ( .B1(n15517), .B2(n12909), .A(n12908), .ZN(n12975) );
  MUX2_X1 U15136 ( .A(n12910), .B(n12975), .S(n15547), .Z(n12911) );
  OAI21_X1 U15137 ( .B1(n12978), .B2(n12957), .A(n12911), .ZN(P3_U3483) );
  INV_X1 U15138 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12915) );
  INV_X1 U15139 ( .A(n12912), .ZN(n12914) );
  AOI21_X1 U15140 ( .B1(n15517), .B2(n12914), .A(n12913), .ZN(n12979) );
  MUX2_X1 U15141 ( .A(n12915), .B(n12979), .S(n15547), .Z(n12916) );
  OAI21_X1 U15142 ( .B1(n12982), .B2(n12957), .A(n12916), .ZN(P3_U3482) );
  NAND2_X1 U15143 ( .A1(n12917), .A2(n15497), .ZN(n12918) );
  NAND2_X1 U15144 ( .A1(n12919), .A2(n12918), .ZN(n12983) );
  MUX2_X1 U15145 ( .A(P3_REG1_REG_22__SCAN_IN), .B(n12983), .S(n15547), .Z(
        n12920) );
  AOI21_X1 U15146 ( .B1(n12951), .B2(n12985), .A(n12920), .ZN(n12921) );
  INV_X1 U15147 ( .A(n12921), .ZN(P3_U3481) );
  NAND2_X1 U15148 ( .A1(n12922), .A2(n15497), .ZN(n12923) );
  NAND2_X1 U15149 ( .A1(n12924), .A2(n12923), .ZN(n12987) );
  MUX2_X1 U15150 ( .A(P3_REG1_REG_21__SCAN_IN), .B(n12987), .S(n15547), .Z(
        n12925) );
  AOI21_X1 U15151 ( .B1(n12951), .B2(n12989), .A(n12925), .ZN(n12926) );
  INV_X1 U15152 ( .A(n12926), .ZN(P3_U3480) );
  INV_X1 U15153 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13313) );
  NAND3_X1 U15154 ( .A1(n12928), .A2(n15497), .A3(n12927), .ZN(n12930) );
  NAND2_X1 U15155 ( .A1(n12930), .A2(n12929), .ZN(n12931) );
  NOR2_X1 U15156 ( .A1(n12932), .A2(n12931), .ZN(n12991) );
  MUX2_X1 U15157 ( .A(n13313), .B(n12991), .S(n15547), .Z(n12933) );
  INV_X1 U15158 ( .A(n12933), .ZN(P3_U3479) );
  NAND2_X1 U15159 ( .A1(n12934), .A2(n15497), .ZN(n12935) );
  NAND2_X1 U15160 ( .A1(n12936), .A2(n12935), .ZN(n12994) );
  MUX2_X1 U15161 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n12994), .S(n15547), .Z(
        n12937) );
  INV_X1 U15162 ( .A(n12937), .ZN(n12938) );
  OAI21_X1 U15163 ( .B1(n12957), .B2(n12997), .A(n12938), .ZN(P3_U3478) );
  AOI21_X1 U15164 ( .B1(n12940), .B2(n15497), .A(n12939), .ZN(n12998) );
  MUX2_X1 U15165 ( .A(n12941), .B(n12998), .S(n15547), .Z(n12942) );
  OAI21_X1 U15166 ( .B1(n13001), .B2(n12957), .A(n12942), .ZN(P3_U3477) );
  AOI21_X1 U15167 ( .B1(n12944), .B2(n15497), .A(n12943), .ZN(n13002) );
  MUX2_X1 U15168 ( .A(n12945), .B(n13002), .S(n15547), .Z(n12946) );
  OAI21_X1 U15169 ( .B1(n13005), .B2(n12957), .A(n12946), .ZN(P3_U3476) );
  NAND2_X1 U15170 ( .A1(n12947), .A2(n15497), .ZN(n12948) );
  NAND2_X1 U15171 ( .A1(n12949), .A2(n12948), .ZN(n13006) );
  MUX2_X1 U15172 ( .A(n13006), .B(P3_REG1_REG_16__SCAN_IN), .S(n15544), .Z(
        n12950) );
  AOI21_X1 U15173 ( .B1(n12951), .B2(n13008), .A(n12950), .ZN(n12952) );
  INV_X1 U15174 ( .A(n12952), .ZN(P3_U3475) );
  AOI21_X1 U15175 ( .B1(n15497), .B2(n12954), .A(n12953), .ZN(n13011) );
  MUX2_X1 U15176 ( .A(n12955), .B(n13011), .S(n15547), .Z(n12956) );
  OAI21_X1 U15177 ( .B1(n13015), .B2(n12957), .A(n12956), .ZN(P3_U3474) );
  INV_X1 U15178 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n12958) );
  MUX2_X1 U15179 ( .A(n14786), .B(n12958), .S(n15526), .Z(n12959) );
  OAI21_X1 U15180 ( .B1(n12960), .B2(n13014), .A(n12959), .ZN(P3_U3458) );
  INV_X1 U15181 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n12962) );
  INV_X1 U15182 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n12965) );
  INV_X1 U15183 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12968) );
  MUX2_X1 U15184 ( .A(n12968), .B(n12967), .S(n15528), .Z(n12969) );
  OAI21_X1 U15185 ( .B1(n12970), .B2(n13014), .A(n12969), .ZN(P3_U3453) );
  INV_X1 U15186 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n12972) );
  MUX2_X1 U15187 ( .A(n12972), .B(n12971), .S(n15528), .Z(n12973) );
  OAI21_X1 U15188 ( .B1(n12974), .B2(n13014), .A(n12973), .ZN(P3_U3452) );
  INV_X1 U15189 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n12976) );
  MUX2_X1 U15190 ( .A(n12976), .B(n12975), .S(n15528), .Z(n12977) );
  OAI21_X1 U15191 ( .B1(n12978), .B2(n13014), .A(n12977), .ZN(P3_U3451) );
  INV_X1 U15192 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n12980) );
  MUX2_X1 U15193 ( .A(n12980), .B(n12979), .S(n15528), .Z(n12981) );
  OAI21_X1 U15194 ( .B1(n12982), .B2(n13014), .A(n12981), .ZN(P3_U3450) );
  MUX2_X1 U15195 ( .A(P3_REG0_REG_22__SCAN_IN), .B(n12983), .S(n15528), .Z(
        n12984) );
  AOI21_X1 U15196 ( .B1(n13009), .B2(n12985), .A(n12984), .ZN(n12986) );
  INV_X1 U15197 ( .A(n12986), .ZN(P3_U3449) );
  MUX2_X1 U15198 ( .A(P3_REG0_REG_21__SCAN_IN), .B(n12987), .S(n15528), .Z(
        n12988) );
  AOI21_X1 U15199 ( .B1(n13009), .B2(n12989), .A(n12988), .ZN(n12990) );
  INV_X1 U15200 ( .A(n12990), .ZN(P3_U3448) );
  INV_X1 U15201 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n12992) );
  MUX2_X1 U15202 ( .A(n12992), .B(n12991), .S(n15528), .Z(n12993) );
  INV_X1 U15203 ( .A(n12993), .ZN(P3_U3447) );
  MUX2_X1 U15204 ( .A(n12994), .B(P3_REG0_REG_19__SCAN_IN), .S(n15526), .Z(
        n12995) );
  INV_X1 U15205 ( .A(n12995), .ZN(n12996) );
  OAI21_X1 U15206 ( .B1(n13014), .B2(n12997), .A(n12996), .ZN(P3_U3446) );
  INV_X1 U15207 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n12999) );
  MUX2_X1 U15208 ( .A(n12999), .B(n12998), .S(n15528), .Z(n13000) );
  OAI21_X1 U15209 ( .B1(n13001), .B2(n13014), .A(n13000), .ZN(P3_U3444) );
  INV_X1 U15210 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13003) );
  MUX2_X1 U15211 ( .A(n13003), .B(n13002), .S(n15528), .Z(n13004) );
  OAI21_X1 U15212 ( .B1(n13005), .B2(n13014), .A(n13004), .ZN(P3_U3441) );
  MUX2_X1 U15213 ( .A(n13006), .B(P3_REG0_REG_16__SCAN_IN), .S(n15526), .Z(
        n13007) );
  AOI21_X1 U15214 ( .B1(n13009), .B2(n13008), .A(n13007), .ZN(n13010) );
  INV_X1 U15215 ( .A(n13010), .ZN(P3_U3438) );
  INV_X1 U15216 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13012) );
  MUX2_X1 U15217 ( .A(n13012), .B(n13011), .S(n15528), .Z(n13013) );
  OAI21_X1 U15218 ( .B1(n13015), .B2(n13014), .A(n13013), .ZN(P3_U3435) );
  MUX2_X1 U15219 ( .A(n13016), .B(P3_D_REG_1__SCAN_IN), .S(n13017), .Z(
        P3_U3377) );
  MUX2_X1 U15220 ( .A(n13018), .B(P3_D_REG_0__SCAN_IN), .S(n13017), .Z(
        P3_U3376) );
  NAND3_X1 U15221 ( .A1(n13019), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n13021) );
  OAI22_X1 U15222 ( .A1(n13022), .A2(n13021), .B1(n13020), .B2(n14721), .ZN(
        n13023) );
  AOI21_X1 U15223 ( .B1(n13024), .B2(n13381), .A(n13023), .ZN(n13025) );
  INV_X1 U15224 ( .A(n13025), .ZN(P3_U3264) );
  INV_X1 U15225 ( .A(n13026), .ZN(n13029) );
  OAI222_X1 U15226 ( .A1(n14721), .A2(n13030), .B1(n14722), .B2(n13029), .C1(
        P3_U3151), .C2(n13027), .ZN(P3_U3266) );
  OAI22_X1 U15227 ( .A1(P2_REG2_REG_20__SCAN_IN), .A2(keyinput27), .B1(
        keyinput95), .B2(P1_REG2_REG_3__SCAN_IN), .ZN(n13031) );
  AOI221_X1 U15228 ( .B1(P2_REG2_REG_20__SCAN_IN), .B2(keyinput27), .C1(
        P1_REG2_REG_3__SCAN_IN), .C2(keyinput95), .A(n13031), .ZN(n13038) );
  OAI22_X1 U15229 ( .A1(P2_D_REG_8__SCAN_IN), .A2(keyinput96), .B1(keyinput46), 
        .B2(P2_ADDR_REG_2__SCAN_IN), .ZN(n13032) );
  AOI221_X1 U15230 ( .B1(P2_D_REG_8__SCAN_IN), .B2(keyinput96), .C1(
        P2_ADDR_REG_2__SCAN_IN), .C2(keyinput46), .A(n13032), .ZN(n13037) );
  OAI22_X1 U15231 ( .A1(SI_8_), .A2(keyinput94), .B1(P1_D_REG_15__SCAN_IN), 
        .B2(keyinput41), .ZN(n13033) );
  AOI221_X1 U15232 ( .B1(SI_8_), .B2(keyinput94), .C1(keyinput41), .C2(
        P1_D_REG_15__SCAN_IN), .A(n13033), .ZN(n13036) );
  OAI22_X1 U15233 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(keyinput44), .B1(
        keyinput25), .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n13034) );
  AOI221_X1 U15234 ( .B1(P1_IR_REG_27__SCAN_IN), .B2(keyinput44), .C1(
        P3_DATAO_REG_13__SCAN_IN), .C2(keyinput25), .A(n13034), .ZN(n13035) );
  NAND4_X1 U15235 ( .A1(n13038), .A2(n13037), .A3(n13036), .A4(n13035), .ZN(
        n13066) );
  OAI22_X1 U15236 ( .A1(P2_D_REG_26__SCAN_IN), .A2(keyinput42), .B1(keyinput88), .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n13039) );
  AOI221_X1 U15237 ( .B1(P2_D_REG_26__SCAN_IN), .B2(keyinput42), .C1(
        P1_DATAO_REG_13__SCAN_IN), .C2(keyinput88), .A(n13039), .ZN(n13046) );
  OAI22_X1 U15238 ( .A1(P2_REG2_REG_26__SCAN_IN), .A2(keyinput115), .B1(
        P3_REG0_REG_4__SCAN_IN), .B2(keyinput101), .ZN(n13040) );
  AOI221_X1 U15239 ( .B1(P2_REG2_REG_26__SCAN_IN), .B2(keyinput115), .C1(
        keyinput101), .C2(P3_REG0_REG_4__SCAN_IN), .A(n13040), .ZN(n13045) );
  OAI22_X1 U15240 ( .A1(P3_D_REG_25__SCAN_IN), .A2(keyinput19), .B1(
        P3_D_REG_3__SCAN_IN), .B2(keyinput104), .ZN(n13041) );
  AOI221_X1 U15241 ( .B1(P3_D_REG_25__SCAN_IN), .B2(keyinput19), .C1(
        keyinput104), .C2(P3_D_REG_3__SCAN_IN), .A(n13041), .ZN(n13044) );
  OAI22_X1 U15242 ( .A1(P2_REG0_REG_8__SCAN_IN), .A2(keyinput91), .B1(
        keyinput9), .B2(P3_REG1_REG_7__SCAN_IN), .ZN(n13042) );
  AOI221_X1 U15243 ( .B1(P2_REG0_REG_8__SCAN_IN), .B2(keyinput91), .C1(
        P3_REG1_REG_7__SCAN_IN), .C2(keyinput9), .A(n13042), .ZN(n13043) );
  NAND4_X1 U15244 ( .A1(n13046), .A2(n13045), .A3(n13044), .A4(n13043), .ZN(
        n13065) );
  OAI22_X1 U15245 ( .A1(P3_REG3_REG_26__SCAN_IN), .A2(keyinput36), .B1(
        P1_REG2_REG_6__SCAN_IN), .B2(keyinput58), .ZN(n13047) );
  AOI221_X1 U15246 ( .B1(P3_REG3_REG_26__SCAN_IN), .B2(keyinput36), .C1(
        keyinput58), .C2(P1_REG2_REG_6__SCAN_IN), .A(n13047), .ZN(n13054) );
  OAI22_X1 U15247 ( .A1(SI_11_), .A2(keyinput122), .B1(keyinput53), .B2(
        P1_REG1_REG_21__SCAN_IN), .ZN(n13048) );
  AOI221_X1 U15248 ( .B1(SI_11_), .B2(keyinput122), .C1(
        P1_REG1_REG_21__SCAN_IN), .C2(keyinput53), .A(n13048), .ZN(n13053) );
  OAI22_X1 U15249 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput82), .B1(
        P1_REG1_REG_24__SCAN_IN), .B2(keyinput17), .ZN(n13049) );
  AOI221_X1 U15250 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput82), .C1(
        keyinput17), .C2(P1_REG1_REG_24__SCAN_IN), .A(n13049), .ZN(n13052) );
  OAI22_X1 U15251 ( .A1(P3_REG3_REG_5__SCAN_IN), .A2(keyinput113), .B1(
        keyinput110), .B2(P1_D_REG_4__SCAN_IN), .ZN(n13050) );
  AOI221_X1 U15252 ( .B1(P3_REG3_REG_5__SCAN_IN), .B2(keyinput113), .C1(
        P1_D_REG_4__SCAN_IN), .C2(keyinput110), .A(n13050), .ZN(n13051) );
  NAND4_X1 U15253 ( .A1(n13054), .A2(n13053), .A3(n13052), .A4(n13051), .ZN(
        n13064) );
  OAI22_X1 U15254 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(keyinput10), .B1(
        keyinput74), .B2(P1_D_REG_30__SCAN_IN), .ZN(n13055) );
  AOI221_X1 U15255 ( .B1(P3_REG1_REG_10__SCAN_IN), .B2(keyinput10), .C1(
        P1_D_REG_30__SCAN_IN), .C2(keyinput74), .A(n13055), .ZN(n13062) );
  OAI22_X1 U15256 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(keyinput55), .B1(
        keyinput64), .B2(P1_REG3_REG_16__SCAN_IN), .ZN(n13056) );
  AOI221_X1 U15257 ( .B1(P3_IR_REG_14__SCAN_IN), .B2(keyinput55), .C1(
        P1_REG3_REG_16__SCAN_IN), .C2(keyinput64), .A(n13056), .ZN(n13061) );
  OAI22_X1 U15258 ( .A1(P2_REG1_REG_23__SCAN_IN), .A2(keyinput8), .B1(
        P1_REG2_REG_27__SCAN_IN), .B2(keyinput39), .ZN(n13057) );
  AOI221_X1 U15259 ( .B1(P2_REG1_REG_23__SCAN_IN), .B2(keyinput8), .C1(
        keyinput39), .C2(P1_REG2_REG_27__SCAN_IN), .A(n13057), .ZN(n13060) );
  OAI22_X1 U15260 ( .A1(P3_REG2_REG_28__SCAN_IN), .A2(keyinput16), .B1(
        keyinput18), .B2(P3_REG1_REG_3__SCAN_IN), .ZN(n13058) );
  AOI221_X1 U15261 ( .B1(P3_REG2_REG_28__SCAN_IN), .B2(keyinput16), .C1(
        P3_REG1_REG_3__SCAN_IN), .C2(keyinput18), .A(n13058), .ZN(n13059) );
  NAND4_X1 U15262 ( .A1(n13062), .A2(n13061), .A3(n13060), .A4(n13059), .ZN(
        n13063) );
  NOR4_X1 U15263 ( .A1(n13066), .A2(n13065), .A3(n13064), .A4(n13063), .ZN(
        n13379) );
  AOI22_X1 U15264 ( .A1(P3_DATAO_REG_15__SCAN_IN), .A2(keyinput189), .B1(
        P1_REG1_REG_21__SCAN_IN), .B2(keyinput181), .ZN(n13067) );
  OAI221_X1 U15265 ( .B1(P3_DATAO_REG_15__SCAN_IN), .B2(keyinput189), .C1(
        P1_REG1_REG_21__SCAN_IN), .C2(keyinput181), .A(n13067), .ZN(n13074) );
  AOI22_X1 U15266 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(keyinput221), .B1(
        P3_D_REG_11__SCAN_IN), .B2(keyinput187), .ZN(n13068) );
  OAI221_X1 U15267 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(keyinput221), .C1(
        P3_D_REG_11__SCAN_IN), .C2(keyinput187), .A(n13068), .ZN(n13073) );
  AOI22_X1 U15268 ( .A1(P3_REG2_REG_28__SCAN_IN), .A2(keyinput144), .B1(
        P3_REG3_REG_5__SCAN_IN), .B2(keyinput241), .ZN(n13069) );
  OAI221_X1 U15269 ( .B1(P3_REG2_REG_28__SCAN_IN), .B2(keyinput144), .C1(
        P3_REG3_REG_5__SCAN_IN), .C2(keyinput241), .A(n13069), .ZN(n13072) );
  AOI22_X1 U15270 ( .A1(SI_1_), .A2(keyinput143), .B1(P2_IR_REG_17__SCAN_IN), 
        .B2(keyinput205), .ZN(n13070) );
  OAI221_X1 U15271 ( .B1(SI_1_), .B2(keyinput143), .C1(P2_IR_REG_17__SCAN_IN), 
        .C2(keyinput205), .A(n13070), .ZN(n13071) );
  NOR4_X1 U15272 ( .A1(n13074), .A2(n13073), .A3(n13072), .A4(n13071), .ZN(
        n13102) );
  AOI22_X1 U15273 ( .A1(P3_IR_REG_23__SCAN_IN), .A2(keyinput198), .B1(
        P2_REG0_REG_13__SCAN_IN), .B2(keyinput217), .ZN(n13075) );
  OAI221_X1 U15274 ( .B1(P3_IR_REG_23__SCAN_IN), .B2(keyinput198), .C1(
        P2_REG0_REG_13__SCAN_IN), .C2(keyinput217), .A(n13075), .ZN(n13082) );
  AOI22_X1 U15275 ( .A1(P3_ADDR_REG_10__SCAN_IN), .A2(keyinput248), .B1(
        P1_REG1_REG_0__SCAN_IN), .B2(keyinput156), .ZN(n13076) );
  OAI221_X1 U15276 ( .B1(P3_ADDR_REG_10__SCAN_IN), .B2(keyinput248), .C1(
        P1_REG1_REG_0__SCAN_IN), .C2(keyinput156), .A(n13076), .ZN(n13081) );
  AOI22_X1 U15277 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(keyinput192), .B1(
        P3_REG0_REG_11__SCAN_IN), .B2(keyinput228), .ZN(n13077) );
  OAI221_X1 U15278 ( .B1(P1_REG3_REG_16__SCAN_IN), .B2(keyinput192), .C1(
        P3_REG0_REG_11__SCAN_IN), .C2(keyinput228), .A(n13077), .ZN(n13080) );
  AOI22_X1 U15279 ( .A1(P3_REG1_REG_20__SCAN_IN), .A2(keyinput177), .B1(
        P3_REG2_REG_13__SCAN_IN), .B2(keyinput251), .ZN(n13078) );
  OAI221_X1 U15280 ( .B1(P3_REG1_REG_20__SCAN_IN), .B2(keyinput177), .C1(
        P3_REG2_REG_13__SCAN_IN), .C2(keyinput251), .A(n13078), .ZN(n13079) );
  NOR4_X1 U15281 ( .A1(n13082), .A2(n13081), .A3(n13080), .A4(n13079), .ZN(
        n13101) );
  AOI22_X1 U15282 ( .A1(P1_REG2_REG_3__SCAN_IN), .A2(keyinput223), .B1(
        P1_REG2_REG_16__SCAN_IN), .B2(keyinput131), .ZN(n13083) );
  OAI221_X1 U15283 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(keyinput223), .C1(
        P1_REG2_REG_16__SCAN_IN), .C2(keyinput131), .A(n13083), .ZN(n13090) );
  AOI22_X1 U15284 ( .A1(P3_REG0_REG_4__SCAN_IN), .A2(keyinput229), .B1(
        P2_REG2_REG_26__SCAN_IN), .B2(keyinput243), .ZN(n13084) );
  OAI221_X1 U15285 ( .B1(P3_REG0_REG_4__SCAN_IN), .B2(keyinput229), .C1(
        P2_REG2_REG_26__SCAN_IN), .C2(keyinput243), .A(n13084), .ZN(n13089) );
  AOI22_X1 U15286 ( .A1(P3_DATAO_REG_13__SCAN_IN), .A2(keyinput153), .B1(
        P2_REG2_REG_20__SCAN_IN), .B2(keyinput155), .ZN(n13085) );
  OAI221_X1 U15287 ( .B1(P3_DATAO_REG_13__SCAN_IN), .B2(keyinput153), .C1(
        P2_REG2_REG_20__SCAN_IN), .C2(keyinput155), .A(n13085), .ZN(n13088) );
  AOI22_X1 U15288 ( .A1(P1_REG0_REG_25__SCAN_IN), .A2(keyinput220), .B1(
        P3_REG0_REG_14__SCAN_IN), .B2(keyinput152), .ZN(n13086) );
  OAI221_X1 U15289 ( .B1(P1_REG0_REG_25__SCAN_IN), .B2(keyinput220), .C1(
        P3_REG0_REG_14__SCAN_IN), .C2(keyinput152), .A(n13086), .ZN(n13087) );
  NOR4_X1 U15290 ( .A1(n13090), .A2(n13089), .A3(n13088), .A4(n13087), .ZN(
        n13100) );
  AOI22_X1 U15291 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(keyinput211), .B1(
        P2_REG1_REG_17__SCAN_IN), .B2(keyinput239), .ZN(n13091) );
  OAI221_X1 U15292 ( .B1(P3_ADDR_REG_6__SCAN_IN), .B2(keyinput211), .C1(
        P2_REG1_REG_17__SCAN_IN), .C2(keyinput239), .A(n13091), .ZN(n13098) );
  AOI22_X1 U15293 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(keyinput247), .B1(
        P1_IR_REG_30__SCAN_IN), .B2(keyinput201), .ZN(n13092) );
  OAI221_X1 U15294 ( .B1(P1_REG3_REG_28__SCAN_IN), .B2(keyinput247), .C1(
        P1_IR_REG_30__SCAN_IN), .C2(keyinput201), .A(n13092), .ZN(n13097) );
  AOI22_X1 U15295 ( .A1(P1_REG1_REG_25__SCAN_IN), .A2(keyinput249), .B1(
        P2_REG1_REG_23__SCAN_IN), .B2(keyinput136), .ZN(n13093) );
  OAI221_X1 U15296 ( .B1(P1_REG1_REG_25__SCAN_IN), .B2(keyinput249), .C1(
        P2_REG1_REG_23__SCAN_IN), .C2(keyinput136), .A(n13093), .ZN(n13096) );
  AOI22_X1 U15297 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(keyinput159), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(keyinput128), .ZN(n13094) );
  OAI221_X1 U15298 ( .B1(P2_DATAO_REG_20__SCAN_IN), .B2(keyinput159), .C1(
        P2_DATAO_REG_4__SCAN_IN), .C2(keyinput128), .A(n13094), .ZN(n13095) );
  NOR4_X1 U15299 ( .A1(n13098), .A2(n13097), .A3(n13096), .A4(n13095), .ZN(
        n13099) );
  NAND4_X1 U15300 ( .A1(n13102), .A2(n13101), .A3(n13100), .A4(n13099), .ZN(
        n13233) );
  AOI22_X1 U15301 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(keyinput174), .B1(
        P1_REG2_REG_6__SCAN_IN), .B2(keyinput186), .ZN(n13103) );
  OAI221_X1 U15302 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(keyinput174), .C1(
        P1_REG2_REG_6__SCAN_IN), .C2(keyinput186), .A(n13103), .ZN(n13110) );
  AOI22_X1 U15303 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(keyinput231), .B1(
        P3_IR_REG_14__SCAN_IN), .B2(keyinput183), .ZN(n13104) );
  OAI221_X1 U15304 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(keyinput231), .C1(
        P3_IR_REG_14__SCAN_IN), .C2(keyinput183), .A(n13104), .ZN(n13109) );
  AOI22_X1 U15305 ( .A1(P3_DATAO_REG_28__SCAN_IN), .A2(keyinput134), .B1(
        P2_D_REG_21__SCAN_IN), .B2(keyinput197), .ZN(n13105) );
  OAI221_X1 U15306 ( .B1(P3_DATAO_REG_28__SCAN_IN), .B2(keyinput134), .C1(
        P2_D_REG_21__SCAN_IN), .C2(keyinput197), .A(n13105), .ZN(n13108) );
  AOI22_X1 U15307 ( .A1(P2_D_REG_25__SCAN_IN), .A2(keyinput148), .B1(
        P2_IR_REG_14__SCAN_IN), .B2(keyinput132), .ZN(n13106) );
  OAI221_X1 U15308 ( .B1(P2_D_REG_25__SCAN_IN), .B2(keyinput148), .C1(
        P2_IR_REG_14__SCAN_IN), .C2(keyinput132), .A(n13106), .ZN(n13107) );
  NOR4_X1 U15309 ( .A1(n13110), .A2(n13109), .A3(n13108), .A4(n13107), .ZN(
        n13138) );
  AOI22_X1 U15310 ( .A1(P2_REG1_REG_7__SCAN_IN), .A2(keyinput233), .B1(
        P2_D_REG_13__SCAN_IN), .B2(keyinput230), .ZN(n13111) );
  OAI221_X1 U15311 ( .B1(P2_REG1_REG_7__SCAN_IN), .B2(keyinput233), .C1(
        P2_D_REG_13__SCAN_IN), .C2(keyinput230), .A(n13111), .ZN(n13118) );
  AOI22_X1 U15312 ( .A1(P1_REG1_REG_24__SCAN_IN), .A2(keyinput145), .B1(
        P3_REG1_REG_4__SCAN_IN), .B2(keyinput165), .ZN(n13112) );
  OAI221_X1 U15313 ( .B1(P1_REG1_REG_24__SCAN_IN), .B2(keyinput145), .C1(
        P3_REG1_REG_4__SCAN_IN), .C2(keyinput165), .A(n13112), .ZN(n13117) );
  AOI22_X1 U15314 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(keyinput138), .B1(
        P2_D_REG_6__SCAN_IN), .B2(keyinput149), .ZN(n13113) );
  OAI221_X1 U15315 ( .B1(P3_REG1_REG_10__SCAN_IN), .B2(keyinput138), .C1(
        P2_D_REG_6__SCAN_IN), .C2(keyinput149), .A(n13113), .ZN(n13116) );
  AOI22_X1 U15316 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(keyinput216), .B1(
        P2_D_REG_1__SCAN_IN), .B2(keyinput135), .ZN(n13114) );
  OAI221_X1 U15317 ( .B1(P1_DATAO_REG_13__SCAN_IN), .B2(keyinput216), .C1(
        P2_D_REG_1__SCAN_IN), .C2(keyinput135), .A(n13114), .ZN(n13115) );
  NOR4_X1 U15318 ( .A1(n13118), .A2(n13117), .A3(n13116), .A4(n13115), .ZN(
        n13137) );
  AOI22_X1 U15319 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(keyinput154), .B1(
        P2_D_REG_8__SCAN_IN), .B2(keyinput224), .ZN(n13119) );
  OAI221_X1 U15320 ( .B1(P1_IR_REG_10__SCAN_IN), .B2(keyinput154), .C1(
        P2_D_REG_8__SCAN_IN), .C2(keyinput224), .A(n13119), .ZN(n13126) );
  AOI22_X1 U15321 ( .A1(P3_DATAO_REG_18__SCAN_IN), .A2(keyinput204), .B1(
        P1_REG0_REG_27__SCAN_IN), .B2(keyinput173), .ZN(n13120) );
  OAI221_X1 U15322 ( .B1(P3_DATAO_REG_18__SCAN_IN), .B2(keyinput204), .C1(
        P1_REG0_REG_27__SCAN_IN), .C2(keyinput173), .A(n13120), .ZN(n13125) );
  AOI22_X1 U15323 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(keyinput240), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(keyinput237), .ZN(n13121) );
  OAI221_X1 U15324 ( .B1(P1_DATAO_REG_7__SCAN_IN), .B2(keyinput240), .C1(
        P1_DATAO_REG_9__SCAN_IN), .C2(keyinput237), .A(n13121), .ZN(n13124) );
  AOI22_X1 U15325 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(keyinput199), .B1(SI_11_), 
        .B2(keyinput250), .ZN(n13122) );
  OAI221_X1 U15326 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(keyinput199), .C1(SI_11_), .C2(keyinput250), .A(n13122), .ZN(n13123) );
  NOR4_X1 U15327 ( .A1(n13126), .A2(n13125), .A3(n13124), .A4(n13123), .ZN(
        n13136) );
  AOI22_X1 U15328 ( .A1(P1_REG2_REG_27__SCAN_IN), .A2(keyinput167), .B1(
        P3_D_REG_10__SCAN_IN), .B2(keyinput209), .ZN(n13127) );
  OAI221_X1 U15329 ( .B1(P1_REG2_REG_27__SCAN_IN), .B2(keyinput167), .C1(
        P3_D_REG_10__SCAN_IN), .C2(keyinput209), .A(n13127), .ZN(n13134) );
  AOI22_X1 U15330 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(keyinput139), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(keyinput175), .ZN(n13128) );
  OAI221_X1 U15331 ( .B1(P1_IR_REG_26__SCAN_IN), .B2(keyinput139), .C1(
        P2_DATAO_REG_3__SCAN_IN), .C2(keyinput175), .A(n13128), .ZN(n13133) );
  AOI22_X1 U15332 ( .A1(P2_REG0_REG_8__SCAN_IN), .A2(keyinput219), .B1(
        P2_REG0_REG_19__SCAN_IN), .B2(keyinput166), .ZN(n13129) );
  OAI221_X1 U15333 ( .B1(P2_REG0_REG_8__SCAN_IN), .B2(keyinput219), .C1(
        P2_REG0_REG_19__SCAN_IN), .C2(keyinput166), .A(n13129), .ZN(n13132) );
  AOI22_X1 U15334 ( .A1(P1_REG2_REG_25__SCAN_IN), .A2(keyinput157), .B1(
        P3_REG3_REG_9__SCAN_IN), .B2(keyinput188), .ZN(n13130) );
  OAI221_X1 U15335 ( .B1(P1_REG2_REG_25__SCAN_IN), .B2(keyinput157), .C1(
        P3_REG3_REG_9__SCAN_IN), .C2(keyinput188), .A(n13130), .ZN(n13131) );
  NOR4_X1 U15336 ( .A1(n13134), .A2(n13133), .A3(n13132), .A4(n13131), .ZN(
        n13135) );
  NAND4_X1 U15337 ( .A1(n13138), .A2(n13137), .A3(n13136), .A4(n13135), .ZN(
        n13232) );
  AOI22_X1 U15338 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(keyinput163), .B1(
        P3_REG1_REG_31__SCAN_IN), .B2(keyinput225), .ZN(n13139) );
  OAI221_X1 U15339 ( .B1(P1_REG3_REG_9__SCAN_IN), .B2(keyinput163), .C1(
        P3_REG1_REG_31__SCAN_IN), .C2(keyinput225), .A(n13139), .ZN(n13146) );
  AOI22_X1 U15340 ( .A1(P1_D_REG_15__SCAN_IN), .A2(keyinput169), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(keyinput253), .ZN(n13140) );
  OAI221_X1 U15341 ( .B1(P1_D_REG_15__SCAN_IN), .B2(keyinput169), .C1(
        P2_DATAO_REG_13__SCAN_IN), .C2(keyinput253), .A(n13140), .ZN(n13145)
         );
  AOI22_X1 U15342 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(keyinput191), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(keyinput193), .ZN(n13141) );
  OAI221_X1 U15343 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(keyinput191), .C1(
        P2_DATAO_REG_0__SCAN_IN), .C2(keyinput193), .A(n13141), .ZN(n13144) );
  AOI22_X1 U15344 ( .A1(P2_REG0_REG_31__SCAN_IN), .A2(keyinput245), .B1(
        P2_D_REG_0__SCAN_IN), .B2(keyinput180), .ZN(n13142) );
  OAI221_X1 U15345 ( .B1(P2_REG0_REG_31__SCAN_IN), .B2(keyinput245), .C1(
        P2_D_REG_0__SCAN_IN), .C2(keyinput180), .A(n13142), .ZN(n13143) );
  NOR4_X1 U15346 ( .A1(n13146), .A2(n13145), .A3(n13144), .A4(n13143), .ZN(
        n13185) );
  AOI22_X1 U15347 ( .A1(P2_REG0_REG_10__SCAN_IN), .A2(keyinput171), .B1(
        P2_REG1_REG_26__SCAN_IN), .B2(keyinput160), .ZN(n13147) );
  OAI221_X1 U15348 ( .B1(P2_REG0_REG_10__SCAN_IN), .B2(keyinput171), .C1(
        P2_REG1_REG_26__SCAN_IN), .C2(keyinput160), .A(n13147), .ZN(n13157) );
  AOI22_X1 U15349 ( .A1(P1_REG0_REG_28__SCAN_IN), .A2(keyinput214), .B1(n13149), .B2(keyinput196), .ZN(n13148) );
  OAI221_X1 U15350 ( .B1(P1_REG0_REG_28__SCAN_IN), .B2(keyinput214), .C1(
        n13149), .C2(keyinput196), .A(n13148), .ZN(n13156) );
  AOI22_X1 U15351 ( .A1(n13151), .A2(keyinput185), .B1(n8844), .B2(keyinput227), .ZN(n13150) );
  OAI221_X1 U15352 ( .B1(n13151), .B2(keyinput185), .C1(n8844), .C2(
        keyinput227), .A(n13150), .ZN(n13155) );
  INV_X1 U15353 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n15131) );
  AOI22_X1 U15354 ( .A1(n13153), .A2(keyinput133), .B1(n15131), .B2(
        keyinput202), .ZN(n13152) );
  OAI221_X1 U15355 ( .B1(n13153), .B2(keyinput133), .C1(n15131), .C2(
        keyinput202), .A(n13152), .ZN(n13154) );
  NOR4_X1 U15356 ( .A1(n13157), .A2(n13156), .A3(n13155), .A4(n13154), .ZN(
        n13184) );
  AOI22_X1 U15357 ( .A1(n13159), .A2(keyinput164), .B1(keyinput140), .B2(
        n13275), .ZN(n13158) );
  OAI221_X1 U15358 ( .B1(n13159), .B2(keyinput164), .C1(n13275), .C2(
        keyinput140), .A(n13158), .ZN(n13160) );
  INV_X1 U15359 ( .A(n13160), .ZN(n13172) );
  INV_X1 U15360 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n13163) );
  INV_X1 U15361 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n13162) );
  AOI22_X1 U15362 ( .A1(n13163), .A2(keyinput203), .B1(n13162), .B2(
        keyinput129), .ZN(n13161) );
  OAI221_X1 U15363 ( .B1(n13163), .B2(keyinput203), .C1(n13162), .C2(
        keyinput129), .A(n13161), .ZN(n13164) );
  INV_X1 U15364 ( .A(n13164), .ZN(n13171) );
  XNOR2_X1 U15365 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(keyinput212), .ZN(n13167)
         );
  XNOR2_X1 U15366 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput208), .ZN(n13166) );
  XNOR2_X1 U15367 ( .A(keyinput146), .B(P3_REG1_REG_3__SCAN_IN), .ZN(n13165)
         );
  AND3_X1 U15368 ( .A1(n13167), .A2(n13166), .A3(n13165), .ZN(n13170) );
  INV_X1 U15369 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n15132) );
  INV_X1 U15370 ( .A(keyinput194), .ZN(n13168) );
  XNOR2_X1 U15371 ( .A(n15132), .B(n13168), .ZN(n13169) );
  AND4_X1 U15372 ( .A1(n13172), .A2(n13171), .A3(n13170), .A4(n13169), .ZN(
        n13183) );
  INV_X1 U15373 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n15148) );
  AOI22_X1 U15374 ( .A1(n10691), .A2(keyinput252), .B1(keyinput182), .B2(
        n15148), .ZN(n13173) );
  OAI221_X1 U15375 ( .B1(n10691), .B2(keyinput252), .C1(n15148), .C2(
        keyinput182), .A(n13173), .ZN(n13181) );
  AOI22_X1 U15376 ( .A1(n7695), .A2(keyinput190), .B1(keyinput200), .B2(n10022), .ZN(n13174) );
  OAI221_X1 U15377 ( .B1(n7695), .B2(keyinput190), .C1(n10022), .C2(
        keyinput200), .A(n13174), .ZN(n13180) );
  XOR2_X1 U15378 ( .A(n9943), .B(keyinput161), .Z(n13178) );
  XOR2_X1 U15379 ( .A(n15540), .B(keyinput137), .Z(n13177) );
  XNOR2_X1 U15380 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput234), .ZN(n13176) );
  XNOR2_X1 U15381 ( .A(SI_8_), .B(keyinput222), .ZN(n13175) );
  NAND4_X1 U15382 ( .A1(n13178), .A2(n13177), .A3(n13176), .A4(n13175), .ZN(
        n13179) );
  NOR3_X1 U15383 ( .A1(n13181), .A2(n13180), .A3(n13179), .ZN(n13182) );
  NAND4_X1 U15384 ( .A1(n13185), .A2(n13184), .A3(n13183), .A4(n13182), .ZN(
        n13231) );
  INV_X1 U15385 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n13288) );
  INV_X1 U15386 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n13187) );
  AOI22_X1 U15387 ( .A1(n13288), .A2(keyinput130), .B1(n13187), .B2(
        keyinput184), .ZN(n13186) );
  OAI221_X1 U15388 ( .B1(n13288), .B2(keyinput130), .C1(n13187), .C2(
        keyinput184), .A(n13186), .ZN(n13196) );
  AOI22_X1 U15389 ( .A1(n9687), .A2(keyinput195), .B1(n13189), .B2(keyinput210), .ZN(n13188) );
  OAI221_X1 U15390 ( .B1(n9687), .B2(keyinput195), .C1(n13189), .C2(
        keyinput210), .A(n13188), .ZN(n13195) );
  XOR2_X1 U15391 ( .A(n13312), .B(keyinput254), .Z(n13192) );
  XNOR2_X1 U15392 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput151), .ZN(n13191) );
  XNOR2_X1 U15393 ( .A(P2_IR_REG_2__SCAN_IN), .B(keyinput150), .ZN(n13190) );
  NAND3_X1 U15394 ( .A1(n13192), .A2(n13191), .A3(n13190), .ZN(n13194) );
  XNOR2_X1 U15395 ( .A(n15026), .B(keyinput255), .ZN(n13193) );
  NOR4_X1 U15396 ( .A1(n13196), .A2(n13195), .A3(n13194), .A4(n13193), .ZN(
        n13229) );
  AOI22_X1 U15397 ( .A1(n9728), .A2(keyinput226), .B1(keyinput246), .B2(n13247), .ZN(n13197) );
  OAI221_X1 U15398 ( .B1(n9728), .B2(keyinput226), .C1(n13247), .C2(
        keyinput246), .A(n13197), .ZN(n13205) );
  INV_X1 U15399 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n15134) );
  INV_X1 U15400 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n15296) );
  AOI22_X1 U15401 ( .A1(n15134), .A2(keyinput162), .B1(n15296), .B2(
        keyinput178), .ZN(n13198) );
  OAI221_X1 U15402 ( .B1(n15134), .B2(keyinput162), .C1(n15296), .C2(
        keyinput178), .A(n13198), .ZN(n13204) );
  INV_X1 U15403 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n15141) );
  AOI22_X1 U15404 ( .A1(n15141), .A2(keyinput179), .B1(n13302), .B2(
        keyinput168), .ZN(n13199) );
  OAI221_X1 U15405 ( .B1(n15141), .B2(keyinput179), .C1(n13302), .C2(
        keyinput168), .A(n13199), .ZN(n13203) );
  XNOR2_X1 U15406 ( .A(P2_IR_REG_20__SCAN_IN), .B(keyinput235), .ZN(n13201) );
  XNOR2_X1 U15407 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(keyinput215), .ZN(n13200)
         );
  NAND2_X1 U15408 ( .A1(n13201), .A2(n13200), .ZN(n13202) );
  NOR4_X1 U15409 ( .A1(n13205), .A2(n13204), .A3(n13203), .A4(n13202), .ZN(
        n13228) );
  INV_X1 U15410 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n15294) );
  AOI22_X1 U15411 ( .A1(n15294), .A2(keyinput170), .B1(keyinput176), .B2(
        n14367), .ZN(n13206) );
  OAI221_X1 U15412 ( .B1(n15294), .B2(keyinput170), .C1(n14367), .C2(
        keyinput176), .A(n13206), .ZN(n13215) );
  AOI22_X1 U15413 ( .A1(n13208), .A2(keyinput232), .B1(keyinput244), .B2(
        n10162), .ZN(n13207) );
  OAI221_X1 U15414 ( .B1(n13208), .B2(keyinput232), .C1(n10162), .C2(
        keyinput244), .A(n13207), .ZN(n13214) );
  INV_X1 U15415 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n15157) );
  AOI22_X1 U15416 ( .A1(n11492), .A2(keyinput242), .B1(keyinput238), .B2(
        n15157), .ZN(n13209) );
  OAI221_X1 U15417 ( .B1(n11492), .B2(keyinput242), .C1(n15157), .C2(
        keyinput238), .A(n13209), .ZN(n13213) );
  XNOR2_X1 U15418 ( .A(P3_REG0_REG_25__SCAN_IN), .B(keyinput141), .ZN(n13211)
         );
  XNOR2_X1 U15419 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput172), .ZN(n13210) );
  NAND2_X1 U15420 ( .A1(n13211), .A2(n13210), .ZN(n13212) );
  NOR4_X1 U15421 ( .A1(n13215), .A2(n13214), .A3(n13213), .A4(n13212), .ZN(
        n13227) );
  INV_X1 U15422 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n13267) );
  AOI22_X1 U15423 ( .A1(n13261), .A2(keyinput142), .B1(keyinput213), .B2(
        n13267), .ZN(n13216) );
  OAI221_X1 U15424 ( .B1(n13261), .B2(keyinput142), .C1(n13267), .C2(
        keyinput213), .A(n13216), .ZN(n13225) );
  XNOR2_X1 U15425 ( .A(n13297), .B(keyinput218), .ZN(n13224) );
  XNOR2_X1 U15426 ( .A(n13217), .B(keyinput147), .ZN(n13223) );
  XNOR2_X1 U15427 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput158), .ZN(n13221)
         );
  XNOR2_X1 U15428 ( .A(P3_IR_REG_7__SCAN_IN), .B(keyinput207), .ZN(n13220) );
  XNOR2_X1 U15429 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput206), .ZN(n13219)
         );
  XNOR2_X1 U15430 ( .A(keyinput236), .B(P1_REG2_REG_11__SCAN_IN), .ZN(n13218)
         );
  NAND4_X1 U15431 ( .A1(n13221), .A2(n13220), .A3(n13219), .A4(n13218), .ZN(
        n13222) );
  NOR4_X1 U15432 ( .A1(n13225), .A2(n13224), .A3(n13223), .A4(n13222), .ZN(
        n13226) );
  NAND4_X1 U15433 ( .A1(n13229), .A2(n13228), .A3(n13227), .A4(n13226), .ZN(
        n13230) );
  NOR4_X1 U15434 ( .A1(n13233), .A2(n13232), .A3(n13231), .A4(n13230), .ZN(
        n13340) );
  INV_X1 U15435 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14815) );
  AOI22_X1 U15436 ( .A1(n14863), .A2(keyinput111), .B1(keyinput100), .B2(
        n14815), .ZN(n13234) );
  OAI221_X1 U15437 ( .B1(n14863), .B2(keyinput111), .C1(n14815), .C2(
        keyinput100), .A(n13234), .ZN(n13244) );
  INV_X1 U15438 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n13236) );
  AOI22_X1 U15439 ( .A1(n13237), .A2(keyinput38), .B1(keyinput29), .B2(n13236), 
        .ZN(n13235) );
  OAI221_X1 U15440 ( .B1(n13237), .B2(keyinput38), .C1(n13236), .C2(keyinput29), .A(n13235), .ZN(n13243) );
  XOR2_X1 U15441 ( .A(P1_REG2_REG_11__SCAN_IN), .B(keyinput108), .Z(n13241) );
  XNOR2_X1 U15442 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput80), .ZN(n13240) );
  XNOR2_X1 U15443 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(keyinput112), .ZN(n13239)
         );
  XNOR2_X1 U15444 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(keyinput84), .ZN(n13238)
         );
  NAND4_X1 U15445 ( .A1(n13241), .A2(n13240), .A3(n13239), .A4(n13238), .ZN(
        n13242) );
  NOR3_X1 U15446 ( .A1(n13244), .A2(n13243), .A3(n13242), .ZN(n13286) );
  AOI22_X1 U15447 ( .A1(n11492), .A2(keyinput114), .B1(keyinput51), .B2(n15141), .ZN(n13245) );
  OAI221_X1 U15448 ( .B1(n11492), .B2(keyinput114), .C1(n15141), .C2(
        keyinput51), .A(n13245), .ZN(n13255) );
  INV_X1 U15449 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n13248) );
  AOI22_X1 U15450 ( .A1(n13248), .A2(keyinput121), .B1(keyinput118), .B2(
        n13247), .ZN(n13246) );
  OAI221_X1 U15451 ( .B1(n13248), .B2(keyinput121), .C1(n13247), .C2(
        keyinput118), .A(n13246), .ZN(n13254) );
  INV_X1 U15452 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n15376) );
  XOR2_X1 U15453 ( .A(n15376), .B(keyinput43), .Z(n13252) );
  XNOR2_X1 U15454 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput11), .ZN(n13251) );
  XNOR2_X1 U15455 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput106), .ZN(n13250) );
  XNOR2_X1 U15456 ( .A(P2_REG1_REG_26__SCAN_IN), .B(keyinput32), .ZN(n13249)
         );
  NAND4_X1 U15457 ( .A1(n13252), .A2(n13251), .A3(n13250), .A4(n13249), .ZN(
        n13253) );
  NOR3_X1 U15458 ( .A1(n13255), .A2(n13254), .A3(n13253), .ZN(n13285) );
  XNOR2_X1 U15459 ( .A(n13256), .B(keyinput70), .ZN(n13260) );
  XNOR2_X1 U15460 ( .A(n13257), .B(keyinput78), .ZN(n13259) );
  XNOR2_X1 U15461 ( .A(keyinput116), .B(n10162), .ZN(n13258) );
  NOR3_X1 U15462 ( .A1(n13260), .A2(n13259), .A3(n13258), .ZN(n13264) );
  XOR2_X1 U15463 ( .A(n13261), .B(keyinput14), .Z(n13263) );
  XNOR2_X1 U15464 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(keyinput109), .ZN(n13262)
         );
  NAND3_X1 U15465 ( .A1(n13264), .A2(n13263), .A3(n13262), .ZN(n13271) );
  AOI22_X1 U15466 ( .A1(n13267), .A2(keyinput85), .B1(keyinput83), .B2(n13266), 
        .ZN(n13265) );
  OAI221_X1 U15467 ( .B1(n13267), .B2(keyinput85), .C1(n13266), .C2(keyinput83), .A(n13265), .ZN(n13270) );
  XNOR2_X1 U15468 ( .A(n13268), .B(keyinput76), .ZN(n13269) );
  NOR3_X1 U15469 ( .A1(n13271), .A2(n13270), .A3(n13269), .ZN(n13284) );
  AOI22_X1 U15470 ( .A1(n9728), .A2(keyinput98), .B1(n15132), .B2(keyinput66), 
        .ZN(n13272) );
  OAI221_X1 U15471 ( .B1(n9728), .B2(keyinput98), .C1(n15132), .C2(keyinput66), 
        .A(n13272), .ZN(n13282) );
  INV_X1 U15472 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n13274) );
  AOI22_X1 U15473 ( .A1(n13275), .A2(keyinput12), .B1(keyinput45), .B2(n13274), 
        .ZN(n13273) );
  OAI221_X1 U15474 ( .B1(n13275), .B2(keyinput12), .C1(n13274), .C2(keyinput45), .A(n13273), .ZN(n13281) );
  INV_X1 U15475 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n15295) );
  AOI22_X1 U15476 ( .A1(n15295), .A2(keyinput69), .B1(n15299), .B2(keyinput52), 
        .ZN(n13276) );
  OAI221_X1 U15477 ( .B1(n15295), .B2(keyinput69), .C1(n15299), .C2(keyinput52), .A(n13276), .ZN(n13280) );
  AOI22_X1 U15478 ( .A1(n9523), .A2(keyinput105), .B1(n13278), .B2(keyinput87), 
        .ZN(n13277) );
  OAI221_X1 U15479 ( .B1(n9523), .B2(keyinput105), .C1(n13278), .C2(keyinput87), .A(n13277), .ZN(n13279) );
  NOR4_X1 U15480 ( .A1(n13282), .A2(n13281), .A3(n13280), .A4(n13279), .ZN(
        n13283) );
  NAND4_X1 U15481 ( .A1(n13286), .A2(n13285), .A3(n13284), .A4(n13283), .ZN(
        n13339) );
  INV_X1 U15482 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n13289) );
  AOI22_X1 U15483 ( .A1(n13289), .A2(keyinput35), .B1(keyinput2), .B2(n13288), 
        .ZN(n13287) );
  OAI221_X1 U15484 ( .B1(n13289), .B2(keyinput35), .C1(n13288), .C2(keyinput2), 
        .A(n13287), .ZN(n13300) );
  INV_X1 U15485 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15534) );
  AOI22_X1 U15486 ( .A1(n15534), .A2(keyinput37), .B1(n13291), .B2(keyinput31), 
        .ZN(n13290) );
  OAI221_X1 U15487 ( .B1(n15534), .B2(keyinput37), .C1(n13291), .C2(keyinput31), .A(n13290), .ZN(n13295) );
  INV_X1 U15488 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n14686) );
  XNOR2_X1 U15489 ( .A(n14686), .B(keyinput73), .ZN(n13294) );
  XNOR2_X1 U15490 ( .A(n13292), .B(keyinput59), .ZN(n13293) );
  OR3_X1 U15491 ( .A1(n13295), .A2(n13294), .A3(n13293), .ZN(n13299) );
  AOI22_X1 U15492 ( .A1(n15134), .A2(keyinput34), .B1(keyinput90), .B2(n13297), 
        .ZN(n13296) );
  OAI221_X1 U15493 ( .B1(n15134), .B2(keyinput34), .C1(n13297), .C2(keyinput90), .A(n13296), .ZN(n13298) );
  NOR3_X1 U15494 ( .A1(n13300), .A2(n13299), .A3(n13298), .ZN(n13337) );
  AOI22_X1 U15495 ( .A1(n13302), .A2(keyinput40), .B1(keyinput71), .B2(n14310), 
        .ZN(n13301) );
  OAI221_X1 U15496 ( .B1(n13302), .B2(keyinput40), .C1(n14310), .C2(keyinput71), .A(n13301), .ZN(n13310) );
  AOI22_X1 U15497 ( .A1(n9687), .A2(keyinput67), .B1(keyinput62), .B2(n7695), 
        .ZN(n13303) );
  OAI221_X1 U15498 ( .B1(n9687), .B2(keyinput67), .C1(n7695), .C2(keyinput62), 
        .A(n13303), .ZN(n13309) );
  XOR2_X1 U15499 ( .A(n8729), .B(keyinput89), .Z(n13307) );
  XNOR2_X1 U15500 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(keyinput47), .ZN(n13306)
         );
  XNOR2_X1 U15501 ( .A(P1_REG0_REG_28__SCAN_IN), .B(keyinput86), .ZN(n13305)
         );
  XNOR2_X1 U15502 ( .A(P2_IR_REG_20__SCAN_IN), .B(keyinput107), .ZN(n13304) );
  NAND4_X1 U15503 ( .A1(n13307), .A2(n13306), .A3(n13305), .A4(n13304), .ZN(
        n13308) );
  NOR3_X1 U15504 ( .A1(n13310), .A2(n13309), .A3(n13308), .ZN(n13336) );
  AOI22_X1 U15505 ( .A1(n13313), .A2(keyinput49), .B1(n13312), .B2(keyinput126), .ZN(n13311) );
  OAI221_X1 U15506 ( .B1(n13313), .B2(keyinput49), .C1(n13312), .C2(
        keyinput126), .A(n13311), .ZN(n13322) );
  AOI22_X1 U15507 ( .A1(n15148), .A2(keyinput54), .B1(n13315), .B2(keyinput26), 
        .ZN(n13314) );
  OAI221_X1 U15508 ( .B1(n15148), .B2(keyinput54), .C1(n13315), .C2(keyinput26), .A(n13314), .ZN(n13321) );
  XOR2_X1 U15509 ( .A(n15552), .B(keyinput63), .Z(n13318) );
  XNOR2_X1 U15510 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput23), .ZN(n13317) );
  XNOR2_X1 U15511 ( .A(SI_1_), .B(keyinput15), .ZN(n13316) );
  NAND3_X1 U15512 ( .A1(n13318), .A2(n13317), .A3(n13316), .ZN(n13320) );
  INV_X1 U15513 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n15420) );
  XNOR2_X1 U15514 ( .A(n15420), .B(keyinput120), .ZN(n13319) );
  NOR4_X1 U15515 ( .A1(n13322), .A2(n13321), .A3(n13320), .A4(n13319), .ZN(
        n13335) );
  INV_X1 U15516 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n15297) );
  AOI22_X1 U15517 ( .A1(n13324), .A2(keyinput97), .B1(n15297), .B2(keyinput21), 
        .ZN(n13323) );
  OAI221_X1 U15518 ( .B1(n13324), .B2(keyinput97), .C1(n15297), .C2(keyinput21), .A(n13323), .ZN(n13333) );
  AOI22_X1 U15519 ( .A1(n14367), .A2(keyinput48), .B1(n13326), .B2(keyinput60), 
        .ZN(n13325) );
  OAI221_X1 U15520 ( .B1(n14367), .B2(keyinput48), .C1(n13326), .C2(keyinput60), .A(n13325), .ZN(n13332) );
  XNOR2_X1 U15521 ( .A(P2_IR_REG_14__SCAN_IN), .B(keyinput4), .ZN(n13330) );
  XNOR2_X1 U15522 ( .A(P3_REG2_REG_31__SCAN_IN), .B(keyinput1), .ZN(n13329) );
  XNOR2_X1 U15523 ( .A(P3_IR_REG_7__SCAN_IN), .B(keyinput79), .ZN(n13328) );
  XNOR2_X1 U15524 ( .A(P1_REG3_REG_24__SCAN_IN), .B(keyinput93), .ZN(n13327)
         );
  NAND4_X1 U15525 ( .A1(n13330), .A2(n13329), .A3(n13328), .A4(n13327), .ZN(
        n13331) );
  NOR3_X1 U15526 ( .A1(n13333), .A2(n13332), .A3(n13331), .ZN(n13334) );
  NAND4_X1 U15527 ( .A1(n13337), .A2(n13336), .A3(n13335), .A4(n13334), .ZN(
        n13338) );
  NOR3_X1 U15528 ( .A1(n13340), .A2(n13339), .A3(n13338), .ZN(n13378) );
  OAI22_X1 U15529 ( .A1(P2_D_REG_13__SCAN_IN), .A2(keyinput102), .B1(
        P3_REG2_REG_8__SCAN_IN), .B2(keyinput103), .ZN(n13341) );
  AOI221_X1 U15530 ( .B1(P2_D_REG_13__SCAN_IN), .B2(keyinput102), .C1(
        keyinput103), .C2(P3_REG2_REG_8__SCAN_IN), .A(n13341), .ZN(n13348) );
  OAI22_X1 U15531 ( .A1(P2_D_REG_1__SCAN_IN), .A2(keyinput7), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(keyinput68), .ZN(n13342) );
  AOI221_X1 U15532 ( .B1(P2_D_REG_1__SCAN_IN), .B2(keyinput7), .C1(keyinput68), 
        .C2(P2_DATAO_REG_9__SCAN_IN), .A(n13342), .ZN(n13347) );
  OAI22_X1 U15533 ( .A1(P3_REG0_REG_25__SCAN_IN), .A2(keyinput13), .B1(
        keyinput33), .B2(P1_REG3_REG_3__SCAN_IN), .ZN(n13343) );
  AOI221_X1 U15534 ( .B1(P3_REG0_REG_25__SCAN_IN), .B2(keyinput13), .C1(
        P1_REG3_REG_3__SCAN_IN), .C2(keyinput33), .A(n13343), .ZN(n13346) );
  OAI22_X1 U15535 ( .A1(P2_D_REG_25__SCAN_IN), .A2(keyinput20), .B1(keyinput28), .B2(P1_REG1_REG_0__SCAN_IN), .ZN(n13344) );
  AOI221_X1 U15536 ( .B1(P2_D_REG_25__SCAN_IN), .B2(keyinput20), .C1(
        P1_REG1_REG_0__SCAN_IN), .C2(keyinput28), .A(n13344), .ZN(n13345) );
  NAND4_X1 U15537 ( .A1(n13348), .A2(n13347), .A3(n13346), .A4(n13345), .ZN(
        n13376) );
  OAI22_X1 U15538 ( .A1(P2_D_REG_18__SCAN_IN), .A2(keyinput50), .B1(keyinput56), .B2(P3_REG1_REG_29__SCAN_IN), .ZN(n13349) );
  AOI221_X1 U15539 ( .B1(P2_D_REG_18__SCAN_IN), .B2(keyinput50), .C1(
        P3_REG1_REG_29__SCAN_IN), .C2(keyinput56), .A(n13349), .ZN(n13356) );
  OAI22_X1 U15540 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(keyinput99), .B1(
        keyinput127), .B2(P1_ADDR_REG_13__SCAN_IN), .ZN(n13350) );
  AOI221_X1 U15541 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(keyinput99), .C1(
        P1_ADDR_REG_13__SCAN_IN), .C2(keyinput127), .A(n13350), .ZN(n13355) );
  OAI22_X1 U15542 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(keyinput65), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(keyinput72), .ZN(n13351) );
  AOI221_X1 U15543 ( .B1(P2_DATAO_REG_0__SCAN_IN), .B2(keyinput65), .C1(
        keyinput72), .C2(P3_REG3_REG_2__SCAN_IN), .A(n13351), .ZN(n13354) );
  OAI22_X1 U15544 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(keyinput75), .B1(keyinput6), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n13352) );
  AOI221_X1 U15545 ( .B1(P1_IR_REG_8__SCAN_IN), .B2(keyinput75), .C1(
        P3_DATAO_REG_28__SCAN_IN), .C2(keyinput6), .A(n13352), .ZN(n13353) );
  NAND4_X1 U15546 ( .A1(n13356), .A2(n13355), .A3(n13354), .A4(n13353), .ZN(
        n13375) );
  OAI22_X1 U15547 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(keyinput77), .B1(
        keyinput123), .B2(P3_REG2_REG_13__SCAN_IN), .ZN(n13357) );
  AOI221_X1 U15548 ( .B1(P2_IR_REG_17__SCAN_IN), .B2(keyinput77), .C1(
        P3_REG2_REG_13__SCAN_IN), .C2(keyinput123), .A(n13357), .ZN(n13364) );
  OAI22_X1 U15549 ( .A1(P3_REG0_REG_14__SCAN_IN), .A2(keyinput24), .B1(
        keyinput117), .B2(P2_REG0_REG_31__SCAN_IN), .ZN(n13358) );
  AOI221_X1 U15550 ( .B1(P3_REG0_REG_14__SCAN_IN), .B2(keyinput24), .C1(
        P2_REG0_REG_31__SCAN_IN), .C2(keyinput117), .A(n13358), .ZN(n13363) );
  OAI22_X1 U15551 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(keyinput3), .B1(
        keyinput5), .B2(P3_ADDR_REG_16__SCAN_IN), .ZN(n13359) );
  AOI221_X1 U15552 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(keyinput3), .C1(
        P3_ADDR_REG_16__SCAN_IN), .C2(keyinput5), .A(n13359), .ZN(n13362) );
  OAI22_X1 U15553 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(keyinput124), .B1(
        P1_REG0_REG_25__SCAN_IN), .B2(keyinput92), .ZN(n13360) );
  AOI221_X1 U15554 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(keyinput124), .C1(
        keyinput92), .C2(P1_REG0_REG_25__SCAN_IN), .A(n13360), .ZN(n13361) );
  NAND4_X1 U15555 ( .A1(n13364), .A2(n13363), .A3(n13362), .A4(n13361), .ZN(
        n13374) );
  OAI22_X1 U15556 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(keyinput22), .B1(keyinput81), .B2(P3_D_REG_10__SCAN_IN), .ZN(n13365) );
  AOI221_X1 U15557 ( .B1(P2_IR_REG_2__SCAN_IN), .B2(keyinput22), .C1(
        P3_D_REG_10__SCAN_IN), .C2(keyinput81), .A(n13365), .ZN(n13372) );
  OAI22_X1 U15558 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput30), .B1(
        P3_D_REG_2__SCAN_IN), .B2(keyinput57), .ZN(n13366) );
  AOI221_X1 U15559 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput30), .C1(
        keyinput57), .C2(P3_D_REG_2__SCAN_IN), .A(n13366), .ZN(n13371) );
  OAI22_X1 U15560 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(keyinput125), .B1(
        keyinput0), .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n13367) );
  AOI221_X1 U15561 ( .B1(P2_DATAO_REG_13__SCAN_IN), .B2(keyinput125), .C1(
        P2_DATAO_REG_4__SCAN_IN), .C2(keyinput0), .A(n13367), .ZN(n13370) );
  OAI22_X1 U15562 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(keyinput119), .B1(
        P3_DATAO_REG_15__SCAN_IN), .B2(keyinput61), .ZN(n13368) );
  AOI221_X1 U15563 ( .B1(P1_REG3_REG_28__SCAN_IN), .B2(keyinput119), .C1(
        keyinput61), .C2(P3_DATAO_REG_15__SCAN_IN), .A(n13368), .ZN(n13369) );
  NAND4_X1 U15564 ( .A1(n13372), .A2(n13371), .A3(n13370), .A4(n13369), .ZN(
        n13373) );
  NOR4_X1 U15565 ( .A1(n13376), .A2(n13375), .A3(n13374), .A4(n13373), .ZN(
        n13377) );
  NAND3_X1 U15566 ( .A1(n13379), .A2(n13378), .A3(n13377), .ZN(n13384) );
  AOI222_X1 U15567 ( .A1(n13382), .A2(n13381), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10150), .C1(SI_3_), .C2(n13380), .ZN(n13383) );
  XOR2_X1 U15568 ( .A(n13384), .B(n13383), .Z(P3_U3292) );
  XNOR2_X1 U15569 ( .A(n13386), .B(n13385), .ZN(n13394) );
  INV_X1 U15570 ( .A(n13598), .ZN(n13391) );
  NAND2_X1 U15571 ( .A1(n13475), .A2(n13509), .ZN(n13389) );
  OR2_X1 U15572 ( .A1(n13492), .A2(n13387), .ZN(n13388) );
  NAND2_X1 U15573 ( .A1(n13389), .A2(n13388), .ZN(n13594) );
  AOI22_X1 U15574 ( .A1(n13496), .A2(n13594), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13390) );
  OAI21_X1 U15575 ( .B1(n13391), .B2(n13498), .A(n13390), .ZN(n13392) );
  AOI21_X1 U15576 ( .B1(n13773), .B2(n13501), .A(n13392), .ZN(n13393) );
  OAI21_X1 U15577 ( .B1(n13394), .B2(n13503), .A(n13393), .ZN(P2_U3186) );
  OAI21_X1 U15578 ( .B1(n13396), .B2(n13395), .A(n13448), .ZN(n13397) );
  NAND2_X1 U15579 ( .A1(n13397), .A2(n13454), .ZN(n13403) );
  OAI22_X1 U15580 ( .A1(n13399), .A2(n13495), .B1(n13398), .B2(n13492), .ZN(
        n13652) );
  INV_X1 U15581 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13400) );
  OAI22_X1 U15582 ( .A1(n13498), .A2(n13654), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13400), .ZN(n13401) );
  AOI21_X1 U15583 ( .B1(n13652), .B2(n13496), .A(n13401), .ZN(n13402) );
  OAI211_X1 U15584 ( .C1(n7316), .C2(n13461), .A(n13403), .B(n13402), .ZN(
        P2_U3188) );
  NOR2_X1 U15585 ( .A1(n13404), .A2(n6781), .ZN(n13405) );
  XNOR2_X1 U15586 ( .A(n13406), .B(n13405), .ZN(n13411) );
  AOI22_X1 U15587 ( .A1(n13515), .A2(n13474), .B1(n13475), .B2(n13517), .ZN(
        n13714) );
  NAND2_X1 U15588 ( .A1(n13467), .A2(n13718), .ZN(n13408) );
  OAI211_X1 U15589 ( .C1(n13714), .C2(n13476), .A(n13408), .B(n13407), .ZN(
        n13409) );
  AOI21_X1 U15590 ( .B1(n13818), .B2(n13501), .A(n13409), .ZN(n13410) );
  OAI21_X1 U15591 ( .B1(n13411), .B2(n13503), .A(n13410), .ZN(P2_U3191) );
  XNOR2_X1 U15592 ( .A(n13413), .B(n13412), .ZN(n13418) );
  AND2_X1 U15593 ( .A1(n13515), .A2(n13475), .ZN(n13414) );
  AOI21_X1 U15594 ( .B1(n13513), .B2(n13474), .A(n13414), .ZN(n13690) );
  AOI22_X1 U15595 ( .A1(n13682), .A2(n13467), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13415) );
  OAI21_X1 U15596 ( .B1(n13690), .B2(n13476), .A(n13415), .ZN(n13416) );
  AOI21_X1 U15597 ( .B1(n13804), .B2(n13501), .A(n13416), .ZN(n13417) );
  OAI21_X1 U15598 ( .B1(n13418), .B2(n13503), .A(n13417), .ZN(P2_U3195) );
  XNOR2_X1 U15599 ( .A(n13420), .B(n13419), .ZN(n13428) );
  INV_X1 U15600 ( .A(n13631), .ZN(n13425) );
  NAND2_X1 U15601 ( .A1(n13475), .A2(n13511), .ZN(n13423) );
  OR2_X1 U15602 ( .A1(n13421), .A2(n13492), .ZN(n13422) );
  NAND2_X1 U15603 ( .A1(n13423), .A2(n13422), .ZN(n13623) );
  AOI22_X1 U15604 ( .A1(n13496), .A2(n13623), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13424) );
  OAI21_X1 U15605 ( .B1(n13425), .B2(n13498), .A(n13424), .ZN(n13426) );
  AOI21_X1 U15606 ( .B1(n13785), .B2(n13501), .A(n13426), .ZN(n13427) );
  OAI21_X1 U15607 ( .B1(n13428), .B2(n13503), .A(n13427), .ZN(P2_U3197) );
  OAI21_X1 U15608 ( .B1(n13431), .B2(n13430), .A(n13429), .ZN(n13432) );
  NAND2_X1 U15609 ( .A1(n13432), .A2(n13454), .ZN(n13437) );
  INV_X1 U15610 ( .A(n13747), .ZN(n13435) );
  AOI22_X1 U15611 ( .A1(n13518), .A2(n13474), .B1(n13475), .B2(n13520), .ZN(
        n13744) );
  OAI21_X1 U15612 ( .B1(n13744), .B2(n13476), .A(n13433), .ZN(n13434) );
  AOI21_X1 U15613 ( .B1(n13435), .B2(n13467), .A(n13434), .ZN(n13436) );
  OAI211_X1 U15614 ( .C1(n14868), .C2(n13461), .A(n13437), .B(n13436), .ZN(
        P2_U3198) );
  OAI21_X1 U15615 ( .B1(n13440), .B2(n13439), .A(n13438), .ZN(n13441) );
  NAND2_X1 U15616 ( .A1(n13441), .A2(n13454), .ZN(n13447) );
  INV_X1 U15617 ( .A(n13442), .ZN(n13445) );
  NAND2_X1 U15618 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n15268)
         );
  OAI21_X1 U15619 ( .B1(n13443), .B2(n13476), .A(n15268), .ZN(n13444) );
  AOI21_X1 U15620 ( .B1(n13445), .B2(n13467), .A(n13444), .ZN(n13446) );
  OAI211_X1 U15621 ( .C1(n14859), .C2(n13461), .A(n13447), .B(n13446), .ZN(
        P2_U3200) );
  INV_X1 U15622 ( .A(n13448), .ZN(n13452) );
  INV_X1 U15623 ( .A(n13449), .ZN(n13451) );
  NOR3_X1 U15624 ( .A1(n13452), .A2(n13451), .A3(n13450), .ZN(n13456) );
  INV_X1 U15625 ( .A(n13453), .ZN(n13455) );
  OAI21_X1 U15626 ( .B1(n13456), .B2(n13455), .A(n13454), .ZN(n13460) );
  AOI22_X1 U15627 ( .A1(n13474), .A2(n13510), .B1(n13475), .B2(n13512), .ZN(
        n13638) );
  OAI22_X1 U15628 ( .A1(n13476), .A2(n13638), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13457), .ZN(n13458) );
  AOI21_X1 U15629 ( .B1(n13642), .B2(n13467), .A(n13458), .ZN(n13459) );
  OAI211_X1 U15630 ( .C1(n13644), .C2(n13461), .A(n13460), .B(n13459), .ZN(
        P2_U3201) );
  NAND2_X1 U15631 ( .A1(n7492), .A2(n13463), .ZN(n13464) );
  XNOR2_X1 U15632 ( .A(n13465), .B(n13464), .ZN(n13471) );
  AOI22_X1 U15633 ( .A1(n13514), .A2(n13474), .B1(n13475), .B2(n13516), .ZN(
        n13701) );
  INV_X1 U15634 ( .A(n13466), .ZN(n13705) );
  AOI22_X1 U15635 ( .A1(n13467), .A2(n13705), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13468) );
  OAI21_X1 U15636 ( .B1(n13701), .B2(n13476), .A(n13468), .ZN(n13469) );
  AOI21_X1 U15637 ( .B1(n13813), .B2(n13501), .A(n13469), .ZN(n13470) );
  OAI21_X1 U15638 ( .B1(n13471), .B2(n13503), .A(n13470), .ZN(P2_U3205) );
  XNOR2_X1 U15639 ( .A(n13473), .B(n13472), .ZN(n13481) );
  AOI22_X1 U15640 ( .A1(n13514), .A2(n13475), .B1(n13474), .B2(n13512), .ZN(
        n13665) );
  NOR2_X1 U15641 ( .A1(n13665), .A2(n13476), .ZN(n13479) );
  OAI22_X1 U15642 ( .A1(n13669), .A2(n13498), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13477), .ZN(n13478) );
  AOI211_X1 U15643 ( .C1(n13800), .C2(n13501), .A(n13479), .B(n13478), .ZN(
        n13480) );
  OAI21_X1 U15644 ( .B1(n13481), .B2(n13503), .A(n13480), .ZN(P2_U3207) );
  XNOR2_X1 U15645 ( .A(n13483), .B(n13482), .ZN(n13489) );
  OAI22_X1 U15646 ( .A1(n13485), .A2(n13492), .B1(n13484), .B2(n13495), .ZN(
        n13725) );
  AOI22_X1 U15647 ( .A1(n13725), .A2(n13496), .B1(P2_REG3_REG_18__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13486) );
  OAI21_X1 U15648 ( .B1(n13730), .B2(n13498), .A(n13486), .ZN(n13487) );
  AOI21_X1 U15649 ( .B1(n13822), .B2(n13501), .A(n13487), .ZN(n13488) );
  OAI21_X1 U15650 ( .B1(n13489), .B2(n13503), .A(n13488), .ZN(P2_U3210) );
  INV_X1 U15651 ( .A(n13614), .ZN(n13499) );
  OAI22_X1 U15652 ( .A1(n13495), .A2(n13494), .B1(n13493), .B2(n13492), .ZN(
        n13608) );
  AOI22_X1 U15653 ( .A1(n13496), .A2(n13608), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13497) );
  OAI21_X1 U15654 ( .B1(n13499), .B2(n13498), .A(n13497), .ZN(n13500) );
  AOI21_X1 U15655 ( .B1(n13779), .B2(n13501), .A(n13500), .ZN(n13502) );
  OAI21_X1 U15656 ( .B1(n13504), .B2(n13503), .A(n13502), .ZN(P2_U3212) );
  INV_X2 U15657 ( .A(P2_U3947), .ZN(n13534) );
  MUX2_X1 U15658 ( .A(n13564), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13534), .Z(
        P2_U3562) );
  MUX2_X1 U15659 ( .A(n13505), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13534), .Z(
        P2_U3561) );
  MUX2_X1 U15660 ( .A(n13506), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13534), .Z(
        P2_U3560) );
  MUX2_X1 U15661 ( .A(n13507), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13534), .Z(
        P2_U3559) );
  MUX2_X1 U15662 ( .A(n13508), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13534), .Z(
        P2_U3558) );
  MUX2_X1 U15663 ( .A(n13509), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13534), .Z(
        P2_U3557) );
  MUX2_X1 U15664 ( .A(n13510), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13534), .Z(
        P2_U3556) );
  MUX2_X1 U15665 ( .A(n13511), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13534), .Z(
        P2_U3555) );
  MUX2_X1 U15666 ( .A(n13512), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13534), .Z(
        P2_U3554) );
  MUX2_X1 U15667 ( .A(n13513), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13534), .Z(
        P2_U3553) );
  MUX2_X1 U15668 ( .A(n13514), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13534), .Z(
        P2_U3552) );
  MUX2_X1 U15669 ( .A(n13515), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13534), .Z(
        P2_U3551) );
  MUX2_X1 U15670 ( .A(n13516), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13534), .Z(
        P2_U3550) );
  MUX2_X1 U15671 ( .A(n13517), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13534), .Z(
        P2_U3549) );
  MUX2_X1 U15672 ( .A(n13518), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13534), .Z(
        P2_U3548) );
  MUX2_X1 U15673 ( .A(n13519), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13534), .Z(
        P2_U3547) );
  MUX2_X1 U15674 ( .A(n13520), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13534), .Z(
        P2_U3546) );
  MUX2_X1 U15675 ( .A(n13521), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13534), .Z(
        P2_U3545) );
  MUX2_X1 U15676 ( .A(n13522), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13534), .Z(
        P2_U3543) );
  MUX2_X1 U15677 ( .A(n13523), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13534), .Z(
        P2_U3542) );
  MUX2_X1 U15678 ( .A(n13524), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13534), .Z(
        P2_U3541) );
  MUX2_X1 U15679 ( .A(n13525), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13534), .Z(
        P2_U3540) );
  MUX2_X1 U15680 ( .A(n13526), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13534), .Z(
        P2_U3539) );
  MUX2_X1 U15681 ( .A(n13527), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13534), .Z(
        P2_U3538) );
  MUX2_X1 U15682 ( .A(n13528), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13534), .Z(
        P2_U3537) );
  MUX2_X1 U15683 ( .A(n13529), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13534), .Z(
        P2_U3536) );
  MUX2_X1 U15684 ( .A(n13530), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13534), .Z(
        P2_U3535) );
  MUX2_X1 U15685 ( .A(n13531), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13534), .Z(
        P2_U3534) );
  MUX2_X1 U15686 ( .A(n13532), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13534), .Z(
        P2_U3533) );
  MUX2_X1 U15687 ( .A(n13533), .B(n6866), .S(n13534), .Z(P2_U3532) );
  MUX2_X1 U15688 ( .A(n8463), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13534), .Z(
        P2_U3531) );
  XOR2_X1 U15689 ( .A(n13536), .B(n13535), .Z(n13537) );
  AOI22_X1 U15690 ( .A1(n6858), .A2(n15254), .B1(n15264), .B2(n13537), .ZN(
        n13546) );
  MUX2_X1 U15691 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n9413), .S(n13538), .Z(
        n13539) );
  NAND3_X1 U15692 ( .A1(n15206), .A2(n13540), .A3(n13539), .ZN(n13541) );
  NAND3_X1 U15693 ( .A1(n15271), .A2(n13542), .A3(n13541), .ZN(n13545) );
  NAND2_X1 U15694 ( .A1(n15270), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n13544) );
  NAND2_X1 U15695 ( .A1(P2_U3088), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n13543) );
  NAND4_X1 U15696 ( .A1(n13546), .A2(n13545), .A3(n13544), .A4(n13543), .ZN(
        P2_U3216) );
  OAI22_X1 U15697 ( .A1(n15250), .A2(n8366), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13547), .ZN(n13548) );
  AOI21_X1 U15698 ( .B1(n13554), .B2(n15254), .A(n13548), .ZN(n13562) );
  MUX2_X1 U15699 ( .A(n9523), .B(P2_REG1_REG_7__SCAN_IN), .S(n13554), .Z(
        n13549) );
  NAND3_X1 U15700 ( .A1(n13551), .A2(n13550), .A3(n13549), .ZN(n13552) );
  NAND3_X1 U15701 ( .A1(n15264), .A2(n13553), .A3(n13552), .ZN(n13561) );
  MUX2_X1 U15702 ( .A(n10297), .B(P2_REG2_REG_7__SCAN_IN), .S(n13554), .Z(
        n13555) );
  NAND3_X1 U15703 ( .A1(n13557), .A2(n13556), .A3(n13555), .ZN(n13558) );
  NAND3_X1 U15704 ( .A1(n15271), .A2(n13559), .A3(n13558), .ZN(n13560) );
  NAND3_X1 U15705 ( .A1(n13562), .A2(n13561), .A3(n13560), .ZN(P2_U3221) );
  XNOR2_X1 U15706 ( .A(n13571), .B(n13566), .ZN(n13563) );
  NAND2_X1 U15707 ( .A1(n13563), .A2(n14852), .ZN(n13756) );
  NAND2_X1 U15708 ( .A1(n13565), .A2(n13564), .ZN(n13758) );
  NOR2_X1 U15709 ( .A1(n15292), .A2(n13758), .ZN(n13575) );
  INV_X1 U15710 ( .A(n13566), .ZN(n13757) );
  NOR2_X1 U15711 ( .A1(n13757), .A2(n15282), .ZN(n13567) );
  AOI211_X1 U15712 ( .C1(n15292), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13575), 
        .B(n13567), .ZN(n13568) );
  OAI21_X1 U15713 ( .B1(n13756), .B2(n13685), .A(n13568), .ZN(P2_U3234) );
  INV_X1 U15714 ( .A(n13570), .ZN(n13573) );
  INV_X1 U15715 ( .A(n13571), .ZN(n13572) );
  OAI211_X1 U15716 ( .C1(n13760), .C2(n13573), .A(n13572), .B(n14852), .ZN(
        n13759) );
  NOR2_X1 U15717 ( .A1(n13760), .A2(n15282), .ZN(n13574) );
  AOI211_X1 U15718 ( .C1(n15292), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13575), 
        .B(n13574), .ZN(n13576) );
  OAI21_X1 U15719 ( .B1(n13685), .B2(n13759), .A(n13576), .ZN(P2_U3235) );
  OAI21_X1 U15720 ( .B1(n13578), .B2(n13579), .A(n13577), .ZN(n13770) );
  AOI21_X1 U15721 ( .B1(n13580), .B2(n13579), .A(n14819), .ZN(n13583) );
  AOI21_X1 U15722 ( .B1(n13583), .B2(n13582), .A(n13581), .ZN(n13769) );
  AOI21_X1 U15723 ( .B1(n13767), .B2(n13596), .A(n13728), .ZN(n13585) );
  AND2_X1 U15724 ( .A1(n13585), .A2(n13584), .ZN(n13766) );
  AOI22_X1 U15725 ( .A1(n13766), .A2(n13587), .B1(n15279), .B2(n13586), .ZN(
        n13588) );
  AOI21_X1 U15726 ( .B1(n13769), .B2(n13588), .A(n15292), .ZN(n13589) );
  INV_X1 U15727 ( .A(n13589), .ZN(n13591) );
  AOI22_X1 U15728 ( .A1(n13767), .A2(n14844), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n15292), .ZN(n13590) );
  OAI211_X1 U15729 ( .C1(n13738), .C2(n13770), .A(n13591), .B(n13590), .ZN(
        P2_U3237) );
  XNOR2_X1 U15730 ( .A(n13593), .B(n13592), .ZN(n13595) );
  AOI21_X1 U15731 ( .B1(n13595), .B2(n14841), .A(n13594), .ZN(n13777) );
  AOI21_X1 U15732 ( .B1(n13773), .B2(n13612), .A(n13728), .ZN(n13597) );
  NAND2_X1 U15733 ( .A1(n13597), .A2(n13596), .ZN(n13776) );
  AOI22_X1 U15734 ( .A1(n15292), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n13598), 
        .B2(n15279), .ZN(n13600) );
  NAND2_X1 U15735 ( .A1(n13773), .A2(n14844), .ZN(n13599) );
  OAI211_X1 U15736 ( .C1(n13776), .C2(n13685), .A(n13600), .B(n13599), .ZN(
        n13601) );
  INV_X1 U15737 ( .A(n13601), .ZN(n13605) );
  OR2_X1 U15738 ( .A1(n13603), .A2(n13602), .ZN(n13772) );
  NAND3_X1 U15739 ( .A1(n13772), .A2(n13771), .A3(n15288), .ZN(n13604) );
  OAI211_X1 U15740 ( .C1(n13777), .C2(n15292), .A(n13605), .B(n13604), .ZN(
        P2_U3238) );
  XNOR2_X1 U15741 ( .A(n13607), .B(n13606), .ZN(n13609) );
  AOI21_X1 U15742 ( .B1(n13609), .B2(n14841), .A(n13608), .ZN(n13781) );
  XNOR2_X1 U15743 ( .A(n13611), .B(n13610), .ZN(n13782) );
  INV_X1 U15744 ( .A(n13782), .ZN(n13619) );
  AOI21_X1 U15745 ( .B1(n13628), .B2(n13779), .A(n13728), .ZN(n13613) );
  AND2_X1 U15746 ( .A1(n13613), .A2(n13612), .ZN(n13778) );
  NAND2_X1 U15747 ( .A1(n13778), .A2(n15285), .ZN(n13616) );
  AOI22_X1 U15748 ( .A1(n15292), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n13614), 
        .B2(n15279), .ZN(n13615) );
  OAI211_X1 U15749 ( .C1(n13617), .C2(n15282), .A(n13616), .B(n13615), .ZN(
        n13618) );
  AOI21_X1 U15750 ( .B1(n13619), .B2(n15288), .A(n13618), .ZN(n13620) );
  OAI21_X1 U15751 ( .B1(n13781), .B2(n15292), .A(n13620), .ZN(P2_U3239) );
  XNOR2_X1 U15752 ( .A(n13622), .B(n13621), .ZN(n13624) );
  AOI21_X1 U15753 ( .B1(n13624), .B2(n14841), .A(n13623), .ZN(n13787) );
  OAI21_X1 U15754 ( .B1(n13627), .B2(n13626), .A(n13625), .ZN(n13783) );
  INV_X1 U15755 ( .A(n13641), .ZN(n13630) );
  INV_X1 U15756 ( .A(n13628), .ZN(n13629) );
  AOI211_X1 U15757 ( .C1(n13785), .C2(n13630), .A(n13728), .B(n13629), .ZN(
        n13784) );
  NAND2_X1 U15758 ( .A1(n13784), .A2(n15285), .ZN(n13633) );
  AOI22_X1 U15759 ( .A1(n15292), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n13631), 
        .B2(n15279), .ZN(n13632) );
  OAI211_X1 U15760 ( .C1(n13634), .C2(n15282), .A(n13633), .B(n13632), .ZN(
        n13635) );
  AOI21_X1 U15761 ( .B1(n13783), .B2(n15288), .A(n13635), .ZN(n13636) );
  OAI21_X1 U15762 ( .B1(n13787), .B2(n15292), .A(n13636), .ZN(P2_U3240) );
  XNOR2_X1 U15763 ( .A(n13637), .B(n13645), .ZN(n13640) );
  INV_X1 U15764 ( .A(n13638), .ZN(n13639) );
  AOI21_X1 U15765 ( .B1(n13640), .B2(n14841), .A(n13639), .ZN(n13792) );
  AOI211_X1 U15766 ( .C1(n13790), .C2(n13656), .A(n13728), .B(n13641), .ZN(
        n13789) );
  AOI22_X1 U15767 ( .A1(n15292), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n13642), 
        .B2(n15279), .ZN(n13643) );
  OAI21_X1 U15768 ( .B1(n13644), .B2(n15282), .A(n13643), .ZN(n13648) );
  XNOR2_X1 U15769 ( .A(n13646), .B(n13645), .ZN(n13793) );
  NOR2_X1 U15770 ( .A1(n13793), .A2(n13738), .ZN(n13647) );
  AOI211_X1 U15771 ( .C1(n13789), .C2(n15285), .A(n13648), .B(n13647), .ZN(
        n13649) );
  OAI21_X1 U15772 ( .B1(n15292), .B2(n13792), .A(n13649), .ZN(P2_U3241) );
  XNOR2_X1 U15773 ( .A(n6684), .B(n13651), .ZN(n13798) );
  XOR2_X1 U15774 ( .A(n13651), .B(n13650), .Z(n13653) );
  AOI21_X1 U15775 ( .B1(n13653), .B2(n14841), .A(n13652), .ZN(n13797) );
  OAI21_X1 U15776 ( .B1(n13654), .B2(n14827), .A(n13797), .ZN(n13655) );
  NAND2_X1 U15777 ( .A1(n13655), .A2(n13748), .ZN(n13661) );
  INV_X1 U15778 ( .A(n13656), .ZN(n13657) );
  AOI211_X1 U15779 ( .C1(n13795), .C2(n13667), .A(n13728), .B(n13657), .ZN(
        n13794) );
  INV_X1 U15780 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n13658) );
  OAI22_X1 U15781 ( .A1(n7316), .A2(n15282), .B1(n13748), .B2(n13658), .ZN(
        n13659) );
  AOI21_X1 U15782 ( .B1(n13794), .B2(n15285), .A(n13659), .ZN(n13660) );
  OAI211_X1 U15783 ( .C1(n13738), .C2(n13798), .A(n13661), .B(n13660), .ZN(
        P2_U3242) );
  OAI211_X1 U15784 ( .C1(n13664), .C2(n13663), .A(n13662), .B(n14841), .ZN(
        n13666) );
  INV_X1 U15785 ( .A(n13667), .ZN(n13668) );
  AOI211_X1 U15786 ( .C1(n13800), .C2(n13681), .A(n13728), .B(n13668), .ZN(
        n13799) );
  INV_X1 U15787 ( .A(n13669), .ZN(n13670) );
  AOI22_X1 U15788 ( .A1(n13670), .A2(n15279), .B1(P2_REG2_REG_22__SCAN_IN), 
        .B2(n15292), .ZN(n13671) );
  OAI21_X1 U15789 ( .B1(n7269), .B2(n15282), .A(n13671), .ZN(n13677) );
  NOR2_X1 U15790 ( .A1(n13673), .A2(n13672), .ZN(n13674) );
  OR2_X1 U15791 ( .A1(n13675), .A2(n13674), .ZN(n13803) );
  NOR2_X1 U15792 ( .A1(n13803), .A2(n13738), .ZN(n13676) );
  AOI211_X1 U15793 ( .C1(n13799), .C2(n15285), .A(n13677), .B(n13676), .ZN(
        n13678) );
  OAI21_X1 U15794 ( .B1(n15292), .B2(n13802), .A(n13678), .ZN(P2_U3243) );
  XNOR2_X1 U15795 ( .A(n6911), .B(n6850), .ZN(n13807) );
  NAND2_X1 U15796 ( .A1(n13804), .A2(n13703), .ZN(n13680) );
  NAND3_X1 U15797 ( .A1(n13681), .A2(n14852), .A3(n13680), .ZN(n13806) );
  AOI22_X1 U15798 ( .A1(n13682), .A2(n15279), .B1(n15292), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n13684) );
  NAND2_X1 U15799 ( .A1(n13804), .A2(n14844), .ZN(n13683) );
  OAI211_X1 U15800 ( .C1(n13806), .C2(n13685), .A(n13684), .B(n13683), .ZN(
        n13694) );
  NOR2_X1 U15801 ( .A1(n13687), .A2(n13686), .ZN(n13688) );
  OR2_X1 U15802 ( .A1(n13689), .A2(n13688), .ZN(n13692) );
  INV_X1 U15803 ( .A(n13690), .ZN(n13691) );
  AOI21_X1 U15804 ( .B1(n13692), .B2(n14841), .A(n13691), .ZN(n13810) );
  NOR2_X1 U15805 ( .A1(n13810), .A2(n15292), .ZN(n13693) );
  AOI211_X1 U15806 ( .C1(n13807), .C2(n15288), .A(n13694), .B(n13693), .ZN(
        n13695) );
  INV_X1 U15807 ( .A(n13695), .ZN(P2_U3244) );
  XOR2_X1 U15808 ( .A(n13696), .B(n13700), .Z(n13815) );
  INV_X1 U15809 ( .A(n13697), .ZN(n13698) );
  AOI21_X1 U15810 ( .B1(n13700), .B2(n13699), .A(n13698), .ZN(n13702) );
  OAI21_X1 U15811 ( .B1(n13702), .B2(n14819), .A(n13701), .ZN(n13811) );
  INV_X1 U15812 ( .A(n13813), .ZN(n13708) );
  AOI21_X1 U15813 ( .B1(n13813), .B2(n13717), .A(n13728), .ZN(n13704) );
  AND2_X1 U15814 ( .A1(n13704), .A2(n13703), .ZN(n13812) );
  NAND2_X1 U15815 ( .A1(n13812), .A2(n15285), .ZN(n13707) );
  AOI22_X1 U15816 ( .A1(n15292), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13705), 
        .B2(n15279), .ZN(n13706) );
  OAI211_X1 U15817 ( .C1(n13708), .C2(n15282), .A(n13707), .B(n13706), .ZN(
        n13709) );
  AOI21_X1 U15818 ( .B1(n13811), .B2(n13748), .A(n13709), .ZN(n13710) );
  OAI21_X1 U15819 ( .B1(n13738), .B2(n13815), .A(n13710), .ZN(P2_U3245) );
  XNOR2_X1 U15820 ( .A(n13711), .B(n13713), .ZN(n13820) );
  XOR2_X1 U15821 ( .A(n13713), .B(n13712), .Z(n13715) );
  OAI21_X1 U15822 ( .B1(n13715), .B2(n14819), .A(n13714), .ZN(n13816) );
  OR2_X1 U15823 ( .A1(n13721), .A2(n13727), .ZN(n13716) );
  AND3_X1 U15824 ( .A1(n13717), .A2(n13716), .A3(n14852), .ZN(n13817) );
  NAND2_X1 U15825 ( .A1(n13817), .A2(n15285), .ZN(n13720) );
  AOI22_X1 U15826 ( .A1(n15292), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13718), 
        .B2(n15279), .ZN(n13719) );
  OAI211_X1 U15827 ( .C1(n13721), .C2(n15282), .A(n13720), .B(n13719), .ZN(
        n13722) );
  AOI21_X1 U15828 ( .B1(n13816), .B2(n13748), .A(n13722), .ZN(n13723) );
  OAI21_X1 U15829 ( .B1(n13738), .B2(n13820), .A(n13723), .ZN(P2_U3246) );
  XOR2_X1 U15830 ( .A(n13737), .B(n13724), .Z(n13726) );
  AOI21_X1 U15831 ( .B1(n13726), .B2(n14841), .A(n13725), .ZN(n13824) );
  AOI211_X1 U15832 ( .C1(n13822), .C2(n13729), .A(n13728), .B(n13727), .ZN(
        n13821) );
  INV_X1 U15833 ( .A(n13822), .ZN(n13733) );
  INV_X1 U15834 ( .A(n13730), .ZN(n13731) );
  AOI22_X1 U15835 ( .A1(n15292), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13731), 
        .B2(n15279), .ZN(n13732) );
  OAI21_X1 U15836 ( .B1(n13733), .B2(n15282), .A(n13732), .ZN(n13740) );
  INV_X1 U15837 ( .A(n13734), .ZN(n13735) );
  AOI21_X1 U15838 ( .B1(n13737), .B2(n13736), .A(n13735), .ZN(n13825) );
  NOR2_X1 U15839 ( .A1(n13825), .A2(n13738), .ZN(n13739) );
  AOI211_X1 U15840 ( .C1(n13821), .C2(n15285), .A(n13740), .B(n13739), .ZN(
        n13741) );
  OAI21_X1 U15841 ( .B1(n15292), .B2(n13824), .A(n13741), .ZN(P2_U3247) );
  OAI211_X1 U15842 ( .C1(n13743), .C2(n13751), .A(n13742), .B(n14841), .ZN(
        n13745) );
  NAND2_X1 U15843 ( .A1(n13745), .A2(n13744), .ZN(n14869) );
  OAI211_X1 U15844 ( .C1(n14817), .C2(n14868), .A(n14852), .B(n13746), .ZN(
        n14866) );
  OAI22_X1 U15845 ( .A1(n14866), .A2(n6843), .B1(n14827), .B2(n13747), .ZN(
        n13749) );
  OAI21_X1 U15846 ( .B1(n14869), .B2(n13749), .A(n13748), .ZN(n13755) );
  AOI22_X1 U15847 ( .A1(n13750), .A2(n14844), .B1(P2_REG2_REG_16__SCAN_IN), 
        .B2(n15292), .ZN(n13754) );
  NAND2_X1 U15848 ( .A1(n13752), .A2(n13751), .ZN(n14864) );
  NAND3_X1 U15849 ( .A1(n14865), .A2(n14864), .A3(n15288), .ZN(n13753) );
  NAND3_X1 U15850 ( .A1(n13755), .A2(n13754), .A3(n13753), .ZN(P2_U3249) );
  OAI211_X1 U15851 ( .C1(n13757), .C2(n15380), .A(n13756), .B(n13758), .ZN(
        n13826) );
  MUX2_X1 U15852 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13826), .S(n15401), .Z(
        P2_U3530) );
  OAI211_X1 U15853 ( .C1(n13760), .C2(n15380), .A(n13759), .B(n13758), .ZN(
        n13827) );
  MUX2_X1 U15854 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13827), .S(n15401), .Z(
        P2_U3529) );
  AOI21_X1 U15855 ( .B1(n15368), .B2(n13762), .A(n13761), .ZN(n13763) );
  OAI211_X1 U15856 ( .C1(n15350), .C2(n13765), .A(n13764), .B(n13763), .ZN(
        n13828) );
  MUX2_X1 U15857 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13828), .S(n15401), .Z(
        P2_U3528) );
  AOI21_X1 U15858 ( .B1(n15368), .B2(n13767), .A(n13766), .ZN(n13768) );
  MUX2_X1 U15859 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13829), .S(n15401), .Z(
        P2_U3527) );
  NAND3_X1 U15860 ( .A1(n13772), .A2(n13771), .A3(n15377), .ZN(n13775) );
  NAND2_X1 U15861 ( .A1(n13773), .A2(n15368), .ZN(n13774) );
  NAND4_X1 U15862 ( .A1(n13777), .A2(n13776), .A3(n13775), .A4(n13774), .ZN(
        n13830) );
  MUX2_X1 U15863 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13830), .S(n15401), .Z(
        P2_U3526) );
  AOI21_X1 U15864 ( .B1(n15368), .B2(n13779), .A(n13778), .ZN(n13780) );
  OAI211_X1 U15865 ( .C1(n15350), .C2(n13782), .A(n13781), .B(n13780), .ZN(
        n13831) );
  MUX2_X1 U15866 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13831), .S(n15401), .Z(
        P2_U3525) );
  INV_X1 U15867 ( .A(n13783), .ZN(n13788) );
  AOI21_X1 U15868 ( .B1(n15368), .B2(n13785), .A(n13784), .ZN(n13786) );
  OAI211_X1 U15869 ( .C1(n15350), .C2(n13788), .A(n13787), .B(n13786), .ZN(
        n13832) );
  MUX2_X1 U15870 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13832), .S(n15401), .Z(
        P2_U3524) );
  AOI21_X1 U15871 ( .B1(n15368), .B2(n13790), .A(n13789), .ZN(n13791) );
  OAI211_X1 U15872 ( .C1(n15350), .C2(n13793), .A(n13792), .B(n13791), .ZN(
        n13833) );
  MUX2_X1 U15873 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13833), .S(n15401), .Z(
        P2_U3523) );
  AOI21_X1 U15874 ( .B1(n15368), .B2(n13795), .A(n13794), .ZN(n13796) );
  OAI211_X1 U15875 ( .C1(n15350), .C2(n13798), .A(n13797), .B(n13796), .ZN(
        n13834) );
  MUX2_X1 U15876 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13834), .S(n15401), .Z(
        P2_U3522) );
  AOI21_X1 U15877 ( .B1(n15368), .B2(n13800), .A(n13799), .ZN(n13801) );
  OAI211_X1 U15878 ( .C1(n15350), .C2(n13803), .A(n13802), .B(n13801), .ZN(
        n13835) );
  MUX2_X1 U15879 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13835), .S(n15401), .Z(
        P2_U3521) );
  NAND2_X1 U15880 ( .A1(n13804), .A2(n15368), .ZN(n13805) );
  AND2_X1 U15881 ( .A1(n13806), .A2(n13805), .ZN(n13809) );
  NAND2_X1 U15882 ( .A1(n13807), .A2(n15377), .ZN(n13808) );
  NAND3_X1 U15883 ( .A1(n13810), .A2(n13809), .A3(n13808), .ZN(n13836) );
  MUX2_X1 U15884 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13836), .S(n15401), .Z(
        P2_U3520) );
  AOI211_X1 U15885 ( .C1(n15368), .C2(n13813), .A(n13812), .B(n13811), .ZN(
        n13814) );
  OAI21_X1 U15886 ( .B1(n15350), .B2(n13815), .A(n13814), .ZN(n13837) );
  MUX2_X1 U15887 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13837), .S(n15401), .Z(
        P2_U3519) );
  AOI211_X1 U15888 ( .C1(n15368), .C2(n13818), .A(n13817), .B(n13816), .ZN(
        n13819) );
  OAI21_X1 U15889 ( .B1(n15350), .B2(n13820), .A(n13819), .ZN(n13838) );
  MUX2_X1 U15890 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13838), .S(n15401), .Z(
        P2_U3518) );
  AOI21_X1 U15891 ( .B1(n15368), .B2(n13822), .A(n13821), .ZN(n13823) );
  OAI211_X1 U15892 ( .C1(n13825), .C2(n15350), .A(n13824), .B(n13823), .ZN(
        n13839) );
  MUX2_X1 U15893 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13839), .S(n15401), .Z(
        P2_U3517) );
  MUX2_X1 U15894 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13826), .S(n15387), .Z(
        P2_U3498) );
  MUX2_X1 U15895 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13827), .S(n15387), .Z(
        P2_U3497) );
  MUX2_X1 U15896 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n13828), .S(n15387), .Z(
        P2_U3496) );
  MUX2_X1 U15897 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13829), .S(n15387), .Z(
        P2_U3495) );
  MUX2_X1 U15898 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13830), .S(n15387), .Z(
        P2_U3494) );
  MUX2_X1 U15899 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13831), .S(n15387), .Z(
        P2_U3493) );
  MUX2_X1 U15900 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13832), .S(n15387), .Z(
        P2_U3492) );
  MUX2_X1 U15901 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13833), .S(n15387), .Z(
        P2_U3491) );
  MUX2_X1 U15902 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13834), .S(n15387), .Z(
        P2_U3490) );
  MUX2_X1 U15903 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13835), .S(n15387), .Z(
        P2_U3489) );
  MUX2_X1 U15904 ( .A(n13836), .B(P2_REG0_REG_21__SCAN_IN), .S(n15385), .Z(
        P2_U3488) );
  MUX2_X1 U15905 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13837), .S(n15387), .Z(
        P2_U3487) );
  MUX2_X1 U15906 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13838), .S(n15387), .Z(
        P2_U3486) );
  MUX2_X1 U15907 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13839), .S(n15387), .Z(
        P2_U3484) );
  INV_X1 U15908 ( .A(n14692), .ZN(n13843) );
  INV_X1 U15909 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n13840) );
  NOR4_X1 U15910 ( .A1(n7641), .A2(P2_IR_REG_30__SCAN_IN), .A3(n13840), .A4(
        P2_U3088), .ZN(n13841) );
  AOI21_X1 U15911 ( .B1(n13848), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n13841), 
        .ZN(n13842) );
  OAI21_X1 U15912 ( .B1(n13843), .B2(n13854), .A(n13842), .ZN(P2_U3296) );
  OAI222_X1 U15913 ( .A1(n13852), .A2(n13846), .B1(n13854), .B2(n13845), .C1(
        n13844), .C2(P2_U3088), .ZN(P2_U3298) );
  AOI21_X1 U15914 ( .B1(n13848), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13847), 
        .ZN(n13849) );
  OAI21_X1 U15915 ( .B1(n13850), .B2(n13854), .A(n13849), .ZN(P2_U3299) );
  INV_X1 U15916 ( .A(n13851), .ZN(n14697) );
  OAI222_X1 U15917 ( .A1(n13855), .A2(P2_U3088), .B1(n13854), .B2(n14697), 
        .C1(n13853), .C2(n13852), .ZN(P2_U3301) );
  INV_X1 U15918 ( .A(n13856), .ZN(n13857) );
  MUX2_X1 U15919 ( .A(n13857), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  XOR2_X1 U15920 ( .A(n13859), .B(n13858), .Z(n13866) );
  INV_X1 U15921 ( .A(n14392), .ZN(n13863) );
  NAND2_X1 U15922 ( .A1(n14424), .A2(n14571), .ZN(n13861) );
  NAND2_X1 U15923 ( .A1(n14262), .A2(n14573), .ZN(n13860) );
  NAND2_X1 U15924 ( .A1(n13861), .A2(n13860), .ZN(n14607) );
  AOI22_X1 U15925 ( .A1(n13987), .A2(n14607), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13862) );
  OAI21_X1 U15926 ( .B1(n14941), .B2(n13863), .A(n13862), .ZN(n13864) );
  AOI21_X1 U15927 ( .B1(n14608), .B2(n14937), .A(n13864), .ZN(n13865) );
  OAI21_X1 U15928 ( .B1(n13866), .B2(n14932), .A(n13865), .ZN(P1_U3214) );
  NAND2_X1 U15929 ( .A1(n13950), .A2(n13867), .ZN(n13868) );
  XOR2_X1 U15930 ( .A(n13869), .B(n13868), .Z(n13876) );
  NAND2_X1 U15931 ( .A1(n14497), .A2(n14571), .ZN(n13871) );
  NAND2_X1 U15932 ( .A1(n14423), .A2(n14573), .ZN(n13870) );
  AND2_X1 U15933 ( .A1(n13871), .A2(n13870), .ZN(n14630) );
  OAI22_X1 U15934 ( .A1(n13918), .A2(n14630), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13872), .ZN(n13874) );
  NOR2_X1 U15935 ( .A1(n14461), .A2(n14005), .ZN(n13873) );
  AOI211_X1 U15936 ( .C1(n14459), .C2(n14001), .A(n13874), .B(n13873), .ZN(
        n13875) );
  OAI21_X1 U15937 ( .B1(n13876), .B2(n14932), .A(n13875), .ZN(P1_U3216) );
  AOI21_X1 U15938 ( .B1(n13878), .B2(n13877), .A(n14932), .ZN(n13879) );
  NAND2_X1 U15939 ( .A1(n13879), .A2(n13887), .ZN(n13885) );
  NOR2_X1 U15940 ( .A1(n13880), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14355) );
  AOI21_X1 U15941 ( .B1(n13997), .B2(n14498), .A(n14355), .ZN(n13881) );
  OAI21_X1 U15942 ( .B1(n14530), .B2(n14925), .A(n13881), .ZN(n13882) );
  AOI21_X1 U15943 ( .B1(n13883), .B2(n14001), .A(n13882), .ZN(n13884) );
  OAI211_X1 U15944 ( .C1(n14534), .C2(n14005), .A(n13885), .B(n13884), .ZN(
        P1_U3219) );
  NAND2_X1 U15945 ( .A1(n13887), .A2(n13886), .ZN(n13947) );
  NAND2_X1 U15946 ( .A1(n13947), .A2(n13932), .ZN(n13931) );
  NAND2_X1 U15947 ( .A1(n13931), .A2(n13888), .ZN(n13890) );
  NOR2_X1 U15948 ( .A1(n13890), .A2(n13891), .ZN(n13889) );
  AOI21_X1 U15949 ( .B1(n13891), .B2(n13890), .A(n13889), .ZN(n13896) );
  NAND2_X1 U15950 ( .A1(n14001), .A2(n14491), .ZN(n13893) );
  AOI22_X1 U15951 ( .A1(n13997), .A2(n14497), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13892) );
  OAI211_X1 U15952 ( .C1(n14532), .C2(n14925), .A(n13893), .B(n13892), .ZN(
        n13894) );
  AOI21_X1 U15953 ( .B1(n14644), .B2(n14937), .A(n13894), .ZN(n13895) );
  OAI21_X1 U15954 ( .B1(n13896), .B2(n14932), .A(n13895), .ZN(P1_U3223) );
  AOI211_X1 U15955 ( .C1(n13898), .C2(n13897), .A(n14932), .B(n6769), .ZN(
        n13899) );
  INV_X1 U15956 ( .A(n13899), .ZN(n13905) );
  NAND2_X1 U15957 ( .A1(n14270), .A2(n14571), .ZN(n13901) );
  NAND2_X1 U15958 ( .A1(n14268), .A2(n14573), .ZN(n13900) );
  AND2_X1 U15959 ( .A1(n13901), .A2(n13900), .ZN(n14733) );
  OAI21_X1 U15960 ( .B1(n13918), .B2(n14733), .A(n13902), .ZN(n13903) );
  AOI21_X1 U15961 ( .B1(n14001), .B2(n14736), .A(n13903), .ZN(n13904) );
  OAI211_X1 U15962 ( .C1(n14746), .C2(n14005), .A(n13905), .B(n13904), .ZN(
        P1_U3224) );
  XOR2_X1 U15963 ( .A(n13907), .B(n13906), .Z(n13913) );
  NAND2_X1 U15964 ( .A1(n14001), .A2(n14427), .ZN(n13909) );
  AOI22_X1 U15965 ( .A1(n13964), .A2(n14423), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13908) );
  OAI211_X1 U15966 ( .C1(n13910), .C2(n14926), .A(n13909), .B(n13908), .ZN(
        n13911) );
  AOI21_X1 U15967 ( .B1(n14431), .B2(n14937), .A(n13911), .ZN(n13912) );
  OAI21_X1 U15968 ( .B1(n13913), .B2(n14932), .A(n13912), .ZN(P1_U3225) );
  OAI21_X1 U15969 ( .B1(n13916), .B2(n13915), .A(n13914), .ZN(n13917) );
  NAND2_X1 U15970 ( .A1(n13917), .A2(n13994), .ZN(n13921) );
  AOI22_X1 U15971 ( .A1(n14265), .A2(n14573), .B1(n14571), .B2(n14266), .ZN(
        n14559) );
  NAND2_X1 U15972 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n15084)
         );
  OAI21_X1 U15973 ( .B1(n13918), .B2(n14559), .A(n15084), .ZN(n13919) );
  AOI21_X1 U15974 ( .B1(n14001), .B2(n14562), .A(n13919), .ZN(n13920) );
  OAI211_X1 U15975 ( .C1(n14944), .C2(n14005), .A(n13921), .B(n13920), .ZN(
        P1_U3228) );
  XOR2_X1 U15976 ( .A(n13923), .B(n13922), .Z(n13930) );
  NAND2_X1 U15977 ( .A1(n14470), .A2(n14571), .ZN(n13925) );
  NAND2_X1 U15978 ( .A1(n14264), .A2(n14573), .ZN(n13924) );
  NAND2_X1 U15979 ( .A1(n13925), .A2(n13924), .ZN(n14437) );
  AOI22_X1 U15980 ( .A1(n13987), .A2(n14437), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13926) );
  OAI21_X1 U15981 ( .B1(n14941), .B2(n13927), .A(n13926), .ZN(n13928) );
  AOI21_X1 U15982 ( .B1(n14626), .B2(n14937), .A(n13928), .ZN(n13929) );
  OAI21_X1 U15983 ( .B1(n13930), .B2(n14932), .A(n13929), .ZN(P1_U3229) );
  OAI211_X1 U15984 ( .C1(n13947), .C2(n13932), .A(n13931), .B(n13994), .ZN(
        n13936) );
  AOI22_X1 U15985 ( .A1(n13997), .A2(n14506), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13933) );
  OAI21_X1 U15986 ( .B1(n13966), .B2(n14925), .A(n13933), .ZN(n13934) );
  AOI21_X1 U15987 ( .B1(n14509), .B2(n14001), .A(n13934), .ZN(n13935) );
  OAI211_X1 U15988 ( .C1(n14518), .C2(n14005), .A(n13936), .B(n13935), .ZN(
        P1_U3233) );
  NAND2_X1 U15989 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n15024)
         );
  NAND2_X1 U15990 ( .A1(n13987), .A2(n13937), .ZN(n13938) );
  OAI211_X1 U15991 ( .C1(n14941), .C2(n13939), .A(n15024), .B(n13938), .ZN(
        n13944) );
  INV_X1 U15992 ( .A(n13940), .ZN(n14904) );
  AOI211_X1 U15993 ( .C1(n13942), .C2(n13941), .A(n14932), .B(n14904), .ZN(
        n13943) );
  AOI211_X1 U15994 ( .C1(n14112), .C2(n14937), .A(n13944), .B(n13943), .ZN(
        n13945) );
  INV_X1 U15995 ( .A(n13945), .ZN(P1_U3234) );
  NAND2_X1 U15996 ( .A1(n13947), .A2(n13946), .ZN(n13949) );
  AND2_X1 U15997 ( .A1(n13949), .A2(n13948), .ZN(n13951) );
  OAI21_X1 U15998 ( .B1(n13952), .B2(n13951), .A(n13950), .ZN(n13953) );
  NAND2_X1 U15999 ( .A1(n13953), .A2(n13994), .ZN(n13960) );
  NOR2_X1 U16000 ( .A1(n14925), .A2(n13954), .ZN(n13958) );
  OAI22_X1 U16001 ( .A1(n14926), .A2(n13956), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13955), .ZN(n13957) );
  AOI211_X1 U16002 ( .C1(n14473), .C2(n14001), .A(n13958), .B(n13957), .ZN(
        n13959) );
  OAI211_X1 U16003 ( .C1(n14005), .C2(n13961), .A(n13960), .B(n13959), .ZN(
        P1_U3235) );
  XOR2_X1 U16004 ( .A(n13963), .B(n13962), .Z(n13970) );
  NAND2_X1 U16005 ( .A1(n13964), .A2(n14574), .ZN(n13965) );
  NAND2_X1 U16006 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n15102)
         );
  OAI211_X1 U16007 ( .C1(n13966), .C2(n14926), .A(n13965), .B(n15102), .ZN(
        n13967) );
  AOI21_X1 U16008 ( .B1(n14549), .B2(n14001), .A(n13967), .ZN(n13969) );
  NAND2_X1 U16009 ( .A1(n14667), .A2(n14937), .ZN(n13968) );
  OAI211_X1 U16010 ( .C1(n13970), .C2(n14932), .A(n13969), .B(n13968), .ZN(
        P1_U3238) );
  OAI211_X1 U16011 ( .C1(n13973), .C2(n13972), .A(n13971), .B(n13994), .ZN(
        n13982) );
  INV_X1 U16012 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n13974) );
  OAI22_X1 U16013 ( .A1(n14926), .A2(n14088), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13974), .ZN(n13976) );
  NOR2_X1 U16014 ( .A1(n14925), .A2(n6897), .ZN(n13975) );
  NOR2_X1 U16015 ( .A1(n13976), .A2(n13975), .ZN(n13981) );
  OR2_X1 U16016 ( .A1(n14941), .A2(n13977), .ZN(n13980) );
  OR2_X1 U16017 ( .A1(n14005), .A2(n13978), .ZN(n13979) );
  NAND4_X1 U16018 ( .A1(n13982), .A2(n13981), .A3(n13980), .A4(n13979), .ZN(
        P1_U3239) );
  XOR2_X1 U16019 ( .A(n13984), .B(n13983), .Z(n13992) );
  INV_X1 U16020 ( .A(n14407), .ZN(n13989) );
  OAI22_X1 U16021 ( .A1(n13986), .A2(n14531), .B1(n13985), .B2(n14533), .ZN(
        n14404) );
  AOI22_X1 U16022 ( .A1(n13987), .A2(n14404), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13988) );
  OAI21_X1 U16023 ( .B1(n14941), .B2(n13989), .A(n13988), .ZN(n13990) );
  AOI21_X1 U16024 ( .B1(n14614), .B2(n14937), .A(n13990), .ZN(n13991) );
  OAI21_X1 U16025 ( .B1(n13992), .B2(n14932), .A(n13991), .ZN(P1_U3240) );
  OAI211_X1 U16026 ( .C1(n13996), .C2(n13995), .A(n13993), .B(n13994), .ZN(
        n14004) );
  NAND2_X1 U16027 ( .A1(n13997), .A2(n14266), .ZN(n13998) );
  NAND2_X1 U16028 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n15054)
         );
  OAI211_X1 U16029 ( .C1(n13999), .C2(n14925), .A(n13998), .B(n15054), .ZN(
        n14000) );
  AOI21_X1 U16030 ( .B1(n14002), .B2(n14001), .A(n14000), .ZN(n14003) );
  OAI211_X1 U16031 ( .C1(n14006), .C2(n14005), .A(n14004), .B(n14003), .ZN(
        P1_U3241) );
  NAND2_X1 U16032 ( .A1(n14007), .A2(n14579), .ZN(n14009) );
  INV_X1 U16033 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n14015) );
  NAND2_X1 U16034 ( .A1(n14011), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n14014) );
  NAND2_X1 U16035 ( .A1(n14012), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n14013) );
  OAI211_X1 U16036 ( .C1(n14016), .C2(n14015), .A(n14014), .B(n14013), .ZN(
        n14359) );
  INV_X1 U16037 ( .A(n14359), .ZN(n14211) );
  AND2_X1 U16038 ( .A1(n6639), .A2(n14211), .ZN(n14210) );
  NAND2_X1 U16039 ( .A1(n14692), .A2(n14017), .ZN(n14019) );
  INV_X1 U16040 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n14687) );
  OR2_X1 U16041 ( .A1(n6648), .A2(n14687), .ZN(n14018) );
  NAND2_X1 U16042 ( .A1(n14187), .A2(n14359), .ZN(n14206) );
  NAND2_X1 U16043 ( .A1(n14007), .A2(n14020), .ZN(n14021) );
  NAND2_X1 U16044 ( .A1(n14022), .A2(n14021), .ZN(n14024) );
  AND2_X1 U16045 ( .A1(n14024), .A2(n14023), .ZN(n14214) );
  OAI21_X1 U16046 ( .B1(n14361), .B2(n14206), .A(n14214), .ZN(n14205) );
  OR2_X1 U16047 ( .A1(n14026), .A2(n14025), .ZN(n14029) );
  OR2_X1 U16048 ( .A1(n6649), .A2(n14027), .ZN(n14028) );
  INV_X1 U16049 ( .A(n14030), .ZN(n14031) );
  OAI21_X1 U16050 ( .B1(n14359), .B2(n14031), .A(n14260), .ZN(n14032) );
  MUX2_X1 U16051 ( .A(n14366), .B(n14032), .S(n14187), .Z(n14200) );
  INV_X1 U16052 ( .A(n14200), .ZN(n14204) );
  MUX2_X1 U16053 ( .A(n14271), .B(n14097), .S(n6639), .Z(n14102) );
  NAND3_X1 U16054 ( .A1(n14041), .A2(n14033), .A3(n14044), .ZN(n14037) );
  INV_X1 U16055 ( .A(n14033), .ZN(n14035) );
  NAND3_X1 U16056 ( .A1(n14035), .A2(n6639), .A3(n14034), .ZN(n14036) );
  NAND2_X1 U16057 ( .A1(n14037), .A2(n14036), .ZN(n14040) );
  NAND2_X1 U16058 ( .A1(n14219), .A2(n14038), .ZN(n14039) );
  MUX2_X1 U16059 ( .A(n14034), .B(n14041), .S(n14198), .Z(n14042) );
  NOR2_X1 U16060 ( .A1(n14044), .A2(n6840), .ZN(n14046) );
  AND2_X1 U16061 ( .A1(n14044), .A2(n6840), .ZN(n14045) );
  MUX2_X1 U16062 ( .A(n14053), .B(n14278), .S(n14044), .Z(n14057) );
  NAND2_X1 U16063 ( .A1(n14056), .A2(n14057), .ZN(n14055) );
  MUX2_X1 U16064 ( .A(n14278), .B(n14053), .S(n14187), .Z(n14054) );
  NAND2_X1 U16065 ( .A1(n14055), .A2(n14054), .ZN(n14061) );
  INV_X1 U16066 ( .A(n14056), .ZN(n14059) );
  INV_X1 U16067 ( .A(n14057), .ZN(n14058) );
  NAND2_X1 U16068 ( .A1(n14059), .A2(n14058), .ZN(n14060) );
  MUX2_X1 U16069 ( .A(n14277), .B(n14062), .S(n14187), .Z(n14066) );
  NAND2_X1 U16070 ( .A1(n14065), .A2(n14066), .ZN(n14064) );
  MUX2_X1 U16071 ( .A(n14062), .B(n14277), .S(n14187), .Z(n14063) );
  NAND2_X1 U16072 ( .A1(n14064), .A2(n14063), .ZN(n14070) );
  INV_X1 U16073 ( .A(n14065), .ZN(n14068) );
  INV_X1 U16074 ( .A(n14066), .ZN(n14067) );
  MUX2_X1 U16075 ( .A(n14071), .B(n14276), .S(n14187), .Z(n14073) );
  MUX2_X1 U16076 ( .A(n14276), .B(n14071), .S(n14187), .Z(n14072) );
  MUX2_X1 U16077 ( .A(n14074), .B(n14274), .S(n14187), .Z(n14086) );
  XNOR2_X1 U16078 ( .A(n14075), .B(n14273), .ZN(n14090) );
  NAND3_X1 U16079 ( .A1(n14091), .A2(n14086), .A3(n14090), .ZN(n14085) );
  MUX2_X1 U16080 ( .A(n14273), .B(n14075), .S(n14187), .Z(n14077) );
  NOR2_X1 U16081 ( .A1(n14077), .A2(n14076), .ZN(n14083) );
  OAI21_X1 U16082 ( .B1(n14272), .B2(n14187), .A(n14078), .ZN(n14082) );
  OAI21_X1 U16083 ( .B1(n14198), .B2(n14080), .A(n14079), .ZN(n14081) );
  AOI22_X1 U16084 ( .A1(n14083), .A2(n14091), .B1(n14082), .B2(n14081), .ZN(
        n14084) );
  OAI21_X1 U16085 ( .B1(n14094), .B2(n14085), .A(n14084), .ZN(n14096) );
  INV_X1 U16086 ( .A(n14086), .ZN(n14093) );
  MUX2_X1 U16087 ( .A(n14088), .B(n14087), .S(n14187), .Z(n14089) );
  NAND3_X1 U16088 ( .A1(n14091), .A2(n14090), .A3(n14089), .ZN(n14092) );
  AOI21_X1 U16089 ( .B1(n14094), .B2(n14093), .A(n14092), .ZN(n14095) );
  MUX2_X1 U16090 ( .A(n14271), .B(n14097), .S(n14187), .Z(n14098) );
  NAND2_X1 U16091 ( .A1(n14099), .A2(n14098), .ZN(n14100) );
  MUX2_X1 U16092 ( .A(n14270), .B(n14938), .S(n14187), .Z(n14106) );
  MUX2_X1 U16093 ( .A(n14270), .B(n14938), .S(n6639), .Z(n14103) );
  INV_X1 U16094 ( .A(n14105), .ZN(n14108) );
  INV_X1 U16095 ( .A(n14106), .ZN(n14107) );
  NAND2_X1 U16096 ( .A1(n14108), .A2(n14107), .ZN(n14109) );
  MUX2_X1 U16097 ( .A(n14269), .B(n14738), .S(n14198), .Z(n14111) );
  MUX2_X1 U16098 ( .A(n14269), .B(n14738), .S(n14187), .Z(n14110) );
  MUX2_X1 U16099 ( .A(n14268), .B(n14112), .S(n14187), .Z(n14114) );
  MUX2_X1 U16100 ( .A(n14901), .B(n7609), .S(n14198), .Z(n14113) );
  NAND2_X1 U16101 ( .A1(n14115), .A2(n14114), .ZN(n14116) );
  AND2_X1 U16102 ( .A1(n14124), .A2(n14118), .ZN(n14121) );
  AND2_X1 U16103 ( .A1(n14123), .A2(n14119), .ZN(n14120) );
  MUX2_X1 U16104 ( .A(n14121), .B(n14120), .S(n14187), .Z(n14122) );
  MUX2_X1 U16105 ( .A(n14124), .B(n14123), .S(n14198), .Z(n14125) );
  NAND2_X1 U16106 ( .A1(n14142), .A2(n14913), .ZN(n14127) );
  NOR2_X1 U16107 ( .A1(n14921), .A2(n14187), .ZN(n14137) );
  INV_X1 U16108 ( .A(n14137), .ZN(n14126) );
  AOI21_X1 U16109 ( .B1(n14127), .B2(n14126), .A(n14565), .ZN(n14135) );
  NAND2_X1 U16110 ( .A1(n14142), .A2(n14574), .ZN(n14129) );
  AND2_X1 U16111 ( .A1(n14187), .A2(n14128), .ZN(n14138) );
  INV_X1 U16112 ( .A(n14138), .ZN(n14131) );
  AOI21_X1 U16113 ( .B1(n14129), .B2(n14131), .A(n14944), .ZN(n14134) );
  AND2_X1 U16114 ( .A1(n14198), .A2(n14574), .ZN(n14136) );
  INV_X1 U16115 ( .A(n14136), .ZN(n14130) );
  OR2_X1 U16116 ( .A1(n14921), .A2(n14130), .ZN(n14133) );
  OR2_X1 U16117 ( .A1(n14131), .A2(n14574), .ZN(n14132) );
  NAND2_X1 U16118 ( .A1(n14133), .A2(n14132), .ZN(n14141) );
  AOI21_X1 U16119 ( .B1(n14142), .B2(n14137), .A(n14136), .ZN(n14145) );
  NAND2_X1 U16120 ( .A1(n14142), .A2(n14138), .ZN(n14139) );
  OAI21_X1 U16121 ( .B1(n6639), .B2(n14574), .A(n14139), .ZN(n14140) );
  NAND2_X1 U16122 ( .A1(n14140), .A2(n14565), .ZN(n14144) );
  NAND2_X1 U16123 ( .A1(n14142), .A2(n14141), .ZN(n14143) );
  OAI211_X1 U16124 ( .C1(n14145), .C2(n14565), .A(n14144), .B(n14143), .ZN(
        n14146) );
  MUX2_X1 U16125 ( .A(n14148), .B(n14147), .S(n6639), .Z(n14149) );
  NAND2_X1 U16126 ( .A1(n14662), .A2(n14198), .ZN(n14151) );
  OR2_X1 U16127 ( .A1(n14662), .A2(n14198), .ZN(n14150) );
  MUX2_X1 U16128 ( .A(n14151), .B(n14150), .S(n14545), .Z(n14152) );
  MUX2_X1 U16129 ( .A(n14532), .B(n14518), .S(n14187), .Z(n14155) );
  MUX2_X1 U16130 ( .A(n14498), .B(n14652), .S(n14198), .Z(n14154) );
  NAND2_X1 U16131 ( .A1(n14156), .A2(n14155), .ZN(n14160) );
  MUX2_X1 U16132 ( .A(n14506), .B(n14644), .S(n6639), .Z(n14158) );
  MUX2_X1 U16133 ( .A(n14506), .B(n14644), .S(n14187), .Z(n14157) );
  INV_X1 U16134 ( .A(n14158), .ZN(n14159) );
  MUX2_X1 U16135 ( .A(n14497), .B(n14639), .S(n14187), .Z(n14165) );
  NAND2_X1 U16136 ( .A1(n14164), .A2(n14165), .ZN(n14163) );
  MUX2_X1 U16137 ( .A(n14497), .B(n14639), .S(n14198), .Z(n14162) );
  NAND2_X1 U16138 ( .A1(n14163), .A2(n14162), .ZN(n14169) );
  INV_X1 U16139 ( .A(n14164), .ZN(n14167) );
  INV_X1 U16140 ( .A(n14165), .ZN(n14166) );
  MUX2_X1 U16141 ( .A(n14470), .B(n14633), .S(n6639), .Z(n14171) );
  MUX2_X1 U16142 ( .A(n14470), .B(n14633), .S(n14187), .Z(n14170) );
  MUX2_X1 U16143 ( .A(n14423), .B(n14626), .S(n14187), .Z(n14175) );
  NAND2_X1 U16144 ( .A1(n14174), .A2(n14175), .ZN(n14173) );
  MUX2_X1 U16145 ( .A(n14423), .B(n14626), .S(n6639), .Z(n14172) );
  INV_X1 U16146 ( .A(n14174), .ZN(n14177) );
  INV_X1 U16147 ( .A(n14175), .ZN(n14176) );
  MUX2_X1 U16148 ( .A(n14264), .B(n14431), .S(n6639), .Z(n14179) );
  MUX2_X1 U16149 ( .A(n14264), .B(n14431), .S(n14187), .Z(n14178) );
  MUX2_X1 U16150 ( .A(n14424), .B(n14614), .S(n14187), .Z(n14183) );
  NAND2_X1 U16151 ( .A1(n14182), .A2(n14183), .ZN(n14181) );
  MUX2_X1 U16152 ( .A(n14424), .B(n14614), .S(n14198), .Z(n14180) );
  MUX2_X1 U16153 ( .A(n14263), .B(n14608), .S(n6639), .Z(n14186) );
  MUX2_X1 U16154 ( .A(n14263), .B(n14608), .S(n14187), .Z(n14185) );
  MUX2_X1 U16155 ( .A(n14262), .B(n14384), .S(n14187), .Z(n14188) );
  MUX2_X1 U16156 ( .A(n14262), .B(n14384), .S(n14198), .Z(n14190) );
  MUX2_X1 U16157 ( .A(n14191), .B(n14593), .S(n6639), .Z(n14192) );
  MUX2_X1 U16158 ( .A(n14191), .B(n14593), .S(n14187), .Z(n14193) );
  INV_X1 U16159 ( .A(n14260), .ZN(n14197) );
  AOI22_X1 U16160 ( .A1(n14198), .A2(n14359), .B1(n14195), .B2(n14194), .ZN(
        n14196) );
  OAI22_X1 U16161 ( .A1(n14366), .A2(n6639), .B1(n14197), .B2(n14196), .ZN(
        n14199) );
  OAI21_X1 U16162 ( .B1(n14201), .B2(n14200), .A(n14199), .ZN(n14202) );
  NAND2_X1 U16163 ( .A1(n14359), .A2(n14214), .ZN(n14207) );
  MUX2_X1 U16164 ( .A(n14214), .B(n14207), .S(n14206), .Z(n14218) );
  INV_X1 U16165 ( .A(n14214), .ZN(n14208) );
  XNOR2_X1 U16166 ( .A(n14361), .B(n14359), .ZN(n14247) );
  NAND3_X1 U16167 ( .A1(n14209), .A2(n14208), .A3(n14247), .ZN(n14217) );
  INV_X1 U16168 ( .A(n14210), .ZN(n14213) );
  NAND3_X1 U16169 ( .A1(n14213), .A2(n14211), .A3(n14214), .ZN(n14212) );
  OAI21_X1 U16170 ( .B1(n14214), .B2(n14213), .A(n14212), .ZN(n14215) );
  AOI21_X1 U16171 ( .B1(n14361), .B2(n14215), .A(n14249), .ZN(n14216) );
  NAND3_X1 U16172 ( .A1(n14221), .A2(n14220), .A3(n14219), .ZN(n14223) );
  NOR4_X1 U16173 ( .A1(n15108), .A2(n14224), .A3(n14223), .A4(n14222), .ZN(
        n14228) );
  NAND4_X1 U16174 ( .A1(n14228), .A2(n14227), .A3(n14226), .A4(n14225), .ZN(
        n14230) );
  NOR4_X1 U16175 ( .A1(n14231), .A2(n14730), .A3(n14230), .A4(n14229), .ZN(
        n14235) );
  NAND4_X1 U16176 ( .A1(n14235), .A2(n14234), .A3(n14233), .A4(n14232), .ZN(
        n14236) );
  NOR4_X1 U16177 ( .A1(n14557), .A2(n14238), .A3(n14237), .A4(n14236), .ZN(
        n14239) );
  NAND4_X1 U16178 ( .A1(n14515), .A2(n7545), .A3(n14239), .A4(n14524), .ZN(
        n14240) );
  NOR3_X1 U16179 ( .A1(n14469), .A2(n14241), .A3(n14240), .ZN(n14242) );
  NAND4_X1 U16180 ( .A1(n14420), .A2(n14242), .A3(n14440), .A4(n14455), .ZN(
        n14243) );
  NOR4_X1 U16181 ( .A1(n14373), .A2(n14398), .A3(n14410), .A4(n14243), .ZN(
        n14246) );
  XNOR2_X1 U16182 ( .A(n14587), .B(n14260), .ZN(n14244) );
  NAND4_X1 U16183 ( .A1(n14247), .A2(n14246), .A3(n14245), .A4(n14244), .ZN(
        n14248) );
  XNOR2_X1 U16184 ( .A(n14248), .B(n14352), .ZN(n14251) );
  INV_X1 U16185 ( .A(n14249), .ZN(n14250) );
  INV_X1 U16186 ( .A(n14253), .ZN(n14259) );
  NOR3_X1 U16187 ( .A1(n14255), .A2(n14254), .A3(n14531), .ZN(n14257) );
  OAI21_X1 U16188 ( .B1(n14258), .B2(n14699), .A(P1_B_REG_SCAN_IN), .ZN(n14256) );
  OAI22_X1 U16189 ( .A1(n14259), .A2(n14258), .B1(n14257), .B2(n14256), .ZN(
        P1_U3242) );
  MUX2_X1 U16190 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14359), .S(n14282), .Z(
        P1_U3591) );
  MUX2_X1 U16191 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14260), .S(n14282), .Z(
        P1_U3590) );
  MUX2_X1 U16192 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14261), .S(n14282), .Z(
        P1_U3589) );
  MUX2_X1 U16193 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14262), .S(n14282), .Z(
        P1_U3588) );
  MUX2_X1 U16194 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14263), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16195 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14424), .S(n14282), .Z(
        P1_U3586) );
  MUX2_X1 U16196 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14264), .S(n14282), .Z(
        P1_U3585) );
  MUX2_X1 U16197 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14423), .S(n14282), .Z(
        P1_U3584) );
  MUX2_X1 U16198 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14470), .S(n14282), .Z(
        P1_U3583) );
  MUX2_X1 U16199 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14497), .S(n14282), .Z(
        P1_U3582) );
  MUX2_X1 U16200 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14506), .S(n14282), .Z(
        P1_U3581) );
  MUX2_X1 U16201 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14498), .S(n14282), .Z(
        P1_U3580) );
  MUX2_X1 U16202 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14545), .S(n14282), .Z(
        P1_U3579) );
  MUX2_X1 U16203 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14265), .S(n14282), .Z(
        P1_U3578) );
  MUX2_X1 U16204 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14574), .S(n14282), .Z(
        P1_U3577) );
  MUX2_X1 U16205 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14266), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U16206 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14572), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16207 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14267), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U16208 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14268), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16209 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14269), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U16210 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14270), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U16211 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14271), .S(n14282), .Z(
        P1_U3570) );
  MUX2_X1 U16212 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14272), .S(n14282), .Z(
        P1_U3569) );
  MUX2_X1 U16213 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14273), .S(n14282), .Z(
        P1_U3568) );
  MUX2_X1 U16214 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14274), .S(n14282), .Z(
        P1_U3567) );
  MUX2_X1 U16215 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14276), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U16216 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14277), .S(n14282), .Z(
        P1_U3565) );
  MUX2_X1 U16217 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14278), .S(n14282), .Z(
        P1_U3564) );
  MUX2_X1 U16218 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14279), .S(n14282), .Z(
        P1_U3563) );
  MUX2_X1 U16219 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14280), .S(n14282), .Z(
        P1_U3562) );
  MUX2_X1 U16220 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6932), .S(n14282), .Z(
        P1_U3561) );
  MUX2_X1 U16221 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9935), .S(n14282), .Z(
        P1_U3560) );
  OAI22_X1 U16222 ( .A1(n15104), .A2(n6834), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14283), .ZN(n14284) );
  AOI21_X1 U16223 ( .B1(n14285), .B2(n15068), .A(n14284), .ZN(n14294) );
  OAI211_X1 U16224 ( .C1(n14288), .C2(n14287), .A(n15091), .B(n14286), .ZN(
        n14293) );
  OAI211_X1 U16225 ( .C1(n14291), .C2(n14290), .A(n15096), .B(n14289), .ZN(
        n14292) );
  NAND3_X1 U16226 ( .A1(n14294), .A2(n14293), .A3(n14292), .ZN(P1_U3244) );
  INV_X1 U16227 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n14295) );
  OAI22_X1 U16228 ( .A1(n15104), .A2(n7274), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14295), .ZN(n14296) );
  AOI21_X1 U16229 ( .B1(n14297), .B2(n15068), .A(n14296), .ZN(n14306) );
  OAI211_X1 U16230 ( .C1(n14300), .C2(n14299), .A(n15096), .B(n14298), .ZN(
        n14305) );
  OAI211_X1 U16231 ( .C1(n14303), .C2(n14302), .A(n15091), .B(n14301), .ZN(
        n14304) );
  NAND4_X1 U16232 ( .A1(n14307), .A2(n14306), .A3(n14305), .A4(n14304), .ZN(
        P1_U3245) );
  INV_X1 U16233 ( .A(n14308), .ZN(n14312) );
  NAND2_X1 U16234 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n14309) );
  OAI21_X1 U16235 ( .B1(n15104), .B2(n14310), .A(n14309), .ZN(n14311) );
  AOI21_X1 U16236 ( .B1(n14312), .B2(n15068), .A(n14311), .ZN(n14321) );
  OAI211_X1 U16237 ( .C1(n14315), .C2(n14314), .A(n15096), .B(n14313), .ZN(
        n14320) );
  OAI211_X1 U16238 ( .C1(n14318), .C2(n14317), .A(n15091), .B(n14316), .ZN(
        n14319) );
  NAND3_X1 U16239 ( .A1(n14321), .A2(n14320), .A3(n14319), .ZN(P1_U3246) );
  INV_X1 U16240 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n14322) );
  MUX2_X1 U16241 ( .A(P1_REG2_REG_16__SCAN_IN), .B(n14322), .S(n15067), .Z(
        n14323) );
  INV_X1 U16242 ( .A(n14323), .ZN(n15063) );
  INV_X1 U16243 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n14324) );
  MUX2_X1 U16244 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n14324), .S(n15023), .Z(
        n14325) );
  INV_X1 U16245 ( .A(n14325), .ZN(n15016) );
  OAI21_X1 U16246 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n14337), .A(n14326), 
        .ZN(n15017) );
  NOR2_X1 U16247 ( .A1(n15016), .A2(n15017), .ZN(n15015) );
  MUX2_X1 U16248 ( .A(n11412), .B(P1_REG2_REG_14__SCAN_IN), .S(n14338), .Z(
        n15029) );
  NAND2_X1 U16249 ( .A1(n14327), .A2(n15052), .ZN(n14329) );
  XNOR2_X1 U16250 ( .A(n15052), .B(n14328), .ZN(n15044) );
  INV_X1 U16251 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n15043) );
  NAND2_X1 U16252 ( .A1(n15044), .A2(n15043), .ZN(n15042) );
  NAND2_X1 U16253 ( .A1(n14329), .A2(n15042), .ZN(n15064) );
  INV_X1 U16254 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14330) );
  MUX2_X1 U16255 ( .A(n14330), .B(P1_REG2_REG_17__SCAN_IN), .S(n14343), .Z(
        n15074) );
  NOR2_X1 U16256 ( .A1(n14331), .A2(n15099), .ZN(n14332) );
  INV_X1 U16257 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n15093) );
  XNOR2_X1 U16258 ( .A(n15099), .B(n14331), .ZN(n15094) );
  NOR2_X1 U16259 ( .A1(n15093), .A2(n15094), .ZN(n15092) );
  NOR2_X1 U16260 ( .A1(n14332), .A2(n15092), .ZN(n14333) );
  XNOR2_X1 U16261 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n14333), .ZN(n14351) );
  INV_X1 U16262 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n15088) );
  INV_X1 U16263 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n14334) );
  MUX2_X1 U16264 ( .A(n14334), .B(P1_REG1_REG_16__SCAN_IN), .S(n15067), .Z(
        n15059) );
  INV_X1 U16265 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n14335) );
  MUX2_X1 U16266 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n14335), .S(n14338), .Z(
        n15033) );
  OAI21_X1 U16267 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n14337), .A(n14336), 
        .ZN(n15020) );
  MUX2_X1 U16268 ( .A(n11477), .B(P1_REG1_REG_13__SCAN_IN), .S(n15023), .Z(
        n15019) );
  NOR2_X1 U16269 ( .A1(n15020), .A2(n15019), .ZN(n15018) );
  NAND2_X1 U16270 ( .A1(n15033), .A2(n15032), .ZN(n15031) );
  OAI21_X1 U16271 ( .B1(n14338), .B2(P1_REG1_REG_14__SCAN_IN), .A(n15031), 
        .ZN(n14339) );
  NAND2_X1 U16272 ( .A1(n15052), .A2(n14339), .ZN(n14341) );
  INV_X1 U16273 ( .A(n14339), .ZN(n14340) );
  INV_X1 U16274 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n15047) );
  NAND2_X1 U16275 ( .A1(n15048), .A2(n15047), .ZN(n15046) );
  NAND2_X1 U16276 ( .A1(n14341), .A2(n15046), .ZN(n15060) );
  INV_X1 U16277 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n14342) );
  MUX2_X1 U16278 ( .A(n14342), .B(P1_REG1_REG_17__SCAN_IN), .S(n14343), .Z(
        n15078) );
  XNOR2_X1 U16279 ( .A(n15099), .B(n14344), .ZN(n15089) );
  NOR2_X1 U16280 ( .A1(n15088), .A2(n15089), .ZN(n15087) );
  NOR2_X1 U16281 ( .A1(n14344), .A2(n15099), .ZN(n14345) );
  NOR2_X1 U16282 ( .A1(n15087), .A2(n14345), .ZN(n14347) );
  INV_X1 U16283 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14346) );
  XOR2_X1 U16284 ( .A(n14347), .B(n14346), .Z(n14350) );
  INV_X1 U16285 ( .A(n14350), .ZN(n14348) );
  NAND2_X1 U16286 ( .A1(n14348), .A2(n15091), .ZN(n14349) );
  AOI22_X1 U16287 ( .A1(n14351), .A2(n15096), .B1(n15091), .B2(n14350), .ZN(
        n14353) );
  MUX2_X1 U16288 ( .A(n14354), .B(n14353), .S(n14352), .Z(n14357) );
  INV_X1 U16289 ( .A(n14355), .ZN(n14356) );
  OAI211_X1 U16290 ( .C1(n7779), .C2(n15104), .A(n14357), .B(n14356), .ZN(
        P1_U3262) );
  XOR2_X1 U16291 ( .A(n14364), .B(n14361), .Z(n14358) );
  NAND2_X1 U16292 ( .A1(n14358), .A2(n15120), .ZN(n14585) );
  NAND2_X1 U16293 ( .A1(n14360), .A2(n14359), .ZN(n14589) );
  NOR2_X1 U16294 ( .A1(n15129), .A2(n14589), .ZN(n14368) );
  INV_X1 U16295 ( .A(n14361), .ZN(n14586) );
  NOR2_X1 U16296 ( .A1(n14586), .A2(n15116), .ZN(n14362) );
  AOI211_X1 U16297 ( .C1(n15129), .C2(P1_REG2_REG_31__SCAN_IN), .A(n14368), 
        .B(n14362), .ZN(n14363) );
  OAI21_X1 U16298 ( .B1(n14585), .B2(n14519), .A(n14363), .ZN(P1_U3263) );
  OAI21_X1 U16299 ( .B1(n14366), .B2(n14365), .A(n14364), .ZN(n14590) );
  NOR2_X1 U16300 ( .A1(n14552), .A2(n14367), .ZN(n14369) );
  AOI211_X1 U16301 ( .C1(n14587), .C2(n14737), .A(n14369), .B(n14368), .ZN(
        n14370) );
  OAI21_X1 U16302 ( .B1(n14590), .B2(n14371), .A(n14370), .ZN(P1_U3264) );
  XNOR2_X1 U16303 ( .A(n14372), .B(n14373), .ZN(n14605) );
  AOI21_X1 U16304 ( .B1(n14376), .B2(n14375), .A(n14374), .ZN(n14603) );
  NAND2_X1 U16305 ( .A1(n14384), .A2(n14390), .ZN(n14377) );
  NAND2_X1 U16306 ( .A1(n14377), .A2(n15120), .ZN(n14378) );
  NOR2_X1 U16307 ( .A1(n14379), .A2(n14378), .ZN(n14602) );
  NAND2_X1 U16308 ( .A1(n14602), .A2(n15125), .ZN(n14386) );
  NAND2_X1 U16309 ( .A1(n15129), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n14382) );
  NAND2_X1 U16310 ( .A1(n15114), .A2(n14380), .ZN(n14381) );
  OAI211_X1 U16311 ( .C1(n15129), .C2(n14599), .A(n14382), .B(n14381), .ZN(
        n14383) );
  AOI21_X1 U16312 ( .B1(n14384), .B2(n14737), .A(n14383), .ZN(n14385) );
  NAND2_X1 U16313 ( .A1(n14386), .A2(n14385), .ZN(n14387) );
  AOI21_X1 U16314 ( .B1(n14603), .B2(n14516), .A(n14387), .ZN(n14388) );
  OAI21_X1 U16315 ( .B1(n14605), .B2(n14483), .A(n14388), .ZN(P1_U3265) );
  XNOR2_X1 U16316 ( .A(n14389), .B(n14398), .ZN(n14612) );
  AOI211_X1 U16317 ( .C1(n14608), .C2(n14406), .A(n15161), .B(n14391), .ZN(
        n14606) );
  INV_X1 U16318 ( .A(n14608), .ZN(n14395) );
  AOI22_X1 U16319 ( .A1(n14552), .A2(n14607), .B1(n14392), .B2(n15114), .ZN(
        n14394) );
  NAND2_X1 U16320 ( .A1(n15129), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n14393) );
  OAI211_X1 U16321 ( .C1(n14395), .C2(n15116), .A(n14394), .B(n14393), .ZN(
        n14396) );
  AOI21_X1 U16322 ( .B1(n14606), .B2(n15125), .A(n14396), .ZN(n14401) );
  OAI21_X1 U16323 ( .B1(n14399), .B2(n14398), .A(n14397), .ZN(n14609) );
  NAND2_X1 U16324 ( .A1(n14609), .A2(n14516), .ZN(n14400) );
  OAI211_X1 U16325 ( .C1(n14612), .C2(n14483), .A(n14401), .B(n14400), .ZN(
        P1_U3266) );
  XNOR2_X1 U16326 ( .A(n14403), .B(n14402), .ZN(n14405) );
  AOI21_X1 U16327 ( .B1(n14405), .B2(n14971), .A(n14404), .ZN(n14616) );
  AOI211_X1 U16328 ( .C1(n14614), .C2(n14421), .A(n15161), .B(n7210), .ZN(
        n14613) );
  INV_X1 U16329 ( .A(n14614), .ZN(n14409) );
  AOI22_X1 U16330 ( .A1(n15129), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n14407), 
        .B2(n15114), .ZN(n14408) );
  OAI21_X1 U16331 ( .B1(n14409), .B2(n15116), .A(n14408), .ZN(n14413) );
  XNOR2_X1 U16332 ( .A(n14411), .B(n14410), .ZN(n14617) );
  NOR2_X1 U16333 ( .A1(n14617), .A2(n14584), .ZN(n14412) );
  AOI211_X1 U16334 ( .C1(n14613), .C2(n15125), .A(n14413), .B(n14412), .ZN(
        n14414) );
  OAI21_X1 U16335 ( .B1(n14616), .B2(n15129), .A(n14414), .ZN(P1_U3267) );
  OAI21_X1 U16336 ( .B1(n14417), .B2(n14416), .A(n14415), .ZN(n14624) );
  OAI21_X1 U16337 ( .B1(n7618), .B2(n14420), .A(n14419), .ZN(n14622) );
  AOI21_X1 U16338 ( .B1(n14431), .B2(n14443), .A(n15161), .ZN(n14422) );
  NAND2_X1 U16339 ( .A1(n14422), .A2(n14421), .ZN(n14619) );
  NAND2_X1 U16340 ( .A1(n14423), .A2(n14571), .ZN(n14426) );
  NAND2_X1 U16341 ( .A1(n14424), .A2(n14573), .ZN(n14425) );
  AND2_X1 U16342 ( .A1(n14426), .A2(n14425), .ZN(n14618) );
  NAND2_X1 U16343 ( .A1(n15129), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n14429) );
  NAND2_X1 U16344 ( .A1(n15114), .A2(n14427), .ZN(n14428) );
  OAI211_X1 U16345 ( .C1(n15129), .C2(n14618), .A(n14429), .B(n14428), .ZN(
        n14430) );
  AOI21_X1 U16346 ( .B1(n14431), .B2(n14737), .A(n14430), .ZN(n14432) );
  OAI21_X1 U16347 ( .B1(n14619), .B2(n14519), .A(n14432), .ZN(n14433) );
  AOI21_X1 U16348 ( .B1(n14622), .B2(n14505), .A(n14433), .ZN(n14434) );
  OAI21_X1 U16349 ( .B1(n14584), .B2(n14624), .A(n14434), .ZN(P1_U3268) );
  AOI21_X1 U16350 ( .B1(n14436), .B2(n14435), .A(n15109), .ZN(n14439) );
  AOI21_X1 U16351 ( .B1(n14439), .B2(n14438), .A(n14437), .ZN(n14628) );
  AND2_X1 U16352 ( .A1(n14441), .A2(n14440), .ZN(n14442) );
  NOR2_X1 U16353 ( .A1(n6692), .A2(n14442), .ZN(n14629) );
  INV_X1 U16354 ( .A(n14629), .ZN(n14450) );
  AOI21_X1 U16355 ( .B1(n14626), .B2(n14453), .A(n15161), .ZN(n14444) );
  AND2_X1 U16356 ( .A1(n14444), .A2(n14443), .ZN(n14625) );
  NAND2_X1 U16357 ( .A1(n14625), .A2(n15125), .ZN(n14447) );
  AOI22_X1 U16358 ( .A1(n15129), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n14445), 
        .B2(n15114), .ZN(n14446) );
  OAI211_X1 U16359 ( .C1(n14448), .C2(n15116), .A(n14447), .B(n14446), .ZN(
        n14449) );
  AOI21_X1 U16360 ( .B1(n14450), .B2(n14516), .A(n14449), .ZN(n14451) );
  OAI21_X1 U16361 ( .B1(n14628), .B2(n15129), .A(n14451), .ZN(P1_U3269) );
  XNOR2_X1 U16362 ( .A(n14452), .B(n14455), .ZN(n14636) );
  INV_X1 U16363 ( .A(n14480), .ZN(n14454) );
  AOI211_X1 U16364 ( .C1(n14633), .C2(n14454), .A(n15161), .B(n7205), .ZN(
        n14631) );
  INV_X1 U16365 ( .A(n14631), .ZN(n14458) );
  XNOR2_X1 U16366 ( .A(n14456), .B(n14455), .ZN(n14457) );
  NAND2_X1 U16367 ( .A1(n14457), .A2(n14971), .ZN(n14635) );
  OAI211_X1 U16368 ( .C1(n14579), .C2(n14458), .A(n14635), .B(n14630), .ZN(
        n14463) );
  AOI22_X1 U16369 ( .A1(n15129), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n14459), 
        .B2(n15114), .ZN(n14460) );
  OAI21_X1 U16370 ( .B1(n14461), .B2(n15116), .A(n14460), .ZN(n14462) );
  AOI21_X1 U16371 ( .B1(n14463), .B2(n14552), .A(n14462), .ZN(n14464) );
  OAI21_X1 U16372 ( .B1(n14584), .B2(n14636), .A(n14464), .ZN(P1_U3270) );
  XNOR2_X1 U16373 ( .A(n14465), .B(n14469), .ZN(n14640) );
  INV_X1 U16374 ( .A(n14466), .ZN(n14467) );
  AOI21_X1 U16375 ( .B1(n14469), .B2(n14468), .A(n14467), .ZN(n14643) );
  NAND2_X1 U16376 ( .A1(n14506), .A2(n14571), .ZN(n14472) );
  NAND2_X1 U16377 ( .A1(n14470), .A2(n14573), .ZN(n14471) );
  NAND2_X1 U16378 ( .A1(n14472), .A2(n14471), .ZN(n14638) );
  INV_X1 U16379 ( .A(n14638), .ZN(n14476) );
  NAND2_X1 U16380 ( .A1(n15129), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n14475) );
  NAND2_X1 U16381 ( .A1(n15114), .A2(n14473), .ZN(n14474) );
  OAI211_X1 U16382 ( .C1(n15129), .C2(n14476), .A(n14475), .B(n14474), .ZN(
        n14477) );
  AOI21_X1 U16383 ( .B1(n14639), .B2(n14737), .A(n14477), .ZN(n14482) );
  NAND2_X1 U16384 ( .A1(n14489), .A2(n14639), .ZN(n14478) );
  NAND2_X1 U16385 ( .A1(n14478), .A2(n15120), .ZN(n14479) );
  NOR2_X1 U16386 ( .A1(n14480), .A2(n14479), .ZN(n14637) );
  NAND2_X1 U16387 ( .A1(n14637), .A2(n15125), .ZN(n14481) );
  OAI211_X1 U16388 ( .C1(n14643), .C2(n14483), .A(n14482), .B(n14481), .ZN(
        n14484) );
  AOI21_X1 U16389 ( .B1(n14516), .B2(n14640), .A(n14484), .ZN(n14485) );
  INV_X1 U16390 ( .A(n14485), .ZN(P1_U3271) );
  NAND2_X1 U16391 ( .A1(n14486), .A2(n14495), .ZN(n14487) );
  INV_X1 U16392 ( .A(n14489), .ZN(n14490) );
  AOI21_X1 U16393 ( .B1(n14644), .B2(n14517), .A(n14490), .ZN(n14645) );
  INV_X1 U16394 ( .A(n14644), .ZN(n14493) );
  AOI22_X1 U16395 ( .A1(n15129), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n14491), 
        .B2(n15114), .ZN(n14492) );
  OAI21_X1 U16396 ( .B1(n14493), .B2(n15116), .A(n14492), .ZN(n14502) );
  OAI211_X1 U16397 ( .C1(n14496), .C2(n14495), .A(n14494), .B(n14971), .ZN(
        n14500) );
  AOI22_X1 U16398 ( .A1(n14498), .A2(n14571), .B1(n14573), .B2(n14497), .ZN(
        n14499) );
  AND2_X1 U16399 ( .A1(n14500), .A2(n14499), .ZN(n14647) );
  NOR2_X1 U16400 ( .A1(n14647), .A2(n15129), .ZN(n14501) );
  AOI211_X1 U16401 ( .C1(n14645), .C2(n14503), .A(n14502), .B(n14501), .ZN(
        n14504) );
  OAI21_X1 U16402 ( .B1(n14648), .B2(n14584), .A(n14504), .ZN(P1_U3272) );
  OR2_X1 U16403 ( .A1(n6764), .A2(n14515), .ZN(n14650) );
  NAND3_X1 U16404 ( .A1(n14650), .A2(n14649), .A3(n14505), .ZN(n14523) );
  NAND2_X1 U16405 ( .A1(n14545), .A2(n14571), .ZN(n14508) );
  NAND2_X1 U16406 ( .A1(n14506), .A2(n14573), .ZN(n14507) );
  NAND2_X1 U16407 ( .A1(n14508), .A2(n14507), .ZN(n14651) );
  INV_X1 U16408 ( .A(n14651), .ZN(n14512) );
  NAND2_X1 U16409 ( .A1(n15129), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n14511) );
  NAND2_X1 U16410 ( .A1(n15114), .A2(n14509), .ZN(n14510) );
  OAI211_X1 U16411 ( .C1(n15129), .C2(n14512), .A(n14511), .B(n14510), .ZN(
        n14513) );
  AOI21_X1 U16412 ( .B1(n14652), .B2(n14737), .A(n14513), .ZN(n14522) );
  NAND2_X1 U16413 ( .A1(n14514), .A2(n14515), .ZN(n14653) );
  NAND3_X1 U16414 ( .A1(n14654), .A2(n14653), .A3(n14516), .ZN(n14521) );
  OAI211_X1 U16415 ( .C1(n14518), .C2(n14535), .A(n15120), .B(n14517), .ZN(
        n14655) );
  OR2_X1 U16416 ( .A1(n14655), .A2(n14519), .ZN(n14520) );
  NAND4_X1 U16417 ( .A1(n14523), .A2(n14522), .A3(n14521), .A4(n14520), .ZN(
        P1_U3273) );
  XNOR2_X1 U16418 ( .A(n14525), .B(n14524), .ZN(n14664) );
  AOI21_X1 U16419 ( .B1(n14528), .B2(n14527), .A(n14526), .ZN(n14529) );
  OAI222_X1 U16420 ( .A1(n14533), .A2(n14532), .B1(n14531), .B2(n14530), .C1(
        n15109), .C2(n14529), .ZN(n14660) );
  OAI21_X1 U16421 ( .B1(n14548), .B2(n14534), .A(n15120), .ZN(n14536) );
  OR2_X1 U16422 ( .A1(n14536), .A2(n14535), .ZN(n14659) );
  OAI22_X1 U16423 ( .A1(n14659), .A2(n14579), .B1(n14578), .B2(n14537), .ZN(
        n14538) );
  OAI21_X1 U16424 ( .B1(n14660), .B2(n14538), .A(n14552), .ZN(n14540) );
  AOI22_X1 U16425 ( .A1(n14662), .A2(n14737), .B1(P1_REG2_REG_19__SCAN_IN), 
        .B2(n15129), .ZN(n14539) );
  OAI211_X1 U16426 ( .C1(n14664), .C2(n14584), .A(n14540), .B(n14539), .ZN(
        P1_U3274) );
  XNOR2_X1 U16427 ( .A(n14542), .B(n14541), .ZN(n14669) );
  OAI211_X1 U16428 ( .C1(n14544), .C2(n7545), .A(n14543), .B(n14971), .ZN(
        n14547) );
  AOI22_X1 U16429 ( .A1(n14571), .A2(n14574), .B1(n14545), .B2(n14573), .ZN(
        n14546) );
  NAND2_X1 U16430 ( .A1(n14547), .A2(n14546), .ZN(n14665) );
  AOI211_X1 U16431 ( .C1(n14667), .C2(n6765), .A(n15161), .B(n14548), .ZN(
        n14666) );
  INV_X1 U16432 ( .A(n14666), .ZN(n14551) );
  INV_X1 U16433 ( .A(n14549), .ZN(n14550) );
  OAI22_X1 U16434 ( .A1(n14551), .A2(n14579), .B1(n14578), .B2(n14550), .ZN(
        n14553) );
  OAI21_X1 U16435 ( .B1(n14665), .B2(n14553), .A(n14552), .ZN(n14555) );
  AOI22_X1 U16436 ( .A1(n14667), .A2(n14737), .B1(n15129), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n14554) );
  OAI211_X1 U16437 ( .C1(n14584), .C2(n14669), .A(n14555), .B(n14554), .ZN(
        P1_U3275) );
  XOR2_X1 U16438 ( .A(n14557), .B(n14556), .Z(n14942) );
  OAI211_X1 U16439 ( .C1(n7678), .C2(n11781), .A(n14971), .B(n14558), .ZN(
        n14560) );
  NAND2_X1 U16440 ( .A1(n14560), .A2(n14559), .ZN(n14945) );
  AOI21_X1 U16441 ( .B1(n14576), .B2(n14565), .A(n15161), .ZN(n14561) );
  NAND2_X1 U16442 ( .A1(n14561), .A2(n6765), .ZN(n14943) );
  INV_X1 U16443 ( .A(n14562), .ZN(n14563) );
  OAI22_X1 U16444 ( .A1(n14943), .A2(n14579), .B1(n14578), .B2(n14563), .ZN(
        n14564) );
  OAI21_X1 U16445 ( .B1(n14945), .B2(n14564), .A(n14552), .ZN(n14567) );
  AOI22_X1 U16446 ( .A1(n14565), .A2(n14737), .B1(n15129), .B2(
        P1_REG2_REG_17__SCAN_IN), .ZN(n14566) );
  OAI211_X1 U16447 ( .C1(n14942), .C2(n14584), .A(n14567), .B(n14566), .ZN(
        P1_U3276) );
  XNOR2_X1 U16448 ( .A(n14568), .B(n14570), .ZN(n14948) );
  OAI21_X1 U16449 ( .B1(n6746), .B2(n14570), .A(n14569), .ZN(n14575) );
  AOI222_X1 U16450 ( .A1(n14971), .A2(n14575), .B1(n14574), .B2(n14573), .C1(
        n14572), .C2(n14571), .ZN(n14950) );
  INV_X1 U16451 ( .A(n14950), .ZN(n14581) );
  OAI211_X1 U16452 ( .C1(n14577), .C2(n14951), .A(n15120), .B(n14576), .ZN(
        n14949) );
  OAI22_X1 U16453 ( .A1(n14949), .A2(n14579), .B1(n14578), .B2(n14923), .ZN(
        n14580) );
  OAI21_X1 U16454 ( .B1(n14581), .B2(n14580), .A(n14552), .ZN(n14583) );
  AOI22_X1 U16455 ( .A1(n14921), .A2(n14737), .B1(n15129), .B2(
        P1_REG2_REG_16__SCAN_IN), .ZN(n14582) );
  OAI211_X1 U16456 ( .C1(n14948), .C2(n14584), .A(n14583), .B(n14582), .ZN(
        P1_U3277) );
  OAI211_X1 U16457 ( .C1(n14586), .C2(n15187), .A(n14585), .B(n14589), .ZN(
        n14672) );
  MUX2_X1 U16458 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14672), .S(n15202), .Z(
        P1_U3559) );
  NAND2_X1 U16459 ( .A1(n14587), .A2(n14955), .ZN(n14588) );
  OAI211_X1 U16460 ( .C1(n14590), .C2(n15161), .A(n14589), .B(n14588), .ZN(
        n14673) );
  MUX2_X1 U16461 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14673), .S(n15202), .Z(
        P1_U3558) );
  OAI211_X1 U16462 ( .C1(n14593), .C2(n15187), .A(n14592), .B(n14591), .ZN(
        n14594) );
  AOI21_X1 U16463 ( .B1(n14595), .B2(n15120), .A(n14594), .ZN(n14596) );
  OAI21_X1 U16464 ( .B1(n14600), .B2(n15187), .A(n14599), .ZN(n14601) );
  OAI21_X1 U16465 ( .B1(n14605), .B2(n15109), .A(n14604), .ZN(n14675) );
  MUX2_X1 U16466 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14675), .S(n15202), .Z(
        P1_U3556) );
  NAND2_X1 U16467 ( .A1(n14609), .A2(n15191), .ZN(n14610) );
  OAI211_X1 U16468 ( .C1(n14612), .C2(n15109), .A(n14611), .B(n14610), .ZN(
        n14676) );
  MUX2_X1 U16469 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14676), .S(n15202), .Z(
        P1_U3555) );
  AOI21_X1 U16470 ( .B1(n14614), .B2(n14955), .A(n14613), .ZN(n14615) );
  OAI211_X1 U16471 ( .C1(n14670), .C2(n14617), .A(n14616), .B(n14615), .ZN(
        n14677) );
  MUX2_X1 U16472 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14677), .S(n15202), .Z(
        P1_U3554) );
  OAI211_X1 U16473 ( .C1(n14620), .C2(n15187), .A(n14619), .B(n14618), .ZN(
        n14621) );
  AOI21_X1 U16474 ( .B1(n14622), .B2(n14971), .A(n14621), .ZN(n14623) );
  OAI21_X1 U16475 ( .B1(n14670), .B2(n14624), .A(n14623), .ZN(n14678) );
  MUX2_X1 U16476 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14678), .S(n15202), .Z(
        P1_U3553) );
  AOI21_X1 U16477 ( .B1(n14626), .B2(n14955), .A(n14625), .ZN(n14627) );
  OAI211_X1 U16478 ( .C1(n14670), .C2(n14629), .A(n14628), .B(n14627), .ZN(
        n14679) );
  MUX2_X1 U16479 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14679), .S(n15202), .Z(
        P1_U3552) );
  INV_X1 U16480 ( .A(n14630), .ZN(n14632) );
  AOI211_X1 U16481 ( .C1(n14633), .C2(n14955), .A(n14632), .B(n14631), .ZN(
        n14634) );
  OAI211_X1 U16482 ( .C1(n14670), .C2(n14636), .A(n14635), .B(n14634), .ZN(
        n14680) );
  MUX2_X1 U16483 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14680), .S(n15202), .Z(
        P1_U3551) );
  AOI211_X1 U16484 ( .C1(n14639), .C2(n14955), .A(n14638), .B(n14637), .ZN(
        n14642) );
  NAND2_X1 U16485 ( .A1(n14640), .A2(n15191), .ZN(n14641) );
  OAI211_X1 U16486 ( .C1(n14643), .C2(n15109), .A(n14642), .B(n14641), .ZN(
        n14681) );
  MUX2_X1 U16487 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14681), .S(n15202), .Z(
        P1_U3550) );
  AOI22_X1 U16488 ( .A1(n14645), .A2(n15120), .B1(n14644), .B2(n14955), .ZN(
        n14646) );
  OAI211_X1 U16489 ( .C1(n14670), .C2(n14648), .A(n14647), .B(n14646), .ZN(
        n14682) );
  MUX2_X1 U16490 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14682), .S(n15202), .Z(
        P1_U3549) );
  NAND3_X1 U16491 ( .A1(n14650), .A2(n14649), .A3(n14971), .ZN(n14658) );
  AOI21_X1 U16492 ( .B1(n14652), .B2(n14955), .A(n14651), .ZN(n14657) );
  NAND3_X1 U16493 ( .A1(n14654), .A2(n14653), .A3(n15191), .ZN(n14656) );
  NAND4_X1 U16494 ( .A1(n14658), .A2(n14657), .A3(n14656), .A4(n14655), .ZN(
        n14683) );
  MUX2_X1 U16495 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14683), .S(n15202), .Z(
        P1_U3548) );
  INV_X1 U16496 ( .A(n14659), .ZN(n14661) );
  AOI211_X1 U16497 ( .C1(n14662), .C2(n14955), .A(n14661), .B(n14660), .ZN(
        n14663) );
  OAI21_X1 U16498 ( .B1(n14670), .B2(n14664), .A(n14663), .ZN(n14684) );
  MUX2_X1 U16499 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14684), .S(n15202), .Z(
        P1_U3547) );
  AOI211_X1 U16500 ( .C1(n14667), .C2(n14955), .A(n14666), .B(n14665), .ZN(
        n14668) );
  OAI21_X1 U16501 ( .B1(n14670), .B2(n14669), .A(n14668), .ZN(n14685) );
  MUX2_X1 U16502 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14685), .S(n15202), .Z(
        P1_U3546) );
  MUX2_X1 U16503 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n14671), .S(n15202), .Z(
        P1_U3528) );
  MUX2_X1 U16504 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14672), .S(n15194), .Z(
        P1_U3527) );
  MUX2_X1 U16505 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14673), .S(n15194), .Z(
        P1_U3526) );
  MUX2_X1 U16506 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14674), .S(n15194), .Z(
        P1_U3525) );
  MUX2_X1 U16507 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14675), .S(n15194), .Z(
        P1_U3524) );
  MUX2_X1 U16508 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14676), .S(n15194), .Z(
        P1_U3523) );
  MUX2_X1 U16509 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14677), .S(n15194), .Z(
        P1_U3522) );
  MUX2_X1 U16510 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14678), .S(n15194), .Z(
        P1_U3521) );
  MUX2_X1 U16511 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14679), .S(n15194), .Z(
        P1_U3520) );
  MUX2_X1 U16512 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14680), .S(n15194), .Z(
        P1_U3519) );
  MUX2_X1 U16513 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14681), .S(n15194), .Z(
        P1_U3518) );
  MUX2_X1 U16514 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14682), .S(n15194), .Z(
        P1_U3517) );
  MUX2_X1 U16515 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14683), .S(n15194), .Z(
        P1_U3516) );
  MUX2_X1 U16516 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14684), .S(n15194), .Z(
        P1_U3515) );
  MUX2_X1 U16517 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14685), .S(n15194), .Z(
        P1_U3513) );
  NAND3_X1 U16518 ( .A1(n14686), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n14688) );
  OAI22_X1 U16519 ( .A1(n14689), .A2(n14688), .B1(n14687), .B2(n14694), .ZN(
        n14690) );
  AOI21_X1 U16520 ( .B1(n14692), .B2(n14691), .A(n14690), .ZN(n14693) );
  INV_X1 U16521 ( .A(n14693), .ZN(P1_U3324) );
  OAI222_X1 U16522 ( .A1(n11910), .A2(n14697), .B1(P1_U3086), .B2(n14696), 
        .C1(n14695), .C2(n14694), .ZN(P1_U3329) );
  MUX2_X1 U16523 ( .A(n14699), .B(n14698), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U16524 ( .A(n14700), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AOI21_X1 U16525 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14704) );
  OAI21_X1 U16526 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14704), 
        .ZN(U28) );
  AOI21_X1 U16527 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14705) );
  OAI21_X1 U16528 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14705), 
        .ZN(U29) );
  OAI21_X1 U16529 ( .B1(n14708), .B2(n14707), .A(n14706), .ZN(n14709) );
  XNOR2_X1 U16530 ( .A(n14709), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  AOI21_X1 U16531 ( .B1(n14712), .B2(n14711), .A(n14710), .ZN(SUB_1596_U57) );
  AOI21_X1 U16532 ( .B1(n14715), .B2(n14714), .A(n14713), .ZN(n14716) );
  XOR2_X1 U16533 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n14716), .Z(SUB_1596_U55) );
  AOI21_X1 U16534 ( .B1(n14719), .B2(n14718), .A(n14717), .ZN(n14720) );
  XOR2_X1 U16535 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n14720), .Z(SUB_1596_U54) );
  OAI22_X1 U16536 ( .A1(n14723), .A2(n14722), .B1(SI_22_), .B2(n14721), .ZN(
        n14724) );
  AOI21_X1 U16537 ( .B1(P3_STATE_REG_SCAN_IN), .B2(n14725), .A(n14724), .ZN(
        P3_U3273) );
  AOI21_X1 U16538 ( .B1(n14728), .B2(n14727), .A(n14726), .ZN(n14729) );
  XOR2_X1 U16539 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n14729), .Z(SUB_1596_U70)
         );
  XNOR2_X1 U16540 ( .A(n14731), .B(n14730), .ZN(n14750) );
  XNOR2_X1 U16541 ( .A(n14732), .B(n7384), .ZN(n14734) );
  OAI21_X1 U16542 ( .B1(n14734), .B2(n15109), .A(n14733), .ZN(n14735) );
  AOI21_X1 U16543 ( .B1(n15183), .B2(n14750), .A(n14735), .ZN(n14747) );
  AOI222_X1 U16544 ( .A1(n14738), .A2(n14737), .B1(n14736), .B2(n15114), .C1(
        P1_REG2_REG_12__SCAN_IN), .C2(n15129), .ZN(n14744) );
  INV_X1 U16545 ( .A(n14739), .ZN(n14741) );
  OAI211_X1 U16546 ( .C1(n14741), .C2(n14746), .A(n15120), .B(n14740), .ZN(
        n14745) );
  INV_X1 U16547 ( .A(n14745), .ZN(n14742) );
  AOI22_X1 U16548 ( .A1(n14750), .A2(n15126), .B1(n15125), .B2(n14742), .ZN(
        n14743) );
  OAI211_X1 U16549 ( .C1(n15129), .C2(n14747), .A(n14744), .B(n14743), .ZN(
        P1_U3281) );
  OAI21_X1 U16550 ( .B1(n14746), .B2(n15187), .A(n14745), .ZN(n14749) );
  INV_X1 U16551 ( .A(n14747), .ZN(n14748) );
  AOI211_X1 U16552 ( .C1(n15173), .C2(n14750), .A(n14749), .B(n14748), .ZN(
        n14753) );
  INV_X1 U16553 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14751) );
  AOI22_X1 U16554 ( .A1(n15194), .A2(n14753), .B1(n14751), .B2(n15192), .ZN(
        P1_U3495) );
  AOI22_X1 U16555 ( .A1(n15202), .A2(n14753), .B1(n14752), .B2(n15200), .ZN(
        P1_U3540) );
  AOI21_X1 U16556 ( .B1(n14756), .B2(n14755), .A(n14754), .ZN(n14757) );
  XOR2_X1 U16557 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n14757), .Z(SUB_1596_U63)
         );
  XNOR2_X1 U16558 ( .A(n14758), .B(n7451), .ZN(n14797) );
  XNOR2_X1 U16559 ( .A(n14760), .B(n14759), .ZN(n14761) );
  OAI222_X1 U16560 ( .A1(n15448), .A2(n14763), .B1(n15450), .B2(n14762), .C1(
        n14761), .C2(n15456), .ZN(n14795) );
  AOI21_X1 U16561 ( .B1(n14797), .B2(n14779), .A(n14795), .ZN(n14767) );
  NOR2_X1 U16562 ( .A1(n14764), .A2(n15521), .ZN(n14796) );
  AOI22_X1 U16563 ( .A1(n14782), .A2(n14796), .B1(n15473), .B2(n14765), .ZN(
        n14766) );
  OAI221_X1 U16564 ( .B1(n12871), .B2(n14767), .C1(n15477), .C2(n11868), .A(
        n14766), .ZN(P3_U3220) );
  XNOR2_X1 U16565 ( .A(n14769), .B(n14768), .ZN(n14801) );
  NAND2_X1 U16566 ( .A1(n14771), .A2(n14770), .ZN(n14773) );
  NAND2_X1 U16567 ( .A1(n14773), .A2(n14772), .ZN(n14775) );
  XNOR2_X1 U16568 ( .A(n14775), .B(n14774), .ZN(n14776) );
  OAI222_X1 U16569 ( .A1(n15448), .A2(n14778), .B1(n15450), .B2(n14777), .C1(
        n14776), .C2(n15456), .ZN(n14799) );
  AOI21_X1 U16570 ( .B1(n14801), .B2(n14779), .A(n14799), .ZN(n14785) );
  NOR2_X1 U16571 ( .A1(n14780), .A2(n15521), .ZN(n14800) );
  AOI22_X1 U16572 ( .A1(n14782), .A2(n14800), .B1(n15473), .B2(n14781), .ZN(
        n14783) );
  OAI221_X1 U16573 ( .B1(n12871), .B2(n14785), .C1(n15477), .C2(n14784), .A(
        n14783), .ZN(P3_U3221) );
  OAI21_X1 U16574 ( .B1(n14787), .B2(n15521), .A(n14786), .ZN(n14807) );
  OAI22_X1 U16575 ( .A1(n15544), .A2(n14807), .B1(P3_REG1_REG_30__SCAN_IN), 
        .B2(n15547), .ZN(n14788) );
  INV_X1 U16576 ( .A(n14788), .ZN(P3_U3489) );
  OAI22_X1 U16577 ( .A1(n14791), .A2(n14790), .B1(n15521), .B2(n14789), .ZN(
        n14792) );
  NOR2_X1 U16578 ( .A1(n14793), .A2(n14792), .ZN(n14810) );
  INV_X1 U16579 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n14794) );
  AOI22_X1 U16580 ( .A1(n15547), .A2(n14810), .B1(n14794), .B2(n15544), .ZN(
        P3_U3473) );
  AOI211_X1 U16581 ( .C1(n14797), .C2(n15497), .A(n14796), .B(n14795), .ZN(
        n14812) );
  AOI22_X1 U16582 ( .A1(n15547), .A2(n14812), .B1(n14798), .B2(n15544), .ZN(
        P3_U3472) );
  AOI211_X1 U16583 ( .C1(n14801), .C2(n15497), .A(n14800), .B(n14799), .ZN(
        n14814) );
  AOI22_X1 U16584 ( .A1(n15547), .A2(n14814), .B1(n14802), .B2(n15544), .ZN(
        P3_U3471) );
  AOI211_X1 U16585 ( .C1(n15497), .C2(n14805), .A(n14804), .B(n14803), .ZN(
        n14816) );
  AOI22_X1 U16586 ( .A1(n15547), .A2(n14816), .B1(n14806), .B2(n15544), .ZN(
        P3_U3470) );
  OAI22_X1 U16587 ( .A1(n15526), .A2(n14807), .B1(P3_REG0_REG_30__SCAN_IN), 
        .B2(n15528), .ZN(n14808) );
  INV_X1 U16588 ( .A(n14808), .ZN(P3_U3457) );
  INV_X1 U16589 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n14809) );
  AOI22_X1 U16590 ( .A1(n15528), .A2(n14810), .B1(n14809), .B2(n15526), .ZN(
        P3_U3432) );
  INV_X1 U16591 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14811) );
  AOI22_X1 U16592 ( .A1(n15528), .A2(n14812), .B1(n14811), .B2(n15526), .ZN(
        P3_U3429) );
  INV_X1 U16593 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14813) );
  AOI22_X1 U16594 ( .A1(n15528), .A2(n14814), .B1(n14813), .B2(n15526), .ZN(
        P3_U3426) );
  AOI22_X1 U16595 ( .A1(n15528), .A2(n14816), .B1(n14815), .B2(n15526), .ZN(
        P3_U3423) );
  OAI21_X1 U16596 ( .B1(n14851), .B2(n14874), .A(n14852), .ZN(n14818) );
  OR2_X1 U16597 ( .A1(n14818), .A2(n14817), .ZN(n14872) );
  AOI21_X1 U16598 ( .B1(n14820), .B2(n14835), .A(n14819), .ZN(n14824) );
  INV_X1 U16599 ( .A(n14821), .ZN(n14822) );
  AOI21_X1 U16600 ( .B1(n14824), .B2(n14823), .A(n14822), .ZN(n14873) );
  INV_X1 U16601 ( .A(n14825), .ZN(n14829) );
  NOR2_X1 U16602 ( .A1(n14827), .A2(n14826), .ZN(n14828) );
  AOI21_X1 U16603 ( .B1(n14830), .B2(n14829), .A(n14828), .ZN(n14831) );
  OAI211_X1 U16604 ( .C1(n6843), .C2(n14872), .A(n14873), .B(n14831), .ZN(
        n14833) );
  INV_X1 U16605 ( .A(n14833), .ZN(n14837) );
  OAI21_X1 U16606 ( .B1(n6659), .B2(n14835), .A(n14834), .ZN(n14876) );
  AOI22_X1 U16607 ( .A1(n14876), .A2(n15288), .B1(P2_REG2_REG_15__SCAN_IN), 
        .B2(n15292), .ZN(n14836) );
  OAI21_X1 U16608 ( .B1(n15292), .B2(n14837), .A(n14836), .ZN(P2_U3250) );
  XNOR2_X1 U16609 ( .A(n14839), .B(n14838), .ZN(n14842) );
  AOI21_X1 U16610 ( .B1(n14842), .B2(n14841), .A(n14840), .ZN(n14879) );
  AOI222_X1 U16611 ( .A1(n14849), .A2(n14844), .B1(P2_REG2_REG_14__SCAN_IN), 
        .B2(n15292), .C1(n14843), .C2(n15279), .ZN(n14856) );
  INV_X1 U16612 ( .A(n14845), .ZN(n14846) );
  AOI21_X1 U16613 ( .B1(n14848), .B2(n14847), .A(n14846), .ZN(n14882) );
  INV_X1 U16614 ( .A(n14849), .ZN(n14878) );
  INV_X1 U16615 ( .A(n14851), .ZN(n14853) );
  OAI211_X1 U16616 ( .C1(n14878), .C2(n7324), .A(n14853), .B(n14852), .ZN(
        n14877) );
  INV_X1 U16617 ( .A(n14877), .ZN(n14854) );
  AOI22_X1 U16618 ( .A1(n14882), .A2(n15288), .B1(n14854), .B2(n15285), .ZN(
        n14855) );
  OAI211_X1 U16619 ( .C1(n15292), .C2(n14879), .A(n14856), .B(n14855), .ZN(
        P2_U3251) );
  INV_X1 U16620 ( .A(n14857), .ZN(n14862) );
  OAI21_X1 U16621 ( .B1(n14859), .B2(n15380), .A(n14858), .ZN(n14861) );
  AOI211_X1 U16622 ( .C1(n14862), .C2(n15377), .A(n14861), .B(n14860), .ZN(
        n14893) );
  AOI22_X1 U16623 ( .A1(n15401), .A2(n14893), .B1(n14863), .B2(n15399), .ZN(
        P2_U3516) );
  NAND3_X1 U16624 ( .A1(n14865), .A2(n14864), .A3(n15377), .ZN(n14867) );
  OAI211_X1 U16625 ( .C1(n14868), .C2(n15380), .A(n14867), .B(n14866), .ZN(
        n14870) );
  NOR2_X1 U16626 ( .A1(n14870), .A2(n14869), .ZN(n14895) );
  AOI22_X1 U16627 ( .A1(n15401), .A2(n14895), .B1(n14871), .B2(n15399), .ZN(
        P2_U3515) );
  OAI211_X1 U16628 ( .C1(n14874), .C2(n15380), .A(n14873), .B(n14872), .ZN(
        n14875) );
  AOI21_X1 U16629 ( .B1(n15377), .B2(n14876), .A(n14875), .ZN(n14897) );
  AOI22_X1 U16630 ( .A1(n15401), .A2(n14897), .B1(n10706), .B2(n15399), .ZN(
        P2_U3514) );
  OAI21_X1 U16631 ( .B1(n14878), .B2(n15380), .A(n14877), .ZN(n14881) );
  INV_X1 U16632 ( .A(n14879), .ZN(n14880) );
  AOI211_X1 U16633 ( .C1(n14882), .C2(n15377), .A(n14881), .B(n14880), .ZN(
        n14899) );
  AOI22_X1 U16634 ( .A1(n15401), .A2(n14899), .B1(n14883), .B2(n15399), .ZN(
        P2_U3513) );
  AND2_X1 U16635 ( .A1(n14884), .A2(n15377), .ZN(n14890) );
  NAND2_X1 U16636 ( .A1(n14885), .A2(n15368), .ZN(n14886) );
  NAND2_X1 U16637 ( .A1(n14887), .A2(n14886), .ZN(n14888) );
  NOR3_X1 U16638 ( .A1(n14890), .A2(n14889), .A3(n14888), .ZN(n14900) );
  INV_X1 U16639 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n14891) );
  AOI22_X1 U16640 ( .A1(n15401), .A2(n14900), .B1(n14891), .B2(n15399), .ZN(
        P2_U3512) );
  INV_X1 U16641 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n14892) );
  AOI22_X1 U16642 ( .A1(n15387), .A2(n14893), .B1(n14892), .B2(n15385), .ZN(
        P2_U3481) );
  INV_X1 U16643 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n14894) );
  AOI22_X1 U16644 ( .A1(n15387), .A2(n14895), .B1(n14894), .B2(n15385), .ZN(
        P2_U3478) );
  INV_X1 U16645 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n14896) );
  AOI22_X1 U16646 ( .A1(n15387), .A2(n14897), .B1(n14896), .B2(n15385), .ZN(
        P2_U3475) );
  INV_X1 U16647 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n14898) );
  AOI22_X1 U16648 ( .A1(n15387), .A2(n14899), .B1(n14898), .B2(n15385), .ZN(
        P2_U3472) );
  AOI22_X1 U16649 ( .A1(n15387), .A2(n14900), .B1(n8729), .B2(n15385), .ZN(
        P2_U3469) );
  OAI22_X1 U16650 ( .A1(n14901), .A2(n14925), .B1(n14926), .B2(n14912), .ZN(
        n14908) );
  OAI21_X1 U16651 ( .B1(n14904), .B2(n14903), .A(n14902), .ZN(n14906) );
  AOI21_X1 U16652 ( .B1(n14906), .B2(n14905), .A(n14932), .ZN(n14907) );
  AOI211_X1 U16653 ( .C1(n14909), .C2(n14937), .A(n14908), .B(n14907), .ZN(
        n14910) );
  NAND2_X1 U16654 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n15039)
         );
  OAI211_X1 U16655 ( .C1(n14941), .C2(n14911), .A(n14910), .B(n15039), .ZN(
        P1_U3215) );
  OAI22_X1 U16656 ( .A1(n14913), .A2(n14926), .B1(n14925), .B2(n14912), .ZN(
        n14920) );
  AOI21_X1 U16657 ( .B1(n13993), .B2(n14915), .A(n14914), .ZN(n14916) );
  INV_X1 U16658 ( .A(n14916), .ZN(n14918) );
  AOI21_X1 U16659 ( .B1(n14918), .B2(n14917), .A(n14932), .ZN(n14919) );
  AOI211_X1 U16660 ( .C1(n14921), .C2(n14937), .A(n14920), .B(n14919), .ZN(
        n14922) );
  NAND2_X1 U16661 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n15069)
         );
  OAI211_X1 U16662 ( .C1(n14941), .C2(n14923), .A(n14922), .B(n15069), .ZN(
        P1_U3226) );
  OAI22_X1 U16663 ( .A1(n14927), .A2(n14926), .B1(n14925), .B2(n14924), .ZN(
        n14936) );
  AOI21_X1 U16664 ( .B1(n14930), .B2(n14929), .A(n14928), .ZN(n14931) );
  INV_X1 U16665 ( .A(n14931), .ZN(n14934) );
  AOI21_X1 U16666 ( .B1(n14934), .B2(n14933), .A(n14932), .ZN(n14935) );
  AOI211_X1 U16667 ( .C1(n14938), .C2(n14937), .A(n14936), .B(n14935), .ZN(
        n14939) );
  NAND2_X1 U16668 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n15012)
         );
  OAI211_X1 U16669 ( .C1(n14941), .C2(n14940), .A(n14939), .B(n15012), .ZN(
        P1_U3236) );
  INV_X1 U16670 ( .A(n14942), .ZN(n14947) );
  OAI21_X1 U16671 ( .B1(n14944), .B2(n15187), .A(n14943), .ZN(n14946) );
  AOI211_X1 U16672 ( .C1(n14947), .C2(n15191), .A(n14946), .B(n14945), .ZN(
        n14974) );
  AOI22_X1 U16673 ( .A1(n15202), .A2(n14974), .B1(n14342), .B2(n15200), .ZN(
        P1_U3545) );
  INV_X1 U16674 ( .A(n14948), .ZN(n14953) );
  OAI211_X1 U16675 ( .C1(n14951), .C2(n15187), .A(n14950), .B(n14949), .ZN(
        n14952) );
  AOI21_X1 U16676 ( .B1(n14953), .B2(n15191), .A(n14952), .ZN(n14976) );
  AOI22_X1 U16677 ( .A1(n15202), .A2(n14976), .B1(n14334), .B2(n15200), .ZN(
        P1_U3544) );
  AOI21_X1 U16678 ( .B1(n14956), .B2(n14955), .A(n14954), .ZN(n14957) );
  OAI21_X1 U16679 ( .B1(n14958), .B2(n15161), .A(n14957), .ZN(n14962) );
  NOR3_X1 U16680 ( .A1(n14960), .A2(n14959), .A3(n15109), .ZN(n14961) );
  AOI211_X1 U16681 ( .C1(n15191), .C2(n14963), .A(n14962), .B(n14961), .ZN(
        n14978) );
  AOI22_X1 U16682 ( .A1(n15202), .A2(n14978), .B1(n15047), .B2(n15200), .ZN(
        P1_U3543) );
  AND3_X1 U16683 ( .A1(n14965), .A2(n15191), .A3(n14964), .ZN(n14970) );
  OAI211_X1 U16684 ( .C1(n14968), .C2(n15187), .A(n14967), .B(n14966), .ZN(
        n14969) );
  AOI211_X1 U16685 ( .C1(n14972), .C2(n11791), .A(n14970), .B(n14969), .ZN(
        n14980) );
  AOI22_X1 U16686 ( .A1(n15202), .A2(n14980), .B1(n14335), .B2(n15200), .ZN(
        P1_U3542) );
  INV_X1 U16687 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n14973) );
  AOI22_X1 U16688 ( .A1(n15194), .A2(n14974), .B1(n14973), .B2(n15192), .ZN(
        P1_U3510) );
  INV_X1 U16689 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n14975) );
  AOI22_X1 U16690 ( .A1(n15194), .A2(n14976), .B1(n14975), .B2(n15192), .ZN(
        P1_U3507) );
  INV_X1 U16691 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n14977) );
  AOI22_X1 U16692 ( .A1(n15194), .A2(n14978), .B1(n14977), .B2(n15192), .ZN(
        P1_U3504) );
  INV_X1 U16693 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14979) );
  AOI22_X1 U16694 ( .A1(n15194), .A2(n14980), .B1(n14979), .B2(n15192), .ZN(
        P1_U3501) );
  OAI21_X1 U16695 ( .B1(n14983), .B2(n14982), .A(n14981), .ZN(n14984) );
  XNOR2_X1 U16696 ( .A(n14984), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  OAI222_X1 U16697 ( .A1(n15251), .A2(n14988), .B1(n15251), .B2(n14987), .C1(
        n14986), .C2(n14985), .ZN(SUB_1596_U68) );
  OAI21_X1 U16698 ( .B1(n14991), .B2(n14990), .A(n14989), .ZN(SUB_1596_U67) );
  OAI21_X1 U16699 ( .B1(n14994), .B2(n14993), .A(n14992), .ZN(SUB_1596_U66) );
  OAI21_X1 U16700 ( .B1(n14997), .B2(n14996), .A(n14995), .ZN(SUB_1596_U65) );
  AOI21_X1 U16701 ( .B1(n15000), .B2(n14999), .A(n14998), .ZN(n15001) );
  XOR2_X1 U16702 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n15001), .Z(SUB_1596_U64)
         );
  INV_X1 U16703 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n15014) );
  OAI21_X1 U16704 ( .B1(n15004), .B2(n15003), .A(n15002), .ZN(n15011) );
  NOR2_X1 U16705 ( .A1(n15100), .A2(n15005), .ZN(n15010) );
  AOI211_X1 U16706 ( .C1(n15008), .C2(n15007), .A(n15061), .B(n15006), .ZN(
        n15009) );
  AOI211_X1 U16707 ( .C1(n15091), .C2(n15011), .A(n15010), .B(n15009), .ZN(
        n15013) );
  OAI211_X1 U16708 ( .C1(n15014), .C2(n15104), .A(n15013), .B(n15012), .ZN(
        P1_U3254) );
  AOI211_X1 U16709 ( .C1(n15017), .C2(n15016), .A(n15015), .B(n15061), .ZN(
        n15022) );
  AOI211_X1 U16710 ( .C1(n15020), .C2(n15019), .A(n15018), .B(n15057), .ZN(
        n15021) );
  AOI211_X1 U16711 ( .C1(n15068), .C2(n15023), .A(n15022), .B(n15021), .ZN(
        n15025) );
  OAI211_X1 U16712 ( .C1(n15026), .C2(n15104), .A(n15025), .B(n15024), .ZN(
        P1_U3256) );
  INV_X1 U16713 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n15041) );
  AOI21_X1 U16714 ( .B1(n15029), .B2(n15028), .A(n15027), .ZN(n15030) );
  NAND2_X1 U16715 ( .A1(n15096), .A2(n15030), .ZN(n15036) );
  OAI21_X1 U16716 ( .B1(n15033), .B2(n15032), .A(n15031), .ZN(n15034) );
  NAND2_X1 U16717 ( .A1(n15091), .A2(n15034), .ZN(n15035) );
  OAI211_X1 U16718 ( .C1(n15100), .C2(n15037), .A(n15036), .B(n15035), .ZN(
        n15038) );
  INV_X1 U16719 ( .A(n15038), .ZN(n15040) );
  OAI211_X1 U16720 ( .C1(n15041), .C2(n15104), .A(n15040), .B(n15039), .ZN(
        P1_U3257) );
  OAI21_X1 U16721 ( .B1(n15044), .B2(n15043), .A(n15042), .ZN(n15045) );
  NAND2_X1 U16722 ( .A1(n15096), .A2(n15045), .ZN(n15051) );
  OAI21_X1 U16723 ( .B1(n15048), .B2(n15047), .A(n15046), .ZN(n15049) );
  NAND2_X1 U16724 ( .A1(n15091), .A2(n15049), .ZN(n15050) );
  OAI211_X1 U16725 ( .C1(n15100), .C2(n15052), .A(n15051), .B(n15050), .ZN(
        n15053) );
  INV_X1 U16726 ( .A(n15053), .ZN(n15055) );
  OAI211_X1 U16727 ( .C1(n15056), .C2(n15104), .A(n15055), .B(n15054), .ZN(
        P1_U3258) );
  AOI211_X1 U16728 ( .C1(n15060), .C2(n15059), .A(n15058), .B(n15057), .ZN(
        n15066) );
  AOI211_X1 U16729 ( .C1(n15064), .C2(n15063), .A(n15062), .B(n15061), .ZN(
        n15065) );
  AOI211_X1 U16730 ( .C1(n15068), .C2(n15067), .A(n15066), .B(n15065), .ZN(
        n15070) );
  OAI211_X1 U16731 ( .C1(n15071), .C2(n15104), .A(n15070), .B(n15069), .ZN(
        P1_U3259) );
  AOI21_X1 U16732 ( .B1(n15074), .B2(n15073), .A(n15072), .ZN(n15075) );
  NAND2_X1 U16733 ( .A1(n15096), .A2(n15075), .ZN(n15081) );
  AOI21_X1 U16734 ( .B1(n15078), .B2(n15077), .A(n15076), .ZN(n15079) );
  NAND2_X1 U16735 ( .A1(n15091), .A2(n15079), .ZN(n15080) );
  OAI211_X1 U16736 ( .C1(n15100), .C2(n15082), .A(n15081), .B(n15080), .ZN(
        n15083) );
  INV_X1 U16737 ( .A(n15083), .ZN(n15085) );
  OAI211_X1 U16738 ( .C1(n15086), .C2(n15104), .A(n15085), .B(n15084), .ZN(
        P1_U3260) );
  INV_X1 U16739 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n15105) );
  AOI21_X1 U16740 ( .B1(n15089), .B2(n15088), .A(n15087), .ZN(n15090) );
  NAND2_X1 U16741 ( .A1(n15091), .A2(n15090), .ZN(n15098) );
  AOI21_X1 U16742 ( .B1(n15094), .B2(n15093), .A(n15092), .ZN(n15095) );
  NAND2_X1 U16743 ( .A1(n15096), .A2(n15095), .ZN(n15097) );
  OAI211_X1 U16744 ( .C1(n15100), .C2(n15099), .A(n15098), .B(n15097), .ZN(
        n15101) );
  INV_X1 U16745 ( .A(n15101), .ZN(n15103) );
  OAI211_X1 U16746 ( .C1(n15105), .C2(n15104), .A(n15103), .B(n15102), .ZN(
        P1_U3261) );
  XNOR2_X1 U16747 ( .A(n15106), .B(n15108), .ZN(n15172) );
  XNOR2_X1 U16748 ( .A(n15108), .B(n15107), .ZN(n15110) );
  NOR2_X1 U16749 ( .A1(n15110), .A2(n15109), .ZN(n15111) );
  AOI211_X1 U16750 ( .C1(n15172), .C2(n15183), .A(n15112), .B(n15111), .ZN(
        n15169) );
  AOI22_X1 U16751 ( .A1(n15129), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n15114), .ZN(n15115) );
  OAI21_X1 U16752 ( .B1(n15116), .B2(n6840), .A(n15115), .ZN(n15117) );
  INV_X1 U16753 ( .A(n15117), .ZN(n15128) );
  NAND2_X1 U16754 ( .A1(n15119), .A2(n15118), .ZN(n15121) );
  NAND2_X1 U16755 ( .A1(n15121), .A2(n15120), .ZN(n15123) );
  OR2_X1 U16756 ( .A1(n15123), .A2(n15122), .ZN(n15168) );
  INV_X1 U16757 ( .A(n15168), .ZN(n15124) );
  AOI22_X1 U16758 ( .A1(n15126), .A2(n15172), .B1(n15125), .B2(n15124), .ZN(
        n15127) );
  OAI211_X1 U16759 ( .C1(n15129), .C2(n15169), .A(n15128), .B(n15127), .ZN(
        P1_U3291) );
  INV_X1 U16760 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n15130) );
  NOR2_X1 U16761 ( .A1(n15160), .A2(n15130), .ZN(P1_U3294) );
  NOR2_X1 U16762 ( .A1(n15160), .A2(n15131), .ZN(P1_U3295) );
  NOR2_X1 U16763 ( .A1(n15160), .A2(n15132), .ZN(P1_U3296) );
  INV_X1 U16764 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n15133) );
  NOR2_X1 U16765 ( .A1(n15160), .A2(n15133), .ZN(P1_U3297) );
  NOR2_X1 U16766 ( .A1(n15160), .A2(n15134), .ZN(P1_U3298) );
  INV_X1 U16767 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n15135) );
  NOR2_X1 U16768 ( .A1(n15160), .A2(n15135), .ZN(P1_U3299) );
  INV_X1 U16769 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n15136) );
  NOR2_X1 U16770 ( .A1(n15160), .A2(n15136), .ZN(P1_U3300) );
  INV_X1 U16771 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n15137) );
  NOR2_X1 U16772 ( .A1(n15160), .A2(n15137), .ZN(P1_U3301) );
  INV_X1 U16773 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n15138) );
  NOR2_X1 U16774 ( .A1(n15160), .A2(n15138), .ZN(P1_U3302) );
  INV_X1 U16775 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n15139) );
  NOR2_X1 U16776 ( .A1(n15160), .A2(n15139), .ZN(P1_U3303) );
  INV_X1 U16777 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n15140) );
  NOR2_X1 U16778 ( .A1(n15160), .A2(n15140), .ZN(P1_U3304) );
  NOR2_X1 U16779 ( .A1(n15160), .A2(n15141), .ZN(P1_U3305) );
  INV_X1 U16780 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n15142) );
  NOR2_X1 U16781 ( .A1(n15160), .A2(n15142), .ZN(P1_U3306) );
  INV_X1 U16782 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n15143) );
  NOR2_X1 U16783 ( .A1(n15160), .A2(n15143), .ZN(P1_U3307) );
  INV_X1 U16784 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n15144) );
  NOR2_X1 U16785 ( .A1(n15160), .A2(n15144), .ZN(P1_U3308) );
  INV_X1 U16786 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n15145) );
  NOR2_X1 U16787 ( .A1(n15160), .A2(n15145), .ZN(P1_U3309) );
  INV_X1 U16788 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n15146) );
  NOR2_X1 U16789 ( .A1(n15160), .A2(n15146), .ZN(P1_U3310) );
  INV_X1 U16790 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n15147) );
  NOR2_X1 U16791 ( .A1(n15160), .A2(n15147), .ZN(P1_U3311) );
  NOR2_X1 U16792 ( .A1(n15160), .A2(n15148), .ZN(P1_U3312) );
  INV_X1 U16793 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n15149) );
  NOR2_X1 U16794 ( .A1(n15160), .A2(n15149), .ZN(P1_U3313) );
  INV_X1 U16795 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n15150) );
  NOR2_X1 U16796 ( .A1(n15160), .A2(n15150), .ZN(P1_U3314) );
  INV_X1 U16797 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n15151) );
  NOR2_X1 U16798 ( .A1(n15160), .A2(n15151), .ZN(P1_U3315) );
  INV_X1 U16799 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n15152) );
  NOR2_X1 U16800 ( .A1(n15160), .A2(n15152), .ZN(P1_U3316) );
  INV_X1 U16801 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n15153) );
  NOR2_X1 U16802 ( .A1(n15160), .A2(n15153), .ZN(P1_U3317) );
  INV_X1 U16803 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n15154) );
  NOR2_X1 U16804 ( .A1(n15160), .A2(n15154), .ZN(P1_U3318) );
  INV_X1 U16805 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n15155) );
  NOR2_X1 U16806 ( .A1(n15160), .A2(n15155), .ZN(P1_U3319) );
  INV_X1 U16807 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n15156) );
  NOR2_X1 U16808 ( .A1(n15160), .A2(n15156), .ZN(P1_U3320) );
  NOR2_X1 U16809 ( .A1(n15160), .A2(n15157), .ZN(P1_U3321) );
  INV_X1 U16810 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n15158) );
  NOR2_X1 U16811 ( .A1(n15160), .A2(n15158), .ZN(P1_U3322) );
  INV_X1 U16812 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n15159) );
  NOR2_X1 U16813 ( .A1(n15160), .A2(n15159), .ZN(P1_U3323) );
  OAI22_X1 U16814 ( .A1(n15162), .A2(n15161), .B1(n9972), .B2(n15187), .ZN(
        n15165) );
  INV_X1 U16815 ( .A(n15163), .ZN(n15164) );
  AOI211_X1 U16816 ( .C1(n15166), .C2(n15191), .A(n15165), .B(n15164), .ZN(
        n15196) );
  INV_X1 U16817 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n15167) );
  AOI22_X1 U16818 ( .A1(n15194), .A2(n15196), .B1(n15167), .B2(n15192), .ZN(
        P1_U3462) );
  OAI21_X1 U16819 ( .B1(n6840), .B2(n15187), .A(n15168), .ZN(n15171) );
  INV_X1 U16820 ( .A(n15169), .ZN(n15170) );
  AOI211_X1 U16821 ( .C1(n15173), .C2(n15172), .A(n15171), .B(n15170), .ZN(
        n15198) );
  INV_X1 U16822 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n15174) );
  AOI22_X1 U16823 ( .A1(n15194), .A2(n15198), .B1(n15174), .B2(n15192), .ZN(
        P1_U3465) );
  NOR2_X1 U16824 ( .A1(n15176), .A2(n15175), .ZN(n15181) );
  OAI211_X1 U16825 ( .C1(n15179), .C2(n15187), .A(n15178), .B(n15177), .ZN(
        n15180) );
  AOI211_X1 U16826 ( .C1(n15183), .C2(n15182), .A(n15181), .B(n15180), .ZN(
        n15199) );
  INV_X1 U16827 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n15184) );
  AOI22_X1 U16828 ( .A1(n15194), .A2(n15199), .B1(n15184), .B2(n15192), .ZN(
        P1_U3468) );
  OAI211_X1 U16829 ( .C1(n15188), .C2(n15187), .A(n15186), .B(n15185), .ZN(
        n15189) );
  AOI21_X1 U16830 ( .B1(n15191), .B2(n15190), .A(n15189), .ZN(n15201) );
  INV_X1 U16831 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n15193) );
  AOI22_X1 U16832 ( .A1(n15194), .A2(n15201), .B1(n15193), .B2(n15192), .ZN(
        P1_U3489) );
  AOI22_X1 U16833 ( .A1(n15202), .A2(n15196), .B1(n15195), .B2(n15200), .ZN(
        P1_U3529) );
  AOI22_X1 U16834 ( .A1(n15202), .A2(n15198), .B1(n15197), .B2(n15200), .ZN(
        P1_U3530) );
  AOI22_X1 U16835 ( .A1(n15202), .A2(n15199), .B1(n9304), .B2(n15200), .ZN(
        P1_U3531) );
  AOI22_X1 U16836 ( .A1(n15202), .A2(n15201), .B1(n9906), .B2(n15200), .ZN(
        P1_U3538) );
  NOR2_X1 U16837 ( .A1(n15270), .A2(P2_U3947), .ZN(P2_U3087) );
  OAI21_X1 U16838 ( .B1(n15204), .B2(n15203), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15205) );
  OAI21_X1 U16839 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n15205), .ZN(n15215) );
  OAI211_X1 U16840 ( .C1(n15208), .C2(n15207), .A(n15271), .B(n15206), .ZN(
        n15214) );
  OAI211_X1 U16841 ( .C1(n15211), .C2(n15210), .A(n15264), .B(n15209), .ZN(
        n15213) );
  NAND2_X1 U16842 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n15270), .ZN(n15212) );
  NAND4_X1 U16843 ( .A1(n15215), .A2(n15214), .A3(n15213), .A4(n15212), .ZN(
        P2_U3215) );
  NAND2_X1 U16844 ( .A1(n15270), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n15216) );
  OAI211_X1 U16845 ( .C1(n15278), .C2(n15218), .A(n15217), .B(n15216), .ZN(
        n15219) );
  INV_X1 U16846 ( .A(n15219), .ZN(n15232) );
  AOI21_X1 U16847 ( .B1(n15222), .B2(n15221), .A(n15220), .ZN(n15224) );
  NAND2_X1 U16848 ( .A1(n15224), .A2(n15223), .ZN(n15231) );
  AOI21_X1 U16849 ( .B1(n15227), .B2(n15226), .A(n15225), .ZN(n15229) );
  NAND2_X1 U16850 ( .A1(n15229), .A2(n15228), .ZN(n15230) );
  NAND3_X1 U16851 ( .A1(n15232), .A2(n15231), .A3(n15230), .ZN(P2_U3224) );
  INV_X1 U16852 ( .A(n15233), .ZN(n15235) );
  NAND3_X1 U16853 ( .A1(n15236), .A2(n15235), .A3(n15234), .ZN(n15237) );
  NAND2_X1 U16854 ( .A1(n15238), .A2(n15237), .ZN(n15239) );
  NAND2_X1 U16855 ( .A1(n15239), .A2(n15271), .ZN(n15245) );
  OAI21_X1 U16856 ( .B1(n15242), .B2(n15241), .A(n15240), .ZN(n15243) );
  NAND2_X1 U16857 ( .A1(n15243), .A2(n15264), .ZN(n15244) );
  OAI211_X1 U16858 ( .C1(n15278), .C2(n15246), .A(n15245), .B(n15244), .ZN(
        n15247) );
  INV_X1 U16859 ( .A(n15247), .ZN(n15249) );
  OAI211_X1 U16860 ( .C1(n15251), .C2(n15250), .A(n15249), .B(n15248), .ZN(
        P2_U3226) );
  AOI22_X1 U16861 ( .A1(n15270), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n15262) );
  NAND2_X1 U16862 ( .A1(n15254), .A2(n15253), .ZN(n15261) );
  OAI211_X1 U16863 ( .C1(n15256), .C2(P2_REG2_REG_15__SCAN_IN), .A(n15271), 
        .B(n15255), .ZN(n15260) );
  XNOR2_X1 U16864 ( .A(n15257), .B(P2_REG1_REG_15__SCAN_IN), .ZN(n15258) );
  NAND2_X1 U16865 ( .A1(n15258), .A2(n15264), .ZN(n15259) );
  NAND4_X1 U16866 ( .A1(n15262), .A2(n15261), .A3(n15260), .A4(n15259), .ZN(
        P2_U3229) );
  OAI211_X1 U16867 ( .C1(n15266), .C2(n15265), .A(n15264), .B(n15263), .ZN(
        n15267) );
  NAND2_X1 U16868 ( .A1(n15268), .A2(n15267), .ZN(n15269) );
  AOI21_X1 U16869 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(n15270), .A(n15269), 
        .ZN(n15276) );
  OAI211_X1 U16870 ( .C1(n15274), .C2(n15273), .A(n15272), .B(n15271), .ZN(
        n15275) );
  OAI211_X1 U16871 ( .C1(n15278), .C2(n15277), .A(n15276), .B(n15275), .ZN(
        P2_U3231) );
  AOI22_X1 U16872 ( .A1(n15292), .A2(P2_REG2_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(n15279), .ZN(n15280) );
  OAI21_X1 U16873 ( .B1(n15282), .B2(n15281), .A(n15280), .ZN(n15283) );
  INV_X1 U16874 ( .A(n15283), .ZN(n15290) );
  INV_X1 U16875 ( .A(n15284), .ZN(n15286) );
  AOI22_X1 U16876 ( .A1(n15288), .A2(n15287), .B1(n15286), .B2(n15285), .ZN(
        n15289) );
  OAI211_X1 U16877 ( .C1(n15292), .C2(n15291), .A(n15290), .B(n15289), .ZN(
        P2_U3263) );
  NOR2_X1 U16878 ( .A1(n15293), .A2(n15302), .ZN(n15301) );
  AND2_X1 U16879 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15298), .ZN(P2_U3266) );
  AND2_X1 U16880 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15298), .ZN(P2_U3267) );
  AND2_X1 U16881 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15298), .ZN(P2_U3268) );
  AND2_X1 U16882 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15298), .ZN(P2_U3269) );
  AND2_X1 U16883 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15298), .ZN(P2_U3270) );
  NOR2_X1 U16884 ( .A1(n15301), .A2(n15294), .ZN(P2_U3271) );
  AND2_X1 U16885 ( .A1(n15298), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3272) );
  AND2_X1 U16886 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15298), .ZN(P2_U3273) );
  AND2_X1 U16887 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15298), .ZN(P2_U3274) );
  AND2_X1 U16888 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15298), .ZN(P2_U3275) );
  NOR2_X1 U16889 ( .A1(n15301), .A2(n15295), .ZN(P2_U3276) );
  AND2_X1 U16890 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15298), .ZN(P2_U3277) );
  AND2_X1 U16891 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15298), .ZN(P2_U3278) );
  NOR2_X1 U16892 ( .A1(n15301), .A2(n15296), .ZN(P2_U3279) );
  AND2_X1 U16893 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15298), .ZN(P2_U3280) );
  AND2_X1 U16894 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15298), .ZN(P2_U3281) );
  AND2_X1 U16895 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15298), .ZN(P2_U3282) );
  AND2_X1 U16896 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15298), .ZN(P2_U3283) );
  AND2_X1 U16897 ( .A1(n15298), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3284) );
  AND2_X1 U16898 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15298), .ZN(P2_U3285) );
  AND2_X1 U16899 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15298), .ZN(P2_U3286) );
  AND2_X1 U16900 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15298), .ZN(P2_U3287) );
  AND2_X1 U16901 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15298), .ZN(P2_U3288) );
  AND2_X1 U16902 ( .A1(n15298), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3289) );
  AND2_X1 U16903 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15298), .ZN(P2_U3290) );
  NOR2_X1 U16904 ( .A1(n15301), .A2(n15297), .ZN(P2_U3291) );
  AND2_X1 U16905 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15298), .ZN(P2_U3292) );
  AND2_X1 U16906 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15298), .ZN(P2_U3293) );
  AND2_X1 U16907 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15298), .ZN(P2_U3294) );
  AND2_X1 U16908 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15298), .ZN(P2_U3295) );
  AOI22_X1 U16909 ( .A1(n15301), .A2(n15300), .B1(n15299), .B2(n15298), .ZN(
        P2_U3416) );
  AOI22_X1 U16910 ( .A1(n15305), .A2(n15304), .B1(n15303), .B2(n15302), .ZN(
        P2_U3417) );
  OAI22_X1 U16911 ( .A1(n15308), .A2(n15372), .B1(n15307), .B2(n15306), .ZN(
        n15309) );
  NOR2_X1 U16912 ( .A1(n15310), .A2(n15309), .ZN(n15389) );
  INV_X1 U16913 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n15311) );
  AOI22_X1 U16914 ( .A1(n15387), .A2(n15389), .B1(n15311), .B2(n15385), .ZN(
        P2_U3430) );
  INV_X1 U16915 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n15312) );
  AOI22_X1 U16916 ( .A1(n15387), .A2(n15313), .B1(n15312), .B2(n15385), .ZN(
        P2_U3433) );
  INV_X1 U16917 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n15314) );
  AOI22_X1 U16918 ( .A1(n15387), .A2(n15315), .B1(n15314), .B2(n15385), .ZN(
        P2_U3436) );
  NOR2_X1 U16919 ( .A1(n15316), .A2(n15350), .ZN(n15321) );
  OAI21_X1 U16920 ( .B1(n6842), .B2(n15380), .A(n15317), .ZN(n15318) );
  NOR4_X1 U16921 ( .A1(n15321), .A2(n15320), .A3(n15319), .A4(n15318), .ZN(
        n15390) );
  INV_X1 U16922 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n15322) );
  AOI22_X1 U16923 ( .A1(n15387), .A2(n15390), .B1(n15322), .B2(n15385), .ZN(
        P2_U3439) );
  AOI21_X1 U16924 ( .B1(n15368), .B2(n15324), .A(n15323), .ZN(n15326) );
  OAI211_X1 U16925 ( .C1(n15372), .C2(n15327), .A(n15326), .B(n15325), .ZN(
        n15328) );
  INV_X1 U16926 ( .A(n15328), .ZN(n15391) );
  INV_X1 U16927 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n15329) );
  AOI22_X1 U16928 ( .A1(n15387), .A2(n15391), .B1(n15329), .B2(n15385), .ZN(
        P2_U3442) );
  INV_X1 U16929 ( .A(n15330), .ZN(n15332) );
  OAI211_X1 U16930 ( .C1(n15333), .C2(n15380), .A(n15332), .B(n15331), .ZN(
        n15336) );
  AOI21_X1 U16931 ( .B1(n15372), .B2(n15342), .A(n15334), .ZN(n15335) );
  NOR2_X1 U16932 ( .A1(n15336), .A2(n15335), .ZN(n15392) );
  INV_X1 U16933 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n15337) );
  AOI22_X1 U16934 ( .A1(n15387), .A2(n15392), .B1(n15337), .B2(n15385), .ZN(
        P2_U3445) );
  INV_X1 U16935 ( .A(n15338), .ZN(n15340) );
  OAI211_X1 U16936 ( .C1(n7314), .C2(n15380), .A(n15340), .B(n15339), .ZN(
        n15344) );
  AOI21_X1 U16937 ( .B1(n15372), .B2(n15342), .A(n15341), .ZN(n15343) );
  NOR2_X1 U16938 ( .A1(n15344), .A2(n15343), .ZN(n15393) );
  INV_X1 U16939 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n15345) );
  AOI22_X1 U16940 ( .A1(n15387), .A2(n15393), .B1(n15345), .B2(n15385), .ZN(
        P2_U3448) );
  AOI21_X1 U16941 ( .B1(n15368), .B2(n15347), .A(n15346), .ZN(n15349) );
  OAI211_X1 U16942 ( .C1(n15351), .C2(n15350), .A(n15349), .B(n15348), .ZN(
        n15352) );
  INV_X1 U16943 ( .A(n15352), .ZN(n15394) );
  INV_X1 U16944 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n15353) );
  AOI22_X1 U16945 ( .A1(n15387), .A2(n15394), .B1(n15353), .B2(n15385), .ZN(
        P2_U3451) );
  OAI21_X1 U16946 ( .B1(n15355), .B2(n15380), .A(n15354), .ZN(n15358) );
  INV_X1 U16947 ( .A(n15356), .ZN(n15357) );
  AOI211_X1 U16948 ( .C1(n9570), .C2(n15359), .A(n15358), .B(n15357), .ZN(
        n15395) );
  INV_X1 U16949 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n15360) );
  AOI22_X1 U16950 ( .A1(n15387), .A2(n15395), .B1(n15360), .B2(n15385), .ZN(
        P2_U3454) );
  NAND2_X1 U16951 ( .A1(n15361), .A2(n15368), .ZN(n15362) );
  OAI211_X1 U16952 ( .C1(n15364), .C2(n15372), .A(n15363), .B(n15362), .ZN(
        n15365) );
  NOR2_X1 U16953 ( .A1(n15366), .A2(n15365), .ZN(n15396) );
  INV_X1 U16954 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n15367) );
  AOI22_X1 U16955 ( .A1(n15387), .A2(n15396), .B1(n15367), .B2(n15385), .ZN(
        P2_U3457) );
  NAND2_X1 U16956 ( .A1(n15369), .A2(n15368), .ZN(n15370) );
  OAI211_X1 U16957 ( .C1(n15373), .C2(n15372), .A(n15371), .B(n15370), .ZN(
        n15374) );
  NOR2_X1 U16958 ( .A1(n15375), .A2(n15374), .ZN(n15398) );
  AOI22_X1 U16959 ( .A1(n15387), .A2(n15398), .B1(n15376), .B2(n15385), .ZN(
        P2_U3460) );
  AND2_X1 U16960 ( .A1(n15378), .A2(n15377), .ZN(n15384) );
  OAI21_X1 U16961 ( .B1(n15381), .B2(n15380), .A(n15379), .ZN(n15382) );
  NOR3_X1 U16962 ( .A1(n15384), .A2(n15383), .A3(n15382), .ZN(n15400) );
  INV_X1 U16963 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n15386) );
  AOI22_X1 U16964 ( .A1(n15387), .A2(n15400), .B1(n15386), .B2(n15385), .ZN(
        P2_U3463) );
  INV_X1 U16965 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n15388) );
  AOI22_X1 U16966 ( .A1(n15401), .A2(n15389), .B1(n15388), .B2(n15399), .ZN(
        P2_U3499) );
  AOI22_X1 U16967 ( .A1(n15401), .A2(n15390), .B1(n9397), .B2(n15399), .ZN(
        P2_U3502) );
  AOI22_X1 U16968 ( .A1(n15401), .A2(n15391), .B1(n9426), .B2(n15399), .ZN(
        P2_U3503) );
  AOI22_X1 U16969 ( .A1(n15401), .A2(n15392), .B1(n9427), .B2(n15399), .ZN(
        P2_U3504) );
  AOI22_X1 U16970 ( .A1(n15401), .A2(n15393), .B1(n9522), .B2(n15399), .ZN(
        P2_U3505) );
  AOI22_X1 U16971 ( .A1(n15401), .A2(n15394), .B1(n9523), .B2(n15399), .ZN(
        P2_U3506) );
  AOI22_X1 U16972 ( .A1(n15401), .A2(n15395), .B1(n9527), .B2(n15399), .ZN(
        P2_U3507) );
  AOI22_X1 U16973 ( .A1(n15401), .A2(n15396), .B1(n9530), .B2(n15399), .ZN(
        P2_U3508) );
  AOI22_X1 U16974 ( .A1(n15401), .A2(n15398), .B1(n15397), .B2(n15399), .ZN(
        P2_U3509) );
  AOI22_X1 U16975 ( .A1(n15401), .A2(n15400), .B1(n9534), .B2(n15399), .ZN(
        P2_U3510) );
  NOR2_X1 U16976 ( .A1(P3_U3897), .A2(n15405), .ZN(P3_U3150) );
  AOI22_X1 U16977 ( .A1(n15404), .A2(n15403), .B1(n7353), .B2(n15402), .ZN(
        n15413) );
  AOI22_X1 U16978 ( .A1(P3_ADDR_REG_0__SCAN_IN), .A2(n15405), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n15412) );
  NAND3_X1 U16979 ( .A1(n15438), .A2(n15425), .A3(n15434), .ZN(n15408) );
  INV_X1 U16980 ( .A(n15406), .ZN(n15407) );
  AOI22_X1 U16981 ( .A1(n15430), .A2(P3_IR_REG_0__SCAN_IN), .B1(n15408), .B2(
        n15407), .ZN(n15411) );
  OR3_X1 U16982 ( .A1(n15434), .A2(P3_IR_REG_0__SCAN_IN), .A3(n15409), .ZN(
        n15410) );
  NAND4_X1 U16983 ( .A1(n15413), .A2(n15412), .A3(n15411), .A4(n15410), .ZN(
        P3_U3182) );
  AOI21_X1 U16984 ( .B1(n15416), .B2(n15415), .A(n15414), .ZN(n15439) );
  INV_X1 U16985 ( .A(n15417), .ZN(n15429) );
  INV_X1 U16986 ( .A(n15418), .ZN(n15419) );
  OAI21_X1 U16987 ( .B1(n15421), .B2(n15420), .A(n15419), .ZN(n15428) );
  AOI21_X1 U16988 ( .B1(n15424), .B2(n15423), .A(n15422), .ZN(n15426) );
  NOR2_X1 U16989 ( .A1(n15426), .A2(n15425), .ZN(n15427) );
  AOI211_X1 U16990 ( .C1(n15430), .C2(n15429), .A(n15428), .B(n15427), .ZN(
        n15437) );
  AOI21_X1 U16991 ( .B1(n15433), .B2(n15432), .A(n15431), .ZN(n15435) );
  OR2_X1 U16992 ( .A1(n15435), .A2(n15434), .ZN(n15436) );
  OAI211_X1 U16993 ( .C1(n15439), .C2(n15438), .A(n15437), .B(n15436), .ZN(
        P3_U3192) );
  OAI21_X1 U16994 ( .B1(n15441), .B2(n15446), .A(n15440), .ZN(n15485) );
  NOR2_X1 U16995 ( .A1(n15442), .A2(n15521), .ZN(n15484) );
  INV_X1 U16996 ( .A(n15484), .ZN(n15445) );
  OAI22_X1 U16997 ( .A1(n15445), .A2(n15444), .B1(n10022), .B2(n15443), .ZN(
        n15457) );
  XNOR2_X1 U16998 ( .A(n15447), .B(n15446), .ZN(n15455) );
  OAI22_X1 U16999 ( .A1(n15451), .A2(n15450), .B1(n15449), .B2(n15448), .ZN(
        n15452) );
  AOI21_X1 U17000 ( .B1(n15485), .B2(n15453), .A(n15452), .ZN(n15454) );
  OAI21_X1 U17001 ( .B1(n15456), .B2(n15455), .A(n15454), .ZN(n15483) );
  AOI211_X1 U17002 ( .C1(n15458), .C2(n15485), .A(n15457), .B(n15483), .ZN(
        n15459) );
  AOI22_X1 U17003 ( .A1(n12871), .A2(n10148), .B1(n15459), .B2(n15477), .ZN(
        P3_U3231) );
  NOR2_X1 U17004 ( .A1(n7796), .A2(n15521), .ZN(n15480) );
  XNOR2_X1 U17005 ( .A(n15460), .B(n10025), .ZN(n15472) );
  AOI22_X1 U17006 ( .A1(n15464), .A2(n15463), .B1(n15462), .B2(n15461), .ZN(
        n15469) );
  XNOR2_X1 U17007 ( .A(n10025), .B(n15465), .ZN(n15467) );
  NAND2_X1 U17008 ( .A1(n15467), .A2(n15466), .ZN(n15468) );
  OAI211_X1 U17009 ( .C1(n15472), .C2(n15470), .A(n15469), .B(n15468), .ZN(
        n15479) );
  AOI21_X1 U17010 ( .B1(n15480), .B2(n15471), .A(n15479), .ZN(n15478) );
  INV_X1 U17011 ( .A(n15472), .ZN(n15481) );
  AOI22_X1 U17012 ( .A1(n15481), .A2(n15474), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15473), .ZN(n15475) );
  OAI221_X1 U17013 ( .B1(n12871), .B2(n15478), .C1(n15477), .C2(n15476), .A(
        n15475), .ZN(P3_U3232) );
  AOI211_X1 U17014 ( .C1(n15517), .C2(n15481), .A(n15480), .B(n15479), .ZN(
        n15530) );
  INV_X1 U17015 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15482) );
  AOI22_X1 U17016 ( .A1(n15528), .A2(n15530), .B1(n15482), .B2(n15526), .ZN(
        P3_U3393) );
  AOI211_X1 U17017 ( .C1(n15517), .C2(n15485), .A(n15484), .B(n15483), .ZN(
        n15531) );
  INV_X1 U17018 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15486) );
  AOI22_X1 U17019 ( .A1(n15528), .A2(n15531), .B1(n15486), .B2(n15526), .ZN(
        P3_U3396) );
  AOI22_X1 U17020 ( .A1(n15489), .A2(n15517), .B1(n15488), .B2(n15487), .ZN(
        n15490) );
  AND2_X1 U17021 ( .A1(n15491), .A2(n15490), .ZN(n15533) );
  INV_X1 U17022 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15492) );
  AOI22_X1 U17023 ( .A1(n15528), .A2(n15533), .B1(n15492), .B2(n15526), .ZN(
        P3_U3399) );
  INV_X1 U17024 ( .A(n15493), .ZN(n15498) );
  INV_X1 U17025 ( .A(n15494), .ZN(n15495) );
  AOI211_X1 U17026 ( .C1(n15498), .C2(n15497), .A(n15496), .B(n15495), .ZN(
        n15535) );
  INV_X1 U17027 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15499) );
  AOI22_X1 U17028 ( .A1(n15528), .A2(n15535), .B1(n15499), .B2(n15526), .ZN(
        P3_U3402) );
  INV_X1 U17029 ( .A(n15500), .ZN(n15503) );
  AOI211_X1 U17030 ( .C1(n15503), .C2(n15517), .A(n15502), .B(n15501), .ZN(
        n15537) );
  INV_X1 U17031 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15504) );
  AOI22_X1 U17032 ( .A1(n15528), .A2(n15537), .B1(n15504), .B2(n15526), .ZN(
        P3_U3405) );
  AOI211_X1 U17033 ( .C1(n15517), .C2(n15507), .A(n15506), .B(n15505), .ZN(
        n15539) );
  INV_X1 U17034 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15508) );
  AOI22_X1 U17035 ( .A1(n15528), .A2(n15539), .B1(n15508), .B2(n15526), .ZN(
        P3_U3408) );
  OAI22_X1 U17036 ( .A1(n15510), .A2(n15522), .B1(n15521), .B2(n15509), .ZN(
        n15511) );
  NOR2_X1 U17037 ( .A1(n15512), .A2(n15511), .ZN(n15541) );
  INV_X1 U17038 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15513) );
  AOI22_X1 U17039 ( .A1(n15528), .A2(n15541), .B1(n15513), .B2(n15526), .ZN(
        P3_U3411) );
  INV_X1 U17040 ( .A(n15514), .ZN(n15518) );
  AOI211_X1 U17041 ( .C1(n15518), .C2(n15517), .A(n15516), .B(n15515), .ZN(
        n15543) );
  INV_X1 U17042 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15519) );
  AOI22_X1 U17043 ( .A1(n15528), .A2(n15543), .B1(n15519), .B2(n15526), .ZN(
        P3_U3414) );
  OAI22_X1 U17044 ( .A1(n15523), .A2(n15522), .B1(n15521), .B2(n15520), .ZN(
        n15524) );
  NOR2_X1 U17045 ( .A1(n15525), .A2(n15524), .ZN(n15546) );
  INV_X1 U17046 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15527) );
  AOI22_X1 U17047 ( .A1(n15528), .A2(n15546), .B1(n15527), .B2(n15526), .ZN(
        P3_U3420) );
  AOI22_X1 U17048 ( .A1(n15547), .A2(n15530), .B1(n15529), .B2(n15544), .ZN(
        P3_U3460) );
  AOI22_X1 U17049 ( .A1(n15547), .A2(n15531), .B1(n10162), .B2(n15544), .ZN(
        P3_U3461) );
  AOI22_X1 U17050 ( .A1(n15547), .A2(n15533), .B1(n15532), .B2(n15544), .ZN(
        P3_U3462) );
  AOI22_X1 U17051 ( .A1(n15547), .A2(n15535), .B1(n15534), .B2(n15544), .ZN(
        P3_U3463) );
  AOI22_X1 U17052 ( .A1(n15547), .A2(n15537), .B1(n15536), .B2(n15544), .ZN(
        P3_U3464) );
  INV_X1 U17053 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15538) );
  AOI22_X1 U17054 ( .A1(n15547), .A2(n15539), .B1(n15538), .B2(n15544), .ZN(
        P3_U3465) );
  AOI22_X1 U17055 ( .A1(n15547), .A2(n15541), .B1(n15540), .B2(n15544), .ZN(
        P3_U3466) );
  INV_X1 U17056 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15542) );
  AOI22_X1 U17057 ( .A1(n15547), .A2(n15543), .B1(n15542), .B2(n15544), .ZN(
        P3_U3467) );
  INV_X1 U17058 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n15545) );
  AOI22_X1 U17059 ( .A1(n15547), .A2(n15546), .B1(n15545), .B2(n15544), .ZN(
        P3_U3469) );
  OAI21_X1 U17060 ( .B1(n15550), .B2(n15549), .A(n15548), .ZN(SUB_1596_U59) );
  OAI21_X1 U17061 ( .B1(n15553), .B2(n15552), .A(n15551), .ZN(SUB_1596_U58) );
  XOR2_X1 U17062 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15554), .Z(SUB_1596_U53) );
  OAI21_X1 U17063 ( .B1(n15557), .B2(n15556), .A(n15555), .ZN(SUB_1596_U56) );
  AOI21_X1 U17064 ( .B1(n15560), .B2(n15559), .A(n15558), .ZN(n15561) );
  XOR2_X1 U17065 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15561), .Z(SUB_1596_U60) );
  AOI21_X1 U17066 ( .B1(n15564), .B2(n15563), .A(n15562), .ZN(SUB_1596_U5) );
  INV_X2 U7528 ( .A(n8456), .ZN(n8439) );
  AND4_X4 U10841 ( .A1(n8469), .A2(n8468), .A3(n8467), .A4(n8466), .ZN(n9646)
         );
  CLKBUF_X1 U7389 ( .A(n8128), .Z(n6846) );
  INV_X1 U7421 ( .A(n12161), .ZN(n12171) );
  CLKBUF_X1 U7439 ( .A(n12379), .Z(n6823) );
  CLKBUF_X1 U7506 ( .A(n6820), .Z(n6650) );
  CLKBUF_X1 U7893 ( .A(n8460), .Z(n6637) );
  CLKBUF_X2 U7969 ( .A(n8481), .Z(n9035) );
  NAND2_X1 U8053 ( .A1(n8460), .A2(n10827), .ZN(n10184) );
  CLKBUF_X2 U8069 ( .A(n11759), .Z(n6649) );
  CLKBUF_X1 U9766 ( .A(n7880), .Z(n7908) );
endmodule

