

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput0, keyinput1, keyinput2, 
        keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, 
        keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, 
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, 
        keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, 
        keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, 
        keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, 
        keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, 
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, 
        keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, 
        keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, 
        keyinput63 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2957, n2958, n2959, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668;

  AND2_X1 U3405 ( .A1(n4100), .A2(n5149), .ZN(n5138) );
  INV_X1 U3406 ( .A(n5965), .ZN(n5948) );
  AND2_X1 U3407 ( .A1(n4181), .A2(n4180), .ZN(n3106) );
  OAI21_X1 U3408 ( .B1(n4729), .B2(n4175), .A(n4147), .ZN(n4149) );
  AOI21_X1 U3409 ( .B1(n4646), .B2(n6530), .A(n3317), .ZN(n3368) );
  NAND2_X2 U3410 ( .A1(n4003), .A2(n4248), .ZN(n4087) );
  CLKBUF_X2 U3411 ( .A(n3207), .Z(n3879) );
  NAND2_X1 U3412 ( .A1(n3293), .A2(n3291), .ZN(n3298) );
  CLKBUF_X2 U3413 ( .A(n3386), .Z(n3843) );
  CLKBUF_X2 U3414 ( .A(n3217), .Z(n3885) );
  CLKBUF_X2 U3415 ( .A(n3179), .Z(n3380) );
  CLKBUF_X2 U3416 ( .A(n3201), .Z(n3860) );
  CLKBUF_X2 U3417 ( .A(n3396), .Z(n3387) );
  BUF_X2 U3418 ( .A(n3188), .Z(n3884) );
  CLKBUF_X2 U3419 ( .A(n3281), .Z(n3787) );
  CLKBUF_X1 U3420 ( .A(n3178), .Z(n4685) );
  NAND4_X2 U3421 ( .A1(n3200), .A2(n3199), .A3(n3198), .A4(n3197), .ZN(n3236)
         );
  AND4_X1 U3422 ( .A1(n3131), .A2(n3130), .A3(n3129), .A4(n3128), .ZN(n3137)
         );
  AND4_X1 U3423 ( .A1(n3117), .A2(n3116), .A3(n3115), .A4(n3114), .ZN(n3127)
         );
  NOR2_X1 U3424 ( .A1(n3268), .A2(n3978), .ZN(n2975) );
  NOR2_X1 U3425 ( .A1(n2975), .A2(n4669), .ZN(n3026) );
  CLKBUF_X2 U3426 ( .A(n3206), .Z(n3837) );
  AND2_X1 U3427 ( .A1(n3247), .A2(n4523), .ZN(n3263) );
  AND4_X1 U3428 ( .A1(n3125), .A2(n3124), .A3(n3123), .A4(n3122), .ZN(n3126)
         );
  AND2_X1 U3429 ( .A1(n3268), .A2(n2985), .ZN(n4163) );
  AND2_X1 U3430 ( .A1(n3294), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3930) );
  OR2_X1 U3431 ( .A1(n3904), .A2(n3236), .ZN(n4273) );
  AND2_X1 U3432 ( .A1(n4059), .A2(n3020), .ZN(n5118) );
  OR2_X1 U3433 ( .A1(n4729), .A2(n3612), .ZN(n3367) );
  INV_X1 U3434 ( .A(n2991), .ZN(n5587) );
  NAND2_X1 U3435 ( .A1(n3361), .A2(n3360), .ZN(n4729) );
  NAND2_X2 U3436 ( .A1(n3961), .A2(n3960), .ZN(n4540) );
  INV_X1 U3437 ( .A(n5899), .ZN(n4228) );
  INV_X1 U3438 ( .A(n2979), .ZN(n5310) );
  OAI21_X1 U3440 ( .B1(n5496), .B2(n5599), .A(n5495), .ZN(n5497) );
  NAND2_X1 U3441 ( .A1(n4254), .A2(n4253), .ZN(n4292) );
  OAI21_X1 U3442 ( .B1(n5209), .B2(n5208), .A(n5207), .ZN(n5496) );
  XOR2_X1 U3443 ( .A(n3099), .B(n4202), .Z(n2957) );
  AND4_X1 U3444 ( .A1(n3155), .A2(n3154), .A3(n3153), .A4(n3152), .ZN(n2958)
         );
  AND2_X2 U34450 ( .A1(n3137), .A2(n3136), .ZN(n2959) );
  NOR2_X1 U34460 ( .A1(n3243), .A2(n4681), .ZN(n4484) );
  OAI22_X1 U34470 ( .A1(n5584), .A2(n4189), .B1(n5587), .B2(n4188), .ZN(n5567)
         );
  AND4_X2 U34480 ( .A1(n3055), .A2(n3054), .A3(n3053), .A4(n3030), .ZN(n5584)
         );
  NOR2_X2 U3449 ( .A1(n5211), .A2(n3993), .ZN(n5202) );
  OR2_X2 U34510 ( .A1(n3106), .A2(n3107), .ZN(n3004) );
  NOR2_X2 U34530 ( .A1(n5674), .A2(n4426), .ZN(n5662) );
  OAI22_X1 U3454 ( .A1(n5567), .A2(n4191), .B1(n4190), .B2(n2992), .ZN(n3052)
         );
  NAND2_X2 U34550 ( .A1(n3338), .A2(n3337), .ZN(n4771) );
  NAND2_X1 U34560 ( .A1(n3299), .A2(n3298), .ZN(n3320) );
  OR2_X1 U3458 ( .A1(n4274), .A2(n4256), .ZN(n4527) );
  AND2_X2 U34590 ( .A1(n3242), .A2(n2990), .ZN(n2974) );
  CLKBUF_X1 U34600 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n2983) );
  AOI21_X1 U34610 ( .B1(n4443), .B2(n6104), .A(n3105), .ZN(n4447) );
  AND2_X1 U34620 ( .A1(n4211), .A2(n4210), .ZN(n4212) );
  AOI21_X1 U34630 ( .B1(n3098), .B2(n2994), .A(n4200), .ZN(n5487) );
  OAI21_X1 U34640 ( .B1(n4450), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n5587), .ZN(n2978) );
  OR2_X1 U34650 ( .A1(n4449), .A2(n5509), .ZN(n4450) );
  NAND2_X1 U3466 ( .A1(n4234), .A2(n4233), .ZN(n4446) );
  OR2_X1 U3467 ( .A1(n5542), .A2(n2981), .ZN(n2980) );
  NOR2_X1 U34680 ( .A1(n4475), .A2(n4474), .ZN(n4473) );
  AOI211_X1 U34690 ( .C1(REIP_REG_27__SCAN_IN), .C2(n5221), .A(n5217), .B(
        n5216), .ZN(n5218) );
  OAI21_X1 U34700 ( .B1(n3076), .B2(n3073), .A(n3009), .ZN(n3072) );
  NAND2_X1 U34710 ( .A1(n2964), .A2(n2961), .ZN(n3062) );
  XNOR2_X1 U34720 ( .A(n4092), .B(n4218), .ZN(n5196) );
  NAND2_X1 U34730 ( .A1(n2964), .A2(n3103), .ZN(n2963) );
  NOR2_X1 U34740 ( .A1(n4193), .A2(n3079), .ZN(n3078) );
  AND2_X1 U3475 ( .A1(n4162), .A2(n3103), .ZN(n2961) );
  AND2_X1 U3476 ( .A1(n4488), .A2(n3083), .ZN(n5199) );
  OR2_X1 U3477 ( .A1(n5052), .A2(n4186), .ZN(n3054) );
  INV_X1 U3478 ( .A(n3066), .ZN(n2965) );
  NOR3_X1 U3479 ( .A1(n3095), .A2(n3857), .A3(n3098), .ZN(n3094) );
  XNOR2_X1 U3480 ( .A(n4161), .B(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3066)
         );
  NAND2_X1 U3481 ( .A1(n4152), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3103)
         );
  AND2_X1 U3482 ( .A1(n3004), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4186)
         );
  XNOR2_X1 U3483 ( .A(n2991), .B(n5773), .ZN(n5023) );
  AND3_X1 U3484 ( .A1(n5305), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .ZN(n5273) );
  INV_X1 U3485 ( .A(n3106), .ZN(n2992) );
  NAND2_X1 U3486 ( .A1(n3367), .A2(n3366), .ZN(n4586) );
  XNOR2_X1 U3487 ( .A(n4149), .B(n4148), .ZN(n4633) );
  AND2_X1 U3488 ( .A1(n5975), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5392) );
  CLKBUF_X1 U3489 ( .A(n4653), .Z(n6172) );
  OR2_X1 U3490 ( .A1(n3359), .A2(n4771), .ZN(n3361) );
  NOR2_X1 U3491 ( .A1(n5011), .A2(n5028), .ZN(n5027) );
  NAND2_X1 U3492 ( .A1(n5610), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4141)
         );
  AND2_X1 U3493 ( .A1(n3417), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4568) );
  CLKBUF_X1 U3494 ( .A(n4658), .Z(n6307) );
  NAND3_X1 U3495 ( .A1(n3958), .A2(n3957), .A3(n3956), .ZN(n3961) );
  NAND2_X1 U3496 ( .A1(n3412), .A2(n3297), .ZN(n3372) );
  NAND2_X1 U3497 ( .A1(n2967), .A2(n3304), .ZN(n3318) );
  NAND2_X1 U3498 ( .A1(n3237), .A2(STATE2_REG_0__SCAN_IN), .ZN(n2969) );
  NAND2_X1 U3499 ( .A1(n3321), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n2967) );
  NAND2_X1 U3500 ( .A1(n4005), .A2(n4004), .ZN(n4007) );
  NAND2_X1 U3501 ( .A1(n3964), .A2(n3242), .ZN(n4105) );
  OR2_X1 U3502 ( .A1(n3414), .A2(n3413), .ZN(n3415) );
  NAND2_X1 U3503 ( .A1(n4237), .A2(n2974), .ZN(n3247) );
  CLKBUF_X2 U3504 ( .A(n4012), .Z(n4576) );
  INV_X1 U3505 ( .A(n2974), .ZN(n6662) );
  NOR2_X1 U3506 ( .A1(n4527), .A2(n2972), .ZN(n4528) );
  AND2_X1 U3507 ( .A1(n4104), .A2(n3908), .ZN(n3935) );
  NAND2_X1 U3508 ( .A1(n3306), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3923) );
  AND2_X1 U3509 ( .A1(n3156), .A2(n3258), .ZN(n3241) );
  CLKBUF_X1 U3510 ( .A(n3258), .Z(n4661) );
  AND2_X1 U3511 ( .A1(n3006), .A2(STATE2_REG_0__SCAN_IN), .ZN(n2966) );
  NAND2_X1 U3512 ( .A1(n3230), .A2(n2986), .ZN(n3904) );
  NAND2_X1 U3513 ( .A1(n4250), .A2(n2986), .ZN(n3065) );
  NAND2_X1 U3514 ( .A1(n3001), .A2(n2958), .ZN(n3258) );
  BUF_X2 U3515 ( .A(n3248), .Z(n4674) );
  OR2_X1 U3516 ( .A1(n3393), .A2(n3392), .ZN(n4130) );
  OR2_X1 U3517 ( .A1(n3407), .A2(n3406), .ZN(n4182) );
  NAND2_X1 U3518 ( .A1(n3147), .A2(n3146), .ZN(n3248) );
  AND4_X1 U3519 ( .A1(n3205), .A2(n3204), .A3(n3203), .A4(n3202), .ZN(n3225)
         );
  AND4_X1 U3520 ( .A1(n3192), .A2(n3191), .A3(n3190), .A4(n3189), .ZN(n3198)
         );
  AND4_X1 U3521 ( .A1(n3196), .A2(n3195), .A3(n3194), .A4(n3193), .ZN(n3197)
         );
  AND4_X1 U3522 ( .A1(n3141), .A2(n3140), .A3(n3139), .A4(n3138), .ZN(n3147)
         );
  AND4_X1 U3523 ( .A1(n3183), .A2(n3182), .A3(n3181), .A4(n3180), .ZN(n3200)
         );
  AND4_X1 U3524 ( .A1(n3216), .A2(n3215), .A3(n3214), .A4(n3213), .ZN(n3223)
         );
  AND4_X1 U3525 ( .A1(n3187), .A2(n3186), .A3(n3185), .A4(n3184), .ZN(n3199)
         );
  AND4_X1 U3526 ( .A1(n3145), .A2(n3144), .A3(n3143), .A4(n3142), .ZN(n3146)
         );
  BUF_X2 U3527 ( .A(n3379), .Z(n3779) );
  INV_X1 U3528 ( .A(n2970), .ZN(n5160) );
  AND2_X2 U3529 ( .A1(n3064), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3119)
         );
  AND2_X2 U3530 ( .A1(n3090), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3120)
         );
  AND2_X2 U3531 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4720) );
  NAND2_X1 U3532 ( .A1(n2962), .A2(n4162), .ZN(n4886) );
  NAND2_X1 U3533 ( .A1(n2965), .A2(n2963), .ZN(n2962) );
  XNOR2_X1 U3534 ( .A(n2965), .B(n2963), .ZN(n6143) );
  NAND2_X1 U3535 ( .A1(n4623), .A2(n4624), .ZN(n2964) );
  NAND2_X1 U3536 ( .A1(n3237), .A2(n2966), .ZN(n3299) );
  NAND3_X1 U3537 ( .A1(n3320), .A2(n3319), .A3(n3318), .ZN(n4722) );
  NAND2_X2 U3538 ( .A1(n2969), .A2(n2968), .ZN(n3319) );
  AOI21_X2 U3539 ( .B1(n3252), .B2(n3016), .A(n3253), .ZN(n2968) );
  CLKBUF_X1 U3540 ( .A(n2971), .Z(n2970) );
  AND2_X4 U3541 ( .A1(n3118), .A2(n2971), .ZN(n3280) );
  AND2_X2 U3542 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n2971) );
  NAND2_X1 U3543 ( .A1(n2970), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4707) );
  NAND2_X1 U3544 ( .A1(n2970), .A2(n3425), .ZN(n5157) );
  AND2_X2 U3545 ( .A1(n2971), .A2(n4720), .ZN(n3217) );
  AND2_X2 U3546 ( .A1(n3121), .A2(n2971), .ZN(n3179) );
  AND2_X2 U3547 ( .A1(n3120), .A2(n2971), .ZN(n3188) );
  NAND2_X1 U3548 ( .A1(n2973), .A2(n5160), .ZN(n2972) );
  INV_X1 U3549 ( .A(n4526), .ZN(n2973) );
  AOI21_X1 U3550 ( .B1(n2974), .B2(n3261), .A(n6538), .ZN(n3262) );
  OAI211_X1 U3551 ( .C1(n2975), .C2(n2985), .A(n4534), .B(n3267), .ZN(n3249)
         );
  NAND2_X1 U3552 ( .A1(n4633), .A2(n4634), .ZN(n4151) );
  NAND2_X1 U3553 ( .A1(n2978), .A2(n2976), .ZN(n4451) );
  NAND3_X1 U3554 ( .A1(n2977), .A2(n2992), .A3(n2980), .ZN(n2976) );
  NAND2_X1 U3555 ( .A1(n4449), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n2977) );
  NOR2_X2 U3556 ( .A1(n5542), .A2(n5718), .ZN(n5509) );
  AND2_X4 U3557 ( .A1(n5321), .A2(n5322), .ZN(n2979) );
  OR2_X1 U3558 ( .A1(n5718), .A2(n2982), .ZN(n2981) );
  INV_X1 U3559 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n2982) );
  NOR2_X2 U3560 ( .A1(n3264), .A2(n4273), .ZN(n3964) );
  AND2_X2 U3561 ( .A1(n3119), .A2(n4720), .ZN(n3379) );
  AND2_X2 U3562 ( .A1(n3119), .A2(n3118), .ZN(n3279) );
  AOI21_X1 U3563 ( .B1(n3206), .B2(INSTQUEUE_REG_4__1__SCAN_IN), .A(n3212), 
        .ZN(n3224) );
  BUF_X2 U3564 ( .A(n3279), .Z(n3394) );
  AND2_X2 U3565 ( .A1(n3120), .A2(n4532), .ZN(n3396) );
  AND2_X2 U3566 ( .A1(n4532), .A2(n4720), .ZN(n3201) );
  INV_X1 U3567 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4529) );
  NOR2_X2 U3568 ( .A1(n5041), .A2(n3086), .ZN(n5313) );
  INV_X1 U3569 ( .A(n6662), .ZN(n2984) );
  BUF_X2 U3570 ( .A(n3244), .Z(n3268) );
  AND4_X1 U3571 ( .A1(n3221), .A2(n3220), .A3(n3219), .A4(n3218), .ZN(n3222)
         );
  INV_X1 U3572 ( .A(n2959), .ZN(n2985) );
  NAND2_X1 U3573 ( .A1(n3137), .A2(n3136), .ZN(n2986) );
  NAND2_X2 U3574 ( .A1(n3257), .A2(n2986), .ZN(n3228) );
  INV_X2 U3575 ( .A(n3178), .ZN(n3257) );
  INV_X1 U3576 ( .A(n2987), .ZN(n4246) );
  AND2_X2 U3577 ( .A1(n4102), .A2(n3232), .ZN(n2987) );
  NAND2_X1 U3578 ( .A1(n4151), .A2(n4150), .ZN(n4623) );
  CLKBUF_X1 U3579 ( .A(n4722), .Z(n2988) );
  INV_X1 U3580 ( .A(n4771), .ZN(n2989) );
  AND2_X1 U3581 ( .A1(n4771), .A2(n3092), .ZN(n3027) );
  AOI21_X4 U3582 ( .B1(n5337), .B2(n3614), .A(n3613), .ZN(n5321) );
  OR2_X1 U3583 ( .A1(n3228), .A2(n3248), .ZN(n3157) );
  NAND2_X2 U3584 ( .A1(n3569), .A2(n3568), .ZN(n5337) );
  AND2_X4 U3585 ( .A1(n4526), .A2(n4720), .ZN(n3386) );
  NOR2_X4 U3586 ( .A1(n4840), .A2(n3503), .ZN(n5007) );
  NAND4_X1 U3587 ( .A1(n3200), .A2(n3199), .A3(n3198), .A4(n3197), .ZN(n2990)
         );
  INV_X2 U3588 ( .A(n3236), .ZN(n4669) );
  NOR2_X2 U3589 ( .A1(n3265), .A2(n4262), .ZN(n4102) );
  INV_X1 U3590 ( .A(n3106), .ZN(n2991) );
  INV_X1 U3591 ( .A(n3352), .ZN(n3351) );
  OR2_X1 U3592 ( .A1(n5242), .A2(n3856), .ZN(n3857) );
  INV_X1 U3593 ( .A(n3584), .ZN(n3612) );
  AND2_X1 U3594 ( .A1(n4802), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4201) );
  INV_X1 U3595 ( .A(n3455), .ZN(n3726) );
  NOR2_X1 U3596 ( .A1(n4685), .A2(n4802), .ZN(n3584) );
  NAND2_X1 U3597 ( .A1(n4802), .A2(n6432), .ZN(n3832) );
  NAND2_X1 U3598 ( .A1(n3244), .A2(n3243), .ZN(n4214) );
  NAND2_X1 U3599 ( .A1(n4099), .A2(n3104), .ZN(n5149) );
  INV_X1 U3600 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4333) );
  AND2_X1 U3601 ( .A1(n3534), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3550)
         );
  AND2_X1 U3602 ( .A1(n3109), .A2(n3068), .ZN(n3067) );
  INV_X1 U3603 ( .A(n5129), .ZN(n3068) );
  NAND2_X1 U3604 ( .A1(n2991), .A2(n4232), .ZN(n4233) );
  OAI21_X1 U3605 ( .B1(n5952), .B2(n5423), .A(n3045), .ZN(n3044) );
  AOI22_X1 U3606 ( .A1(n5732), .A2(n5927), .B1(n5960), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3045) );
  NAND2_X1 U3607 ( .A1(n4208), .A2(n3013), .ZN(n5965) );
  INV_X1 U3608 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3090) );
  INV_X1 U3609 ( .A(n4204), .ZN(n3303) );
  OAI21_X1 U3610 ( .B1(n3947), .B2(n4823), .A(n3448), .ZN(n3458) );
  AND2_X1 U3611 ( .A1(n3471), .A2(n3470), .ZN(n3477) );
  AND2_X1 U3612 ( .A1(n3350), .A2(n3349), .ZN(n3352) );
  NOR2_X1 U3613 ( .A1(n3248), .A2(n3178), .ZN(n3232) );
  OR2_X1 U3614 ( .A1(n5269), .A2(n4576), .ZN(n4083) );
  INV_X1 U3615 ( .A(n5241), .ZN(n3096) );
  NOR2_X1 U3616 ( .A1(n5529), .A2(n3033), .ZN(n3032) );
  NOR2_X1 U3617 ( .A1(n4333), .A2(n3036), .ZN(n3035) );
  INV_X1 U3618 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3036) );
  INV_X1 U3619 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3051) );
  NAND2_X1 U3620 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3426) );
  INV_X1 U3621 ( .A(n3832), .ZN(n3903) );
  NAND2_X1 U3622 ( .A1(n3018), .A2(n4039), .ZN(n3089) );
  INV_X1 U3623 ( .A(n5765), .ZN(n4039) );
  INV_X1 U3624 ( .A(n5023), .ZN(n3030) );
  INV_X1 U3625 ( .A(n5058), .ZN(n4029) );
  INV_X1 U3626 ( .A(n4920), .ZN(n3082) );
  NAND2_X1 U3627 ( .A1(n4888), .A2(n4921), .ZN(n4920) );
  INV_X1 U3628 ( .A(n4630), .ZN(n4018) );
  INV_X1 U3629 ( .A(n4083), .ZN(n4074) );
  NAND2_X1 U3630 ( .A1(n3268), .A2(n4669), .ZN(n4534) );
  INV_X1 U3631 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6306) );
  AND2_X1 U3632 ( .A1(n6504), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6206)
         );
  INV_X1 U3633 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6504) );
  NAND2_X1 U3634 ( .A1(n2987), .A2(n4248), .ZN(n3963) );
  INV_X1 U3635 ( .A(n5939), .ZN(n5381) );
  AND2_X1 U3636 ( .A1(n2959), .A2(n4484), .ZN(n3226) );
  XNOR2_X1 U3637 ( .A(n3976), .B(n4225), .ZN(n4208) );
  AND2_X1 U3638 ( .A1(n3733), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3874)
         );
  INV_X1 U3639 ( .A(n3695), .ZN(n3696) );
  NAND2_X1 U3640 ( .A1(n3696), .A2(n3032), .ZN(n3731) );
  OR2_X1 U3641 ( .A1(n3667), .A2(n3666), .ZN(n3695) );
  INV_X1 U3642 ( .A(n3626), .ZN(n3627) );
  NAND2_X1 U3643 ( .A1(n2993), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3626)
         );
  AND2_X1 U3644 ( .A1(n3567), .A2(n3566), .ZN(n5873) );
  NOR2_X1 U3645 ( .A1(n3520), .A2(n3519), .ZN(n3534) );
  NAND2_X1 U3646 ( .A1(n4540), .A2(n4545), .ZN(n4548) );
  NOR2_X1 U3647 ( .A1(n5490), .A2(n3070), .ZN(n5164) );
  NAND2_X1 U3648 ( .A1(n5587), .A2(n5638), .ZN(n3070) );
  NOR2_X1 U3649 ( .A1(n4064), .A2(n5283), .ZN(n3081) );
  AND2_X1 U3650 ( .A1(n4066), .A2(n4065), .ZN(n5253) );
  NAND2_X1 U3651 ( .A1(n4059), .A2(n2996), .ZN(n5256) );
  AOI21_X1 U3652 ( .B1(n5750), .B2(n3078), .A(n3028), .ZN(n5528) );
  NAND2_X1 U3653 ( .A1(n3076), .A2(n3029), .ZN(n3028) );
  NAND2_X1 U3654 ( .A1(n2992), .A2(n4231), .ZN(n3029) );
  INV_X1 U3655 ( .A(n3017), .ZN(n3075) );
  AND2_X1 U3656 ( .A1(n4051), .A2(n4050), .ZN(n5323) );
  NAND2_X1 U3657 ( .A1(n5810), .A2(n5814), .ZN(n5737) );
  NAND2_X1 U3658 ( .A1(n4161), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4162)
         );
  INV_X1 U3659 ( .A(n3248), .ZN(n4256) );
  CLKBUF_X1 U3660 ( .A(n4646), .Z(n4647) );
  NAND2_X1 U3661 ( .A1(n6530), .A2(n4659), .ZN(n6312) );
  NOR2_X1 U3662 ( .A1(n4291), .A2(n3242), .ZN(n6499) );
  AND2_X1 U3663 ( .A1(n6172), .A2(n2989), .ZN(n6277) );
  AND2_X1 U3664 ( .A1(n4652), .A2(n5062), .ZN(n5063) );
  AND2_X1 U3665 ( .A1(n5963), .A2(n4647), .ZN(n6437) );
  AND2_X1 U3666 ( .A1(n4647), .A2(n4520), .ZN(n6274) );
  INV_X1 U3667 ( .A(n6312), .ZN(n4852) );
  AND2_X1 U3668 ( .A1(n4654), .A2(n6172), .ZN(n4662) );
  OR2_X1 U3669 ( .A1(n4239), .A2(n3904), .ZN(n6517) );
  OR2_X1 U3670 ( .A1(n4246), .A2(n6662), .ZN(n6527) );
  INV_X1 U3671 ( .A(n5960), .ZN(n5908) );
  AND2_X1 U3672 ( .A1(n5392), .A2(n4095), .ZN(n5927) );
  OR2_X1 U3673 ( .A1(n6528), .A2(n3973), .ZN(n3974) );
  INV_X1 U3674 ( .A(n5961), .ZN(n5952) );
  OR2_X1 U3675 ( .A1(n5987), .A2(n4492), .ZN(n4493) );
  NAND2_X1 U3676 ( .A1(n5987), .A2(n3231), .ZN(n5433) );
  INV_X1 U3677 ( .A(n5991), .ZN(n5473) );
  OAI21_X1 U3678 ( .B1(n5170), .B2(n3855), .A(n2994), .ZN(n5178) );
  NAND2_X1 U3679 ( .A1(n4436), .A2(n4098), .ZN(n4100) );
  OR2_X1 U3680 ( .A1(n5660), .A2(n6100), .ZN(n4480) );
  NAND2_X1 U3681 ( .A1(n6112), .A2(n5611), .ZN(n5594) );
  OR2_X1 U3682 ( .A1(n6647), .A2(n6543), .ZN(n6122) );
  NAND2_X1 U3683 ( .A1(n4203), .A2(n6380), .ZN(n5599) );
  INV_X1 U3684 ( .A(n5594), .ZN(n6105) );
  NAND2_X1 U3685 ( .A1(n4091), .A2(n4090), .ZN(n4092) );
  NAND2_X1 U3686 ( .A1(n5199), .A2(n4213), .ZN(n4091) );
  OR2_X1 U3687 ( .A1(n5199), .A2(n3245), .ZN(n4090) );
  XNOR2_X1 U3688 ( .A(n4466), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5137)
         );
  NAND2_X1 U3689 ( .A1(n3002), .A2(n4464), .ZN(n4466) );
  XNOR2_X1 U3690 ( .A(n3031), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5669)
         );
  OAI22_X1 U3691 ( .A1(n4446), .A2(n4445), .B1(n5511), .B2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3031) );
  INV_X1 U3692 ( .A(n6307), .ZN(n5062) );
  NOR2_X2 U3693 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6380) );
  INV_X1 U3694 ( .A(n6380), .ZN(n6435) );
  OR2_X1 U3695 ( .A1(n4766), .A2(n5062), .ZN(n4898) );
  NAND2_X1 U3696 ( .A1(n3241), .A2(n4256), .ZN(n4237) );
  INV_X1 U3697 ( .A(n3905), .ZN(n3920) );
  NAND2_X1 U3698 ( .A1(n3927), .A2(n3926), .ZN(n3945) );
  XNOR2_X1 U3699 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3944) );
  NAND2_X1 U3700 ( .A1(n3228), .A2(n4674), .ZN(n3267) );
  AND2_X1 U3701 ( .A1(n3351), .A2(n3458), .ZN(n3092) );
  INV_X1 U3702 ( .A(n3360), .ZN(n3093) );
  OR2_X1 U3703 ( .A1(n3447), .A2(n3446), .ZN(n4157) );
  OR2_X1 U3704 ( .A1(n3348), .A2(n3347), .ZN(n4154) );
  OR2_X1 U3705 ( .A1(n3316), .A2(n3315), .ZN(n4123) );
  INV_X1 U3706 ( .A(n4123), .ZN(n4116) );
  AOI22_X1 U3707 ( .A1(n3395), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3132) );
  OR2_X1 U3708 ( .A1(n3336), .A2(n3335), .ZN(n4146) );
  INV_X1 U3709 ( .A(n3306), .ZN(n3294) );
  NAND2_X1 U3710 ( .A1(n3930), .A2(n4163), .ZN(n3938) );
  NAND2_X1 U3711 ( .A1(n3256), .A2(n3255), .ZN(n3293) );
  AOI22_X1 U3712 ( .A1(n3208), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3201), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3151) );
  INV_X1 U3713 ( .A(n4199), .ZN(n3095) );
  NOR2_X1 U3714 ( .A1(n3826), .A2(n4440), .ZN(n3812) );
  AND2_X1 U3715 ( .A1(n5285), .A2(n3101), .ZN(n3100) );
  NOR2_X1 U3716 ( .A1(n5300), .A2(n5312), .ZN(n3101) );
  NOR2_X1 U3717 ( .A1(n3042), .A2(n3040), .ZN(n3039) );
  NOR2_X1 U3718 ( .A1(n4527), .A2(n6530), .ZN(n3900) );
  AND2_X1 U3719 ( .A1(n5008), .A2(n5018), .ZN(n3091) );
  INV_X1 U3720 ( .A(n3426), .ZN(n3362) );
  INV_X1 U3721 ( .A(n4196), .ZN(n3073) );
  INV_X1 U3722 ( .A(n5751), .ZN(n3079) );
  INV_X1 U3723 ( .A(n3077), .ZN(n3076) );
  OAI21_X1 U3724 ( .B1(n4193), .B2(n3017), .A(n4192), .ZN(n3077) );
  INV_X1 U3725 ( .A(n5013), .ZN(n4033) );
  NAND2_X1 U3726 ( .A1(n3066), .A2(n4162), .ZN(n3061) );
  INV_X1 U3727 ( .A(n4130), .ZN(n4135) );
  NAND2_X1 U3728 ( .A1(n3288), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3289) );
  NAND2_X1 U3729 ( .A1(n3246), .A2(n3245), .ZN(n4523) );
  INV_X1 U3730 ( .A(n3904), .ZN(n3246) );
  INV_X1 U3731 ( .A(n3964), .ZN(n4291) );
  AND2_X1 U3732 ( .A1(n3252), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3321) );
  NAND4_X2 U3733 ( .A1(n3225), .A2(n3224), .A3(n3223), .A4(n3222), .ZN(n3244)
         );
  AOI22_X1 U3734 ( .A1(n3279), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3201), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3116) );
  INV_X1 U3735 ( .A(n3938), .ZN(n3959) );
  INV_X1 U3736 ( .A(n3923), .ZN(n3955) );
  AND2_X1 U3737 ( .A1(n3954), .A2(n3953), .ZN(n3965) );
  OR2_X1 U3738 ( .A1(n3952), .A2(n3951), .ZN(n3954) );
  AND2_X1 U3739 ( .A1(n6162), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3951)
         );
  OR2_X1 U3740 ( .A1(n6647), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4204) );
  INV_X1 U3741 ( .A(n4012), .ZN(n4483) );
  OR2_X1 U3742 ( .A1(n4658), .A2(n4274), .ZN(n3417) );
  INV_X1 U3743 ( .A(n3878), .ZN(n3975) );
  NAND2_X1 U3744 ( .A1(n3874), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3875)
         );
  OR2_X1 U3745 ( .A1(n3875), .A2(n5484), .ZN(n3878) );
  NOR2_X1 U3746 ( .A1(n3857), .A2(n3098), .ZN(n3097) );
  AND2_X1 U3747 ( .A1(n3732), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3733)
         );
  INV_X1 U3748 ( .A(n3815), .ZN(n3732) );
  NAND2_X1 U3749 ( .A1(n3812), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3815)
         );
  NAND2_X1 U3750 ( .A1(n3696), .A2(n2999), .ZN(n3824) );
  OR2_X1 U3751 ( .A1(n3824), .A2(n5514), .ZN(n3826) );
  NAND2_X1 U3752 ( .A1(n3665), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3667)
         );
  INV_X1 U3753 ( .A(n3664), .ZN(n3665) );
  INV_X1 U3754 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3666) );
  NAND2_X1 U3755 ( .A1(n3627), .A2(n3038), .ZN(n3664) );
  AND2_X1 U3756 ( .A1(n3039), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3038)
         );
  CLKBUF_X1 U3757 ( .A(n5039), .Z(n5040) );
  NAND2_X1 U3758 ( .A1(n3514), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3520)
         );
  AND3_X1 U3759 ( .A1(n3500), .A2(n3499), .A3(n3498), .ZN(n5047) );
  AND2_X1 U3760 ( .A1(n3482), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3514)
         );
  AND2_X1 U3761 ( .A1(n3050), .A2(n3048), .ZN(n3482) );
  NOR2_X1 U3762 ( .A1(n3051), .A2(n3049), .ZN(n3048) );
  NOR2_X1 U3763 ( .A1(n3450), .A2(n3426), .ZN(n3050) );
  CLKBUF_X1 U3764 ( .A(n4840), .Z(n4841) );
  NOR2_X1 U3765 ( .A1(n3426), .A2(n3051), .ZN(n3047) );
  INV_X1 U3766 ( .A(n3450), .ZN(n3046) );
  NAND2_X1 U3767 ( .A1(n3362), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3451)
         );
  CLKBUF_X1 U3768 ( .A(n4585), .Z(n4749) );
  NOR2_X1 U3769 ( .A1(n5179), .A2(n3084), .ZN(n3083) );
  OR2_X1 U3770 ( .A1(n5214), .A2(n3085), .ZN(n3084) );
  INV_X1 U3771 ( .A(n5152), .ZN(n3085) );
  NAND2_X1 U3772 ( .A1(n5199), .A2(n5198), .ZN(n5197) );
  NOR2_X1 U3773 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n5587), .ZN(n4460)
         );
  AND2_X1 U3774 ( .A1(n4077), .A2(n4076), .ZN(n5119) );
  NAND2_X1 U3776 ( .A1(n3087), .A2(n4052), .ZN(n3086) );
  INV_X1 U3777 ( .A(n3089), .ZN(n3087) );
  NOR2_X1 U3778 ( .A1(n5041), .A2(n3089), .ZN(n5430) );
  NAND2_X1 U3779 ( .A1(n3088), .A2(n4039), .ZN(n5360) );
  INV_X1 U3780 ( .A(n5041), .ZN(n3088) );
  NAND2_X1 U3781 ( .A1(n3058), .A2(n3060), .ZN(n3053) );
  NOR2_X1 U3782 ( .A1(n4186), .A2(n3059), .ZN(n3058) );
  NAND2_X1 U3783 ( .A1(n2995), .A2(n3063), .ZN(n3059) );
  NAND2_X1 U3784 ( .A1(n4927), .A2(n3056), .ZN(n3055) );
  INV_X1 U3785 ( .A(n4745), .ZN(n3080) );
  NAND2_X1 U3786 ( .A1(n5737), .A2(n6151), .ZN(n5694) );
  NAND2_X1 U3787 ( .A1(n4615), .A2(n4142), .ZN(n4593) );
  OR2_X1 U3788 ( .A1(n5737), .A2(n5767), .ZN(n5696) );
  XNOR2_X1 U3789 ( .A(n4141), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4616)
         );
  CLKBUF_X1 U3790 ( .A(n4519), .Z(n4520) );
  OR2_X1 U3791 ( .A1(n4729), .A2(n6172), .ZN(n6382) );
  NAND2_X1 U3792 ( .A1(n3359), .A2(n4771), .ZN(n3360) );
  NAND2_X1 U3793 ( .A1(n6377), .A2(n5061), .ZN(n6337) );
  AND2_X1 U3794 ( .A1(n4652), .A2(n6307), .ZN(n6376) );
  INV_X1 U3795 ( .A(n6382), .ZN(n6377) );
  AND3_X1 U3796 ( .A1(n5061), .A2(n4771), .A3(n6172), .ZN(n4777) );
  INV_X1 U3797 ( .A(n4670), .ZN(n4690) );
  INV_X1 U3798 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n4725) );
  INV_X1 U3799 ( .A(n5904), .ZN(n5907) );
  AND2_X1 U3800 ( .A1(n5392), .A2(n3997), .ZN(n5961) );
  INV_X1 U3801 ( .A(n5507), .ZN(n5448) );
  OAI21_X1 U3802 ( .B1(n4536), .B2(n4108), .A(n4545), .ZN(n4109) );
  AND2_X1 U3803 ( .A1(n4521), .A2(n4485), .ZN(n4108) );
  INV_X1 U3804 ( .A(n5988), .ZN(n5476) );
  AND2_X1 U3805 ( .A1(n4551), .A2(n4550), .ZN(n6022) );
  NAND2_X1 U3806 ( .A1(n6092), .A2(n4549), .ZN(n4551) );
  INV_X1 U3807 ( .A(n6037), .ZN(n6086) );
  INV_X1 U3808 ( .A(n6092), .ZN(n6085) );
  INV_X1 U3809 ( .A(n6083), .ZN(n6090) );
  OAI21_X1 U3810 ( .B1(n2984), .B2(n6660), .A(n4514), .ZN(n6089) );
  OR2_X1 U3811 ( .A1(n4548), .A2(n6527), .ZN(n6092) );
  INV_X1 U3812 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5514) );
  XNOR2_X1 U3813 ( .A(n4446), .B(n4236), .ZN(n5519) );
  INV_X1 U3814 ( .A(n4235), .ZN(n4236) );
  NAND2_X1 U3815 ( .A1(n3696), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3697)
         );
  INV_X1 U3816 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5529) );
  NAND2_X1 U3817 ( .A1(n3627), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3645)
         );
  NAND2_X1 U3818 ( .A1(n3550), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3551)
         );
  INV_X1 U3819 ( .A(n6112), .ZN(n6094) );
  INV_X1 U3820 ( .A(n6100), .ZN(n6107) );
  INV_X2 U3821 ( .A(n5599), .ZN(n6104) );
  NAND2_X1 U3822 ( .A1(n3071), .A2(n3069), .ZN(n4198) );
  NOR2_X1 U3823 ( .A1(n4301), .A2(n4300), .ZN(n4302) );
  AND2_X1 U3824 ( .A1(n4059), .A2(n3081), .ZN(n5254) );
  NAND2_X1 U3825 ( .A1(n4059), .A2(n4058), .ZN(n5268) );
  XNOR2_X1 U3826 ( .A(n4451), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5707)
         );
  INV_X1 U3827 ( .A(n4450), .ZN(n5536) );
  OR2_X1 U3828 ( .A1(n5808), .A2(n5766), .ZN(n5816) );
  AND2_X1 U3829 ( .A1(n4934), .A2(n4933), .ZN(n6121) );
  INV_X1 U3830 ( .A(n5696), .ZN(n6153) );
  INV_X1 U3831 ( .A(n6142), .ZN(n6155) );
  INV_X1 U3833 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6162) );
  OAI21_X1 U3834 ( .B1(n4728), .B2(n6630), .A(n6312), .ZN(n6161) );
  NAND2_X1 U3835 ( .A1(n4725), .A2(n3238), .ZN(n6647) );
  INV_X1 U3836 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3425) );
  INV_X1 U3837 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4823) );
  NOR2_X1 U3838 ( .A1(n4801), .A2(n4800), .ZN(n4839) );
  OR2_X1 U3839 ( .A1(n4765), .A2(n4764), .ZN(n6163) );
  INV_X1 U3840 ( .A(n6199), .ZN(n4968) );
  OAI21_X1 U3841 ( .B1(n4942), .B2(n4943), .A(n5073), .ZN(n4966) );
  AND2_X1 U3842 ( .A1(n6184), .A2(n5063), .ZN(n6199) );
  OAI21_X1 U3843 ( .B1(n6183), .B2(n6182), .A(n6181), .ZN(n6201) );
  AND2_X1 U3844 ( .A1(n6184), .A2(n6376), .ZN(n6209) );
  INV_X1 U3845 ( .A(n6298), .ZN(n6270) );
  OAI211_X1 U3846 ( .C1(n6264), .C2(n3238), .A(n4978), .B(n6509), .ZN(n6267)
         );
  AND2_X1 U3847 ( .A1(n6277), .A2(n5063), .ZN(n6298) );
  INV_X1 U3848 ( .A(n6336), .ZN(n6310) );
  NOR2_X2 U3849 ( .A1(n6337), .A2(n6307), .ZN(n6369) );
  NAND2_X1 U3850 ( .A1(n6377), .A2(n5063), .ZN(n6400) );
  INV_X1 U3851 ( .A(n6400), .ZN(n6418) );
  INV_X1 U3852 ( .A(n6348), .ZN(n6431) );
  INV_X1 U3853 ( .A(n5079), .ZN(n6446) );
  INV_X1 U3854 ( .A(n6351), .ZN(n6447) );
  INV_X1 U3855 ( .A(n5068), .ZN(n6452) );
  INV_X1 U3856 ( .A(n6355), .ZN(n6453) );
  INV_X1 U3857 ( .A(n6358), .ZN(n6459) );
  INV_X1 U3858 ( .A(n5105), .ZN(n6464) );
  INV_X1 U3859 ( .A(n6361), .ZN(n6465) );
  INV_X1 U3860 ( .A(n5089), .ZN(n6470) );
  INV_X1 U3861 ( .A(n6364), .ZN(n6471) );
  INV_X1 U3862 ( .A(n5099), .ZN(n6476) );
  INV_X1 U3863 ( .A(n6367), .ZN(n6477) );
  INV_X1 U3864 ( .A(n5084), .ZN(n6483) );
  OAI21_X1 U3865 ( .B1(n4775), .B2(n4774), .A(n4773), .ZN(n4793) );
  AND2_X1 U3866 ( .A1(n4777), .A2(n5062), .ZN(n6486) );
  AND2_X1 U3867 ( .A1(n6104), .A2(DATAI_16_), .ZN(n6442) );
  AND2_X1 U3868 ( .A1(n6104), .A2(DATAI_17_), .ZN(n6448) );
  AND2_X1 U3869 ( .A1(n6104), .A2(DATAI_18_), .ZN(n6454) );
  AND2_X1 U3870 ( .A1(n6104), .A2(DATAI_20_), .ZN(n6466) );
  AND2_X1 U3871 ( .A1(n6104), .A2(DATAI_21_), .ZN(n6472) );
  AND2_X1 U3872 ( .A1(n6104), .A2(DATAI_22_), .ZN(n6478) );
  AND2_X1 U3873 ( .A1(n6104), .A2(DATAI_23_), .ZN(n6487) );
  AND2_X1 U3874 ( .A1(n6104), .A2(DATAI_24_), .ZN(n6379) );
  AND2_X1 U3875 ( .A1(n6104), .A2(DATAI_25_), .ZN(n6393) );
  NAND2_X1 U3876 ( .A1(DATAI_1_), .A2(n4852), .ZN(n6351) );
  AND2_X1 U3877 ( .A1(n6104), .A2(DATAI_26_), .ZN(n6352) );
  NAND2_X1 U3878 ( .A1(DATAI_2_), .A2(n4852), .ZN(n6355) );
  NAND2_X1 U3879 ( .A1(DATAI_3_), .A2(n4852), .ZN(n6358) );
  AND2_X1 U3880 ( .A1(n6104), .A2(DATAI_28_), .ZN(n6405) );
  NAND2_X1 U3881 ( .A1(DATAI_4_), .A2(n4852), .ZN(n6361) );
  AND2_X1 U3882 ( .A1(n6104), .A2(DATAI_29_), .ZN(n6409) );
  NAND2_X1 U3883 ( .A1(DATAI_6_), .A2(n4852), .ZN(n6367) );
  NAND2_X1 U3884 ( .A1(DATAI_7_), .A2(n4852), .ZN(n6374) );
  AND2_X1 U3885 ( .A1(n4662), .A2(n5062), .ZN(n4882) );
  AND2_X1 U3886 ( .A1(n6104), .A2(DATAI_31_), .ZN(n6419) );
  NAND2_X1 U3887 ( .A1(n4540), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6531) );
  NAND2_X1 U3888 ( .A1(n3962), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6537) );
  NOR2_X1 U3889 ( .A1(n6613), .A2(n5840), .ZN(n6629) );
  INV_X1 U3890 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6549) );
  INV_X1 U3891 ( .A(READY_N), .ZN(n6660) );
  NOR2_X1 U3892 ( .A1(n6565), .A2(n6668), .ZN(n6622) );
  INV_X1 U3893 ( .A(n6613), .ZN(n6668) );
  NAND2_X1 U3894 ( .A1(n2957), .A2(n4228), .ZN(n4229) );
  OAI21_X1 U3895 ( .B1(n5466), .B2(n5899), .A(n3008), .ZN(n3043) );
  INV_X1 U3896 ( .A(n5138), .ZN(n4496) );
  OAI21_X1 U3897 ( .B1(n5652), .B2(n5433), .A(n4493), .ZN(n4494) );
  OAI21_X1 U3898 ( .B1(n5175), .B2(n5594), .A(n5174), .ZN(n5176) );
  AOI21_X1 U3899 ( .B1(n5494), .B2(n6105), .A(n5493), .ZN(n5495) );
  NAND2_X1 U3900 ( .A1(n5138), .A2(n6104), .ZN(n4482) );
  OAI21_X1 U3901 ( .B1(n5669), .B2(n6100), .A(n4447), .ZN(U2962) );
  OAI211_X1 U3902 ( .C1(n5196), .C2(n6149), .A(n5134), .B(n5133), .ZN(n5135)
         );
  AND2_X1 U3903 ( .A1(n3550), .A2(n2997), .ZN(n2993) );
  OR2_X1 U3904 ( .A1(n5241), .A2(n3857), .ZN(n2994) );
  NAND2_X1 U3905 ( .A1(n2979), .A2(n3649), .ZN(n5299) );
  NAND2_X1 U3906 ( .A1(n4170), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n2995)
         );
  NAND2_X1 U3907 ( .A1(n4488), .A2(n5152), .ZN(n5151) );
  INV_X2 U3908 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n4802) );
  NAND2_X1 U3909 ( .A1(n4587), .A2(n4589), .ZN(n4588) );
  AND2_X1 U3910 ( .A1(n3081), .A2(n5253), .ZN(n2996) );
  AND2_X1 U3911 ( .A1(n3035), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n2997)
         );
  AND2_X1 U3912 ( .A1(n3091), .A2(n3549), .ZN(n2998) );
  AND2_X1 U3913 ( .A1(n3032), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n2999)
         );
  NAND2_X2 U3914 ( .A1(n4087), .A2(n5269), .ZN(n4016) );
  AND2_X1 U3915 ( .A1(n2979), .A2(n3101), .ZN(n5284) );
  AND2_X1 U3916 ( .A1(n5007), .A2(n5008), .ZN(n3000) );
  AND2_X1 U3917 ( .A1(n2979), .A2(n3100), .ZN(n4452) );
  AND4_X1 U3918 ( .A1(n3151), .A2(n3150), .A3(n3149), .A4(n3148), .ZN(n3001)
         );
  NAND2_X1 U3919 ( .A1(n5490), .A2(n3067), .ZN(n3002) );
  AND2_X1 U3920 ( .A1(n4018), .A2(n4589), .ZN(n3003) );
  XNOR2_X1 U3921 ( .A(n4200), .B(n4199), .ZN(n5192) );
  INV_X1 U3922 ( .A(n4681), .ZN(n4250) );
  OR2_X1 U3923 ( .A1(n5150), .A2(n4098), .ZN(n3005) );
  OR2_X1 U3924 ( .A1(n3253), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3006)
         );
  OR2_X1 U3925 ( .A1(n5196), .A2(n5968), .ZN(n3007) );
  NOR2_X1 U3926 ( .A1(n5320), .A2(n3044), .ZN(n3008) );
  OR2_X1 U3927 ( .A1(n5587), .A2(n4195), .ZN(n3009) );
  OR2_X1 U3928 ( .A1(n5151), .A2(n5214), .ZN(n3010) );
  OR2_X1 U3929 ( .A1(n3244), .A2(n2990), .ZN(n4104) );
  INV_X1 U3930 ( .A(n4104), .ZN(n3227) );
  AND2_X1 U3931 ( .A1(n3067), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3011)
         );
  AND3_X1 U3932 ( .A1(n3003), .A2(n4587), .A3(n3080), .ZN(n4744) );
  AND2_X1 U3933 ( .A1(n5007), .A2(n3091), .ZN(n3012) );
  AND2_X1 U3934 ( .A1(n4744), .A2(n4889), .ZN(n4888) );
  INV_X1 U3935 ( .A(n5200), .ZN(n3098) );
  NAND2_X1 U3936 ( .A1(n3003), .A2(n4587), .ZN(n4628) );
  AND2_X1 U3937 ( .A1(n5975), .A2(STATE2_REG_1__SCAN_IN), .ZN(n3013) );
  NAND2_X1 U3938 ( .A1(n3082), .A2(n4029), .ZN(n5012) );
  NOR2_X1 U3939 ( .A1(n5229), .A2(n5228), .ZN(n3014) );
  NAND2_X1 U3940 ( .A1(n3627), .A2(n3039), .ZN(n3015) );
  AND2_X1 U3941 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        STATE2_REG_0__SCAN_IN), .ZN(n3016) );
  INV_X1 U3942 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6530) );
  NAND2_X1 U3943 ( .A1(n5027), .A2(n5042), .ZN(n5041) );
  INV_X1 U3944 ( .A(n5283), .ZN(n4058) );
  INV_X1 U3945 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5345) );
  INV_X1 U3946 ( .A(n5312), .ZN(n3649) );
  OR2_X1 U3947 ( .A1(n5587), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3017)
         );
  AND2_X1 U3948 ( .A1(n5359), .A2(n5351), .ZN(n3018) );
  AND2_X1 U3949 ( .A1(n5118), .A2(n4078), .ZN(n4489) );
  AND2_X1 U3950 ( .A1(n4489), .A2(n4490), .ZN(n4488) );
  AND2_X1 U3951 ( .A1(n4455), .A2(n3100), .ZN(n3019) );
  AND2_X1 U3952 ( .A1(n2996), .A2(n3014), .ZN(n3020) );
  AND2_X1 U3953 ( .A1(n4029), .A2(n4033), .ZN(n3021) );
  AND2_X1 U3954 ( .A1(STATE2_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3022) );
  AND2_X1 U3955 ( .A1(n3550), .A2(n3035), .ZN(n3023) );
  INV_X1 U3956 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3040) );
  AND2_X1 U3957 ( .A1(n4602), .A2(n4603), .ZN(n4587) );
  AND2_X1 U3958 ( .A1(n3047), .A2(n3046), .ZN(n3024) );
  INV_X1 U3959 ( .A(n5038), .ZN(n3549) );
  AOI21_X1 U3960 ( .B1(n4575), .B2(n4483), .A(n4007), .ZN(n4602) );
  INV_X1 U3961 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3049) );
  INV_X1 U3962 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3037) );
  INV_X1 U3963 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3033) );
  INV_X1 U3964 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3041) );
  INV_X1 U3965 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3064) );
  NAND2_X1 U3966 ( .A1(n2987), .A2(n3026), .ZN(n3025) );
  NAND3_X1 U3967 ( .A1(n3025), .A2(n4105), .A3(n4260), .ZN(n3237) );
  NAND2_X1 U3968 ( .A1(n3359), .A2(n3027), .ZN(n3476) );
  NOR2_X2 U3969 ( .A1(n3370), .A2(n3368), .ZN(n3359) );
  NAND2_X2 U3970 ( .A1(n3052), .A2(n5568), .ZN(n5750) );
  NAND3_X1 U3971 ( .A1(n3055), .A2(n3054), .A3(n3053), .ZN(n5022) );
  NAND2_X1 U3972 ( .A1(n4177), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3063)
         );
  INV_X1 U3973 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3034) );
  INV_X1 U3974 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3042) );
  OR2_X1 U3975 ( .A1(n5319), .A2(n3043), .ZN(U2810) );
  AOI21_X2 U3976 ( .B1(n5750), .B2(n5751), .A(n3075), .ZN(n5550) );
  NOR2_X1 U3977 ( .A1(n4186), .A2(n3057), .ZN(n3056) );
  INV_X1 U3978 ( .A(n3063), .ZN(n3057) );
  OAI21_X1 U3979 ( .B1(n4926), .B2(n4927), .A(n3063), .ZN(n5051) );
  AND2_X1 U3980 ( .A1(n3060), .A2(n2995), .ZN(n4926) );
  NAND3_X1 U3981 ( .A1(n3062), .A2(n3061), .A3(n4887), .ZN(n3060) );
  NAND2_X1 U3982 ( .A1(n3065), .A2(n4003), .ZN(n3229) );
  AOI21_X1 U3983 ( .B1(n4138), .B2(n4137), .A(n3065), .ZN(n4139) );
  NAND2_X1 U3984 ( .A1(n3252), .A2(n3022), .ZN(n3256) );
  NAND2_X1 U3985 ( .A1(n5490), .A2(n3109), .ZN(n5489) );
  NAND2_X1 U3986 ( .A1(n5490), .A2(n3011), .ZN(n3071) );
  NAND2_X1 U3987 ( .A1(n5164), .A2(n4197), .ZN(n3069) );
  AOI21_X1 U3988 ( .B1(n5750), .B2(n3074), .A(n3072), .ZN(n4475) );
  AND2_X1 U3989 ( .A1(n3078), .A2(n4196), .ZN(n3074) );
  NAND2_X1 U3990 ( .A1(n3082), .A2(n3021), .ZN(n5011) );
  NAND2_X1 U3991 ( .A1(n5007), .A2(n2998), .ZN(n5039) );
  NAND2_X1 U3992 ( .A1(n3093), .A2(n3351), .ZN(n3457) );
  NAND2_X1 U3993 ( .A1(n3096), .A2(n3094), .ZN(n3099) );
  AND2_X1 U3994 ( .A1(n3096), .A2(n3097), .ZN(n4200) );
  NAND2_X1 U3995 ( .A1(n2979), .A2(n3019), .ZN(n4453) );
  INV_X1 U3996 ( .A(n5497), .ZN(n5498) );
  NOR2_X1 U3997 ( .A1(n5528), .A2(n5527), .ZN(n5526) );
  OAI21_X1 U3998 ( .B1(n5192), .B2(n5599), .A(n4470), .ZN(n4471) );
  OAI21_X1 U3999 ( .B1(n5192), .B2(n5899), .A(n4001), .ZN(n4002) );
  AOI22_X1 U4000 ( .A1(n3280), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3206), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3139) );
  AOI22_X1 U4001 ( .A1(n3379), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3386), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3143) );
  AND2_X1 U4002 ( .A1(n4164), .A2(n4163), .ZN(n4181) );
  OR2_X1 U4003 ( .A1(n4432), .A2(n4431), .ZN(n3102) );
  INV_X1 U4004 ( .A(n6138), .ZN(n6149) );
  INV_X2 U4005 ( .A(n5989), .ZN(n5477) );
  AND2_X1 U4006 ( .A1(n5991), .A2(n4110), .ZN(n5989) );
  AND2_X1 U4007 ( .A1(n3457), .A2(n3353), .ZN(n4115) );
  NOR2_X1 U4008 ( .A1(n4435), .A2(n4098), .ZN(n3104) );
  OR2_X1 U4009 ( .A1(n4442), .A2(n4441), .ZN(n3105) );
  AND2_X1 U4010 ( .A1(n3823), .A2(n3822), .ZN(n4435) );
  NOR2_X1 U4011 ( .A1(n4184), .A2(n4183), .ZN(n3107) );
  INV_X1 U4012 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4232) );
  INV_X1 U4013 ( .A(n5499), .ZN(n4462) );
  NOR2_X1 U4014 ( .A1(n4888), .A2(n4890), .ZN(n3108) );
  AND2_X1 U4015 ( .A1(n5500), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3109)
         );
  INV_X1 U4016 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6509) );
  AND2_X1 U4017 ( .A1(n4439), .A2(n4438), .ZN(n3110) );
  AND2_X1 U4018 ( .A1(n4113), .A2(n4112), .ZN(n3111) );
  AND2_X1 U4019 ( .A1(n4458), .A2(n4457), .ZN(n3112) );
  NOR2_X1 U4020 ( .A1(n4661), .A2(n4802), .ZN(n3481) );
  NAND2_X1 U4021 ( .A1(n5232), .A2(n5234), .ZN(n5233) );
  OR2_X1 U4022 ( .A1(n3287), .A2(n3286), .ZN(n4134) );
  AOI22_X1 U4023 ( .A1(n3385), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3125) );
  NOR2_X1 U4024 ( .A1(n4709), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3943)
         );
  BUF_X1 U4025 ( .A(n3208), .Z(n3838) );
  NAND2_X1 U4026 ( .A1(n4674), .A2(n3236), .ZN(n3306) );
  AOI21_X1 U4027 ( .B1(n3945), .B2(n3944), .A(n3943), .ZN(n3950) );
  INV_X1 U4028 ( .A(n5873), .ZN(n3568) );
  NOR2_X1 U4029 ( .A1(n4179), .A2(n6530), .ZN(n4180) );
  OR2_X1 U4030 ( .A1(n3469), .A2(n3468), .ZN(n4172) );
  INV_X1 U4031 ( .A(n3930), .ZN(n3947) );
  AND2_X1 U4032 ( .A1(n3950), .A2(n3946), .ZN(n3966) );
  INV_X1 U4033 ( .A(n3254), .ZN(n3255) );
  INV_X1 U4035 ( .A(n3481), .ZN(n3455) );
  INV_X1 U4036 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4440) );
  INV_X1 U4037 ( .A(n3248), .ZN(n3230) );
  AND2_X1 U4038 ( .A1(n4045), .A2(n4044), .ZN(n5351) );
  OR2_X1 U4039 ( .A1(n4277), .A2(n2959), .ZN(n4706) );
  NAND2_X1 U4040 ( .A1(n3418), .A2(n6530), .ZN(n3412) );
  OR4_X1 U4041 ( .A1(n3969), .A2(n3968), .A3(n3967), .A4(n3966), .ZN(n3970) );
  OR2_X1 U4042 ( .A1(n5220), .A2(n3980), .ZN(n5211) );
  OR2_X1 U4043 ( .A1(n5272), .A2(n3989), .ZN(n5121) );
  NAND2_X1 U4044 ( .A1(n3975), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n3976)
         );
  AND2_X1 U4045 ( .A1(n5429), .A2(n5323), .ZN(n4052) );
  NOR2_X1 U4046 ( .A1(n4524), .A2(n4279), .ZN(n4281) );
  INV_X1 U4047 ( .A(n3900), .ZN(n3872) );
  OR2_X1 U4048 ( .A1(n4548), .A2(n4700), .ZN(n4549) );
  INV_X1 U4049 ( .A(n3817), .ZN(n4098) );
  INV_X1 U4050 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3519) );
  OR2_X1 U4051 ( .A1(n5199), .A2(n4214), .ZN(n4217) );
  INV_X1 U4052 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4709) );
  AND2_X1 U4053 ( .A1(n6437), .A2(n6207), .ZN(n6235) );
  NAND2_X1 U4054 ( .A1(n3326), .A2(n3325), .ZN(n6436) );
  NAND2_X1 U4055 ( .A1(n3959), .A2(n3965), .ZN(n3960) );
  AOI21_X1 U4056 ( .B1(n4000), .B2(n4221), .A(n3999), .ZN(n4001) );
  AND2_X1 U4057 ( .A1(n4080), .A2(n4079), .ZN(n4490) );
  AND2_X1 U4058 ( .A1(n4061), .A2(n4060), .ZN(n5282) );
  AND2_X1 U4059 ( .A1(n4685), .A2(n4661), .ZN(n4265) );
  NOR2_X1 U4060 ( .A1(n5358), .A2(n5357), .ZN(n5356) );
  INV_X1 U4061 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4465) );
  AND2_X1 U4062 ( .A1(n5662), .A2(n4428), .ZN(n5636) );
  OR2_X1 U4063 ( .A1(n4548), .A2(n4252), .ZN(n4253) );
  OAI21_X1 U4064 ( .B1(n6663), .B2(n4735), .A(n6531), .ZN(n4659) );
  INV_X1 U4065 ( .A(n6309), .ZN(n6338) );
  INV_X1 U4066 ( .A(n6172), .ZN(n5793) );
  AND2_X1 U4067 ( .A1(n4729), .A2(n5793), .ZN(n6184) );
  OR2_X1 U4068 ( .A1(n6337), .A2(n5062), .ZN(n5114) );
  INV_X1 U4069 ( .A(n4652), .ZN(n5061) );
  NAND2_X1 U4070 ( .A1(n4662), .A2(n6307), .ZN(n4834) );
  NOR2_X1 U4071 ( .A1(n4208), .A2(n4725), .ZN(n3977) );
  AND2_X1 U4072 ( .A1(n5939), .A2(n5377), .ZN(n5904) );
  INV_X1 U4073 ( .A(n5918), .ZN(n5933) );
  AND2_X1 U4074 ( .A1(n5975), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5960) );
  INV_X1 U4075 ( .A(n5433), .ZN(n5979) );
  AND2_X1 U4076 ( .A1(n5991), .A2(n4111), .ZN(n5468) );
  NAND2_X1 U4077 ( .A1(n4583), .A2(n4582), .ZN(n5988) );
  INV_X1 U4078 ( .A(n5992), .ZN(n6001) );
  OR2_X1 U4079 ( .A1(n4548), .A2(n3963), .ZN(n4513) );
  INV_X1 U4080 ( .A(n6544), .ZN(n4203) );
  NAND2_X1 U4081 ( .A1(n5519), .A2(n6155), .ZN(n4303) );
  AND2_X1 U4082 ( .A1(n4292), .A2(n4261), .ZN(n6138) );
  INV_X1 U4083 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n3238) );
  INV_X1 U4084 ( .A(n6537), .ZN(n4545) );
  INV_X1 U4085 ( .A(n4918), .ZN(n6164) );
  INV_X1 U4086 ( .A(n4898), .ZN(n6166) );
  INV_X1 U4087 ( .A(n4940), .ZN(n6175) );
  OR2_X1 U4088 ( .A1(n6212), .A2(n6211), .ZN(n6230) );
  NOR2_X2 U4089 ( .A1(n6213), .A2(n5062), .ZN(n6266) );
  NOR2_X1 U4090 ( .A1(n4645), .A2(n6435), .ZN(n6308) );
  OR3_X1 U4091 ( .A1(n6316), .A2(n6315), .A3(n6314), .ZN(n6333) );
  OAI21_X1 U4092 ( .B1(n6345), .B2(n6344), .A(n6343), .ZN(n6371) );
  INV_X1 U4093 ( .A(n5114), .ZN(n6370) );
  OAI21_X1 U4094 ( .B1(n6389), .B2(n6386), .A(n6385), .ZN(n6421) );
  OR2_X1 U4095 ( .A1(n6441), .A2(n6440), .ZN(n6488) );
  INV_X1 U4096 ( .A(n5094), .ZN(n6458) );
  INV_X1 U4097 ( .A(n6374), .ZN(n6485) );
  AND2_X1 U4098 ( .A1(n6104), .A2(DATAI_19_), .ZN(n6460) );
  AND2_X1 U4099 ( .A1(n4803), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4973) );
  INV_X1 U4100 ( .A(n6463), .ZN(n6401) );
  INV_X1 U4101 ( .A(n6481), .ZN(n6413) );
  AND2_X1 U4102 ( .A1(n4725), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3962) );
  NOR2_X1 U4103 ( .A1(n4725), .A2(n4802), .ZN(n4735) );
  INV_X1 U4104 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6559) );
  INV_X1 U4105 ( .A(n6624), .ZN(n6618) );
  NAND2_X1 U4106 ( .A1(n4513), .A2(n5802), .ZN(n6658) );
  INV_X1 U4107 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6432) );
  NAND2_X1 U4108 ( .A1(n6559), .A2(STATE_REG_1__SCAN_IN), .ZN(n6657) );
  INV_X1 U4109 ( .A(n4002), .ZN(n4096) );
  INV_X1 U4110 ( .A(n5927), .ZN(n5968) );
  NAND2_X1 U4111 ( .A1(n5975), .A2(n3977), .ZN(n5899) );
  OR2_X1 U4112 ( .A1(n6658), .A2(n3974), .ZN(n5975) );
  INV_X1 U4113 ( .A(n4494), .ZN(n4495) );
  AND2_X2 U4114 ( .A1(n4487), .A2(n4545), .ZN(n5987) );
  NAND2_X1 U4115 ( .A1(n6083), .A2(n4109), .ZN(n5991) );
  NAND2_X1 U4116 ( .A1(n6022), .A2(n4248), .ZN(n5992) );
  INV_X1 U4117 ( .A(n6022), .ZN(n6035) );
  INV_X1 U4118 ( .A(n6089), .ZN(n6037) );
  OR2_X1 U4119 ( .A1(n4513), .A2(n4101), .ZN(n6083) );
  AND2_X1 U4120 ( .A1(n4480), .A2(n4479), .ZN(n4481) );
  NAND2_X1 U4121 ( .A1(n6100), .A2(n4205), .ZN(n6112) );
  OR2_X2 U4122 ( .A1(n4548), .A2(n6517), .ZN(n6100) );
  NAND2_X1 U4123 ( .A1(n4303), .A2(n4302), .ZN(n4420) );
  INV_X1 U4124 ( .A(n5816), .ZN(n6119) );
  NAND2_X1 U4125 ( .A1(n4292), .A2(n4259), .ZN(n6142) );
  INV_X1 U4126 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6378) );
  OR2_X1 U4127 ( .A1(n4766), .A2(n6307), .ZN(n4918) );
  AOI22_X1 U4128 ( .A1(n6179), .A2(n6182), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6178), .ZN(n6204) );
  INV_X1 U4129 ( .A(n6209), .ZN(n6233) );
  AOI22_X1 U4130 ( .A1(n6239), .A2(n6237), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6242), .ZN(n6262) );
  INV_X1 U4131 ( .A(n6276), .ZN(n6302) );
  NAND2_X1 U4132 ( .A1(n6277), .A2(n6376), .ZN(n6336) );
  INV_X1 U4133 ( .A(n6340), .ZN(n6375) );
  AOI22_X1 U4134 ( .A1(n5071), .A2(n6383), .B1(n5066), .B2(n5065), .ZN(n5117)
         );
  INV_X1 U4135 ( .A(n6379), .ZN(n6445) );
  INV_X1 U4136 ( .A(n6352), .ZN(n6457) );
  NAND2_X1 U4137 ( .A1(n6377), .A2(n6376), .ZN(n6491) );
  NAND2_X1 U4138 ( .A1(n4777), .A2(n6307), .ZN(n4879) );
  NAND2_X1 U4139 ( .A1(DATAI_0_), .A2(n4852), .ZN(n6348) );
  NAND2_X1 U4140 ( .A1(DATAI_5_), .A2(n4852), .ZN(n6364) );
  NOR2_X1 U4141 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6663) );
  INV_X1 U4142 ( .A(n6629), .ZN(n6548) );
  INV_X1 U4143 ( .A(n6657), .ZN(n6613) );
  INV_X1 U4144 ( .A(n6622), .ZN(n6620) );
  OAI21_X1 U4145 ( .B1(n4496), .B2(n5438), .A(n4495), .ZN(U2834) );
  NAND2_X1 U4146 ( .A1(n4114), .A2(n3111), .ZN(U2866) );
  NAND2_X1 U4147 ( .A1(n4482), .A2(n4481), .ZN(U2961) );
  NOR2_X4 U4148 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4526) );
  AND2_X4 U4149 ( .A1(n4526), .A2(n3120), .ZN(n3207) );
  AND2_X4 U4150 ( .A1(n4529), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4532)
         );
  NOR2_X4 U4151 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3121) );
  AND2_X4 U4152 ( .A1(n4532), .A2(n3121), .ZN(n3208) );
  AOI22_X1 U4153 ( .A1(n3207), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3208), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3117) );
  INV_X1 U4154 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3113) );
  AND2_X4 U4155 ( .A1(n3113), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3118)
         );
  AND2_X4 U4156 ( .A1(n3120), .A2(n3119), .ZN(n3395) );
  AND2_X4 U4157 ( .A1(n4526), .A2(n3121), .ZN(n3281) );
  AOI22_X1 U4158 ( .A1(n3395), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3115) );
  AND2_X4 U4159 ( .A1(n3118), .A2(n4526), .ZN(n3206) );
  AOI22_X1 U4160 ( .A1(n3280), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3206), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3114) );
  AND2_X4 U4161 ( .A1(n4532), .A2(n3118), .ZN(n3385) );
  AOI22_X1 U4162 ( .A1(n3379), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3386), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3124) );
  AND2_X4 U4163 ( .A1(n3119), .A2(n3121), .ZN(n3274) );
  AOI22_X1 U4164 ( .A1(n3274), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3217), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3123) );
  AOI22_X1 U4165 ( .A1(n3396), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3179), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3122) );
  NAND2_X2 U4166 ( .A1(n3127), .A2(n3126), .ZN(n3178) );
  AOI22_X1 U4167 ( .A1(n3279), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3201), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3131) );
  AOI22_X1 U4168 ( .A1(n3379), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3386), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3130) );
  AOI22_X1 U4169 ( .A1(n3385), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3206), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3129) );
  AOI22_X1 U4170 ( .A1(n3179), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3217), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3128) );
  AOI22_X1 U4171 ( .A1(n3396), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3274), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3135) );
  AOI22_X1 U4172 ( .A1(n3207), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3280), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3134) );
  AOI22_X1 U4173 ( .A1(n3208), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3133) );
  AOI22_X1 U4175 ( .A1(n3207), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3208), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3141) );
  AOI22_X1 U4176 ( .A1(n3279), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3201), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3140) );
  AOI22_X1 U4177 ( .A1(n3395), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3138) );
  AOI22_X1 U4178 ( .A1(n3385), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3145) );
  AOI22_X1 U4179 ( .A1(n3396), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3179), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3144) );
  AOI22_X1 U4180 ( .A1(n3274), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3217), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3142) );
  NAND2_X1 U4181 ( .A1(n2959), .A2(n3178), .ZN(n3156) );
  AOI22_X1 U4182 ( .A1(n3379), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3150) );
  AOI22_X1 U4183 ( .A1(n3395), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3149) );
  AOI22_X1 U4184 ( .A1(n3396), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3217), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3148) );
  AOI22_X1 U4185 ( .A1(n3207), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3206), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3155) );
  AOI22_X1 U4186 ( .A1(n3279), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3280), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3154) );
  AOI22_X1 U4187 ( .A1(n3385), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3386), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3153) );
  AOI22_X1 U4188 ( .A1(n3274), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3179), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3152) );
  NAND2_X1 U4189 ( .A1(n3157), .A2(n3241), .ZN(n3265) );
  AOI22_X1 U4190 ( .A1(n3395), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3161) );
  AOI22_X1 U4191 ( .A1(n3385), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3160) );
  AOI22_X1 U4192 ( .A1(n3201), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3206), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3159) );
  AOI22_X1 U4193 ( .A1(n3274), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3386), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3158) );
  AND4_X2 U4194 ( .A1(n3161), .A2(n3160), .A3(n3159), .A4(n3158), .ZN(n3167)
         );
  AOI22_X1 U4195 ( .A1(n3279), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3280), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3165) );
  AOI22_X1 U4196 ( .A1(n3208), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3164) );
  AOI22_X1 U4197 ( .A1(n3396), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3179), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3163) );
  AOI22_X1 U4198 ( .A1(n3379), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3217), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3162) );
  AND4_X2 U4199 ( .A1(n3165), .A2(n3164), .A3(n3163), .A4(n3162), .ZN(n3166)
         );
  NAND2_X4 U4200 ( .A1(n3167), .A2(n3166), .ZN(n4681) );
  AOI22_X1 U4201 ( .A1(n3279), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3201), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3171) );
  AOI22_X1 U4202 ( .A1(n3207), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3208), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3170) );
  AOI22_X1 U4203 ( .A1(n3280), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3206), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3169) );
  AOI22_X1 U4204 ( .A1(n3395), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3168) );
  NAND4_X1 U4205 ( .A1(n3171), .A2(n3170), .A3(n3169), .A4(n3168), .ZN(n3177)
         );
  AOI22_X1 U4206 ( .A1(n3385), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3175) );
  AOI22_X1 U4207 ( .A1(n3379), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3386), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3174) );
  AOI22_X1 U4208 ( .A1(n3396), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3179), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3173) );
  AOI22_X1 U4209 ( .A1(n3274), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3217), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3172) );
  NAND4_X1 U4210 ( .A1(n3175), .A2(n3174), .A3(n3173), .A4(n3172), .ZN(n3176)
         );
  OR2_X2 U4211 ( .A1(n3177), .A2(n3176), .ZN(n3243) );
  NAND2_X1 U4212 ( .A1(n4250), .A2(n3243), .ZN(n4262) );
  NAND2_X1 U4213 ( .A1(n3396), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3183) );
  NAND2_X1 U4214 ( .A1(n3274), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3182) );
  NAND2_X1 U4215 ( .A1(n3217), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3181)
         );
  NAND2_X1 U4216 ( .A1(n3179), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3180) );
  NAND2_X1 U4217 ( .A1(n3201), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3187)
         );
  NAND2_X1 U4218 ( .A1(n3279), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3186) );
  NAND2_X1 U4219 ( .A1(n3206), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3185) );
  NAND2_X1 U4220 ( .A1(n3280), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3184) );
  NAND2_X1 U4221 ( .A1(n3385), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3192) );
  NAND2_X1 U4222 ( .A1(n3188), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3191)
         );
  NAND2_X1 U4223 ( .A1(n3379), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3190)
         );
  NAND2_X1 U4224 ( .A1(n3386), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3189)
         );
  NAND2_X1 U4225 ( .A1(n3208), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3196) );
  NAND2_X1 U4226 ( .A1(n3395), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3195)
         );
  NAND2_X1 U4227 ( .A1(n3207), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3194) );
  NAND2_X1 U4228 ( .A1(n3281), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3193) );
  NAND2_X1 U4229 ( .A1(n3201), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3205)
         );
  NAND2_X1 U4230 ( .A1(n3395), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3204)
         );
  NAND2_X1 U4231 ( .A1(n3279), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3203) );
  NAND2_X1 U4232 ( .A1(n3281), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3202) );
  NAND2_X1 U4233 ( .A1(n3207), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3211) );
  NAND2_X1 U4234 ( .A1(n3208), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3210) );
  NAND2_X1 U4235 ( .A1(n3280), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3209) );
  NAND3_X1 U4236 ( .A1(n3211), .A2(n3210), .A3(n3209), .ZN(n3212) );
  NAND2_X1 U4237 ( .A1(n3379), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3216)
         );
  NAND2_X1 U4238 ( .A1(n3396), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3215) );
  NAND2_X1 U4239 ( .A1(n3385), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3214) );
  NAND2_X1 U4240 ( .A1(n3179), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3213) );
  NAND2_X1 U4241 ( .A1(n3188), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3221)
         );
  NAND2_X1 U4242 ( .A1(n3274), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3220) );
  NAND2_X1 U4243 ( .A1(n3386), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3219)
         );
  NAND2_X1 U4244 ( .A1(n3217), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3218)
         );
  XNOR2_X1 U4245 ( .A(n6549), .B(STATE_REG_2__SCAN_IN), .ZN(n3978) );
  AND2_X2 U4246 ( .A1(n3227), .A2(n3226), .ZN(n4521) );
  NAND2_X1 U4247 ( .A1(n4521), .A2(n4265), .ZN(n4260) );
  NAND2_X1 U4249 ( .A1(n3229), .A2(n3228), .ZN(n3235) );
  NAND2_X1 U4250 ( .A1(n3904), .A2(n4681), .ZN(n3234) );
  INV_X1 U4251 ( .A(n3258), .ZN(n3231) );
  NOR2_X1 U4252 ( .A1(n3232), .A2(n3231), .ZN(n3233) );
  NAND3_X2 U4253 ( .A1(n3235), .A2(n3234), .A3(n3233), .ZN(n3264) );
  INV_X2 U4254 ( .A(n3244), .ZN(n3242) );
  XNOR2_X1 U4255 ( .A(n6504), .B(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6305)
         );
  NAND2_X1 U4256 ( .A1(n3303), .A2(n6305), .ZN(n3240) );
  INV_X1 U4257 ( .A(n3962), .ZN(n3302) );
  NAND2_X1 U4258 ( .A1(n3302), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3239) );
  NAND2_X1 U4259 ( .A1(n3240), .A2(n3239), .ZN(n3253) );
  NAND2_X1 U4260 ( .A1(n3264), .A2(n4669), .ZN(n3251) );
  INV_X2 U4261 ( .A(n4214), .ZN(n3245) );
  INV_X1 U4262 ( .A(n3249), .ZN(n3250) );
  NAND4_X1 U4263 ( .A1(n3251), .A2(n3263), .A3(n3250), .A4(n4102), .ZN(n3252)
         );
  NAND2_X1 U4264 ( .A1(n3299), .A2(n3319), .ZN(n3273) );
  MUX2_X1 U4265 ( .A(n3302), .B(n3303), .S(n6378), .Z(n3254) );
  NAND2_X1 U4266 ( .A1(n3257), .A2(n3258), .ZN(n4274) );
  INV_X1 U4267 ( .A(n4527), .ZN(n6496) );
  INV_X1 U4268 ( .A(n4484), .ZN(n3259) );
  NOR2_X1 U4269 ( .A1(n3259), .A2(n4248), .ZN(n3260) );
  NAND2_X1 U4270 ( .A1(n6496), .A2(n3260), .ZN(n4277) );
  NAND2_X1 U4271 ( .A1(n3228), .A2(n3243), .ZN(n3261) );
  OR2_X1 U4272 ( .A1(n6647), .A2(n6530), .ZN(n6538) );
  OAI211_X1 U4273 ( .C1(n4669), .C2(n4681), .A(n4273), .B(n4104), .ZN(n4268)
         );
  AND3_X1 U4274 ( .A1(n4277), .A2(n3262), .A3(n4268), .ZN(n3271) );
  NAND2_X1 U4275 ( .A1(n3264), .A2(n3227), .ZN(n4270) );
  NAND2_X1 U4277 ( .A1(n3267), .A2(n3243), .ZN(n3269) );
  OAI21_X1 U4278 ( .B1(n3266), .B2(n3269), .A(n3268), .ZN(n3270) );
  NAND4_X1 U4279 ( .A1(n3271), .A2(n3263), .A3(n4270), .A4(n3270), .ZN(n3291)
         );
  INV_X1 U4280 ( .A(n3298), .ZN(n3272) );
  XNOR2_X1 U4281 ( .A(n3273), .B(n3272), .ZN(n4519) );
  NAND2_X1 U4282 ( .A1(n4519), .A2(n6530), .ZN(n3290) );
  AOI22_X1 U4283 ( .A1(n3378), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3208), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3278) );
  AOI22_X1 U4284 ( .A1(n3779), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3884), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3277) );
  BUF_X1 U4285 ( .A(n3274), .Z(n3441) );
  AOI22_X1 U4286 ( .A1(n3387), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3441), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3276) );
  AOI22_X1 U4287 ( .A1(n3860), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3206), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3275) );
  NAND4_X1 U4288 ( .A1(n3278), .A2(n3277), .A3(n3276), .A4(n3275), .ZN(n3287)
         );
  INV_X1 U4289 ( .A(n3280), .ZN(n4708) );
  AOI22_X1 U4290 ( .A1(n3394), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3280), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3285) );
  AOI22_X1 U4291 ( .A1(n3207), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3284) );
  AOI22_X1 U4292 ( .A1(n3397), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3843), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3283) );
  AOI22_X1 U4293 ( .A1(n3380), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3885), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3282) );
  NAND4_X1 U4294 ( .A1(n3285), .A2(n3284), .A3(n3283), .A4(n3282), .ZN(n3286)
         );
  AND2_X1 U4295 ( .A1(n4256), .A2(n4134), .ZN(n3288) );
  NAND2_X1 U4296 ( .A1(n3290), .A2(n3289), .ZN(n3371) );
  INV_X1 U4297 ( .A(n3291), .ZN(n3292) );
  XNOR2_X1 U4298 ( .A(n3293), .B(n3292), .ZN(n3418) );
  NAND2_X1 U4299 ( .A1(n4669), .A2(n4134), .ZN(n3295) );
  NAND2_X1 U4300 ( .A1(n3295), .A2(n4674), .ZN(n3296) );
  AOI22_X1 U4301 ( .A1(n3930), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3296), 
        .B2(STATE2_REG_0__SCAN_IN), .ZN(n3297) );
  NAND2_X1 U4302 ( .A1(n3371), .A2(n3372), .ZN(n3370) );
  NAND2_X1 U4303 ( .A1(n3320), .A2(n3319), .ZN(n3305) );
  NAND2_X1 U4304 ( .A1(n6306), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5067) );
  MUX2_X1 U4305 ( .A(n5067), .B(n6306), .S(n6378), .Z(n3301) );
  INV_X1 U4306 ( .A(n6206), .ZN(n3300) );
  NAND2_X1 U4307 ( .A1(n3301), .A2(n3300), .ZN(n4803) );
  AOI22_X1 U4308 ( .A1(n4803), .A2(n3303), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3302), .ZN(n3304) );
  XNOR2_X1 U4309 ( .A(n3305), .B(n3318), .ZN(n4646) );
  INV_X1 U4310 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4827) );
  AOI22_X1 U4311 ( .A1(n3860), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3280), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3310) );
  AOI22_X1 U4312 ( .A1(n3274), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3884), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3309) );
  AOI22_X1 U4313 ( .A1(n3378), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3206), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3308) );
  AOI22_X1 U4314 ( .A1(n3387), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3885), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3307) );
  NAND4_X1 U4315 ( .A1(n3310), .A2(n3309), .A3(n3308), .A4(n3307), .ZN(n3316)
         );
  AOI22_X1 U4316 ( .A1(n3394), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3314) );
  AOI22_X1 U4317 ( .A1(n3838), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3787), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3313) );
  AOI22_X1 U4318 ( .A1(n3397), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3843), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3312) );
  AOI22_X1 U4319 ( .A1(n3779), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3311) );
  NAND4_X1 U4320 ( .A1(n3314), .A2(n3313), .A3(n3312), .A4(n3311), .ZN(n3315)
         );
  OAI22_X1 U4321 ( .A1(n4827), .A2(n3947), .B1(n3923), .B2(n4116), .ZN(n3317)
         );
  NAND2_X1 U4322 ( .A1(n3321), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3326) );
  NAND3_X1 U4323 ( .A1(n6509), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6279) );
  INV_X1 U4324 ( .A(n6279), .ZN(n3322) );
  NAND2_X1 U4325 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3322), .ZN(n6273) );
  NAND2_X1 U4326 ( .A1(n6509), .A2(n6273), .ZN(n3323) );
  NAND3_X1 U4327 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4850) );
  INV_X1 U4328 ( .A(n4850), .ZN(n4649) );
  NAND2_X1 U4329 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4649), .ZN(n4691) );
  NAND2_X1 U4330 ( .A1(n3323), .A2(n4691), .ZN(n6304) );
  OAI22_X1 U4331 ( .A1(n4204), .A2(n6304), .B1(n3962), .B2(n6509), .ZN(n3324)
         );
  INV_X1 U4332 ( .A(n3324), .ZN(n3325) );
  XNOR2_X2 U4333 ( .A(n4722), .B(n6436), .ZN(n4645) );
  NAND2_X1 U4334 ( .A1(n4645), .A2(n6530), .ZN(n3338) );
  AOI22_X1 U4335 ( .A1(n3394), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3330) );
  AOI22_X1 U4336 ( .A1(n3879), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3838), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3329) );
  INV_X1 U4337 ( .A(n4708), .ZN(n3459) );
  AOI22_X1 U4338 ( .A1(n3459), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3206), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3328) );
  AOI22_X1 U4339 ( .A1(n3378), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3787), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3327) );
  NAND4_X1 U4340 ( .A1(n3330), .A2(n3329), .A3(n3328), .A4(n3327), .ZN(n3336)
         );
  AOI22_X1 U4341 ( .A1(n3397), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3884), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3334) );
  AOI22_X1 U4342 ( .A1(n3779), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3843), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3333) );
  AOI22_X1 U4343 ( .A1(n3387), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3332) );
  AOI22_X1 U4344 ( .A1(n3441), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3885), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3331) );
  NAND4_X1 U4345 ( .A1(n3334), .A2(n3333), .A3(n3332), .A4(n3331), .ZN(n3335)
         );
  AOI22_X1 U4346 ( .A1(INSTQUEUE_REG_0__3__SCAN_IN), .A2(n3930), .B1(n3955), 
        .B2(n4146), .ZN(n3337) );
  NAND2_X1 U4347 ( .A1(n3930), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3350) );
  AOI22_X1 U4348 ( .A1(n3394), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3342) );
  AOI22_X1 U4349 ( .A1(n3397), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3441), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3341) );
  AOI22_X1 U4350 ( .A1(n3459), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3787), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3340) );
  AOI22_X1 U4351 ( .A1(n3387), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3339) );
  NAND4_X1 U4352 ( .A1(n3342), .A2(n3341), .A3(n3340), .A4(n3339), .ZN(n3348)
         );
  AOI22_X1 U4353 ( .A1(n3378), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3838), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3346) );
  AOI22_X1 U4354 ( .A1(n3879), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3345) );
  AOI22_X1 U4355 ( .A1(n3884), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3843), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3344) );
  AOI22_X1 U4356 ( .A1(n3779), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3885), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3343) );
  NAND4_X1 U4357 ( .A1(n3346), .A2(n3345), .A3(n3344), .A4(n3343), .ZN(n3347)
         );
  NAND2_X1 U4358 ( .A1(n3955), .A2(n4154), .ZN(n3349) );
  NAND2_X1 U4359 ( .A1(n3360), .A2(n3352), .ZN(n3353) );
  AND2_X1 U4360 ( .A1(n4265), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3419) );
  INV_X1 U4361 ( .A(n3419), .ZN(n3429) );
  INV_X1 U4362 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4723) );
  NAND2_X1 U4363 ( .A1(n4802), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3355)
         );
  NAND2_X1 U4364 ( .A1(n3726), .A2(EAX_REG_4__SCAN_IN), .ZN(n3354) );
  OAI211_X1 U4365 ( .C1(n3429), .C2(n4723), .A(n3355), .B(n3354), .ZN(n3357)
         );
  INV_X1 U4366 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3356) );
  XNOR2_X1 U4367 ( .A(n3451), .B(n3356), .ZN(n5934) );
  MUX2_X1 U4368 ( .A(n3357), .B(n5934), .S(n3903), .Z(n3358) );
  AOI21_X1 U4369 ( .B1(n4115), .B2(n3584), .A(n3358), .ZN(n4750) );
  INV_X1 U4370 ( .A(n4750), .ZN(n3436) );
  OAI21_X1 U4371 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3362), .A(n3451), 
        .ZN(n5946) );
  AOI22_X1 U4372 ( .A1(n3903), .A2(n5946), .B1(n4201), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3364) );
  NAND2_X1 U4373 ( .A1(n3726), .A2(EAX_REG_3__SCAN_IN), .ZN(n3363) );
  OAI211_X1 U4374 ( .C1(n3429), .C2(n4709), .A(n3364), .B(n3363), .ZN(n3365)
         );
  INV_X1 U4375 ( .A(n3365), .ZN(n3366) );
  INV_X1 U4376 ( .A(n3368), .ZN(n3369) );
  XNOR2_X1 U4377 ( .A(n3370), .B(n3369), .ZN(n4653) );
  AOI21_X1 U4378 ( .B1(n4653), .B2(n3584), .A(n4201), .ZN(n3430) );
  INV_X1 U4379 ( .A(n3371), .ZN(n3373) );
  XNOR2_X2 U4380 ( .A(n3373), .B(n3372), .ZN(n4651) );
  NAND2_X1 U4381 ( .A1(n4651), .A2(n3584), .ZN(n3377) );
  AOI22_X1 U4382 ( .A1(n3481), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n4802), .ZN(n3375) );
  NAND2_X1 U4383 ( .A1(n3419), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3374) );
  AND2_X1 U4384 ( .A1(n3375), .A2(n3374), .ZN(n3376) );
  NAND2_X1 U4385 ( .A1(n3377), .A2(n3376), .ZN(n4572) );
  INV_X1 U4386 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4807) );
  AOI22_X1 U4387 ( .A1(n3394), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3280), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3384) );
  BUF_X1 U4388 ( .A(n3395), .Z(n3378) );
  AOI22_X1 U4389 ( .A1(n3378), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3884), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3383) );
  AOI22_X1 U4390 ( .A1(n3208), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3206), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3382) );
  AOI22_X1 U4391 ( .A1(n3779), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3381) );
  NAND4_X1 U4392 ( .A1(n3384), .A2(n3383), .A3(n3382), .A4(n3381), .ZN(n3393)
         );
  AOI22_X1 U4393 ( .A1(n3207), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3391) );
  BUF_X1 U4394 ( .A(n3385), .Z(n3397) );
  AOI22_X1 U4395 ( .A1(n3397), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3787), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3390) );
  AOI22_X1 U4396 ( .A1(n3441), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3386), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3389) );
  AOI22_X1 U4397 ( .A1(n3387), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3217), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3388) );
  NAND4_X1 U4398 ( .A1(n3391), .A2(n3390), .A3(n3389), .A4(n3388), .ZN(n3392)
         );
  AOI21_X1 U4399 ( .B1(n4669), .B2(n4130), .A(n6530), .ZN(n3408) );
  AOI22_X1 U4400 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n3394), .B1(n3207), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3401) );
  AOI22_X1 U4401 ( .A1(n3378), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3208), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3400) );
  AOI22_X1 U4402 ( .A1(INSTQUEUE_REG_10__7__SCAN_IN), .A2(n3387), .B1(n3441), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3399) );
  AOI22_X1 U4403 ( .A1(n3397), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3386), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3398) );
  NAND4_X1 U4404 ( .A1(n3401), .A2(n3400), .A3(n3399), .A4(n3398), .ZN(n3407)
         );
  AOI22_X1 U4405 ( .A1(INSTQUEUE_REG_12__7__SCAN_IN), .A2(n3884), .B1(n3779), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3405) );
  AOI22_X1 U4406 ( .A1(n3860), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3280), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3404) );
  AOI22_X1 U4407 ( .A1(n3206), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3403) );
  AOI22_X1 U4408 ( .A1(n3380), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3217), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3402) );
  NAND4_X1 U4409 ( .A1(n3405), .A2(n3404), .A3(n3403), .A4(n3402), .ZN(n3406)
         );
  NAND2_X1 U4410 ( .A1(n4256), .A2(n4182), .ZN(n4179) );
  OAI211_X1 U4411 ( .C1(n3947), .C2(n4807), .A(n3408), .B(n4179), .ZN(n3414)
         );
  XNOR2_X1 U4412 ( .A(n4135), .B(n4182), .ZN(n3410) );
  NOR2_X1 U4413 ( .A1(n4674), .A2(n6530), .ZN(n3409) );
  NAND2_X1 U4414 ( .A1(n3410), .A2(n3409), .ZN(n3413) );
  AND2_X1 U4415 ( .A1(n3414), .A2(n3413), .ZN(n3411) );
  NAND2_X1 U4416 ( .A1(n3412), .A2(n3411), .ZN(n3416) );
  NAND2_X1 U4417 ( .A1(n3416), .A2(n3415), .ZN(n4658) );
  NAND2_X1 U4418 ( .A1(n6495), .A2(n3584), .ZN(n3423) );
  AOI22_X1 U4419 ( .A1(n3481), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n4802), .ZN(n3421) );
  NAND2_X1 U4420 ( .A1(n3419), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3420) );
  AND2_X1 U4421 ( .A1(n3421), .A2(n3420), .ZN(n3422) );
  NAND2_X1 U4422 ( .A1(n3423), .A2(n3422), .ZN(n4567) );
  NAND2_X1 U4423 ( .A1(n4568), .A2(n4567), .ZN(n4566) );
  OR2_X1 U4424 ( .A1(n4567), .A2(n3832), .ZN(n3424) );
  NAND2_X1 U4425 ( .A1(n4566), .A2(n3424), .ZN(n4571) );
  NAND2_X1 U4426 ( .A1(n4572), .A2(n4571), .ZN(n4573) );
  NAND2_X1 U4427 ( .A1(n3430), .A2(n4573), .ZN(n4580) );
  OAI21_X1 U4428 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A(n3426), .ZN(n5393) );
  AOI22_X1 U4429 ( .A1(n3903), .A2(n5393), .B1(n4201), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3428) );
  NAND2_X1 U4430 ( .A1(n3726), .A2(EAX_REG_2__SCAN_IN), .ZN(n3427) );
  OAI211_X1 U4431 ( .C1(n3429), .C2(n3425), .A(n3428), .B(n3427), .ZN(n4579)
         );
  NAND2_X1 U4432 ( .A1(n4580), .A2(n4579), .ZN(n3434) );
  INV_X1 U4433 ( .A(n4573), .ZN(n3432) );
  INV_X1 U4434 ( .A(n3430), .ZN(n3431) );
  NAND2_X1 U4435 ( .A1(n3432), .A2(n3431), .ZN(n3433) );
  NAND2_X1 U4436 ( .A1(n3434), .A2(n3433), .ZN(n4578) );
  NAND2_X1 U4437 ( .A1(n4586), .A2(n4578), .ZN(n4585) );
  INV_X1 U4438 ( .A(n4585), .ZN(n3435) );
  NAND2_X1 U4439 ( .A1(n3436), .A2(n3435), .ZN(n4740) );
  AOI22_X1 U4440 ( .A1(n3394), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3440) );
  AOI22_X1 U4441 ( .A1(n3879), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3838), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3439) );
  AOI22_X1 U4442 ( .A1(n3459), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3438) );
  AOI22_X1 U4443 ( .A1(n3378), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3437) );
  NAND4_X1 U4444 ( .A1(n3440), .A2(n3439), .A3(n3438), .A4(n3437), .ZN(n3447)
         );
  AOI22_X1 U4445 ( .A1(n3397), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3884), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3445) );
  INV_X1 U4446 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4359) );
  AOI22_X1 U4447 ( .A1(n3779), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3843), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3444) );
  AOI22_X1 U4448 ( .A1(n3387), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3443) );
  AOI22_X1 U4449 ( .A1(n3441), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3885), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3442) );
  NAND4_X1 U4450 ( .A1(n3445), .A2(n3444), .A3(n3443), .A4(n3442), .ZN(n3446)
         );
  NAND2_X1 U4451 ( .A1(n3955), .A2(n4157), .ZN(n3448) );
  XNOR2_X1 U4452 ( .A(n3457), .B(n3458), .ZN(n4153) );
  INV_X1 U4453 ( .A(EAX_REG_5__SCAN_IN), .ZN(n3454) );
  INV_X1 U4454 ( .A(n3451), .ZN(n3449) );
  AOI21_X1 U4455 ( .B1(n3449), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3452) );
  NAND2_X1 U4456 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3450) );
  OR2_X1 U4457 ( .A1(n3452), .A2(n3024), .ZN(n5925) );
  AOI22_X1 U4458 ( .A1(n5925), .A2(n3903), .B1(n4201), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3453) );
  OAI21_X1 U4459 ( .B1(n3455), .B2(n3454), .A(n3453), .ZN(n3456) );
  AOI21_X1 U4460 ( .B1(n4153), .B2(n3584), .A(n3456), .ZN(n4741) );
  NOR2_X2 U4461 ( .A1(n4740), .A2(n4741), .ZN(n4742) );
  NAND2_X1 U4462 ( .A1(n3930), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3471) );
  AOI22_X1 U4463 ( .A1(n3378), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3463) );
  AOI22_X1 U4464 ( .A1(n3394), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3462) );
  AOI22_X1 U4465 ( .A1(n3884), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3843), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3461) );
  AOI22_X1 U4466 ( .A1(n3441), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3885), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3460) );
  NAND4_X1 U4467 ( .A1(n3463), .A2(n3462), .A3(n3461), .A4(n3460), .ZN(n3469)
         );
  AOI22_X1 U4468 ( .A1(n3397), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3467) );
  AOI22_X1 U4469 ( .A1(n3860), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3466) );
  AOI22_X1 U4470 ( .A1(n3838), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3787), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3465) );
  AOI22_X1 U4471 ( .A1(n3387), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3464) );
  NAND4_X1 U4472 ( .A1(n3467), .A2(n3466), .A3(n3465), .A4(n3464), .ZN(n3468)
         );
  NAND2_X1 U4473 ( .A1(n3955), .A2(n4172), .ZN(n3470) );
  NAND2_X1 U4474 ( .A1(n3476), .A2(n3477), .ZN(n4165) );
  NAND2_X1 U4475 ( .A1(n4165), .A2(n3584), .ZN(n3475) );
  NOR2_X1 U4476 ( .A1(n3024), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3472)
         );
  OR2_X1 U4477 ( .A1(n3482), .A2(n3472), .ZN(n5914) );
  INV_X1 U4478 ( .A(n5914), .ZN(n6106) );
  AOI22_X1 U4479 ( .A1(n3726), .A2(EAX_REG_6__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n4802), .ZN(n3473) );
  MUX2_X1 U4480 ( .A(n6106), .B(n3473), .S(n3832), .Z(n3474) );
  NAND2_X1 U4481 ( .A1(n3475), .A2(n3474), .ZN(n4842) );
  NAND2_X1 U4482 ( .A1(n4742), .A2(n4842), .ZN(n4840) );
  INV_X1 U4483 ( .A(n3476), .ZN(n3479) );
  INV_X1 U4484 ( .A(n3477), .ZN(n3478) );
  NAND2_X1 U4485 ( .A1(n3479), .A2(n3478), .ZN(n4164) );
  AOI22_X1 U4486 ( .A1(INSTQUEUE_REG_0__7__SCAN_IN), .A2(n3930), .B1(n3955), 
        .B2(n4182), .ZN(n3480) );
  XNOR2_X1 U4487 ( .A(n4164), .B(n3480), .ZN(n4176) );
  INV_X1 U4488 ( .A(n4176), .ZN(n3487) );
  INV_X1 U4489 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3485) );
  NOR2_X1 U4490 ( .A1(n3482), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3483)
         );
  OR2_X1 U4491 ( .A1(n3514), .A2(n3483), .ZN(n5898) );
  AOI22_X1 U4492 ( .A1(n5898), .A2(n3903), .B1(n4201), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3484) );
  OAI21_X1 U4493 ( .B1(n3455), .B2(n3485), .A(n3484), .ZN(n3486) );
  AOI21_X1 U4494 ( .B1(n3487), .B2(n3584), .A(n3486), .ZN(n4919) );
  INV_X1 U4495 ( .A(n4919), .ZN(n3502) );
  AOI22_X1 U4496 ( .A1(n3395), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3491) );
  AOI22_X1 U4497 ( .A1(n3387), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3441), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3490) );
  AOI22_X1 U4498 ( .A1(n3860), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3489) );
  AOI22_X1 U4499 ( .A1(n3837), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3787), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3488) );
  NAND4_X1 U4500 ( .A1(n3491), .A2(n3490), .A3(n3489), .A4(n3488), .ZN(n3497)
         );
  AOI22_X1 U4501 ( .A1(n3394), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3495) );
  AOI22_X1 U4502 ( .A1(n3838), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3884), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3494) );
  AOI22_X1 U4503 ( .A1(n3397), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3843), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3493) );
  AOI22_X1 U4504 ( .A1(n3380), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3885), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3492) );
  NAND4_X1 U4505 ( .A1(n3495), .A2(n3494), .A3(n3493), .A4(n3492), .ZN(n3496)
         );
  OAI21_X1 U4506 ( .B1(n3497), .B2(n3496), .A(n3584), .ZN(n3500) );
  XOR2_X1 U4507 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3514), .Z(n5888) );
  INV_X1 U4508 ( .A(n5888), .ZN(n5054) );
  AOI22_X1 U4509 ( .A1(n4201), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n3903), 
        .B2(n5054), .ZN(n3499) );
  NAND2_X1 U4510 ( .A1(n3726), .A2(EAX_REG_8__SCAN_IN), .ZN(n3498) );
  INV_X1 U4511 ( .A(n5047), .ZN(n3501) );
  NAND2_X1 U4512 ( .A1(n3502), .A2(n3501), .ZN(n3503) );
  AOI22_X1 U4513 ( .A1(n3394), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3838), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3507) );
  AOI22_X1 U4514 ( .A1(n3378), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3884), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3506) );
  AOI22_X1 U4515 ( .A1(n3397), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3843), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3505) );
  AOI22_X1 U4516 ( .A1(n3779), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3504) );
  NAND4_X1 U4517 ( .A1(n3507), .A2(n3506), .A3(n3505), .A4(n3504), .ZN(n3513)
         );
  AOI22_X1 U4518 ( .A1(n3860), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3511) );
  AOI22_X1 U4519 ( .A1(n3879), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3510) );
  AOI22_X1 U4520 ( .A1(n3441), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3787), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3509) );
  AOI22_X1 U4521 ( .A1(n3387), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3885), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3508) );
  NAND4_X1 U4522 ( .A1(n3511), .A2(n3510), .A3(n3509), .A4(n3508), .ZN(n3512)
         );
  NOR2_X1 U4523 ( .A1(n3513), .A2(n3512), .ZN(n3518) );
  INV_X1 U4524 ( .A(n3520), .ZN(n3515) );
  XNOR2_X1 U4525 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3515), .ZN(n5385) );
  AOI22_X1 U4526 ( .A1(n3903), .A2(n5385), .B1(n4201), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3517) );
  NAND2_X1 U4527 ( .A1(n3726), .A2(EAX_REG_9__SCAN_IN), .ZN(n3516) );
  OAI211_X1 U4528 ( .C1(n3612), .C2(n3518), .A(n3517), .B(n3516), .ZN(n5008)
         );
  XOR2_X1 U4529 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3534), .Z(n5880) );
  AOI22_X1 U4530 ( .A1(n3394), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3524) );
  AOI22_X1 U4531 ( .A1(n3378), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3884), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3523) );
  AOI22_X1 U4532 ( .A1(n3397), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3843), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3522) );
  AOI22_X1 U4533 ( .A1(n3441), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3885), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3521) );
  NAND4_X1 U4534 ( .A1(n3524), .A2(n3523), .A3(n3522), .A4(n3521), .ZN(n3530)
         );
  AOI22_X1 U4535 ( .A1(n3860), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3528) );
  AOI22_X1 U4536 ( .A1(n3838), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3527) );
  AOI22_X1 U4537 ( .A1(n3779), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3787), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3526) );
  AOI22_X1 U4538 ( .A1(n3387), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3525) );
  NAND4_X1 U4539 ( .A1(n3528), .A2(n3527), .A3(n3526), .A4(n3525), .ZN(n3529)
         );
  OR2_X1 U4540 ( .A1(n3530), .A2(n3529), .ZN(n3531) );
  AOI22_X1 U4541 ( .A1(n3584), .A2(n3531), .B1(n4201), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3533) );
  NAND2_X1 U4542 ( .A1(n3726), .A2(EAX_REG_10__SCAN_IN), .ZN(n3532) );
  OAI211_X1 U4543 ( .C1(n5880), .C2(n3832), .A(n3533), .B(n3532), .ZN(n5018)
         );
  XNOR2_X1 U4544 ( .A(n3550), .B(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5593)
         );
  AOI22_X1 U4545 ( .A1(n3779), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3884), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3538) );
  AOI22_X1 U4546 ( .A1(n3860), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3537) );
  AOI22_X1 U4547 ( .A1(n3378), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3787), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3536) );
  AOI22_X1 U4548 ( .A1(n3387), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3535) );
  NAND4_X1 U4549 ( .A1(n3538), .A2(n3537), .A3(n3536), .A4(n3535), .ZN(n3544)
         );
  AOI22_X1 U4550 ( .A1(n3879), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3838), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3542) );
  AOI22_X1 U4551 ( .A1(n3394), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3541) );
  AOI22_X1 U4552 ( .A1(n3397), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3843), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3540) );
  AOI22_X1 U4553 ( .A1(n3441), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3885), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3539) );
  NAND4_X1 U4554 ( .A1(n3542), .A2(n3541), .A3(n3540), .A4(n3539), .ZN(n3543)
         );
  NOR2_X1 U4555 ( .A1(n3544), .A2(n3543), .ZN(n3547) );
  NAND2_X1 U4556 ( .A1(n3726), .A2(EAX_REG_11__SCAN_IN), .ZN(n3546) );
  NAND2_X1 U4557 ( .A1(n4201), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3545)
         );
  OAI211_X1 U4558 ( .C1(n3612), .C2(n3547), .A(n3546), .B(n3545), .ZN(n3548)
         );
  AOI21_X1 U4559 ( .B1(n5593), .B2(n3903), .A(n3548), .ZN(n5038) );
  INV_X1 U4560 ( .A(n5039), .ZN(n3569) );
  AOI21_X1 U4561 ( .B1(n4333), .B2(n3551), .A(n3023), .ZN(n6096) );
  OR2_X1 U4562 ( .A1(n6096), .A2(n3832), .ZN(n3567) );
  AOI22_X1 U4563 ( .A1(n3395), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3555) );
  AOI22_X1 U4564 ( .A1(n3387), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3554) );
  AOI22_X1 U4565 ( .A1(n3394), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3553) );
  AOI22_X1 U4566 ( .A1(n3884), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3843), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3552) );
  NAND4_X1 U4567 ( .A1(n3555), .A2(n3554), .A3(n3553), .A4(n3552), .ZN(n3561)
         );
  AOI22_X1 U4568 ( .A1(n3397), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3441), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3559) );
  AOI22_X1 U4569 ( .A1(n3860), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3558) );
  AOI22_X1 U4570 ( .A1(n3838), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3787), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3557) );
  AOI22_X1 U4571 ( .A1(n3380), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3885), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3556) );
  NAND4_X1 U4572 ( .A1(n3559), .A2(n3558), .A3(n3557), .A4(n3556), .ZN(n3560)
         );
  NOR2_X1 U4573 ( .A1(n3561), .A2(n3560), .ZN(n3564) );
  NAND2_X1 U4574 ( .A1(n3726), .A2(EAX_REG_12__SCAN_IN), .ZN(n3563) );
  NAND2_X1 U4575 ( .A1(n4201), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3562)
         );
  OAI211_X1 U4576 ( .C1(n3612), .C2(n3564), .A(n3563), .B(n3562), .ZN(n3565)
         );
  INV_X1 U4577 ( .A(n3565), .ZN(n3566) );
  XNOR2_X1 U4578 ( .A(n3023), .B(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5579)
         );
  NAND2_X1 U4579 ( .A1(n5579), .A2(n3903), .ZN(n3572) );
  INV_X1 U4580 ( .A(n4201), .ZN(n3819) );
  NOR2_X1 U4581 ( .A1(n3819), .A2(n3037), .ZN(n3570) );
  AOI21_X1 U4582 ( .B1(n3726), .B2(EAX_REG_13__SCAN_IN), .A(n3570), .ZN(n3571)
         );
  NAND2_X1 U4583 ( .A1(n3572), .A2(n3571), .ZN(n5339) );
  AOI22_X1 U4584 ( .A1(n3441), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3576) );
  AOI22_X1 U4585 ( .A1(n3394), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3838), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3575) );
  AOI22_X1 U4586 ( .A1(n3378), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3574) );
  AOI22_X1 U4587 ( .A1(n3397), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3573) );
  NAND4_X1 U4588 ( .A1(n3576), .A2(n3575), .A3(n3574), .A4(n3573), .ZN(n3582)
         );
  AOI22_X1 U4589 ( .A1(n3879), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3884), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3580) );
  AOI22_X1 U4590 ( .A1(n3387), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3579) );
  AOI22_X1 U4591 ( .A1(n3459), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3885), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3578) );
  AOI22_X1 U4592 ( .A1(n3787), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3843), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3577) );
  NAND4_X1 U4593 ( .A1(n3580), .A2(n3579), .A3(n3578), .A4(n3577), .ZN(n3581)
         );
  OR2_X1 U4594 ( .A1(n3582), .A2(n3581), .ZN(n3583) );
  AND2_X1 U4595 ( .A1(n3584), .A2(n3583), .ZN(n5338) );
  NAND2_X1 U4596 ( .A1(n5339), .A2(n5338), .ZN(n3614) );
  AOI22_X1 U4597 ( .A1(n3860), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3588) );
  AOI22_X1 U4598 ( .A1(INSTQUEUE_REG_4__7__SCAN_IN), .A2(n3441), .B1(n3884), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3587) );
  AOI22_X1 U4599 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n3208), .B1(n3837), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3586) );
  AOI22_X1 U4600 ( .A1(n3387), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3885), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3585) );
  NAND4_X1 U4601 ( .A1(n3588), .A2(n3587), .A3(n3586), .A4(n3585), .ZN(n3594)
         );
  AOI22_X1 U4602 ( .A1(n3394), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3592) );
  AOI22_X1 U4603 ( .A1(INSTQUEUE_REG_12__7__SCAN_IN), .A2(n3395), .B1(n3787), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3591) );
  AOI22_X1 U4604 ( .A1(n3385), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3843), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3590) );
  AOI22_X1 U4605 ( .A1(INSTQUEUE_REG_0__7__SCAN_IN), .A2(n3779), .B1(n3380), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3589) );
  NAND4_X1 U4606 ( .A1(n3592), .A2(n3591), .A3(n3590), .A4(n3589), .ZN(n3593)
         );
  NOR2_X1 U4607 ( .A1(n3594), .A2(n3593), .ZN(n3598) );
  XOR2_X1 U4608 ( .A(n3040), .B(n3626), .Z(n5866) );
  INV_X1 U4609 ( .A(n5866), .ZN(n3595) );
  AOI22_X1 U4610 ( .A1(n4201), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n3903), 
        .B2(n3595), .ZN(n3597) );
  NAND2_X1 U4611 ( .A1(n3726), .A2(EAX_REG_15__SCAN_IN), .ZN(n3596) );
  OAI211_X1 U4612 ( .C1(n3612), .C2(n3598), .A(n3597), .B(n3596), .ZN(n5426)
         );
  AOI22_X1 U4613 ( .A1(n3879), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3602) );
  AOI22_X1 U4614 ( .A1(n3838), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3884), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3601) );
  AOI22_X1 U4615 ( .A1(n3397), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3843), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3600) );
  AOI22_X1 U4616 ( .A1(n3387), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3885), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3599) );
  NAND4_X1 U4617 ( .A1(n3602), .A2(n3601), .A3(n3600), .A4(n3599), .ZN(n3608)
         );
  AOI22_X1 U4618 ( .A1(n3395), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3606) );
  AOI22_X1 U4619 ( .A1(n3394), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3605) );
  AOI22_X1 U4620 ( .A1(n3837), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3787), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3604) );
  AOI22_X1 U4621 ( .A1(n3441), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3603) );
  NAND4_X1 U4622 ( .A1(n3606), .A2(n3605), .A3(n3604), .A4(n3603), .ZN(n3607)
         );
  NOR2_X1 U4623 ( .A1(n3608), .A2(n3607), .ZN(n3611) );
  XNOR2_X1 U4624 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n2993), .ZN(n5573)
         );
  AOI22_X1 U4625 ( .A1(n3903), .A2(n5573), .B1(n4201), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3610) );
  NAND2_X1 U4626 ( .A1(n3726), .A2(EAX_REG_14__SCAN_IN), .ZN(n3609) );
  OAI211_X1 U4627 ( .C1(n3612), .C2(n3611), .A(n3610), .B(n3609), .ZN(n5341)
         );
  OAI211_X1 U4628 ( .C1(n5339), .C2(n5338), .A(n5426), .B(n5341), .ZN(n3613)
         );
  AOI22_X1 U4629 ( .A1(n3879), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3618) );
  AOI22_X1 U4630 ( .A1(n3779), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3884), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3617) );
  AOI22_X1 U4631 ( .A1(n3387), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3274), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3616) );
  AOI22_X1 U4632 ( .A1(n3838), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3787), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3615) );
  NAND4_X1 U4633 ( .A1(n3618), .A2(n3617), .A3(n3616), .A4(n3615), .ZN(n3624)
         );
  AOI22_X1 U4634 ( .A1(n3394), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3622) );
  AOI22_X1 U4635 ( .A1(n3378), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3621) );
  AOI22_X1 U4636 ( .A1(n3385), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3843), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3620) );
  AOI22_X1 U4637 ( .A1(n3380), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3885), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3619) );
  NAND4_X1 U4638 ( .A1(n3622), .A2(n3621), .A3(n3620), .A4(n3619), .ZN(n3623)
         );
  OR2_X1 U4639 ( .A1(n3624), .A2(n3623), .ZN(n3625) );
  NAND2_X1 U4640 ( .A1(n3900), .A2(n3625), .ZN(n3630) );
  XNOR2_X1 U4641 ( .A(n3645), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5565)
         );
  OAI22_X1 U4642 ( .A1(n5565), .A2(n3832), .B1(n3819), .B2(n3042), .ZN(n3628)
         );
  AOI21_X1 U4643 ( .B1(n3726), .B2(EAX_REG_16__SCAN_IN), .A(n3628), .ZN(n3629)
         );
  NAND2_X1 U4644 ( .A1(n3630), .A2(n3629), .ZN(n5322) );
  AOI22_X1 U4645 ( .A1(n3394), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3634) );
  AOI22_X1 U4646 ( .A1(n3879), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3633) );
  AOI22_X1 U4647 ( .A1(n3884), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3843), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3632) );
  AOI22_X1 U4648 ( .A1(n3779), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3631) );
  NAND4_X1 U4649 ( .A1(n3634), .A2(n3633), .A3(n3632), .A4(n3631), .ZN(n3640)
         );
  AOI22_X1 U4650 ( .A1(n3385), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3441), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3638) );
  AOI22_X1 U4651 ( .A1(n3208), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3637) );
  AOI22_X1 U4652 ( .A1(n3395), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3787), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3636) );
  AOI22_X1 U4653 ( .A1(n3387), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3885), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3635) );
  NAND4_X1 U4654 ( .A1(n3638), .A2(n3637), .A3(n3636), .A4(n3635), .ZN(n3639)
         );
  NOR2_X1 U4655 ( .A1(n3640), .A2(n3639), .ZN(n3644) );
  OAI21_X1 U4656 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6432), .A(n4802), 
        .ZN(n3641) );
  INV_X1 U4657 ( .A(n3641), .ZN(n3642) );
  AOI21_X1 U4658 ( .B1(n3726), .B2(EAX_REG_17__SCAN_IN), .A(n3642), .ZN(n3643)
         );
  OAI21_X1 U4659 ( .B1(n3872), .B2(n3644), .A(n3643), .ZN(n3648) );
  NAND2_X1 U4660 ( .A1(n3015), .A2(n3041), .ZN(n3646) );
  AND2_X1 U4661 ( .A1(n3664), .A2(n3646), .ZN(n5318) );
  NAND2_X1 U4662 ( .A1(n5318), .A2(n3903), .ZN(n3647) );
  NAND2_X1 U4663 ( .A1(n3648), .A2(n3647), .ZN(n5312) );
  XNOR2_X1 U4664 ( .A(n3664), .B(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5544)
         );
  AOI22_X1 U4665 ( .A1(n3394), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3838), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3653) );
  AOI22_X1 U4666 ( .A1(n3378), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3884), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3652) );
  AOI22_X1 U4667 ( .A1(n3385), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3651) );
  AOI22_X1 U4668 ( .A1(n3380), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3885), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3650) );
  NAND4_X1 U4669 ( .A1(n3653), .A2(n3652), .A3(n3651), .A4(n3650), .ZN(n3659)
         );
  AOI22_X1 U4670 ( .A1(n3860), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3280), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3657) );
  AOI22_X1 U4671 ( .A1(n3387), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3441), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3656) );
  AOI22_X1 U4672 ( .A1(n3879), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3655) );
  AOI22_X1 U4673 ( .A1(n3787), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3843), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3654) );
  NAND4_X1 U4674 ( .A1(n3657), .A2(n3656), .A3(n3655), .A4(n3654), .ZN(n3658)
         );
  OR2_X1 U4675 ( .A1(n3659), .A2(n3658), .ZN(n3662) );
  INV_X1 U4676 ( .A(EAX_REG_18__SCAN_IN), .ZN(n3660) );
  INV_X1 U4677 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5546) );
  OAI22_X1 U4678 ( .A1(n3455), .A2(n3660), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5546), .ZN(n3661) );
  AOI21_X1 U4679 ( .B1(n3900), .B2(n3662), .A(n3661), .ZN(n3663) );
  MUX2_X1 U4680 ( .A(n5544), .B(n3663), .S(n3832), .Z(n5300) );
  NAND2_X1 U4681 ( .A1(n3667), .A2(n3666), .ZN(n3668) );
  NAND2_X1 U4682 ( .A1(n3695), .A2(n3668), .ZN(n5537) );
  AOI22_X1 U4683 ( .A1(n3879), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3838), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3672) );
  AOI22_X1 U4684 ( .A1(n3378), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3884), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3671) );
  AOI22_X1 U4685 ( .A1(n3394), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3670) );
  AOI22_X1 U4686 ( .A1(n3779), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3885), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3669) );
  NAND4_X1 U4687 ( .A1(n3672), .A2(n3671), .A3(n3670), .A4(n3669), .ZN(n3678)
         );
  AOI22_X1 U4688 ( .A1(n3860), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3280), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3676) );
  AOI22_X1 U4689 ( .A1(n3397), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3787), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3675) );
  AOI22_X1 U4690 ( .A1(n3441), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3843), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3674) );
  AOI22_X1 U4691 ( .A1(n3387), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3673) );
  NAND4_X1 U4692 ( .A1(n3676), .A2(n3675), .A3(n3674), .A4(n3673), .ZN(n3677)
         );
  NOR2_X1 U4693 ( .A1(n3678), .A2(n3677), .ZN(n3680) );
  AOI22_X1 U4694 ( .A1(n3726), .A2(EAX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n4802), .ZN(n3679) );
  OAI21_X1 U4695 ( .B1(n3872), .B2(n3680), .A(n3679), .ZN(n3681) );
  MUX2_X1 U4696 ( .A(n5537), .B(n3681), .S(n3832), .Z(n5285) );
  XNOR2_X1 U4697 ( .A(n3695), .B(n3033), .ZN(n5274) );
  AOI22_X1 U4698 ( .A1(n3879), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3397), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3685) );
  AOI22_X1 U4699 ( .A1(n3274), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3684) );
  AOI22_X1 U4700 ( .A1(n3280), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3683) );
  AOI22_X1 U4701 ( .A1(n3380), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3885), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3682) );
  NAND4_X1 U4702 ( .A1(n3685), .A2(n3684), .A3(n3683), .A4(n3682), .ZN(n3691)
         );
  AOI22_X1 U4703 ( .A1(n3394), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3689) );
  AOI22_X1 U4704 ( .A1(n3395), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3884), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3688) );
  AOI22_X1 U4705 ( .A1(n3838), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3787), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3687) );
  AOI22_X1 U4706 ( .A1(n3387), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3843), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3686) );
  NAND4_X1 U4707 ( .A1(n3689), .A2(n3688), .A3(n3687), .A4(n3686), .ZN(n3690)
         );
  NOR2_X1 U4708 ( .A1(n3691), .A2(n3690), .ZN(n3693) );
  AOI22_X1 U4709 ( .A1(n3726), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n4802), .ZN(n3692) );
  OAI21_X1 U4710 ( .B1(n3872), .B2(n3693), .A(n3692), .ZN(n3694) );
  MUX2_X1 U4711 ( .A(n5274), .B(n3694), .S(n3832), .Z(n4455) );
  INV_X1 U4712 ( .A(n4453), .ZN(n3714) );
  NAND2_X1 U4713 ( .A1(n3697), .A2(n5529), .ZN(n3698) );
  AND2_X1 U4714 ( .A1(n3731), .A2(n3698), .ZN(n5533) );
  AOI22_X1 U4715 ( .A1(n3394), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3702) );
  AOI22_X1 U4716 ( .A1(n3208), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3701) );
  AOI22_X1 U4717 ( .A1(n3395), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3787), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3700) );
  AOI22_X1 U4718 ( .A1(n3274), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3699) );
  NAND4_X1 U4719 ( .A1(n3702), .A2(n3701), .A3(n3700), .A4(n3699), .ZN(n3708)
         );
  AOI22_X1 U4720 ( .A1(n3385), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3884), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3706) );
  AOI22_X1 U4721 ( .A1(n3879), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3705) );
  AOI22_X1 U4722 ( .A1(n3779), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3843), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3704) );
  AOI22_X1 U4723 ( .A1(n3387), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3885), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3703) );
  NAND4_X1 U4724 ( .A1(n3706), .A2(n3705), .A3(n3704), .A4(n3703), .ZN(n3707)
         );
  OR2_X1 U4725 ( .A1(n3708), .A2(n3707), .ZN(n3711) );
  INV_X1 U4726 ( .A(EAX_REG_21__SCAN_IN), .ZN(n3709) );
  OAI22_X1 U4727 ( .A1(n3455), .A2(n3709), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5529), .ZN(n3710) );
  AOI21_X1 U4728 ( .B1(n3900), .B2(n3711), .A(n3710), .ZN(n3712) );
  MUX2_X1 U4729 ( .A(n5533), .B(n3712), .S(n3832), .Z(n5257) );
  INV_X1 U4730 ( .A(n5257), .ZN(n3713) );
  NAND2_X2 U4731 ( .A1(n3714), .A2(n3713), .ZN(n5241) );
  AOI22_X1 U4732 ( .A1(n3394), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3718) );
  AOI22_X1 U4733 ( .A1(n3879), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3838), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3717) );
  AOI22_X1 U4734 ( .A1(n3459), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3716) );
  AOI22_X1 U4735 ( .A1(n3395), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3787), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3715) );
  NAND4_X1 U4736 ( .A1(n3718), .A2(n3717), .A3(n3716), .A4(n3715), .ZN(n3724)
         );
  AOI22_X1 U4737 ( .A1(n3385), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3722) );
  AOI22_X1 U4738 ( .A1(n3779), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3843), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3721) );
  AOI22_X1 U4739 ( .A1(n3387), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3720) );
  AOI22_X1 U4740 ( .A1(n3274), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3885), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3719) );
  NAND4_X1 U4741 ( .A1(n3722), .A2(n3721), .A3(n3720), .A4(n3719), .ZN(n3723)
         );
  NOR2_X1 U4742 ( .A1(n3724), .A2(n3723), .ZN(n3728) );
  AOI21_X1 U4743 ( .B1(n3034), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3725) );
  AOI21_X1 U4744 ( .B1(n3726), .B2(EAX_REG_22__SCAN_IN), .A(n3725), .ZN(n3727)
         );
  OAI21_X1 U4745 ( .B1(n3872), .B2(n3728), .A(n3727), .ZN(n3730) );
  XNOR2_X1 U4746 ( .A(n3731), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5522)
         );
  NAND2_X1 U4747 ( .A1(n5522), .A2(n3903), .ZN(n3729) );
  NAND2_X1 U4748 ( .A1(n3730), .A2(n3729), .ZN(n5242) );
  INV_X1 U4749 ( .A(n3733), .ZN(n3734) );
  INV_X1 U4750 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5492) );
  AOI21_X1 U4751 ( .B1(n3734), .B2(n5492), .A(n3874), .ZN(n5494) );
  AOI22_X1 U4752 ( .A1(n3394), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3738) );
  AOI22_X1 U4753 ( .A1(n3879), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3838), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3737) );
  AOI22_X1 U4754 ( .A1(n3459), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3736) );
  AOI22_X1 U4755 ( .A1(n3378), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3787), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3735) );
  NAND4_X1 U4756 ( .A1(n3738), .A2(n3737), .A3(n3736), .A4(n3735), .ZN(n3744)
         );
  AOI22_X1 U4757 ( .A1(n3397), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3884), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3742) );
  AOI22_X1 U4758 ( .A1(n3779), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3843), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3741) );
  AOI22_X1 U4759 ( .A1(n3387), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3740) );
  AOI22_X1 U4760 ( .A1(n3441), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3885), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3739) );
  NAND4_X1 U4761 ( .A1(n3742), .A2(n3741), .A3(n3740), .A4(n3739), .ZN(n3743)
         );
  OR2_X1 U4762 ( .A1(n3744), .A2(n3743), .ZN(n3835) );
  AOI22_X1 U4763 ( .A1(n3394), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3838), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3748) );
  AOI22_X1 U4764 ( .A1(n3397), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3747) );
  AOI22_X1 U4765 ( .A1(n3779), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3843), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3746) );
  AOI22_X1 U4766 ( .A1(n3380), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3885), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3745) );
  NAND4_X1 U4767 ( .A1(n3748), .A2(n3747), .A3(n3746), .A4(n3745), .ZN(n3754)
         );
  AOI22_X1 U4768 ( .A1(n3860), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3752) );
  AOI22_X1 U4769 ( .A1(n3378), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3884), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3751) );
  AOI22_X1 U4770 ( .A1(n3387), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3274), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3750) );
  AOI22_X1 U4771 ( .A1(n3879), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3749) );
  NAND4_X1 U4772 ( .A1(n3752), .A2(n3751), .A3(n3750), .A4(n3749), .ZN(n3753)
         );
  NOR2_X1 U4773 ( .A1(n3754), .A2(n3753), .ZN(n3802) );
  AOI22_X1 U4774 ( .A1(n3394), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3758) );
  AOI22_X1 U4775 ( .A1(n3879), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3838), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3757) );
  AOI22_X1 U4776 ( .A1(n3459), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3756) );
  AOI22_X1 U4777 ( .A1(n3378), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3787), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3755) );
  NAND4_X1 U4778 ( .A1(n3758), .A2(n3757), .A3(n3756), .A4(n3755), .ZN(n3764)
         );
  AOI22_X1 U4779 ( .A1(n3397), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3884), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3762) );
  AOI22_X1 U4780 ( .A1(n3779), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3843), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3761) );
  AOI22_X1 U4781 ( .A1(n3387), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3760) );
  AOI22_X1 U4782 ( .A1(n3441), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3885), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3759) );
  NAND4_X1 U4783 ( .A1(n3762), .A2(n3761), .A3(n3760), .A4(n3759), .ZN(n3763)
         );
  OR2_X1 U4784 ( .A1(n3764), .A2(n3763), .ZN(n3818) );
  INV_X1 U4785 ( .A(n3818), .ZN(n3786) );
  AOI22_X1 U4786 ( .A1(n3394), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3768) );
  AOI22_X1 U4787 ( .A1(n3879), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3838), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3767) );
  AOI22_X1 U4788 ( .A1(n3459), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3766) );
  INV_X1 U4789 ( .A(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4370) );
  AOI22_X1 U4790 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n3378), .B1(n3281), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3765) );
  NAND4_X1 U4791 ( .A1(n3768), .A2(n3767), .A3(n3766), .A4(n3765), .ZN(n3774)
         );
  AOI22_X1 U4792 ( .A1(INSTQUEUE_REG_8__7__SCAN_IN), .A2(n3397), .B1(n3884), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3772) );
  AOI22_X1 U4793 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n3779), .B1(n3843), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3771) );
  AOI22_X1 U4794 ( .A1(n3387), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3770) );
  AOI22_X1 U4795 ( .A1(n3441), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3885), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3769) );
  NAND4_X1 U4796 ( .A1(n3772), .A2(n3771), .A3(n3770), .A4(n3769), .ZN(n3773)
         );
  OR2_X1 U4797 ( .A1(n3774), .A2(n3773), .ZN(n3828) );
  AOI22_X1 U4798 ( .A1(n3394), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4799 ( .A1(n3879), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3838), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3777) );
  AOI22_X1 U4800 ( .A1(n3459), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3776) );
  AOI22_X1 U4801 ( .A1(n3378), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3787), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3775) );
  NAND4_X1 U4802 ( .A1(n3778), .A2(n3777), .A3(n3776), .A4(n3775), .ZN(n3785)
         );
  AOI22_X1 U4803 ( .A1(n3397), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3884), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3783) );
  AOI22_X1 U4804 ( .A1(n3779), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3843), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3782) );
  AOI22_X1 U4805 ( .A1(n3387), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3781) );
  AOI22_X1 U4806 ( .A1(n3441), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3885), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3780) );
  NAND4_X1 U4807 ( .A1(n3783), .A2(n3782), .A3(n3781), .A4(n3780), .ZN(n3784)
         );
  OR2_X1 U4808 ( .A1(n3785), .A2(n3784), .ZN(n3829) );
  NAND2_X1 U4809 ( .A1(n3828), .A2(n3829), .ZN(n3827) );
  NOR2_X1 U4810 ( .A1(n3786), .A2(n3827), .ZN(n3808) );
  AOI22_X1 U4811 ( .A1(n3394), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3791) );
  AOI22_X1 U4812 ( .A1(n3879), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3838), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3790) );
  AOI22_X1 U4813 ( .A1(n3459), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3789) );
  INV_X1 U4814 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4367) );
  AOI22_X1 U4815 ( .A1(n3378), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3787), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3788) );
  NAND4_X1 U4816 ( .A1(n3791), .A2(n3790), .A3(n3789), .A4(n3788), .ZN(n3797)
         );
  AOI22_X1 U4817 ( .A1(n3397), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3884), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3795) );
  AOI22_X1 U4818 ( .A1(n3779), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3843), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4819 ( .A1(n3387), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4820 ( .A1(n3441), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3885), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3792) );
  NAND4_X1 U4821 ( .A1(n3795), .A2(n3794), .A3(n3793), .A4(n3792), .ZN(n3796)
         );
  OR2_X1 U4822 ( .A1(n3797), .A2(n3796), .ZN(n3809) );
  NAND2_X1 U4823 ( .A1(n3808), .A2(n3809), .ZN(n3803) );
  NOR2_X1 U4824 ( .A1(n3802), .A2(n3803), .ZN(n3836) );
  XOR2_X1 U4825 ( .A(n3835), .B(n3836), .Z(n3800) );
  INV_X1 U4826 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4553) );
  NOR2_X1 U4827 ( .A1(n6432), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3798)
         );
  OAI22_X1 U4828 ( .A1(n3455), .A2(n4553), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3798), .ZN(n3799) );
  AOI21_X1 U4829 ( .B1(n3800), .B2(n3900), .A(n3799), .ZN(n3801) );
  AOI21_X1 U4830 ( .B1(n3903), .B2(n5494), .A(n3801), .ZN(n5208) );
  XOR2_X1 U4831 ( .A(n3803), .B(n3802), .Z(n3806) );
  INV_X1 U4832 ( .A(EAX_REG_26__SCAN_IN), .ZN(n3804) );
  INV_X1 U4833 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5505) );
  OAI22_X1 U4834 ( .A1(n3455), .A2(n3804), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5505), .ZN(n3805) );
  AOI21_X1 U4835 ( .B1(n3806), .B2(n3900), .A(n3805), .ZN(n3807) );
  XNOR2_X1 U4836 ( .A(n3815), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5503)
         );
  MUX2_X1 U4837 ( .A(n3807), .B(n5503), .S(n3903), .Z(n5150) );
  XNOR2_X1 U4838 ( .A(n3809), .B(n3808), .ZN(n3811) );
  AOI22_X1 U4839 ( .A1(n3726), .A2(EAX_REG_25__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n4802), .ZN(n3810) );
  OAI21_X1 U4840 ( .B1(n3872), .B2(n3811), .A(n3810), .ZN(n3816) );
  INV_X1 U4841 ( .A(n3812), .ZN(n3813) );
  INV_X1 U4842 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4476) );
  NAND2_X1 U4843 ( .A1(n3813), .A2(n4476), .ZN(n3814) );
  NAND2_X1 U4844 ( .A1(n3815), .A2(n3814), .ZN(n5141) );
  MUX2_X1 U4845 ( .A(n3816), .B(n5141), .S(n3903), .Z(n3817) );
  XNOR2_X1 U4846 ( .A(n3827), .B(n3818), .ZN(n3821) );
  INV_X1 U4847 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4515) );
  OAI22_X1 U4848 ( .A1(n3455), .A2(n4515), .B1(n3819), .B2(n4440), .ZN(n3820)
         );
  AOI21_X1 U4849 ( .B1(n3900), .B2(n3821), .A(n3820), .ZN(n3823) );
  XNOR2_X1 U4850 ( .A(n3826), .B(n4440), .ZN(n5124) );
  NAND2_X1 U4851 ( .A1(n5124), .A2(n3903), .ZN(n3822) );
  NOR2_X1 U4852 ( .A1(n3005), .A2(n4435), .ZN(n5147) );
  AND2_X1 U4853 ( .A1(n5208), .A2(n5147), .ZN(n3834) );
  NAND2_X1 U4854 ( .A1(n3824), .A2(n5514), .ZN(n3825) );
  NAND2_X1 U4855 ( .A1(n3826), .A2(n3825), .ZN(n5513) );
  OAI21_X1 U4856 ( .B1(n3829), .B2(n3828), .A(n3827), .ZN(n3831) );
  AOI22_X1 U4857 ( .A1(n3726), .A2(EAX_REG_23__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n4802), .ZN(n3830) );
  OAI21_X1 U4858 ( .B1(n3872), .B2(n3831), .A(n3830), .ZN(n3833) );
  MUX2_X1 U4859 ( .A(n5513), .B(n3833), .S(n3832), .Z(n5234) );
  AND2_X1 U4860 ( .A1(n3834), .A2(n5234), .ZN(n5168) );
  NAND2_X1 U4861 ( .A1(n3836), .A2(n3835), .ZN(n3858) );
  AOI22_X1 U4862 ( .A1(n3441), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3884), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3842) );
  AOI22_X1 U4863 ( .A1(n3860), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3841) );
  AOI22_X1 U4864 ( .A1(n3838), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3787), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4865 ( .A1(n3387), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3885), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3839) );
  NAND4_X1 U4866 ( .A1(n3842), .A2(n3841), .A3(n3840), .A4(n3839), .ZN(n3849)
         );
  AOI22_X1 U4867 ( .A1(n3378), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3847) );
  AOI22_X1 U4868 ( .A1(n3394), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3846) );
  AOI22_X1 U4869 ( .A1(n3397), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3843), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4870 ( .A1(n3779), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3844) );
  NAND4_X1 U4871 ( .A1(n3847), .A2(n3846), .A3(n3845), .A4(n3844), .ZN(n3848)
         );
  NOR2_X1 U4872 ( .A1(n3849), .A2(n3848), .ZN(n3859) );
  XOR2_X1 U4873 ( .A(n3858), .B(n3859), .Z(n3852) );
  INV_X1 U4874 ( .A(EAX_REG_28__SCAN_IN), .ZN(n3850) );
  INV_X1 U4875 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5172) );
  OAI22_X1 U4876 ( .A1(n3455), .A2(n3850), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5172), .ZN(n3851) );
  AOI21_X1 U4877 ( .B1(n3852), .B2(n3900), .A(n3851), .ZN(n3854) );
  INV_X1 U4878 ( .A(n3874), .ZN(n3853) );
  XNOR2_X1 U4879 ( .A(n3853), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5183)
         );
  MUX2_X1 U4880 ( .A(n3854), .B(n5183), .S(n3903), .Z(n5169) );
  INV_X1 U4881 ( .A(n5169), .ZN(n3855) );
  NAND2_X1 U4882 ( .A1(n5168), .A2(n3855), .ZN(n3856) );
  NOR2_X1 U4883 ( .A1(n3859), .A2(n3858), .ZN(n3894) );
  AOI22_X1 U4884 ( .A1(n3394), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3864) );
  AOI22_X1 U4885 ( .A1(n3879), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3208), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4886 ( .A1(n3459), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4887 ( .A1(n3378), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3787), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3861) );
  NAND4_X1 U4888 ( .A1(n3864), .A2(n3863), .A3(n3862), .A4(n3861), .ZN(n3870)
         );
  AOI22_X1 U4889 ( .A1(n3385), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3884), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3868) );
  AOI22_X1 U4890 ( .A1(n3779), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3843), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3867) );
  AOI22_X1 U4891 ( .A1(n3387), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3866) );
  AOI22_X1 U4892 ( .A1(n3274), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3885), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3865) );
  NAND4_X1 U4893 ( .A1(n3868), .A2(n3867), .A3(n3866), .A4(n3865), .ZN(n3869)
         );
  OR2_X1 U4894 ( .A1(n3870), .A2(n3869), .ZN(n3893) );
  XNOR2_X1 U4895 ( .A(n3894), .B(n3893), .ZN(n3873) );
  AOI22_X1 U4896 ( .A1(n3726), .A2(EAX_REG_29__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n4802), .ZN(n3871) );
  OAI21_X1 U4897 ( .B1(n3873), .B2(n3872), .A(n3871), .ZN(n3877) );
  INV_X1 U4898 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5484) );
  NAND2_X1 U4899 ( .A1(n3875), .A2(n5484), .ZN(n3876) );
  NAND2_X1 U4900 ( .A1(n3878), .A2(n3876), .ZN(n5483) );
  MUX2_X1 U4901 ( .A(n3877), .B(n5483), .S(n3903), .Z(n5200) );
  XOR2_X1 U4902 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .B(n3975), .Z(n4469) );
  AOI22_X1 U4903 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n3860), .B1(n3280), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3883) );
  AOI22_X1 U4904 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n3387), .B1(n3274), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3882) );
  AOI22_X1 U4905 ( .A1(n3879), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3837), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3881) );
  AOI22_X1 U4906 ( .A1(n3208), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3843), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3880) );
  NAND4_X1 U4907 ( .A1(n3883), .A2(n3882), .A3(n3881), .A4(n3880), .ZN(n3892)
         );
  AOI22_X1 U4908 ( .A1(n3378), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3884), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4909 ( .A1(n3385), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3889) );
  AOI22_X1 U4910 ( .A1(n3394), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3787), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3888) );
  AOI22_X1 U4911 ( .A1(n3380), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3885), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3887) );
  NAND4_X1 U4912 ( .A1(n3890), .A2(n3889), .A3(n3888), .A4(n3887), .ZN(n3891)
         );
  NOR2_X1 U4913 ( .A1(n3892), .A2(n3891), .ZN(n3896) );
  NAND2_X1 U4914 ( .A1(n3894), .A2(n3893), .ZN(n3895) );
  XOR2_X1 U4915 ( .A(n3896), .B(n3895), .Z(n3901) );
  INV_X1 U4916 ( .A(EAX_REG_30__SCAN_IN), .ZN(n3898) );
  OAI21_X1 U4917 ( .B1(n6432), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n4802), 
        .ZN(n3897) );
  OAI21_X1 U4918 ( .B1(n3455), .B2(n3898), .A(n3897), .ZN(n3899) );
  AOI21_X1 U4919 ( .B1(n3901), .B2(n3900), .A(n3899), .ZN(n3902) );
  AOI21_X1 U4920 ( .B1(n4469), .B2(n3903), .A(n3902), .ZN(n4199) );
  NAND2_X1 U4921 ( .A1(n6378), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3905) );
  XNOR2_X1 U4922 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3919) );
  XNOR2_X1 U4923 ( .A(n3920), .B(n3919), .ZN(n3967) );
  OAI21_X1 U4924 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6378), .A(n3905), 
        .ZN(n3910) );
  INV_X1 U4925 ( .A(n3910), .ZN(n3906) );
  NAND2_X1 U4926 ( .A1(n3904), .A2(n3906), .ZN(n3907) );
  NAND2_X1 U4927 ( .A1(n3907), .A2(n4248), .ZN(n3909) );
  NAND2_X1 U4928 ( .A1(n3242), .A2(n2985), .ZN(n3908) );
  NAND2_X1 U4929 ( .A1(n3909), .A2(n3935), .ZN(n3914) );
  OAI21_X1 U4930 ( .B1(n3923), .B2(n3242), .A(n2985), .ZN(n3916) );
  INV_X1 U4931 ( .A(n3967), .ZN(n3915) );
  NOR2_X1 U4932 ( .A1(n3923), .A2(n3910), .ZN(n3911) );
  OAI211_X1 U4933 ( .C1(n3916), .C2(n3915), .A(n3911), .B(n3914), .ZN(n3912)
         );
  NAND2_X1 U4934 ( .A1(n3912), .A2(n3938), .ZN(n3913) );
  OAI21_X1 U4935 ( .B1(n3967), .B2(n3914), .A(n3913), .ZN(n3918) );
  NAND3_X1 U4936 ( .A1(n3916), .A2(STATE2_REG_0__SCAN_IN), .A3(n3915), .ZN(
        n3917) );
  NAND2_X1 U4937 ( .A1(n3918), .A2(n3917), .ZN(n3933) );
  NAND2_X1 U4938 ( .A1(n3920), .A2(n3919), .ZN(n3922) );
  NAND2_X1 U4939 ( .A1(n6504), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3921) );
  NAND2_X1 U4940 ( .A1(n3922), .A2(n3921), .ZN(n3925) );
  XNOR2_X1 U4941 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3924) );
  XNOR2_X1 U4942 ( .A(n3925), .B(n3924), .ZN(n3968) );
  OAI21_X1 U4943 ( .B1(n3923), .B2(n3968), .A(n3935), .ZN(n3929) );
  NAND2_X1 U4944 ( .A1(n3925), .A2(n3924), .ZN(n3927) );
  NAND2_X1 U4945 ( .A1(n6306), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3926) );
  XNOR2_X1 U4946 ( .A(n3945), .B(n3944), .ZN(n3969) );
  INV_X1 U4947 ( .A(n3969), .ZN(n3928) );
  NAND2_X1 U4948 ( .A1(n3929), .A2(n3928), .ZN(n3934) );
  NAND2_X1 U4949 ( .A1(n3930), .A2(n3968), .ZN(n3931) );
  NAND2_X1 U4950 ( .A1(n3934), .A2(n3931), .ZN(n3932) );
  NAND2_X1 U4951 ( .A1(n3933), .A2(n3932), .ZN(n3942) );
  INV_X1 U4952 ( .A(n3934), .ZN(n3940) );
  INV_X1 U4953 ( .A(n3935), .ZN(n3937) );
  INV_X1 U4954 ( .A(n3968), .ZN(n3936) );
  AND3_X1 U4955 ( .A1(n3937), .A2(n3955), .A3(n3936), .ZN(n3939) );
  AOI22_X1 U4956 ( .A1(n3940), .A2(n3939), .B1(n3959), .B2(n3969), .ZN(n3941)
         );
  NAND2_X1 U4957 ( .A1(n3942), .A2(n3941), .ZN(n3949) );
  NOR2_X1 U4958 ( .A1(n6162), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3946)
         );
  NAND2_X1 U4959 ( .A1(n3947), .A2(n3966), .ZN(n3948) );
  NAND2_X1 U4960 ( .A1(n3949), .A2(n3948), .ZN(n3958) );
  AOI22_X1 U4961 ( .A1(n3959), .A2(n3966), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6530), .ZN(n3957) );
  INV_X1 U4962 ( .A(n3950), .ZN(n3952) );
  NAND2_X1 U4963 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n4723), .ZN(n3953) );
  NAND2_X1 U4964 ( .A1(n3955), .A2(n3965), .ZN(n3956) );
  INV_X1 U4965 ( .A(n3965), .ZN(n3971) );
  NAND2_X1 U4966 ( .A1(n3971), .A2(n3970), .ZN(n4509) );
  NOR2_X1 U4967 ( .A1(n4291), .A2(n4509), .ZN(n4500) );
  NAND2_X1 U4968 ( .A1(n4500), .A2(n4545), .ZN(n5802) );
  INV_X1 U4969 ( .A(n6663), .ZN(n6532) );
  NOR3_X1 U4970 ( .A1(n6530), .A2(n3238), .A3(n6532), .ZN(n6528) );
  NAND2_X1 U4971 ( .A1(n6530), .A2(n4802), .ZN(n6543) );
  NOR3_X1 U4972 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n6543), .A3(n4725), .ZN(
        n6539) );
  INV_X1 U4973 ( .A(n6539), .ZN(n3972) );
  NAND2_X1 U4974 ( .A1(n6122), .A2(n3972), .ZN(n3973) );
  INV_X1 U4975 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4225) );
  INV_X1 U4976 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6594) );
  NAND2_X1 U4977 ( .A1(n3268), .A2(n6660), .ZN(n4101) );
  NAND2_X1 U4978 ( .A1(n3978), .A2(n6559), .ZN(n6556) );
  OR2_X1 U4979 ( .A1(READY_N), .A2(n6556), .ZN(n4537) );
  NAND2_X1 U4980 ( .A1(n4101), .A2(n4537), .ZN(n4538) );
  AND3_X1 U4981 ( .A1(n4538), .A2(n6432), .A3(n4248), .ZN(n3979) );
  AND2_X2 U4982 ( .A1(n5392), .A2(n3979), .ZN(n5939) );
  INV_X1 U4983 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6592) );
  INV_X1 U4984 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6590) );
  INV_X1 U4985 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6587) );
  INV_X1 U4986 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6583) );
  INV_X1 U4987 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6572) );
  NAND3_X1 U4988 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n5937) );
  NOR2_X1 U4989 ( .A1(n6572), .A2(n5937), .ZN(n5915) );
  NAND2_X1 U4990 ( .A1(REIP_REG_5__SCAN_IN), .A2(n5915), .ZN(n5379) );
  NAND4_X1 U4991 ( .A1(REIP_REG_9__SCAN_IN), .A2(REIP_REG_8__SCAN_IN), .A3(
        REIP_REG_7__SCAN_IN), .A4(REIP_REG_6__SCAN_IN), .ZN(n5878) );
  NOR3_X1 U4992 ( .A1(n6583), .A2(n5379), .A3(n5878), .ZN(n5369) );
  NAND2_X1 U4993 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5369), .ZN(n5362) );
  NOR2_X1 U4994 ( .A1(n6587), .A2(n5362), .ZN(n5363) );
  NAND2_X1 U4995 ( .A1(REIP_REG_13__SCAN_IN), .A2(n5363), .ZN(n5350) );
  NOR2_X1 U4996 ( .A1(n6590), .A2(n5350), .ZN(n5329) );
  NAND2_X1 U4997 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5329), .ZN(n5325) );
  NOR2_X1 U4998 ( .A1(n6592), .A2(n5325), .ZN(n3983) );
  NAND2_X1 U4999 ( .A1(n5939), .A2(n3983), .ZN(n5317) );
  NOR2_X1 U5000 ( .A1(n6594), .A2(n5317), .ZN(n5305) );
  NAND2_X1 U5001 ( .A1(REIP_REG_20__SCAN_IN), .A2(n5273), .ZN(n5260) );
  INV_X1 U5002 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6605) );
  INV_X1 U5003 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6603) );
  NOR2_X1 U5004 ( .A1(n6605), .A2(n6603), .ZN(n5243) );
  NAND2_X1 U5005 ( .A1(REIP_REG_23__SCAN_IN), .A2(n5243), .ZN(n3988) );
  NOR2_X1 U5006 ( .A1(n5260), .A2(n3988), .ZN(n5122) );
  NAND2_X1 U5007 ( .A1(n5122), .A2(REIP_REG_24__SCAN_IN), .ZN(n5220) );
  AND2_X1 U5008 ( .A1(REIP_REG_26__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n3990) );
  INV_X1 U5009 ( .A(n3990), .ZN(n3980) );
  NAND2_X1 U5010 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n3993) );
  INV_X1 U5011 ( .A(n5202), .ZN(n3982) );
  INV_X1 U5012 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6621) );
  INV_X1 U5013 ( .A(REIP_REG_30__SCAN_IN), .ZN(n3981) );
  OAI21_X1 U5014 ( .B1(n3982), .B2(n6621), .A(n3981), .ZN(n4000) );
  NAND2_X1 U5015 ( .A1(n3983), .A2(REIP_REG_17__SCAN_IN), .ZN(n3984) );
  NAND2_X1 U5016 ( .A1(n5939), .A2(n3984), .ZN(n3985) );
  AND2_X1 U5017 ( .A1(n3985), .A2(n5975), .ZN(n5316) );
  INV_X1 U5018 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6596) );
  INV_X1 U5019 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6598) );
  NOR2_X1 U5020 ( .A1(n6596), .A2(n6598), .ZN(n5290) );
  NAND2_X1 U5021 ( .A1(n5290), .A2(REIP_REG_20__SCAN_IN), .ZN(n3986) );
  NAND2_X1 U5022 ( .A1(n5939), .A2(n3986), .ZN(n3987) );
  NAND2_X1 U5023 ( .A1(n5316), .A2(n3987), .ZN(n5272) );
  NAND2_X1 U5024 ( .A1(n5381), .A2(n5975), .ZN(n5928) );
  AND2_X1 U5025 ( .A1(n5928), .A2(n3988), .ZN(n3989) );
  NAND2_X1 U5026 ( .A1(n3990), .A2(REIP_REG_24__SCAN_IN), .ZN(n3991) );
  AND2_X1 U5027 ( .A1(n5928), .A2(n3991), .ZN(n3992) );
  NOR2_X1 U5028 ( .A1(n5121), .A2(n3992), .ZN(n5210) );
  NAND2_X1 U5029 ( .A1(n5939), .A2(n3993), .ZN(n3994) );
  AND2_X1 U5030 ( .A1(n5210), .A2(n3994), .ZN(n5181) );
  OAI211_X1 U5031 ( .C1(REIP_REG_29__SCAN_IN), .C2(n5381), .A(n5181), .B(
        REIP_REG_30__SCAN_IN), .ZN(n4221) );
  NAND2_X1 U5032 ( .A1(n6432), .A2(n6660), .ZN(n4093) );
  OR2_X1 U5033 ( .A1(n6556), .A2(n4093), .ZN(n6526) );
  AND2_X1 U5034 ( .A1(n2984), .A2(n6526), .ZN(n4222) );
  INV_X1 U5035 ( .A(n4222), .ZN(n3996) );
  INV_X1 U5036 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5410) );
  NAND3_X1 U5037 ( .A1(n4248), .A2(n4093), .A3(n5410), .ZN(n3995) );
  NAND2_X1 U5038 ( .A1(n3996), .A2(n3995), .ZN(n3997) );
  INV_X1 U5039 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5195) );
  AOI22_X1 U5040 ( .A1(n4469), .A2(n5948), .B1(n5960), .B2(
        PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n3998) );
  OAI21_X1 U5041 ( .B1(n5952), .B2(n5195), .A(n3998), .ZN(n3999) );
  NAND2_X1 U5042 ( .A1(n4248), .A2(n3268), .ZN(n4012) );
  INV_X1 U5043 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4577) );
  OR2_X1 U5045 ( .A1(n4016), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4004)
         );
  INV_X1 U5046 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4006) );
  OAI22_X1 U5047 ( .A1(n4087), .A2(n4006), .B1(n5269), .B2(EBX_REG_0__SCAN_IN), 
        .ZN(n4569) );
  XNOR2_X1 U5048 ( .A(n4007), .B(n4569), .ZN(n4575) );
  OR2_X1 U5049 ( .A1(n4008), .A2(EBX_REG_2__SCAN_IN), .ZN(n4011) );
  NAND2_X1 U5050 ( .A1(n5269), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4009)
         );
  OAI211_X1 U5051 ( .C1(n4576), .C2(EBX_REG_2__SCAN_IN), .A(n4087), .B(n4009), 
        .ZN(n4010) );
  AND2_X1 U5052 ( .A1(n4011), .A2(n4010), .ZN(n4603) );
  INV_X1 U5053 ( .A(EBX_REG_3__SCAN_IN), .ZN(n5953) );
  NAND2_X1 U5054 ( .A1(n4074), .A2(n5953), .ZN(n4015) );
  INV_X1 U5055 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4148) );
  NAND2_X1 U5056 ( .A1(n4087), .A2(n4148), .ZN(n4013) );
  INV_X4 U5057 ( .A(n3245), .ZN(n5269) );
  OAI211_X1 U5058 ( .C1(n4576), .C2(EBX_REG_3__SCAN_IN), .A(n4013), .B(n5269), 
        .ZN(n4014) );
  NAND2_X1 U5059 ( .A1(n4015), .A2(n4014), .ZN(n4589) );
  MUX2_X1 U5060 ( .A(n4008), .B(n5269), .S(EBX_REG_4__SCAN_IN), .Z(n4017) );
  OAI21_X1 U5061 ( .B1(n4016), .B2(INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4017), 
        .ZN(n4630) );
  NAND2_X1 U5062 ( .A1(n5269), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4019)
         );
  AND2_X1 U5063 ( .A1(n4087), .A2(n4019), .ZN(n4021) );
  NOR2_X1 U5064 ( .A1(n4576), .A2(EBX_REG_5__SCAN_IN), .ZN(n4020) );
  MUX2_X1 U5065 ( .A(n4021), .B(n5269), .S(n4020), .Z(n4745) );
  OR2_X1 U5066 ( .A1(n4016), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4024)
         );
  INV_X1 U5067 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4022) );
  MUX2_X1 U5068 ( .A(n5269), .B(n4008), .S(n4022), .Z(n4023) );
  AND2_X1 U5069 ( .A1(n4024), .A2(n4023), .ZN(n4889) );
  INV_X1 U5070 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4923) );
  NAND2_X1 U5071 ( .A1(n4074), .A2(n4923), .ZN(n4027) );
  INV_X1 U5072 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4178) );
  NAND2_X1 U5073 ( .A1(n4087), .A2(n4178), .ZN(n4025) );
  OAI211_X1 U5074 ( .C1(n4576), .C2(EBX_REG_7__SCAN_IN), .A(n4025), .B(n5269), 
        .ZN(n4026) );
  NAND2_X1 U5075 ( .A1(n4027), .A2(n4026), .ZN(n4921) );
  MUX2_X1 U5076 ( .A(n4008), .B(n5269), .S(EBX_REG_8__SCAN_IN), .Z(n4028) );
  OAI21_X1 U5077 ( .B1(n4016), .B2(INSTADDRPOINTER_REG_8__SCAN_IN), .A(n4028), 
        .ZN(n5058) );
  INV_X1 U5078 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5015) );
  NAND2_X1 U5079 ( .A1(n4074), .A2(n5015), .ZN(n4032) );
  INV_X1 U5080 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5773) );
  NAND2_X1 U5081 ( .A1(n4087), .A2(n5773), .ZN(n4030) );
  OAI211_X1 U5082 ( .C1(n4576), .C2(EBX_REG_9__SCAN_IN), .A(n4030), .B(n5269), 
        .ZN(n4031) );
  AND2_X1 U5083 ( .A1(n4032), .A2(n4031), .ZN(n5013) );
  INV_X1 U5084 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5030) );
  MUX2_X1 U5085 ( .A(n5269), .B(n4008), .S(n5030), .Z(n4034) );
  OAI21_X1 U5086 ( .B1(n4016), .B2(INSTADDRPOINTER_REG_10__SCAN_IN), .A(n4034), 
        .ZN(n5028) );
  INV_X1 U5087 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5373) );
  NAND2_X1 U5088 ( .A1(n4074), .A2(n5373), .ZN(n4037) );
  INV_X1 U5089 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U5090 ( .A1(n4087), .A2(n5588), .ZN(n4035) );
  OAI211_X1 U5091 ( .C1(n4576), .C2(EBX_REG_11__SCAN_IN), .A(n4035), .B(n5269), 
        .ZN(n4036) );
  NAND2_X1 U5092 ( .A1(n4037), .A2(n4036), .ZN(n5042) );
  MUX2_X1 U5093 ( .A(n4008), .B(n5269), .S(EBX_REG_12__SCAN_IN), .Z(n4038) );
  OAI21_X1 U5094 ( .B1(n4016), .B2(INSTADDRPOINTER_REG_12__SCAN_IN), .A(n4038), 
        .ZN(n5765) );
  NAND2_X1 U5095 ( .A1(n5269), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4040) );
  NAND2_X1 U5096 ( .A1(n4087), .A2(n4040), .ZN(n4042) );
  NOR2_X1 U5097 ( .A1(n4576), .A2(EBX_REG_13__SCAN_IN), .ZN(n4041) );
  MUX2_X1 U5098 ( .A(n4042), .B(n3245), .S(n4041), .Z(n5359) );
  OR2_X1 U5099 ( .A1(n4008), .A2(EBX_REG_14__SCAN_IN), .ZN(n4045) );
  NAND2_X1 U5100 ( .A1(n5269), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4043) );
  OAI211_X1 U5101 ( .C1(n4576), .C2(EBX_REG_14__SCAN_IN), .A(n4087), .B(n4043), 
        .ZN(n4044) );
  NAND2_X1 U5102 ( .A1(n4016), .A2(EBX_REG_15__SCAN_IN), .ZN(n4047) );
  NAND2_X1 U5103 ( .A1(n4576), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4046) );
  NAND2_X1 U5104 ( .A1(n4047), .A2(n4046), .ZN(n4048) );
  XNOR2_X1 U5105 ( .A(n4048), .B(n5269), .ZN(n5429) );
  OR2_X1 U5106 ( .A1(n4008), .A2(EBX_REG_16__SCAN_IN), .ZN(n4051) );
  NAND2_X1 U5107 ( .A1(n5269), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4049) );
  OAI211_X1 U5108 ( .C1(n4576), .C2(EBX_REG_16__SCAN_IN), .A(n4087), .B(n4049), 
        .ZN(n4050) );
  NAND2_X1 U5109 ( .A1(n5269), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4053) );
  NAND2_X1 U5110 ( .A1(n4087), .A2(n4053), .ZN(n4055) );
  NOR2_X1 U5111 ( .A1(n4576), .A2(EBX_REG_17__SCAN_IN), .ZN(n4054) );
  MUX2_X1 U5112 ( .A(n4055), .B(n3245), .S(n4054), .Z(n5315) );
  NAND2_X1 U5113 ( .A1(n5313), .A2(n5315), .ZN(n5281) );
  INV_X2 U5114 ( .A(n5281), .ZN(n4059) );
  MUX2_X1 U5115 ( .A(n4008), .B(n5269), .S(EBX_REG_19__SCAN_IN), .Z(n4057) );
  OR2_X1 U5116 ( .A1(n4016), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4056)
         );
  NAND2_X1 U5117 ( .A1(n4057), .A2(n4056), .ZN(n5283) );
  NAND2_X1 U5118 ( .A1(n4016), .A2(EBX_REG_18__SCAN_IN), .ZN(n4061) );
  NAND2_X1 U5119 ( .A1(n4576), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4060) );
  INV_X1 U5120 ( .A(n5282), .ZN(n4063) );
  OAI22_X1 U5121 ( .A1(n4016), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        EBX_REG_20__SCAN_IN), .B2(n4576), .ZN(n5270) );
  MUX2_X1 U5122 ( .A(n5269), .B(n5282), .S(n5270), .Z(n4062) );
  OAI21_X1 U5123 ( .B1(n3245), .B2(n4063), .A(n4062), .ZN(n4064) );
  MUX2_X1 U5124 ( .A(n4008), .B(n5269), .S(EBX_REG_21__SCAN_IN), .Z(n4066) );
  OR2_X1 U5125 ( .A1(n4016), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4065)
         );
  NAND2_X1 U5126 ( .A1(n5269), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4067) );
  AND2_X1 U5127 ( .A1(n4087), .A2(n4067), .ZN(n4069) );
  NOR2_X1 U5128 ( .A1(n4576), .A2(EBX_REG_22__SCAN_IN), .ZN(n4068) );
  MUX2_X1 U5129 ( .A(n4069), .B(n5269), .S(n4068), .Z(n5229) );
  OR2_X1 U5130 ( .A1(n4008), .A2(EBX_REG_23__SCAN_IN), .ZN(n4072) );
  NAND2_X1 U5131 ( .A1(n5269), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4070) );
  OAI211_X1 U5132 ( .C1(n4576), .C2(EBX_REG_23__SCAN_IN), .A(n4087), .B(n4070), 
        .ZN(n4071) );
  NAND2_X1 U5133 ( .A1(n4072), .A2(n4071), .ZN(n5228) );
  INV_X1 U5134 ( .A(EBX_REG_24__SCAN_IN), .ZN(n4073) );
  NAND2_X1 U5135 ( .A1(n4074), .A2(n4073), .ZN(n4077) );
  INV_X1 U5136 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5663) );
  NAND2_X1 U5137 ( .A1(n4087), .A2(n5663), .ZN(n4075) );
  OAI211_X1 U5138 ( .C1(EBX_REG_24__SCAN_IN), .C2(n4576), .A(n4075), .B(n5269), 
        .ZN(n4076) );
  INV_X1 U5139 ( .A(n5119), .ZN(n4078) );
  MUX2_X1 U5140 ( .A(n4008), .B(n5269), .S(EBX_REG_25__SCAN_IN), .Z(n4080) );
  OR2_X1 U5141 ( .A1(n4016), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4079)
         );
  INV_X1 U5142 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5647) );
  NAND2_X1 U5143 ( .A1(n4087), .A2(n5647), .ZN(n4081) );
  OAI211_X1 U5144 ( .C1(EBX_REG_26__SCAN_IN), .C2(n4576), .A(n4081), .B(n5269), 
        .ZN(n4082) );
  OAI21_X1 U5145 ( .B1(EBX_REG_26__SCAN_IN), .B2(n4083), .A(n4082), .ZN(n5152)
         );
  MUX2_X1 U5146 ( .A(n4008), .B(n5269), .S(EBX_REG_27__SCAN_IN), .Z(n4085) );
  OR2_X1 U5147 ( .A1(n4016), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4084)
         );
  NAND2_X1 U5148 ( .A1(n4085), .A2(n4084), .ZN(n5214) );
  NAND2_X1 U5149 ( .A1(n5269), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4086) );
  AND2_X1 U5150 ( .A1(n4087), .A2(n4086), .ZN(n4089) );
  NOR2_X1 U5151 ( .A1(n4576), .A2(EBX_REG_28__SCAN_IN), .ZN(n4088) );
  MUX2_X1 U5152 ( .A(n4089), .B(n5269), .S(n4088), .Z(n5179) );
  OAI22_X1 U5153 ( .A1(n4016), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        EBX_REG_29__SCAN_IN), .B2(n4576), .ZN(n4213) );
  AOI22_X1 U5154 ( .A1(n4016), .A2(EBX_REG_30__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n4576), .ZN(n4218) );
  NAND2_X1 U5155 ( .A1(n4093), .A2(EBX_REG_31__SCAN_IN), .ZN(n4094) );
  NOR2_X1 U5156 ( .A1(n4576), .A2(n4094), .ZN(n4095) );
  NAND2_X1 U5157 ( .A1(n4096), .A2(n3007), .ZN(U2797) );
  NOR2_X4 U5158 ( .A1(n5241), .A2(n5242), .ZN(n5232) );
  INV_X1 U5159 ( .A(n4435), .ZN(n4097) );
  NAND2_X1 U5160 ( .A1(n5148), .A2(n4097), .ZN(n4436) );
  INV_X1 U5161 ( .A(n5233), .ZN(n4099) );
  OAI21_X1 U5162 ( .B1(n4527), .B2(n2959), .A(n4669), .ZN(n4103) );
  NAND2_X1 U5163 ( .A1(n4102), .A2(n4103), .ZN(n4239) );
  NOR2_X1 U5164 ( .A1(n4239), .A2(n4104), .ZN(n4696) );
  NAND2_X1 U5165 ( .A1(n4540), .A2(n4696), .ZN(n4107) );
  INV_X1 U5166 ( .A(n4105), .ZN(n4726) );
  NOR2_X1 U5167 ( .A1(READY_N), .A2(n4509), .ZN(n4241) );
  NAND2_X1 U5168 ( .A1(n4726), .A2(n4241), .ZN(n4106) );
  NAND2_X1 U5169 ( .A1(n4107), .A2(n4106), .ZN(n4536) );
  AND3_X1 U5170 ( .A1(n4256), .A2(n3231), .A3(n4685), .ZN(n4485) );
  AND2_X1 U5171 ( .A1(n2959), .A2(n4661), .ZN(n4111) );
  NOR2_X1 U5172 ( .A1(n4111), .A2(n4265), .ZN(n4110) );
  NAND2_X1 U5173 ( .A1(n5138), .A2(n5989), .ZN(n4114) );
  AND2_X1 U5174 ( .A1(n5991), .A2(n4265), .ZN(n5467) );
  AOI22_X1 U5175 ( .A1(n5467), .A2(DATAI_25_), .B1(n5473), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n4113) );
  NAND2_X1 U5176 ( .A1(n5468), .A2(DATAI_9_), .ZN(n4112) );
  NAND2_X1 U5177 ( .A1(n4115), .A2(n4163), .ZN(n4119) );
  NAND2_X1 U5178 ( .A1(n4134), .A2(n4130), .ZN(n4122) );
  NAND2_X1 U5179 ( .A1(n4122), .A2(n4116), .ZN(n4145) );
  NAND2_X1 U5180 ( .A1(n4145), .A2(n4146), .ZN(n4156) );
  XNOR2_X1 U5181 ( .A(n4156), .B(n4154), .ZN(n4117) );
  NAND2_X1 U5182 ( .A1(n4117), .A2(n2984), .ZN(n4118) );
  NAND2_X1 U5183 ( .A1(n4119), .A2(n4118), .ZN(n4152) );
  INV_X1 U5184 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4120) );
  XNOR2_X1 U5185 ( .A(n4152), .B(n4120), .ZN(n4624) );
  NAND2_X1 U5186 ( .A1(n4653), .A2(n4163), .ZN(n4128) );
  INV_X1 U5187 ( .A(n4122), .ZN(n4121) );
  NOR2_X1 U5188 ( .A1(n6662), .A2(n4121), .ZN(n4138) );
  NOR2_X1 U5189 ( .A1(n6662), .A2(n4122), .ZN(n4124) );
  MUX2_X1 U5190 ( .A(n4138), .B(n4124), .S(n4123), .Z(n4126) );
  NAND2_X1 U5191 ( .A1(n4669), .A2(n3243), .ZN(n4129) );
  INV_X1 U5192 ( .A(n4129), .ZN(n4125) );
  NOR2_X1 U5193 ( .A1(n4126), .A2(n4125), .ZN(n4127) );
  NAND2_X1 U5194 ( .A1(n4128), .A2(n4127), .ZN(n4592) );
  NAND2_X1 U5195 ( .A1(n4658), .A2(n4163), .ZN(n4133) );
  OAI21_X1 U5196 ( .B1(n6662), .B2(n4130), .A(n4129), .ZN(n4131) );
  INV_X1 U5197 ( .A(n4131), .ZN(n4132) );
  NAND2_X1 U5198 ( .A1(n4133), .A2(n4132), .ZN(n5610) );
  NAND2_X1 U5199 ( .A1(n4651), .A2(n4163), .ZN(n4140) );
  INV_X1 U5200 ( .A(n4134), .ZN(n4136) );
  NAND2_X1 U5201 ( .A1(n4136), .A2(n4135), .ZN(n4137) );
  NAND2_X1 U5202 ( .A1(n4140), .A2(n4139), .ZN(n4617) );
  NAND2_X1 U5203 ( .A1(n4616), .A2(n4617), .ZN(n4615) );
  INV_X1 U5204 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6159) );
  OR2_X1 U5205 ( .A1(n4141), .A2(n6159), .ZN(n4142) );
  OAI21_X1 U5206 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n4592), .A(n4593), 
        .ZN(n4144) );
  NAND2_X1 U5207 ( .A1(n4592), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4143)
         );
  NAND2_X1 U5208 ( .A1(n4144), .A2(n4143), .ZN(n4634) );
  INV_X1 U5209 ( .A(n4163), .ZN(n4175) );
  OAI211_X1 U5210 ( .C1(n4146), .C2(n4145), .A(n4156), .B(n2984), .ZN(n4147)
         );
  NAND2_X1 U5211 ( .A1(n4149), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4150)
         );
  NAND2_X1 U5212 ( .A1(n4153), .A2(n4163), .ZN(n4160) );
  INV_X1 U5213 ( .A(n4154), .ZN(n4155) );
  NOR2_X1 U5214 ( .A1(n4156), .A2(n4155), .ZN(n4158) );
  NAND2_X1 U5215 ( .A1(n4158), .A2(n4157), .ZN(n4171) );
  OAI211_X1 U5216 ( .C1(n4158), .C2(n4157), .A(n4171), .B(n2984), .ZN(n4159)
         );
  NAND2_X1 U5217 ( .A1(n4160), .A2(n4159), .ZN(n4161) );
  NAND2_X1 U5218 ( .A1(n4181), .A2(n4165), .ZN(n4168) );
  XNOR2_X1 U5219 ( .A(n4171), .B(n4172), .ZN(n4166) );
  NAND2_X1 U5220 ( .A1(n4166), .A2(n2984), .ZN(n4167) );
  NAND2_X1 U5221 ( .A1(n4168), .A2(n4167), .ZN(n4170) );
  INV_X1 U5222 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4169) );
  XNOR2_X1 U5223 ( .A(n4170), .B(n4169), .ZN(n4887) );
  INV_X1 U5224 ( .A(n4171), .ZN(n4173) );
  NAND2_X1 U5225 ( .A1(n4173), .A2(n4172), .ZN(n4184) );
  XOR2_X1 U5226 ( .A(n4182), .B(n4184), .Z(n4174) );
  OAI22_X1 U5227 ( .A1(n4176), .A2(n4175), .B1(n4174), .B2(n6662), .ZN(n4177)
         );
  XNOR2_X1 U5228 ( .A(n4177), .B(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4927)
         );
  NAND2_X1 U5229 ( .A1(n2984), .A2(n4182), .ZN(n4183) );
  INV_X1 U5230 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4185) );
  NOR4_X1 U5231 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(INSTADDRPOINTER_REG_11__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4187) );
  NOR2_X1 U5232 ( .A1(n2992), .A2(n4187), .ZN(n4189) );
  AND2_X1 U5233 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4188) );
  AOI21_X1 U5234 ( .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A(n5587), .ZN(n4191) );
  NOR2_X1 U5235 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4190) );
  INV_X1 U5236 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5569) );
  NAND2_X1 U5237 ( .A1(n2992), .A2(n5569), .ZN(n5568) );
  NAND2_X1 U5238 ( .A1(n5587), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5751) );
  NOR2_X1 U5239 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5700) );
  INV_X1 U5240 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5718) );
  INV_X1 U5241 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5727) );
  INV_X1 U5242 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5729) );
  AND3_X1 U5243 ( .A1(n5718), .A2(n5727), .A3(n5729), .ZN(n4448) );
  AOI21_X1 U5244 ( .B1(n5700), .B2(n4448), .A(n2992), .ZN(n4193) );
  NAND2_X1 U5245 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4284) );
  OAI21_X1 U5246 ( .B1(n5718), .B2(n4284), .A(n2992), .ZN(n4192) );
  NOR2_X1 U5247 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4299) );
  INV_X1 U5248 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5675) );
  NAND3_X1 U5249 ( .A1(n4299), .A2(n5663), .A3(n5675), .ZN(n4194) );
  NAND2_X1 U5250 ( .A1(n5587), .A2(n4194), .ZN(n4196) );
  AND2_X1 U5251 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5699) );
  AND2_X1 U5252 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4422) );
  AND2_X1 U5253 ( .A1(n5699), .A2(n4422), .ZN(n5676) );
  AND2_X1 U5254 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4425) );
  NAND2_X1 U5255 ( .A1(n5676), .A2(n4425), .ZN(n4421) );
  INV_X1 U5256 ( .A(n4421), .ZN(n4195) );
  XOR2_X1 U5257 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .B(n2992), .Z(n4474) );
  INV_X1 U5258 ( .A(n4473), .ZN(n5490) );
  NOR2_X1 U5259 ( .A1(n5587), .A2(n5647), .ZN(n5500) );
  INV_X1 U5260 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5656) );
  AND2_X1 U5261 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5617) );
  NAND2_X1 U5262 ( .A1(n5617), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5129) );
  NOR4_X1 U5263 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .A3(INSTADDRPOINTER_REG_26__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4197) );
  XNOR2_X1 U5264 ( .A(n4198), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4434)
         );
  AOI22_X1 U5265 ( .A1(n3726), .A2(EAX_REG_31__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n4201), .ZN(n4202) );
  NAND3_X1 U5266 ( .A1(n6530), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6544) );
  NAND2_X1 U5267 ( .A1(n2957), .A2(n6104), .ZN(n4211) );
  NAND2_X1 U5268 ( .A1(n6435), .A2(n4204), .ZN(n6659) );
  NAND2_X1 U5269 ( .A1(n6659), .A2(n6530), .ZN(n4205) );
  INV_X1 U5270 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6625) );
  NOR2_X1 U5271 ( .A1(n6122), .A2(n6625), .ZN(n4431) );
  NAND2_X1 U5272 ( .A1(n6530), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4207) );
  NAND2_X1 U5273 ( .A1(n6432), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4206) );
  NAND2_X1 U5274 ( .A1(n4207), .A2(n4206), .ZN(n5611) );
  NOR2_X1 U5275 ( .A1(n5594), .A2(n4208), .ZN(n4209) );
  AOI211_X1 U5276 ( .C1(n6094), .C2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n4431), 
        .B(n4209), .ZN(n4210) );
  OAI21_X1 U5277 ( .B1(n4434), .B2(n6100), .A(n4212), .ZN(U2955) );
  INV_X1 U5278 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5412) );
  NOR2_X1 U5279 ( .A1(n5269), .A2(n5412), .ZN(n4215) );
  AOI21_X1 U5280 ( .B1(n4213), .B2(n5269), .A(n4215), .ZN(n5198) );
  INV_X1 U5281 ( .A(n4215), .ZN(n4216) );
  OAI211_X1 U5282 ( .C1(n5197), .C2(n4218), .A(n4217), .B(n4216), .ZN(n4220)
         );
  AOI22_X1 U5283 ( .A1(n4016), .A2(EBX_REG_31__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4576), .ZN(n4219) );
  XNOR2_X1 U5284 ( .A(n4220), .B(n4219), .ZN(n5409) );
  AND3_X1 U5285 ( .A1(n4221), .A2(REIP_REG_31__SCAN_IN), .A3(n5928), .ZN(n4227) );
  NAND4_X1 U5286 ( .A1(n5202), .A2(REIP_REG_30__SCAN_IN), .A3(
        REIP_REG_29__SCAN_IN), .A4(n6625), .ZN(n4224) );
  NAND3_X1 U5287 ( .A1(n5392), .A2(EBX_REG_31__SCAN_IN), .A3(n4222), .ZN(n4223) );
  OAI211_X1 U5288 ( .C1(n5908), .C2(n4225), .A(n4224), .B(n4223), .ZN(n4226)
         );
  AOI211_X1 U5289 ( .C1(n5409), .C2(n5927), .A(n4227), .B(n4226), .ZN(n4230)
         );
  NAND2_X1 U5290 ( .A1(n4230), .A2(n4229), .ZN(U2796) );
  INV_X1 U5291 ( .A(n5699), .ZN(n4231) );
  XNOR2_X1 U5292 ( .A(n5587), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5527)
         );
  INV_X1 U5293 ( .A(n5526), .ZN(n4234) );
  NOR2_X1 U5294 ( .A1(n2992), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4444)
         );
  AOI21_X1 U5295 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n2991), .A(n4444), 
        .ZN(n4235) );
  NOR2_X1 U5296 ( .A1(n4527), .A2(n3242), .ZN(n4280) );
  INV_X1 U5297 ( .A(n4280), .ZN(n4244) );
  NAND2_X1 U5298 ( .A1(n4237), .A2(n4248), .ZN(n4238) );
  MUX2_X1 U5299 ( .A(n6662), .B(n4238), .S(n3228), .Z(n4272) );
  INV_X1 U5300 ( .A(n4272), .ZN(n4240) );
  OAI21_X1 U5301 ( .B1(n4240), .B2(n4239), .A(n4291), .ZN(n4533) );
  NAND2_X1 U5302 ( .A1(n3268), .A2(n6556), .ZN(n4242) );
  NAND3_X1 U5303 ( .A1(n4242), .A2(n4241), .A3(n4681), .ZN(n4243) );
  OAI211_X1 U5304 ( .C1(n4540), .C2(n4244), .A(n4533), .B(n4243), .ZN(n4245)
         );
  NAND2_X1 U5305 ( .A1(n4245), .A2(n4545), .ZN(n4254) );
  INV_X1 U5306 ( .A(n4538), .ZN(n4249) );
  INV_X1 U5307 ( .A(n4265), .ZN(n4247) );
  OAI211_X1 U5308 ( .C1(n4246), .C2(n4249), .A(n4248), .B(n4247), .ZN(n4251)
         );
  NAND2_X1 U5309 ( .A1(n4251), .A2(n4250), .ZN(n4252) );
  INV_X1 U5310 ( .A(n6517), .ZN(n4255) );
  NOR2_X1 U5311 ( .A1(n4255), .A2(n4696), .ZN(n4505) );
  OAI22_X1 U5312 ( .A1(n4246), .A2(n4576), .B1(n4256), .B2(n4260), .ZN(n4257)
         );
  INV_X1 U5313 ( .A(n4257), .ZN(n4258) );
  NAND3_X1 U5314 ( .A1(n4505), .A2(n4258), .A3(n4105), .ZN(n4259) );
  XNOR2_X1 U5315 ( .A(n5256), .B(n5229), .ZN(n5416) );
  OAI21_X1 U5316 ( .B1(n4260), .B2(n4674), .A(n6527), .ZN(n4261) );
  NAND2_X1 U5317 ( .A1(n4016), .A2(n4262), .ZN(n4264) );
  INV_X1 U5318 ( .A(n4534), .ZN(n5391) );
  NAND2_X1 U5319 ( .A1(n5391), .A2(n4484), .ZN(n4263) );
  OAI211_X1 U5320 ( .C1(n4250), .C2(n4265), .A(n4264), .B(n4263), .ZN(n4266)
         );
  INV_X1 U5321 ( .A(n4266), .ZN(n4269) );
  NAND2_X1 U5322 ( .A1(n3266), .A2(n3245), .ZN(n4267) );
  AND4_X1 U5323 ( .A1(n4270), .A2(n4269), .A3(n4268), .A4(n4267), .ZN(n4271)
         );
  NAND2_X1 U5324 ( .A1(n4272), .A2(n4271), .ZN(n4524) );
  INV_X1 U5325 ( .A(n4273), .ZN(n4276) );
  INV_X1 U5326 ( .A(n4274), .ZN(n4275) );
  AOI22_X1 U5327 ( .A1(n3245), .A2(n4276), .B1(n4521), .B2(n4275), .ZN(n4278)
         );
  NAND2_X1 U5328 ( .A1(n4278), .A2(n4706), .ZN(n4279) );
  NAND2_X1 U5329 ( .A1(n4281), .A2(n4280), .ZN(n4698) );
  INV_X1 U5330 ( .A(n4698), .ZN(n4506) );
  NAND2_X2 U5331 ( .A1(n4292), .A2(n4506), .ZN(n4601) );
  INV_X2 U5332 ( .A(n6122), .ZN(n6095) );
  NOR2_X1 U5333 ( .A1(n6095), .A2(n4292), .ZN(n5785) );
  INV_X1 U5334 ( .A(n4281), .ZN(n4282) );
  NAND2_X1 U5335 ( .A1(n4292), .A2(n4282), .ZN(n5810) );
  AND2_X1 U5336 ( .A1(n4601), .A2(n5810), .ZN(n5811) );
  NOR2_X1 U5337 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5811), .ZN(n5782)
         );
  NOR2_X1 U5338 ( .A1(n5785), .A2(n5782), .ZN(n6160) );
  AND2_X1 U5339 ( .A1(n4601), .A2(n6160), .ZN(n5735) );
  INV_X1 U5340 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4283) );
  NAND2_X1 U5341 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5822) );
  NOR2_X1 U5342 ( .A1(n4283), .A2(n5822), .ZN(n5817) );
  AND2_X1 U5343 ( .A1(n5817), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5742)
         );
  NAND2_X1 U5344 ( .A1(n5742), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5745) );
  OR2_X1 U5345 ( .A1(n5745), .A2(n4284), .ZN(n5720) );
  INV_X1 U5346 ( .A(n5720), .ZN(n4285) );
  AOI21_X1 U5347 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n4598) );
  NOR2_X2 U5348 ( .A1(n4598), .A2(n4601), .ZN(n6133) );
  NOR2_X1 U5349 ( .A1(n4120), .A2(n4148), .ZN(n6132) );
  NAND2_X1 U5350 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6132), .ZN(n4893)
         );
  NOR2_X1 U5351 ( .A1(n4169), .A2(n4893), .ZN(n4288) );
  NAND2_X1 U5352 ( .A1(n6133), .A2(n4288), .ZN(n4931) );
  NOR2_X1 U5353 ( .A1(n4185), .A2(n4178), .ZN(n6130) );
  NAND3_X1 U5354 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n6130), .ZN(n4289) );
  NOR2_X2 U5355 ( .A1(n4931), .A2(n4289), .ZN(n5808) );
  NAND2_X1 U5356 ( .A1(n4285), .A2(n5808), .ZN(n5689) );
  NAND2_X1 U5357 ( .A1(n5699), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4286) );
  NOR2_X1 U5358 ( .A1(n5689), .A2(n4286), .ZN(n4287) );
  OR2_X1 U5359 ( .A1(n5735), .A2(n4287), .ZN(n4295) );
  INV_X1 U5360 ( .A(n4288), .ZN(n4928) );
  NAND2_X1 U5361 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4626) );
  OR2_X1 U5362 ( .A1(n4928), .A2(n4626), .ZN(n4932) );
  NOR2_X1 U5363 ( .A1(n4289), .A2(n4932), .ZN(n4297) );
  NOR2_X1 U5364 ( .A1(n5745), .A2(n5729), .ZN(n4290) );
  NAND2_X1 U5365 ( .A1(n4297), .A2(n4290), .ZN(n5691) );
  NAND3_X1 U5366 ( .A1(n5699), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4293) );
  NAND2_X1 U5367 ( .A1(n4292), .A2(n6499), .ZN(n5814) );
  OAI21_X1 U5368 ( .B1(n5691), .B2(n4293), .A(n5737), .ZN(n4294) );
  NAND2_X1 U5369 ( .A1(n4295), .A2(n4294), .ZN(n5681) );
  NOR2_X1 U5370 ( .A1(n6122), .A2(n6605), .ZN(n5521) );
  AOI21_X1 U5371 ( .B1(n5681), .B2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n5521), 
        .ZN(n4296) );
  OAI21_X1 U5372 ( .B1(n5416), .B2(n6149), .A(n4296), .ZN(n4301) );
  INV_X1 U5373 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6641) );
  NAND2_X1 U5374 ( .A1(n5814), .A2(n6641), .ZN(n6151) );
  INV_X1 U5375 ( .A(n4297), .ZN(n5736) );
  NOR2_X1 U5376 ( .A1(n5694), .A2(n5736), .ZN(n5766) );
  NOR2_X1 U5377 ( .A1(n5720), .A2(n5718), .ZN(n4298) );
  NAND2_X1 U5378 ( .A1(n5816), .A2(n4298), .ZN(n5716) );
  INV_X1 U5379 ( .A(n5716), .ZN(n5702) );
  NAND2_X1 U5380 ( .A1(n5702), .A2(n5699), .ZN(n5680) );
  NOR3_X1 U5381 ( .A1(n5680), .A2(n4299), .A3(n4422), .ZN(n4300) );
  INV_X1 U5382 ( .A(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n6170) );
  NOR4_X1 U5383 ( .A1(INSTQUEUE_REG_4__6__SCAN_IN), .A2(
        INSTQUEUE_REG_8__6__SCAN_IN), .A3(n4370), .A4(n6170), .ZN(n4306) );
  NOR4_X1 U5384 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(READY_N), .A3(
        INSTQUEUE_REG_7__2__SCAN_IN), .A4(n4367), .ZN(n4305) );
  NOR3_X1 U5385 ( .A1(INSTQUEUE_REG_4__2__SCAN_IN), .A2(FLUSH_REG_SCAN_IN), 
        .A3(DATAO_REG_19__SCAN_IN), .ZN(n4304) );
  NAND4_X1 U5386 ( .A1(n4306), .A2(n4305), .A3(DATAI_22_), .A4(n4304), .ZN(
        n4323) );
  NOR4_X1 U5387 ( .A1(DATAI_13_), .A2(DATAI_7_), .A3(LWORD_REG_13__SCAN_IN), 
        .A4(BS16_N), .ZN(n4310) );
  INV_X1 U5388 ( .A(LWORD_REG_7__SCAN_IN), .ZN(n6021) );
  NOR4_X1 U5389 ( .A1(EBX_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .A3(UWORD_REG_8__SCAN_IN), .A4(n6021), .ZN(n4309) );
  INV_X1 U5390 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4335) );
  NOR4_X1 U5391 ( .A1(ADDRESS_REG_11__SCAN_IN), .A2(DATAI_6_), .A3(
        DATAO_REG_6__SCAN_IN), .A4(n4335), .ZN(n4308) );
  NOR4_X1 U5392 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(
        ADDRESS_REG_17__SCAN_IN), .A3(n4333), .A4(n5484), .ZN(n4307) );
  NAND4_X1 U5393 ( .A1(n4310), .A2(n4309), .A3(n4308), .A4(n4307), .ZN(n4322)
         );
  NOR3_X1 U5394 ( .A1(EBX_REG_30__SCAN_IN), .A2(LWORD_REG_14__SCAN_IN), .A3(
        DATAO_REG_8__SCAN_IN), .ZN(n4313) );
  INV_X1 U5395 ( .A(EAX_REG_17__SCAN_IN), .ZN(n6041) );
  NOR4_X1 U5396 ( .A1(DATAO_REG_18__SCAN_IN), .A2(ADDRESS_REG_26__SCAN_IN), 
        .A3(DATAO_REG_30__SCAN_IN), .A4(n6041), .ZN(n4312) );
  INV_X1 U5397 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4531) );
  INV_X1 U5398 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6030) );
  NOR4_X1 U5399 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(n4476), .A3(n4531), 
        .A4(n6030), .ZN(n4311) );
  NAND4_X1 U5400 ( .A1(DATAO_REG_22__SCAN_IN), .A2(n4313), .A3(n4312), .A4(
        n4311), .ZN(n4321) );
  INV_X1 U5401 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4595) );
  INV_X1 U5402 ( .A(EBX_REG_2__SCAN_IN), .ZN(n5986) );
  NAND4_X1 U5403 ( .A1(EBX_REG_5__SCAN_IN), .A2(EBX_REG_6__SCAN_IN), .A3(n4595), .A4(n5986), .ZN(n4315) );
  NAND4_X1 U5404 ( .A1(EAX_REG_25__SCAN_IN), .A2(EAX_REG_1__SCAN_IN), .A3(
        REIP_REG_10__SCAN_IN), .A4(REIP_REG_21__SCAN_IN), .ZN(n4314) );
  OR4_X1 U5405 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(
        INSTQUEUE_REG_8__3__SCAN_IN), .A3(n4315), .A4(n4314), .ZN(n4319) );
  INV_X1 U5406 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n4399) );
  NAND4_X1 U5407 ( .A1(EAX_REG_12__SCAN_IN), .A2(ADDRESS_REG_23__SCAN_IN), 
        .A3(UWORD_REG_11__SCAN_IN), .A4(n4399), .ZN(n4318) );
  NOR2_X1 U5408 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n5845) );
  INV_X1 U5409 ( .A(n5845), .ZN(n4317) );
  INV_X1 U5410 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4369) );
  NAND4_X1 U5411 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(
        INSTQUEUE_REG_15__4__SCAN_IN), .A3(n4369), .A4(n6159), .ZN(n4316) );
  OR4_X1 U5412 ( .A1(n4319), .A2(n4318), .A3(n4317), .A4(n4316), .ZN(n4320) );
  NOR4_X1 U5413 ( .A1(n4323), .A2(n4322), .A3(n4321), .A4(n4320), .ZN(n4384)
         );
  INV_X1 U5414 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5978) );
  NOR4_X1 U5415 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(
        INSTQUEUE_REG_12__1__SCAN_IN), .A3(n4232), .A4(n5978), .ZN(n4383) );
  INV_X1 U5416 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n6019) );
  AOI22_X1 U5417 ( .A1(n6019), .A2(keyinput22), .B1(n5195), .B2(keyinput29), 
        .ZN(n4324) );
  OAI221_X1 U5418 ( .B1(n6019), .B2(keyinput22), .C1(n5195), .C2(keyinput29), 
        .A(n4324), .ZN(n4331) );
  INV_X1 U5419 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n5998) );
  AOI22_X1 U5420 ( .A1(n5998), .A2(keyinput44), .B1(n6041), .B2(keyinput7), 
        .ZN(n4325) );
  OAI221_X1 U5421 ( .B1(n5998), .B2(keyinput44), .C1(n6041), .C2(keyinput7), 
        .A(n4325), .ZN(n4330) );
  INV_X1 U5422 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n6614) );
  AOI22_X1 U5423 ( .A1(n4022), .A2(keyinput13), .B1(keyinput57), .B2(n6614), 
        .ZN(n4326) );
  OAI221_X1 U5424 ( .B1(n4022), .B2(keyinput13), .C1(n6614), .C2(keyinput57), 
        .A(n4326), .ZN(n4329) );
  INV_X1 U5425 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n6003) );
  AOI22_X1 U5426 ( .A1(n6159), .A2(keyinput14), .B1(keyinput19), .B2(n6003), 
        .ZN(n4327) );
  OAI221_X1 U5427 ( .B1(n6159), .B2(keyinput14), .C1(n6003), .C2(keyinput19), 
        .A(n4327), .ZN(n4328) );
  OR4_X1 U5428 ( .A1(n4331), .A2(n4330), .A3(n4329), .A4(n4328), .ZN(n4382) );
  AOI22_X1 U5429 ( .A1(n5484), .A2(keyinput17), .B1(keyinput8), .B2(n4333), 
        .ZN(n4332) );
  OAI221_X1 U5430 ( .B1(n5484), .B2(keyinput17), .C1(n4333), .C2(keyinput8), 
        .A(n4332), .ZN(n4340) );
  AOI22_X1 U5431 ( .A1(n4335), .A2(keyinput1), .B1(n3049), .B2(keyinput10), 
        .ZN(n4334) );
  OAI221_X1 U5432 ( .B1(n4335), .B2(keyinput1), .C1(n3049), .C2(keyinput10), 
        .A(n4334), .ZN(n4339) );
  INV_X1 U5433 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4337) );
  INV_X1 U5434 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5191) );
  AOI22_X1 U5435 ( .A1(n4337), .A2(keyinput45), .B1(keyinput56), .B2(n5191), 
        .ZN(n4336) );
  OAI221_X1 U5436 ( .B1(n4337), .B2(keyinput45), .C1(n5191), .C2(keyinput56), 
        .A(n4336), .ZN(n4338) );
  NOR3_X1 U5437 ( .A1(n4340), .A2(n4339), .A3(n4338), .ZN(n4343) );
  INV_X1 U5438 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n6597) );
  XOR2_X1 U5439 ( .A(keyinput31), .B(n6597), .Z(n4342) );
  INV_X1 U5440 ( .A(DATAWIDTH_REG_24__SCAN_IN), .ZN(n6547) );
  XOR2_X1 U5441 ( .A(keyinput46), .B(n6547), .Z(n4341) );
  NAND3_X1 U5442 ( .A1(n4343), .A2(n4342), .A3(n4341), .ZN(n4356) );
  INV_X1 U5443 ( .A(EAX_REG_25__SCAN_IN), .ZN(n6049) );
  INV_X1 U5444 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6032) );
  AOI22_X1 U5445 ( .A1(n6049), .A2(keyinput50), .B1(keyinput2), .B2(n6032), 
        .ZN(n4344) );
  OAI221_X1 U5446 ( .B1(n6049), .B2(keyinput50), .C1(n6032), .C2(keyinput2), 
        .A(n4344), .ZN(n4355) );
  INV_X1 U5447 ( .A(UWORD_REG_8__SCAN_IN), .ZN(n5996) );
  INV_X1 U5448 ( .A(DATAI_6_), .ZN(n6068) );
  AOI22_X1 U5449 ( .A1(n5996), .A2(keyinput48), .B1(keyinput37), .B2(n6068), 
        .ZN(n4345) );
  OAI221_X1 U5450 ( .B1(n5996), .B2(keyinput48), .C1(n6068), .C2(keyinput37), 
        .A(n4345), .ZN(n4354) );
  INV_X1 U5451 ( .A(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4347) );
  AOI22_X1 U5452 ( .A1(n4347), .A2(keyinput47), .B1(keyinput12), .B2(n6021), 
        .ZN(n4346) );
  OAI221_X1 U5453 ( .B1(n4347), .B2(keyinput47), .C1(n6021), .C2(keyinput12), 
        .A(n4346), .ZN(n4352) );
  INV_X1 U5454 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5638) );
  AOI22_X1 U5455 ( .A1(n5638), .A2(keyinput59), .B1(keyinput36), .B2(n4232), 
        .ZN(n4348) );
  OAI221_X1 U5456 ( .B1(n5638), .B2(keyinput59), .C1(n4232), .C2(keyinput36), 
        .A(n4348), .ZN(n4351) );
  XOR2_X1 U5457 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .B(keyinput3), .Z(n4350)
         );
  XOR2_X1 U5458 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .B(keyinput21), .Z(n4349)
         );
  OR4_X1 U5459 ( .A1(n4352), .A2(n4351), .A3(n4350), .A4(n4349), .ZN(n4353) );
  NOR4_X1 U5460 ( .A1(n4356), .A2(n4355), .A3(n4354), .A4(n4353), .ZN(n4380)
         );
  INV_X1 U5461 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n6586) );
  XOR2_X1 U5462 ( .A(keyinput28), .B(n6586), .Z(n4379) );
  INV_X1 U5463 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n4358) );
  INV_X1 U5464 ( .A(DATAWIDTH_REG_27__SCAN_IN), .ZN(n6546) );
  AOI22_X1 U5465 ( .A1(n4358), .A2(keyinput18), .B1(n6546), .B2(keyinput24), 
        .ZN(n4357) );
  OAI221_X1 U5466 ( .B1(n4358), .B2(keyinput18), .C1(n6546), .C2(keyinput24), 
        .A(n4357), .ZN(n4363) );
  XOR2_X1 U5467 ( .A(INSTQUEUE_REG_1__0__SCAN_IN), .B(keyinput49), .Z(n4362)
         );
  XOR2_X1 U5468 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .B(keyinput42), .Z(n4361)
         );
  XNOR2_X1 U5469 ( .A(keyinput23), .B(n4359), .ZN(n4360) );
  NOR4_X1 U5470 ( .A1(n4363), .A2(n4362), .A3(n4361), .A4(n4360), .ZN(n4378)
         );
  INV_X1 U5471 ( .A(LWORD_REG_14__SCAN_IN), .ZN(n6006) );
  INV_X1 U5472 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4365) );
  AOI22_X1 U5473 ( .A1(n6006), .A2(keyinput41), .B1(n4365), .B2(keyinput5), 
        .ZN(n4364) );
  OAI221_X1 U5474 ( .B1(n6006), .B2(keyinput41), .C1(n4365), .C2(keyinput5), 
        .A(n4364), .ZN(n4376) );
  AOI22_X1 U5475 ( .A1(n5986), .A2(keyinput6), .B1(n4367), .B2(keyinput53), 
        .ZN(n4366) );
  OAI221_X1 U5476 ( .B1(n5986), .B2(keyinput6), .C1(n4367), .C2(keyinput53), 
        .A(n4366), .ZN(n4375) );
  AOI22_X1 U5477 ( .A1(n4370), .A2(keyinput40), .B1(n4369), .B2(keyinput30), 
        .ZN(n4368) );
  OAI221_X1 U5478 ( .B1(n4370), .B2(keyinput40), .C1(n4369), .C2(keyinput30), 
        .A(n4368), .ZN(n4374) );
  INV_X1 U5479 ( .A(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4372) );
  AOI22_X1 U5480 ( .A1(n6603), .A2(keyinput52), .B1(n4372), .B2(keyinput33), 
        .ZN(n4371) );
  OAI221_X1 U5481 ( .B1(n6603), .B2(keyinput52), .C1(n4372), .C2(keyinput33), 
        .A(n4371), .ZN(n4373) );
  NOR4_X1 U5482 ( .A1(n4376), .A2(n4375), .A3(n4374), .A4(n4373), .ZN(n4377)
         );
  NAND4_X1 U5483 ( .A1(n4380), .A2(n4379), .A3(n4378), .A4(n4377), .ZN(n4381)
         );
  AOI211_X1 U5484 ( .C1(n4384), .C2(n4383), .A(n4382), .B(n4381), .ZN(n4418)
         );
  INV_X1 U5485 ( .A(UWORD_REG_11__SCAN_IN), .ZN(n4517) );
  INV_X1 U5486 ( .A(EBX_REG_5__SCAN_IN), .ZN(n5920) );
  AOI22_X1 U5487 ( .A1(n4517), .A2(keyinput54), .B1(n5920), .B2(keyinput51), 
        .ZN(n4385) );
  OAI221_X1 U5488 ( .B1(n4517), .B2(keyinput54), .C1(n5920), .C2(keyinput51), 
        .A(n4385), .ZN(n4394) );
  INV_X1 U5489 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6081) );
  INV_X1 U5490 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n6608) );
  AOI22_X1 U5491 ( .A1(n6081), .A2(keyinput4), .B1(keyinput15), .B2(n6608), 
        .ZN(n4386) );
  OAI221_X1 U5492 ( .B1(n6081), .B2(keyinput4), .C1(n6608), .C2(keyinput15), 
        .A(n4386), .ZN(n4393) );
  INV_X1 U5493 ( .A(LWORD_REG_13__SCAN_IN), .ZN(n4389) );
  INV_X1 U5494 ( .A(BS16_N), .ZN(n4388) );
  AOI22_X1 U5495 ( .A1(n4389), .A2(keyinput39), .B1(keyinput60), .B2(n4388), 
        .ZN(n4387) );
  OAI221_X1 U5496 ( .B1(n4389), .B2(keyinput39), .C1(n4388), .C2(keyinput60), 
        .A(n4387), .ZN(n4392) );
  INV_X1 U5497 ( .A(DATAI_13_), .ZN(n6084) );
  INV_X1 U5498 ( .A(DATAI_7_), .ZN(n6070) );
  AOI22_X1 U5499 ( .A1(n6084), .A2(keyinput34), .B1(keyinput55), .B2(n6070), 
        .ZN(n4390) );
  OAI221_X1 U5500 ( .B1(n6084), .B2(keyinput34), .C1(n6070), .C2(keyinput55), 
        .A(n4390), .ZN(n4391) );
  NOR4_X1 U5501 ( .A1(n4394), .A2(n4393), .A3(n4392), .A4(n4391), .ZN(n4417)
         );
  INV_X1 U5502 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n5994) );
  AOI22_X1 U5503 ( .A1(n5994), .A2(keyinput35), .B1(n4476), .B2(keyinput32), 
        .ZN(n4395) );
  OAI221_X1 U5504 ( .B1(n5994), .B2(keyinput35), .C1(n4476), .C2(keyinput32), 
        .A(n4395), .ZN(n4403) );
  INV_X1 U5505 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6552) );
  AOI22_X1 U5506 ( .A1(n6552), .A2(keyinput16), .B1(n4595), .B2(keyinput43), 
        .ZN(n4396) );
  OAI221_X1 U5507 ( .B1(n6552), .B2(keyinput16), .C1(n4595), .C2(keyinput43), 
        .A(n4396), .ZN(n4402) );
  AOI22_X1 U5508 ( .A1(n6170), .A2(keyinput11), .B1(keyinput26), .B2(n6030), 
        .ZN(n4397) );
  OAI221_X1 U5509 ( .B1(n6170), .B2(keyinput11), .C1(n6030), .C2(keyinput26), 
        .A(n4397), .ZN(n4401) );
  AOI22_X1 U5510 ( .A1(n4531), .A2(keyinput62), .B1(keyinput9), .B2(n4399), 
        .ZN(n4398) );
  OAI221_X1 U5511 ( .B1(n4531), .B2(keyinput62), .C1(n4399), .C2(keyinput9), 
        .A(n4398), .ZN(n4400) );
  NOR4_X1 U5512 ( .A1(n4403), .A2(n4402), .A3(n4401), .A4(n4400), .ZN(n4416)
         );
  INV_X1 U5513 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4405) );
  AOI22_X1 U5514 ( .A1(n4405), .A2(keyinput61), .B1(keyinput63), .B2(n6660), 
        .ZN(n4404) );
  OAI221_X1 U5515 ( .B1(n4405), .B2(keyinput61), .C1(n6660), .C2(keyinput63), 
        .A(n4404), .ZN(n4414) );
  INV_X1 U5516 ( .A(DATAI_22_), .ZN(n4407) );
  AOI22_X1 U5517 ( .A1(n4407), .A2(keyinput25), .B1(n5978), .B2(keyinput58), 
        .ZN(n4406) );
  OAI221_X1 U5518 ( .B1(n4407), .B2(keyinput25), .C1(n5978), .C2(keyinput58), 
        .A(n4406), .ZN(n4413) );
  INV_X1 U5519 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5842) );
  INV_X1 U5520 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4409) );
  AOI22_X1 U5521 ( .A1(n5842), .A2(keyinput27), .B1(n4409), .B2(keyinput0), 
        .ZN(n4408) );
  OAI221_X1 U5522 ( .B1(n5842), .B2(keyinput27), .C1(n4409), .C2(keyinput0), 
        .A(n4408), .ZN(n4412) );
  INV_X1 U5523 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n6000) );
  AOI22_X1 U5524 ( .A1(n6000), .A2(keyinput20), .B1(keyinput38), .B2(n6583), 
        .ZN(n4410) );
  OAI221_X1 U5525 ( .B1(n6000), .B2(keyinput20), .C1(n6583), .C2(keyinput38), 
        .A(n4410), .ZN(n4411) );
  NOR4_X1 U5526 ( .A1(n4414), .A2(n4413), .A3(n4412), .A4(n4411), .ZN(n4415)
         );
  NAND4_X1 U5527 ( .A1(n4418), .A2(n4417), .A3(n4416), .A4(n4415), .ZN(n4419)
         );
  XNOR2_X1 U5528 ( .A(n4420), .B(n4419), .ZN(U2996) );
  NOR2_X1 U5529 ( .A1(n5716), .A2(n4421), .ZN(n5657) );
  AND2_X1 U5530 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4427) );
  NAND2_X1 U5531 ( .A1(n5657), .A2(n4427), .ZN(n5630) );
  NOR3_X1 U5532 ( .A1(n5630), .A2(n5129), .A3(n4465), .ZN(n4430) );
  INV_X1 U5533 ( .A(n4601), .ZN(n5767) );
  INV_X1 U5534 ( .A(n4422), .ZN(n4423) );
  AND2_X1 U5535 ( .A1(n5696), .A2(n4423), .ZN(n4424) );
  OR2_X2 U5536 ( .A1(n4424), .A2(n5681), .ZN(n5674) );
  AOI21_X1 U5537 ( .B1(n5694), .B2(n4601), .A(n4425), .ZN(n4426) );
  INV_X1 U5538 ( .A(n4427), .ZN(n5644) );
  NAND2_X1 U5539 ( .A1(n5696), .A2(n5644), .ZN(n4428) );
  OAI21_X1 U5540 ( .B1(n5617), .B2(n6153), .A(n5636), .ZN(n5616) );
  AOI21_X1 U5541 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_29__SCAN_IN), .A(n6153), .ZN(n4429) );
  OR2_X1 U5542 ( .A1(n5616), .A2(n4429), .ZN(n5130) );
  MUX2_X1 U5543 ( .A(n4430), .B(n5130), .S(INSTADDRPOINTER_REG_31__SCAN_IN), 
        .Z(n4432) );
  AOI21_X1 U5544 ( .B1(n5409), .B2(n6138), .A(n3102), .ZN(n4433) );
  OAI21_X1 U5545 ( .B1(n4434), .B2(n6142), .A(n4433), .ZN(U2987) );
  OAI21_X2 U5546 ( .B1(n4097), .B2(n4099), .A(n4436), .ZN(n4437) );
  INV_X1 U5547 ( .A(n4437), .ZN(n4443) );
  AOI22_X1 U5548 ( .A1(n5467), .A2(DATAI_24_), .B1(n5473), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n4439) );
  NAND2_X1 U5549 ( .A1(n5468), .A2(DATAI_8_), .ZN(n4438) );
  OAI21_X1 U5550 ( .B1(n4437), .B2(n5477), .A(n3110), .ZN(U2867) );
  NOR2_X1 U5551 ( .A1(n5594), .A2(n5124), .ZN(n4442) );
  NAND2_X1 U5552 ( .A1(n6095), .A2(REIP_REG_24__SCAN_IN), .ZN(n5661) );
  OAI21_X1 U5553 ( .B1(n6112), .B2(n4440), .A(n5661), .ZN(n4441) );
  NAND3_X1 U5554 ( .A1(n2992), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4445) );
  NAND2_X1 U5555 ( .A1(n5526), .A2(n4444), .ZN(n5511) );
  NAND2_X1 U5556 ( .A1(n2992), .A2(n5729), .ZN(n5559) );
  NAND3_X1 U5557 ( .A1(n5550), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5559), .ZN(n5542) );
  INV_X1 U5558 ( .A(n5550), .ZN(n5561) );
  AOI21_X1 U5559 ( .B1(n5561), .B2(n4448), .A(n2992), .ZN(n4449) );
  NAND2_X1 U5560 ( .A1(n5707), .A2(n6107), .ZN(n4459) );
  BUF_X1 U5561 ( .A(n4453), .Z(n4454) );
  OAI21_X1 U5562 ( .B1(n4452), .B2(n4455), .A(n4454), .ZN(n5458) );
  OR2_X1 U5563 ( .A1(n5458), .A2(n5599), .ZN(n4458) );
  INV_X1 U5564 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6601) );
  NOR2_X1 U5565 ( .A1(n6122), .A2(n6601), .ZN(n5698) );
  NOR2_X1 U5566 ( .A1(n5594), .A2(n5274), .ZN(n4456) );
  AOI211_X1 U5567 ( .C1(n6094), .C2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n5698), 
        .B(n4456), .ZN(n4457) );
  NAND2_X1 U5568 ( .A1(n4459), .A2(n3112), .ZN(U2966) );
  NOR2_X1 U5569 ( .A1(n4473), .A2(n4460), .ZN(n5501) );
  NAND2_X1 U5570 ( .A1(n5587), .A2(n5647), .ZN(n5499) );
  NOR2_X1 U5571 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4461) );
  NAND2_X1 U5572 ( .A1(n4462), .A2(n4461), .ZN(n4463) );
  NOR2_X1 U5573 ( .A1(n5501), .A2(n4463), .ZN(n5481) );
  INV_X1 U5574 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5620) );
  NAND2_X1 U5575 ( .A1(n5481), .A2(n5620), .ZN(n4464) );
  INV_X1 U5576 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4467) );
  NAND2_X1 U5577 ( .A1(n6095), .A2(REIP_REG_30__SCAN_IN), .ZN(n5134) );
  OAI21_X1 U5578 ( .B1(n6112), .B2(n4467), .A(n5134), .ZN(n4468) );
  AOI21_X1 U5579 ( .B1(n4469), .B2(n6105), .A(n4468), .ZN(n4470) );
  INV_X1 U5580 ( .A(n4471), .ZN(n4472) );
  OAI21_X1 U5581 ( .B1(n5137), .B2(n6100), .A(n4472), .ZN(U2956) );
  AOI21_X1 U5582 ( .B1(n4475), .B2(n4474), .A(n4473), .ZN(n5660) );
  NOR2_X1 U5583 ( .A1(n5594), .A2(n5141), .ZN(n4478) );
  NAND2_X1 U5584 ( .A1(n6095), .A2(REIP_REG_25__SCAN_IN), .ZN(n5653) );
  OAI21_X1 U5585 ( .B1(n6112), .B2(n4476), .A(n5653), .ZN(n4477) );
  NOR2_X1 U5586 ( .A1(n4478), .A2(n4477), .ZN(n4479) );
  NAND4_X1 U5587 ( .A1(n4485), .A2(n2959), .A3(n4484), .A4(n4483), .ZN(n4486)
         );
  OAI21_X1 U5588 ( .B1(n4540), .B2(n4698), .A(n4486), .ZN(n4487) );
  NAND2_X2 U5589 ( .A1(n5987), .A2(n4661), .ZN(n5438) );
  NOR2_X1 U5590 ( .A1(n4489), .A2(n4490), .ZN(n4491) );
  OR2_X1 U5591 ( .A1(n4488), .A2(n4491), .ZN(n5652) );
  INV_X1 U5592 ( .A(EBX_REG_25__SCAN_IN), .ZN(n4492) );
  AND2_X1 U5593 ( .A1(n6380), .A2(n4725), .ZN(n5289) );
  INV_X1 U5594 ( .A(n5289), .ZN(n4497) );
  NAND2_X1 U5595 ( .A1(n4513), .A2(n4497), .ZN(n5801) );
  NOR2_X1 U5596 ( .A1(n5801), .A2(READREQUEST_REG_SCAN_IN), .ZN(n4498) );
  AND2_X1 U5597 ( .A1(n4498), .A2(n5802), .ZN(n4499) );
  OR2_X1 U5598 ( .A1(n2984), .A2(n5391), .ZN(n4504) );
  OAI22_X1 U5599 ( .A1(n4499), .A2(n4504), .B1(n4498), .B2(n6658), .ZN(U3474)
         );
  OR2_X1 U5600 ( .A1(n4540), .A2(n3227), .ZN(n4503) );
  INV_X1 U5601 ( .A(n4500), .ZN(n4501) );
  NAND2_X1 U5602 ( .A1(n4501), .A2(n3963), .ZN(n4502) );
  NAND2_X1 U5603 ( .A1(n4503), .A2(n4502), .ZN(n5837) );
  AOI21_X1 U5604 ( .B1(n4504), .B2(n6556), .A(READY_N), .ZN(n6661) );
  NOR2_X1 U5605 ( .A1(n5837), .A2(n6661), .ZN(n6515) );
  OR2_X1 U5606 ( .A1(n6515), .A2(n6537), .ZN(n4510) );
  INV_X1 U5607 ( .A(n4510), .ZN(n5843) );
  INV_X1 U5608 ( .A(MORE_REG_SCAN_IN), .ZN(n4512) );
  NAND2_X1 U5609 ( .A1(n4505), .A2(n3963), .ZN(n4507) );
  MUX2_X1 U5610 ( .A(n4507), .B(n4506), .S(n4540), .Z(n4508) );
  AOI21_X1 U5611 ( .B1(n3964), .B2(n4509), .A(n4508), .ZN(n6518) );
  OR2_X1 U5612 ( .A1(n6518), .A2(n4510), .ZN(n4511) );
  OAI21_X1 U5613 ( .B1(n5843), .B2(n4512), .A(n4511), .ZN(U3471) );
  INV_X1 U5614 ( .A(DATAI_8_), .ZN(n4516) );
  INV_X1 U5615 ( .A(n4513), .ZN(n4514) );
  OAI222_X1 U5616 ( .A1(n4516), .A2(n6083), .B1(n6037), .B2(n5996), .C1(n4515), 
        .C2(n6092), .ZN(U2932) );
  INV_X1 U5617 ( .A(DATAI_11_), .ZN(n4518) );
  OAI222_X1 U5618 ( .A1(n4518), .A2(n6083), .B1(n6037), .B2(n4517), .C1(n4553), 
        .C2(n6092), .ZN(U2935) );
  INV_X1 U5619 ( .A(n4520), .ZN(n5963) );
  INV_X1 U5620 ( .A(n4521), .ZN(n4522) );
  NAND4_X1 U5621 ( .A1(n4523), .A2(n4105), .A3(n4246), .A4(n4522), .ZN(n4525)
         );
  NOR2_X1 U5622 ( .A1(n4525), .A2(n4524), .ZN(n6493) );
  AOI21_X1 U5623 ( .B1(n6499), .B2(n4529), .A(n4528), .ZN(n4530) );
  OAI21_X1 U5624 ( .B1(n5963), .B2(n6493), .A(n4530), .ZN(n6502) );
  INV_X1 U5625 ( .A(n6647), .ZN(n6635) );
  AOI22_X1 U5626 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4531), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6159), .ZN(n5156) );
  NOR2_X1 U5627 ( .A1(n4725), .A2(n6641), .ZN(n5154) );
  INV_X1 U5628 ( .A(n6531), .ZN(n6634) );
  AOI222_X1 U5629 ( .A1(n6502), .A2(n6635), .B1(n5156), .B2(n5154), .C1(n4532), 
        .C2(n6634), .ZN(n4547) );
  OAI21_X1 U5630 ( .B1(n4534), .B2(n4681), .A(n4533), .ZN(n4535) );
  NOR2_X1 U5631 ( .A1(n4536), .A2(n4535), .ZN(n4543) );
  NAND2_X1 U5632 ( .A1(n3963), .A2(n4537), .ZN(n4539) );
  OAI211_X1 U5633 ( .C1(n6499), .C2(n2987), .A(n4539), .B(n4538), .ZN(n4541)
         );
  MUX2_X1 U5634 ( .A(n4698), .B(n4541), .S(n4540), .Z(n4542) );
  NAND2_X1 U5635 ( .A1(n4543), .A2(n4542), .ZN(n6501) );
  NAND2_X1 U5636 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4735), .ZN(n6630) );
  NOR2_X1 U5637 ( .A1(n6630), .A2(n5842), .ZN(n4544) );
  AOI21_X1 U5638 ( .B1(n6501), .B2(n4545), .A(n4544), .ZN(n5835) );
  NAND2_X1 U5639 ( .A1(n6530), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6631) );
  NAND2_X1 U5640 ( .A1(n5835), .A2(n6631), .ZN(n6645) );
  INV_X1 U5641 ( .A(n6645), .ZN(n5162) );
  NOR2_X1 U5642 ( .A1(n6531), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6640)
         );
  OAI21_X1 U5643 ( .B1(n5162), .B2(n6640), .A(n2983), .ZN(n4546) );
  OAI21_X1 U5644 ( .B1(n4547), .B2(n5162), .A(n4546), .ZN(U3460) );
  INV_X1 U5645 ( .A(n6499), .ZN(n4700) );
  INV_X1 U5646 ( .A(n6556), .ZN(n4550) );
  NAND2_X1 U5647 ( .A1(n4735), .A2(n6530), .ZN(n6523) );
  INV_X2 U5648 ( .A(n6523), .ZN(n6016) );
  NOR2_X4 U5649 ( .A1(n6022), .A2(n6016), .ZN(n6033) );
  AOI22_X1 U5650 ( .A1(UWORD_REG_11__SCAN_IN), .A2(n6016), .B1(n6033), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4552) );
  OAI21_X1 U5651 ( .B1(n4553), .B2(n5992), .A(n4552), .ZN(U2896) );
  AOI22_X1 U5652 ( .A1(n6016), .A2(UWORD_REG_9__SCAN_IN), .B1(n6033), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4554) );
  OAI21_X1 U5653 ( .B1(n6049), .B2(n5992), .A(n4554), .ZN(U2898) );
  INV_X1 U5654 ( .A(EAX_REG_16__SCAN_IN), .ZN(n6039) );
  AOI22_X1 U5655 ( .A1(n6016), .A2(UWORD_REG_0__SCAN_IN), .B1(n6033), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4555) );
  OAI21_X1 U5656 ( .B1(n6039), .B2(n5992), .A(n4555), .ZN(U2907) );
  AOI22_X1 U5657 ( .A1(n6016), .A2(UWORD_REG_1__SCAN_IN), .B1(n6033), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4556) );
  OAI21_X1 U5658 ( .B1(n6041), .B2(n5992), .A(n4556), .ZN(U2906) );
  AOI22_X1 U5659 ( .A1(n6016), .A2(UWORD_REG_5__SCAN_IN), .B1(n6033), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4557) );
  OAI21_X1 U5660 ( .B1(n3709), .B2(n5992), .A(n4557), .ZN(U2902) );
  AOI22_X1 U5661 ( .A1(n6016), .A2(UWORD_REG_12__SCAN_IN), .B1(n6033), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4558) );
  OAI21_X1 U5662 ( .B1(n3850), .B2(n5992), .A(n4558), .ZN(U2895) );
  INV_X1 U5663 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4560) );
  AOI22_X1 U5664 ( .A1(n6016), .A2(UWORD_REG_7__SCAN_IN), .B1(n6033), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4559) );
  OAI21_X1 U5665 ( .B1(n4560), .B2(n5992), .A(n4559), .ZN(U2900) );
  INV_X1 U5666 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4562) );
  AOI22_X1 U5667 ( .A1(n6016), .A2(UWORD_REG_4__SCAN_IN), .B1(n6033), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4561) );
  OAI21_X1 U5668 ( .B1(n4562), .B2(n5992), .A(n4561), .ZN(U2903) );
  AOI22_X1 U5669 ( .A1(n6016), .A2(UWORD_REG_10__SCAN_IN), .B1(n6033), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4563) );
  OAI21_X1 U5670 ( .B1(n3804), .B2(n5992), .A(n4563), .ZN(U2897) );
  INV_X1 U5671 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4565) );
  AOI22_X1 U5672 ( .A1(n6016), .A2(UWORD_REG_13__SCAN_IN), .B1(n6033), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4564) );
  OAI21_X1 U5673 ( .B1(n4565), .B2(n5992), .A(n4564), .ZN(U2894) );
  OAI21_X1 U5674 ( .B1(n4568), .B2(n4567), .A(n4566), .ZN(n5608) );
  NOR2_X1 U5675 ( .A1(n4016), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4570)
         );
  OR2_X1 U5676 ( .A1(n4570), .A2(n4569), .ZN(n5780) );
  OAI222_X1 U5677 ( .A1(n5608), .A2(n5438), .B1(n4006), .B2(n5987), .C1(n5780), 
        .C2(n5433), .ZN(U2859) );
  OR2_X1 U5678 ( .A1(n4572), .A2(n4571), .ZN(n4574) );
  NAND2_X1 U5679 ( .A1(n4574), .A2(n4573), .ZN(n5962) );
  XNOR2_X1 U5680 ( .A(n4575), .B(n4576), .ZN(n6148) );
  OAI222_X1 U5681 ( .A1(n5962), .A2(n5438), .B1(n4577), .B2(n5987), .C1(n5433), 
        .C2(n6148), .ZN(U2858) );
  NOR2_X1 U5682 ( .A1(n4580), .A2(n4579), .ZN(n4581) );
  OR2_X1 U5683 ( .A1(n4578), .A2(n4581), .ZN(n5983) );
  INV_X1 U5684 ( .A(n5467), .ZN(n4583) );
  INV_X1 U5685 ( .A(n5468), .ZN(n4582) );
  AOI22_X1 U5686 ( .A1(n5988), .A2(DATAI_2_), .B1(EAX_REG_2__SCAN_IN), .B2(
        n5473), .ZN(n4584) );
  OAI21_X1 U5687 ( .B1(n5983), .B2(n5477), .A(n4584), .ZN(U2889) );
  OAI21_X1 U5688 ( .B1(n4578), .B2(n4586), .A(n4749), .ZN(n5945) );
  OAI21_X1 U5689 ( .B1(n4587), .B2(n4589), .A(n4588), .ZN(n5951) );
  INV_X1 U5690 ( .A(n5951), .ZN(n4590) );
  INV_X1 U5691 ( .A(n5987), .ZN(n5436) );
  AOI22_X1 U5692 ( .A1(n5979), .A2(n4590), .B1(EBX_REG_3__SCAN_IN), .B2(n5436), 
        .ZN(n4591) );
  OAI21_X1 U5693 ( .B1(n5945), .B2(n5438), .A(n4591), .ZN(U2856) );
  XOR2_X1 U5694 ( .A(n4592), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n4594) );
  XNOR2_X1 U5695 ( .A(n4594), .B(n4593), .ZN(n4614) );
  NAND2_X1 U5696 ( .A1(n5737), .A2(n4626), .ZN(n4625) );
  OAI21_X1 U5697 ( .B1(n5767), .B2(n6160), .A(n4625), .ZN(n4597) );
  NOR2_X1 U5698 ( .A1(n5694), .A2(n6159), .ZN(n4596) );
  MUX2_X1 U5699 ( .A(n4597), .B(n4596), .S(n4595), .Z(n4607) );
  NOR2_X1 U5700 ( .A1(n6641), .A2(n6159), .ZN(n4599) );
  AOI21_X1 U5701 ( .B1(n4599), .B2(INSTADDRPOINTER_REG_2__SCAN_IN), .A(n4598), 
        .ZN(n4600) );
  NOR2_X1 U5702 ( .A1(n4601), .A2(n4600), .ZN(n4606) );
  NOR2_X1 U5703 ( .A1(n4602), .A2(n4603), .ZN(n4604) );
  OR2_X1 U5704 ( .A1(n4587), .A2(n4604), .ZN(n5982) );
  INV_X1 U5705 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6568) );
  OAI22_X1 U5706 ( .A1(n6149), .A2(n5982), .B1(n6568), .B2(n6122), .ZN(n4605)
         );
  NOR3_X1 U5707 ( .A1(n4607), .A2(n4606), .A3(n4605), .ZN(n4608) );
  OAI21_X1 U5708 ( .B1(n6142), .B2(n4614), .A(n4608), .ZN(U3016) );
  INV_X1 U5709 ( .A(DATAI_0_), .ZN(n6056) );
  INV_X1 U5710 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6036) );
  OAI222_X1 U5711 ( .A1(n5608), .A2(n5477), .B1(n5476), .B2(n6056), .C1(n5991), 
        .C2(n6036), .ZN(U2891) );
  INV_X1 U5712 ( .A(DATAI_1_), .ZN(n6058) );
  OAI222_X1 U5713 ( .A1(n5962), .A2(n5477), .B1(n5476), .B2(n6058), .C1(n5991), 
        .C2(n6032), .ZN(U2890) );
  INV_X1 U5714 ( .A(DATAI_3_), .ZN(n6062) );
  INV_X1 U5715 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6028) );
  OAI222_X1 U5716 ( .A1(n5945), .A2(n5477), .B1(n5476), .B2(n6062), .C1(n5991), 
        .C2(n6028), .ZN(U2888) );
  INV_X1 U5717 ( .A(n5983), .ZN(n4612) );
  NOR2_X1 U5718 ( .A1(n5594), .A2(n5393), .ZN(n4611) );
  INV_X1 U5719 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n4609) );
  OAI22_X1 U5720 ( .A1(n6112), .A2(n4609), .B1(n6122), .B2(n6568), .ZN(n4610)
         );
  AOI211_X1 U5721 ( .C1(n4612), .C2(n6104), .A(n4611), .B(n4610), .ZN(n4613)
         );
  OAI21_X1 U5722 ( .B1(n6100), .B2(n4614), .A(n4613), .ZN(U2984) );
  OAI21_X1 U5723 ( .B1(n4617), .B2(n4616), .A(n4615), .ZN(n4618) );
  INV_X1 U5724 ( .A(n4618), .ZN(n6156) );
  INV_X1 U5725 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4620) );
  NAND2_X1 U5726 ( .A1(n6105), .A2(n4620), .ZN(n4619) );
  NAND2_X1 U5727 ( .A1(n6095), .A2(REIP_REG_1__SCAN_IN), .ZN(n6147) );
  OAI211_X1 U5728 ( .C1(n6112), .C2(n4620), .A(n4619), .B(n6147), .ZN(n4621)
         );
  AOI21_X1 U5729 ( .B1(n6156), .B2(n6107), .A(n4621), .ZN(n4622) );
  OAI21_X1 U5730 ( .B1(n5599), .B2(n5962), .A(n4622), .ZN(U2985) );
  XNOR2_X1 U5731 ( .A(n4623), .B(n4624), .ZN(n4756) );
  OAI21_X1 U5732 ( .B1(n6133), .B2(n5735), .A(n4625), .ZN(n4892) );
  NOR2_X1 U5733 ( .A1(n4626), .A2(n5694), .ZN(n6131) );
  NOR2_X1 U5734 ( .A1(n6133), .A2(n6131), .ZN(n4929) );
  AOI211_X1 U5735 ( .C1(n4120), .C2(n4148), .A(n4929), .B(n6132), .ZN(n4627)
         );
  AOI21_X1 U5736 ( .B1(INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n4892), .A(n4627), 
        .ZN(n4632) );
  INV_X1 U5737 ( .A(n4628), .ZN(n4629) );
  AOI21_X1 U5738 ( .B1(n4630), .B2(n4588), .A(n4629), .ZN(n5926) );
  NOR2_X1 U5739 ( .A1(n6122), .A2(n6572), .ZN(n4752) );
  AOI21_X1 U5740 ( .B1(n5926), .B2(n6138), .A(n4752), .ZN(n4631) );
  OAI211_X1 U5741 ( .C1(n6142), .C2(n4756), .A(n4632), .B(n4631), .ZN(U3014)
         );
  XOR2_X1 U5742 ( .A(n4634), .B(n4633), .Z(n4639) );
  NAND2_X1 U5743 ( .A1(n6095), .A2(REIP_REG_3__SCAN_IN), .ZN(n4640) );
  OAI21_X1 U5744 ( .B1(n6149), .B2(n5951), .A(n4640), .ZN(n4637) );
  INV_X1 U5745 ( .A(n4929), .ZN(n4635) );
  MUX2_X1 U5746 ( .A(n4635), .B(n4892), .S(INSTADDRPOINTER_REG_3__SCAN_IN), 
        .Z(n4636) );
  AOI211_X1 U5747 ( .C1(n6155), .C2(n4639), .A(n4637), .B(n4636), .ZN(n4638)
         );
  INV_X1 U5748 ( .A(n4638), .ZN(U3015) );
  NAND2_X1 U5749 ( .A1(n4639), .A2(n6107), .ZN(n4644) );
  INV_X1 U5750 ( .A(n4640), .ZN(n4642) );
  NOR2_X1 U5751 ( .A1(n5594), .A2(n5946), .ZN(n4641) );
  AOI211_X1 U5752 ( .C1(n6094), .C2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n4642), 
        .B(n4641), .ZN(n4643) );
  OAI211_X1 U5753 ( .C1(n5599), .C2(n5945), .A(n4644), .B(n4643), .ZN(U2983)
         );
  AND2_X1 U5754 ( .A1(n4645), .A2(n6495), .ZN(n6339) );
  INV_X1 U5755 ( .A(n4691), .ZN(n4648) );
  AOI21_X1 U5756 ( .B1(n6339), .B2(n6274), .A(n4648), .ZN(n4656) );
  INV_X1 U5757 ( .A(n4656), .ZN(n4650) );
  AOI22_X1 U5758 ( .A1(n4650), .A2(n6380), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4649), .ZN(n4695) );
  AOI21_X1 U5759 ( .B1(n6378), .B2(STATE2_REG_3__SCAN_IN), .A(n6312), .ZN(
        n6240) );
  AND2_X1 U5760 ( .A1(n4652), .A2(n4771), .ZN(n4654) );
  NAND2_X1 U5761 ( .A1(n6380), .A2(n6432), .ZN(n6208) );
  OAI21_X1 U5762 ( .B1(n4662), .B2(n5599), .A(n6208), .ZN(n4655) );
  AOI22_X1 U5763 ( .A1(n4656), .A2(n4655), .B1(n4850), .B2(n6435), .ZN(n4657)
         );
  NAND2_X1 U5764 ( .A1(n6240), .A2(n4657), .ZN(n4689) );
  NAND2_X1 U5765 ( .A1(n4689), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4665)
         );
  INV_X1 U5766 ( .A(n6631), .ZN(n4660) );
  NAND2_X1 U5767 ( .A1(n4660), .A2(n4659), .ZN(n4670) );
  NAND2_X1 U5768 ( .A1(n4690), .A2(n4661), .ZN(n5084) );
  INV_X1 U5769 ( .A(n6487), .ZN(n6424) );
  OAI22_X1 U5770 ( .A1(n5084), .A2(n4691), .B1(n6424), .B2(n4834), .ZN(n4663)
         );
  AOI21_X1 U5771 ( .B1(n6419), .B2(n4882), .A(n4663), .ZN(n4664) );
  OAI211_X1 U5772 ( .C1(n4695), .C2(n6374), .A(n4665), .B(n4664), .ZN(U3147)
         );
  NAND2_X1 U5773 ( .A1(n4689), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4668)
         );
  NAND2_X1 U5774 ( .A1(n6104), .A2(DATAI_27_), .ZN(n6463) );
  NAND2_X1 U5775 ( .A1(n4690), .A2(n3243), .ZN(n5094) );
  INV_X1 U5776 ( .A(n6460), .ZN(n6404) );
  OAI22_X1 U5777 ( .A1(n5094), .A2(n4691), .B1(n6404), .B2(n4834), .ZN(n4666)
         );
  AOI21_X1 U5778 ( .B1(n6401), .B2(n4882), .A(n4666), .ZN(n4667) );
  OAI211_X1 U5779 ( .C1(n4695), .C2(n6358), .A(n4668), .B(n4667), .ZN(U3143)
         );
  NAND2_X1 U5780 ( .A1(n4689), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4673)
         );
  NOR2_X2 U5781 ( .A1(n4670), .A2(n4669), .ZN(n6430) );
  INV_X1 U5782 ( .A(n6430), .ZN(n4947) );
  INV_X1 U5783 ( .A(n6442), .ZN(n6392) );
  OAI22_X1 U5784 ( .A1(n4947), .A2(n4691), .B1(n6392), .B2(n4834), .ZN(n4671)
         );
  AOI21_X1 U5785 ( .B1(n6379), .B2(n4882), .A(n4671), .ZN(n4672) );
  OAI211_X1 U5786 ( .C1(n4695), .C2(n6348), .A(n4673), .B(n4672), .ZN(U3140)
         );
  NAND2_X1 U5787 ( .A1(n4689), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4677)
         );
  NAND2_X1 U5788 ( .A1(n4690), .A2(n4674), .ZN(n5105) );
  INV_X1 U5789 ( .A(n6466), .ZN(n6408) );
  OAI22_X1 U5790 ( .A1(n5105), .A2(n4691), .B1(n6408), .B2(n4834), .ZN(n4675)
         );
  AOI21_X1 U5791 ( .B1(n6405), .B2(n4882), .A(n4675), .ZN(n4676) );
  OAI211_X1 U5792 ( .C1(n4695), .C2(n6361), .A(n4677), .B(n4676), .ZN(U3144)
         );
  NAND2_X1 U5793 ( .A1(n4689), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4680)
         );
  NAND2_X1 U5794 ( .A1(n4690), .A2(n2985), .ZN(n5089) );
  INV_X1 U5795 ( .A(n6472), .ZN(n6412) );
  OAI22_X1 U5796 ( .A1(n5089), .A2(n4691), .B1(n6412), .B2(n4834), .ZN(n4678)
         );
  AOI21_X1 U5797 ( .B1(n6409), .B2(n4882), .A(n4678), .ZN(n4679) );
  OAI211_X1 U5798 ( .C1(n4695), .C2(n6364), .A(n4680), .B(n4679), .ZN(U3145)
         );
  NAND2_X1 U5799 ( .A1(n4689), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4684)
         );
  NAND2_X1 U5800 ( .A1(n4690), .A2(n4681), .ZN(n5068) );
  INV_X1 U5801 ( .A(n6454), .ZN(n5076) );
  OAI22_X1 U5802 ( .A1(n5068), .A2(n4691), .B1(n5076), .B2(n4834), .ZN(n4682)
         );
  AOI21_X1 U5803 ( .B1(n6352), .B2(n4882), .A(n4682), .ZN(n4683) );
  OAI211_X1 U5804 ( .C1(n4695), .C2(n6355), .A(n4684), .B(n4683), .ZN(U3142)
         );
  NAND2_X1 U5805 ( .A1(n4689), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4688)
         );
  NAND2_X1 U5806 ( .A1(n6104), .A2(DATAI_30_), .ZN(n6481) );
  NAND2_X1 U5807 ( .A1(n4690), .A2(n4685), .ZN(n5099) );
  INV_X1 U5808 ( .A(n6478), .ZN(n6416) );
  OAI22_X1 U5809 ( .A1(n5099), .A2(n4691), .B1(n6416), .B2(n4834), .ZN(n4686)
         );
  AOI21_X1 U5810 ( .B1(n6413), .B2(n4882), .A(n4686), .ZN(n4687) );
  OAI211_X1 U5811 ( .C1(n4695), .C2(n6367), .A(n4688), .B(n4687), .ZN(U3146)
         );
  NAND2_X1 U5812 ( .A1(n4689), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4694)
         );
  NAND2_X1 U5813 ( .A1(n4690), .A2(n3268), .ZN(n5079) );
  INV_X1 U5814 ( .A(n6448), .ZN(n6396) );
  OAI22_X1 U5815 ( .A1(n5079), .A2(n4691), .B1(n6396), .B2(n4834), .ZN(n4692)
         );
  AOI21_X1 U5816 ( .B1(n6393), .B2(n4882), .A(n4692), .ZN(n4693) );
  OAI211_X1 U5817 ( .C1(n4695), .C2(n6351), .A(n4694), .B(n4693), .ZN(U3141)
         );
  INV_X1 U5818 ( .A(n4696), .ZN(n4697) );
  NAND2_X1 U5819 ( .A1(n4698), .A2(n4697), .ZN(n4716) );
  NAND2_X1 U5820 ( .A1(n5160), .A2(n3425), .ZN(n4713) );
  NAND2_X1 U5821 ( .A1(n4713), .A2(n4707), .ZN(n4703) );
  XNOR2_X1 U5822 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n2983), .ZN(n4699)
         );
  OAI22_X1 U5823 ( .A1(n4700), .A2(n4699), .B1(n4706), .B2(n4703), .ZN(n4702)
         );
  INV_X1 U5824 ( .A(n4647), .ZN(n5795) );
  NOR2_X1 U5825 ( .A1(n5795), .A2(n6493), .ZN(n4701) );
  AOI211_X1 U5826 ( .C1(n4716), .C2(n4703), .A(n4702), .B(n4701), .ZN(n5153)
         );
  MUX2_X1 U5827 ( .A(n3425), .B(n5153), .S(n6501), .Z(n6507) );
  NOR2_X1 U5828 ( .A1(n6507), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4721) );
  INV_X1 U5829 ( .A(n4645), .ZN(n5950) );
  NAND2_X1 U5830 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4704) );
  INV_X1 U5831 ( .A(n4704), .ZN(n4705) );
  MUX2_X1 U5832 ( .A(n4705), .B(n4704), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4712) );
  INV_X1 U5833 ( .A(n4706), .ZN(n4711) );
  INV_X1 U5834 ( .A(n4707), .ZN(n4710) );
  OAI21_X1 U5835 ( .B1(n4710), .B2(n4709), .A(n4708), .ZN(n6633) );
  AOI22_X1 U5836 ( .A1(n6499), .A2(n4712), .B1(n4711), .B2(n6633), .ZN(n4718)
         );
  INV_X1 U5837 ( .A(n4713), .ZN(n4714) );
  XNOR2_X1 U5838 ( .A(n4714), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4715)
         );
  NAND2_X1 U5839 ( .A1(n4716), .A2(n4715), .ZN(n4717) );
  OAI211_X1 U5840 ( .C1(n5950), .C2(n6493), .A(n4718), .B(n4717), .ZN(n6636)
         );
  MUX2_X1 U5841 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6636), .S(n6501), 
        .Z(n6508) );
  AND2_X1 U5842 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5842), .ZN(n4719) );
  AOI22_X1 U5843 ( .A1(n4721), .A2(n6508), .B1(n4720), .B2(n4719), .ZN(n6514)
         );
  NOR2_X1 U5844 ( .A1(n6514), .A2(n4526), .ZN(n4737) );
  MUX2_X1 U5845 ( .A(FLUSH_REG_SCAN_IN), .B(n6501), .S(n4725), .Z(n4727) );
  INV_X1 U5846 ( .A(n6436), .ZN(n6207) );
  NOR2_X1 U5847 ( .A1(n2988), .A2(n6207), .ZN(n4724) );
  XNOR2_X1 U5848 ( .A(n4724), .B(n4723), .ZN(n5930) );
  NAND3_X1 U5849 ( .A1(n5930), .A2(n4726), .A3(n4725), .ZN(n5832) );
  OAI21_X1 U5850 ( .B1(n4723), .B2(n4727), .A(n5832), .ZN(n6521) );
  NOR3_X1 U5851 ( .A1(n4737), .A2(n6521), .A3(FLUSH_REG_SCAN_IN), .ZN(n4728)
         );
  NAND2_X1 U5852 ( .A1(n4652), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6381) );
  MUX2_X1 U5853 ( .A(n4652), .B(n6381), .S(n2989), .Z(n4730) );
  OAI21_X1 U5854 ( .B1(n5793), .B2(n4730), .A(n6382), .ZN(n4731) );
  NAND2_X1 U5855 ( .A1(n4731), .A2(n6380), .ZN(n6174) );
  INV_X1 U5856 ( .A(n6174), .ZN(n4733) );
  AND2_X1 U5857 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n3238), .ZN(n5794) );
  OAI22_X1 U5858 ( .A1(n4729), .A2(n6208), .B1(n5950), .B2(n5794), .ZN(n4732)
         );
  OAI21_X1 U5859 ( .B1(n4733), .B2(n4732), .A(n6161), .ZN(n4734) );
  OAI21_X1 U5860 ( .B1(n6161), .B2(n6509), .A(n4734), .ZN(U3462) );
  INV_X1 U5861 ( .A(n4735), .ZN(n4736) );
  NOR3_X1 U5862 ( .A1(n4737), .A2(n6521), .A3(n4736), .ZN(n6529) );
  INV_X1 U5863 ( .A(n6495), .ZN(n4759) );
  OAI22_X1 U5864 ( .A1(n5062), .A2(n6435), .B1(n4759), .B2(n5794), .ZN(n4738)
         );
  OAI21_X1 U5865 ( .B1(n6529), .B2(n4738), .A(n6161), .ZN(n4739) );
  OAI21_X1 U5866 ( .B1(n6161), .B2(n6378), .A(n4739), .ZN(U3465) );
  AND2_X1 U5867 ( .A1(n4740), .A2(n4741), .ZN(n4743) );
  OR2_X1 U5868 ( .A1(n4743), .A2(n4742), .ZN(n4846) );
  INV_X1 U5869 ( .A(DATAI_5_), .ZN(n6066) );
  OAI222_X1 U5870 ( .A1(n4846), .A2(n5477), .B1(n5476), .B2(n6066), .C1(n5991), 
        .C2(n3454), .ZN(U2886) );
  AND2_X1 U5871 ( .A1(n4628), .A2(n4745), .ZN(n4746) );
  NOR2_X1 U5872 ( .A1(n4744), .A2(n4746), .ZN(n6139) );
  INV_X1 U5873 ( .A(n6139), .ZN(n4747) );
  OAI222_X1 U5874 ( .A1(n4846), .A2(n5438), .B1(n5987), .B2(n5920), .C1(n4747), 
        .C2(n5433), .ZN(U2854) );
  INV_X1 U5875 ( .A(n4740), .ZN(n4748) );
  AOI21_X1 U5876 ( .B1(n4750), .B2(n4749), .A(n4748), .ZN(n5936) );
  INV_X1 U5877 ( .A(n5936), .ZN(n4757) );
  AOI22_X1 U5878 ( .A1(n5926), .A2(n5979), .B1(EBX_REG_4__SCAN_IN), .B2(n5436), 
        .ZN(n4751) );
  OAI21_X1 U5879 ( .B1(n4757), .B2(n5438), .A(n4751), .ZN(U2855) );
  AOI21_X1 U5880 ( .B1(n6094), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n4752), 
        .ZN(n4753) );
  OAI21_X1 U5881 ( .B1(n5934), .B2(n5594), .A(n4753), .ZN(n4754) );
  AOI21_X1 U5882 ( .B1(n5936), .B2(n6104), .A(n4754), .ZN(n4755) );
  OAI21_X1 U5883 ( .B1(n6100), .B2(n4756), .A(n4755), .ZN(U2982) );
  INV_X1 U5884 ( .A(DATAI_4_), .ZN(n6064) );
  INV_X1 U5885 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6026) );
  OAI222_X1 U5886 ( .A1(n4757), .A2(n5477), .B1(n5476), .B2(n6064), .C1(n5991), 
        .C2(n6026), .ZN(U2887) );
  NAND3_X1 U5887 ( .A1(n4729), .A2(n5793), .A3(n5061), .ZN(n4766) );
  OR2_X1 U5888 ( .A1(n4766), .A2(n6432), .ZN(n4758) );
  NAND2_X1 U5889 ( .A1(n4758), .A2(n6380), .ZN(n4762) );
  NOR2_X1 U5890 ( .A1(n4645), .A2(n4759), .ZN(n6275) );
  OR2_X1 U5891 ( .A1(n4647), .A2(n4520), .ZN(n6309) );
  NAND3_X1 U5892 ( .A1(n6509), .A2(n6306), .A3(n6504), .ZN(n4798) );
  NOR2_X1 U5893 ( .A1(n6378), .A2(n4798), .ZN(n6165) );
  AOI21_X1 U5894 ( .B1(n6275), .B2(n6338), .A(n6165), .ZN(n4760) );
  OAI22_X1 U5895 ( .A1(n4762), .A2(n4760), .B1(n4798), .B2(n4802), .ZN(n6167)
         );
  INV_X1 U5896 ( .A(n6167), .ZN(n4770) );
  INV_X1 U5897 ( .A(n4760), .ZN(n4761) );
  NOR2_X1 U5898 ( .A1(n4762), .A2(n4761), .ZN(n4765) );
  INV_X1 U5899 ( .A(n4798), .ZN(n4763) );
  OAI21_X1 U5900 ( .B1(n6380), .B2(n4763), .A(n6240), .ZN(n4764) );
  AOI22_X1 U5901 ( .A1(n6379), .A2(n6164), .B1(n6430), .B2(n6165), .ZN(n4767)
         );
  OAI21_X1 U5902 ( .B1(n6392), .B2(n4898), .A(n4767), .ZN(n4768) );
  AOI21_X1 U5903 ( .B1(INSTQUEUE_REG_1__0__SCAN_IN), .B2(n6163), .A(n4768), 
        .ZN(n4769) );
  OAI21_X1 U5904 ( .B1(n4770), .B2(n6348), .A(n4769), .ZN(U3028) );
  NAND2_X1 U5905 ( .A1(n4777), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4772) );
  NAND2_X1 U5906 ( .A1(n6380), .A2(n4772), .ZN(n4775) );
  NAND2_X1 U5907 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6206), .ZN(n6429) );
  NOR2_X1 U5908 ( .A1(n6378), .A2(n6429), .ZN(n4794) );
  AOI21_X1 U5909 ( .B1(n6339), .B2(n6437), .A(n4794), .ZN(n4776) );
  INV_X1 U5910 ( .A(n4776), .ZN(n4774) );
  INV_X1 U5911 ( .A(n6240), .ZN(n6384) );
  AOI21_X1 U5912 ( .B1(n6435), .B2(n6429), .A(n6384), .ZN(n4773) );
  OAI22_X1 U5913 ( .A1(n4776), .A2(n4775), .B1(n4802), .B2(n6429), .ZN(n4792)
         );
  AOI22_X1 U5914 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4793), .B1(n6477), 
        .B2(n4792), .ZN(n4779) );
  AOI22_X1 U5915 ( .A1(n6476), .A2(n4794), .B1(n6413), .B2(n6486), .ZN(n4778)
         );
  OAI211_X1 U5916 ( .C1(n6416), .C2(n4879), .A(n4779), .B(n4778), .ZN(U3130)
         );
  AOI22_X1 U5917 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4793), .B1(n6471), 
        .B2(n4792), .ZN(n4781) );
  AOI22_X1 U5918 ( .A1(n6470), .A2(n4794), .B1(n6409), .B2(n6486), .ZN(n4780)
         );
  OAI211_X1 U5919 ( .C1(n6412), .C2(n4879), .A(n4781), .B(n4780), .ZN(U3129)
         );
  AOI22_X1 U5920 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4793), .B1(n6465), 
        .B2(n4792), .ZN(n4783) );
  AOI22_X1 U5921 ( .A1(n6464), .A2(n4794), .B1(n6405), .B2(n6486), .ZN(n4782)
         );
  OAI211_X1 U5922 ( .C1(n6408), .C2(n4879), .A(n4783), .B(n4782), .ZN(U3128)
         );
  AOI22_X1 U5923 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4793), .B1(n6459), 
        .B2(n4792), .ZN(n4785) );
  AOI22_X1 U5924 ( .A1(n6458), .A2(n4794), .B1(n6401), .B2(n6486), .ZN(n4784)
         );
  OAI211_X1 U5925 ( .C1(n6404), .C2(n4879), .A(n4785), .B(n4784), .ZN(U3127)
         );
  AOI22_X1 U5926 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4793), .B1(n6431), 
        .B2(n4792), .ZN(n4787) );
  AOI22_X1 U5927 ( .A1(n6430), .A2(n4794), .B1(n6379), .B2(n6486), .ZN(n4786)
         );
  OAI211_X1 U5928 ( .C1(n4879), .C2(n6392), .A(n4787), .B(n4786), .ZN(U3124)
         );
  AOI22_X1 U5929 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4793), .B1(n6447), 
        .B2(n4792), .ZN(n4789) );
  AOI22_X1 U5930 ( .A1(n6446), .A2(n4794), .B1(n6393), .B2(n6486), .ZN(n4788)
         );
  OAI211_X1 U5931 ( .C1(n6396), .C2(n4879), .A(n4789), .B(n4788), .ZN(U3125)
         );
  AOI22_X1 U5932 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4793), .B1(n6485), 
        .B2(n4792), .ZN(n4791) );
  AOI22_X1 U5933 ( .A1(n6483), .A2(n4794), .B1(n6419), .B2(n6486), .ZN(n4790)
         );
  OAI211_X1 U5934 ( .C1(n6424), .C2(n4879), .A(n4791), .B(n4790), .ZN(U3131)
         );
  AOI22_X1 U5935 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4793), .B1(n6453), 
        .B2(n4792), .ZN(n4796) );
  AOI22_X1 U5936 ( .A1(n6452), .A2(n4794), .B1(n6352), .B2(n6486), .ZN(n4795)
         );
  OAI211_X1 U5937 ( .C1(n5076), .C2(n4879), .A(n4796), .B(n4795), .ZN(U3126)
         );
  NAND3_X1 U5938 ( .A1(n4918), .A2(n6380), .A3(n4834), .ZN(n4797) );
  AOI22_X1 U5939 ( .A1(n4797), .A2(n6208), .B1(n5950), .B2(n6338), .ZN(n4801)
         );
  NOR2_X1 U5940 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4798), .ZN(n4832)
         );
  INV_X1 U5941 ( .A(n4973), .ZN(n6426) );
  INV_X1 U5942 ( .A(n6304), .ZN(n4799) );
  OR2_X1 U5943 ( .A1(n6305), .A2(n4799), .ZN(n6205) );
  AOI21_X1 U5944 ( .B1(n6205), .B2(STATE2_REG_2__SCAN_IN), .A(n6312), .ZN(
        n6210) );
  OAI211_X1 U5945 ( .C1(n3238), .C2(n4832), .A(n6426), .B(n6210), .ZN(n4800)
         );
  INV_X1 U5946 ( .A(n6308), .ZN(n6313) );
  NOR2_X1 U5947 ( .A1(n4803), .A2(n4802), .ZN(n5066) );
  INV_X1 U5948 ( .A(n5066), .ZN(n6439) );
  OAI22_X1 U5949 ( .A1(n6313), .A2(n6309), .B1(n6439), .B2(n6205), .ZN(n4836)
         );
  AOI22_X1 U5950 ( .A1(n6442), .A2(n6164), .B1(n6430), .B2(n4832), .ZN(n4804)
         );
  OAI21_X1 U5951 ( .B1(n6445), .B2(n4834), .A(n4804), .ZN(n4805) );
  AOI21_X1 U5952 ( .B1(n6431), .B2(n4836), .A(n4805), .ZN(n4806) );
  OAI21_X1 U5953 ( .B1(n4839), .B2(n4807), .A(n4806), .ZN(U3020) );
  INV_X1 U5954 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4811) );
  INV_X1 U5955 ( .A(n6405), .ZN(n6469) );
  AOI22_X1 U5956 ( .A1(n6464), .A2(n4832), .B1(n6164), .B2(n6466), .ZN(n4808)
         );
  OAI21_X1 U5957 ( .B1(n6469), .B2(n4834), .A(n4808), .ZN(n4809) );
  AOI21_X1 U5958 ( .B1(n6465), .B2(n4836), .A(n4809), .ZN(n4810) );
  OAI21_X1 U5959 ( .B1(n4839), .B2(n4811), .A(n4810), .ZN(U3024) );
  INV_X1 U5960 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4815) );
  INV_X1 U5961 ( .A(n6419), .ZN(n6492) );
  AOI22_X1 U5962 ( .A1(n6483), .A2(n4832), .B1(n6164), .B2(n6487), .ZN(n4812)
         );
  OAI21_X1 U5963 ( .B1(n6492), .B2(n4834), .A(n4812), .ZN(n4813) );
  AOI21_X1 U5964 ( .B1(n6485), .B2(n4836), .A(n4813), .ZN(n4814) );
  OAI21_X1 U5965 ( .B1(n4839), .B2(n4815), .A(n4814), .ZN(U3027) );
  INV_X1 U5966 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4819) );
  INV_X1 U5967 ( .A(n6393), .ZN(n6451) );
  AOI22_X1 U5968 ( .A1(n6446), .A2(n4832), .B1(n6164), .B2(n6448), .ZN(n4816)
         );
  OAI21_X1 U5969 ( .B1(n6451), .B2(n4834), .A(n4816), .ZN(n4817) );
  AOI21_X1 U5970 ( .B1(n6447), .B2(n4836), .A(n4817), .ZN(n4818) );
  OAI21_X1 U5971 ( .B1(n4839), .B2(n4819), .A(n4818), .ZN(U3021) );
  INV_X1 U5972 ( .A(n6409), .ZN(n6475) );
  AOI22_X1 U5973 ( .A1(n6470), .A2(n4832), .B1(n6164), .B2(n6472), .ZN(n4820)
         );
  OAI21_X1 U5974 ( .B1(n6475), .B2(n4834), .A(n4820), .ZN(n4821) );
  AOI21_X1 U5975 ( .B1(n6471), .B2(n4836), .A(n4821), .ZN(n4822) );
  OAI21_X1 U5976 ( .B1(n4839), .B2(n4823), .A(n4822), .ZN(U3025) );
  AOI22_X1 U5977 ( .A1(n6452), .A2(n4832), .B1(n6164), .B2(n6454), .ZN(n4824)
         );
  OAI21_X1 U5978 ( .B1(n6457), .B2(n4834), .A(n4824), .ZN(n4825) );
  AOI21_X1 U5979 ( .B1(n6453), .B2(n4836), .A(n4825), .ZN(n4826) );
  OAI21_X1 U5980 ( .B1(n4839), .B2(n4827), .A(n4826), .ZN(U3022) );
  INV_X1 U5981 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4831) );
  AOI22_X1 U5982 ( .A1(n6476), .A2(n4832), .B1(n6164), .B2(n6478), .ZN(n4828)
         );
  OAI21_X1 U5983 ( .B1(n6481), .B2(n4834), .A(n4828), .ZN(n4829) );
  AOI21_X1 U5984 ( .B1(n6477), .B2(n4836), .A(n4829), .ZN(n4830) );
  OAI21_X1 U5985 ( .B1(n4839), .B2(n4831), .A(n4830), .ZN(U3026) );
  INV_X1 U5986 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4838) );
  AOI22_X1 U5987 ( .A1(n6458), .A2(n4832), .B1(n6164), .B2(n6460), .ZN(n4833)
         );
  OAI21_X1 U5988 ( .B1(n6463), .B2(n4834), .A(n4833), .ZN(n4835) );
  AOI21_X1 U5989 ( .B1(n6459), .B2(n4836), .A(n4835), .ZN(n4837) );
  OAI21_X1 U5990 ( .B1(n4839), .B2(n4838), .A(n4837), .ZN(U3023) );
  OR2_X1 U5991 ( .A1(n4742), .A2(n4842), .ZN(n4843) );
  AND2_X1 U5992 ( .A1(n4841), .A2(n4843), .ZN(n6103) );
  INV_X1 U5993 ( .A(n6103), .ZN(n4845) );
  AOI22_X1 U5994 ( .A1(n5988), .A2(DATAI_6_), .B1(EAX_REG_6__SCAN_IN), .B2(
        n5473), .ZN(n4844) );
  OAI21_X1 U5995 ( .B1(n4845), .B2(n5477), .A(n4844), .ZN(U2885) );
  INV_X1 U5996 ( .A(n4846), .ZN(n5923) );
  INV_X1 U5997 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6574) );
  NOR2_X1 U5998 ( .A1(n6122), .A2(n6574), .ZN(n6137) );
  AOI21_X1 U5999 ( .B1(n6094), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n6137), 
        .ZN(n4847) );
  OAI21_X1 U6000 ( .B1(n5925), .B2(n5594), .A(n4847), .ZN(n4848) );
  AOI21_X1 U6001 ( .B1(n5923), .B2(n6104), .A(n4848), .ZN(n4849) );
  OAI21_X1 U6002 ( .B1(n6143), .B2(n6100), .A(n4849), .ZN(U2981) );
  NOR2_X1 U6003 ( .A1(n5950), .A2(n6435), .ZN(n6303) );
  INV_X1 U6004 ( .A(n6305), .ZN(n4938) );
  NOR2_X1 U6005 ( .A1(n4938), .A2(n6509), .ZN(n5065) );
  AOI22_X1 U6006 ( .A1(n6303), .A2(n6274), .B1(n4973), .B2(n5065), .ZN(n4885)
         );
  OR2_X1 U6007 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4850), .ZN(n4880)
         );
  OAI22_X1 U6008 ( .A1(n4947), .A2(n4880), .B1(n6445), .B2(n4879), .ZN(n4851)
         );
  AOI21_X1 U6009 ( .B1(n6442), .B2(n4882), .A(n4851), .ZN(n4859) );
  OAI21_X1 U6010 ( .B1(n6305), .B2(n4802), .A(n4852), .ZN(n4975) );
  NOR2_X1 U6011 ( .A1(n5066), .A2(n4975), .ZN(n4857) );
  AOI21_X1 U6012 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n4880), .A(n6509), .ZN(
        n4856) );
  INV_X1 U6013 ( .A(n4879), .ZN(n4853) );
  OAI21_X1 U6014 ( .B1(n4853), .B2(n4882), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4854) );
  NOR2_X1 U6015 ( .A1(n6274), .A2(n6435), .ZN(n4977) );
  NAND2_X1 U6016 ( .A1(n4854), .A2(n4977), .ZN(n4855) );
  NAND3_X1 U6017 ( .A1(n4857), .A2(n4856), .A3(n4855), .ZN(n4878) );
  NAND2_X1 U6018 ( .A1(n4878), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4858)
         );
  OAI211_X1 U6019 ( .C1(n4885), .C2(n6348), .A(n4859), .B(n4858), .ZN(U3132)
         );
  NAND2_X1 U6020 ( .A1(n4878), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4862)
         );
  OAI22_X1 U6021 ( .A1(n5094), .A2(n4880), .B1(n6463), .B2(n4879), .ZN(n4860)
         );
  AOI21_X1 U6022 ( .B1(n6460), .B2(n4882), .A(n4860), .ZN(n4861) );
  OAI211_X1 U6023 ( .C1(n4885), .C2(n6358), .A(n4862), .B(n4861), .ZN(U3135)
         );
  NAND2_X1 U6024 ( .A1(n4878), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4865)
         );
  OAI22_X1 U6025 ( .A1(n5079), .A2(n4880), .B1(n6451), .B2(n4879), .ZN(n4863)
         );
  AOI21_X1 U6026 ( .B1(n6448), .B2(n4882), .A(n4863), .ZN(n4864) );
  OAI211_X1 U6027 ( .C1(n4885), .C2(n6351), .A(n4865), .B(n4864), .ZN(U3133)
         );
  NAND2_X1 U6028 ( .A1(n4878), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4868)
         );
  OAI22_X1 U6029 ( .A1(n5089), .A2(n4880), .B1(n6475), .B2(n4879), .ZN(n4866)
         );
  AOI21_X1 U6030 ( .B1(n6472), .B2(n4882), .A(n4866), .ZN(n4867) );
  OAI211_X1 U6031 ( .C1(n4885), .C2(n6364), .A(n4868), .B(n4867), .ZN(U3137)
         );
  NAND2_X1 U6032 ( .A1(n4878), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4871)
         );
  OAI22_X1 U6033 ( .A1(n5105), .A2(n4880), .B1(n6469), .B2(n4879), .ZN(n4869)
         );
  AOI21_X1 U6034 ( .B1(n6466), .B2(n4882), .A(n4869), .ZN(n4870) );
  OAI211_X1 U6035 ( .C1(n4885), .C2(n6361), .A(n4871), .B(n4870), .ZN(U3136)
         );
  NAND2_X1 U6036 ( .A1(n4878), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4874)
         );
  OAI22_X1 U6037 ( .A1(n5084), .A2(n4880), .B1(n6492), .B2(n4879), .ZN(n4872)
         );
  AOI21_X1 U6038 ( .B1(n6487), .B2(n4882), .A(n4872), .ZN(n4873) );
  OAI211_X1 U6039 ( .C1(n4885), .C2(n6374), .A(n4874), .B(n4873), .ZN(U3139)
         );
  NAND2_X1 U6040 ( .A1(n4878), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4877)
         );
  OAI22_X1 U6041 ( .A1(n5068), .A2(n4880), .B1(n6457), .B2(n4879), .ZN(n4875)
         );
  AOI21_X1 U6042 ( .B1(n6454), .B2(n4882), .A(n4875), .ZN(n4876) );
  OAI211_X1 U6043 ( .C1(n4885), .C2(n6355), .A(n4877), .B(n4876), .ZN(U3134)
         );
  NAND2_X1 U6044 ( .A1(n4878), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4884)
         );
  OAI22_X1 U6045 ( .A1(n5099), .A2(n4880), .B1(n6481), .B2(n4879), .ZN(n4881)
         );
  AOI21_X1 U6046 ( .B1(n6478), .B2(n4882), .A(n4881), .ZN(n4883) );
  OAI211_X1 U6047 ( .C1(n4885), .C2(n6367), .A(n4884), .B(n4883), .ZN(U3138)
         );
  XNOR2_X1 U6048 ( .A(n4887), .B(n4886), .ZN(n6102) );
  NOR2_X1 U6049 ( .A1(n4744), .A2(n4889), .ZN(n4890) );
  AND2_X1 U6051 ( .A1(n5696), .A2(n4893), .ZN(n4891) );
  OR2_X1 U6052 ( .A1(n4892), .A2(n4891), .ZN(n6136) );
  INV_X1 U6053 ( .A(n6136), .ZN(n4894) );
  OAI33_X1 U6054 ( .A1(1'b0), .A2(n4894), .A3(n4169), .B1(
        INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n4929), .B3(n4893), .ZN(n4896) );
  INV_X1 U6055 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6576) );
  NOR2_X1 U6056 ( .A1(n6122), .A2(n6576), .ZN(n6109) );
  AOI211_X1 U6057 ( .C1(n3108), .C2(n6138), .A(n4896), .B(n6109), .ZN(n4897)
         );
  OAI21_X1 U6058 ( .B1(n6102), .B2(n6142), .A(n4897), .ZN(U3012) );
  INV_X1 U6059 ( .A(n6165), .ZN(n4915) );
  AOI22_X1 U6060 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n6163), .B1(n6459), 
        .B2(n6167), .ZN(n4899) );
  OAI21_X1 U6061 ( .B1(n5094), .B2(n4915), .A(n4899), .ZN(n4900) );
  AOI21_X1 U6062 ( .B1(n6460), .B2(n6166), .A(n4900), .ZN(n4901) );
  OAI21_X1 U6063 ( .B1(n6463), .B2(n4918), .A(n4901), .ZN(U3031) );
  AOI22_X1 U6064 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n6163), .B1(n6453), 
        .B2(n6167), .ZN(n4902) );
  OAI21_X1 U6065 ( .B1(n5068), .B2(n4915), .A(n4902), .ZN(n4903) );
  AOI21_X1 U6066 ( .B1(n6454), .B2(n6166), .A(n4903), .ZN(n4904) );
  OAI21_X1 U6067 ( .B1(n6457), .B2(n4918), .A(n4904), .ZN(U3030) );
  AOI22_X1 U6068 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n6163), .B1(n6471), 
        .B2(n6167), .ZN(n4905) );
  OAI21_X1 U6069 ( .B1(n5089), .B2(n4915), .A(n4905), .ZN(n4906) );
  AOI21_X1 U6070 ( .B1(n6472), .B2(n6166), .A(n4906), .ZN(n4907) );
  OAI21_X1 U6071 ( .B1(n6475), .B2(n4918), .A(n4907), .ZN(U3033) );
  AOI22_X1 U6072 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n6163), .B1(n6477), 
        .B2(n6167), .ZN(n4908) );
  OAI21_X1 U6073 ( .B1(n5099), .B2(n4915), .A(n4908), .ZN(n4909) );
  AOI21_X1 U6074 ( .B1(n6478), .B2(n6166), .A(n4909), .ZN(n4910) );
  OAI21_X1 U6075 ( .B1(n6481), .B2(n4918), .A(n4910), .ZN(U3034) );
  AOI22_X1 U6076 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n6163), .B1(n6485), 
        .B2(n6167), .ZN(n4911) );
  OAI21_X1 U6077 ( .B1(n5084), .B2(n4915), .A(n4911), .ZN(n4912) );
  AOI21_X1 U6078 ( .B1(n6487), .B2(n6166), .A(n4912), .ZN(n4913) );
  OAI21_X1 U6079 ( .B1(n6492), .B2(n4918), .A(n4913), .ZN(U3035) );
  AOI22_X1 U6080 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n6163), .B1(n6447), 
        .B2(n6167), .ZN(n4914) );
  OAI21_X1 U6081 ( .B1(n5079), .B2(n4915), .A(n4914), .ZN(n4916) );
  AOI21_X1 U6082 ( .B1(n6448), .B2(n6166), .A(n4916), .ZN(n4917) );
  OAI21_X1 U6083 ( .B1(n6451), .B2(n4918), .A(n4917), .ZN(U3029) );
  NOR2_X1 U6084 ( .A1(n4841), .A2(n4919), .ZN(n5046) );
  AOI21_X1 U6085 ( .B1(n4919), .B2(n4841), .A(n5046), .ZN(n5004) );
  INV_X1 U6086 ( .A(n5438), .ZN(n5980) );
  OR2_X1 U6087 ( .A1(n4888), .A2(n4921), .ZN(n4922) );
  NAND2_X1 U6088 ( .A1(n4920), .A2(n4922), .ZN(n5897) );
  OAI22_X1 U6089 ( .A1(n5897), .A2(n5433), .B1(n4923), .B2(n5987), .ZN(n4924)
         );
  AOI21_X1 U6090 ( .B1(n5004), .B2(n5980), .A(n4924), .ZN(n4925) );
  INV_X1 U6091 ( .A(n4925), .ZN(U2852) );
  XNOR2_X1 U6092 ( .A(n4926), .B(n4927), .ZN(n5006) );
  NOR2_X1 U6093 ( .A1(n4929), .A2(n4928), .ZN(n6120) );
  INV_X1 U6094 ( .A(n5735), .ZN(n4930) );
  NAND2_X1 U6095 ( .A1(n4931), .A2(n4930), .ZN(n4934) );
  NAND2_X1 U6096 ( .A1(n5737), .A2(n4932), .ZN(n4933) );
  NOR2_X1 U6097 ( .A1(n6121), .A2(n4178), .ZN(n4936) );
  NAND2_X1 U6098 ( .A1(n6095), .A2(REIP_REG_7__SCAN_IN), .ZN(n5001) );
  OAI21_X1 U6099 ( .B1(n5897), .B2(n6149), .A(n5001), .ZN(n4935) );
  AOI211_X1 U6100 ( .C1(n6120), .C2(n4178), .A(n4936), .B(n4935), .ZN(n4937)
         );
  OAI21_X1 U6101 ( .B1(n5006), .B2(n6142), .A(n4937), .ZN(U3011) );
  OR2_X1 U6102 ( .A1(n5963), .A2(n4647), .ZN(n4940) );
  NOR2_X1 U6103 ( .A1(n4938), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4974)
         );
  AOI22_X1 U6104 ( .A1(n6308), .A2(n6175), .B1(n4974), .B2(n5066), .ZN(n4972)
         );
  OAI21_X1 U6105 ( .B1(n6166), .B2(n6199), .A(n6208), .ZN(n4939) );
  OAI21_X1 U6106 ( .B1(n4940), .B2(n4645), .A(n4939), .ZN(n4941) );
  AND2_X1 U6107 ( .A1(n4941), .A2(n3238), .ZN(n4942) );
  OR2_X1 U6108 ( .A1(n5067), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6180)
         );
  NOR2_X1 U6109 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6180), .ZN(n4943)
         );
  NOR2_X1 U6110 ( .A1(n4973), .A2(n4975), .ZN(n5073) );
  NAND2_X1 U6111 ( .A1(n4966), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4946) );
  INV_X1 U6112 ( .A(n4943), .ZN(n4967) );
  OAI22_X1 U6113 ( .A1(n4968), .A2(n6396), .B1(n5079), .B2(n4967), .ZN(n4944)
         );
  AOI21_X1 U6114 ( .B1(n6393), .B2(n6166), .A(n4944), .ZN(n4945) );
  OAI211_X1 U6115 ( .C1(n4972), .C2(n6351), .A(n4946), .B(n4945), .ZN(U3037)
         );
  NAND2_X1 U6116 ( .A1(n4966), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4950) );
  OAI22_X1 U6117 ( .A1(n4947), .A2(n4967), .B1(n6392), .B2(n4968), .ZN(n4948)
         );
  AOI21_X1 U6118 ( .B1(n6379), .B2(n6166), .A(n4948), .ZN(n4949) );
  OAI211_X1 U6119 ( .C1(n4972), .C2(n6348), .A(n4950), .B(n4949), .ZN(U3036)
         );
  NAND2_X1 U6120 ( .A1(n4966), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4953) );
  OAI22_X1 U6121 ( .A1(n4968), .A2(n6404), .B1(n5094), .B2(n4967), .ZN(n4951)
         );
  AOI21_X1 U6122 ( .B1(n6401), .B2(n6166), .A(n4951), .ZN(n4952) );
  OAI211_X1 U6123 ( .C1(n4972), .C2(n6358), .A(n4953), .B(n4952), .ZN(U3039)
         );
  NAND2_X1 U6124 ( .A1(n4966), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4956) );
  OAI22_X1 U6125 ( .A1(n4968), .A2(n6408), .B1(n5105), .B2(n4967), .ZN(n4954)
         );
  AOI21_X1 U6126 ( .B1(n6405), .B2(n6166), .A(n4954), .ZN(n4955) );
  OAI211_X1 U6127 ( .C1(n4972), .C2(n6361), .A(n4956), .B(n4955), .ZN(U3040)
         );
  NAND2_X1 U6128 ( .A1(n4966), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4959) );
  OAI22_X1 U6129 ( .A1(n4968), .A2(n6424), .B1(n5084), .B2(n4967), .ZN(n4957)
         );
  AOI21_X1 U6130 ( .B1(n6419), .B2(n6166), .A(n4957), .ZN(n4958) );
  OAI211_X1 U6131 ( .C1(n4972), .C2(n6374), .A(n4959), .B(n4958), .ZN(U3043)
         );
  NAND2_X1 U6132 ( .A1(n4966), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4962) );
  OAI22_X1 U6133 ( .A1(n4968), .A2(n5076), .B1(n5068), .B2(n4967), .ZN(n4960)
         );
  AOI21_X1 U6134 ( .B1(n6352), .B2(n6166), .A(n4960), .ZN(n4961) );
  OAI211_X1 U6135 ( .C1(n4972), .C2(n6355), .A(n4962), .B(n4961), .ZN(U3038)
         );
  NAND2_X1 U6136 ( .A1(n4966), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4965) );
  OAI22_X1 U6137 ( .A1(n4968), .A2(n6412), .B1(n5089), .B2(n4967), .ZN(n4963)
         );
  AOI21_X1 U6138 ( .B1(n6409), .B2(n6166), .A(n4963), .ZN(n4964) );
  OAI211_X1 U6139 ( .C1(n4972), .C2(n6364), .A(n4965), .B(n4964), .ZN(U3041)
         );
  NAND2_X1 U6140 ( .A1(n4966), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4971) );
  OAI22_X1 U6141 ( .A1(n4968), .A2(n6416), .B1(n5099), .B2(n4967), .ZN(n4969)
         );
  AOI21_X1 U6142 ( .B1(n6413), .B2(n6166), .A(n4969), .ZN(n4970) );
  OAI211_X1 U6143 ( .C1(n4972), .C2(n6367), .A(n4971), .B(n4970), .ZN(U3042)
         );
  INV_X1 U6144 ( .A(n5004), .ZN(n5900) );
  OAI222_X1 U6145 ( .A1(n5900), .A2(n5477), .B1(n5476), .B2(n6070), .C1(n5991), 
        .C2(n3485), .ZN(U2884) );
  AOI22_X1 U6146 ( .A1(n6308), .A2(n6274), .B1(n4974), .B2(n4973), .ZN(n6263)
         );
  NOR2_X1 U6147 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6279), .ZN(n6264)
         );
  NAND3_X1 U6148 ( .A1(n5061), .A2(n6172), .A3(n2989), .ZN(n6213) );
  OAI21_X1 U6149 ( .B1(n6266), .B2(n6298), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4976) );
  AOI211_X1 U6150 ( .C1(n4977), .C2(n4976), .A(n5066), .B(n4975), .ZN(n4978)
         );
  NAND2_X1 U6151 ( .A1(n6267), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4981) );
  INV_X1 U6152 ( .A(n6264), .ZN(n4997) );
  OAI22_X1 U6153 ( .A1(n5099), .A2(n4997), .B1(n6270), .B2(n6416), .ZN(n4979)
         );
  AOI21_X1 U6154 ( .B1(n6266), .B2(n6413), .A(n4979), .ZN(n4980) );
  OAI211_X1 U6155 ( .C1(n6263), .C2(n6367), .A(n4981), .B(n4980), .ZN(U3074)
         );
  NAND2_X1 U6156 ( .A1(n6267), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4984) );
  OAI22_X1 U6157 ( .A1(n5105), .A2(n4997), .B1(n6270), .B2(n6408), .ZN(n4982)
         );
  AOI21_X1 U6158 ( .B1(n6266), .B2(n6405), .A(n4982), .ZN(n4983) );
  OAI211_X1 U6159 ( .C1(n6263), .C2(n6361), .A(n4984), .B(n4983), .ZN(U3072)
         );
  NAND2_X1 U6160 ( .A1(n6267), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4987) );
  OAI22_X1 U6161 ( .A1(n5084), .A2(n4997), .B1(n6270), .B2(n6424), .ZN(n4985)
         );
  AOI21_X1 U6162 ( .B1(n6266), .B2(n6419), .A(n4985), .ZN(n4986) );
  OAI211_X1 U6163 ( .C1(n6263), .C2(n6374), .A(n4987), .B(n4986), .ZN(U3075)
         );
  NAND2_X1 U6164 ( .A1(n6267), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4990) );
  OAI22_X1 U6165 ( .A1(n5068), .A2(n4997), .B1(n6270), .B2(n5076), .ZN(n4988)
         );
  AOI21_X1 U6166 ( .B1(n6266), .B2(n6352), .A(n4988), .ZN(n4989) );
  OAI211_X1 U6167 ( .C1(n6263), .C2(n6355), .A(n4990), .B(n4989), .ZN(U3070)
         );
  NAND2_X1 U6168 ( .A1(n6267), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4993) );
  OAI22_X1 U6169 ( .A1(n5079), .A2(n4997), .B1(n6270), .B2(n6396), .ZN(n4991)
         );
  AOI21_X1 U6170 ( .B1(n6266), .B2(n6393), .A(n4991), .ZN(n4992) );
  OAI211_X1 U6171 ( .C1(n6263), .C2(n6351), .A(n4993), .B(n4992), .ZN(U3069)
         );
  NAND2_X1 U6172 ( .A1(n6267), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4996) );
  OAI22_X1 U6173 ( .A1(n5094), .A2(n4997), .B1(n6270), .B2(n6404), .ZN(n4994)
         );
  AOI21_X1 U6174 ( .B1(n6266), .B2(n6401), .A(n4994), .ZN(n4995) );
  OAI211_X1 U6175 ( .C1(n6263), .C2(n6358), .A(n4996), .B(n4995), .ZN(U3071)
         );
  NAND2_X1 U6176 ( .A1(n6267), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n5000) );
  OAI22_X1 U6177 ( .A1(n5089), .A2(n4997), .B1(n6270), .B2(n6412), .ZN(n4998)
         );
  AOI21_X1 U6178 ( .B1(n6266), .B2(n6409), .A(n4998), .ZN(n4999) );
  OAI211_X1 U6179 ( .C1(n6263), .C2(n6364), .A(n5000), .B(n4999), .ZN(U3073)
         );
  NAND2_X1 U6180 ( .A1(n6094), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5002)
         );
  OAI211_X1 U6181 ( .C1(n5594), .C2(n5898), .A(n5002), .B(n5001), .ZN(n5003)
         );
  AOI21_X1 U6182 ( .B1(n5004), .B2(n6104), .A(n5003), .ZN(n5005) );
  OAI21_X1 U6183 ( .B1(n5006), .B2(n6100), .A(n5005), .ZN(U2979) );
  NOR2_X1 U6184 ( .A1(n5007), .A2(n5008), .ZN(n5009) );
  OR2_X1 U6185 ( .A1(n3000), .A2(n5009), .ZN(n5386) );
  AOI22_X1 U6186 ( .A1(n5988), .A2(DATAI_9_), .B1(EAX_REG_9__SCAN_IN), .B2(
        n5473), .ZN(n5010) );
  OAI21_X1 U6187 ( .B1(n5386), .B2(n5477), .A(n5010), .ZN(U2882) );
  INV_X1 U6188 ( .A(n5386), .ZN(n5035) );
  NAND2_X1 U6189 ( .A1(n5012), .A2(n5013), .ZN(n5014) );
  NAND2_X1 U6190 ( .A1(n5011), .A2(n5014), .ZN(n5384) );
  OAI22_X1 U6191 ( .A1(n5384), .A2(n5433), .B1(n5015), .B2(n5987), .ZN(n5016)
         );
  AOI21_X1 U6192 ( .B1(n5035), .B2(n5980), .A(n5016), .ZN(n5017) );
  INV_X1 U6193 ( .A(n5017), .ZN(U2850) );
  INV_X1 U6194 ( .A(n5018), .ZN(n5020) );
  INV_X1 U6195 ( .A(n3000), .ZN(n5019) );
  AOI21_X1 U6196 ( .B1(n5020), .B2(n5019), .A(n3012), .ZN(n5881) );
  INV_X1 U6197 ( .A(n5881), .ZN(n5031) );
  AOI22_X1 U6198 ( .A1(n5988), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n5473), .ZN(n5021) );
  OAI21_X1 U6199 ( .B1(n5031), .B2(n5477), .A(n5021), .ZN(U2881) );
  XNOR2_X1 U6200 ( .A(n5023), .B(n5022), .ZN(n5037) );
  OAI21_X1 U6201 ( .B1(n6130), .B2(n6153), .A(n6121), .ZN(n5775) );
  NAND2_X1 U6202 ( .A1(n6095), .A2(REIP_REG_9__SCAN_IN), .ZN(n5032) );
  OAI21_X1 U6203 ( .B1(n5384), .B2(n6149), .A(n5032), .ZN(n5025) );
  NAND2_X1 U6204 ( .A1(n6130), .A2(n6120), .ZN(n5772) );
  NOR2_X1 U6205 ( .A1(n5772), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5024)
         );
  AOI211_X1 U6206 ( .C1(n5775), .C2(INSTADDRPOINTER_REG_9__SCAN_IN), .A(n5025), 
        .B(n5024), .ZN(n5026) );
  OAI21_X1 U6207 ( .B1(n5037), .B2(n6142), .A(n5026), .ZN(U3009) );
  AOI21_X1 U6208 ( .B1(n5028), .B2(n5011), .A(n5027), .ZN(n5877) );
  INV_X1 U6209 ( .A(n5877), .ZN(n5029) );
  OAI222_X1 U6210 ( .A1(n5031), .A2(n5438), .B1(n5030), .B2(n5987), .C1(n5433), 
        .C2(n5029), .ZN(U2849) );
  NAND2_X1 U6211 ( .A1(n6094), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5033)
         );
  OAI211_X1 U6212 ( .C1(n5594), .C2(n5385), .A(n5033), .B(n5032), .ZN(n5034)
         );
  AOI21_X1 U6213 ( .B1(n5035), .B2(n6104), .A(n5034), .ZN(n5036) );
  OAI21_X1 U6214 ( .B1(n5037), .B2(n6100), .A(n5036), .ZN(U2977) );
  OAI21_X1 U6215 ( .B1(n3012), .B2(n3549), .A(n5040), .ZN(n5598) );
  OAI21_X1 U6216 ( .B1(n5027), .B2(n5042), .A(n5041), .ZN(n5043) );
  INV_X1 U6217 ( .A(n5043), .ZN(n6114) );
  AOI22_X1 U6218 ( .A1(n6114), .A2(n5979), .B1(EBX_REG_11__SCAN_IN), .B2(n5436), .ZN(n5044) );
  OAI21_X1 U6219 ( .B1(n5598), .B2(n5438), .A(n5044), .ZN(U2848) );
  AOI22_X1 U6220 ( .A1(n5988), .A2(DATAI_11_), .B1(EAX_REG_11__SCAN_IN), .B2(
        n5473), .ZN(n5045) );
  OAI21_X1 U6221 ( .B1(n5598), .B2(n5477), .A(n5045), .ZN(U2880) );
  INV_X1 U6222 ( .A(n5046), .ZN(n5048) );
  AND2_X1 U6223 ( .A1(n5048), .A2(n5047), .ZN(n5049) );
  NOR2_X1 U6224 ( .A1(n5007), .A2(n5049), .ZN(n5889) );
  INV_X1 U6225 ( .A(n5889), .ZN(n5060) );
  AOI22_X1 U6226 ( .A1(n5988), .A2(DATAI_8_), .B1(EAX_REG_8__SCAN_IN), .B2(
        n5473), .ZN(n5050) );
  OAI21_X1 U6227 ( .B1(n5060), .B2(n5477), .A(n5050), .ZN(U2883) );
  XNOR2_X1 U6228 ( .A(n5051), .B(n5052), .ZN(n6124) );
  AOI22_X1 U6229 ( .A1(n6094), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n6095), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n5053) );
  OAI21_X1 U6230 ( .B1(n5594), .B2(n5054), .A(n5053), .ZN(n5055) );
  AOI21_X1 U6231 ( .B1(n5889), .B2(n6104), .A(n5055), .ZN(n5056) );
  OAI21_X1 U6232 ( .B1(n6124), .B2(n6100), .A(n5056), .ZN(U2978) );
  INV_X1 U6233 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5059) );
  INV_X1 U6234 ( .A(n5012), .ZN(n5057) );
  AOI21_X1 U6235 ( .B1(n5058), .B2(n4920), .A(n5057), .ZN(n5887) );
  INV_X1 U6236 ( .A(n5887), .ZN(n6123) );
  OAI222_X1 U6237 ( .A1(n5060), .A2(n5438), .B1(n5059), .B2(n5987), .C1(n5433), 
        .C2(n6123), .ZN(U2851) );
  NAND2_X1 U6238 ( .A1(n5114), .A2(n6400), .ZN(n5064) );
  AOI21_X1 U6239 ( .B1(n5064), .B2(STATEBS16_REG_SCAN_IN), .A(n6435), .ZN(
        n5071) );
  AND2_X1 U6240 ( .A1(n6175), .A2(n4645), .ZN(n6383) );
  OR2_X1 U6241 ( .A1(n5067), .A2(n6509), .ZN(n6387) );
  NOR2_X1 U6242 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6387), .ZN(n5111)
         );
  INV_X1 U6243 ( .A(n5111), .ZN(n5104) );
  OR2_X1 U6244 ( .A1(n5068), .A2(n5104), .ZN(n5075) );
  INV_X1 U6245 ( .A(n6383), .ZN(n5070) );
  NOR2_X1 U6246 ( .A1(n5111), .A2(n3238), .ZN(n5069) );
  AOI21_X1 U6247 ( .B1(n5071), .B2(n5070), .A(n5069), .ZN(n5072) );
  OAI211_X1 U6248 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n4802), .A(n5073), .B(n5072), .ZN(n5110) );
  NAND2_X1 U6249 ( .A1(INSTQUEUE_REG_10__2__SCAN_IN), .A2(n5110), .ZN(n5074)
         );
  OAI211_X1 U6250 ( .C1(n6400), .C2(n5076), .A(n5075), .B(n5074), .ZN(n5077)
         );
  AOI21_X1 U6251 ( .B1(n6352), .B2(n6370), .A(n5077), .ZN(n5078) );
  OAI21_X1 U6252 ( .B1(n5117), .B2(n6355), .A(n5078), .ZN(U3102) );
  OR2_X1 U6253 ( .A1(n5079), .A2(n5104), .ZN(n5081) );
  NAND2_X1 U6254 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(n5110), .ZN(n5080)
         );
  OAI211_X1 U6255 ( .C1(n6400), .C2(n6396), .A(n5081), .B(n5080), .ZN(n5082)
         );
  AOI21_X1 U6256 ( .B1(n6393), .B2(n6370), .A(n5082), .ZN(n5083) );
  OAI21_X1 U6257 ( .B1(n5117), .B2(n6351), .A(n5083), .ZN(U3101) );
  OR2_X1 U6258 ( .A1(n5084), .A2(n5104), .ZN(n5086) );
  NAND2_X1 U6259 ( .A1(INSTQUEUE_REG_10__7__SCAN_IN), .A2(n5110), .ZN(n5085)
         );
  OAI211_X1 U6260 ( .C1(n6400), .C2(n6424), .A(n5086), .B(n5085), .ZN(n5087)
         );
  AOI21_X1 U6261 ( .B1(n6419), .B2(n6370), .A(n5087), .ZN(n5088) );
  OAI21_X1 U6262 ( .B1(n5117), .B2(n6374), .A(n5088), .ZN(U3107) );
  OR2_X1 U6263 ( .A1(n5089), .A2(n5104), .ZN(n5091) );
  NAND2_X1 U6264 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(n5110), .ZN(n5090)
         );
  OAI211_X1 U6265 ( .C1(n6400), .C2(n6412), .A(n5091), .B(n5090), .ZN(n5092)
         );
  AOI21_X1 U6266 ( .B1(n6409), .B2(n6370), .A(n5092), .ZN(n5093) );
  OAI21_X1 U6267 ( .B1(n5117), .B2(n6364), .A(n5093), .ZN(U3105) );
  OR2_X1 U6268 ( .A1(n5094), .A2(n5104), .ZN(n5096) );
  NAND2_X1 U6269 ( .A1(INSTQUEUE_REG_10__3__SCAN_IN), .A2(n5110), .ZN(n5095)
         );
  OAI211_X1 U6270 ( .C1(n6400), .C2(n6404), .A(n5096), .B(n5095), .ZN(n5097)
         );
  AOI21_X1 U6271 ( .B1(n6401), .B2(n6370), .A(n5097), .ZN(n5098) );
  OAI21_X1 U6272 ( .B1(n5117), .B2(n6358), .A(n5098), .ZN(U3103) );
  OR2_X1 U6273 ( .A1(n5099), .A2(n5104), .ZN(n5101) );
  NAND2_X1 U6274 ( .A1(INSTQUEUE_REG_10__6__SCAN_IN), .A2(n5110), .ZN(n5100)
         );
  OAI211_X1 U6275 ( .C1(n6400), .C2(n6416), .A(n5101), .B(n5100), .ZN(n5102)
         );
  AOI21_X1 U6276 ( .B1(n6413), .B2(n6370), .A(n5102), .ZN(n5103) );
  OAI21_X1 U6277 ( .B1(n5117), .B2(n6367), .A(n5103), .ZN(U3106) );
  OR2_X1 U6278 ( .A1(n5105), .A2(n5104), .ZN(n5107) );
  NAND2_X1 U6279 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n5110), .ZN(n5106)
         );
  OAI211_X1 U6280 ( .C1(n6400), .C2(n6408), .A(n5107), .B(n5106), .ZN(n5108)
         );
  AOI21_X1 U6281 ( .B1(n6405), .B2(n6370), .A(n5108), .ZN(n5109) );
  OAI21_X1 U6282 ( .B1(n5117), .B2(n6361), .A(n5109), .ZN(U3104) );
  AOI22_X1 U6283 ( .A1(n6430), .A2(n5111), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5110), .ZN(n5113) );
  OR2_X1 U6284 ( .A1(n6400), .A2(n6392), .ZN(n5112) );
  OAI211_X1 U6285 ( .C1(n5114), .C2(n6445), .A(n5113), .B(n5112), .ZN(n5115)
         );
  INV_X1 U6286 ( .A(n5115), .ZN(n5116) );
  OAI21_X1 U6287 ( .B1(n5117), .B2(n6348), .A(n5116), .ZN(U3100) );
  INV_X1 U6288 ( .A(n5118), .ZN(n5230) );
  AOI21_X1 U6289 ( .B1(n5119), .B2(n5230), .A(n4489), .ZN(n5667) );
  AOI22_X1 U6290 ( .A1(n5667), .A2(n5979), .B1(EBX_REG_24__SCAN_IN), .B2(n5436), .ZN(n5120) );
  OAI21_X1 U6291 ( .B1(n4437), .B2(n5438), .A(n5120), .ZN(U2835) );
  INV_X1 U6292 ( .A(n5121), .ZN(n5236) );
  INV_X1 U6293 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6607) );
  NAND2_X1 U6294 ( .A1(n5122), .A2(n6607), .ZN(n5142) );
  NAND2_X1 U6295 ( .A1(n5960), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5123)
         );
  OAI211_X1 U6296 ( .C1(n5965), .C2(n5124), .A(n5142), .B(n5123), .ZN(n5125)
         );
  AOI21_X1 U6297 ( .B1(n5961), .B2(EBX_REG_24__SCAN_IN), .A(n5125), .ZN(n5126)
         );
  OAI21_X1 U6298 ( .B1(n5236), .B2(n6607), .A(n5126), .ZN(n5127) );
  AOI21_X1 U6299 ( .B1(n5667), .B2(n5927), .A(n5127), .ZN(n5128) );
  OAI21_X1 U6300 ( .B1(n4437), .B2(n5899), .A(n5128), .ZN(U2803) );
  NOR2_X1 U6301 ( .A1(n5630), .A2(n5129), .ZN(n5131) );
  MUX2_X1 U6302 ( .A(n5131), .B(n5130), .S(INSTADDRPOINTER_REG_30__SCAN_IN), 
        .Z(n5132) );
  INV_X1 U6303 ( .A(n5132), .ZN(n5133) );
  INV_X1 U6304 ( .A(n5135), .ZN(n5136) );
  OAI21_X1 U6305 ( .B1(n5137), .B2(n6142), .A(n5136), .ZN(U2988) );
  NAND2_X1 U6306 ( .A1(n5138), .A2(n4228), .ZN(n5146) );
  INV_X1 U6307 ( .A(n5220), .ZN(n5139) );
  INV_X1 U6308 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6609) );
  AOI22_X1 U6309 ( .A1(n5960), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .B1(n5139), 
        .B2(n6609), .ZN(n5140) );
  OAI21_X1 U6310 ( .B1(n5965), .B2(n5141), .A(n5140), .ZN(n5144) );
  AOI21_X1 U6311 ( .B1(n5236), .B2(n5142), .A(n6609), .ZN(n5143) );
  AOI211_X1 U6312 ( .C1(EBX_REG_25__SCAN_IN), .C2(n5961), .A(n5144), .B(n5143), 
        .ZN(n5145) );
  OAI211_X1 U6313 ( .C1(n5652), .C2(n5968), .A(n5146), .B(n5145), .ZN(U2802)
         );
  AND2_X1 U6314 ( .A1(n5232), .A2(n5234), .ZN(n5148) );
  AND2_X2 U6315 ( .A1(n5148), .A2(n5147), .ZN(n5209) );
  AOI21_X2 U6316 ( .B1(n5150), .B2(n5149), .A(n5209), .ZN(n5507) );
  INV_X1 U6317 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5225) );
  OAI21_X1 U6318 ( .B1(n4488), .B2(n5152), .A(n5151), .ZN(n5219) );
  OAI222_X1 U6319 ( .A1(n5448), .A2(n5438), .B1(n5225), .B2(n5987), .C1(n5219), 
        .C2(n5433), .ZN(U2833) );
  INV_X1 U6320 ( .A(n5153), .ZN(n5159) );
  INV_X1 U6321 ( .A(n5154), .ZN(n5155) );
  OAI22_X1 U6322 ( .A1(n6531), .A2(n5157), .B1(n5156), .B2(n5155), .ZN(n5158)
         );
  AOI21_X1 U6323 ( .B1(n5159), .B2(n6635), .A(n5158), .ZN(n5163) );
  AOI21_X1 U6324 ( .B1(n6634), .B2(n5160), .A(n5162), .ZN(n5161) );
  OAI22_X1 U6325 ( .A1(n5163), .A2(n5162), .B1(n5161), .B2(n3425), .ZN(U3459)
         );
  INV_X1 U6326 ( .A(n5489), .ZN(n5165) );
  OAI22_X1 U6327 ( .A1(n5165), .A2(n5164), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5647), .ZN(n5167) );
  INV_X1 U6328 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5166) );
  XNOR2_X1 U6329 ( .A(n5167), .B(n5166), .ZN(n5634) );
  NAND2_X1 U6330 ( .A1(n5232), .A2(n5168), .ZN(n5207) );
  INV_X1 U6331 ( .A(n5207), .ZN(n5170) );
  NOR2_X1 U6332 ( .A1(n5178), .A2(n5599), .ZN(n5171) );
  INV_X1 U6333 ( .A(n5183), .ZN(n5175) );
  NAND2_X1 U6334 ( .A1(n6095), .A2(REIP_REG_28__SCAN_IN), .ZN(n5628) );
  OAI21_X1 U6335 ( .B1(n6112), .B2(n5172), .A(n5628), .ZN(n5173) );
  INV_X1 U6336 ( .A(n5173), .ZN(n5174) );
  NOR2_X1 U6337 ( .A1(n5171), .A2(n5176), .ZN(n5177) );
  OAI21_X1 U6338 ( .B1(n5634), .B2(n6100), .A(n5177), .ZN(U2958) );
  AND2_X1 U6339 ( .A1(n3010), .A2(n5179), .ZN(n5180) );
  OR2_X1 U6340 ( .A1(n5180), .A2(n5199), .ZN(n5190) );
  INV_X1 U6341 ( .A(n5190), .ZN(n5632) );
  INV_X1 U6342 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6615) );
  NOR2_X1 U6343 ( .A1(n5211), .A2(n6615), .ZN(n5182) );
  INV_X1 U6344 ( .A(n5181), .ZN(n5201) );
  MUX2_X1 U6345 ( .A(n5182), .B(n5201), .S(REIP_REG_28__SCAN_IN), .Z(n5186) );
  AOI22_X1 U6346 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n5960), .B1(n5948), 
        .B2(n5183), .ZN(n5184) );
  OAI21_X1 U6347 ( .B1(n5952), .B2(n5191), .A(n5184), .ZN(n5185) );
  AOI211_X1 U6348 ( .C1(n5632), .C2(n5927), .A(n5186), .B(n5185), .ZN(n5187)
         );
  OAI21_X1 U6349 ( .B1(n5178), .B2(n5899), .A(n5187), .ZN(U2799) );
  AOI22_X1 U6350 ( .A1(n5467), .A2(DATAI_28_), .B1(n5473), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5189) );
  NAND2_X1 U6351 ( .A1(n5468), .A2(DATAI_12_), .ZN(n5188) );
  OAI211_X1 U6352 ( .C1(n5178), .C2(n5477), .A(n5189), .B(n5188), .ZN(U2863)
         );
  OAI222_X1 U6353 ( .A1(n5178), .A2(n5438), .B1(n5191), .B2(n5987), .C1(n5190), 
        .C2(n5433), .ZN(U2831) );
  AOI22_X1 U6354 ( .A1(n5467), .A2(DATAI_30_), .B1(n5473), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5194) );
  NAND2_X1 U6355 ( .A1(n5468), .A2(DATAI_14_), .ZN(n5193) );
  OAI211_X1 U6356 ( .C1(n5192), .C2(n5477), .A(n5194), .B(n5193), .ZN(U2861)
         );
  OAI222_X1 U6357 ( .A1(n5438), .A2(n5192), .B1(n5433), .B2(n5196), .C1(n5195), 
        .C2(n5987), .ZN(U2829) );
  OAI21_X1 U6358 ( .B1(n5199), .B2(n5198), .A(n5197), .ZN(n5615) );
  NAND2_X1 U6359 ( .A1(n5487), .A2(n4228), .ZN(n5206) );
  OAI22_X1 U6360 ( .A1(n5484), .A2(n5908), .B1(n5965), .B2(n5483), .ZN(n5204)
         );
  MUX2_X1 U6361 ( .A(n5202), .B(n5201), .S(REIP_REG_29__SCAN_IN), .Z(n5203) );
  AOI211_X1 U6362 ( .C1(n5961), .C2(EBX_REG_29__SCAN_IN), .A(n5204), .B(n5203), 
        .ZN(n5205) );
  OAI211_X1 U6363 ( .C1(n5615), .C2(n5968), .A(n5206), .B(n5205), .ZN(U2798)
         );
  INV_X1 U6364 ( .A(n5210), .ZN(n5221) );
  INV_X1 U6365 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5413) );
  OAI22_X1 U6366 ( .A1(n5908), .A2(n5492), .B1(REIP_REG_27__SCAN_IN), .B2(
        n5211), .ZN(n5212) );
  AOI21_X1 U6367 ( .B1(n5494), .B2(n5948), .A(n5212), .ZN(n5213) );
  OAI21_X1 U6368 ( .B1(n5952), .B2(n5413), .A(n5213), .ZN(n5217) );
  NAND2_X1 U6369 ( .A1(n5151), .A2(n5214), .ZN(n5215) );
  NAND2_X1 U6370 ( .A1(n3010), .A2(n5215), .ZN(n5640) );
  NOR2_X1 U6371 ( .A1(n5640), .A2(n5968), .ZN(n5216) );
  OAI21_X1 U6372 ( .B1(n5496), .B2(n5899), .A(n5218), .ZN(U2800) );
  INV_X1 U6373 ( .A(n5219), .ZN(n5649) );
  NOR2_X1 U6374 ( .A1(n5220), .A2(n6609), .ZN(n5222) );
  OAI21_X1 U6375 ( .B1(REIP_REG_26__SCAN_IN), .B2(n5222), .A(n5221), .ZN(n5224) );
  AOI22_X1 U6376 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n5960), .B1(n5948), 
        .B2(n5503), .ZN(n5223) );
  OAI211_X1 U6377 ( .C1(n5225), .C2(n5952), .A(n5224), .B(n5223), .ZN(n5226)
         );
  AOI21_X1 U6378 ( .B1(n5649), .B2(n5927), .A(n5226), .ZN(n5227) );
  OAI21_X1 U6379 ( .B1(n5448), .B2(n5899), .A(n5227), .ZN(U2801) );
  OAI21_X1 U6380 ( .B1(n5256), .B2(n5229), .A(n5228), .ZN(n5231) );
  NAND2_X1 U6381 ( .A1(n5231), .A2(n5230), .ZN(n5671) );
  OAI21_X1 U6382 ( .B1(n5232), .B2(n5234), .A(n5233), .ZN(n5451) );
  INV_X1 U6383 ( .A(n5451), .ZN(n5517) );
  NAND2_X1 U6384 ( .A1(n5517), .A2(n4228), .ZN(n5240) );
  OAI22_X1 U6385 ( .A1(n5514), .A2(n5908), .B1(n5965), .B2(n5513), .ZN(n5238)
         );
  INV_X1 U6386 ( .A(n5260), .ZN(n5245) );
  AOI21_X1 U6387 ( .B1(n5245), .B2(n5243), .A(REIP_REG_23__SCAN_IN), .ZN(n5235) );
  NOR2_X1 U6388 ( .A1(n5236), .A2(n5235), .ZN(n5237) );
  AOI211_X1 U6389 ( .C1(n5961), .C2(EBX_REG_23__SCAN_IN), .A(n5238), .B(n5237), 
        .ZN(n5239) );
  OAI211_X1 U6390 ( .C1(n5671), .C2(n5968), .A(n5240), .B(n5239), .ZN(U2804)
         );
  AOI21_X1 U6391 ( .B1(n5242), .B2(n5241), .A(n5232), .ZN(n5415) );
  NAND2_X1 U6392 ( .A1(n5415), .A2(n4228), .ZN(n5252) );
  NAND2_X1 U6393 ( .A1(n5961), .A2(EBX_REG_22__SCAN_IN), .ZN(n5249) );
  NAND2_X1 U6394 ( .A1(n5960), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5248)
         );
  NAND2_X1 U6395 ( .A1(n5948), .A2(n5522), .ZN(n5247) );
  INV_X1 U6396 ( .A(n5243), .ZN(n5244) );
  OAI211_X1 U6397 ( .C1(REIP_REG_22__SCAN_IN), .C2(REIP_REG_21__SCAN_IN), .A(
        n5245), .B(n5244), .ZN(n5246) );
  NAND4_X1 U6398 ( .A1(n5249), .A2(n5248), .A3(n5247), .A4(n5246), .ZN(n5250)
         );
  AOI21_X1 U6399 ( .B1(n5272), .B2(REIP_REG_22__SCAN_IN), .A(n5250), .ZN(n5251) );
  OAI211_X1 U6400 ( .C1(n5416), .C2(n5968), .A(n5252), .B(n5251), .ZN(U2805)
         );
  OR2_X1 U6401 ( .A1(n5254), .A2(n5253), .ZN(n5255) );
  NAND2_X1 U6402 ( .A1(n5256), .A2(n5255), .ZN(n5684) );
  INV_X1 U6403 ( .A(n4454), .ZN(n5258) );
  OAI21_X1 U6404 ( .B1(n5258), .B2(n3713), .A(n5241), .ZN(n5530) );
  INV_X1 U6405 ( .A(n5530), .ZN(n5259) );
  NAND2_X1 U6406 ( .A1(n5259), .A2(n4228), .ZN(n5267) );
  INV_X1 U6407 ( .A(n5533), .ZN(n5264) );
  NAND2_X1 U6408 ( .A1(n5961), .A2(EBX_REG_21__SCAN_IN), .ZN(n5263) );
  NOR2_X1 U6409 ( .A1(n5260), .A2(REIP_REG_21__SCAN_IN), .ZN(n5261) );
  AOI21_X1 U6410 ( .B1(n5960), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n5261), 
        .ZN(n5262) );
  OAI211_X1 U6411 ( .C1(n5965), .C2(n5264), .A(n5263), .B(n5262), .ZN(n5265)
         );
  AOI21_X1 U6412 ( .B1(n5272), .B2(REIP_REG_21__SCAN_IN), .A(n5265), .ZN(n5266) );
  OAI211_X1 U6413 ( .C1(n5684), .C2(n5968), .A(n5267), .B(n5266), .ZN(U2806)
         );
  MUX2_X1 U6414 ( .A(n5282), .B(n5269), .S(n5268), .Z(n5271) );
  XNOR2_X1 U6415 ( .A(n5271), .B(n5270), .ZN(n5705) );
  INV_X1 U6416 ( .A(n5705), .ZN(n5279) );
  INV_X1 U6417 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5419) );
  OAI21_X1 U6418 ( .B1(REIP_REG_20__SCAN_IN), .B2(n5273), .A(n5272), .ZN(n5277) );
  INV_X1 U6419 ( .A(n5274), .ZN(n5275) );
  AOI22_X1 U6420 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n5960), .B1(n5948), 
        .B2(n5275), .ZN(n5276) );
  OAI211_X1 U6421 ( .C1(n5952), .C2(n5419), .A(n5277), .B(n5276), .ZN(n5278)
         );
  AOI21_X1 U6422 ( .B1(n5279), .B2(n5927), .A(n5278), .ZN(n5280) );
  OAI21_X1 U6423 ( .B1(n5458), .B2(n5899), .A(n5280), .ZN(U2807) );
  XNOR2_X1 U6424 ( .A(n5282), .B(n5269), .ZN(n5303) );
  OR2_X1 U6425 ( .A1(n5314), .A2(n5303), .ZN(n5301) );
  XNOR2_X1 U6426 ( .A(n5301), .B(n5283), .ZN(n5710) );
  NOR2_X1 U6427 ( .A1(n5284), .A2(n5285), .ZN(n5286) );
  OR2_X1 U6428 ( .A1(n4452), .A2(n5286), .ZN(n5541) );
  INV_X1 U6429 ( .A(n5541), .ZN(n5287) );
  NAND2_X1 U6430 ( .A1(n5287), .A2(n4228), .ZN(n5298) );
  INV_X1 U6431 ( .A(n5316), .ZN(n5296) );
  INV_X1 U6432 ( .A(n5537), .ZN(n5288) );
  AOI22_X1 U6433 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n5960), .B1(n5948), 
        .B2(n5288), .ZN(n5294) );
  NAND2_X1 U6434 ( .A1(n5961), .A2(EBX_REG_19__SCAN_IN), .ZN(n5293) );
  NAND2_X1 U6435 ( .A1(n5975), .A2(n5289), .ZN(n5918) );
  AOI21_X1 U6436 ( .B1(n6596), .B2(n6598), .A(n5290), .ZN(n5291) );
  NAND2_X1 U6437 ( .A1(n5291), .A2(n5305), .ZN(n5292) );
  NAND4_X1 U6438 ( .A1(n5294), .A2(n5293), .A3(n5918), .A4(n5292), .ZN(n5295)
         );
  AOI21_X1 U6439 ( .B1(n5296), .B2(REIP_REG_19__SCAN_IN), .A(n5295), .ZN(n5297) );
  OAI211_X1 U6440 ( .C1(n5710), .C2(n5968), .A(n5298), .B(n5297), .ZN(U2808)
         );
  AOI21_X1 U6441 ( .B1(n5300), .B2(n5299), .A(n5284), .ZN(n5548) );
  INV_X1 U6442 ( .A(n5548), .ZN(n5463) );
  INV_X1 U6443 ( .A(n5301), .ZN(n5302) );
  AOI21_X1 U6444 ( .B1(n5303), .B2(n5314), .A(n5302), .ZN(n5723) );
  AOI21_X1 U6445 ( .B1(n5948), .B2(n5544), .A(n5933), .ZN(n5304) );
  OAI21_X1 U6446 ( .B1(n5546), .B2(n5908), .A(n5304), .ZN(n5308) );
  AOI22_X1 U6447 ( .A1(EBX_REG_18__SCAN_IN), .A2(n5961), .B1(n5305), .B2(n6598), .ZN(n5306) );
  OAI21_X1 U6448 ( .B1(n5316), .B2(n6598), .A(n5306), .ZN(n5307) );
  AOI211_X1 U6449 ( .C1(n5723), .C2(n5927), .A(n5308), .B(n5307), .ZN(n5309)
         );
  OAI21_X1 U6450 ( .B1(n5463), .B2(n5899), .A(n5309), .ZN(U2809) );
  INV_X1 U6451 ( .A(n5299), .ZN(n5311) );
  AOI21_X1 U6452 ( .B1(n5312), .B2(n5310), .A(n5311), .ZN(n5557) );
  INV_X1 U6453 ( .A(n5557), .ZN(n5466) );
  OAI21_X1 U6454 ( .B1(n5313), .B2(n5315), .A(n5314), .ZN(n5422) );
  INV_X1 U6455 ( .A(n5422), .ZN(n5732) );
  AOI21_X1 U6456 ( .B1(n6594), .B2(n5317), .A(n5316), .ZN(n5320) );
  INV_X1 U6457 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5423) );
  INV_X1 U6458 ( .A(n5318), .ZN(n5555) );
  OAI21_X1 U6459 ( .B1(n5965), .B2(n5555), .A(n5918), .ZN(n5319) );
  OAI21_X1 U6460 ( .B1(n5321), .B2(n5322), .A(n5310), .ZN(n5562) );
  AOI21_X1 U6461 ( .B1(n5430), .B2(n5429), .A(n5323), .ZN(n5324) );
  OR2_X1 U6462 ( .A1(n5313), .A2(n5324), .ZN(n5744) );
  INV_X1 U6463 ( .A(n5744), .ZN(n5335) );
  INV_X1 U6464 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5328) );
  NOR3_X1 U6465 ( .A1(n5381), .A2(REIP_REG_16__SCAN_IN), .A3(n5325), .ZN(n5326) );
  AOI21_X1 U6466 ( .B1(n5948), .B2(n5565), .A(n5326), .ZN(n5327) );
  OAI21_X1 U6467 ( .B1(n5952), .B2(n5328), .A(n5327), .ZN(n5334) );
  INV_X1 U6468 ( .A(n5329), .ZN(n5331) );
  NOR2_X1 U6469 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5331), .ZN(n5330) );
  AND2_X1 U6470 ( .A1(n5939), .A2(n5330), .ZN(n5863) );
  NAND2_X1 U6471 ( .A1(n5939), .A2(n5331), .ZN(n5349) );
  NAND2_X1 U6472 ( .A1(n5349), .A2(n5975), .ZN(n5860) );
  OAI21_X1 U6473 ( .B1(n5863), .B2(n5860), .A(REIP_REG_16__SCAN_IN), .ZN(n5332) );
  OAI211_X1 U6474 ( .C1(n5908), .C2(n3042), .A(n5918), .B(n5332), .ZN(n5333)
         );
  AOI211_X1 U6475 ( .C1(n5335), .C2(n5927), .A(n5334), .B(n5333), .ZN(n5336)
         );
  OAI21_X1 U6476 ( .B1(n5562), .B2(n5899), .A(n5336), .ZN(U2811) );
  XOR2_X1 U6477 ( .A(n5339), .B(n5337), .Z(n5358) );
  INV_X1 U6478 ( .A(n5338), .ZN(n5357) );
  INV_X1 U6479 ( .A(n5339), .ZN(n5340) );
  NOR2_X1 U6480 ( .A1(n5337), .A2(n5340), .ZN(n5342) );
  OAI21_X1 U6481 ( .B1(n5356), .B2(n5342), .A(n5341), .ZN(n5428) );
  INV_X1 U6482 ( .A(n5428), .ZN(n5344) );
  NOR3_X1 U6483 ( .A1(n5356), .A2(n5342), .A3(n5341), .ZN(n5343) );
  NOR2_X1 U6484 ( .A1(n5344), .A2(n5343), .ZN(n5575) );
  INV_X1 U6485 ( .A(n5575), .ZN(n5475) );
  INV_X1 U6486 ( .A(n5573), .ZN(n5347) );
  INV_X1 U6487 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5432) );
  OAI22_X1 U6488 ( .A1(n5432), .A2(n5952), .B1(n5345), .B2(n5908), .ZN(n5346)
         );
  AOI211_X1 U6489 ( .C1(n5948), .C2(n5347), .A(n5346), .B(n5933), .ZN(n5348)
         );
  OAI21_X1 U6490 ( .B1(n5350), .B2(n5349), .A(n5348), .ZN(n5354) );
  INV_X1 U6491 ( .A(n5360), .ZN(n5764) );
  AOI21_X1 U6492 ( .B1(n5764), .B2(n5359), .A(n5351), .ZN(n5352) );
  OR2_X1 U6493 ( .A1(n5352), .A2(n5430), .ZN(n5805) );
  NOR2_X1 U6494 ( .A1(n5805), .A2(n5968), .ZN(n5353) );
  AOI211_X1 U6495 ( .C1(REIP_REG_14__SCAN_IN), .C2(n5860), .A(n5354), .B(n5353), .ZN(n5355) );
  OAI21_X1 U6496 ( .B1(n5475), .B2(n5899), .A(n5355), .ZN(U2813) );
  AOI21_X1 U6497 ( .B1(n5358), .B2(n5357), .A(n5356), .ZN(n5582) );
  XNOR2_X1 U6498 ( .A(n5360), .B(n5359), .ZN(n5825) );
  AOI22_X1 U6499 ( .A1(EBX_REG_13__SCAN_IN), .A2(n5961), .B1(n5927), .B2(n5825), .ZN(n5361) );
  OAI211_X1 U6500 ( .C1(n5908), .C2(n3037), .A(n5361), .B(n5918), .ZN(n5367)
         );
  NOR3_X1 U6501 ( .A1(n5381), .A2(REIP_REG_12__SCAN_IN), .A3(n5362), .ZN(n5870) );
  NAND2_X1 U6502 ( .A1(n5939), .A2(n5362), .ZN(n5371) );
  NAND2_X1 U6503 ( .A1(n5975), .A2(n5371), .ZN(n5871) );
  OAI21_X1 U6504 ( .B1(n5870), .B2(n5871), .A(REIP_REG_13__SCAN_IN), .ZN(n5365) );
  INV_X1 U6505 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6585) );
  NAND3_X1 U6506 ( .A1(n5939), .A2(n6585), .A3(n5363), .ZN(n5364) );
  OAI211_X1 U6507 ( .C1(n5965), .C2(n5579), .A(n5365), .B(n5364), .ZN(n5366)
         );
  AOI211_X1 U6508 ( .C1(n5582), .C2(n4228), .A(n5367), .B(n5366), .ZN(n5368)
         );
  INV_X1 U6509 ( .A(n5368), .ZN(U2814) );
  INV_X1 U6510 ( .A(n5369), .ZN(n5370) );
  OAI22_X1 U6511 ( .A1(n5371), .A2(n5370), .B1(n5593), .B2(n5965), .ZN(n5375)
         );
  AOI22_X1 U6512 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n5960), .B1(
        REIP_REG_11__SCAN_IN), .B2(n5871), .ZN(n5372) );
  OAI211_X1 U6513 ( .C1(n5952), .C2(n5373), .A(n5372), .B(n5918), .ZN(n5374)
         );
  AOI211_X1 U6514 ( .C1(n6114), .C2(n5927), .A(n5375), .B(n5374), .ZN(n5376)
         );
  OAI21_X1 U6515 ( .B1(n5899), .B2(n5598), .A(n5376), .ZN(U2816) );
  INV_X1 U6516 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6580) );
  INV_X1 U6517 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6578) );
  AND2_X1 U6518 ( .A1(REIP_REG_5__SCAN_IN), .A2(n5915), .ZN(n5377) );
  NOR3_X1 U6519 ( .A1(n6578), .A2(n6576), .A3(n5907), .ZN(n5891) );
  INV_X1 U6520 ( .A(n5891), .ZN(n5378) );
  NOR3_X1 U6521 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6580), .A3(n5378), .ZN(n5882)
         );
  AOI21_X1 U6522 ( .B1(n5960), .B2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n5933), 
        .ZN(n5383) );
  NAND2_X1 U6523 ( .A1(REIP_REG_7__SCAN_IN), .A2(REIP_REG_6__SCAN_IN), .ZN(
        n5903) );
  NOR2_X1 U6524 ( .A1(n6580), .A2(n5903), .ZN(n5380) );
  INV_X1 U6525 ( .A(n5975), .ZN(n5929) );
  OAI21_X1 U6526 ( .B1(n5929), .B2(n5379), .A(n5928), .ZN(n5916) );
  OAI21_X1 U6527 ( .B1(n5381), .B2(n5380), .A(n5916), .ZN(n5890) );
  AOI22_X1 U6528 ( .A1(EBX_REG_9__SCAN_IN), .A2(n5961), .B1(
        REIP_REG_9__SCAN_IN), .B2(n5890), .ZN(n5382) );
  OAI211_X1 U6529 ( .C1(n5968), .C2(n5384), .A(n5383), .B(n5382), .ZN(n5388)
         );
  OAI22_X1 U6530 ( .A1(n5386), .A2(n5899), .B1(n5385), .B2(n5965), .ZN(n5387)
         );
  OR3_X1 U6531 ( .A1(n5882), .A2(n5388), .A3(n5387), .ZN(U2818) );
  NAND2_X1 U6532 ( .A1(n5392), .A2(n3227), .ZN(n5389) );
  NAND2_X1 U6533 ( .A1(n5389), .A2(n5899), .ZN(n5971) );
  INV_X1 U6534 ( .A(n5971), .ZN(n5408) );
  INV_X1 U6535 ( .A(REIP_REG_1__SCAN_IN), .ZN(n5390) );
  NAND2_X1 U6536 ( .A1(n5939), .A2(n5390), .ZN(n5966) );
  NAND2_X1 U6537 ( .A1(n5966), .A2(n5975), .ZN(n5944) );
  NAND2_X1 U6538 ( .A1(n5392), .A2(n5391), .ZN(n5964) );
  INV_X1 U6539 ( .A(n5964), .ZN(n5405) );
  AOI22_X1 U6540 ( .A1(n5405), .A2(n4647), .B1(n5961), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n5399) );
  INV_X1 U6541 ( .A(n5393), .ZN(n5394) );
  AOI22_X1 U6542 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n5960), .B1(n5948), 
        .B2(n5394), .ZN(n5398) );
  NAND3_X1 U6543 ( .A1(n5939), .A2(REIP_REG_1__SCAN_IN), .A3(n6568), .ZN(n5397) );
  INV_X1 U6544 ( .A(n5982), .ZN(n5395) );
  NAND2_X1 U6545 ( .A1(n5927), .A2(n5395), .ZN(n5396) );
  NAND4_X1 U6546 ( .A1(n5399), .A2(n5398), .A3(n5397), .A4(n5396), .ZN(n5400)
         );
  AOI21_X1 U6547 ( .B1(REIP_REG_2__SCAN_IN), .B2(n5944), .A(n5400), .ZN(n5401)
         );
  OAI21_X1 U6548 ( .B1(n5983), .B2(n5408), .A(n5401), .ZN(U2825) );
  INV_X1 U6549 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n5402) );
  AOI21_X1 U6550 ( .B1(n5908), .B2(n5965), .A(n5402), .ZN(n5404) );
  OAI22_X1 U6551 ( .A1(n4006), .A2(n5952), .B1(n5968), .B2(n5780), .ZN(n5403)
         );
  AOI211_X1 U6552 ( .C1(n5405), .C2(n6495), .A(n5404), .B(n5403), .ZN(n5407)
         );
  NAND2_X1 U6553 ( .A1(n5928), .A2(REIP_REG_0__SCAN_IN), .ZN(n5406) );
  OAI211_X1 U6554 ( .C1(n5408), .C2(n5608), .A(n5407), .B(n5406), .ZN(U2827)
         );
  INV_X1 U6555 ( .A(n5409), .ZN(n5411) );
  OAI22_X1 U6556 ( .A1(n5411), .A2(n5433), .B1(n5987), .B2(n5410), .ZN(U2828)
         );
  INV_X1 U6557 ( .A(n5487), .ZN(n5443) );
  OAI222_X1 U6558 ( .A1(n5443), .A2(n5438), .B1(n5412), .B2(n5987), .C1(n5433), 
        .C2(n5615), .ZN(U2830) );
  OAI222_X1 U6559 ( .A1(n5496), .A2(n5438), .B1(n5413), .B2(n5987), .C1(n5640), 
        .C2(n5433), .ZN(U2832) );
  INV_X1 U6560 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5414) );
  OAI222_X1 U6561 ( .A1(n5451), .A2(n5438), .B1(n5414), .B2(n5987), .C1(n5671), 
        .C2(n5433), .ZN(U2836) );
  INV_X1 U6562 ( .A(n5415), .ZN(n5525) );
  INV_X1 U6563 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5417) );
  OAI222_X1 U6564 ( .A1(n5525), .A2(n5438), .B1(n5417), .B2(n5987), .C1(n5433), 
        .C2(n5416), .ZN(U2837) );
  INV_X1 U6565 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5418) );
  OAI222_X1 U6566 ( .A1(n5530), .A2(n5438), .B1(n5418), .B2(n5987), .C1(n5684), 
        .C2(n5433), .ZN(U2838) );
  OAI222_X1 U6567 ( .A1(n5458), .A2(n5438), .B1(n5419), .B2(n5987), .C1(n5705), 
        .C2(n5433), .ZN(U2839) );
  INV_X1 U6568 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5420) );
  OAI222_X1 U6569 ( .A1(n5541), .A2(n5438), .B1(n5420), .B2(n5987), .C1(n5710), 
        .C2(n5433), .ZN(U2840) );
  AOI22_X1 U6570 ( .A1(n5723), .A2(n5979), .B1(EBX_REG_18__SCAN_IN), .B2(n5436), .ZN(n5421) );
  OAI21_X1 U6571 ( .B1(n5463), .B2(n5438), .A(n5421), .ZN(U2841) );
  OAI222_X1 U6572 ( .A1(n5466), .A2(n5438), .B1(n5423), .B2(n5987), .C1(n5422), 
        .C2(n5433), .ZN(U2842) );
  OAI22_X1 U6573 ( .A1(n5744), .A2(n5433), .B1(n5328), .B2(n5987), .ZN(n5424)
         );
  INV_X1 U6574 ( .A(n5424), .ZN(n5425) );
  OAI21_X1 U6575 ( .B1(n5562), .B2(n5438), .A(n5425), .ZN(U2843) );
  INV_X1 U6576 ( .A(n5426), .ZN(n5427) );
  AOI21_X1 U6577 ( .B1(n5428), .B2(n5427), .A(n5321), .ZN(n5864) );
  INV_X1 U6578 ( .A(n5864), .ZN(n5472) );
  XOR2_X1 U6579 ( .A(n5430), .B(n5429), .Z(n5865) );
  AOI22_X1 U6580 ( .A1(n5865), .A2(n5979), .B1(EBX_REG_15__SCAN_IN), .B2(n5436), .ZN(n5431) );
  OAI21_X1 U6581 ( .B1(n5472), .B2(n5438), .A(n5431), .ZN(U2844) );
  OAI22_X1 U6582 ( .A1(n5805), .A2(n5433), .B1(n5432), .B2(n5987), .ZN(n5434)
         );
  AOI21_X1 U6583 ( .B1(n5575), .B2(n5980), .A(n5434), .ZN(n5435) );
  INV_X1 U6584 ( .A(n5435), .ZN(U2845) );
  INV_X1 U6585 ( .A(n5582), .ZN(n5478) );
  AOI22_X1 U6586 ( .A1(n5825), .A2(n5979), .B1(EBX_REG_13__SCAN_IN), .B2(n5436), .ZN(n5437) );
  OAI21_X1 U6587 ( .B1(n5478), .B2(n5438), .A(n5437), .ZN(U2846) );
  NAND3_X1 U6588 ( .A1(n2957), .A2(n3231), .A3(n5991), .ZN(n5440) );
  AOI22_X1 U6589 ( .A1(n5467), .A2(DATAI_31_), .B1(n5473), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n5439) );
  NAND2_X1 U6590 ( .A1(n5440), .A2(n5439), .ZN(U2860) );
  AOI22_X1 U6591 ( .A1(n5467), .A2(DATAI_29_), .B1(n5473), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5442) );
  NAND2_X1 U6592 ( .A1(n5468), .A2(DATAI_13_), .ZN(n5441) );
  OAI211_X1 U6593 ( .C1(n5443), .C2(n5477), .A(n5442), .B(n5441), .ZN(U2862)
         );
  AOI22_X1 U6594 ( .A1(n5467), .A2(DATAI_27_), .B1(n5473), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5445) );
  NAND2_X1 U6595 ( .A1(n5468), .A2(DATAI_11_), .ZN(n5444) );
  OAI211_X1 U6596 ( .C1(n5496), .C2(n5477), .A(n5445), .B(n5444), .ZN(U2864)
         );
  AOI22_X1 U6597 ( .A1(n5467), .A2(DATAI_26_), .B1(n5473), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U6598 ( .A1(n5468), .A2(DATAI_10_), .ZN(n5446) );
  OAI211_X1 U6599 ( .C1(n5448), .C2(n5477), .A(n5447), .B(n5446), .ZN(U2865)
         );
  AOI22_X1 U6600 ( .A1(n5467), .A2(DATAI_23_), .B1(n5473), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5450) );
  NAND2_X1 U6601 ( .A1(n5468), .A2(DATAI_7_), .ZN(n5449) );
  OAI211_X1 U6602 ( .C1(n5451), .C2(n5477), .A(n5450), .B(n5449), .ZN(U2868)
         );
  AOI22_X1 U6603 ( .A1(n5467), .A2(DATAI_22_), .B1(n5473), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5453) );
  NAND2_X1 U6604 ( .A1(n5468), .A2(DATAI_6_), .ZN(n5452) );
  OAI211_X1 U6605 ( .C1(n5525), .C2(n5477), .A(n5453), .B(n5452), .ZN(U2869)
         );
  AOI22_X1 U6606 ( .A1(n5467), .A2(DATAI_21_), .B1(n5473), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5455) );
  NAND2_X1 U6607 ( .A1(n5468), .A2(DATAI_5_), .ZN(n5454) );
  OAI211_X1 U6608 ( .C1(n5530), .C2(n5477), .A(n5455), .B(n5454), .ZN(U2870)
         );
  AOI22_X1 U6609 ( .A1(n5467), .A2(DATAI_20_), .B1(n5473), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5457) );
  NAND2_X1 U6610 ( .A1(n5468), .A2(DATAI_4_), .ZN(n5456) );
  OAI211_X1 U6611 ( .C1(n5458), .C2(n5477), .A(n5457), .B(n5456), .ZN(U2871)
         );
  AOI22_X1 U6612 ( .A1(n5467), .A2(DATAI_19_), .B1(n5473), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5460) );
  NAND2_X1 U6613 ( .A1(n5468), .A2(DATAI_3_), .ZN(n5459) );
  OAI211_X1 U6614 ( .C1(n5541), .C2(n5477), .A(n5460), .B(n5459), .ZN(U2872)
         );
  AOI22_X1 U6615 ( .A1(n5467), .A2(DATAI_18_), .B1(n5473), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5462) );
  NAND2_X1 U6616 ( .A1(n5468), .A2(DATAI_2_), .ZN(n5461) );
  OAI211_X1 U6617 ( .C1(n5463), .C2(n5477), .A(n5462), .B(n5461), .ZN(U2873)
         );
  AOI22_X1 U6618 ( .A1(n5467), .A2(DATAI_17_), .B1(n5473), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5465) );
  NAND2_X1 U6619 ( .A1(n5468), .A2(DATAI_1_), .ZN(n5464) );
  OAI211_X1 U6620 ( .C1(n5466), .C2(n5477), .A(n5465), .B(n5464), .ZN(U2874)
         );
  AOI22_X1 U6621 ( .A1(n5467), .A2(DATAI_16_), .B1(n5473), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U6622 ( .A1(n5468), .A2(DATAI_0_), .ZN(n5469) );
  OAI211_X1 U6623 ( .C1(n5562), .C2(n5477), .A(n5470), .B(n5469), .ZN(U2875)
         );
  AOI22_X1 U6624 ( .A1(n5988), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n5473), .ZN(n5471) );
  OAI21_X1 U6625 ( .B1(n5472), .B2(n5477), .A(n5471), .ZN(U2876) );
  AOI22_X1 U6626 ( .A1(n5988), .A2(DATAI_14_), .B1(EAX_REG_14__SCAN_IN), .B2(
        n5473), .ZN(n5474) );
  OAI21_X1 U6627 ( .B1(n5475), .B2(n5477), .A(n5474), .ZN(U2877) );
  INV_X1 U6628 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6008) );
  OAI222_X1 U6629 ( .A1(n5478), .A2(n5477), .B1(n5476), .B2(n6084), .C1(n6008), 
        .C2(n5991), .ZN(U2878) );
  INV_X1 U6630 ( .A(n5617), .ZN(n5479) );
  NOR2_X1 U6631 ( .A1(n5489), .A2(n5479), .ZN(n5480) );
  NOR2_X1 U6632 ( .A1(n5481), .A2(n5480), .ZN(n5482) );
  XNOR2_X1 U6633 ( .A(n5482), .B(n5620), .ZN(n5625) );
  NOR2_X1 U6634 ( .A1(n5594), .A2(n5483), .ZN(n5486) );
  NAND2_X1 U6635 ( .A1(n6095), .A2(REIP_REG_29__SCAN_IN), .ZN(n5618) );
  OAI21_X1 U6636 ( .B1(n6112), .B2(n5484), .A(n5618), .ZN(n5485) );
  AOI211_X1 U6637 ( .C1(n5487), .C2(n6104), .A(n5486), .B(n5485), .ZN(n5488)
         );
  OAI21_X1 U6638 ( .B1(n5625), .B2(n6100), .A(n5488), .ZN(U2957) );
  OAI21_X1 U6639 ( .B1(n5490), .B2(n5499), .A(n5489), .ZN(n5491) );
  XNOR2_X1 U6640 ( .A(n5491), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5643)
         );
  NAND2_X1 U6641 ( .A1(n6095), .A2(REIP_REG_27__SCAN_IN), .ZN(n5635) );
  OAI21_X1 U6642 ( .B1(n6112), .B2(n5492), .A(n5635), .ZN(n5493) );
  OAI21_X1 U6643 ( .B1(n5643), .B2(n6100), .A(n5498), .ZN(U2959) );
  NOR2_X1 U6644 ( .A1(n4462), .A2(n5500), .ZN(n5502) );
  XOR2_X1 U6645 ( .A(n5502), .B(n5501), .Z(n5651) );
  NAND2_X1 U6646 ( .A1(n6105), .A2(n5503), .ZN(n5504) );
  NAND2_X1 U6647 ( .A1(n6095), .A2(REIP_REG_26__SCAN_IN), .ZN(n5645) );
  OAI211_X1 U6648 ( .C1(n6112), .C2(n5505), .A(n5504), .B(n5645), .ZN(n5506)
         );
  AOI21_X1 U6649 ( .B1(n5507), .B2(n6104), .A(n5506), .ZN(n5508) );
  OAI21_X1 U6650 ( .B1(n5651), .B2(n6100), .A(n5508), .ZN(U2960) );
  NAND3_X1 U6651 ( .A1(n5509), .A2(n5676), .A3(n2991), .ZN(n5510) );
  NAND2_X1 U6652 ( .A1(n5511), .A2(n5510), .ZN(n5512) );
  XNOR2_X1 U6653 ( .A(n5512), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5679)
         );
  NOR2_X1 U6654 ( .A1(n5594), .A2(n5513), .ZN(n5516) );
  NAND2_X1 U6655 ( .A1(n6095), .A2(REIP_REG_23__SCAN_IN), .ZN(n5670) );
  OAI21_X1 U6656 ( .B1(n6112), .B2(n5514), .A(n5670), .ZN(n5515) );
  AOI211_X1 U6657 ( .C1(n5517), .C2(n6104), .A(n5516), .B(n5515), .ZN(n5518)
         );
  OAI21_X1 U6658 ( .B1(n5679), .B2(n6100), .A(n5518), .ZN(U2963) );
  NAND2_X1 U6659 ( .A1(n5519), .A2(n6107), .ZN(n5524) );
  NOR2_X1 U6660 ( .A1(n6112), .A2(n3034), .ZN(n5520) );
  AOI211_X1 U6661 ( .C1(n6105), .C2(n5522), .A(n5521), .B(n5520), .ZN(n5523)
         );
  OAI211_X1 U6662 ( .C1(n5599), .C2(n5525), .A(n5524), .B(n5523), .ZN(U2964)
         );
  AOI21_X1 U6663 ( .B1(n5528), .B2(n5527), .A(n5526), .ZN(n5688) );
  NAND2_X1 U6664 ( .A1(n6095), .A2(REIP_REG_21__SCAN_IN), .ZN(n5683) );
  OAI21_X1 U6665 ( .B1(n6112), .B2(n5529), .A(n5683), .ZN(n5532) );
  NOR2_X1 U6666 ( .A1(n5530), .A2(n5599), .ZN(n5531) );
  AOI211_X1 U6667 ( .C1(n6105), .C2(n5533), .A(n5532), .B(n5531), .ZN(n5534)
         );
  OAI21_X1 U6668 ( .B1(n5688), .B2(n6100), .A(n5534), .ZN(U2965) );
  XNOR2_X1 U6669 ( .A(n2991), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5535)
         );
  XNOR2_X1 U6670 ( .A(n5536), .B(n5535), .ZN(n5709) );
  NAND2_X1 U6671 ( .A1(n5709), .A2(n6107), .ZN(n5540) );
  NOR2_X1 U6672 ( .A1(n6122), .A2(n6596), .ZN(n5712) );
  NOR2_X1 U6673 ( .A1(n5594), .A2(n5537), .ZN(n5538) );
  AOI211_X1 U6674 ( .C1(n6094), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n5712), 
        .B(n5538), .ZN(n5539) );
  OAI211_X1 U6675 ( .C1(n5599), .C2(n5541), .A(n5540), .B(n5539), .ZN(U2967)
         );
  NAND3_X1 U6676 ( .A1(n5561), .A2(n5587), .A3(n5729), .ZN(n5552) );
  OAI22_X1 U6677 ( .A1(n5552), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .B1(n5587), .B2(n5542), .ZN(n5543) );
  XNOR2_X1 U6678 ( .A(n5543), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5725)
         );
  NAND2_X1 U6679 ( .A1(n6105), .A2(n5544), .ZN(n5545) );
  NAND2_X1 U6680 ( .A1(n6095), .A2(REIP_REG_18__SCAN_IN), .ZN(n5717) );
  OAI211_X1 U6681 ( .C1(n6112), .C2(n5546), .A(n5545), .B(n5717), .ZN(n5547)
         );
  AOI21_X1 U6682 ( .B1(n5548), .B2(n6104), .A(n5547), .ZN(n5549) );
  OAI21_X1 U6683 ( .B1(n5725), .B2(n6100), .A(n5549), .ZN(U2968) );
  NAND3_X1 U6684 ( .A1(n5550), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n2992), .ZN(n5551) );
  NAND2_X1 U6685 ( .A1(n5552), .A2(n5551), .ZN(n5553) );
  XNOR2_X1 U6686 ( .A(n5553), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5734)
         );
  NAND2_X1 U6687 ( .A1(n6094), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5554)
         );
  NAND2_X1 U6688 ( .A1(n6095), .A2(REIP_REG_17__SCAN_IN), .ZN(n5726) );
  OAI211_X1 U6689 ( .C1(n5594), .C2(n5555), .A(n5554), .B(n5726), .ZN(n5556)
         );
  AOI21_X1 U6690 ( .B1(n5557), .B2(n6104), .A(n5556), .ZN(n5558) );
  OAI21_X1 U6691 ( .B1(n5734), .B2(n6100), .A(n5558), .ZN(U2969) );
  OAI21_X1 U6692 ( .B1(n5729), .B2(n2992), .A(n5559), .ZN(n5560) );
  XNOR2_X1 U6693 ( .A(n5561), .B(n5560), .ZN(n5749) );
  NAND2_X1 U6694 ( .A1(n6095), .A2(REIP_REG_16__SCAN_IN), .ZN(n5743) );
  OAI21_X1 U6695 ( .B1(n6112), .B2(n3042), .A(n5743), .ZN(n5564) );
  NOR2_X1 U6696 ( .A1(n5562), .A2(n5599), .ZN(n5563) );
  AOI211_X1 U6697 ( .C1(n6105), .C2(n5565), .A(n5564), .B(n5563), .ZN(n5566)
         );
  OAI21_X1 U6698 ( .B1(n5749), .B2(n6100), .A(n5566), .ZN(U2970) );
  INV_X1 U6699 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5761) );
  AOI21_X1 U6700 ( .B1(n2992), .B2(n5761), .A(n5567), .ZN(n5577) );
  XNOR2_X1 U6701 ( .A(n5587), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5578)
         );
  OAI22_X1 U6702 ( .A1(n5577), .A2(n5578), .B1(n5587), .B2(
        INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5571) );
  OAI21_X1 U6703 ( .B1(n2992), .B2(n5569), .A(n5568), .ZN(n5570) );
  XNOR2_X1 U6704 ( .A(n5571), .B(n5570), .ZN(n5804) );
  AOI22_X1 U6705 ( .A1(n6094), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n6095), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n5572) );
  OAI21_X1 U6706 ( .B1(n5573), .B2(n5594), .A(n5572), .ZN(n5574) );
  AOI21_X1 U6707 ( .B1(n5575), .B2(n6104), .A(n5574), .ZN(n5576) );
  OAI21_X1 U6708 ( .B1(n5804), .B2(n6100), .A(n5576), .ZN(U2972) );
  XOR2_X1 U6709 ( .A(n5578), .B(n5577), .Z(n5826) );
  NOR2_X1 U6710 ( .A1(n5594), .A2(n5579), .ZN(n5581) );
  NAND2_X1 U6711 ( .A1(n6095), .A2(REIP_REG_13__SCAN_IN), .ZN(n5823) );
  OAI21_X1 U6712 ( .B1(n6112), .B2(n3037), .A(n5823), .ZN(n5580) );
  AOI211_X1 U6713 ( .C1(n5582), .C2(n6104), .A(n5581), .B(n5580), .ZN(n5583)
         );
  OAI21_X1 U6714 ( .B1(n5826), .B2(n6100), .A(n5583), .ZN(U2973) );
  INV_X1 U6715 ( .A(n5584), .ZN(n5585) );
  OAI21_X1 U6716 ( .B1(n2992), .B2(n5773), .A(n5585), .ZN(n5604) );
  INV_X1 U6717 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5586) );
  NAND2_X1 U6718 ( .A1(n2992), .A2(n5586), .ZN(n5600) );
  AND2_X1 U6719 ( .A1(n5587), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5602)
         );
  AOI21_X1 U6720 ( .B1(n5604), .B2(n5600), .A(n5602), .ZN(n5591) );
  OR2_X1 U6721 ( .A1(n2992), .A2(n5588), .ZN(n5758) );
  NAND2_X1 U6722 ( .A1(n2992), .A2(n5588), .ZN(n5589) );
  NAND2_X1 U6723 ( .A1(n5758), .A2(n5589), .ZN(n5590) );
  NOR2_X1 U6724 ( .A1(n5591), .A2(n5590), .ZN(n5760) );
  AOI21_X1 U6725 ( .B1(n5591), .B2(n5590), .A(n5760), .ZN(n6116) );
  NAND2_X1 U6726 ( .A1(n6116), .A2(n6107), .ZN(n5597) );
  INV_X1 U6727 ( .A(REIP_REG_11__SCAN_IN), .ZN(n5592) );
  NOR2_X1 U6728 ( .A1(n6122), .A2(n5592), .ZN(n6113) );
  NOR2_X1 U6729 ( .A1(n5594), .A2(n5593), .ZN(n5595) );
  AOI211_X1 U6730 ( .C1(n6094), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6113), 
        .B(n5595), .ZN(n5596) );
  OAI211_X1 U6731 ( .C1(n5599), .C2(n5598), .A(n5597), .B(n5596), .ZN(U2975)
         );
  INV_X1 U6732 ( .A(n5600), .ZN(n5601) );
  NOR2_X1 U6733 ( .A1(n5602), .A2(n5601), .ZN(n5603) );
  XNOR2_X1 U6734 ( .A(n5604), .B(n5603), .ZN(n5779) );
  NOR2_X1 U6735 ( .A1(n6122), .A2(n6583), .ZN(n5776) );
  AND2_X1 U6736 ( .A1(n6094), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5605)
         );
  AOI211_X1 U6737 ( .C1(n6105), .C2(n5880), .A(n5776), .B(n5605), .ZN(n5607)
         );
  NAND2_X1 U6738 ( .A1(n5881), .A2(n6104), .ZN(n5606) );
  OAI211_X1 U6739 ( .C1(n5779), .C2(n6100), .A(n5607), .B(n5606), .ZN(U2976)
         );
  INV_X1 U6740 ( .A(n5608), .ZN(n5609) );
  NAND2_X1 U6741 ( .A1(n5609), .A2(n6104), .ZN(n5614) );
  OR2_X1 U6742 ( .A1(n5610), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5787)
         );
  NAND3_X1 U6743 ( .A1(n5787), .A2(n4141), .A3(n6107), .ZN(n5613) );
  NAND2_X1 U6744 ( .A1(n6095), .A2(REIP_REG_0__SCAN_IN), .ZN(n5781) );
  OAI21_X1 U6745 ( .B1(n6094), .B2(n5611), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5612) );
  NAND4_X1 U6746 ( .A1(n5614), .A2(n5613), .A3(n5781), .A4(n5612), .ZN(U2986)
         );
  INV_X1 U6747 ( .A(n5615), .ZN(n5623) );
  INV_X1 U6748 ( .A(n5616), .ZN(n5621) );
  INV_X1 U6749 ( .A(n5630), .ZN(n5639) );
  NAND3_X1 U6750 ( .A1(n5639), .A2(n5617), .A3(n5620), .ZN(n5619) );
  OAI211_X1 U6751 ( .C1(n5621), .C2(n5620), .A(n5619), .B(n5618), .ZN(n5622)
         );
  AOI21_X1 U6752 ( .B1(n5623), .B2(n6138), .A(n5622), .ZN(n5624) );
  OAI21_X1 U6753 ( .B1(n5625), .B2(n6142), .A(n5624), .ZN(U2989) );
  XNOR2_X1 U6754 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .B(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5629) );
  INV_X1 U6755 ( .A(n5636), .ZN(n5626) );
  NAND2_X1 U6756 ( .A1(n5626), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5627) );
  OAI211_X1 U6757 ( .C1(n5630), .C2(n5629), .A(n5628), .B(n5627), .ZN(n5631)
         );
  AOI21_X1 U6758 ( .B1(n5632), .B2(n6138), .A(n5631), .ZN(n5633) );
  OAI21_X1 U6759 ( .B1(n5634), .B2(n6142), .A(n5633), .ZN(U2990) );
  OAI21_X1 U6760 ( .B1(n5636), .B2(n5638), .A(n5635), .ZN(n5637) );
  AOI21_X1 U6761 ( .B1(n5639), .B2(n5638), .A(n5637), .ZN(n5642) );
  OR2_X1 U6762 ( .A1(n5640), .A2(n6149), .ZN(n5641) );
  OAI211_X1 U6763 ( .C1(n5643), .C2(n6142), .A(n5642), .B(n5641), .ZN(U2991)
         );
  OAI211_X1 U6764 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5657), .B(n5644), .ZN(n5646) );
  OAI211_X1 U6765 ( .C1(n5662), .C2(n5647), .A(n5646), .B(n5645), .ZN(n5648)
         );
  AOI21_X1 U6766 ( .B1(n5649), .B2(n6138), .A(n5648), .ZN(n5650) );
  OAI21_X1 U6767 ( .B1(n5651), .B2(n6142), .A(n5650), .ZN(U2992) );
  INV_X1 U6768 ( .A(n5652), .ZN(n5655) );
  OAI21_X1 U6769 ( .B1(n5662), .B2(n5656), .A(n5653), .ZN(n5654) );
  AOI21_X1 U6770 ( .B1(n5655), .B2(n6138), .A(n5654), .ZN(n5659) );
  NAND2_X1 U6771 ( .A1(n5657), .A2(n5656), .ZN(n5658) );
  OAI211_X1 U6772 ( .C1(n5660), .C2(n6142), .A(n5659), .B(n5658), .ZN(U2993)
         );
  INV_X1 U6773 ( .A(n5661), .ZN(n5666) );
  NAND3_X1 U6774 ( .A1(n5702), .A2(n5676), .A3(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5664) );
  AOI21_X1 U6775 ( .B1(n5664), .B2(n5663), .A(n5662), .ZN(n5665) );
  AOI211_X1 U6776 ( .C1(n5667), .C2(n6138), .A(n5666), .B(n5665), .ZN(n5668)
         );
  OAI21_X1 U6777 ( .B1(n5669), .B2(n6142), .A(n5668), .ZN(U2994) );
  INV_X1 U6778 ( .A(n5670), .ZN(n5673) );
  NOR2_X1 U6779 ( .A1(n5671), .A2(n6149), .ZN(n5672) );
  AOI211_X1 U6780 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n5674), .A(n5673), .B(n5672), .ZN(n5678) );
  NAND3_X1 U6781 ( .A1(n5702), .A2(n5676), .A3(n5675), .ZN(n5677) );
  OAI211_X1 U6782 ( .C1(n5679), .C2(n6142), .A(n5678), .B(n5677), .ZN(U2995)
         );
  INV_X1 U6783 ( .A(n5680), .ZN(n5686) );
  NAND2_X1 U6784 ( .A1(n5681), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5682) );
  OAI211_X1 U6785 ( .C1(n5684), .C2(n6149), .A(n5683), .B(n5682), .ZN(n5685)
         );
  AOI21_X1 U6786 ( .B1(n5686), .B2(n4232), .A(n5685), .ZN(n5687) );
  OAI21_X1 U6787 ( .B1(n5688), .B2(n6142), .A(n5687), .ZN(U2997) );
  INV_X1 U6788 ( .A(n5689), .ZN(n5690) );
  OR2_X1 U6789 ( .A1(n5735), .A2(n5690), .ZN(n5693) );
  NAND2_X1 U6790 ( .A1(n5737), .A2(n5691), .ZN(n5692) );
  AND2_X1 U6791 ( .A1(n5693), .A2(n5692), .ZN(n5728) );
  OR2_X1 U6792 ( .A1(n5694), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5695)
         );
  AND2_X1 U6793 ( .A1(n5728), .A2(n5695), .ZN(n5719) );
  NAND2_X1 U6794 ( .A1(n5696), .A2(n5718), .ZN(n5697) );
  NAND2_X1 U6795 ( .A1(n5719), .A2(n5697), .ZN(n5713) );
  AOI21_X1 U6796 ( .B1(n5713), .B2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5698), 
        .ZN(n5704) );
  NOR2_X1 U6797 ( .A1(n5700), .A2(n5699), .ZN(n5701) );
  NAND2_X1 U6798 ( .A1(n5702), .A2(n5701), .ZN(n5703) );
  OAI211_X1 U6799 ( .C1(n5705), .C2(n6149), .A(n5704), .B(n5703), .ZN(n5706)
         );
  AOI21_X1 U6800 ( .B1(n5707), .B2(n6155), .A(n5706), .ZN(n5708) );
  INV_X1 U6801 ( .A(n5708), .ZN(U2998) );
  NAND2_X1 U6802 ( .A1(n5709), .A2(n6155), .ZN(n5715) );
  NOR2_X1 U6803 ( .A1(n5710), .A2(n6149), .ZN(n5711) );
  AOI211_X1 U6804 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n5713), .A(n5712), .B(n5711), .ZN(n5714) );
  OAI211_X1 U6805 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n5716), .A(n5715), .B(n5714), .ZN(U2999) );
  OAI21_X1 U6806 ( .B1(n5719), .B2(n5718), .A(n5717), .ZN(n5722) );
  NOR3_X1 U6807 ( .A1(n6119), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n5720), 
        .ZN(n5721) );
  AOI211_X1 U6808 ( .C1(n6138), .C2(n5723), .A(n5722), .B(n5721), .ZN(n5724)
         );
  OAI21_X1 U6809 ( .B1(n5725), .B2(n6142), .A(n5724), .ZN(U3000) );
  OAI21_X1 U6810 ( .B1(n5728), .B2(n5727), .A(n5726), .ZN(n5731) );
  NOR4_X1 U6811 ( .A1(n6119), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5729), 
        .A4(n5745), .ZN(n5730) );
  AOI211_X1 U6812 ( .C1(n6138), .C2(n5732), .A(n5731), .B(n5730), .ZN(n5733)
         );
  OAI21_X1 U6813 ( .B1(n5734), .B2(n6142), .A(n5733), .ZN(U3001) );
  OR2_X1 U6814 ( .A1(n5808), .A2(n5735), .ZN(n5739) );
  NAND2_X1 U6815 ( .A1(n5737), .A2(n5736), .ZN(n5738) );
  NAND2_X1 U6816 ( .A1(n5739), .A2(n5738), .ZN(n6115) );
  INV_X1 U6817 ( .A(n6115), .ZN(n5741) );
  INV_X1 U6818 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5740) );
  NAND3_X1 U6819 ( .A1(n5816), .A2(n5742), .A3(n5740), .ZN(n5753) );
  OAI211_X1 U6820 ( .C1(n5742), .C2(n6153), .A(n5741), .B(n5753), .ZN(n5754)
         );
  OAI21_X1 U6821 ( .B1(n5744), .B2(n6149), .A(n5743), .ZN(n5747) );
  NOR3_X1 U6822 ( .A1(n6119), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5745), 
        .ZN(n5746) );
  AOI211_X1 U6823 ( .C1(INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n5754), .A(n5747), .B(n5746), .ZN(n5748) );
  OAI21_X1 U6824 ( .B1(n5749), .B2(n6142), .A(n5748), .ZN(U3002) );
  NAND2_X1 U6825 ( .A1(n3017), .A2(n5751), .ZN(n5752) );
  XNOR2_X1 U6826 ( .A(n5750), .B(n5752), .ZN(n5800) );
  AOI22_X1 U6827 ( .A1(n5865), .A2(n6138), .B1(n6095), .B2(
        REIP_REG_15__SCAN_IN), .ZN(n5757) );
  INV_X1 U6828 ( .A(n5753), .ZN(n5755) );
  OAI21_X1 U6829 ( .B1(n5755), .B2(INSTADDRPOINTER_REG_15__SCAN_IN), .A(n5754), 
        .ZN(n5756) );
  OAI211_X1 U6830 ( .C1(n5800), .C2(n6142), .A(n5757), .B(n5756), .ZN(U3003)
         );
  INV_X1 U6831 ( .A(n5758), .ZN(n5759) );
  NOR2_X1 U6832 ( .A1(n5760), .A2(n5759), .ZN(n5763) );
  XNOR2_X1 U6833 ( .A(n2992), .B(n5761), .ZN(n5762) );
  XNOR2_X1 U6834 ( .A(n5763), .B(n5762), .ZN(n6101) );
  AOI21_X1 U6835 ( .B1(n5765), .B2(n5041), .A(n5764), .ZN(n5976) );
  AOI22_X1 U6836 ( .A1(n5976), .A2(n6138), .B1(n6095), .B2(
        REIP_REG_12__SCAN_IN), .ZN(n5771) );
  AOI221_X1 U6837 ( .B1(n5767), .B2(n5822), .C1(n5766), .C2(n5822), .A(n6115), 
        .ZN(n5769) );
  AOI21_X1 U6838 ( .B1(n5816), .B2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5768) );
  OR2_X1 U6839 ( .A1(n5769), .A2(n5768), .ZN(n5770) );
  OAI211_X1 U6840 ( .C1(n6101), .C2(n6142), .A(n5771), .B(n5770), .ZN(U3006)
         );
  AOI221_X1 U6841 ( .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n5586), .C2(n5773), .A(n5772), 
        .ZN(n5774) );
  AOI21_X1 U6842 ( .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n5775), .A(n5774), 
        .ZN(n5778) );
  AOI21_X1 U6843 ( .B1(n5877), .B2(n6138), .A(n5776), .ZN(n5777) );
  OAI211_X1 U6844 ( .C1(n5779), .C2(n6142), .A(n5778), .B(n5777), .ZN(U3008)
         );
  INV_X1 U6845 ( .A(n5780), .ZN(n5784) );
  INV_X1 U6846 ( .A(n5781), .ZN(n5783) );
  AOI211_X1 U6847 ( .C1(n6138), .C2(n5784), .A(n5783), .B(n5782), .ZN(n5790)
         );
  INV_X1 U6848 ( .A(n5814), .ZN(n5786) );
  OAI21_X1 U6849 ( .B1(n5786), .B2(n5785), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5789) );
  NAND3_X1 U6850 ( .A1(n5787), .A2(n4141), .A3(n6155), .ZN(n5788) );
  NAND3_X1 U6851 ( .A1(n5790), .A2(n5789), .A3(n5788), .ZN(U3018) );
  OAI211_X1 U6852 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n4652), .A(n6381), .B(
        n6380), .ZN(n5791) );
  OAI21_X1 U6853 ( .B1(n5794), .B2(n5963), .A(n5791), .ZN(n5792) );
  MUX2_X1 U6854 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5792), .S(n6161), 
        .Z(U3464) );
  XNOR2_X1 U6855 ( .A(n5793), .B(n6381), .ZN(n5796) );
  OAI22_X1 U6856 ( .A1(n5796), .A2(n6435), .B1(n5795), .B2(n5794), .ZN(n5797)
         );
  MUX2_X1 U6857 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5797), .S(n6161), 
        .Z(U3463) );
  AOI22_X1 U6858 ( .A1(n6095), .A2(REIP_REG_15__SCAN_IN), .B1(n6094), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5799) );
  AOI22_X1 U6859 ( .A1(n5864), .A2(n6104), .B1(n5866), .B2(n6105), .ZN(n5798)
         );
  OAI211_X1 U6860 ( .C1(n6100), .C2(n5800), .A(n5799), .B(n5798), .ZN(U2971)
         );
  AND2_X1 U6861 ( .A1(n6033), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI21_X1 U6862 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(n5802), .A(n5801), .ZN(
        n5803) );
  INV_X1 U6863 ( .A(n5803), .ZN(U2788) );
  INV_X1 U6864 ( .A(n5804), .ZN(n5807) );
  INV_X1 U6865 ( .A(n5805), .ZN(n5806) );
  AOI22_X1 U6866 ( .A1(n5807), .A2(n6155), .B1(n6138), .B2(n5806), .ZN(n5821)
         );
  NAND2_X1 U6867 ( .A1(n6095), .A2(REIP_REG_14__SCAN_IN), .ZN(n5820) );
  INV_X1 U6868 ( .A(n5808), .ZN(n5809) );
  AOI21_X1 U6869 ( .B1(n5810), .B2(n5809), .A(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5815) );
  INV_X1 U6870 ( .A(n5811), .ZN(n5812) );
  AOI21_X1 U6871 ( .B1(n5822), .B2(n5812), .A(n6115), .ZN(n5813) );
  OAI21_X1 U6872 ( .B1(n5817), .B2(n5814), .A(n5813), .ZN(n5827) );
  OAI21_X1 U6873 ( .B1(n5815), .B2(n5827), .A(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n5819) );
  NAND3_X1 U6874 ( .A1(n5817), .A2(n5569), .A3(n5816), .ZN(n5818) );
  NAND4_X1 U6875 ( .A1(n5821), .A2(n5820), .A3(n5819), .A4(n5818), .ZN(U3004)
         );
  OR2_X1 U6876 ( .A1(n5822), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5831)
         );
  INV_X1 U6877 ( .A(n5823), .ZN(n5824) );
  AOI21_X1 U6878 ( .B1(n5825), .B2(n6138), .A(n5824), .ZN(n5830) );
  INV_X1 U6879 ( .A(n5826), .ZN(n5828) );
  AOI22_X1 U6880 ( .A1(n5828), .A2(n6155), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5827), .ZN(n5829) );
  OAI211_X1 U6881 ( .C1(n6119), .C2(n5831), .A(n5830), .B(n5829), .ZN(U3005)
         );
  INV_X1 U6882 ( .A(n5832), .ZN(n5833) );
  NAND2_X1 U6883 ( .A1(n5833), .A2(n3238), .ZN(n5834) );
  OAI22_X1 U6884 ( .A1(n5835), .A2(n5834), .B1(n4723), .B2(n6645), .ZN(U3455)
         );
  INV_X1 U6885 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6565) );
  AOI21_X1 U6886 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6565), .A(n6559), .ZN(n5840) );
  INV_X1 U6887 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5836) );
  AOI21_X1 U6888 ( .B1(n5840), .B2(n5836), .A(n6613), .ZN(U2789) );
  OAI21_X1 U6889 ( .B1(n5837), .B2(n6537), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5838) );
  OAI21_X1 U6890 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6538), .A(n5838), .ZN(
        U2790) );
  NOR2_X1 U6891 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5841) );
  OAI21_X1 U6892 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5841), .A(n6668), .ZN(n5839)
         );
  OAI21_X1 U6893 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6657), .A(n5839), .ZN(
        U2791) );
  OAI21_X1 U6894 ( .B1(BS16_N), .B2(n5841), .A(n6629), .ZN(n6627) );
  OAI21_X1 U6895 ( .B1(n6629), .B2(n6432), .A(n6627), .ZN(U2792) );
  OAI21_X1 U6896 ( .B1(n5843), .B2(n5842), .A(n6100), .ZN(U2793) );
  INV_X1 U6897 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5846) );
  INV_X1 U6898 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6628) );
  NOR4_X1 U6899 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(DATAWIDTH_REG_3__SCAN_IN), 
        .A3(DATAWIDTH_REG_4__SCAN_IN), .A4(DATAWIDTH_REG_5__SCAN_IN), .ZN(
        n5844) );
  OAI211_X1 U6900 ( .C1(n5846), .C2(n6628), .A(n5845), .B(n5844), .ZN(n5854)
         );
  OR4_X1 U6901 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(DATAWIDTH_REG_11__SCAN_IN), .A3(DATAWIDTH_REG_12__SCAN_IN), .A4(DATAWIDTH_REG_13__SCAN_IN), .ZN(n5853)
         );
  OR4_X1 U6902 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), 
        .A3(DATAWIDTH_REG_8__SCAN_IN), .A4(DATAWIDTH_REG_9__SCAN_IN), .ZN(
        n5852) );
  NOR4_X1 U6903 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(
        DATAWIDTH_REG_19__SCAN_IN), .A3(DATAWIDTH_REG_20__SCAN_IN), .A4(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n5850) );
  NOR4_X1 U6904 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_14__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_17__SCAN_IN), .ZN(n5849) );
  NOR4_X1 U6905 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_29__SCAN_IN), .A4(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n5848) );
  NOR4_X1 U6906 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_23__SCAN_IN), .A3(DATAWIDTH_REG_25__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5847) );
  NAND4_X1 U6907 ( .A1(n5850), .A2(n5849), .A3(n5848), .A4(n5847), .ZN(n5851)
         );
  NOR4_X2 U6908 ( .A1(n5854), .A2(n5853), .A3(n5852), .A4(n5851), .ZN(n6655)
         );
  INV_X1 U6909 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5856) );
  NOR3_X1 U6910 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5857) );
  OAI21_X1 U6911 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5857), .A(n6655), .ZN(n5855)
         );
  OAI21_X1 U6912 ( .B1(n6655), .B2(n5856), .A(n5855), .ZN(U2794) );
  AOI21_X1 U6913 ( .B1(n5390), .B2(n6628), .A(n5857), .ZN(n5859) );
  INV_X1 U6914 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5858) );
  INV_X1 U6915 ( .A(n6655), .ZN(n6650) );
  AOI22_X1 U6916 ( .A1(n6655), .A2(n5859), .B1(n5858), .B2(n6650), .ZN(U2795)
         );
  AOI22_X1 U6917 ( .A1(EBX_REG_15__SCAN_IN), .A2(n5961), .B1(
        REIP_REG_15__SCAN_IN), .B2(n5860), .ZN(n5861) );
  OAI211_X1 U6918 ( .C1(n5908), .C2(n3040), .A(n5861), .B(n5918), .ZN(n5862)
         );
  AOI211_X1 U6919 ( .C1(n5864), .C2(n4228), .A(n5863), .B(n5862), .ZN(n5868)
         );
  AOI22_X1 U6920 ( .A1(n5866), .A2(n5948), .B1(n5927), .B2(n5865), .ZN(n5867)
         );
  NAND2_X1 U6921 ( .A1(n5868), .A2(n5867), .ZN(U2812) );
  AOI22_X1 U6922 ( .A1(PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n5960), .B1(n5927), 
        .B2(n5976), .ZN(n5876) );
  NOR2_X1 U6923 ( .A1(n5978), .A2(n5952), .ZN(n5869) );
  AOI211_X1 U6924 ( .C1(REIP_REG_12__SCAN_IN), .C2(n5871), .A(n5870), .B(n5869), .ZN(n5875) );
  INV_X1 U6925 ( .A(n5337), .ZN(n5872) );
  AOI21_X1 U6926 ( .B1(n5873), .B2(n5040), .A(n5872), .ZN(n6097) );
  AOI22_X1 U6927 ( .A1(n6097), .A2(n4228), .B1(n5948), .B2(n6096), .ZN(n5874)
         );
  NAND4_X1 U6928 ( .A1(n5876), .A2(n5875), .A3(n5874), .A4(n5918), .ZN(U2815)
         );
  AOI22_X1 U6929 ( .A1(EBX_REG_10__SCAN_IN), .A2(n5961), .B1(n5927), .B2(n5877), .ZN(n5886) );
  NOR3_X1 U6930 ( .A1(REIP_REG_10__SCAN_IN), .A2(n5878), .A3(n5907), .ZN(n5879) );
  AOI211_X1 U6931 ( .C1(n5960), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n5933), 
        .B(n5879), .ZN(n5885) );
  AOI22_X1 U6932 ( .A1(n5881), .A2(n4228), .B1(n5948), .B2(n5880), .ZN(n5884)
         );
  OAI21_X1 U6933 ( .B1(n5882), .B2(n5890), .A(REIP_REG_10__SCAN_IN), .ZN(n5883) );
  NAND4_X1 U6934 ( .A1(n5886), .A2(n5885), .A3(n5884), .A4(n5883), .ZN(U2817)
         );
  AOI22_X1 U6935 ( .A1(EBX_REG_8__SCAN_IN), .A2(n5961), .B1(
        PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n5960), .ZN(n5895) );
  AOI21_X1 U6936 ( .B1(n5927), .B2(n5887), .A(n5933), .ZN(n5894) );
  AOI22_X1 U6937 ( .A1(n5889), .A2(n4228), .B1(n5948), .B2(n5888), .ZN(n5893)
         );
  OAI21_X1 U6938 ( .B1(REIP_REG_8__SCAN_IN), .B2(n5891), .A(n5890), .ZN(n5892)
         );
  NAND4_X1 U6939 ( .A1(n5895), .A2(n5894), .A3(n5893), .A4(n5892), .ZN(U2819)
         );
  AOI22_X1 U6940 ( .A1(EBX_REG_7__SCAN_IN), .A2(n5961), .B1(
        PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n5960), .ZN(n5896) );
  OAI211_X1 U6941 ( .C1(n5968), .C2(n5897), .A(n5896), .B(n5918), .ZN(n5902)
         );
  OAI22_X1 U6942 ( .A1(n5900), .A2(n5899), .B1(n5898), .B2(n5965), .ZN(n5901)
         );
  NOR2_X1 U6943 ( .A1(n5902), .A2(n5901), .ZN(n5906) );
  OAI211_X1 U6944 ( .C1(REIP_REG_7__SCAN_IN), .C2(REIP_REG_6__SCAN_IN), .A(
        n5904), .B(n5903), .ZN(n5905) );
  OAI211_X1 U6945 ( .C1(n5916), .C2(n6578), .A(n5906), .B(n5905), .ZN(U2820)
         );
  OAI22_X1 U6946 ( .A1(n5907), .A2(REIP_REG_6__SCAN_IN), .B1(n5916), .B2(n6576), .ZN(n5912) );
  OAI22_X1 U6947 ( .A1(n4022), .A2(n5952), .B1(n3049), .B2(n5908), .ZN(n5909)
         );
  AOI211_X1 U6948 ( .C1(n5927), .C2(n3108), .A(n5933), .B(n5909), .ZN(n5910)
         );
  INV_X1 U6949 ( .A(n5910), .ZN(n5911) );
  AOI211_X1 U6950 ( .C1(n4228), .C2(n6103), .A(n5912), .B(n5911), .ZN(n5913)
         );
  OAI21_X1 U6951 ( .B1(n5914), .B2(n5965), .A(n5913), .ZN(U2821) );
  NAND2_X1 U6952 ( .A1(n5939), .A2(n5915), .ZN(n5917) );
  AOI21_X1 U6953 ( .B1(n6574), .B2(n5917), .A(n5916), .ZN(n5922) );
  AOI22_X1 U6954 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n5960), .B1(n5927), 
        .B2(n6139), .ZN(n5919) );
  OAI211_X1 U6955 ( .C1(n5952), .C2(n5920), .A(n5919), .B(n5918), .ZN(n5921)
         );
  AOI211_X1 U6956 ( .C1(n5923), .C2(n5971), .A(n5922), .B(n5921), .ZN(n5924)
         );
  OAI21_X1 U6957 ( .B1(n5925), .B2(n5965), .A(n5924), .ZN(U2822) );
  AOI22_X1 U6958 ( .A1(EBX_REG_4__SCAN_IN), .A2(n5961), .B1(n5927), .B2(n5926), 
        .ZN(n5943) );
  OAI21_X1 U6959 ( .B1(n5929), .B2(n5937), .A(n5928), .ZN(n5959) );
  INV_X1 U6960 ( .A(n5930), .ZN(n5931) );
  OAI22_X1 U6961 ( .A1(n5959), .A2(n6572), .B1(n5931), .B2(n5964), .ZN(n5932)
         );
  AOI211_X1 U6962 ( .C1(n5960), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n5933), 
        .B(n5932), .ZN(n5942) );
  INV_X1 U6963 ( .A(n5934), .ZN(n5935) );
  AOI22_X1 U6964 ( .A1(n5936), .A2(n5971), .B1(n5935), .B2(n5948), .ZN(n5941)
         );
  INV_X1 U6965 ( .A(n5937), .ZN(n5938) );
  NAND3_X1 U6966 ( .A1(n5939), .A2(n6572), .A3(n5938), .ZN(n5940) );
  NAND4_X1 U6967 ( .A1(n5943), .A2(n5942), .A3(n5941), .A4(n5940), .ZN(U2823)
         );
  INV_X1 U6968 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6570) );
  OR2_X1 U6969 ( .A1(n5944), .A2(n6568), .ZN(n5958) );
  INV_X1 U6970 ( .A(n5945), .ZN(n5956) );
  INV_X1 U6971 ( .A(n5946), .ZN(n5947) );
  AOI22_X1 U6972 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n5960), .B1(n5948), 
        .B2(n5947), .ZN(n5949) );
  OAI21_X1 U6973 ( .B1(n5950), .B2(n5964), .A(n5949), .ZN(n5955) );
  OAI22_X1 U6974 ( .A1(n5953), .A2(n5952), .B1(n5968), .B2(n5951), .ZN(n5954)
         );
  AOI211_X1 U6975 ( .C1(n5956), .C2(n5971), .A(n5955), .B(n5954), .ZN(n5957)
         );
  OAI221_X1 U6976 ( .B1(n5959), .B2(n6570), .C1(n5959), .C2(n5958), .A(n5957), 
        .ZN(U2824) );
  AOI22_X1 U6977 ( .A1(EBX_REG_1__SCAN_IN), .A2(n5961), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n5960), .ZN(n5974) );
  INV_X1 U6978 ( .A(n5962), .ZN(n5972) );
  OAI22_X1 U6979 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n5965), .B1(n5964), 
        .B2(n5963), .ZN(n5970) );
  INV_X1 U6980 ( .A(n4575), .ZN(n5967) );
  OAI21_X1 U6981 ( .B1(n5968), .B2(n5967), .A(n5966), .ZN(n5969) );
  AOI211_X1 U6982 ( .C1(n5972), .C2(n5971), .A(n5970), .B(n5969), .ZN(n5973)
         );
  OAI211_X1 U6983 ( .C1(n5975), .C2(n5390), .A(n5974), .B(n5973), .ZN(U2826)
         );
  AOI22_X1 U6984 ( .A1(n6097), .A2(n5980), .B1(n5979), .B2(n5976), .ZN(n5977)
         );
  OAI21_X1 U6985 ( .B1(n5987), .B2(n5978), .A(n5977), .ZN(U2847) );
  AOI22_X1 U6986 ( .A1(n6103), .A2(n5980), .B1(n5979), .B2(n3108), .ZN(n5981)
         );
  OAI21_X1 U6987 ( .B1(n5987), .B2(n4022), .A(n5981), .ZN(U2853) );
  OAI22_X1 U6988 ( .A1(n5983), .A2(n5438), .B1(n5433), .B2(n5982), .ZN(n5984)
         );
  INV_X1 U6989 ( .A(n5984), .ZN(n5985) );
  OAI21_X1 U6990 ( .B1(n5987), .B2(n5986), .A(n5985), .ZN(U2857) );
  AOI22_X1 U6991 ( .A1(n6097), .A2(n5989), .B1(DATAI_12_), .B2(n5988), .ZN(
        n5990) );
  OAI21_X1 U6992 ( .B1(n6081), .B2(n5991), .A(n5990), .ZN(U2879) );
  INV_X1 U6993 ( .A(n6033), .ZN(n6018) );
  AOI22_X1 U6994 ( .A1(n6001), .A2(EAX_REG_30__SCAN_IN), .B1(n6016), .B2(
        UWORD_REG_14__SCAN_IN), .ZN(n5993) );
  OAI21_X1 U6995 ( .B1(n5994), .B2(n6018), .A(n5993), .ZN(U2893) );
  AOI22_X1 U6996 ( .A1(n6033), .A2(DATAO_REG_24__SCAN_IN), .B1(n6001), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5995) );
  OAI21_X1 U6997 ( .B1(n5996), .B2(n6523), .A(n5995), .ZN(U2899) );
  AOI22_X1 U6998 ( .A1(n6001), .A2(EAX_REG_22__SCAN_IN), .B1(n6016), .B2(
        UWORD_REG_6__SCAN_IN), .ZN(n5997) );
  OAI21_X1 U6999 ( .B1(n5998), .B2(n6018), .A(n5997), .ZN(U2901) );
  AOI22_X1 U7000 ( .A1(n6001), .A2(EAX_REG_19__SCAN_IN), .B1(n6016), .B2(
        UWORD_REG_3__SCAN_IN), .ZN(n5999) );
  OAI21_X1 U7001 ( .B1(n6000), .B2(n6018), .A(n5999), .ZN(U2904) );
  AOI22_X1 U7002 ( .A1(n6001), .A2(EAX_REG_18__SCAN_IN), .B1(n6016), .B2(
        UWORD_REG_2__SCAN_IN), .ZN(n6002) );
  OAI21_X1 U7003 ( .B1(n6003), .B2(n6018), .A(n6002), .ZN(U2905) );
  INV_X1 U7004 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6093) );
  AOI22_X1 U7005 ( .A1(n6016), .A2(LWORD_REG_15__SCAN_IN), .B1(n6033), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6004) );
  OAI21_X1 U7006 ( .B1(n6093), .B2(n6035), .A(n6004), .ZN(U2908) );
  AOI22_X1 U7007 ( .A1(EAX_REG_14__SCAN_IN), .A2(n6022), .B1(n6033), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6005) );
  OAI21_X1 U7008 ( .B1(n6006), .B2(n6523), .A(n6005), .ZN(U2909) );
  AOI22_X1 U7009 ( .A1(LWORD_REG_13__SCAN_IN), .A2(n6016), .B1(n6033), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6007) );
  OAI21_X1 U7010 ( .B1(n6008), .B2(n6035), .A(n6007), .ZN(U2910) );
  AOI22_X1 U7011 ( .A1(n6016), .A2(LWORD_REG_12__SCAN_IN), .B1(n6033), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6009) );
  OAI21_X1 U7012 ( .B1(n6081), .B2(n6035), .A(n6009), .ZN(U2911) );
  INV_X1 U7013 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6011) );
  AOI22_X1 U7014 ( .A1(n6016), .A2(LWORD_REG_11__SCAN_IN), .B1(n6033), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6010) );
  OAI21_X1 U7015 ( .B1(n6011), .B2(n6035), .A(n6010), .ZN(U2912) );
  INV_X1 U7016 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6013) );
  AOI22_X1 U7017 ( .A1(n6016), .A2(LWORD_REG_10__SCAN_IN), .B1(n6033), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6012) );
  OAI21_X1 U7018 ( .B1(n6013), .B2(n6035), .A(n6012), .ZN(U2913) );
  INV_X1 U7019 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6015) );
  AOI22_X1 U7020 ( .A1(n6016), .A2(LWORD_REG_9__SCAN_IN), .B1(n6033), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6014) );
  OAI21_X1 U7021 ( .B1(n6015), .B2(n6035), .A(n6014), .ZN(U2914) );
  AOI22_X1 U7022 ( .A1(EAX_REG_8__SCAN_IN), .A2(n6022), .B1(n6016), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n6017) );
  OAI21_X1 U7023 ( .B1(n6019), .B2(n6018), .A(n6017), .ZN(U2915) );
  AOI22_X1 U7024 ( .A1(EAX_REG_7__SCAN_IN), .A2(n6022), .B1(n6033), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6020) );
  OAI21_X1 U7025 ( .B1(n6021), .B2(n6523), .A(n6020), .ZN(U2916) );
  AOI222_X1 U7026 ( .A1(LWORD_REG_6__SCAN_IN), .A2(n6016), .B1(n6022), .B2(
        EAX_REG_6__SCAN_IN), .C1(n6033), .C2(DATAO_REG_6__SCAN_IN), .ZN(n6023)
         );
  INV_X1 U7027 ( .A(n6023), .ZN(U2917) );
  AOI22_X1 U7028 ( .A1(n6016), .A2(LWORD_REG_5__SCAN_IN), .B1(n6033), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6024) );
  OAI21_X1 U7029 ( .B1(n3454), .B2(n6035), .A(n6024), .ZN(U2918) );
  AOI22_X1 U7030 ( .A1(n6016), .A2(LWORD_REG_4__SCAN_IN), .B1(n6033), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6025) );
  OAI21_X1 U7031 ( .B1(n6026), .B2(n6035), .A(n6025), .ZN(U2919) );
  AOI22_X1 U7032 ( .A1(n6016), .A2(LWORD_REG_3__SCAN_IN), .B1(n6033), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6027) );
  OAI21_X1 U7033 ( .B1(n6028), .B2(n6035), .A(n6027), .ZN(U2920) );
  AOI22_X1 U7034 ( .A1(n6016), .A2(LWORD_REG_2__SCAN_IN), .B1(n6033), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6029) );
  OAI21_X1 U7035 ( .B1(n6030), .B2(n6035), .A(n6029), .ZN(U2921) );
  AOI22_X1 U7036 ( .A1(n6016), .A2(LWORD_REG_1__SCAN_IN), .B1(n6033), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6031) );
  OAI21_X1 U7037 ( .B1(n6032), .B2(n6035), .A(n6031), .ZN(U2922) );
  AOI22_X1 U7038 ( .A1(n6016), .A2(LWORD_REG_0__SCAN_IN), .B1(n6033), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6034) );
  OAI21_X1 U7039 ( .B1(n6036), .B2(n6035), .A(n6034), .ZN(U2923) );
  AOI22_X1 U7040 ( .A1(n6090), .A2(DATAI_0_), .B1(n6086), .B2(
        UWORD_REG_0__SCAN_IN), .ZN(n6038) );
  OAI21_X1 U7041 ( .B1(n6039), .B2(n6092), .A(n6038), .ZN(U2924) );
  AOI22_X1 U7042 ( .A1(n6090), .A2(DATAI_1_), .B1(n6089), .B2(
        UWORD_REG_1__SCAN_IN), .ZN(n6040) );
  OAI21_X1 U7043 ( .B1(n6041), .B2(n6092), .A(n6040), .ZN(U2925) );
  INV_X1 U7044 ( .A(DATAI_2_), .ZN(n6060) );
  AOI22_X1 U7045 ( .A1(n6086), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n6085), .ZN(n6042) );
  OAI21_X1 U7046 ( .B1(n6083), .B2(n6060), .A(n6042), .ZN(U2926) );
  AOI22_X1 U7047 ( .A1(n6089), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n6085), .ZN(n6043) );
  OAI21_X1 U7048 ( .B1(n6083), .B2(n6062), .A(n6043), .ZN(U2927) );
  AOI22_X1 U7049 ( .A1(n6086), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n6085), .ZN(n6044) );
  OAI21_X1 U7050 ( .B1(n6083), .B2(n6064), .A(n6044), .ZN(U2928) );
  AOI22_X1 U7051 ( .A1(n6089), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n6085), .ZN(n6045) );
  OAI21_X1 U7052 ( .B1(n6083), .B2(n6066), .A(n6045), .ZN(U2929) );
  AOI22_X1 U7053 ( .A1(n6086), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n6085), .ZN(n6046) );
  OAI21_X1 U7054 ( .B1(n6068), .B2(n6083), .A(n6046), .ZN(U2930) );
  AOI22_X1 U7055 ( .A1(n6086), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n6085), .ZN(n6047) );
  OAI21_X1 U7056 ( .B1(n6070), .B2(n6083), .A(n6047), .ZN(U2931) );
  AOI22_X1 U7057 ( .A1(n6090), .A2(DATAI_9_), .B1(n6089), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n6048) );
  OAI21_X1 U7058 ( .B1(n6049), .B2(n6092), .A(n6048), .ZN(U2933) );
  AOI22_X1 U7059 ( .A1(n6090), .A2(DATAI_10_), .B1(n6089), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n6050) );
  OAI21_X1 U7060 ( .B1(n3804), .B2(n6092), .A(n6050), .ZN(U2934) );
  INV_X1 U7061 ( .A(DATAI_12_), .ZN(n6051) );
  NOR2_X1 U7062 ( .A1(n6083), .A2(n6051), .ZN(n6079) );
  AOI21_X1 U7063 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n6086), .A(n6079), .ZN(
        n6052) );
  OAI21_X1 U7064 ( .B1(n3850), .B2(n6092), .A(n6052), .ZN(U2936) );
  AOI22_X1 U7065 ( .A1(n6086), .A2(UWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_29__SCAN_IN), .B2(n6085), .ZN(n6053) );
  OAI21_X1 U7066 ( .B1(n6084), .B2(n6083), .A(n6053), .ZN(U2937) );
  AOI22_X1 U7067 ( .A1(n6086), .A2(UWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_30__SCAN_IN), .B2(n6085), .ZN(n6054) );
  NAND2_X1 U7068 ( .A1(n6090), .A2(DATAI_14_), .ZN(n6087) );
  NAND2_X1 U7069 ( .A1(n6054), .A2(n6087), .ZN(U2938) );
  AOI22_X1 U7070 ( .A1(n6086), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n6085), .ZN(n6055) );
  OAI21_X1 U7071 ( .B1(n6083), .B2(n6056), .A(n6055), .ZN(U2939) );
  AOI22_X1 U7072 ( .A1(n6086), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n6085), .ZN(n6057) );
  OAI21_X1 U7073 ( .B1(n6083), .B2(n6058), .A(n6057), .ZN(U2940) );
  AOI22_X1 U7074 ( .A1(n6086), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n6085), .ZN(n6059) );
  OAI21_X1 U7075 ( .B1(n6083), .B2(n6060), .A(n6059), .ZN(U2941) );
  AOI22_X1 U7076 ( .A1(n6086), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n6085), .ZN(n6061) );
  OAI21_X1 U7077 ( .B1(n6083), .B2(n6062), .A(n6061), .ZN(U2942) );
  AOI22_X1 U7078 ( .A1(n6086), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n6085), .ZN(n6063) );
  OAI21_X1 U7079 ( .B1(n6083), .B2(n6064), .A(n6063), .ZN(U2943) );
  AOI22_X1 U7080 ( .A1(n6086), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n6085), .ZN(n6065) );
  OAI21_X1 U7081 ( .B1(n6083), .B2(n6066), .A(n6065), .ZN(U2944) );
  AOI22_X1 U7082 ( .A1(n6086), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n6085), .ZN(n6067) );
  OAI21_X1 U7083 ( .B1(n6068), .B2(n6083), .A(n6067), .ZN(U2945) );
  AOI22_X1 U7084 ( .A1(n6086), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n6085), .ZN(n6069) );
  OAI21_X1 U7085 ( .B1(n6070), .B2(n6083), .A(n6069), .ZN(U2946) );
  AOI22_X1 U7086 ( .A1(n6086), .A2(LWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_8__SCAN_IN), .B2(n6085), .ZN(n6072) );
  NAND2_X1 U7087 ( .A1(n6090), .A2(DATAI_8_), .ZN(n6071) );
  NAND2_X1 U7088 ( .A1(n6072), .A2(n6071), .ZN(U2947) );
  AOI22_X1 U7089 ( .A1(n6086), .A2(LWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_9__SCAN_IN), .B2(n6085), .ZN(n6074) );
  NAND2_X1 U7090 ( .A1(n6090), .A2(DATAI_9_), .ZN(n6073) );
  NAND2_X1 U7091 ( .A1(n6074), .A2(n6073), .ZN(U2948) );
  AOI22_X1 U7092 ( .A1(n6086), .A2(LWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_10__SCAN_IN), .B2(n6085), .ZN(n6076) );
  NAND2_X1 U7093 ( .A1(n6090), .A2(DATAI_10_), .ZN(n6075) );
  NAND2_X1 U7094 ( .A1(n6076), .A2(n6075), .ZN(U2949) );
  AOI22_X1 U7095 ( .A1(n6086), .A2(LWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_11__SCAN_IN), .B2(n6085), .ZN(n6078) );
  NAND2_X1 U7096 ( .A1(n6090), .A2(DATAI_11_), .ZN(n6077) );
  NAND2_X1 U7097 ( .A1(n6078), .A2(n6077), .ZN(U2950) );
  AOI21_X1 U7098 ( .B1(LWORD_REG_12__SCAN_IN), .B2(n6086), .A(n6079), .ZN(
        n6080) );
  OAI21_X1 U7099 ( .B1(n6081), .B2(n6092), .A(n6080), .ZN(U2951) );
  AOI22_X1 U7100 ( .A1(n6086), .A2(LWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_13__SCAN_IN), .B2(n6085), .ZN(n6082) );
  OAI21_X1 U7101 ( .B1(n6084), .B2(n6083), .A(n6082), .ZN(U2952) );
  AOI22_X1 U7102 ( .A1(n6086), .A2(LWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_14__SCAN_IN), .B2(n6085), .ZN(n6088) );
  NAND2_X1 U7103 ( .A1(n6088), .A2(n6087), .ZN(U2953) );
  AOI22_X1 U7104 ( .A1(n6090), .A2(DATAI_15_), .B1(n6089), .B2(
        LWORD_REG_15__SCAN_IN), .ZN(n6091) );
  OAI21_X1 U7105 ( .B1(n6093), .B2(n6092), .A(n6091), .ZN(U2954) );
  AOI22_X1 U7106 ( .A1(n6095), .A2(REIP_REG_12__SCAN_IN), .B1(n6094), .B2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n6099) );
  AOI22_X1 U7107 ( .A1(n6097), .A2(n6104), .B1(n6105), .B2(n6096), .ZN(n6098)
         );
  OAI211_X1 U7108 ( .C1(n6101), .C2(n6100), .A(n6099), .B(n6098), .ZN(U2974)
         );
  INV_X1 U7109 ( .A(n6102), .ZN(n6108) );
  AOI222_X1 U7110 ( .A1(n6108), .A2(n6107), .B1(n6106), .B2(n6105), .C1(n6104), 
        .C2(n6103), .ZN(n6111) );
  INV_X1 U7111 ( .A(n6109), .ZN(n6110) );
  OAI211_X1 U7112 ( .C1(n3049), .C2(n6112), .A(n6111), .B(n6110), .ZN(U2980)
         );
  AOI21_X1 U7113 ( .B1(n6114), .B2(n6138), .A(n6113), .ZN(n6118) );
  AOI22_X1 U7114 ( .A1(n6116), .A2(n6155), .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6115), .ZN(n6117) );
  OAI211_X1 U7115 ( .C1(INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n6119), .A(n6118), .B(n6117), .ZN(U3007) );
  OAI21_X1 U7116 ( .B1(INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .A(n6120), .ZN(n6129) );
  INV_X1 U7117 ( .A(n6121), .ZN(n6127) );
  OAI22_X1 U7118 ( .A1(n6123), .A2(n6149), .B1(n6580), .B2(n6122), .ZN(n6126)
         );
  NOR2_X1 U7119 ( .A1(n6124), .A2(n6142), .ZN(n6125) );
  AOI211_X1 U7120 ( .C1(INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n6127), .A(n6126), 
        .B(n6125), .ZN(n6128) );
  OAI21_X1 U7121 ( .B1(n6130), .B2(n6129), .A(n6128), .ZN(U3010) );
  NAND2_X1 U7122 ( .A1(n6132), .A2(n6131), .ZN(n6146) );
  AOI21_X1 U7123 ( .B1(n6133), .B2(n6132), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n6134) );
  INV_X1 U7124 ( .A(n6134), .ZN(n6135) );
  NAND2_X1 U7125 ( .A1(n6136), .A2(n6135), .ZN(n6141) );
  AOI21_X1 U7126 ( .B1(n6139), .B2(n6138), .A(n6137), .ZN(n6140) );
  OAI211_X1 U7127 ( .C1(n6143), .C2(n6142), .A(n6141), .B(n6140), .ZN(n6144)
         );
  INV_X1 U7128 ( .A(n6144), .ZN(n6145) );
  OAI21_X1 U7129 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n6146), .A(n6145), 
        .ZN(U3013) );
  OAI21_X1 U7130 ( .B1(n6149), .B2(n6148), .A(n6147), .ZN(n6150) );
  INV_X1 U7131 ( .A(n6150), .ZN(n6158) );
  INV_X1 U7132 ( .A(n6151), .ZN(n6152) );
  NOR3_X1 U7133 ( .A1(n6153), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n6152), 
        .ZN(n6154) );
  AOI21_X1 U7134 ( .B1(n6156), .B2(n6155), .A(n6154), .ZN(n6157) );
  OAI211_X1 U7135 ( .C1(n6160), .C2(n6159), .A(n6158), .B(n6157), .ZN(U3017)
         );
  NOR2_X1 U7136 ( .A1(n6162), .A2(n6161), .ZN(U3019) );
  INV_X1 U7137 ( .A(n6163), .ZN(n6171) );
  AOI22_X1 U7138 ( .A1(n6464), .A2(n6165), .B1(n6164), .B2(n6405), .ZN(n6169)
         );
  AOI22_X1 U7139 ( .A1(n6167), .A2(n6465), .B1(n6466), .B2(n6166), .ZN(n6168)
         );
  OAI211_X1 U7140 ( .C1(n6171), .C2(n6170), .A(n6169), .B(n6168), .ZN(U3032)
         );
  OAI21_X1 U7141 ( .B1(n6381), .B2(n6172), .A(n6380), .ZN(n6173) );
  NAND2_X1 U7142 ( .A1(n6174), .A2(n6173), .ZN(n6179) );
  NAND2_X1 U7143 ( .A1(n6275), .A2(n6175), .ZN(n6177) );
  NOR2_X1 U7144 ( .A1(n6378), .A2(n6180), .ZN(n6200) );
  INV_X1 U7145 ( .A(n6200), .ZN(n6176) );
  NAND2_X1 U7146 ( .A1(n6177), .A2(n6176), .ZN(n6182) );
  INV_X1 U7147 ( .A(n6180), .ZN(n6178) );
  AOI22_X1 U7148 ( .A1(n6430), .A2(n6200), .B1(n6199), .B2(n6379), .ZN(n6186)
         );
  INV_X1 U7149 ( .A(n6179), .ZN(n6183) );
  AOI21_X1 U7150 ( .B1(n6435), .B2(n6180), .A(n6384), .ZN(n6181) );
  AOI22_X1 U7151 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6201), .B1(n6442), 
        .B2(n6209), .ZN(n6185) );
  OAI211_X1 U7152 ( .C1(n6204), .C2(n6348), .A(n6186), .B(n6185), .ZN(U3044)
         );
  AOI22_X1 U7153 ( .A1(n6446), .A2(n6200), .B1(n6393), .B2(n6199), .ZN(n6188)
         );
  AOI22_X1 U7154 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6201), .B1(n6448), 
        .B2(n6209), .ZN(n6187) );
  OAI211_X1 U7155 ( .C1(n6204), .C2(n6351), .A(n6188), .B(n6187), .ZN(U3045)
         );
  AOI22_X1 U7156 ( .A1(n6452), .A2(n6200), .B1(n6352), .B2(n6199), .ZN(n6190)
         );
  AOI22_X1 U7157 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6201), .B1(n6454), 
        .B2(n6209), .ZN(n6189) );
  OAI211_X1 U7158 ( .C1(n6204), .C2(n6355), .A(n6190), .B(n6189), .ZN(U3046)
         );
  AOI22_X1 U7159 ( .A1(n6458), .A2(n6200), .B1(n6401), .B2(n6199), .ZN(n6192)
         );
  AOI22_X1 U7160 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6201), .B1(n6460), 
        .B2(n6209), .ZN(n6191) );
  OAI211_X1 U7161 ( .C1(n6204), .C2(n6358), .A(n6192), .B(n6191), .ZN(U3047)
         );
  AOI22_X1 U7162 ( .A1(n6464), .A2(n6200), .B1(n6405), .B2(n6199), .ZN(n6194)
         );
  AOI22_X1 U7163 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6201), .B1(n6466), 
        .B2(n6209), .ZN(n6193) );
  OAI211_X1 U7164 ( .C1(n6204), .C2(n6361), .A(n6194), .B(n6193), .ZN(U3048)
         );
  AOI22_X1 U7165 ( .A1(n6470), .A2(n6200), .B1(n6409), .B2(n6199), .ZN(n6196)
         );
  AOI22_X1 U7166 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6201), .B1(n6472), 
        .B2(n6209), .ZN(n6195) );
  OAI211_X1 U7167 ( .C1(n6204), .C2(n6364), .A(n6196), .B(n6195), .ZN(U3049)
         );
  AOI22_X1 U7168 ( .A1(n6476), .A2(n6200), .B1(n6413), .B2(n6199), .ZN(n6198)
         );
  AOI22_X1 U7169 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6201), .B1(n6478), 
        .B2(n6209), .ZN(n6197) );
  OAI211_X1 U7170 ( .C1(n6204), .C2(n6367), .A(n6198), .B(n6197), .ZN(U3050)
         );
  AOI22_X1 U7171 ( .A1(n6483), .A2(n6200), .B1(n6419), .B2(n6199), .ZN(n6203)
         );
  AOI22_X1 U7172 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6201), .B1(n6487), 
        .B2(n6209), .ZN(n6202) );
  OAI211_X1 U7173 ( .C1(n6204), .C2(n6374), .A(n6203), .B(n6202), .ZN(U3051)
         );
  INV_X1 U7174 ( .A(n6437), .ZN(n6427) );
  OAI22_X1 U7175 ( .A1(n6313), .A2(n6427), .B1(n6426), .B2(n6205), .ZN(n6229)
         );
  NAND2_X1 U7176 ( .A1(n6206), .A2(n6509), .ZN(n6236) );
  NOR2_X1 U7177 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6236), .ZN(n6228)
         );
  AOI22_X1 U7178 ( .A1(n6431), .A2(n6229), .B1(n6430), .B2(n6228), .ZN(n6215)
         );
  OAI21_X1 U7179 ( .B1(n6213), .B2(n6432), .A(n6380), .ZN(n6234) );
  AOI211_X1 U7180 ( .C1(n6209), .C2(n6208), .A(n6235), .B(n6234), .ZN(n6212)
         );
  OAI211_X1 U7181 ( .C1(n3238), .C2(n6228), .A(n6439), .B(n6210), .ZN(n6211)
         );
  NOR2_X2 U7182 ( .A1(n6213), .A2(n6307), .ZN(n6258) );
  AOI22_X1 U7183 ( .A1(n6230), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n6442), 
        .B2(n6258), .ZN(n6214) );
  OAI211_X1 U7184 ( .C1(n6445), .C2(n6233), .A(n6215), .B(n6214), .ZN(U3052)
         );
  AOI22_X1 U7185 ( .A1(n6447), .A2(n6229), .B1(n6446), .B2(n6228), .ZN(n6217)
         );
  AOI22_X1 U7186 ( .A1(n6230), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n6448), 
        .B2(n6258), .ZN(n6216) );
  OAI211_X1 U7187 ( .C1(n6451), .C2(n6233), .A(n6217), .B(n6216), .ZN(U3053)
         );
  AOI22_X1 U7188 ( .A1(n6453), .A2(n6229), .B1(n6452), .B2(n6228), .ZN(n6219)
         );
  AOI22_X1 U7189 ( .A1(n6230), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n6454), 
        .B2(n6258), .ZN(n6218) );
  OAI211_X1 U7190 ( .C1(n6457), .C2(n6233), .A(n6219), .B(n6218), .ZN(U3054)
         );
  AOI22_X1 U7191 ( .A1(n6459), .A2(n6229), .B1(n6458), .B2(n6228), .ZN(n6221)
         );
  AOI22_X1 U7192 ( .A1(n6230), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n6460), 
        .B2(n6258), .ZN(n6220) );
  OAI211_X1 U7193 ( .C1(n6463), .C2(n6233), .A(n6221), .B(n6220), .ZN(U3055)
         );
  AOI22_X1 U7194 ( .A1(n6465), .A2(n6229), .B1(n6464), .B2(n6228), .ZN(n6223)
         );
  AOI22_X1 U7195 ( .A1(n6230), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n6466), 
        .B2(n6258), .ZN(n6222) );
  OAI211_X1 U7196 ( .C1(n6469), .C2(n6233), .A(n6223), .B(n6222), .ZN(U3056)
         );
  AOI22_X1 U7197 ( .A1(n6471), .A2(n6229), .B1(n6470), .B2(n6228), .ZN(n6225)
         );
  AOI22_X1 U7198 ( .A1(n6230), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n6472), 
        .B2(n6258), .ZN(n6224) );
  OAI211_X1 U7199 ( .C1(n6475), .C2(n6233), .A(n6225), .B(n6224), .ZN(U3057)
         );
  AOI22_X1 U7200 ( .A1(n6477), .A2(n6229), .B1(n6476), .B2(n6228), .ZN(n6227)
         );
  AOI22_X1 U7201 ( .A1(n6230), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n6478), 
        .B2(n6258), .ZN(n6226) );
  OAI211_X1 U7202 ( .C1(n6481), .C2(n6233), .A(n6227), .B(n6226), .ZN(U3058)
         );
  AOI22_X1 U7203 ( .A1(n6485), .A2(n6229), .B1(n6483), .B2(n6228), .ZN(n6232)
         );
  AOI22_X1 U7204 ( .A1(n6230), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n6487), 
        .B2(n6258), .ZN(n6231) );
  OAI211_X1 U7205 ( .C1(n6492), .C2(n6233), .A(n6232), .B(n6231), .ZN(U3059)
         );
  INV_X1 U7206 ( .A(n6234), .ZN(n6239) );
  NOR2_X1 U7207 ( .A1(n6378), .A2(n6236), .ZN(n6257) );
  AOI21_X1 U7208 ( .B1(n6235), .B2(n6495), .A(n6257), .ZN(n6238) );
  INV_X1 U7209 ( .A(n6238), .ZN(n6237) );
  INV_X1 U7210 ( .A(n6236), .ZN(n6242) );
  AOI22_X1 U7211 ( .A1(n6430), .A2(n6257), .B1(n6266), .B2(n6442), .ZN(n6244)
         );
  NAND2_X1 U7212 ( .A1(n6239), .A2(n6238), .ZN(n6241) );
  OAI211_X1 U7213 ( .C1(n6380), .C2(n6242), .A(n6241), .B(n6240), .ZN(n6259)
         );
  AOI22_X1 U7214 ( .A1(n6259), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n6379), 
        .B2(n6258), .ZN(n6243) );
  OAI211_X1 U7215 ( .C1(n6262), .C2(n6348), .A(n6244), .B(n6243), .ZN(U3060)
         );
  AOI22_X1 U7216 ( .A1(n6446), .A2(n6257), .B1(n6266), .B2(n6448), .ZN(n6246)
         );
  AOI22_X1 U7217 ( .A1(n6259), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n6393), 
        .B2(n6258), .ZN(n6245) );
  OAI211_X1 U7218 ( .C1(n6262), .C2(n6351), .A(n6246), .B(n6245), .ZN(U3061)
         );
  AOI22_X1 U7219 ( .A1(n6452), .A2(n6257), .B1(n6266), .B2(n6454), .ZN(n6248)
         );
  AOI22_X1 U7220 ( .A1(n6259), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n6352), 
        .B2(n6258), .ZN(n6247) );
  OAI211_X1 U7221 ( .C1(n6262), .C2(n6355), .A(n6248), .B(n6247), .ZN(U3062)
         );
  AOI22_X1 U7222 ( .A1(n6458), .A2(n6257), .B1(n6266), .B2(n6460), .ZN(n6250)
         );
  AOI22_X1 U7223 ( .A1(n6259), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n6401), 
        .B2(n6258), .ZN(n6249) );
  OAI211_X1 U7224 ( .C1(n6262), .C2(n6358), .A(n6250), .B(n6249), .ZN(U3063)
         );
  AOI22_X1 U7225 ( .A1(n6464), .A2(n6257), .B1(n6266), .B2(n6466), .ZN(n6252)
         );
  AOI22_X1 U7226 ( .A1(n6259), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n6405), 
        .B2(n6258), .ZN(n6251) );
  OAI211_X1 U7227 ( .C1(n6262), .C2(n6361), .A(n6252), .B(n6251), .ZN(U3064)
         );
  AOI22_X1 U7228 ( .A1(n6470), .A2(n6257), .B1(n6266), .B2(n6472), .ZN(n6254)
         );
  AOI22_X1 U7229 ( .A1(n6259), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n6409), 
        .B2(n6258), .ZN(n6253) );
  OAI211_X1 U7230 ( .C1(n6262), .C2(n6364), .A(n6254), .B(n6253), .ZN(U3065)
         );
  AOI22_X1 U7231 ( .A1(n6476), .A2(n6257), .B1(n6266), .B2(n6478), .ZN(n6256)
         );
  AOI22_X1 U7232 ( .A1(n6259), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n6413), 
        .B2(n6258), .ZN(n6255) );
  OAI211_X1 U7233 ( .C1(n6262), .C2(n6367), .A(n6256), .B(n6255), .ZN(U3066)
         );
  AOI22_X1 U7234 ( .A1(n6483), .A2(n6257), .B1(n6266), .B2(n6487), .ZN(n6261)
         );
  AOI22_X1 U7235 ( .A1(n6259), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n6419), 
        .B2(n6258), .ZN(n6260) );
  OAI211_X1 U7236 ( .C1(n6262), .C2(n6374), .A(n6261), .B(n6260), .ZN(U3067)
         );
  INV_X1 U7237 ( .A(n6263), .ZN(n6265) );
  AOI22_X1 U7238 ( .A1(n6431), .A2(n6265), .B1(n6430), .B2(n6264), .ZN(n6269)
         );
  AOI22_X1 U7239 ( .A1(n6267), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6379), 
        .B2(n6266), .ZN(n6268) );
  OAI211_X1 U7240 ( .C1(n6392), .C2(n6270), .A(n6269), .B(n6268), .ZN(U3068)
         );
  INV_X1 U7241 ( .A(n6381), .ZN(n6271) );
  NAND2_X1 U7242 ( .A1(n6277), .A2(n6271), .ZN(n6272) );
  NAND2_X1 U7243 ( .A1(n6380), .A2(n6272), .ZN(n6282) );
  INV_X1 U7244 ( .A(n6273), .ZN(n6297) );
  AOI21_X1 U7245 ( .B1(n6275), .B2(n6274), .A(n6297), .ZN(n6278) );
  OAI22_X1 U7246 ( .A1(n4802), .A2(n6279), .B1(n6282), .B2(n6278), .ZN(n6276)
         );
  AOI22_X1 U7247 ( .A1(n6430), .A2(n6297), .B1(n6442), .B2(n6310), .ZN(n6284)
         );
  INV_X1 U7248 ( .A(n6278), .ZN(n6281) );
  AOI21_X1 U7249 ( .B1(n6279), .B2(n6435), .A(n6384), .ZN(n6280) );
  OAI21_X1 U7250 ( .B1(n6282), .B2(n6281), .A(n6280), .ZN(n6299) );
  AOI22_X1 U7251 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6299), .B1(n6379), 
        .B2(n6298), .ZN(n6283) );
  OAI211_X1 U7252 ( .C1(n6302), .C2(n6348), .A(n6284), .B(n6283), .ZN(U3076)
         );
  AOI22_X1 U7253 ( .A1(n6446), .A2(n6297), .B1(n6448), .B2(n6310), .ZN(n6286)
         );
  AOI22_X1 U7254 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6299), .B1(n6393), 
        .B2(n6298), .ZN(n6285) );
  OAI211_X1 U7255 ( .C1(n6302), .C2(n6351), .A(n6286), .B(n6285), .ZN(U3077)
         );
  AOI22_X1 U7256 ( .A1(n6452), .A2(n6297), .B1(n6454), .B2(n6310), .ZN(n6288)
         );
  AOI22_X1 U7257 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6299), .B1(n6352), 
        .B2(n6298), .ZN(n6287) );
  OAI211_X1 U7258 ( .C1(n6302), .C2(n6355), .A(n6288), .B(n6287), .ZN(U3078)
         );
  AOI22_X1 U7259 ( .A1(n6458), .A2(n6297), .B1(n6298), .B2(n6401), .ZN(n6290)
         );
  AOI22_X1 U7260 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6299), .B1(n6460), 
        .B2(n6310), .ZN(n6289) );
  OAI211_X1 U7261 ( .C1(n6302), .C2(n6358), .A(n6290), .B(n6289), .ZN(U3079)
         );
  AOI22_X1 U7262 ( .A1(n6464), .A2(n6297), .B1(n6466), .B2(n6310), .ZN(n6292)
         );
  AOI22_X1 U7263 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6299), .B1(n6405), 
        .B2(n6298), .ZN(n6291) );
  OAI211_X1 U7264 ( .C1(n6302), .C2(n6361), .A(n6292), .B(n6291), .ZN(U3080)
         );
  AOI22_X1 U7265 ( .A1(n6470), .A2(n6297), .B1(n6472), .B2(n6310), .ZN(n6294)
         );
  AOI22_X1 U7266 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6299), .B1(n6409), 
        .B2(n6298), .ZN(n6293) );
  OAI211_X1 U7267 ( .C1(n6302), .C2(n6364), .A(n6294), .B(n6293), .ZN(U3081)
         );
  AOI22_X1 U7268 ( .A1(n6476), .A2(n6297), .B1(n6298), .B2(n6413), .ZN(n6296)
         );
  AOI22_X1 U7269 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6299), .B1(n6478), 
        .B2(n6310), .ZN(n6295) );
  OAI211_X1 U7270 ( .C1(n6302), .C2(n6367), .A(n6296), .B(n6295), .ZN(U3082)
         );
  AOI22_X1 U7271 ( .A1(n6483), .A2(n6297), .B1(n6487), .B2(n6310), .ZN(n6301)
         );
  AOI22_X1 U7272 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6299), .B1(n6419), 
        .B2(n6298), .ZN(n6300) );
  OAI211_X1 U7273 ( .C1(n6302), .C2(n6374), .A(n6301), .B(n6300), .ZN(U3083)
         );
  INV_X1 U7274 ( .A(n6303), .ZN(n6428) );
  OR2_X1 U7275 ( .A1(n6305), .A2(n6304), .ZN(n6425) );
  OAI22_X1 U7276 ( .A1(n6428), .A2(n6309), .B1(n6439), .B2(n6425), .ZN(n6332)
         );
  NAND3_X1 U7277 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6306), .A3(n6504), .ZN(n6342) );
  NOR2_X1 U7278 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6342), .ZN(n6331)
         );
  AOI22_X1 U7279 ( .A1(n6431), .A2(n6332), .B1(n6430), .B2(n6331), .ZN(n6318)
         );
  AOI21_X1 U7280 ( .B1(n6380), .B2(n6309), .A(n6308), .ZN(n6311) );
  NOR3_X1 U7281 ( .A1(n6369), .A2(n6311), .A3(n6310), .ZN(n6316) );
  AOI21_X1 U7282 ( .B1(n6425), .B2(STATE2_REG_2__SCAN_IN), .A(n6312), .ZN(
        n6438) );
  OAI211_X1 U7283 ( .C1(n3238), .C2(n6331), .A(n6426), .B(n6438), .ZN(n6315)
         );
  NOR2_X1 U7284 ( .A1(n6313), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6314) );
  AOI22_X1 U7285 ( .A1(n6333), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n6442), 
        .B2(n6369), .ZN(n6317) );
  OAI211_X1 U7286 ( .C1(n6445), .C2(n6336), .A(n6318), .B(n6317), .ZN(U3084)
         );
  AOI22_X1 U7287 ( .A1(n6447), .A2(n6332), .B1(n6446), .B2(n6331), .ZN(n6320)
         );
  AOI22_X1 U7288 ( .A1(n6333), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n6448), 
        .B2(n6369), .ZN(n6319) );
  OAI211_X1 U7289 ( .C1(n6451), .C2(n6336), .A(n6320), .B(n6319), .ZN(U3085)
         );
  AOI22_X1 U7290 ( .A1(n6453), .A2(n6332), .B1(n6452), .B2(n6331), .ZN(n6322)
         );
  AOI22_X1 U7291 ( .A1(n6333), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n6454), 
        .B2(n6369), .ZN(n6321) );
  OAI211_X1 U7292 ( .C1(n6457), .C2(n6336), .A(n6322), .B(n6321), .ZN(U3086)
         );
  AOI22_X1 U7293 ( .A1(n6459), .A2(n6332), .B1(n6458), .B2(n6331), .ZN(n6324)
         );
  AOI22_X1 U7294 ( .A1(n6333), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n6460), 
        .B2(n6369), .ZN(n6323) );
  OAI211_X1 U7295 ( .C1(n6463), .C2(n6336), .A(n6324), .B(n6323), .ZN(U3087)
         );
  AOI22_X1 U7296 ( .A1(n6465), .A2(n6332), .B1(n6464), .B2(n6331), .ZN(n6326)
         );
  AOI22_X1 U7297 ( .A1(n6333), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n6466), 
        .B2(n6369), .ZN(n6325) );
  OAI211_X1 U7298 ( .C1(n6469), .C2(n6336), .A(n6326), .B(n6325), .ZN(U3088)
         );
  AOI22_X1 U7299 ( .A1(n6471), .A2(n6332), .B1(n6470), .B2(n6331), .ZN(n6328)
         );
  AOI22_X1 U7300 ( .A1(n6333), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n6472), 
        .B2(n6369), .ZN(n6327) );
  OAI211_X1 U7301 ( .C1(n6475), .C2(n6336), .A(n6328), .B(n6327), .ZN(U3089)
         );
  AOI22_X1 U7302 ( .A1(n6477), .A2(n6332), .B1(n6476), .B2(n6331), .ZN(n6330)
         );
  AOI22_X1 U7303 ( .A1(n6333), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n6478), 
        .B2(n6369), .ZN(n6329) );
  OAI211_X1 U7304 ( .C1(n6481), .C2(n6336), .A(n6330), .B(n6329), .ZN(U3090)
         );
  AOI22_X1 U7305 ( .A1(n6485), .A2(n6332), .B1(n6483), .B2(n6331), .ZN(n6335)
         );
  AOI22_X1 U7306 ( .A1(n6333), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n6487), 
        .B2(n6369), .ZN(n6334) );
  OAI211_X1 U7307 ( .C1(n6492), .C2(n6336), .A(n6335), .B(n6334), .ZN(U3091)
         );
  OAI21_X1 U7308 ( .B1(n6337), .B2(n6432), .A(n6380), .ZN(n6345) );
  NOR2_X1 U7309 ( .A1(n6378), .A2(n6342), .ZN(n6368) );
  AOI21_X1 U7310 ( .B1(n6339), .B2(n6338), .A(n6368), .ZN(n6341) );
  OAI22_X1 U7311 ( .A1(n4802), .A2(n6342), .B1(n6345), .B2(n6341), .ZN(n6340)
         );
  AOI22_X1 U7312 ( .A1(n6369), .A2(n6379), .B1(n6430), .B2(n6368), .ZN(n6347)
         );
  INV_X1 U7313 ( .A(n6341), .ZN(n6344) );
  AOI21_X1 U7314 ( .B1(n6435), .B2(n6342), .A(n6384), .ZN(n6343) );
  AOI22_X1 U7315 ( .A1(n6371), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n6442), 
        .B2(n6370), .ZN(n6346) );
  OAI211_X1 U7316 ( .C1(n6375), .C2(n6348), .A(n6347), .B(n6346), .ZN(U3092)
         );
  AOI22_X1 U7317 ( .A1(n6370), .A2(n6448), .B1(n6446), .B2(n6368), .ZN(n6350)
         );
  AOI22_X1 U7318 ( .A1(n6371), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n6393), 
        .B2(n6369), .ZN(n6349) );
  OAI211_X1 U7319 ( .C1(n6375), .C2(n6351), .A(n6350), .B(n6349), .ZN(U3093)
         );
  AOI22_X1 U7320 ( .A1(n6370), .A2(n6454), .B1(n6452), .B2(n6368), .ZN(n6354)
         );
  AOI22_X1 U7321 ( .A1(n6371), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n6352), 
        .B2(n6369), .ZN(n6353) );
  OAI211_X1 U7322 ( .C1(n6375), .C2(n6355), .A(n6354), .B(n6353), .ZN(U3094)
         );
  AOI22_X1 U7323 ( .A1(n6370), .A2(n6460), .B1(n6458), .B2(n6368), .ZN(n6357)
         );
  AOI22_X1 U7324 ( .A1(n6371), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n6401), 
        .B2(n6369), .ZN(n6356) );
  OAI211_X1 U7325 ( .C1(n6375), .C2(n6358), .A(n6357), .B(n6356), .ZN(U3095)
         );
  AOI22_X1 U7326 ( .A1(n6370), .A2(n6466), .B1(n6464), .B2(n6368), .ZN(n6360)
         );
  AOI22_X1 U7327 ( .A1(n6371), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n6405), 
        .B2(n6369), .ZN(n6359) );
  OAI211_X1 U7328 ( .C1(n6375), .C2(n6361), .A(n6360), .B(n6359), .ZN(U3096)
         );
  AOI22_X1 U7329 ( .A1(n6369), .A2(n6409), .B1(n6470), .B2(n6368), .ZN(n6363)
         );
  AOI22_X1 U7330 ( .A1(n6371), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n6472), 
        .B2(n6370), .ZN(n6362) );
  OAI211_X1 U7331 ( .C1(n6375), .C2(n6364), .A(n6363), .B(n6362), .ZN(U3097)
         );
  AOI22_X1 U7332 ( .A1(n6369), .A2(n6413), .B1(n6476), .B2(n6368), .ZN(n6366)
         );
  AOI22_X1 U7333 ( .A1(n6371), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n6478), 
        .B2(n6370), .ZN(n6365) );
  OAI211_X1 U7334 ( .C1(n6375), .C2(n6367), .A(n6366), .B(n6365), .ZN(U3098)
         );
  AOI22_X1 U7335 ( .A1(n6369), .A2(n6419), .B1(n6483), .B2(n6368), .ZN(n6373)
         );
  AOI22_X1 U7336 ( .A1(n6371), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n6487), 
        .B2(n6370), .ZN(n6372) );
  OAI211_X1 U7337 ( .C1(n6375), .C2(n6374), .A(n6373), .B(n6372), .ZN(U3099)
         );
  NOR2_X1 U7338 ( .A1(n6378), .A2(n6387), .ZN(n6417) );
  AOI22_X1 U7339 ( .A1(n6418), .A2(n6379), .B1(n6430), .B2(n6417), .ZN(n6391)
         );
  OAI21_X1 U7340 ( .B1(n6382), .B2(n6381), .A(n6380), .ZN(n6389) );
  AOI21_X1 U7341 ( .B1(n6383), .B2(n6495), .A(n6417), .ZN(n6388) );
  INV_X1 U7342 ( .A(n6388), .ZN(n6386) );
  AOI21_X1 U7343 ( .B1(n6435), .B2(n6387), .A(n6384), .ZN(n6385) );
  OAI22_X1 U7344 ( .A1(n6389), .A2(n6388), .B1(n4802), .B2(n6387), .ZN(n6420)
         );
  AOI22_X1 U7345 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6421), .B1(n6431), 
        .B2(n6420), .ZN(n6390) );
  OAI211_X1 U7346 ( .C1(n6392), .C2(n6491), .A(n6391), .B(n6390), .ZN(U3108)
         );
  AOI22_X1 U7347 ( .A1(n6393), .A2(n6418), .B1(n6446), .B2(n6417), .ZN(n6395)
         );
  AOI22_X1 U7348 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6421), .B1(n6447), 
        .B2(n6420), .ZN(n6394) );
  OAI211_X1 U7349 ( .C1(n6396), .C2(n6491), .A(n6395), .B(n6394), .ZN(U3109)
         );
  INV_X1 U7350 ( .A(n6491), .ZN(n6397) );
  AOI22_X1 U7351 ( .A1(n6454), .A2(n6397), .B1(n6452), .B2(n6417), .ZN(n6399)
         );
  AOI22_X1 U7352 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6421), .B1(n6453), 
        .B2(n6420), .ZN(n6398) );
  OAI211_X1 U7353 ( .C1(n6457), .C2(n6400), .A(n6399), .B(n6398), .ZN(U3110)
         );
  AOI22_X1 U7354 ( .A1(n6401), .A2(n6418), .B1(n6458), .B2(n6417), .ZN(n6403)
         );
  AOI22_X1 U7355 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6421), .B1(n6459), 
        .B2(n6420), .ZN(n6402) );
  OAI211_X1 U7356 ( .C1(n6404), .C2(n6491), .A(n6403), .B(n6402), .ZN(U3111)
         );
  AOI22_X1 U7357 ( .A1(n6405), .A2(n6418), .B1(n6464), .B2(n6417), .ZN(n6407)
         );
  AOI22_X1 U7358 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6421), .B1(n6465), 
        .B2(n6420), .ZN(n6406) );
  OAI211_X1 U7359 ( .C1(n6408), .C2(n6491), .A(n6407), .B(n6406), .ZN(U3112)
         );
  AOI22_X1 U7360 ( .A1(n6409), .A2(n6418), .B1(n6470), .B2(n6417), .ZN(n6411)
         );
  AOI22_X1 U7361 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6421), .B1(n6471), 
        .B2(n6420), .ZN(n6410) );
  OAI211_X1 U7362 ( .C1(n6412), .C2(n6491), .A(n6411), .B(n6410), .ZN(U3113)
         );
  AOI22_X1 U7363 ( .A1(n6413), .A2(n6418), .B1(n6476), .B2(n6417), .ZN(n6415)
         );
  AOI22_X1 U7364 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6421), .B1(n6477), 
        .B2(n6420), .ZN(n6414) );
  OAI211_X1 U7365 ( .C1(n6416), .C2(n6491), .A(n6415), .B(n6414), .ZN(U3114)
         );
  AOI22_X1 U7366 ( .A1(n6419), .A2(n6418), .B1(n6483), .B2(n6417), .ZN(n6423)
         );
  AOI22_X1 U7367 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6421), .B1(n6485), 
        .B2(n6420), .ZN(n6422) );
  OAI211_X1 U7368 ( .C1(n6424), .C2(n6491), .A(n6423), .B(n6422), .ZN(U3115)
         );
  OAI22_X1 U7369 ( .A1(n6428), .A2(n6427), .B1(n6426), .B2(n6425), .ZN(n6484)
         );
  NOR2_X1 U7370 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6429), .ZN(n6482)
         );
  AOI22_X1 U7371 ( .A1(n6431), .A2(n6484), .B1(n6430), .B2(n6482), .ZN(n6444)
         );
  INV_X1 U7372 ( .A(n6486), .ZN(n6433) );
  AOI21_X1 U7373 ( .B1(n6491), .B2(n6433), .A(n6432), .ZN(n6434) );
  AOI211_X1 U7374 ( .C1(n6437), .C2(n6436), .A(n6435), .B(n6434), .ZN(n6441)
         );
  OAI211_X1 U7375 ( .C1(n3238), .C2(n6482), .A(n6439), .B(n6438), .ZN(n6440)
         );
  AOI22_X1 U7376 ( .A1(n6488), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n6442), 
        .B2(n6486), .ZN(n6443) );
  OAI211_X1 U7377 ( .C1(n6445), .C2(n6491), .A(n6444), .B(n6443), .ZN(U3116)
         );
  AOI22_X1 U7378 ( .A1(n6447), .A2(n6484), .B1(n6446), .B2(n6482), .ZN(n6450)
         );
  AOI22_X1 U7379 ( .A1(n6488), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n6448), 
        .B2(n6486), .ZN(n6449) );
  OAI211_X1 U7380 ( .C1(n6451), .C2(n6491), .A(n6450), .B(n6449), .ZN(U3117)
         );
  AOI22_X1 U7381 ( .A1(n6453), .A2(n6484), .B1(n6452), .B2(n6482), .ZN(n6456)
         );
  AOI22_X1 U7382 ( .A1(n6488), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n6454), 
        .B2(n6486), .ZN(n6455) );
  OAI211_X1 U7383 ( .C1(n6457), .C2(n6491), .A(n6456), .B(n6455), .ZN(U3118)
         );
  AOI22_X1 U7384 ( .A1(n6459), .A2(n6484), .B1(n6458), .B2(n6482), .ZN(n6462)
         );
  AOI22_X1 U7385 ( .A1(n6488), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n6460), 
        .B2(n6486), .ZN(n6461) );
  OAI211_X1 U7386 ( .C1(n6463), .C2(n6491), .A(n6462), .B(n6461), .ZN(U3119)
         );
  AOI22_X1 U7387 ( .A1(n6465), .A2(n6484), .B1(n6464), .B2(n6482), .ZN(n6468)
         );
  AOI22_X1 U7388 ( .A1(n6488), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n6466), 
        .B2(n6486), .ZN(n6467) );
  OAI211_X1 U7389 ( .C1(n6469), .C2(n6491), .A(n6468), .B(n6467), .ZN(U3120)
         );
  AOI22_X1 U7390 ( .A1(n6471), .A2(n6484), .B1(n6470), .B2(n6482), .ZN(n6474)
         );
  AOI22_X1 U7391 ( .A1(n6488), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n6472), 
        .B2(n6486), .ZN(n6473) );
  OAI211_X1 U7392 ( .C1(n6475), .C2(n6491), .A(n6474), .B(n6473), .ZN(U3121)
         );
  AOI22_X1 U7393 ( .A1(n6477), .A2(n6484), .B1(n6476), .B2(n6482), .ZN(n6480)
         );
  AOI22_X1 U7394 ( .A1(n6488), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n6478), 
        .B2(n6486), .ZN(n6479) );
  OAI211_X1 U7395 ( .C1(n6481), .C2(n6491), .A(n6480), .B(n6479), .ZN(U3122)
         );
  AOI22_X1 U7396 ( .A1(n6485), .A2(n6484), .B1(n6483), .B2(n6482), .ZN(n6490)
         );
  AOI22_X1 U7397 ( .A1(n6488), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n6487), 
        .B2(n6486), .ZN(n6489) );
  OAI211_X1 U7398 ( .C1(n6492), .C2(n6491), .A(n6490), .B(n6489), .ZN(U3123)
         );
  INV_X1 U7399 ( .A(n6508), .ZN(n6513) );
  INV_X1 U7400 ( .A(n6493), .ZN(n6494) );
  NAND2_X1 U7401 ( .A1(n6495), .A2(n6494), .ZN(n6498) );
  NAND2_X1 U7402 ( .A1(n6496), .A2(n3064), .ZN(n6497) );
  NAND2_X1 U7403 ( .A1(n6498), .A2(n6497), .ZN(n6639) );
  NAND2_X1 U7404 ( .A1(n6499), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6648) );
  NAND2_X1 U7405 ( .A1(n6648), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6500) );
  OR2_X1 U7406 ( .A1(n6639), .A2(n6500), .ZN(n6503) );
  NAND2_X1 U7407 ( .A1(n6503), .A2(n6504), .ZN(n6506) );
  OAI211_X1 U7408 ( .C1(n6504), .C2(n6503), .A(n6502), .B(n6501), .ZN(n6505)
         );
  OAI211_X1 U7409 ( .C1(n6507), .C2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(n6506), .B(n6505), .ZN(n6511) );
  NAND2_X1 U7410 ( .A1(n6507), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6510) );
  AOI22_X1 U7411 ( .A1(n6511), .A2(n6510), .B1(n6509), .B2(n6508), .ZN(n6512)
         );
  AOI211_X1 U7412 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6513), .A(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B(n6512), .ZN(n6522) );
  INV_X1 U7413 ( .A(n6514), .ZN(n6520) );
  OAI21_X1 U7414 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6515), 
        .ZN(n6516) );
  NAND3_X1 U7415 ( .A1(n6518), .A2(n6517), .A3(n6516), .ZN(n6519) );
  NOR4_X1 U7416 ( .A1(n6522), .A2(n6521), .A3(n6520), .A4(n6519), .ZN(n6535)
         );
  INV_X1 U7417 ( .A(n6535), .ZN(n6524) );
  OAI22_X1 U7418 ( .A1(n6524), .A2(n6537), .B1(n6523), .B2(n6660), .ZN(n6525)
         );
  OAI21_X1 U7419 ( .B1(n6527), .B2(n6526), .A(n6525), .ZN(n6632) );
  OAI21_X1 U7420 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6660), .A(n6632), .ZN(
        n6536) );
  AOI221_X1 U7421 ( .B1(n6529), .B2(STATE2_REG_0__SCAN_IN), .C1(n6536), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6528), .ZN(n6534) );
  OAI211_X1 U7422 ( .C1(n6532), .C2(n6531), .A(n6530), .B(n6632), .ZN(n6533)
         );
  OAI211_X1 U7423 ( .C1(n6535), .C2(n6537), .A(n6534), .B(n6533), .ZN(U3148)
         );
  NAND3_X1 U7424 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6543), .A3(n6536), .ZN(
        n6542) );
  OAI21_X1 U7425 ( .B1(READY_N), .B2(n6538), .A(n6537), .ZN(n6540) );
  AOI21_X1 U7426 ( .B1(n6540), .B2(n6632), .A(n6539), .ZN(n6541) );
  NAND2_X1 U7427 ( .A1(n6542), .A2(n6541), .ZN(U3149) );
  OAI211_X1 U7428 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6660), .A(n6543), .B(
        n6630), .ZN(n6545) );
  OAI21_X1 U7429 ( .B1(n6663), .B2(n6545), .A(n6544), .ZN(U3150) );
  AND2_X1 U7430 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6548), .ZN(U3151) );
  AND2_X1 U7431 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6548), .ZN(U3152) );
  AND2_X1 U7432 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6548), .ZN(U3153) );
  AND2_X1 U7433 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6548), .ZN(U3154) );
  NOR2_X1 U7434 ( .A1(n6629), .A2(n6546), .ZN(U3155) );
  AND2_X1 U7435 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6548), .ZN(U3156) );
  AND2_X1 U7436 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6548), .ZN(U3157) );
  NOR2_X1 U7437 ( .A1(n6629), .A2(n6547), .ZN(U3158) );
  AND2_X1 U7438 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6548), .ZN(U3159) );
  AND2_X1 U7439 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6548), .ZN(U3160) );
  AND2_X1 U7440 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6548), .ZN(U3161) );
  AND2_X1 U7441 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6548), .ZN(U3162) );
  AND2_X1 U7442 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6548), .ZN(U3163) );
  AND2_X1 U7443 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6548), .ZN(U3164) );
  AND2_X1 U7444 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6548), .ZN(U3165) );
  AND2_X1 U7445 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6548), .ZN(U3166) );
  AND2_X1 U7446 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6548), .ZN(U3167) );
  AND2_X1 U7447 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6548), .ZN(U3168) );
  AND2_X1 U7448 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6548), .ZN(U3169) );
  AND2_X1 U7449 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6548), .ZN(U3170) );
  AND2_X1 U7450 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6548), .ZN(U3171) );
  AND2_X1 U7451 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6548), .ZN(U3172) );
  AND2_X1 U7452 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6548), .ZN(U3173) );
  AND2_X1 U7453 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6548), .ZN(U3174) );
  AND2_X1 U7454 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6548), .ZN(U3175) );
  AND2_X1 U7455 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6548), .ZN(U3176) );
  AND2_X1 U7456 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6548), .ZN(U3177) );
  AND2_X1 U7457 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6548), .ZN(U3178) );
  AND2_X1 U7458 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6548), .ZN(U3179) );
  AND2_X1 U7459 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6548), .ZN(U3180) );
  NOR2_X1 U7460 ( .A1(n6549), .A2(n6565), .ZN(n6551) );
  NAND2_X1 U7461 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6553) );
  NAND2_X1 U7462 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .ZN(n6563) );
  AND2_X1 U7463 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6554) );
  INV_X1 U7464 ( .A(NA_N), .ZN(n6557) );
  AOI221_X1 U7465 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6557), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6562) );
  AOI221_X1 U7466 ( .B1(n6554), .B2(n6668), .C1(n6552), .C2(n6668), .A(n6562), 
        .ZN(n6550) );
  OAI221_X1 U7467 ( .B1(n6551), .B2(n6553), .C1(n6551), .C2(n6563), .A(n6550), 
        .ZN(U3181) );
  NOR2_X1 U7468 ( .A1(n6559), .A2(n6552), .ZN(n6558) );
  OAI21_X1 U7469 ( .B1(n6558), .B2(n6554), .A(n6553), .ZN(n6555) );
  NAND3_X1 U7470 ( .A1(n6556), .A2(n6563), .A3(n6555), .ZN(U3182) );
  AOI21_X1 U7471 ( .B1(n6558), .B2(n6557), .A(STATE_REG_2__SCAN_IN), .ZN(n6564) );
  AOI221_X1 U7472 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6660), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6560) );
  AOI221_X1 U7473 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6560), .C2(HOLD), .A(n6559), .ZN(n6561) );
  OAI22_X1 U7474 ( .A1(n6564), .A2(n6563), .B1(n6562), .B2(n6561), .ZN(U3183)
         );
  NAND2_X1 U7475 ( .A1(n6565), .A2(n6613), .ZN(n6624) );
  AOI22_X1 U7476 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6618), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6657), .ZN(n6566) );
  OAI21_X1 U7477 ( .B1(n5390), .B2(n6620), .A(n6566), .ZN(U3184) );
  AOI22_X1 U7478 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6618), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6657), .ZN(n6567) );
  OAI21_X1 U7479 ( .B1(n6568), .B2(n6620), .A(n6567), .ZN(U3185) );
  AOI22_X1 U7480 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6618), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6668), .ZN(n6569) );
  OAI21_X1 U7481 ( .B1(n6570), .B2(n6620), .A(n6569), .ZN(U3186) );
  AOI22_X1 U7482 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6618), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6668), .ZN(n6571) );
  OAI21_X1 U7483 ( .B1(n6572), .B2(n6620), .A(n6571), .ZN(U3187) );
  AOI22_X1 U7484 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6618), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6668), .ZN(n6573) );
  OAI21_X1 U7485 ( .B1(n6574), .B2(n6620), .A(n6573), .ZN(U3188) );
  AOI22_X1 U7486 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6618), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6668), .ZN(n6575) );
  OAI21_X1 U7487 ( .B1(n6576), .B2(n6620), .A(n6575), .ZN(U3189) );
  AOI22_X1 U7488 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6618), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6657), .ZN(n6577) );
  OAI21_X1 U7489 ( .B1(n6578), .B2(n6620), .A(n6577), .ZN(U3190) );
  AOI22_X1 U7490 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6618), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6668), .ZN(n6579) );
  OAI21_X1 U7491 ( .B1(n6580), .B2(n6620), .A(n6579), .ZN(U3191) );
  AOI22_X1 U7492 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6622), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6657), .ZN(n6581) );
  OAI21_X1 U7493 ( .B1(n6583), .B2(n6624), .A(n6581), .ZN(U3192) );
  AOI22_X1 U7494 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6618), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6657), .ZN(n6582) );
  OAI21_X1 U7495 ( .B1(n6583), .B2(n6620), .A(n6582), .ZN(U3193) );
  AOI22_X1 U7496 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6622), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6657), .ZN(n6584) );
  OAI21_X1 U7497 ( .B1(n6587), .B2(n6624), .A(n6584), .ZN(U3194) );
  OAI222_X1 U7498 ( .A1(n6620), .A2(n6587), .B1(n6586), .B2(n6613), .C1(n6585), 
        .C2(n6624), .ZN(U3195) );
  AOI22_X1 U7499 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6622), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6657), .ZN(n6588) );
  OAI21_X1 U7500 ( .B1(n6590), .B2(n6624), .A(n6588), .ZN(U3196) );
  AOI22_X1 U7501 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6618), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6657), .ZN(n6589) );
  OAI21_X1 U7502 ( .B1(n6590), .B2(n6620), .A(n6589), .ZN(U3197) );
  AOI22_X1 U7503 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6622), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6657), .ZN(n6591) );
  OAI21_X1 U7504 ( .B1(n6592), .B2(n6624), .A(n6591), .ZN(U3198) );
  AOI22_X1 U7505 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6622), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6657), .ZN(n6593) );
  OAI21_X1 U7506 ( .B1(n6594), .B2(n6624), .A(n6593), .ZN(U3199) );
  AOI22_X1 U7507 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6622), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6657), .ZN(n6595) );
  OAI21_X1 U7508 ( .B1(n6598), .B2(n6624), .A(n6595), .ZN(U3200) );
  OAI222_X1 U7509 ( .A1(n6620), .A2(n6598), .B1(n6597), .B2(n6613), .C1(n6596), 
        .C2(n6624), .ZN(U3201) );
  AOI22_X1 U7510 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6622), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6668), .ZN(n6599) );
  OAI21_X1 U7511 ( .B1(n6601), .B2(n6624), .A(n6599), .ZN(U3202) );
  AOI22_X1 U7512 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6618), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6657), .ZN(n6600) );
  OAI21_X1 U7513 ( .B1(n6601), .B2(n6620), .A(n6600), .ZN(U3203) );
  AOI22_X1 U7514 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6618), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6657), .ZN(n6602) );
  OAI21_X1 U7515 ( .B1(n6603), .B2(n6620), .A(n6602), .ZN(U3204) );
  AOI22_X1 U7516 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6618), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6657), .ZN(n6604) );
  OAI21_X1 U7517 ( .B1(n6605), .B2(n6620), .A(n6604), .ZN(U3205) );
  AOI22_X1 U7518 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6622), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6657), .ZN(n6606) );
  OAI21_X1 U7519 ( .B1(n6607), .B2(n6624), .A(n6606), .ZN(U3206) );
  OAI222_X1 U7520 ( .A1(n6624), .A2(n6609), .B1(n6608), .B2(n6613), .C1(n6607), 
        .C2(n6620), .ZN(U3207) );
  INV_X1 U7521 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6612) );
  AOI22_X1 U7522 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6622), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6668), .ZN(n6610) );
  OAI21_X1 U7523 ( .B1(n6612), .B2(n6624), .A(n6610), .ZN(U3208) );
  AOI22_X1 U7524 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6618), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6657), .ZN(n6611) );
  OAI21_X1 U7525 ( .B1(n6612), .B2(n6620), .A(n6611), .ZN(U3209) );
  INV_X1 U7526 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6617) );
  OAI222_X1 U7527 ( .A1(n6620), .A2(n6615), .B1(n6614), .B2(n6613), .C1(n6617), 
        .C2(n6624), .ZN(U3210) );
  AOI22_X1 U7528 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6618), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6657), .ZN(n6616) );
  OAI21_X1 U7529 ( .B1(n6617), .B2(n6620), .A(n6616), .ZN(U3211) );
  AOI22_X1 U7530 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6618), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6657), .ZN(n6619) );
  OAI21_X1 U7531 ( .B1(n6621), .B2(n6620), .A(n6619), .ZN(U3212) );
  AOI22_X1 U7532 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6622), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6657), .ZN(n6623) );
  OAI21_X1 U7533 ( .B1(n6625), .B2(n6624), .A(n6623), .ZN(U3213) );
  MUX2_X1 U7534 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n6668), .Z(U3445) );
  MUX2_X1 U7535 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6668), .Z(U3446) );
  MUX2_X1 U7536 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6668), .Z(U3447) );
  MUX2_X1 U7537 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6668), .Z(U3448) );
  OAI21_X1 U7538 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6629), .A(n6627), .ZN(
        n6626) );
  INV_X1 U7539 ( .A(n6626), .ZN(U3451) );
  OAI21_X1 U7540 ( .B1(n6629), .B2(n6628), .A(n6627), .ZN(U3452) );
  OAI211_X1 U7541 ( .C1(n6632), .C2(n3238), .A(n6631), .B(n6630), .ZN(U3453)
         );
  AOI22_X1 U7542 ( .A1(n6636), .A2(n6635), .B1(n6634), .B2(n6633), .ZN(n6637)
         );
  INV_X1 U7543 ( .A(n6637), .ZN(n6638) );
  MUX2_X1 U7544 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6638), .S(n6645), 
        .Z(U3456) );
  INV_X1 U7545 ( .A(n6639), .ZN(n6643) );
  AOI21_X1 U7546 ( .B1(STATE2_REG_1__SCAN_IN), .B2(n6641), .A(n6640), .ZN(
        n6642) );
  OAI211_X1 U7547 ( .C1(n6643), .C2(n6647), .A(n6645), .B(n6642), .ZN(n6644)
         );
  OAI21_X1 U7548 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6645), .A(n6644), 
        .ZN(n6646) );
  OAI21_X1 U7549 ( .B1(n6648), .B2(n6647), .A(n6646), .ZN(U3461) );
  AOI21_X1 U7550 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6649) );
  AOI22_X1 U7551 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6649), .B2(n5390), .ZN(n6652) );
  INV_X1 U7552 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6651) );
  AOI22_X1 U7553 ( .A1(n6655), .A2(n6652), .B1(n6651), .B2(n6650), .ZN(U3468)
         );
  INV_X1 U7554 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6654) );
  OAI21_X1 U7555 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6655), .ZN(n6653) );
  OAI21_X1 U7556 ( .B1(n6655), .B2(n6654), .A(n6653), .ZN(U3469) );
  NAND2_X1 U7557 ( .A1(n6657), .A2(W_R_N_REG_SCAN_IN), .ZN(n6656) );
  OAI21_X1 U7558 ( .B1(n6657), .B2(READREQUEST_REG_SCAN_IN), .A(n6656), .ZN(
        U3470) );
  AOI211_X1 U7559 ( .C1(n6016), .C2(n6660), .A(n6659), .B(n6658), .ZN(n6667)
         );
  OAI211_X1 U7560 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6662), .A(n6661), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6664) );
  AOI21_X1 U7561 ( .B1(n6664), .B2(STATE2_REG_0__SCAN_IN), .A(n6663), .ZN(
        n6666) );
  NAND2_X1 U7562 ( .A1(n6667), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6665) );
  OAI21_X1 U7563 ( .B1(n6667), .B2(n6666), .A(n6665), .ZN(U3472) );
  MUX2_X1 U7564 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n6668), .Z(U3473) );
  INV_X1 U4248 ( .A(n3243), .ZN(n4003) );
  NAND2_X2 U4034 ( .A1(n4483), .A2(n5269), .ZN(n4008) );
  MUX2_X1 U5044 ( .A(n4214), .B(n4008), .S(n4577), .Z(n4005) );
  CLKBUF_X1 U3439 ( .A(n3265), .Z(n3266) );
  AND4_X1 U3450 ( .A1(n3135), .A2(n3134), .A3(n3133), .A4(n3132), .ZN(n3136)
         );
  CLKBUF_X1 U34520 ( .A(n4651), .Z(n4652) );
  CLKBUF_X1 U3457 ( .A(n3418), .Z(n6495) );
  CLKBUF_X1 U3775 ( .A(n5281), .Z(n5314) );
  CLKBUF_X1 U3832 ( .A(n3236), .Z(n4248) );
  XNOR2_X1 U4174 ( .A(n3004), .B(n4185), .ZN(n5052) );
endmodule

