
module b14_C_2inp_gates_syn ( 
    DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
    DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
    DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
    DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
    DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
    DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, REG3_REG_27__SCAN_IN,
    REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, REG3_REG_10__SCAN_IN,
    REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, REG3_REG_28__SCAN_IN,
    REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, REG3_REG_21__SCAN_IN,
    REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, REG3_REG_16__SCAN_IN,
    REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, REG3_REG_24__SCAN_IN,
    REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, REG3_REG_0__SCAN_IN,
    REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, IR_REG_0__SCAN_IN,
    IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, IR_REG_3__SCAN_IN,
    IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN,
    IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN,
    IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN,
    IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN,
    IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN,
    IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN,
    IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, IR_REG_24__SCAN_IN,
    IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN,
    IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, IR_REG_30__SCAN_IN,
    IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, D_REG_1__SCAN_IN,
    D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, D_REG_5__SCAN_IN,
    D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
    D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
    D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
    D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
    D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
    D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
    D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
    D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
    D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
    REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
    REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
    REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
    REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
    REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
    REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
    REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
    REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
    REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
    REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
    REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
    REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
    REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
    REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
    REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
    REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
    REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
    REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
    REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
    REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
    REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
    REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
    REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
    REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
    REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
    REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
    REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
    REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
    REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
    REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
    REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
    REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
    ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
    ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
    ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
    ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
    ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
    ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
    DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
    DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
    DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
    DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
    DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
    DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
    DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
    DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
    DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
    DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
    DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
    REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
    REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
    REG3_REG_22__SCAN_IN,
    U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
    U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
    U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
    U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
    U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
    U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
    U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
    U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
    U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
    U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
    U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
    U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
    U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
    U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
    U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
    U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
    U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
    U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
    U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
    U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
    U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
    U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
    U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
    U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
    U3211, U3210, U3149, U3148, U4043  );
  input  DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_,
    DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_,
    DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_,
    DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_,
    DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_,
    DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
    REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
    REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
    REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
    REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
    REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
    REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
    REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
    IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
    IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
    IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
    IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
    IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
    IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
    IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
    IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
    IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
    IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
    IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
    D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN,
    D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN,
    D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN,
    D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN,
    D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN,
    D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN,
    D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN,
    D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN,
    D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN,
    D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN,
    REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN,
    REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN,
    REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN,
    REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN,
    REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN,
    REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN,
    REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN,
    REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN,
    REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN,
    REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN,
    REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN,
    REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN,
    REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN,
    REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN,
    REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN,
    REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN,
    REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN,
    REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN,
    REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN,
    REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN,
    REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN,
    REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN,
    REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN,
    REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN,
    REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN,
    REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN,
    REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN,
    REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN,
    REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN,
    REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN,
    REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN,
    REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN,
    ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN,
    ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN,
    ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN,
    ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN,
    ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN,
    ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN,
    ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
    DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
    DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
    DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
    DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
    DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
    DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
    DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
    DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
    DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
    DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
    B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN,
    REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN,
    REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
    U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
    U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
    U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
    U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
    U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
    U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
    U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
    U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
    U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
    U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
    U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
    U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
    U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
    U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
    U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
    U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
    U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
    U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
    U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
    U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
    U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
    U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
    U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
    U3211, U3210, U3149, U3148, U4043;
  wire n4545, n6589, n5348, n5994, n6725, n7684, n7574, n4360, n6898, n5456,
    n7516, n7712, n4948, n4920, n4716, n7680, n7164, n5372, n5188, n4620,
    n4614, n4358, n4759, n7979, n7309, n7486, n5700, n4730, n7618, n5544,
    n4359, n5804, n6661, n4589, n7282, n5808, n6368, n7252, n5646, n6457,
    n6547, n6456, n4991, n6561, n5859, n5327, n4541, n4543, n7612, n6859,
    n6967, n6345, n6144, n5778, n7617, n7314, n7351, n7394, n7583, n7316,
    n7651, n4711, n4816, n7572, n5496, n6854, n7858, n5688, n4442, n6015,
    n5267, n4891, n4617, n5441, n4616, n5314, n4637, n4965, n4613, n5312,
    n4855, n4768, n4769, n4600, n4789, n4601, n5689, n5665, n4361, n4362,
    n5172, n4918, n4812, n5635, n5502, n5329, n4484, n4483, n4481, n5639,
    n5619, n4516, n4448, n4449, n4450, n4582, n4715, n4694, n4757, n7194,
    n4540, n6136, n7599, n7598, n7571, n7534, n7901, n4404, n7474, n4558,
    n4497, n4519, n5606, n4544, n4406, n4554, n7560, n4426, n4421, n5280,
    n4672, n5862, n4569, n4583, n5021, n7563, n5071, n5018, n5020, n4654,
    n4517, n5959, n5353, n5367, n4523, n4524, n7166, n5331, n4472, n4475,
    n5386, n5393, n4507, n6102, n4508, n6357, n6396, n6516, n4511, n4512,
    n6562, n7379, n7376, n4453, n4454, n7427, n7415, n4444, n7470, n7529,
    n7629, n7645, n7670, n5263, n4574, n4665, n7315, n4584, n4581, n4570,
    n4571, n4572, n6990, n4562, n4565, n4651, n6023, n4413, n7043, n7137,
    n7222, n7246, n5333, n4491, n4489, n4487, n7671, n4417, n4415, n4416,
    n6429, n7398, n4500, n4428, n4430, n6256, n7720, n4551, n4550, n4552,
    n6664, n6074, n6073, n4482, n4532, n4438, n4423, n4468, n4477, n4476,
    n4473, n4527, n4528, n4549, n4433, n4434, n4548, n4402, n4400, n4401,
    n4590, n4419, n4420, n4452, n4418, n4455, n4445, n4542, n5610, n5863,
    n5151, n6878, n5076, n5051, n4557, n6939, n6820, n6919, n5091, n7046,
    n5317, n5357, n4462, n5323, n4465, n4466, n4463, n5377, n4492, n4488,
    n4490, n5521, n5191, n5095, n7365, n6921, n4435, n5574, n5541, n6255,
    n4431, n4432, n4547, n4546, n4399, n6335, n6591, n6595, n4409, n6611,
    n6733, n5572, n7332, n4515, n4514, n7381, n7416, n5570, n7674, n4553,
    n5283, n4609, n4610, n4611, n4705, n5532, n4567, n4568, n4513, n4561,
    n5114, n4578, n4577, n6846, n6845, n6610, n5892, n6954, n6963, n5960,
    n6732, n5155, n4877, n5439, n7083, n7076, n7107, n7150, n4486, n7192,
    n4478, n4533, n7258, n4537, n4536, n4539, n6275, n4505, n4506, n6631,
    n5133, n6723, n4502, n4811, n4622, n7646, n7709, n6299, n4456, n4457,
    n4458, n6518, n4504, n4587, n4607, n4642, n5264, n4770, n4725, n4726,
    n5802, n6991, n5945, n6974, n6979, n6951, n5741, n4563, n7007, n7958,
    n5031, n6840, n7451, n4817, n4686, n4701, n4787, n4439, n7034, n4493,
    n7266, n6620, n4510, n7397, n7632, n6746, n4509, n6634, n4427, n4631,
    n5061, n7747, n7750, n7753, n7768, n7053, n5404, n4767, n7504, n6542,
    n4363, n4364, n4365, n4503, n4886, n5153, n5577, n5567, n5855, n4366,
    n4367, n7446, n4368, n4632, n5943, n5602, n5321, n4647, n5860, n4369,
    n4628, n4370, n4371, n4372, n4373, n4374, n4375, n7468, n4376, n4377,
    n4378, n6309, n4579, n4580, n4379, n4380, n4381, n4382, n4383, n4384,
    n5224, n7377, n6170, n4410, n5972, n5265, n4386, n4387, n7330, n7352,
    n6517, n4429, n4485, n4388, n4389, n4390, n4391, n7443, n4392, n4393,
    n5345, n7676, n4394, n4395, n7514, n4396, n4397, n4398, n4407, n6278,
    n4403, n5660, n4405, n6308, n4408, n5618, n4411, n4412, n5525, n5761,
    n4414, n4422, n4424, n4425, n4556, n7615, n4436, n7472, n5512, n7308,
    n6338, n6375, n4437, n4440, n4441, n4443, n4446, n4447, n4451, n6333,
    n4460, n4459, n5429, n4461, n7126, n4464, n5320, n4467, n4469, n4470,
    n7097, n4471, n4474, n7209, n4480, n4479, n7183, n7181, n7239, n4494,
    n4495, n4499, n4498, n4496, n7154, n7976, n5615, n4501, n6329, n5375,
    n4518, n4520, n4521, n7177, n4522, n7119, n4525, n4526, n4531, n7232,
    n4529, n4530, n5401, n4534, n4535, n4538, n7447, n6279, n4643, n7589,
    n4555, n5026, n6997, n6832, n4559, n4560, n4801, n5736, n4564, n4566,
    n4666, n4573, n4575, n5082, n4576, n5822, n7611, n4657, n4687, n4894,
    n4890, n4585, n4586, n4588, n8005, n4591, n4592, n4593, n4594, n6549,
    n4595, n4596, n7452, n5498, n4597, n6583, n5902, n4598, n5630, n5025,
    n5376, n6532, n6875, n4903, n6152, n5549, n4993, n4754, n5890, n5013,
    n7002, n4873, n5366, n5383, n5392, n6543, n4627, n6879, n5209, n6941,
    n7450, n5609, n5535, n5826, n4848, n7714, n7512, n7706, n5581, n7368,
    n5680, n6966, n6988, n5289, n4681, n7707, n4878, n6955, n7009, n6798,
    n6315, n5969, n5682, n5766, n7985, n7982, n7393, n7277, n7284, n8000,
    n7774, n4599, n4603, n4602, n4605, n4604, n4606, n4703, n4608, n4612,
    n4645, n5281, n4652, n4615, n7722, n7723, n4621, n4619, n4682, n4618,
    n4626, n4624, n4760, n4809, n7546, n4623, n4625, n7503, n4971, n4629,
    n4630, n4664, n4633, n4635, n4636, n4634, n4638, n4639, n6105, n4640,
    n4641, n4644, n5419, n4646, n4648, n4649, n5416, n4650, n4743, n4934,
    n4663, n5774, n4656, n4653, n4655, n4771, n4857, n4658, n7765, n4659,
    n4661, n4660, n4662, n4674, n4667, n4668, n4671, n4669, n4670, n4673,
    n5666, n6216, n5278, n4803, n7784, n4907, n4676, n4675, n4804, n7001,
    n4720, n4678, n4677, n4679, n7553, n4680, n4684, n4683, n4685, n4693,
    n4688, n4689, n4691, n4690, n4692, n4696, n4695, n4723, n4698, n4697,
    n4702, n4700, n7602, n4699, n4710, n4790, n4704, n4706, n7079, n4708,
    n6020, n4707, n4709, n4712, n4722, n4714, n7584, n4713, n4721, n6895,
    n4719, n4717, n4718, n7000, n6909, n4802, n4724, n4732, n4728, n4727,
    n4729, n4731, n4733, n4735, n4734, n4756, n6858, n4737, n4736, n4739,
    n4738, n4748, n4740, n4742, n4741, n5568, n5578, n4746, n4744, n4745,
    n4747, n4750, n4749, n4753, n4752, n4751, n5457, n4755, n4758, n4762,
    n4761, n4766, n4764, n4763, n4765, n4775, n4773, n4772, n4774, n4776,
    n4780, n4778, n7652, n4777, n4779, n4782, n4781, n6980, n4784, n4783,
    n4788, n4786, n4785, n4793, n5352, n4791, n4792, n4794, n4798, n4796,
    n4795, n4797, n4800, n4799, n6833, n6894, n6998, n4806, n4805, n4808,
    n4807, n4815, n4810, n4813, n7521, n4814, n4824, n4818, n4819, n4835,
    n7762, n4820, n4822, n4821, n4823, n4825, n4980, n4827, n4826, n4981,
    n6796, n4829, n4828, n4833, n4831, n7465, n4830, n4832, n4841, n4834,
    n4836, n4837, n7759, n4839, n4838, n4840, n4842, n4983, n4844, n7471,
    n4843, n4984, n4845, n4847, n4846, n4853, n4851, n4849, n4945, n7387,
    n4850, n4852, n4867, n4854, n4856, n4926, n4859, n4858, n4860, n4900,
    n4861, n4862, n4863, n4865, n4864, n4866, n4868, n4915, n4870, n4869,
    n4914, n4895, n7435, n4871, n4872, n4875, n4874, n4876, n4885, n4883,
    n4881, n4879, n5326, n4880, n4882, n4884, n4889, n4888, n4887, n5019,
    n6964, n4893, n4892, n4899, n4896, n6952, n4897, n7407, n4898, n4906,
    n4904, n4902, n4901, n4905, n4909, n7405, n4908, n5017, n4910, n4913,
    n4912, n4911, n6873, n4917, n4916, n4925, n4923, n4919, n6915, n4921,
    n7440, n4922, n4924, n4932, n4927, n7756, n4928, n4930, n4929, n4931,
    n4933, n4937, n4936, n4935, n4938, n4940, n4939, n4941, n6917, n4942,
    n6937, n4944, n4943, n4953, n4951, n4946, n4949, n4947, n7336, n4950,
    n4952, n4959, n4954, n7744, n4955, n4957, n4956, n4958, n4960, n5014,
    n4962, n4961, n4964, n4963, n4970, n4968, n5029, n4966, n7305, n4967,
    n4969, n4976, n4972, n7741, n4974, n4973, n4975, n4977, n4992, n4979,
    n4978, n5023, n4988, n4982, n5856, n4986, n4985, n4987, n4989, n4990,
    n4995, n4994, n4997, n4996, n5001, n4999, n7292, n4998, n5000, n5008,
    n5002, n5003, n5033, n7738, n5004, n5006, n5005, n5007, n5009, n5867,
    n5011, n5010, n5980, n5012, n5016, n5015, n6962, n6872, n5022, n5024,
    n5050, n5028, n5027, n5055, n5877, n5030, n5039, n5032, n5034, n5035,
    n7735, n5037, n5036, n5038, n5040, n5043, n5042, n6598, n5041, n5044,
    n5046, n5045, n5047, n5875, n5048, n5049, n5052, n5889, n5054, n5053,
    n5060, n5897, n5058, n5056, n5057, n5059, n7961, n5066, n5062, n7732,
    n5064, n5063, n5065, n5067, n5070, n5069, n5068, n5887, n5073, n5072,
    n5075, n5074, n5081, n5967, n5079, n5077, n5078, n5080, n7964, n5087,
    n5083, n7729, n5085, n5084, n5086, n5088, n5092, n5090, n5089, n5961,
    n5094, n5093, n5099, n6521, n5097, n5096, n5098, n5177, n5103, n5101,
    n5100, n5102, n5104, n5107, n7967, n5106, n5105, n5108, n5111, n5110,
    n5109, n5112, n5823, n5113, n5929, n5395, n6495, n5121, n5116, n5115,
    n5119, n5117, n5118, n5120, n7970, n5123, n6489, n5122, n5124, n5127,
    n5126, n5621, n5125, n5128, n5837, n5147, n5130, n5129, n5927, n5132,
    n5131, n5138, n5844, n5136, n5134, n5135, n5137, n7973, n5140, n6448,
    n5139, n5141, n5840, n5143, n6437, n5142, n5839, n5144, n5145, n5146,
    n5148, n5150, n5149, n5157, n6423, n5152, n5154, n5156, n5159, n6419,
    n5158, n5160, n5163, n5162, n6410, n5161, n5164, n5168, n5166, n5165,
    n5167, n5944, n5169, n5171, n5170, n5176, n5174, n6399, n5173, n5175,
    n5179, n5815, n5178, n5180, n5185, n5199, n5182, n5181, n5183, n5807,
    n5187, n5184, n5186, n5909, n5190, n5189, n5195, n5193, n5914, n5192,
    n5194, n5197, n5920, n5196, n5198, n5911, n5201, n5200, n5203, n5202,
    n5206, n5204, n5910, n5205, n5208, n5207, n5213, n5271, n6322, n5211,
    n5210, n5212, n5215, n6330, n5214, n5216, n5219, n5218, n5657, n5217,
    n5220, n5697, n5737, n5222, n5221, n5735, n5223, n5270, n5225, n5226,
    n5229, n5227, n5228, n5230, n7721, n5232, n7773, n5231, n5238, n5236,
    n5234, n5233, n5235, n5237, n5254, n5240, n5239, n5244, n5242, n5241,
    n5243, n5252, n5246, n5245, n5250, n5248, n5247, n5249, n5251, n5253,
    n5259, n5256, n5255, n5257, n5258, n5260, n5261, n5672, n5262, n7780,
    n5674, n5679, n5266, n6215, n5343, n5295, n6203, n5268, n5558, n5560,
    n5269, n5288, n5309, n5299, n6301, n5277, n5273, n5272, n5275, n6295,
    n5274, n5276, n7988, n5279, n5286, n5298, n5282, n5346, n5284, n7069,
    n7059, n5307, n5285, n5287, n5453, n5451, n5290, n5450, n5291, n5292,
    n5293, n5294, n5305, n5297, n5296, n6131, n5670, n5303, n5301, n5300,
    n5302, n5304, n5306, n5308, n7124, n7035, n5311, n7029, n5310, n7047,
    n7048, n5313, n5316, n5447, n5315, n5413, n5318, n7096, n5319, n5322,
    n7125, n7143, n5324, n7153, n5325, n5328, n7182, n5330, n7210, n5332,
    n7240, n5335, n5334, n7265, n5337, n5336, n7283, n5339, n5338, n5342,
    n5340, n5341, n5347, n6213, n5396, n5344, n5397, n7018, n7058, n7067,
    n7077, n5405, n7027, n7026, n7066, n5350, n5349, n7042, n7041, n5351,
    n5355, n5354, n5356, n5359, n5358, n7093, n7094, n5361, n5360, n5362,
    n7113, n7120, n5363, n5364, n7122, n5365, n5369, n5368, n7151, n5371,
    n5370, n5373, n7176, n5374, n7204, n7205, n5379, n5378, n5382, n5380,
    n7207, n5381, n5384, n5385, n7220, n7233, n5388, n5387, n7259, n5390,
    n5389, n7273, n7274, n5391, n5394, n7275, n5828, n5398, n7270, n5399,
    n5400, n5403, n7080, n5402, n5406, n5408, n5407, n5410, n5409, n5412,
    n5411, n5415, n5414, n5418, n5417, n5421, n5420, n5423, n5422, n6209,
    n5424, n5426, n5425, n5428, n5427, n5431, n5430, n5433, n5432, n7776,
    n5435, n5434, n5437, n5436, n6826, n5438, n5446, n5440, n5444, n5442,
    n5443, n5445, n5449, n5448, n5452, n6983, n7019, n5461, n5455, n7650,
    n5454, n5459, n7061, n6970, n5458, n5460, n7957, n5463, n5462, n5465,
    n5464, n5467, n5466, n5469, n5468, n5471, n5470, n5473, n5472, n5475,
    n5474, n5477, n5476, n5479, n5478, n5481, n5480, n5483, n5482, n5485,
    n5484, n5487, n5486, n5489, n5488, n5491, n5490, n5493, n5492, n5495,
    n5494, n6133, n6137, n6141, n5497, n7582, n6140, n6147, n5499, n7557,
    n5588, n7558, n6112, n5501, n7496, n7532, n5595, n5500, n6158, n5503,
    n7495, n7473, n6113, n6159, n6157, n6120, n5504, n6118, n7339, n7344,
    n5505, n6129, n5506, n5992, n5607, n7341, n7350, n7343, n5508, n5507,
    n5510, n7367, n5509, n5993, n7310, n5997, n6597, n5999, n5998, n6740,
    n5511, n6594, n6179, n6502, n6084, n6504, n6002, n6477, n6168, n6376,
    n6398, n6070, n5625, n5513, n6111, n6387, n6381, n6167, n5514, n6010,
    n6069, n6356, n6063, n6187, n5518, n6466, n6379, n6008, n6181, n6537,
    n6531, n5898, n5633, n6503, n5515, n6083, n6478, n5516, n6436, n6005,
    n6377, n5517, n6339, n5519, n6310, n6053, n6188, n5722, n6298, n6286,
    n5520, n6280, n6191, n5724, n6264, n5529, n5523, n5522, n5527, n5524,
    n5526, n5528, n7991, n6258, n6049, n6254, n6195, n6050, n6034, n5531,
    n5530, n5540, n5534, n5533, n5536, n5684, n5789, n5538, n6248, n5537,
    n5539, n7994, n5790, n5664, n5663, n5550, n5543, n5542, n5548, n5546,
    n5545, n5547, n6030, n6052, n5553, n5552, n5551, n7678, n5566, n5555,
    n5554, n5557, n5556, n8001, n5559, n6223, n5564, n7668, n7533, n5562,
    n6022, n5561, n5563, n5565, n5687, n5569, n7641, n7570, n5571, n6582,
    n6397, n5573, n6273, n5779, n6231, n5575, n5683, n5576, n5669, n5580,
    n7683, n7685, n5579, n5582, n5583, n5585, n5584, n7591, n7592, n5587,
    n5586, n7556, n5589, n5591, n5590, n7526, n5592, n5594, n5593, n7511,
    n5597, n5596, n7478, n7502, n5598, n5599, n5600, n5601, n5603, n5605,
    n5604, n7340, n5608, n6587, n5636, n5620, n5614, n5611, n6738, n5612,
    n5616, n6736, n5613, n6735, n6590, n5617, n5634, n6458, n6460, n5644,
    n6462, n6459, n6367, n5626, n5624, n5622, n6374, n5623, n5629, n6428,
    n6373, n5627, n6371, n5628, n5649, n5632, n6370, n5631, n5648, n6334,
    n5647, n5645, n5641, n6588, n5637, n5638, n5640, n5643, n5642, n5656,
    n5652, n5651, n6461, n5650, n5654, n5653, n5655, n5658, n5917, n5659,
    n6267, n5661, n6285, n5662, n6014, n6032, n5723, n5667, n7887, n5668,
    n5768, n5671, n5673, n5675, n5767, n5676, n7952, n7954, n5678, n5677,
    n5681, n7608, n7418, n7642, n5685, n5686, n5691, n7698, n7691, n6244,
    n6528, n5690, n5693, n5692, n5694, n5710, n5696, n5695, n5709, n5739,
    n5715, n5699, n5698, n5701, n5705, n5703, n5702, n5704, n5786, n5706,
    n5717, n5707, n5708, n5714, n5712, n5738, n5711, n5716, n5713, n5719,
    n5718, n5720, n5721, n5734, n5730, n5728, n5726, n5725, n5727, n5729,
    n5732, n5731, n5733, n5740, n5751, n5749, n5747, n5745, n5743, n5742,
    n5744, n5746, n5748, n5750, n5753, n5759, n5757, n7997, n5755, n5754,
    n5756, n5758, n6243, n5760, n6240, n5763, n6245, n5762, n5771, n5765,
    n5764, n7900, n7907, n5770, n5769, n5773, n5772, n5776, n5775, n5777,
    n5783, n5781, n5780, n5782, n5787, n5784, n5785, n5788, n5803, n5800,
    n5798, n6251, n5796, n5794, n5792, n5791, n5793, n5795, n5797, n5799,
    n5801, n5806, n5805, n5809, n5821, n5810, n5819, n5812, n5811, n5814,
    n5813, n5817, n5816, n5818, n5820, n5824, n5825, n5836, n5834, n5830,
    n5827, n5829, n5832, n5831, n5833, n5835, n5838, n5928, n5842, n5841,
    n5843, n5854, n6449, n5852, n5848, n5846, n5845, n5847, n5850, n5849,
    n5851, n5853, n5857, n6847, n5858, n6938, n5861, n6935, n6808, n6809,
    n5865, n5864, n5866, n5870, n5869, n5868, n5871, n5979, n5873, n5872,
    n5874, n5876, n5886, n6613, n5884, n5878, n7245, n5880, n5879, n5882,
    n5881, n5883, n5885, n5888, n5895, n5891, n5893, n5894, n5896, n5908,
    n6574, n5906, n5899, n7257, n5901, n6567, n5900, n5904, n5903, n5905,
    n5907, n5912, n5913, n5926, n6360, n5924, n5916, n5915, n5919, n5918,
    n5922, n5921, n5923, n5925, n5930, n5931, n5942, n5932, n5940, n5934,
    n5933, n5936, n5935, n5938, n5937, n5939, n5941, n5946, n5947, n5958,
    n5948, n5956, n5950, n5949, n5952, n5951, n5954, n5953, n5955, n5957,
    n5965, n5963, n5962, n5964, n5966, n5978, n6558, n5976, n5968, n7272,
    n5971, n5970, n5974, n5973, n5975, n5977, n5981, n5991, n5982, n5989,
    n5983, n7231, n5985, n5984, n5987, n5986, n5988, n5990, n5996, n5995,
    n6124, n6000, n6127, n6125, n6001, n6004, n6169, n6003, n6006, n6173,
    n6007, n6009, n6011, n6012, n6013, n6029, n6035, n6027, n6017, n6016,
    n6019, n6018, n6224, n6225, n6043, n6197, n6232, n6021, n6064, n6024,
    n6036, n6025, n6026, n6028, n6040, n6031, n6110, n6033, n6038, n6037,
    n6198, n6039, n6042, n8006, n6233, n6041, n6046, n6062, n6044, n6060,
    n6045, n6047, n6048, n6108, n6051, n6268, n6101, n6282, n7426, n7448,
    n6058, n6312, n7479, n6055, n6132, n6054, n7787, n7703, n6056, n6057,
    n6059, n6099, n6061, n6196, n6342, n6065, n6066, n6097, n6068, n7539,
    n6067, n6072, n6340, n6382, n6071, n6095, n6076, n6075, n6081, n6077,
    n6079, n6078, n6080, n6093, n6082, n6433, n6499, n6089, n6526, n6085,
    n6565, n6087, n7347, n7375, n6086, n6088, n6091, n7614, n6090, n6092,
    n6094, n6096, n6098, n6100, n6103, n6104, n6106, n6107, n6109, n6206,
    n6193, n6185, n6115, n6114, n6155, n6116, n6117, n6119, n6122, n6128,
    n6121, n6123, n6126, n6166, n6130, n6164, n6135, n6134, n6139, n6138,
    n6143, n6142, n6146, n6145, n6150, n6148, n6149, n6154, n6151, n6153,
    n6156, n6162, n6160, n6161, n6163, n6165, n6172, n6174, n6177, n6171,
    n6176, n6175, n6183, n6178, n6180, n6182, n6184, n6186, n6189, n6190,
    n6192, n6194, n6201, n6199, n6200, n6202, n6204, n6205, n6208, n6207,
    n6222, n6210, n6211, n6212, n6214, n6219, n6217, n6218, n6220, n6221,
    n7665, n6230, n6235, n6226, n6621, n6228, n6227, n6229, n6624, n6239,
    n6234, n6625, n6237, n6236, n6238, n6241, n6242, n6247, n7513, n6246,
    n6250, n6249, n6253, n7699, n6252, n6257, n6262, n6260, n6259, n6261,
    n6263, n6265, n6266, n6270, n6632, n6269, n6272, n6271, n6277, n6274,
    n6629, n6276, n6637, n6294, n6281, n6283, n6284, n6292, n7573, n6290,
    n6288, n6287, n6289, n6291, n6293, n6642, n6297, n6296, n6307, n7613,
    n7702, n6305, n6300, n6638, n6303, n6302, n6304, n6306, n6645, n6326,
    n6311, n6313, n6314, n6321, n6319, n6317, n6316, n6318, n6320, n6648,
    n6323, n6324, n6325, n6328, n6327, n6332, n6646, n6331, n6336, n6337,
    n6653, n6353, n6341, n6343, n6344, n6351, n6349, n6347, n6346, n6348,
    n6350, n6352, n6658, n6355, n6354, n6366, n6364, n6359, n6358, n6654,
    n6362, n6361, n6363, n6365, n6369, n6432, n6372, n6393, n6378, n6434,
    n6380, n6406, n6408, n6383, n6384, n6391, n6386, n6385, n6389, n6388,
    n6390, n6392, n6666, n6395, n6394, n6405, n6403, n6422, n6662, n6401,
    n6400, n6402, n6404, n6407, n6409, n6416, n6412, n6411, n6414, n6413,
    n6415, n6672, n6418, n6417, n6427, n6420, n6421, n6670, n6425, n6424,
    n6426, n6431, n6669, n6430, n6677, n6445, n6435, n6443, n6441, n6439,
    n6438, n6440, n6442, n6444, n6682, n6447, n6446, n6455, n6453, n6678,
    n6451, n6450, n6452, n6454, n6548, n6552, n6527, n6475, n6498, n6464,
    n6463, n6473, n7648, n6465, n6472, n6468, n6467, n6470, n6469, n6471,
    n6488, n6474, n6476, n6482, n6479, n6483, n6480, n6481, n6486, n6484,
    n6485, n6487, n6686, n6490, n6685, n6491, n6492, n6494, n6493, n6497,
    n6496, n6501, n6687, n7527, n6500, n6505, n6506, n6507, n6513, n6511,
    n6509, n6508, n6510, n6512, n6695, n6515, n6514, n6525, n6520, n6519,
    n6693, n6523, n6522, n6524, n6530, n6692, n6529, n6533, n6534, n6541,
    n6536, n6535, n6539, n6538, n6540, n6701, n6544, n6700, n6545, n6546,
    n6554, n6550, n6551, n6702, n6553, n6557, n6555, n6556, n6560, n6559,
    n6563, n6564, n6707, n6578, n6566, n6573, n6571, n6569, n6568, n6570,
    n6572, n6710, n6575, n6576, n6577, n6581, n6579, n6580, n6586, n6584,
    n6708, n6585, n7329, n6592, n6593, n6715, n6606, n6596, n6604, n6602,
    n6600, n6599, n6601, n6603, n6605, n6720, n6609, n6607, n6608, n6619,
    n6617, n6612, n6716, n6615, n6614, n6616, n6618, n7883, n6623, n6622,
    n6626, n6749, n6628, n6627, n6630, n6633, n6752, n6636, n6635, n6640,
    n6639, n6641, n6755, n6644, n6643, n6650, n6647, n6649, n6758, n6652,
    n6651, n6656, n6655, n6657, n6761, n6660, n6659, n6663, n6665, n6764,
    n6668, n6667, n6674, n6671, n6673, n6767, n6676, n6675, n6680, n6679,
    n6681, n6770, n6684, n6683, n6689, n7852, n6688, n6773, n6691, n6690,
    n6697, n6694, n6696, n6776, n6699, n6698, n6704, n6703, n6779, n6706,
    n6705, n6712, n6709, n6711, n6782, n6714, n6713, n6718, n6717, n6719,
    n6785, n6722, n6721, n6724, n6731, n6727, n6726, n6729, n6728, n6730,
    n7295, n7289, n6734, n6743, n6737, n7300, n6739, n6741, n7288, n6742,
    n6788, n6745, n6744, n6748, n6747, n6751, n6750, n6754, n6753, n6757,
    n6756, n6760, n6759, n6763, n6762, n6766, n6765, n6769, n6768, n6772,
    n6771, n6775, n6774, n6778, n6777, n6781, n6780, n6784, n6783, n6787,
    n6786, n6790, n6789, n6791, n7118, n6795, n6793, n6792, n6794, n6802,
    n6797, n6800, n6799, n6801, n6803, n7219, n6807, n6805, n6804, n6806,
    n6814, n6810, n6812, n6811, n6813, n6815, n7163, n6819, n6817, n6816,
    n6818, n6825, n6821, n6823, n6822, n6824, n6827, n6831, n6829, n6828,
    n6830, n6838, n6834, n6836, n6835, n6837, n6839, n7136, n6844, n6842,
    n6841, n6843, n6853, n6848, n6849, n6851, n6850, n6852, n7669, n6856,
    n6855, n6866, n6857, n6864, n6860, n6862, n6861, n6863, n6865, n6867,
    n7191, n6871, n6869, n6868, n6870, n6888, n6877, n6874, n6883, n6876,
    n6881, n6880, n6882, n6884, n6886, n6885, n6887, n6889, n7092, n6893,
    n6891, n6890, n6892, n6903, n6896, n6897, n6899, n6901, n6900, n6902,
    n6904, n7075, n6908, n6906, n6905, n6907, n6914, n6910, n6912, n6911,
    n6913, n6916, n7147, n6929, n6918, n6920, n6925, n6923, n6922, n6924,
    n6927, n6926, n6928, n6930, n7203, n6934, n6932, n6931, n6933, n6950,
    n6936, n6945, n6940, n6943, n6942, n6944, n6946, n6948, n6947, n6949,
    n6953, n7175, n6959, n6957, n6956, n6958, n6961, n6960, n6973, n6965,
    n6969, n6968, n6971, n6972, n6978, n6976, n6975, n6977, n6987, n6981,
    n6985, n6982, n6984, n6986, n6989, n7106, n6995, n6993, n6992, n6994,
    n7013, n6996, n7006, n6999, n7004, n7003, n7005, n7008, n7011, n7010,
    n7012, n7014, n7062, n7015, n7016, n7017, n7021, n7020, n7023, n7022,
    n7025, n7024, n7033, n7028, n7031, n7030, n7032, n7038, n7036, n7037,
    n7040, n7039, n7057, n7045, n7044, n7052, n7050, n7049, n7051, n7055,
    n7054, n7056, n7073, n7060, n7065, n7063, n7064, n7072, n7068, n7070,
    n7071, n7089, n7074, n7088, n7078, n7082, n7081, n7086, n7084, n7085,
    n7087, n7090, n7091, n7102, n7095, n7100, n7098, n7099, n7101, n7104,
    n7103, n7105, n7112, n7108, n7110, n7109, n7111, n7116, n7114, n7115,
    n7117, n7132, n7121, n7123, n7130, n7127, n7128, n7129, n7131, n7134,
    n7133, n7135, n7142, n7138, n7140, n7139, n7141, n7146, n7144, n7145,
    n7149, n7148, n7159, n7152, n7157, n7155, n7156, n7158, n7161, n7160,
    n7162, n7171, n7165, n7169, n7167, n7168, n7170, n7173, n7172, n7174,
    n7189, n7178, n7180, n7179, n7187, n7185, n7184, n7186, n7188, n7190,
    n7199, n7193, n7197, n7195, n7196, n7198, n7201, n7200, n7202, n7215,
    n7206, n7208, n7213, n7211, n7212, n7214, n7217, n7216, n7218, n7227,
    n7221, n7225, n7223, n7224, n7226, n7229, n7228, n7230, n7238, n7234,
    n7236, n7235, n7237, n7243, n7241, n7242, n7244, n7251, n7247, n7249,
    n7248, n7250, n7255, n7253, n7254, n7256, n7264, n7262, n7260, n7261,
    n7263, n7269, n7267, n7268, n7271, n7281, n7276, n7279, n7278, n7280,
    n7287, n7285, n7286, n7291, n7290, n7294, n7293, n7296, n7297, n7299,
    n7298, n7902, n7301, n7304, n7302, n7904, n7303, n7307, n7306, n7325,
    n7312, n7311, n7313, n7324, n7322, n7318, n7317, n7320, n7319, n7321,
    n7323, n7906, n7326, n7328, n7327, n7893, n7349, n7335, n7331, n7333,
    n7895, n7334, n7338, n7337, n7361, n7342, n7345, n7346, n7348, n7360,
    n7358, n7356, n7354, n7353, n7355, n7357, n7359, n7897, n7362, n7364,
    n7363, n7366, n7374, n7372, n7370, n7369, n7371, n7373, n7886, n7888,
    n7384, n7378, n7380, n7382, n7884, n7383, n7385, n7386, n7389, n7388,
    n7391, n7390, n7392, n7404, n7402, n7396, n7395, n7400, n7876, n7399,
    n7401, n7403, n7880, n7875, n7406, n7409, n7408, n7410, n7412, n7411,
    n7414, n7413, n7868, n7433, n7417, n7867, n7431, n7422, n7420, n7419,
    n7421, n7425, n7423, n7424, n7430, n7428, n7429, n7872, n7432, n7434,
    n7437, n7436, n7439, n7438, n7442, n7441, n7445, n7859, n7444, n7464,
    n7860, n7462, n7449, n7458, n7456, n7454, n7453, n7455, n7457, n7460,
    n7459, n7864, n7461, n7463, n7467, n7466, n7494, n7469, n7848, n7489,
    n7485, n7483, n7540, n7475, n7476, n7477, n7481, n7851, n7480, n7482,
    n7484, n7488, n7487, n7850, n7490, n7492, n7491, n7493, n7497, n7498,
    n7500, n7499, n7501, n7510, n7508, n7506, n7505, n7507, n7509, n7841,
    n7843, n7518, n7515, n7842, n7517, n7519, n7520, n7523, n7522, n7525,
    n7524, n7833, n7528, n7531, n7836, n7530, n7550, n7538, n7536, n7535,
    n7537, n7545, n7541, n7543, n7542, n7544, n7835, n7547, n7548, n7549,
    n7552, n7551, n7555, n7554, n7581, n7559, n7826, n7569, n7561, n7567,
    n7562, n7565, n7564, n7566, n7568, n7830, n7823, n7575, n7824, n7576,
    n7577, n7579, n7578, n7580, n7588, n7586, n7585, n7587, n7596, n7590,
    n7594, n7816, n7593, n7595, n7818, n7597, n7606, n7600, n7601, n7819,
    n7604, n7603, n7605, n7607, n7610, n7609, n7808, n7627, n7616, n7626,
    n7624, n7622, n7620, n7619, n7621, n7623, n7625, n7813, n7628, n7636,
    n7809, n7631, n7630, n7634, n7633, n7635, n7638, n7637, n7644, n7639,
    n7640, n7800, n7643, n7664, n7801, n7662, n7647, n7660, n7649, n7658,
    n7656, n7654, n7653, n7655, n7657, n7659, n7805, n7661, n7663, n7795,
    n7667, n7666, n7695, n7673, n7672, n7690, n7675, n7677, n7679, n7682,
    n7681, n7688, n7686, n7792, n7687, n7689, n7794, n7692, n7693, n7694,
    n7697, n7696, n7701, n7700, n7705, n7704, n7719, n7708, n7711, n7710,
    n7786, n7713, n7715, n7716, n7717, n7718, n7779, n7724, n7725, n7727,
    n7726, n7728, n7731, n7730, n7734, n7733, n7737, n7736, n7740, n7739,
    n7743, n7742, n7746, n7745, n7749, n7748, n7752, n7751, n7755, n7754,
    n7758, n7757, n7761, n7760, n7764, n7763, n7767, n7766, n7770, n7769,
    n7772, n7771, n7775, n7778, n7781, n7777, n7783, n7782, n7791, n7785,
    n7789, n7788, n7910, n7790, n7799, n7793, n7797, n7796, n7913, n7798,
    n7807, n7803, n7802, n7804, n7916, n7806, n7815, n7811, n7810, n7812,
    n7919, n7814, n7822, n7817, n7820, n7922, n7821, n7832, n7825, n7828,
    n7827, n7829, n7925, n7831, n7840, n7834, n7838, n7837, n7928, n7839,
    n7847, n7845, n7844, n7931, n7846, n7857, n7849, n7855, n7853, n7854,
    n7934, n7856, n7866, n7862, n7861, n7863, n7937, n7865, n7874, n7870,
    n7869, n7871, n7940, n7873, n7882, n7878, n7877, n7879, n7943, n7881,
    n7892, n7885, n7890, n7889, n7946, n7891, n7899, n7894, n7896, n7949,
    n7898, n7909, n7903, n7905, n7953, n7908, n7912, n7911, n7915, n7914,
    n7918, n7917, n7921, n7920, n7924, n7923, n7927, n7926, n7930, n7929,
    n7933, n7932, n7936, n7935, n7939, n7938, n7942, n7941, n7945, n7944,
    n7948, n7947, n7951, n7950, n7956, n7955, n7960, n7959, n7963, n7962,
    n7966, n7965, n7969, n7968, n7972, n7971, n7975, n7974, n7978, n7977,
    n7981, n7980, n7984, n7983, n7987, n7986, n7990, n7989, n7993, n7992,
    n7996, n7995, n7999, n7998, n8004, n8002, n8003, n8008, n8007, n5752;
  assign n4545 = n6309 | n4547;
  assign n6589 = n7376 | n6587;
  assign n5348 = n4726 ^ ~n4725;
  assign n5994 = ~n6725 | ~n7315;
  assign n6725 = ~n7351;
  assign n7684 = ~n6136 | ~n6133;
  assign n7574 = ~n7503;
  assign n4360 = ~n4771;
  assign n6898 = n4715 ^ ~n4716;
  assign n5456 = ~n4748 | ~n4747;
  assign n7516 = ~n4664 | ~n4667;
  assign n7712 = ~n7516;
  assign n4948 = n4920 | n4849;
  assign n4920 = ~n4918 | ~n4848;
  assign n4716 = ~n4696 | ~n4695;
  assign n7680 = ~n4766 | ~n4765;
  assign n7164 = n5372 ^ ~n5326;
  assign n5372 = ~n5371 | ~n5370;
  assign n5188 = ~n5153;
  assign n4620 = n4614 ^ ~n4615;
  assign n4614 = n4616 | n4767;
  assign n4358 = n5312;
  assign n4759 = n6858 | n6859;
  assign n7979 = ~n6345;
  assign n7309 = n5994 & n5997;
  assign n7486 = ~n4817 | ~n4816;
  assign n5700 = ~n4711;
  assign n4730 = ~n5774;
  assign n7618 = ~n4513 | ~n4791;
  assign n5544 = ~n4760;
  assign n4359 = ~n4682;
  assign n5804 = ~n5714 | ~n5713;
  assign n6661 = n4457 ^ ~n4456;
  assign n4589 = n5687 | n5686;
  assign n7282 = ~n5337 & ~n5336;
  assign n5808 = ~n4566 | ~n4567;
  assign n6368 = n6333 & n4590;
  assign n7252 = n7735 ^ ~n5333;
  assign n5646 = n4590 & n5645;
  assign n6457 = n6547 & n4418;
  assign n6547 = n5643 & n5642;
  assign n6456 = n6561 | n5634;
  assign n4991 = ~n5859 & ~n4990;
  assign n6561 = n6587 | n5639;
  assign n5859 = n6937 | n4386;
  assign n5327 = ~n4498 | ~n4497;
  assign n4541 = n4543 & n4382;
  assign n4543 = n5503 | n7473;
  assign n7612 = n4460 & n5582;
  assign n6859 = n4755 & n4754;
  assign n6967 = n4912 | n4911;
  assign n6345 = n5176 & n5175;
  assign n6144 = ~n7582 | ~n7618;
  assign n5778 = n4907;
  assign n7617 = ~n4702 | ~n4701;
  assign n7314 = ~n4953 | ~n4952;
  assign n7351 = ~n4970 | ~n4969;
  assign n7394 = ~n4853 | ~n4852;
  assign n7583 = ~n4686 | ~n4685;
  assign n7316 = ~n5001 | ~n5000;
  assign n7651 = ~n4788 | ~n4787;
  assign n4711 = ~n5688 | ~n5278;
  assign n4816 = n4815 & n4814;
  assign n7572 = n7858 | n7712;
  assign n5496 = ~n4442 | ~n4439;
  assign n6854 = ~n4363 | ~n4374;
  assign n7858 = n5267 | n7784;
  assign n5688 = n5267 | n6105;
  assign n4442 = n4724 & n4443;
  assign n6015 = n4894;
  assign n5267 = n4631 ^ ~IR_REG_20__SCAN_IN;
  assign n4891 = ~n4621 & ~n4461;
  assign n4617 = ~n7722 | ~IR_REG_31__SCAN_IN;
  assign n5441 = n5314 ^ ~n5352;
  assign n4616 = n4613 & n4551;
  assign n5314 = ~n7048 | ~n5313;
  assign n4637 = n4645 & n4632;
  assign n4965 = ~n4948 & ~n4947;
  assign n4613 = n4647 & n4607;
  assign n5312 = n4770 ^ ~n4769;
  assign n4855 = ~IR_REG_6__SCAN_IN & ~IR_REG_7__SCAN_IN;
  assign n4768 = ~IR_REG_0__SCAN_IN & ~IR_REG_1__SCAN_IN;
  assign n4769 = ~IR_REG_2__SCAN_IN;
  assign n4600 = ~IR_REG_16__SCAN_IN & ~IR_REG_20__SCAN_IN;
  assign n4789 = ~IR_REG_3__SCAN_IN;
  assign n4601 = ~IR_REG_18__SCAN_IN & ~IR_REG_17__SCAN_IN;
  assign n5689 = n6052 ^ n5665;
  assign n5665 = n4414 & n4369;
  assign n4361 = ~IR_REG_31__SCAN_IN;
  assign n4362 = n4651 & n4743;
  assign n5172 = n5151 & REG3_REG_21__SCAN_IN;
  assign n4918 = ~n4812 & ~n4811;
  assign n4812 = ~n4622 | ~REG3_REG_4__SCAN_IN;
  assign n5635 = ~n4411 | ~n6595;
  assign n5502 = n7474 & n6158;
  assign n5329 = ~n4484 | ~n4483;
  assign n4484 = ~n7166 | ~n4481;
  assign n4483 = n4479 & n4387;
  assign n4481 = ~n4485 & ~n4482;
  assign n5639 = ~n5620 & ~n5619;
  assign n5619 = n5618 | n5617;
  assign n4516 = ~n5571 | ~n5602;
  assign n4448 = n4449 & n5600;
  assign n4449 = ~n4450 | ~n5599;
  assign n4450 = ~n5598;
  assign n4582 = ~n5961;
  assign n4715 = n4694 ^ ~n5700;
  assign n4694 = ~n4693 | ~n4692;
  assign n4757 = n4733 ^ ~n4711;
  assign n7194 = n5329 ^ ~n5376;
  assign n4540 = n7275 & n4396;
  assign n6136 = n5496 | n7670;
  assign n7599 = n4708 & n4707;
  assign n7598 = ~n7641 & ~n7618;
  assign n7571 = ~n7563;
  assign n7534 = ~n7529;
  assign n7901 = n5296 | n5267;
  assign n4404 = ~n4405 | ~n4408;
  assign n7474 = n5501 | n5500;
  assign n4558 = n4845 & n7002;
  assign n4497 = n4494 & n5325;
  assign n4519 = ~REG2_REG_10__SCAN_IN;
  assign n5606 = n4906 & n6954;
  assign n4544 = n4546 & n6050;
  assign n4406 = ~n4407 | ~n5656;
  assign n4554 = n5511 & n5994;
  assign n7560 = ~n4426 | ~n6147;
  assign n4426 = ~n4424 | ~n4421;
  assign n4421 = n4422 & n4555;
  assign n5280 = n4654 & IR_REG_31__SCAN_IN;
  assign n4672 = n4639 | IR_REG_22__SCAN_IN;
  assign n5862 = n4992 | n4993;
  assign n4569 = ~n5145 & ~n5169;
  assign n4583 = ~n5823;
  assign n5021 = n4915 | n4914;
  assign n7563 = n4691 & n4690;
  assign n5071 = n5069 & n5068;
  assign n5018 = n4905 ^ ~n4711;
  assign n5020 = n4884 ^ ~n5700;
  assign n4654 = ~n4613 | ~n4517;
  assign n4517 = n4645 & n4553;
  assign n5959 = ~n5887 & ~n5892;
  assign n5353 = ~n7041 | ~n5351;
  assign n5367 = ~n4525 | ~n4523;
  assign n4523 = ~n4524 | ~n5365;
  assign n4524 = ~n7120 | ~n5363;
  assign n7166 = n5327 ^ ~n5326;
  assign n5331 = ~n4474 | ~n4472;
  assign n4472 = ~n4473 & ~n4392;
  assign n4475 = ~n4477 & ~n4476;
  assign n5386 = ~n4531 | ~n4529;
  assign n5393 = n7516 ^ ~n5392;
  assign n4507 = n4508 | n6286;
  assign n6102 = n6014 & n6032;
  assign n4508 = n6356 | n5657;
  assign n6357 = ~n6396 | ~n5573;
  assign n6396 = n6516 & n6489;
  assign n6516 = ~n6582 & ~n4511;
  assign n4511 = ~n4365 | ~n5826;
  assign n4512 = ~n6582;
  assign n6562 = n5639 | n5638;
  assign n7379 = n4865 & n4864;
  assign n7376 = ~n4453 | ~n5608;
  assign n4453 = ~n5605 | ~n4454;
  assign n4454 = ~n7398 & ~n4455;
  assign n7427 = ~n4436 | ~n6157;
  assign n7415 = ~n4446 | ~n4444;
  assign n4444 = n4445 & n5601;
  assign n7470 = ~n6840;
  assign n7529 = n4661 & n4660;
  assign n7629 = ~n7618;
  assign n7645 = ~n7685 | ~n5579;
  assign n7670 = n4728 & n4727;
  assign n5263 = ~n4672 | ~IR_REG_31__SCAN_IN;
  assign n4574 = ~n4364 & ~IR_REG_18__SCAN_IN;
  assign n4665 = ~IR_REG_19__SCAN_IN;
  assign n7315 = ~n5610;
  assign n4584 = ~n5960;
  assign n4581 = ~n4582 | ~n5892;
  assign n4570 = ~n5944 & ~n4571;
  assign n4571 = ~n5148;
  assign n4572 = ~n5147 | ~n5146;
  assign n6990 = ~n6974;
  assign n4562 = n4565 & n5205;
  assign n4565 = ~n5735;
  assign n4651 = ~n5688;
  assign n6023 = n5548 & n5547;
  assign n4413 = ~n6015 | ~REG1_REG_16__SCAN_IN;
  assign n7043 = n4358 ^ ~REG2_REG_2__SCAN_IN;
  assign n7137 = n5367 ^ ~n5366;
  assign n7222 = n5331 ^ ~n5383;
  assign n7246 = n5386 ^ ~n7735;
  assign n5333 = ~n4491 | ~n4489;
  assign n4491 = ~n7222 | ~n4487;
  assign n4489 = ~n4490 & ~n4393;
  assign n4487 = ~n4492 & ~n4488;
  assign n7671 = n6203 | n7784;
  assign n4417 = ~n6267 | ~n5661;
  assign n4415 = ~n6102 & ~n4416;
  assign n4416 = ~n5662;
  assign n6429 = n6372 & n6371;
  assign n7398 = n7341 & n7340;
  assign n4500 = ~n7504 & ~n7471;
  assign n4428 = n4430 | n7706;
  assign n4430 = ~n6257 & ~n6256;
  assign n6256 = ~n4545 | ~n4546;
  assign n7720 = ~n5343;
  assign n4551 = n4645 & n4550;
  assign n4550 = n4552 & n4553;
  assign n4552 = ~n4652;
  assign n6664 = n6661 | n7901;
  assign n6074 = ~n7684;
  assign n6073 = ~n6595;
  assign n4482 = ~REG1_REG_10__SCAN_IN;
  assign n4532 = ~n7233;
  assign n4438 = ~n6594 | ~n6073;
  assign n4423 = ~n6137;
  assign n4468 = ~REG1_REG_4__SCAN_IN;
  assign n4477 = ~n7210;
  assign n4476 = ~REG1_REG_12__SCAN_IN;
  assign n4473 = ~n5330 & ~n4477;
  assign n4527 = ~n4532 & ~n4528;
  assign n4528 = ~REG2_REG_14__SCAN_IN;
  assign n4549 = ~n4434 | ~n4433;
  assign n4433 = ~n6188;
  assign n4434 = ~n6309;
  assign n4548 = ~n6191;
  assign n4402 = ~n4404;
  assign n4400 = ~n4401 & ~n4368;
  assign n4401 = ~n4404 & ~n5658;
  assign n4590 = ~n4420 | ~n4419;
  assign n4419 = ~n5644;
  assign n4420 = ~n6457;
  assign n4452 = ~n7376;
  assign n4418 = ~n6549;
  assign n4455 = ~n5604;
  assign n4445 = ~n4448 | ~n4451;
  assign n4542 = ~n7472 | ~n4367;
  assign n5610 = n4974 & n4973;
  assign n5863 = n4995 | n4994;
  assign n5151 = n5133 & REG3_REG_20__SCAN_IN;
  assign n6878 = n4915 & n4914;
  assign n5076 = n5055 & REG3_REG_16__SCAN_IN;
  assign n5051 = n5043 | n5044;
  assign n4557 = ~n6997 | ~n4558;
  assign n6939 = ~n4373 | ~n4595;
  assign n6820 = n4937 | n4938;
  assign n6919 = n6938 | n6917;
  assign n5091 = n5090 & n5089;
  assign n7046 = ~n5311 | ~n5310;
  assign n5317 = ~n5316 | ~n5315;
  assign n5357 = ~n5355 | ~n5354;
  assign n4462 = ~n7107 | ~REG1_REG_6__SCAN_IN;
  assign n5323 = n4466 & n4465;
  assign n4465 = ~n7125;
  assign n4466 = ~n4463 | ~n4462;
  assign n4463 = n5322 & n4464;
  assign n5377 = ~n5375 | ~n5374;
  assign n4492 = ~n7240;
  assign n4488 = ~REG1_REG_14__SCAN_IN;
  assign n4490 = ~n5332 & ~n4492;
  assign n5521 = ~n5271 & ~n5299;
  assign n5191 = n5172 & REG3_REG_22__SCAN_IN;
  assign n5095 = n5076 & REG3_REG_17__SCAN_IN;
  assign n7365 = n7342 & n7341;
  assign n6921 = n4930 & n4929;
  assign n4435 = n6133 & n7674;
  assign n5574 = ~n6275 & ~n5779;
  assign n5541 = ~n5752 & ~n5664;
  assign n6255 = n4432 & n4431;
  assign n4431 = ~n6254;
  assign n4432 = ~n4549 | ~n4548;
  assign n4547 = n6034 | n6188;
  assign n4546 = n4548 | n6034;
  assign n4399 = ~n5655 & ~n4408;
  assign n6335 = n5651 | n5650;
  assign n6591 = ~n4412 | ~n5616;
  assign n6595 = ~n4410 | ~n4409;
  assign n4409 = ~n6179;
  assign n6611 = ~n6733 & ~n5609;
  assign n6733 = ~n5572 | ~n5610;
  assign n5572 = ~n7332;
  assign n7332 = ~n4514 | ~n4515;
  assign n4515 = ~n4516 & ~n7352;
  assign n4514 = ~n7416;
  assign n7381 = ~n7416 & ~n4516;
  assign n7416 = ~n5570 | ~n6921;
  assign n5570 = ~n7443;
  assign n7674 = ~n6854 & ~n5568;
  assign n4553 = ~IR_REG_26__SCAN_IN;
  assign n5283 = ~IR_REG_28__SCAN_IN;
  assign n4609 = ~IR_REG_5__SCAN_IN & ~IR_REG_10__SCAN_IN;
  assign n4610 = ~IR_REG_12__SCAN_IN & ~IR_REG_8__SCAN_IN;
  assign n4611 = ~IR_REG_11__SCAN_IN & ~IR_REG_9__SCAN_IN;
  assign n4705 = ~IR_REG_4__SCAN_IN;
  assign n5532 = n5521 & REG3_REG_26__SCAN_IN;
  assign n4567 = ~n4568 | ~n5168;
  assign n4568 = ~n4570;
  assign n4513 = ~n6020 | ~DATAI_3_;
  assign n4561 = ~n4758;
  assign n5114 = ~n5095 | ~REG3_REG_18__SCAN_IN;
  assign n4578 = ~n4580 | ~n4583;
  assign n4577 = ~n5887 | ~n4582;
  assign n6846 = n4986 | n4985;
  assign n6845 = n4983 | n4984;
  assign n6610 = n5037 & n5036;
  assign n5892 = ~n5073 & ~n5072;
  assign n6954 = n4902 & n4901;
  assign n6963 = n6919 & n6820;
  assign n5960 = n5092 & n5091;
  assign n6732 = n5006 & n5005;
  assign n5155 = n5544 | n6423;
  assign n4877 = n4873 & n4872;
  assign n5439 = n5353 ^ ~n5352;
  assign n7083 = n5357 ^ ~n5413;
  assign n7076 = n5317 ^ ~n7079;
  assign n7107 = n5321 ^ ~n4659;
  assign n7150 = ~n5369 | ~n5368;
  assign n4486 = ~n7166 | ~REG1_REG_10__SCAN_IN;
  assign n7192 = n5377 ^ ~n5376;
  assign n4478 = ~n7194 | ~REG1_REG_12__SCAN_IN;
  assign n4533 = ~n7220 | ~REG2_REG_14__SCAN_IN;
  assign n7258 = ~n5388 & ~n5387;
  assign n4537 = ~n4540 | ~n4395;
  assign n4536 = n7274 & n4539;
  assign n4539 = ~n5393;
  assign n6275 = n6357 | n4505;
  assign n4505 = ~n4506 | ~n6258;
  assign n4506 = ~n4507;
  assign n6631 = ~n4428 | ~n4429;
  assign n5133 = ~n5114 & ~n5395;
  assign n6723 = ~n7308 | ~n5994;
  assign n4502 = ~n4503 | ~n7514;
  assign n4811 = ~REG3_REG_7__SCAN_IN | ~REG3_REG_6__SCAN_IN;
  assign n4622 = REG3_REG_3__SCAN_IN & REG3_REG_5__SCAN_IN;
  assign n7646 = ~n7676 | ~n6136;
  assign n7709 = n7069 & n5558;
  assign n6299 = ~n6357 & ~n4508;
  assign n4456 = ~n6382;
  assign n4457 = ~n4458 | ~n6374;
  assign n4458 = ~n6429 | ~n6373;
  assign n6518 = ~n4512 | ~n4365;
  assign n4504 = ~n4503;
  assign n4587 = n7570 | n7571;
  assign n4607 = ~IR_REG_25__SCAN_IN;
  assign n4642 = ~n5265 | ~IR_REG_31__SCAN_IN;
  assign n5264 = ~n5263;
  assign n4770 = n4768 | n4361;
  assign n4725 = ~IR_REG_1__SCAN_IN;
  assign n4726 = ~IR_REG_31__SCAN_IN | ~IR_REG_0__SCAN_IN;
  assign n5802 = ~n5804 & ~n5785;
  assign n6991 = ~n6951;
  assign n5945 = ~n4572 | ~n5148;
  assign n6974 = n5297 & n7632;
  assign n6979 = ~n4759 | ~n4758;
  assign n6951 = n5298 | n7059;
  assign n5741 = n4563 ^ ~n4388;
  assign n4563 = ~n4564 | ~n5697;
  assign n7007 = n5295 | n5288;
  assign n7958 = ~n5031 | ~n4376;
  assign n5031 = n5028 & n5027;
  assign n6840 = ~n4925 | ~n4924;
  assign n7451 = ~n4833 | ~n4832;
  assign n4817 = n4808 & n4807;
  assign n4686 = n4681 & n4680;
  assign n4701 = n4700 & n4699;
  assign n4787 = n4786 & n4785;
  assign n4439 = n4441 & n4440;
  assign n7034 = n5348 ^ ~REG1_REG_1__SCAN_IN;
  assign n4493 = ~n7222 | ~REG1_REG_14__SCAN_IN;
  assign n7266 = ~n5335 & ~n5334;
  assign n6620 = n4510 ^ ~n6043;
  assign n4510 = ~n6231 & ~n6232;
  assign n7397 = ~n5605 | ~n5604;
  assign n7632 = ~n5670 | ~n7720;
  assign n6746 = ~n4509 | ~n6621;
  assign n4509 = ~n6620 | ~n7883;
  assign n6634 = n4428 & n4427;
  assign n4427 = ~n6630 & ~n6263;
  assign n4631 = ~n4664 | ~IR_REG_31__SCAN_IN;
  assign n5061 = ~n4971 & ~n4630;
  assign n7747 = n4863 ^ ~IR_REG_12__SCAN_IN;
  assign n7750 = n4900 ^ ~IR_REG_11__SCAN_IN;
  assign n7753 = n4879 ^ ~IR_REG_10__SCAN_IN;
  assign n7768 = n4688 ^ ~IR_REG_5__SCAN_IN;
  assign n7053 = ~n4358;
  assign n5404 = n5403 & n5402;
  assign n4767 = ~IR_REG_31__SCAN_IN;
  assign n7504 = ~n7514;
  assign n6542 = ~n4512 | ~n5902;
  assign n4363 = n4737 & n4736;
  assign n4364 = n4630 | IR_REG_17__SCAN_IN;
  assign n4365 = n5972 & n5902;
  assign n4503 = ~n7534 & ~n7571;
  assign n4886 = ~n4881 | ~n4880;
  assign n5153 = ~n4890;
  assign n5577 = n6137 & n6141;
  assign n5567 = n4773 & n4772;
  assign n5855 = n6997 & n7002;
  assign n4366 = n6357 | n4507;
  assign n4367 = n5502 & n7558;
  assign n7446 = ~n4447 | ~n5599;
  assign n4368 = n7988 & n6286;
  assign n4632 = ~n4603 & ~n4602;
  assign n5943 = n4572 & n4570;
  assign n5602 = ~n4886;
  assign n5321 = ~n5320 | ~n5319;
  assign n4647 = n4632 & n4606;
  assign n5860 = n6939 | n4386;
  assign n4369 = n5723 | n5790;
  assign n4628 = ~IR_REG_14__SCAN_IN & ~IR_REG_15__SCAN_IN;
  assign n4370 = n5959 | n5961;
  assign n4371 = n4467 & n7096;
  assign n4372 = ~n5016 | ~n5015;
  assign n4373 = n6873 | n6879;
  assign n4374 = n4739 & n4738;
  assign n4375 = n4398 & n4400;
  assign n7468 = n4839 & n4838;
  assign n4376 = n5030 & n4413;
  assign n4377 = n7617 | n7599;
  assign n4378 = n5917 & n6330;
  assign n6309 = n6338 & n5519;
  assign n4579 = ~n4580;
  assign n4580 = ~n4581 | ~n4584;
  assign n4379 = n4518 & n7176;
  assign n4380 = n4577 & n4579;
  assign n4381 = ~n6456 & ~n5644;
  assign n4382 = n6113 & n6159;
  assign n4383 = ~n6376 & ~n6010;
  assign n4384 = n4582 & n4583;
  assign U3222 = n5309 | n5308;
  assign n5224 = n4642 ^ ~n4641;
  assign n7377 = ~n7416 & ~n4886;
  assign n6170 = n7958 & n6610;
  assign n4410 = ~n6170;
  assign n5972 = n5085 & n5084;
  assign n5265 = ~n5263 | ~n4640;
  assign n4386 = ~n5014 & ~n5013;
  assign n4387 = ~REG1_REG_11__SCAN_IN | ~n7750;
  assign n7330 = n4957 & n4956;
  assign n7352 = ~n7330;
  assign n6517 = ~n5826;
  assign n4429 = ~n6263;
  assign n4485 = ~n7182;
  assign n4388 = n5740 & n5739;
  assign n4389 = n4540 & n7274;
  assign n4390 = ~n7570 & ~n4504;
  assign n4391 = n4543 & n6113;
  assign n7443 = n4501 | n7570;
  assign n4392 = REG1_REG_13__SCAN_IN & n7744;
  assign n4393 = REG1_REG_15__SCAN_IN & n7738;
  assign n5345 = ~n5280 | ~IR_REG_27__SCAN_IN;
  assign n7676 = ~n4435 | ~n6136;
  assign n4394 = REG2_REG_15__SCAN_IN & n7738;
  assign n4395 = ~n5391 | ~n5393;
  assign n7514 = n4822 & n4821;
  assign n4396 = n5391 | n5393;
  assign n4397 = ~n4502 & ~n7570;
  assign U3149 = ~STATE_REG_SCAN_IN;
  assign n4398 = ~n5655 | ~n4402;
  assign n4407 = ~n4399 & ~n4378;
  assign n6278 = ~n4403 | ~n4407;
  assign n4403 = n5656 | n4408;
  assign n5660 = ~n4406 | ~n4375;
  assign n4405 = ~n4378;
  assign n6308 = ~n5656 | ~n5655;
  assign n4408 = ~n5658;
  assign n5618 = ~n5635;
  assign n4411 = ~n6591;
  assign n4412 = ~n5615 | ~n5614;
  assign n5525 = ~n6015;
  assign n5761 = ~n4417 | ~n5662;
  assign n4414 = ~n4417 | ~n4415;
  assign n4422 = ~n7611 | ~n4423;
  assign n4424 = ~n4425 | ~n7611;
  assign n4425 = ~n5497;
  assign n4556 = ~n7615 | ~n7611;
  assign n7615 = ~n5497 | ~n6137;
  assign n4436 = ~n4542 | ~n4541;
  assign n7472 = ~n5499 | ~n5498;
  assign n5512 = ~n7308 | ~n4554;
  assign n7308 = ~n7310 | ~n7309;
  assign n6338 = ~n4438 | ~n4437;
  assign n6375 = ~n4438 | ~n4410;
  assign n4437 = n4383 & n4410;
  assign n4440 = ~n4891 | ~REG2_REG_1__SCAN_IN;
  assign n4441 = ~n4890 | ~REG0_REG_1__SCAN_IN;
  assign n4443 = ~n4894 | ~REG1_REG_1__SCAN_IN;
  assign n4446 = ~n7478 | ~n4448;
  assign n4447 = ~n7478 | ~n5598;
  assign n4451 = ~n5599;
  assign n6333 = ~n4452 | ~n4381;
  assign n4460 = ~n4459 | ~n5580;
  assign n4459 = ~n7645;
  assign n5429 = ~n4621;
  assign n4461 = ~n4620;
  assign n7126 = ~n4462 | ~n5322;
  assign n4464 = ~n7124;
  assign n5320 = ~n4469 | ~n4371;
  assign n4467 = ~n5318 | ~n4468;
  assign n4469 = ~n4470 | ~n5318;
  assign n4470 = ~n7076;
  assign n7097 = ~n4471 | ~n5318;
  assign n4471 = ~n7076 | ~REG1_REG_4__SCAN_IN;
  assign n4474 = ~n7194 | ~n4475;
  assign n7209 = ~n4478 | ~n5330;
  assign n4480 = ~n5328;
  assign n4479 = ~n4480 | ~n7182;
  assign n7183 = ~n7181 | ~n7182;
  assign n7181 = ~n4486 | ~n5328;
  assign n7239 = ~n4493 | ~n5332;
  assign n4494 = ~n4495 | ~n7153;
  assign n4495 = ~n5324;
  assign n4499 = ~n7143 | ~REG1_REG_8__SCAN_IN;
  assign n4498 = ~n7143 | ~n4496;
  assign n4496 = n7153 & REG1_REG_8__SCAN_IN;
  assign n7154 = ~n4499 | ~n5324;
  assign n7976 = ~n5157 | ~n5156;
  assign n5615 = ~n7309 & ~n5613;
  assign n4501 = ~n4503 | ~n4500;
  assign n6329 = ~n6357 & ~n6356;
  assign n5375 = ~n4520 | ~n4379;
  assign n4518 = ~n5373 | ~n4519;
  assign n4520 = ~n4521 | ~n5373;
  assign n4521 = ~n7164;
  assign n7177 = ~n4522 | ~n5373;
  assign n4522 = ~n7164 | ~REG2_REG_10__SCAN_IN;
  assign n7119 = ~n7113 | ~REG2_REG_6__SCAN_IN;
  assign n4525 = ~n7113 | ~n4526;
  assign n4526 = n5365 & REG2_REG_6__SCAN_IN;
  assign n4531 = ~n7220 | ~n4527;
  assign n7232 = ~n4533 | ~n5385;
  assign n4529 = ~n4530 & ~n4394;
  assign n4530 = ~n5385 & ~n4532;
  assign n5401 = ~n4538 | ~n4534;
  assign n4534 = ~n4535 | ~n4537;
  assign n4535 = ~n7273 | ~n4389;
  assign n4538 = ~n7273 | ~n4536;
  assign n7447 = n4542 & n4391;
  assign n6279 = ~n4549;
  assign n4643 = ~n4613 | ~n4645;
  assign n7589 = ~n4556 | ~n6144;
  assign n4555 = n4377 & n6144;
  assign n5026 = ~n4991 | ~n4557;
  assign n6997 = ~n6998 | ~n4586;
  assign n6832 = ~n4559 | ~n4782;
  assign n4559 = ~n4560 | ~n4759;
  assign n4560 = ~n6980 & ~n4561;
  assign n4801 = ~n6832 | ~n6833;
  assign n5736 = ~n5206 | ~n5205;
  assign n4564 = ~n5206 | ~n4562;
  assign n4566 = ~n5147 | ~n4569;
  assign n4666 = ~n4573 | ~IR_REG_31__SCAN_IN;
  assign n4573 = ~n4575 | ~n4574;
  assign n4575 = ~n4971;
  assign n5082 = ~n4971 & ~n4364;
  assign n4576 = ~n5887 | ~n4384;
  assign n5822 = ~n4576 | ~n4578;
  assign n7611 = n6144 & n6140;
  assign n4657 = ~n4608 | ~n4592;
  assign n4687 = n4657;
  assign n4894 = n4461 & n4621;
  assign n4890 = n4620 & n4621;
  assign n4585 = n4743 | n4751;
  assign n4586 = ~n4720 & ~n7000;
  assign n4588 = n7632 | n5684;
  assign n8005 = n8000;
  assign n4591 = n4611 & n4610;
  assign n4592 = n4789 & n4705;
  assign n4593 = ~n4893 | ~n4892;
  assign n4594 = n4894 & REG1_REG_11__SCAN_IN;
  assign n6549 = n5633 & n6504;
  assign n4595 = ~n6820 | ~n5022;
  assign n4596 = n5685 & n4588;
  assign n7452 = ~n6921;
  assign n5498 = ~n7557;
  assign n4597 = n7608 | REG2_REG_29__SCAN_IN;
  assign n6583 = ~n5902;
  assign n5902 = n5064 & n5063;
  assign n4598 = n4855 & n4609;
  assign n5630 = n5624 | n5623;
  assign n5025 = ~n4372 & ~n5024;
  assign n5376 = ~n7747;
  assign n6532 = n6375 | n6502;
  assign n6875 = ~n4913 | ~n6967;
  assign n4903 = n5774 | n6954;
  assign n6152 = ~n7512;
  assign n5549 = ~n6052;
  assign n4993 = n4979 & n4978;
  assign n4754 = n4753 | n4711;
  assign n5890 = n5070 | n5071;
  assign n5013 = n4962 & n4961;
  assign n7002 = n4806 | n4805;
  assign n4873 = ~n4760 | ~n4871;
  assign n5366 = ~n7759;
  assign n5383 = ~n7741;
  assign n5392 = ~REG2_REG_19__SCAN_IN;
  assign n6543 = ~n5972;
  assign n4627 = ~IR_REG_13__SCAN_IN;
  assign n6879 = ~n5021;
  assign n5209 = n5191 & REG3_REG_23__SCAN_IN;
  assign n6941 = n5014 & n5013;
  assign n7450 = ~n7393;
  assign n5609 = ~n6732;
  assign n5535 = n5532 & REG3_REG_27__SCAN_IN;
  assign n5826 = n5101 & n5100;
  assign n4848 = REG3_REG_9__SCAN_IN & REG3_REG_8__SCAN_IN;
  assign n7714 = ~n7671;
  assign n7512 = n5595 & n6112;
  assign n7706 = ~n7678;
  assign n5581 = ~n7680;
  assign n7368 = ~n7379;
  assign n5680 = n5450 & n7720;
  assign n6966 = n5018 | n5017;
  assign n6988 = ~n6955;
  assign n5289 = n5766 & n5679;
  assign n4681 = n5544 | n7553;
  assign n7707 = n5667 | n7712;
  assign n4878 = ~n4859 | ~n4858;
  assign n6955 = n5298 | n7069;
  assign n7009 = ~n6798;
  assign n6798 = n5453 | n5294;
  assign n6315 = n5195 & n5194;
  assign n5969 = n5099 & n5098;
  assign n5682 = n5766 | n5681;
  assign n5766 = n5232 & n5231;
  assign n7985 = n5213 | n5212;
  assign n7982 = ~n6315;
  assign n7393 = n4885;
  assign n7277 = ~n7080;
  assign n7284 = ~n7077;
  assign n8000 = n4743 | n5406;
  assign n7774 = n6215 & STATE_REG_SCAN_IN;
  assign n4599 = ~IR_REG_19__SCAN_IN & ~IR_REG_13__SCAN_IN;
  assign n4603 = ~n4628 | ~n4599;
  assign n4602 = ~n4601 | ~n4600;
  assign n4605 = ~IR_REG_23__SCAN_IN & ~IR_REG_22__SCAN_IN;
  assign n4604 = ~IR_REG_24__SCAN_IN & ~IR_REG_21__SCAN_IN;
  assign n4606 = n4605 & n4604;
  assign n4703 = ~n4768 | ~n4769;
  assign n4608 = ~n4703;
  assign n4612 = ~n4598 | ~n4591;
  assign n4645 = ~n4657 & ~n4612;
  assign n5281 = ~IR_REG_27__SCAN_IN;
  assign n4652 = ~n5281 | ~n5283;
  assign n4615 = ~IR_REG_29__SCAN_IN;
  assign n7722 = ~n4616 | ~n4615;
  assign n7723 = ~IR_REG_30__SCAN_IN;
  assign n4621 = n4617 ^ ~n7723;
  assign n4619 = ~n5188 | ~REG0_REG_6__SCAN_IN;
  assign n4682 = ~n4891;
  assign n4618 = ~n4359 | ~REG2_REG_6__SCAN_IN;
  assign n4626 = n4619 & n4618;
  assign n4624 = ~n6015 | ~REG1_REG_6__SCAN_IN;
  assign n4760 = ~n4621 & ~n4620;
  assign n4809 = ~REG3_REG_6__SCAN_IN;
  assign n7546 = n4812 ^ ~n4809;
  assign n4623 = n5544 | n7546;
  assign n4625 = n4624 & n4623;
  assign n7503 = ~n4626 | ~n4625;
  assign n4971 = ~n4645 | ~n4627;
  assign n4629 = ~IR_REG_16__SCAN_IN;
  assign n4630 = ~n4628 | ~n4629;
  assign n4664 = ~n4666 | ~n4665;
  assign n4633 = n4637 | n4767;
  assign n4635 = ~n4633 | ~IR_REG_21__SCAN_IN;
  assign n4636 = ~IR_REG_21__SCAN_IN;
  assign n4634 = ~n4636 | ~IR_REG_31__SCAN_IN;
  assign n4638 = ~n4635 | ~n4634;
  assign n4639 = ~n4637 | ~n4636;
  assign n6105 = ~n4638 | ~n4639;
  assign n4640 = ~IR_REG_23__SCAN_IN;
  assign n4641 = ~IR_REG_24__SCAN_IN;
  assign n4644 = ~n4643 | ~IR_REG_31__SCAN_IN;
  assign n5419 = n4644 ^ ~IR_REG_26__SCAN_IN;
  assign n4646 = n4645;
  assign n4648 = ~n4646 | ~n4647;
  assign n4649 = ~n4648 | ~IR_REG_31__SCAN_IN;
  assign n5416 = n4649 ^ ~IR_REG_25__SCAN_IN;
  assign n4650 = ~n5419 | ~n5416;
  assign n4743 = n5224 | n4650;
  assign n4934 = n4651 & n4743;
  assign n4663 = ~n7503 | ~n4362;
  assign n5774 = ~n5688 | ~n4743;
  assign n4656 = ~n5345 | ~n4652;
  assign n4653 = ~n4767 & ~IR_REG_28__SCAN_IN;
  assign n4655 = ~n4654 | ~n4653;
  assign n4771 = ~n4656 | ~n4655;
  assign n4857 = ~n4687 & ~IR_REG_5__SCAN_IN;
  assign n4658 = n4857 | n4767;
  assign n7765 = n4658 ^ ~IR_REG_6__SCAN_IN;
  assign n4659 = ~n7765;
  assign n4661 = n4771 | n4659;
  assign n4660 = ~n4771 | ~DATAI_6_;
  assign n4662 = n5774 | n7529;
  assign n4674 = ~n4663 | ~n4662;
  assign n4667 = n4666 | n4665;
  assign n4668 = ~n4639 | ~IR_REG_31__SCAN_IN;
  assign n4671 = ~n4668 | ~IR_REG_22__SCAN_IN;
  assign n4669 = ~IR_REG_22__SCAN_IN;
  assign n4670 = ~n4669 | ~IR_REG_31__SCAN_IN;
  assign n4673 = ~n4671 | ~n4670;
  assign n5666 = ~n4673 | ~n4672;
  assign n6216 = ~n5666;
  assign n5278 = ~n7516 | ~n6216;
  assign n4803 = n4674 ^ ~n5700;
  assign n7784 = ~n5666 | ~n6105;
  assign n4907 = n4730 & n7572;
  assign n4676 = ~n5778 | ~n7503;
  assign n4675 = ~n4934 | ~n7534;
  assign n4804 = n4676 & n4675;
  assign n7001 = n4803 | n4804;
  assign n4720 = ~n7001;
  assign n4678 = ~REG3_REG_5__SCAN_IN;
  assign n4677 = ~REG3_REG_4__SCAN_IN | ~REG3_REG_3__SCAN_IN;
  assign n4679 = ~n4678 | ~n4677;
  assign n7553 = ~n4812 | ~n4679;
  assign n4680 = ~n4894 | ~REG1_REG_5__SCAN_IN;
  assign n4684 = ~n5188 | ~REG0_REG_5__SCAN_IN;
  assign n4683 = ~n4359 | ~REG2_REG_5__SCAN_IN;
  assign n4685 = n4684 & n4683;
  assign n4693 = ~n7583 | ~n4934;
  assign n4688 = ~n4687 | ~IR_REG_31__SCAN_IN;
  assign n4689 = ~n7768;
  assign n4691 = n4771 | n4689;
  assign n4690 = ~n4771 | ~DATAI_5_;
  assign n4692 = n5774 | n7563;
  assign n4696 = ~n5778 | ~n7583;
  assign n4695 = ~n4934 | ~n7571;
  assign n4723 = ~n6898;
  assign n4698 = ~n5188 | ~REG0_REG_4__SCAN_IN;
  assign n4697 = ~n4359 | ~REG2_REG_4__SCAN_IN;
  assign n4702 = n4698 & n4697;
  assign n4700 = ~n6015 | ~REG1_REG_4__SCAN_IN;
  assign n7602 = REG3_REG_4__SCAN_IN ^ ~REG3_REG_3__SCAN_IN;
  assign n4699 = n5544 | n7602;
  assign n4710 = ~n7617 | ~n4934;
  assign n4790 = ~n4703 | ~IR_REG_31__SCAN_IN;
  assign n4704 = ~n4790 | ~n4789;
  assign n4706 = ~n4704 | ~IR_REG_31__SCAN_IN;
  assign n7079 = n4706 ^ ~n4705;
  assign n4708 = n4771 | n7079;
  assign n6020 = ~n4360;
  assign n4707 = ~n6020 | ~DATAI_4_;
  assign n4709 = n5774 | n7599;
  assign n4712 = ~n4710 | ~n4709;
  assign n4722 = n4712 ^ ~n4711;
  assign n4714 = ~n5778 | ~n7617;
  assign n7584 = ~n7599;
  assign n4713 = ~n4362 | ~n7584;
  assign n4721 = ~n4714 | ~n4713;
  assign n6895 = ~n4722 | ~n4721;
  assign n4719 = n4723 | n6895;
  assign n4717 = ~n4715;
  assign n4718 = ~n4717 | ~n4716;
  assign n7000 = ~n4719 | ~n4718;
  assign n6909 = n4722 ^ ~n4721;
  assign n4802 = n6909 | n4723;
  assign n4724 = ~n4760 | ~REG3_REG_1__SCAN_IN;
  assign n4732 = ~n5496 | ~n4362;
  assign n4728 = n4771 | n5348;
  assign n4727 = ~n4771 | ~DATAI_1_;
  assign n4729 = ~n7670;
  assign n4731 = ~n4730 | ~n4729;
  assign n4733 = ~n4732 | ~n4731;
  assign n4735 = ~n4907 | ~n5496;
  assign n4734 = ~n4362 | ~n4729;
  assign n4756 = ~n4735 | ~n4734;
  assign n6858 = n4757 ^ ~n4756;
  assign n4737 = ~n4894 | ~REG1_REG_0__SCAN_IN;
  assign n4736 = ~n4890 | ~REG0_REG_0__SCAN_IN;
  assign n4739 = ~n4760 | ~REG3_REG_0__SCAN_IN;
  assign n4738 = ~n4891 | ~REG2_REG_0__SCAN_IN;
  assign n4748 = ~n4907 | ~n6854;
  assign n4740 = ~IR_REG_0__SCAN_IN;
  assign n4742 = n4771 | n4740;
  assign n4741 = ~n4771 | ~DATAI_0_;
  assign n5568 = n4742 & n4741;
  assign n5578 = ~n5568;
  assign n4746 = ~n4934 | ~n5578;
  assign n4744 = ~n4743;
  assign n4745 = ~n4744 | ~IR_REG_0__SCAN_IN;
  assign n4747 = n4746 & n4745;
  assign n4750 = ~n6854 | ~n4934;
  assign n4749 = ~n4730 | ~n5578;
  assign n4753 = ~n4750 | ~n4749;
  assign n4752 = ~n4753;
  assign n4751 = ~REG1_REG_0__SCAN_IN;
  assign n5457 = ~n4752 | ~n4585;
  assign n4755 = ~n5456 | ~n5457;
  assign n4758 = ~n4757 | ~n4756;
  assign n4762 = ~n4760 | ~REG3_REG_2__SCAN_IN;
  assign n4761 = ~n4894 | ~REG1_REG_2__SCAN_IN;
  assign n4766 = n4762 & n4761;
  assign n4764 = ~n4890 | ~REG0_REG_2__SCAN_IN;
  assign n4763 = ~n4891 | ~REG2_REG_2__SCAN_IN;
  assign n4765 = n4764 & n4763;
  assign n4775 = ~n7680 | ~n4362;
  assign n4773 = n4771 | n4358;
  assign n4772 = ~n4771 | ~DATAI_2_;
  assign n4774 = n5774 | n5567;
  assign n4776 = n4775 & n4774;
  assign n4780 = n4776 ^ ~n4711;
  assign n4778 = ~n4907 | ~n7680;
  assign n7652 = ~n5567;
  assign n4777 = ~n4362 | ~n7652;
  assign n4779 = n4778 & n4777;
  assign n4782 = ~n4780 | ~n4779;
  assign n4781 = n4780 | n4779;
  assign n6980 = ~n4782 | ~n4781;
  assign n4784 = ~n5188 | ~REG0_REG_3__SCAN_IN;
  assign n4783 = ~n4359 | ~REG2_REG_3__SCAN_IN;
  assign n4788 = n4784 & n4783;
  assign n4786 = ~n6015 | ~REG1_REG_3__SCAN_IN;
  assign n4785 = n5544 | REG3_REG_3__SCAN_IN;
  assign n4793 = ~n7651 | ~n4934;
  assign n5352 = n4790 ^ ~n4789;
  assign n4791 = n4771 | n5352;
  assign n4792 = n5774 | n7629;
  assign n4794 = ~n4793 | ~n4792;
  assign n4798 = n4794 ^ ~n4711;
  assign n4796 = ~n5778 | ~n7651;
  assign n4795 = ~n4362 | ~n7618;
  assign n4797 = ~n4796 | ~n4795;
  assign n4800 = n4798 | n4797;
  assign n4799 = ~n4798 | ~n4797;
  assign n6833 = n4800 & n4799;
  assign n6894 = ~n4801 | ~n4800;
  assign n6998 = n4802 | n6894;
  assign n4806 = ~n4803;
  assign n4805 = ~n4804;
  assign n4808 = ~n4890 | ~REG0_REG_7__SCAN_IN;
  assign n4807 = ~n4359 | ~REG2_REG_7__SCAN_IN;
  assign n4815 = ~n6015 | ~REG1_REG_7__SCAN_IN;
  assign n4810 = ~n4812 & ~n4809;
  assign n4813 = ~n4810 & ~REG3_REG_7__SCAN_IN;
  assign n7521 = n4813 | n4918;
  assign n4814 = n5544 | n7521;
  assign n4824 = ~n7486 | ~n4362;
  assign n4818 = ~IR_REG_6__SCAN_IN;
  assign n4819 = ~n4857 | ~n4818;
  assign n4835 = ~n4819 | ~IR_REG_31__SCAN_IN;
  assign n7762 = n4835 ^ ~IR_REG_7__SCAN_IN;
  assign n4820 = ~n7762;
  assign n4822 = n4771 | n4820;
  assign n4821 = ~n4771 | ~DATAI_7_;
  assign n4823 = n5774 | n7514;
  assign n4825 = ~n4824 | ~n4823;
  assign n4980 = n4825 ^ ~n5700;
  assign n4827 = ~n5778 | ~n7486;
  assign n4826 = ~n4934 | ~n7504;
  assign n4981 = ~n4827 | ~n4826;
  assign n6796 = n4980 ^ ~n4981;
  assign n4829 = ~n4890 | ~REG0_REG_8__SCAN_IN;
  assign n4828 = ~n4359 | ~REG2_REG_8__SCAN_IN;
  assign n4833 = n4829 & n4828;
  assign n4831 = ~n6015 | ~REG1_REG_8__SCAN_IN;
  assign n7465 = n4918 ^ ~REG3_REG_8__SCAN_IN;
  assign n4830 = n5544 | n7465;
  assign n4832 = n4831 & n4830;
  assign n4841 = ~n7451 | ~n4362;
  assign n4834 = ~IR_REG_7__SCAN_IN;
  assign n4836 = ~n4835 | ~n4834;
  assign n4837 = ~n4836 | ~IR_REG_31__SCAN_IN;
  assign n7759 = n4837 ^ ~IR_REG_8__SCAN_IN;
  assign n4839 = n4771 | n5366;
  assign n4838 = ~n4771 | ~DATAI_8_;
  assign n4840 = n5774 | n7468;
  assign n4842 = ~n4841 | ~n4840;
  assign n4983 = n4842 ^ ~n4711;
  assign n4844 = ~n5778 | ~n7451;
  assign n7471 = ~n7468;
  assign n4843 = ~n4934 | ~n7471;
  assign n4984 = ~n4844 | ~n4843;
  assign n4845 = n6796 & n6845;
  assign n4847 = ~n5188 | ~REG0_REG_12__SCAN_IN;
  assign n4846 = ~n4359 | ~REG2_REG_12__SCAN_IN;
  assign n4853 = n4847 & n4846;
  assign n4851 = ~n6015 | ~REG1_REG_12__SCAN_IN;
  assign n4849 = ~REG3_REG_11__SCAN_IN | ~REG3_REG_10__SCAN_IN;
  assign n4945 = ~REG3_REG_12__SCAN_IN;
  assign n7387 = n4948 ^ ~n4945;
  assign n4850 = n5544 | n7387;
  assign n4852 = n4851 & n4850;
  assign n4867 = ~n7394 | ~n4362;
  assign n4854 = ~IR_REG_8__SCAN_IN;
  assign n4856 = n4855 & n4854;
  assign n4926 = ~n4857 | ~n4856;
  assign n4859 = ~n4926;
  assign n4858 = ~IR_REG_9__SCAN_IN;
  assign n4860 = ~n4878 & ~IR_REG_10__SCAN_IN;
  assign n4900 = n4860 | n4767;
  assign n4861 = ~IR_REG_11__SCAN_IN;
  assign n4862 = ~n4900 | ~n4861;
  assign n4863 = ~n4862 | ~IR_REG_31__SCAN_IN;
  assign n4865 = ~n7747 | ~n4360;
  assign n4864 = ~n6020 | ~DATAI_12_;
  assign n4866 = n5774 | n7379;
  assign n4868 = ~n4867 | ~n4866;
  assign n4915 = n4868 ^ ~n4711;
  assign n4870 = ~n5778 | ~n7394;
  assign n4869 = ~n4934 | ~n7368;
  assign n4914 = ~n4870 | ~n4869;
  assign n4895 = ~REG3_REG_10__SCAN_IN;
  assign n7435 = n4920 ^ ~n4895;
  assign n4871 = ~n7435;
  assign n4872 = ~n4894 | ~REG1_REG_10__SCAN_IN;
  assign n4875 = ~n5188 | ~REG0_REG_10__SCAN_IN;
  assign n4874 = ~n4359 | ~REG2_REG_10__SCAN_IN;
  assign n4876 = n4875 & n4874;
  assign n4885 = ~n4877 | ~n4876;
  assign n4883 = ~n4885 | ~n4362;
  assign n4881 = ~n6020 | ~DATAI_10_;
  assign n4879 = ~n4878 | ~IR_REG_31__SCAN_IN;
  assign n5326 = ~n7753;
  assign n4880 = n4771 | n5326;
  assign n4882 = ~n4730 | ~n4886;
  assign n4884 = ~n4883 | ~n4882;
  assign n4889 = ~n5020;
  assign n4888 = ~n4907 | ~n4885;
  assign n4887 = ~n4934 | ~n4886;
  assign n5019 = ~n4888 | ~n4887;
  assign n6964 = ~n4889 | ~n5019;
  assign n4893 = ~n4890 | ~REG0_REG_11__SCAN_IN;
  assign n4892 = ~n4891 | ~REG2_REG_11__SCAN_IN;
  assign n4899 = ~n4593 & ~n4594;
  assign n4896 = n4920 | n4895;
  assign n6952 = ~REG3_REG_11__SCAN_IN;
  assign n4897 = ~n4896 | ~n6952;
  assign n7407 = ~n4897 | ~n4948;
  assign n4898 = n5544 | n7407;
  assign n4906 = ~n4899 | ~n4898;
  assign n4904 = ~n4906 | ~n4934;
  assign n4902 = ~n4360 | ~n7750;
  assign n4901 = ~n4771 | ~DATAI_11_;
  assign n4905 = ~n4904 | ~n4903;
  assign n4909 = ~n4907 | ~n4906;
  assign n7405 = ~n6954;
  assign n4908 = ~n4362 | ~n7405;
  assign n5017 = ~n4909 | ~n4908;
  assign n4910 = ~n5018 & ~n5017;
  assign n4913 = n6964 | n4910;
  assign n4912 = ~n5018;
  assign n4911 = ~n5017;
  assign n6873 = ~n6878 & ~n6875;
  assign n4917 = ~n4890 | ~REG0_REG_9__SCAN_IN;
  assign n4916 = ~n4359 | ~REG2_REG_9__SCAN_IN;
  assign n4925 = n4917 & n4916;
  assign n4923 = ~n6015 | ~REG1_REG_9__SCAN_IN;
  assign n4919 = ~n4918 | ~REG3_REG_8__SCAN_IN;
  assign n6915 = ~REG3_REG_9__SCAN_IN;
  assign n4921 = ~n4919 | ~n6915;
  assign n7440 = ~n4921 | ~n4920;
  assign n4922 = n5544 | n7440;
  assign n4924 = n4923 & n4922;
  assign n4932 = ~n6840 | ~n4934;
  assign n4927 = ~n4926 | ~IR_REG_31__SCAN_IN;
  assign n7756 = n4927 ^ ~IR_REG_9__SCAN_IN;
  assign n4928 = ~n7756;
  assign n4930 = n4771 | n4928;
  assign n4929 = ~n6020 | ~DATAI_9_;
  assign n4931 = n5774 | n6921;
  assign n4933 = ~n4932 | ~n4931;
  assign n4937 = n4933 ^ ~n4711;
  assign n4936 = ~n5778 | ~n6840;
  assign n4935 = ~n4362 | ~n7452;
  assign n4938 = ~n4936 | ~n4935;
  assign n4940 = ~n4937;
  assign n4939 = ~n4938;
  assign n4941 = n4940 | n4939;
  assign n6917 = ~n6820 | ~n4941;
  assign n4942 = ~n6917;
  assign n6937 = ~n4373 | ~n4942;
  assign n4944 = ~n5188 | ~REG0_REG_13__SCAN_IN;
  assign n4943 = ~n4359 | ~REG2_REG_13__SCAN_IN;
  assign n4953 = n4944 & n4943;
  assign n4951 = ~n6015 | ~REG1_REG_13__SCAN_IN;
  assign n4946 = ~n4948 & ~n4945;
  assign n4949 = ~n4946 & ~REG3_REG_13__SCAN_IN;
  assign n4947 = ~REG3_REG_12__SCAN_IN | ~REG3_REG_13__SCAN_IN;
  assign n7336 = n4949 | n4965;
  assign n4950 = n5544 | n7336;
  assign n4952 = n4951 & n4950;
  assign n4959 = ~n7314 | ~n4934;
  assign n4954 = n4646 | n4767;
  assign n7744 = n4954 ^ ~IR_REG_13__SCAN_IN;
  assign n4955 = ~n7744;
  assign n4957 = n4771 | n4955;
  assign n4956 = ~n6020 | ~DATAI_13_;
  assign n4958 = n5774 | n7330;
  assign n4960 = ~n4959 | ~n4958;
  assign n5014 = n4960 ^ ~n5700;
  assign n4962 = ~n5778 | ~n7314;
  assign n4961 = ~n4362 | ~n7352;
  assign n4964 = ~n5188 | ~REG0_REG_14__SCAN_IN;
  assign n4963 = ~n4359 | ~REG2_REG_14__SCAN_IN;
  assign n4970 = n4964 & n4963;
  assign n4968 = ~n6015 | ~REG1_REG_14__SCAN_IN;
  assign n5029 = n4965 & REG3_REG_14__SCAN_IN;
  assign n4966 = ~n4965 & ~REG3_REG_14__SCAN_IN;
  assign n7305 = n5029 | n4966;
  assign n4967 = n5544 | n7305;
  assign n4969 = n4968 & n4967;
  assign n4976 = ~n7351 | ~n4934;
  assign n4972 = ~n4971 | ~IR_REG_31__SCAN_IN;
  assign n7741 = n4972 ^ ~IR_REG_14__SCAN_IN;
  assign n4974 = n4771 | n5383;
  assign n4973 = ~n6020 | ~DATAI_14_;
  assign n4975 = n5774 | n5610;
  assign n4977 = ~n4976 | ~n4975;
  assign n4992 = n4977 ^ ~n5700;
  assign n4979 = ~n5778 | ~n7351;
  assign n4978 = ~n4362 | ~n7315;
  assign n5023 = ~n5862;
  assign n4988 = ~n6845;
  assign n4982 = ~n4980;
  assign n5856 = ~n4982 | ~n4981;
  assign n4986 = ~n4983;
  assign n4985 = ~n4984;
  assign n4987 = n5856 & n6846;
  assign n4989 = ~n4988 & ~n4987;
  assign n4990 = n5023 | n4989;
  assign n4995 = ~n4992;
  assign n4994 = ~n4993;
  assign n4997 = ~n5188 | ~REG0_REG_15__SCAN_IN;
  assign n4996 = ~n4359 | ~REG2_REG_15__SCAN_IN;
  assign n5001 = n4997 & n4996;
  assign n4999 = ~n6015 | ~REG1_REG_15__SCAN_IN;
  assign n7292 = n5029 ^ ~REG3_REG_15__SCAN_IN;
  assign n4998 = n5544 | n7292;
  assign n5000 = n4999 & n4998;
  assign n5008 = ~n7316 | ~n4362;
  assign n5002 = ~IR_REG_14__SCAN_IN;
  assign n5003 = ~n4575 | ~n5002;
  assign n5033 = ~n5003 | ~IR_REG_31__SCAN_IN;
  assign n7738 = n5033 ^ ~IR_REG_15__SCAN_IN;
  assign n5004 = ~n7738;
  assign n5006 = n5004 | n4771;
  assign n5005 = ~n6020 | ~DATAI_15_;
  assign n5007 = n5774 | n6732;
  assign n5009 = ~n5008 | ~n5007;
  assign n5867 = n5009 ^ ~n4711;
  assign n5011 = ~n5778 | ~n7316;
  assign n5010 = ~n4362 | ~n5609;
  assign n5980 = ~n5011 | ~n5010;
  assign n5012 = n5867 | n5980;
  assign n5016 = n5863 & n5012;
  assign n5015 = ~n6941 | ~n5862;
  assign n6962 = n5020 ^ ~n5019;
  assign n6872 = n6966 & n6962;
  assign n5022 = n5021 & n6872;
  assign n5024 = ~n5860 & ~n5023;
  assign n5050 = ~n5026 | ~n5025;
  assign n5028 = ~n5188 | ~REG0_REG_16__SCAN_IN;
  assign n5027 = ~n4359 | ~REG2_REG_16__SCAN_IN;
  assign n5055 = n5029 & REG3_REG_15__SCAN_IN;
  assign n5877 = REG3_REG_16__SCAN_IN ^ ~n5055;
  assign n5030 = n5544 | n5877;
  assign n5039 = ~n7958 | ~n4934;
  assign n5032 = ~IR_REG_15__SCAN_IN;
  assign n5034 = ~n5033 | ~n5032;
  assign n5035 = ~n5034 | ~IR_REG_31__SCAN_IN;
  assign n7735 = n5035 ^ ~IR_REG_16__SCAN_IN;
  assign n5037 = ~n7735 | ~n4360;
  assign n5036 = ~n6020 | ~DATAI_16_;
  assign n5038 = n5774 | n6610;
  assign n5040 = ~n5039 | ~n5038;
  assign n5043 = n5040 ^ ~n4711;
  assign n5042 = ~n5778 | ~n7958;
  assign n6598 = ~n6610;
  assign n5041 = ~n4934 | ~n6598;
  assign n5044 = ~n5042 | ~n5041;
  assign n5046 = ~n5043;
  assign n5045 = ~n5044;
  assign n5047 = n5046 | n5045;
  assign n5875 = ~n5051 | ~n5047;
  assign n5048 = n5867 & n5980;
  assign n5049 = ~n5875 & ~n5048;
  assign n5052 = ~n5050 | ~n5049;
  assign n5889 = ~n5052 | ~n5051;
  assign n5054 = ~n5188 | ~REG0_REG_17__SCAN_IN;
  assign n5053 = ~n4359 | ~REG2_REG_17__SCAN_IN;
  assign n5060 = n5054 & n5053;
  assign n5897 = REG3_REG_17__SCAN_IN ^ ~n5076;
  assign n5058 = n5544 | n5897;
  assign n5056 = ~REG1_REG_17__SCAN_IN;
  assign n5057 = n5525 | n5056;
  assign n5059 = n5058 & n5057;
  assign n7961 = ~n5060 | ~n5059;
  assign n5066 = ~n7961 | ~n4362;
  assign n5062 = n5061 | n4767;
  assign n7732 = n5062 ^ ~IR_REG_17__SCAN_IN;
  assign n5064 = ~n4360 | ~n7732;
  assign n5063 = ~n6020 | ~DATAI_17_;
  assign n5065 = n5774 | n5902;
  assign n5067 = ~n5066 | ~n5065;
  assign n5070 = n5067 ^ ~n5700;
  assign n5069 = ~n5778 | ~n7961;
  assign n5068 = ~n4934 | ~n6583;
  assign n5887 = n5889 & n5890;
  assign n5073 = ~n5070;
  assign n5072 = ~n5071;
  assign n5075 = ~n5188 | ~REG0_REG_18__SCAN_IN;
  assign n5074 = ~n4359 | ~REG2_REG_18__SCAN_IN;
  assign n5081 = n5075 & n5074;
  assign n5967 = REG3_REG_18__SCAN_IN ^ ~n5095;
  assign n5079 = n5544 | n5967;
  assign n5077 = ~REG1_REG_18__SCAN_IN;
  assign n5078 = n5525 | n5077;
  assign n5080 = n5079 & n5078;
  assign n7964 = ~n5081 | ~n5080;
  assign n5087 = ~n7964 | ~n4934;
  assign n5083 = n5082 | n4767;
  assign n7729 = n5083 ^ ~IR_REG_18__SCAN_IN;
  assign n5085 = ~n7729 | ~n4360;
  assign n5084 = ~n6020 | ~DATAI_18_;
  assign n5086 = n5774 | n5972;
  assign n5088 = ~n5087 | ~n5086;
  assign n5092 = n5088 ^ ~n5700;
  assign n5090 = ~n5778 | ~n7964;
  assign n5089 = ~n4362 | ~n6543;
  assign n5961 = ~n5092 & ~n5091;
  assign n5094 = ~n5188 | ~REG0_REG_19__SCAN_IN;
  assign n5093 = ~n4359 | ~REG2_REG_19__SCAN_IN;
  assign n5099 = n5094 & n5093;
  assign n6521 = REG3_REG_19__SCAN_IN ^ ~n5114;
  assign n5097 = ~n4760 | ~n6521;
  assign n5096 = ~n6015 | ~REG1_REG_19__SCAN_IN;
  assign n5098 = n5097 & n5096;
  assign n5177 = ~n4934;
  assign n5103 = ~n5969 & ~n5177;
  assign n5101 = n7516 | n4771;
  assign n5100 = ~n6020 | ~DATAI_19_;
  assign n5102 = ~n5826 & ~n5774;
  assign n5104 = ~n5103 & ~n5102;
  assign n5107 = n4711 ^ n5104;
  assign n7967 = ~n5969;
  assign n5106 = ~n5778 | ~n7967;
  assign n5105 = ~n4362 | ~n6517;
  assign n5108 = ~n5106 | ~n5105;
  assign n5111 = ~n5107 | ~n5108;
  assign n5110 = ~n5107;
  assign n5109 = ~n5108;
  assign n5112 = ~n5110 | ~n5109;
  assign n5823 = ~n5111 | ~n5112;
  assign n5113 = ~n5112;
  assign n5929 = ~n5822 & ~n5113;
  assign n5395 = ~REG3_REG_19__SCAN_IN;
  assign n6495 = n5133 ^ ~REG3_REG_20__SCAN_IN;
  assign n5121 = n6495 | n5544;
  assign n5116 = ~n5188 | ~REG0_REG_20__SCAN_IN;
  assign n5115 = ~n4359 | ~REG2_REG_20__SCAN_IN;
  assign n5119 = ~n5116 | ~n5115;
  assign n5117 = ~REG1_REG_20__SCAN_IN;
  assign n5118 = ~n5525 & ~n5117;
  assign n5120 = ~n5119 & ~n5118;
  assign n7970 = ~n5121 | ~n5120;
  assign n5123 = ~n7970 | ~n4934;
  assign n6489 = ~n6020 | ~DATAI_20_;
  assign n5122 = n5774 | n6489;
  assign n5124 = ~n5123 | ~n5122;
  assign n5127 = n5124 ^ ~n5700;
  assign n5126 = ~n7970 | ~n5778;
  assign n5621 = ~n6489;
  assign n5125 = ~n4362 | ~n5621;
  assign n5128 = n5126 & n5125;
  assign n5837 = ~n5127 & ~n5128;
  assign n5147 = n5929 | n5837;
  assign n5130 = ~n5127;
  assign n5129 = ~n5128;
  assign n5927 = n5130 | n5129;
  assign n5132 = ~n4890 | ~REG0_REG_21__SCAN_IN;
  assign n5131 = ~n4359 | ~REG2_REG_21__SCAN_IN;
  assign n5138 = n5132 & n5131;
  assign n5844 = REG3_REG_21__SCAN_IN ^ ~n5151;
  assign n5136 = n5544 | n5844;
  assign n5134 = ~REG1_REG_21__SCAN_IN;
  assign n5135 = n5525 | n5134;
  assign n5137 = n5136 & n5135;
  assign n7973 = ~n5138 | ~n5137;
  assign n5140 = ~n7973 | ~n4934;
  assign n6448 = ~n6020 | ~DATAI_21_;
  assign n5139 = n5774 | n6448;
  assign n5141 = ~n5140 | ~n5139;
  assign n5840 = n5141 ^ ~n4711;
  assign n5143 = ~n5778 | ~n7973;
  assign n6437 = ~n6448;
  assign n5142 = ~n4362 | ~n6437;
  assign n5839 = ~n5143 | ~n5142;
  assign n5144 = n5840 | n5839;
  assign n5145 = ~n5927 | ~n5144;
  assign n5146 = ~n5145;
  assign n5148 = ~n5840 | ~n5839;
  assign n5150 = ~n6015 | ~REG1_REG_22__SCAN_IN;
  assign n5149 = ~n4359 | ~REG2_REG_22__SCAN_IN;
  assign n5157 = n5150 & n5149;
  assign n6423 = REG3_REG_22__SCAN_IN ^ ~n5172;
  assign n5152 = ~REG0_REG_22__SCAN_IN;
  assign n5154 = n5153 | n5152;
  assign n5156 = n5155 & n5154;
  assign n5159 = ~n7976 | ~n4362;
  assign n6419 = ~n6020 | ~DATAI_22_;
  assign n5158 = n5774 | n6419;
  assign n5160 = ~n5159 | ~n5158;
  assign n5163 = n5160 ^ ~n5700;
  assign n5162 = ~n5778 | ~n7976;
  assign n6410 = ~n6419;
  assign n5161 = ~n4934 | ~n6410;
  assign n5164 = n5162 & n5161;
  assign n5168 = ~n5163 | ~n5164;
  assign n5166 = ~n5163;
  assign n5165 = ~n5164;
  assign n5167 = ~n5166 | ~n5165;
  assign n5944 = ~n5168 | ~n5167;
  assign n5169 = ~n5168;
  assign n5171 = ~n4890 | ~REG0_REG_23__SCAN_IN;
  assign n5170 = ~n4359 | ~REG2_REG_23__SCAN_IN;
  assign n5176 = n5171 & n5170;
  assign n5174 = ~n6015 | ~REG1_REG_23__SCAN_IN;
  assign n6399 = REG3_REG_23__SCAN_IN ^ ~n5191;
  assign n5173 = n5544 | n6399;
  assign n5175 = n5174 & n5173;
  assign n5179 = ~n6345 & ~n5177;
  assign n5815 = ~n6020 | ~DATAI_23_;
  assign n5178 = ~n5774 & ~n5815;
  assign n5180 = ~n5179 & ~n5178;
  assign n5185 = n4711 ^ n5180;
  assign n5199 = ~n5778;
  assign n5182 = ~n6345 & ~n5199;
  assign n5181 = ~n5177 & ~n5815;
  assign n5183 = ~n5182 & ~n5181;
  assign n5807 = n5185 ^ ~n5183;
  assign n5187 = ~n5808 | ~n5807;
  assign n5184 = ~n5183;
  assign n5186 = ~n5185 | ~n5184;
  assign n5909 = ~n5187 | ~n5186;
  assign n5190 = ~n5188 | ~REG0_REG_24__SCAN_IN;
  assign n5189 = ~n4359 | ~REG2_REG_24__SCAN_IN;
  assign n5195 = n5190 & n5189;
  assign n5193 = ~n6015 | ~REG1_REG_24__SCAN_IN;
  assign n5914 = REG3_REG_24__SCAN_IN ^ ~n5209;
  assign n5192 = n5544 | n5914;
  assign n5194 = n5193 & n5192;
  assign n5197 = ~n6315 & ~n5177;
  assign n5920 = ~n6020 | ~DATAI_24_;
  assign n5196 = ~n5774 & ~n5920;
  assign n5198 = ~n5197 & ~n5196;
  assign n5911 = n5198 ^ ~n4711;
  assign n5201 = ~n6315 & ~n5199;
  assign n5200 = ~n5177 & ~n5920;
  assign n5203 = ~n5201 & ~n5200;
  assign n5202 = ~n5911 | ~n5203;
  assign n5206 = ~n5909 | ~n5202;
  assign n5204 = ~n5911;
  assign n5910 = ~n5203;
  assign n5205 = ~n5204 | ~n5910;
  assign n5208 = ~n6015 | ~REG1_REG_25__SCAN_IN;
  assign n5207 = ~n5188 | ~REG0_REG_25__SCAN_IN;
  assign n5213 = ~n5208 | ~n5207;
  assign n5271 = ~n5209 | ~REG3_REG_24__SCAN_IN;
  assign n6322 = REG3_REG_25__SCAN_IN ^ ~n5271;
  assign n5211 = ~n4760 | ~n6322;
  assign n5210 = ~n4359 | ~REG2_REG_25__SCAN_IN;
  assign n5212 = ~n5211 | ~n5210;
  assign n5215 = ~n7985 | ~n4934;
  assign n6330 = ~n6020 | ~DATAI_25_;
  assign n5214 = n5774 | n6330;
  assign n5216 = ~n5215 | ~n5214;
  assign n5219 = n5216 ^ ~n5700;
  assign n5218 = ~n5778 | ~n7985;
  assign n5657 = ~n6330;
  assign n5217 = ~n4934 | ~n5657;
  assign n5220 = n5218 & n5217;
  assign n5697 = ~n5219 | ~n5220;
  assign n5737 = ~n5697;
  assign n5222 = ~n5219;
  assign n5221 = ~n5220;
  assign n5735 = n5222 & n5221;
  assign n5223 = ~n5737 & ~n5735;
  assign n5270 = n5736 ^ ~n5223;
  assign n5225 = ~n5416;
  assign n5226 = ~n5224 | ~n5225;
  assign n5229 = ~n5226 | ~B_REG_SCAN_IN;
  assign n5227 = ~B_REG_SCAN_IN;
  assign n5228 = ~n5224 | ~n5227;
  assign n5230 = ~n5229 | ~n5228;
  assign n7721 = ~n5230 | ~n5419;
  assign n5232 = n7721 | D_REG_0__SCAN_IN;
  assign n7773 = ~n5419;
  assign n5231 = ~n5224 | ~n7773;
  assign n5238 = ~D_REG_6__SCAN_IN & ~D_REG_7__SCAN_IN;
  assign n5236 = D_REG_8__SCAN_IN | D_REG_9__SCAN_IN;
  assign n5234 = ~D_REG_10__SCAN_IN & ~D_REG_11__SCAN_IN;
  assign n5233 = ~D_REG_12__SCAN_IN & ~D_REG_13__SCAN_IN;
  assign n5235 = ~n5234 | ~n5233;
  assign n5237 = ~n5236 & ~n5235;
  assign n5254 = ~n5238 | ~n5237;
  assign n5240 = ~D_REG_18__SCAN_IN & ~D_REG_19__SCAN_IN;
  assign n5239 = ~D_REG_20__SCAN_IN & ~D_REG_21__SCAN_IN;
  assign n5244 = ~n5240 | ~n5239;
  assign n5242 = ~D_REG_16__SCAN_IN & ~D_REG_14__SCAN_IN;
  assign n5241 = ~D_REG_15__SCAN_IN & ~D_REG_17__SCAN_IN;
  assign n5243 = ~n5242 | ~n5241;
  assign n5252 = ~n5244 & ~n5243;
  assign n5246 = ~D_REG_26__SCAN_IN & ~D_REG_27__SCAN_IN;
  assign n5245 = ~D_REG_28__SCAN_IN & ~D_REG_31__SCAN_IN;
  assign n5250 = ~n5246 | ~n5245;
  assign n5248 = ~D_REG_22__SCAN_IN & ~D_REG_23__SCAN_IN;
  assign n5247 = ~D_REG_24__SCAN_IN & ~D_REG_25__SCAN_IN;
  assign n5249 = ~n5248 | ~n5247;
  assign n5251 = ~n5250 & ~n5249;
  assign n5253 = ~n5252 | ~n5251;
  assign n5259 = ~n5254 & ~n5253;
  assign n5256 = ~D_REG_2__SCAN_IN & ~D_REG_3__SCAN_IN;
  assign n5255 = ~D_REG_4__SCAN_IN & ~D_REG_5__SCAN_IN;
  assign n5257 = ~n5256 | ~n5255;
  assign n5258 = ~D_REG_30__SCAN_IN & ~n5257;
  assign n5260 = ~n5259 | ~n5258;
  assign n5261 = ~D_REG_29__SCAN_IN & ~n5260;
  assign n5672 = ~n7721 & ~n5261;
  assign n5262 = n7721 | D_REG_1__SCAN_IN;
  assign n7780 = n5419 | n5416;
  assign n5674 = ~n5262 | ~n7780;
  assign n5679 = ~n5672 & ~n5674;
  assign n5266 = ~n5264 | ~IR_REG_23__SCAN_IN;
  assign n6215 = ~n5266 | ~n5265;
  assign n5343 = ~n4743 | ~n7774;
  assign n5295 = ~n5289 | ~n7720;
  assign n6203 = ~n5267;
  assign n5268 = n7516 | n7784;
  assign n5558 = ~n5666 & ~n6105;
  assign n5560 = ~n5558;
  assign n5269 = n5268 & n5560;
  assign n5288 = ~n7671 | ~n5269;
  assign n5309 = ~n5270 & ~n7007;
  assign n5299 = ~REG3_REG_25__SCAN_IN;
  assign n6301 = REG3_REG_26__SCAN_IN ^ n5521;
  assign n5277 = ~n6301 | ~n4760;
  assign n5273 = ~n6015 | ~REG1_REG_26__SCAN_IN;
  assign n5272 = ~n5188 | ~REG0_REG_26__SCAN_IN;
  assign n5275 = ~n5273 | ~n5272;
  assign n6295 = ~REG2_REG_26__SCAN_IN;
  assign n5274 = ~n4682 & ~n6295;
  assign n5276 = ~n5275 & ~n5274;
  assign n7988 = ~n5277 | ~n5276;
  assign n5279 = ~n5688 & ~n5278;
  assign n5286 = n5279 & n7720;
  assign n5298 = ~n5289 | ~n5286;
  assign n5282 = ~n5280;
  assign n5346 = ~n5282 | ~n5281;
  assign n5284 = ~n5346 | ~IR_REG_31__SCAN_IN;
  assign n7069 = n5284 ^ ~n5283;
  assign n7059 = ~n7069;
  assign n5307 = ~n7988 | ~n6991;
  assign n5285 = ~n7671 & ~U3149;
  assign n5287 = ~n5286 & ~n5285;
  assign n5453 = ~n5289 & ~n5287;
  assign n5451 = n5289 | n5288;
  assign n5290 = n5267 | n7712;
  assign n5450 = ~n5290 | ~n5558;
  assign n5291 = n4743 & n6215;
  assign n5292 = n5450 & n5291;
  assign n5293 = ~n5451 | ~n5292;
  assign n5294 = n5293 & STATE_REG_SCAN_IN;
  assign n5305 = ~n6798 | ~n6322;
  assign n5297 = n5295 | n7671;
  assign n5296 = n7516 | n6216;
  assign n6131 = ~n6105;
  assign n5670 = ~n7901 & ~n6131;
  assign n5303 = ~n6974 & ~n6330;
  assign n5301 = ~n6955 & ~n6315;
  assign n5300 = ~STATE_REG_SCAN_IN & ~n5299;
  assign n5302 = n5301 | n5300;
  assign n5304 = ~n5303 & ~n5302;
  assign n5306 = n5305 & n5304;
  assign n5308 = ~n5307 | ~n5306;
  assign n7124 = n7762 & REG1_REG_7__SCAN_IN;
  assign n7035 = IR_REG_0__SCAN_IN & REG1_REG_0__SCAN_IN;
  assign n5311 = ~n7034 | ~n7035;
  assign n7029 = ~n5348;
  assign n5310 = ~n7029 | ~REG1_REG_1__SCAN_IN;
  assign n7047 = n4358 ^ ~REG1_REG_2__SCAN_IN;
  assign n7048 = ~n7046 | ~n7047;
  assign n5313 = ~n7053 | ~REG1_REG_2__SCAN_IN;
  assign n5316 = ~n5441 | ~REG1_REG_3__SCAN_IN;
  assign n5447 = ~n5352;
  assign n5315 = ~n5314 | ~n5447;
  assign n5413 = ~n7079;
  assign n5318 = ~n5317 | ~n5413;
  assign n7096 = REG1_REG_5__SCAN_IN ^ n7768;
  assign n5319 = ~REG1_REG_5__SCAN_IN | ~n7768;
  assign n5322 = ~n7765 | ~n5321;
  assign n7125 = ~n7762 & ~REG1_REG_7__SCAN_IN;
  assign n7143 = n5323 ^ ~n5366;
  assign n5324 = ~n7759 | ~n5323;
  assign n7153 = REG1_REG_9__SCAN_IN ^ n7756;
  assign n5325 = ~REG1_REG_9__SCAN_IN | ~n7756;
  assign n5328 = ~n7753 | ~n5327;
  assign n7182 = REG1_REG_11__SCAN_IN ^ n7750;
  assign n5330 = ~n7747 | ~n5329;
  assign n7210 = REG1_REG_13__SCAN_IN ^ n7744;
  assign n5332 = ~n7741 | ~n5331;
  assign n7240 = REG1_REG_15__SCAN_IN ^ n7738;
  assign n5335 = ~REG1_REG_16__SCAN_IN & ~n7252;
  assign n5334 = ~n7735 & ~n5333;
  assign n7265 = REG1_REG_17__SCAN_IN ^ ~n7732;
  assign n5337 = ~n7266 & ~n7265;
  assign n5336 = ~REG1_REG_17__SCAN_IN & ~n7732;
  assign n7283 = REG1_REG_18__SCAN_IN ^ n7729;
  assign n5339 = ~n7282 | ~n7283;
  assign n5338 = ~REG1_REG_18__SCAN_IN | ~n7729;
  assign n5342 = ~n5339 | ~n5338;
  assign n5340 = ~REG1_REG_19__SCAN_IN;
  assign n5341 = n7516 ^ ~n5340;
  assign n5347 = n5342 ^ ~n5341;
  assign n6213 = n6215 | U3149;
  assign n5396 = ~n5343 | ~n6213;
  assign n5344 = ~n5558 | ~n6215;
  assign n5397 = n5344 & n4771;
  assign n7018 = ~n5396 | ~n5397;
  assign n7058 = ~n5346 | ~n5345;
  assign n7067 = ~n7058;
  assign n7077 = n7018 | n7067;
  assign n5405 = ~n5347 | ~n7284;
  assign n7027 = n5348 ^ ~REG2_REG_1__SCAN_IN;
  assign n7026 = ~IR_REG_0__SCAN_IN | ~REG2_REG_0__SCAN_IN;
  assign n7066 = ~n7026;
  assign n5350 = ~n7027 | ~n7066;
  assign n5349 = ~n7029 | ~REG2_REG_1__SCAN_IN;
  assign n7042 = ~n5350 | ~n5349;
  assign n7041 = ~n7042 | ~n7043;
  assign n5351 = ~n7053 | ~REG2_REG_2__SCAN_IN;
  assign n5355 = ~n5439 | ~REG2_REG_3__SCAN_IN;
  assign n5354 = ~n5353 | ~n5447;
  assign n5356 = ~n7083;
  assign n5359 = ~n5356 | ~REG2_REG_4__SCAN_IN;
  assign n5358 = ~n5357 | ~n5413;
  assign n7093 = ~n5359 | ~n5358;
  assign n7094 = REG2_REG_5__SCAN_IN ^ n7768;
  assign n5361 = ~n7093 | ~n7094;
  assign n5360 = ~REG2_REG_5__SCAN_IN | ~n7768;
  assign n5362 = ~n5361 | ~n5360;
  assign n7113 = n5362 ^ ~n4659;
  assign n7120 = ~n7765 | ~n5362;
  assign n5363 = ~n7762 | ~REG2_REG_7__SCAN_IN;
  assign n5364 = ~n5363;
  assign n7122 = n7762 ^ REG2_REG_7__SCAN_IN;
  assign n5365 = n5364 | n7122;
  assign n5369 = ~n7137 | ~REG2_REG_8__SCAN_IN;
  assign n5368 = ~n7759 | ~n5367;
  assign n7151 = REG2_REG_9__SCAN_IN ^ n7756;
  assign n5371 = ~n7150 | ~n7151;
  assign n5370 = ~REG2_REG_9__SCAN_IN | ~n7756;
  assign n5373 = ~n7753 | ~n5372;
  assign n7176 = REG2_REG_11__SCAN_IN ^ n7750;
  assign n5374 = ~REG2_REG_11__SCAN_IN | ~n7750;
  assign n7204 = ~n7192 | ~REG2_REG_12__SCAN_IN;
  assign n7205 = ~n7747 | ~n5377;
  assign n5379 = ~REG2_REG_13__SCAN_IN | ~n7744;
  assign n5378 = n7205 & n5379;
  assign n5382 = ~n7204 | ~n5378;
  assign n5380 = ~n5379;
  assign n7207 = REG2_REG_13__SCAN_IN ^ n7744;
  assign n5381 = n5380 | n7207;
  assign n5384 = n5382 & n5381;
  assign n5385 = ~n7741 | ~n5384;
  assign n7220 = n5384 ^ ~n5383;
  assign n7233 = REG2_REG_15__SCAN_IN ^ n7738;
  assign n5388 = ~REG2_REG_16__SCAN_IN & ~n7246;
  assign n5387 = ~n7735 & ~n5386;
  assign n7259 = REG2_REG_17__SCAN_IN ^ ~n7732;
  assign n5390 = ~n7258 & ~n7259;
  assign n5389 = ~REG2_REG_17__SCAN_IN & ~n7732;
  assign n7273 = ~n5390 & ~n5389;
  assign n7274 = REG2_REG_18__SCAN_IN ^ n7729;
  assign n5391 = ~REG2_REG_18__SCAN_IN | ~n7729;
  assign n5394 = n7069 | n7058;
  assign n7275 = ~n7018 & ~n5394;
  assign n5828 = ~STATE_REG_SCAN_IN & ~n5395;
  assign n5398 = ~n5396;
  assign n7270 = ~n5398 & ~n5397;
  assign n5399 = n7270 & ADDR_REG_19__SCAN_IN;
  assign n5400 = ~n5828 & ~n5399;
  assign n5403 = n5401 & n5400;
  assign n7080 = n7018 | n7059;
  assign n5402 = ~n7277 | ~n7712;
  assign U3259 = ~n5405 | ~n5404;
  assign n5406 = ~n7774;
  assign U4043 = ~n8000;
  assign n5408 = ~n7029 | ~STATE_REG_SCAN_IN;
  assign n5407 = ~DATAI_1_ | ~U3149;
  assign U3351 = ~n5408 | ~n5407;
  assign n5410 = ~n7053 | ~STATE_REG_SCAN_IN;
  assign n5409 = ~DATAI_2_ | ~U3149;
  assign U3350 = ~n5410 | ~n5409;
  assign n5412 = ~n5447 | ~STATE_REG_SCAN_IN;
  assign n5411 = ~DATAI_3_ | ~U3149;
  assign U3349 = ~n5412 | ~n5411;
  assign n5415 = ~n5413 | ~STATE_REG_SCAN_IN;
  assign n5414 = ~DATAI_4_ | ~U3149;
  assign U3348 = ~n5415 | ~n5414;
  assign n5418 = ~n5416 | ~STATE_REG_SCAN_IN;
  assign n5417 = ~DATAI_25_ | ~U3149;
  assign U3327 = ~n5418 | ~n5417;
  assign n5421 = ~n5419 | ~STATE_REG_SCAN_IN;
  assign n5420 = ~DATAI_26_ | ~U3149;
  assign U3326 = ~n5421 | ~n5420;
  assign n5423 = ~n6131 | ~STATE_REG_SCAN_IN;
  assign n5422 = ~DATAI_21_ | ~U3149;
  assign U3331 = ~n5423 | ~n5422;
  assign n6209 = ~n6216 | ~STATE_REG_SCAN_IN;
  assign n5424 = ~DATAI_22_ | ~U3149;
  assign U3330 = ~n6209 | ~n5424;
  assign n5426 = ~n7067 | ~STATE_REG_SCAN_IN;
  assign n5425 = ~DATAI_27_ | ~U3149;
  assign U3325 = ~n5426 | ~n5425;
  assign n5428 = ~n4461 | ~STATE_REG_SCAN_IN;
  assign n5427 = ~DATAI_29_ | ~U3149;
  assign U3323 = ~n5428 | ~n5427;
  assign n5431 = ~n5429 | ~STATE_REG_SCAN_IN;
  assign n5430 = ~DATAI_30_ | ~U3149;
  assign U3322 = ~n5431 | ~n5430;
  assign n5433 = ~n7059 | ~STATE_REG_SCAN_IN;
  assign n5432 = ~DATAI_28_ | ~U3149;
  assign U3324 = ~n5433 | ~n5432;
  assign n7776 = ~n5224;
  assign n5435 = ~n7776 | ~STATE_REG_SCAN_IN;
  assign n5434 = ~DATAI_24_ | ~U3149;
  assign U3328 = ~n5435 | ~n5434;
  assign n5437 = ~n7712 & ~U3149;
  assign n5436 = ~STATE_REG_SCAN_IN & ~DATAI_19_;
  assign U3333 = ~n5437 & ~n5436;
  assign n6826 = ~REG3_REG_3__SCAN_IN | ~U3149;
  assign n5438 = ~n7270 | ~ADDR_REG_3__SCAN_IN;
  assign n5446 = ~n6826 | ~n5438;
  assign n5440 = n5439 ^ REG2_REG_3__SCAN_IN;
  assign n5444 = ~n5440 | ~n7275;
  assign n5442 = n5441 ^ REG1_REG_3__SCAN_IN;
  assign n5443 = ~n7284 | ~n5442;
  assign n5445 = ~n5444 | ~n5443;
  assign n5449 = ~n5446 & ~n5445;
  assign n5448 = ~n7277 | ~n5447;
  assign U3243 = ~n5449 | ~n5448;
  assign n5452 = ~n5680 | ~n5451;
  assign n6983 = ~n5453 & ~n5452;
  assign n7019 = ~REG3_REG_0__SCAN_IN;
  assign n5461 = ~n6983 & ~n7019;
  assign n5455 = ~n6974 & ~n5568;
  assign n7650 = ~n5496;
  assign n5454 = ~n6951 & ~n7650;
  assign n5459 = ~n5455 & ~n5454;
  assign n7061 = n5457 ^ n5456;
  assign n6970 = ~n7007;
  assign n5458 = ~n7061 | ~n6970;
  assign n5460 = ~n5459 | ~n5458;
  assign U3229 = n5461 | n5460;
  assign n7957 = ~n8005;
  assign U3148 = ~n7270 & ~n7957;
  assign n5463 = ~n7617 | ~n7957;
  assign n5462 = ~n8005 | ~DATAO_REG_4__SCAN_IN;
  assign U3554 = ~n5463 | ~n5462;
  assign n5465 = ~n6854 | ~n7957;
  assign n5464 = ~n8005 | ~DATAO_REG_0__SCAN_IN;
  assign U3550 = ~n5465 | ~n5464;
  assign n5467 = ~n7393 | ~n7957;
  assign n5466 = ~n8000 | ~DATAO_REG_10__SCAN_IN;
  assign U3560 = ~n5467 | ~n5466;
  assign n5469 = ~n7451 | ~n7957;
  assign n5468 = ~n8005 | ~DATAO_REG_8__SCAN_IN;
  assign U3558 = ~n5469 | ~n5468;
  assign n5471 = ~n7394 | ~n7957;
  assign n5470 = ~n8000 | ~DATAO_REG_12__SCAN_IN;
  assign U3562 = ~n5471 | ~n5470;
  assign n5473 = ~n7503 | ~n7957;
  assign n5472 = ~n8005 | ~DATAO_REG_6__SCAN_IN;
  assign U3556 = ~n5473 | ~n5472;
  assign n5475 = ~n7651 | ~n7957;
  assign n5474 = ~n8005 | ~DATAO_REG_3__SCAN_IN;
  assign U3553 = ~n5475 | ~n5474;
  assign n5477 = ~n5496 | ~n7957;
  assign n5476 = ~n8005 | ~DATAO_REG_1__SCAN_IN;
  assign U3551 = ~n5477 | ~n5476;
  assign n5479 = ~n4906 | ~n7957;
  assign n5478 = ~n8000 | ~DATAO_REG_11__SCAN_IN;
  assign U3561 = ~n5479 | ~n5478;
  assign n5481 = ~n7583 | ~n7957;
  assign n5480 = ~n8005 | ~DATAO_REG_5__SCAN_IN;
  assign U3555 = ~n5481 | ~n5480;
  assign n5483 = ~n7680 | ~n7957;
  assign n5482 = ~n8005 | ~DATAO_REG_2__SCAN_IN;
  assign U3552 = ~n5483 | ~n5482;
  assign n5485 = ~n7314 | ~U4043;
  assign n5484 = ~n8000 | ~DATAO_REG_13__SCAN_IN;
  assign U3563 = ~n5485 | ~n5484;
  assign n5487 = ~n6840 | ~U4043;
  assign n5486 = ~n8000 | ~DATAO_REG_9__SCAN_IN;
  assign U3559 = ~n5487 | ~n5486;
  assign n5489 = ~n7316 | ~U4043;
  assign n5488 = ~n8000 | ~DATAO_REG_15__SCAN_IN;
  assign U3565 = ~n5489 | ~n5488;
  assign n5491 = ~n7351 | ~U4043;
  assign n5490 = ~n8000 | ~DATAO_REG_14__SCAN_IN;
  assign U3564 = ~n5491 | ~n5490;
  assign n5493 = ~n7486 | ~U4043;
  assign n5492 = ~n8005 | ~DATAO_REG_7__SCAN_IN;
  assign U3557 = ~n5493 | ~n5492;
  assign n5495 = ~n5267 | ~STATE_REG_SCAN_IN;
  assign n5494 = ~DATAI_20_ | ~U3149;
  assign U3332 = ~n5495 | ~n5494;
  assign n6133 = ~n5496 | ~n7670;
  assign n6137 = ~n5581 | ~n7652;
  assign n6141 = ~n7680 | ~n5567;
  assign n5497 = ~n7646 | ~n5577;
  assign n7582 = ~n7651;
  assign n6140 = ~n7651 | ~n7629;
  assign n6147 = ~n7617 | ~n7599;
  assign n5499 = ~n7560;
  assign n7557 = n7583 & n7563;
  assign n5588 = ~n7583;
  assign n7558 = ~n5588 | ~n7571;
  assign n6112 = ~n7486 | ~n7514;
  assign n5501 = ~n6112;
  assign n7496 = ~n7574 | ~n7534;
  assign n7532 = ~n7486;
  assign n5595 = ~n7532 | ~n7504;
  assign n5500 = n7496 & n5595;
  assign n6158 = n7451 | n7468;
  assign n5503 = ~n5502;
  assign n7495 = ~n7503 | ~n7529;
  assign n7473 = n7495 & n6112;
  assign n6113 = ~n7451 | ~n7468;
  assign n6159 = ~n6840 | ~n6921;
  assign n6157 = ~n7470 | ~n7452;
  assign n6120 = ~n7393 | ~n5602;
  assign n5504 = ~n7427 | ~n6120;
  assign n6118 = ~n7450 | ~n4886;
  assign n7339 = ~n5504 | ~n6118;
  assign n7344 = ~n7394 | ~n7379;
  assign n5505 = ~n7314 | ~n7330;
  assign n6129 = ~n7344 | ~n5505;
  assign n5506 = ~n6129 & ~n5606;
  assign n5992 = ~n7339 | ~n5506;
  assign n5607 = ~n4906;
  assign n7341 = ~n5607 | ~n7405;
  assign n7350 = ~n7394;
  assign n7343 = ~n7350 | ~n7368;
  assign n5508 = ~n7341 | ~n7343;
  assign n5507 = ~n6129;
  assign n5510 = ~n5508 | ~n5507;
  assign n7367 = ~n7314;
  assign n5509 = ~n7367 | ~n7352;
  assign n5993 = n5510 & n5509;
  assign n7310 = ~n5992 | ~n5993;
  assign n5997 = ~n7351 | ~n5610;
  assign n6597 = ~n7316;
  assign n5999 = ~n6597 | ~n5609;
  assign n5998 = ~n7316 | ~n6732;
  assign n6740 = ~n5999 | ~n5998;
  assign n5511 = ~n6740;
  assign n6594 = ~n5512 | ~n5998;
  assign n6179 = ~n7958 & ~n6610;
  assign n6502 = n7961 & n5902;
  assign n6084 = n5969 | n6517;
  assign n6504 = ~n7964 | ~n5972;
  assign n6002 = ~n6084 | ~n6504;
  assign n6477 = n6502 | n6002;
  assign n6168 = n7970 & n6489;
  assign n6376 = n6477 | n6168;
  assign n6398 = ~n5815;
  assign n6070 = ~n6345 & ~n6398;
  assign n5625 = ~n7976 | ~n6419;
  assign n5513 = ~n5625;
  assign n6111 = ~n6070 & ~n5513;
  assign n6387 = ~n7976;
  assign n6381 = ~n6387 | ~n6410;
  assign n6167 = n7973 & n6448;
  assign n5514 = ~n6381 | ~n6167;
  assign n6010 = ~n6111 | ~n5514;
  assign n6069 = ~n6345 | ~n6398;
  assign n6356 = ~n5920;
  assign n6063 = ~n6315 | ~n6356;
  assign n6187 = ~n6069 | ~n6063;
  assign n5518 = ~n6187;
  assign n6466 = ~n7973;
  assign n6379 = ~n6466 | ~n6437;
  assign n6008 = ~n6381 | ~n6379;
  assign n6181 = ~n6008;
  assign n6537 = ~n7961;
  assign n6531 = ~n6537 | ~n6583;
  assign n5898 = ~n7964;
  assign n5633 = ~n5898 | ~n6543;
  assign n6503 = n6531 & n5633;
  assign n5515 = n6002 | n6503;
  assign n6083 = ~n5969 | ~n6517;
  assign n6478 = n5515 & n6083;
  assign n5516 = n6168 | n6478;
  assign n6436 = ~n7970;
  assign n6005 = ~n6436 | ~n5621;
  assign n6377 = n5516 & n6005;
  assign n5517 = n6181 & n6377;
  assign n6339 = n6010 | n5517;
  assign n5519 = n5518 & n6339;
  assign n6310 = ~n7982 | ~n5920;
  assign n6053 = ~n7985 | ~n6330;
  assign n6188 = ~n6310 | ~n6053;
  assign n5722 = ~n7988;
  assign n6298 = ~n6020 | ~DATAI_26_;
  assign n6286 = ~n6298;
  assign n5520 = ~n5722 | ~n6286;
  assign n6280 = n7985 | n6330;
  assign n6191 = ~n5520 | ~n6280;
  assign n5724 = ~REG3_REG_27__SCAN_IN;
  assign n6264 = n5532 ^ ~n5724;
  assign n5529 = ~n6264 | ~n4760;
  assign n5523 = ~n5188 | ~REG0_REG_27__SCAN_IN;
  assign n5522 = ~n4359 | ~REG2_REG_27__SCAN_IN;
  assign n5527 = ~n5523 | ~n5522;
  assign n5524 = ~REG1_REG_27__SCAN_IN;
  assign n5526 = ~n5525 & ~n5524;
  assign n5528 = ~n5527 & ~n5526;
  assign n7991 = ~n5529 | ~n5528;
  assign n6258 = ~n6020 | ~DATAI_27_;
  assign n6049 = n7991 & n6258;
  assign n6254 = ~n5722 & ~n6286;
  assign n6195 = ~n6049 & ~n6254;
  assign n6050 = n7991 | n6258;
  assign n6034 = ~n6195 | ~n6050;
  assign n5531 = ~n6015 | ~REG1_REG_28__SCAN_IN;
  assign n5530 = ~n5188 | ~REG0_REG_28__SCAN_IN;
  assign n5540 = n5531 & n5530;
  assign n5534 = ~REG3_REG_28__SCAN_IN;
  assign n5533 = ~n5535;
  assign n5536 = ~n5534 | ~n5533;
  assign n5684 = ~REG3_REG_28__SCAN_IN | ~n5535;
  assign n5789 = ~n5536 | ~n5684;
  assign n5538 = n5544 | n5789;
  assign n6248 = ~REG2_REG_28__SCAN_IN;
  assign n5537 = n4682 | n6248;
  assign n5539 = n5538 & n5537;
  assign n7994 = ~n5540 | ~n5539;
  assign n5790 = ~n6020 | ~DATAI_28_;
  assign n5664 = n7994 & n5790;
  assign n5663 = ~n7994 & ~n5790;
  assign n5550 = ~n5541 & ~n5663;
  assign n5543 = ~n4890 | ~REG0_REG_29__SCAN_IN;
  assign n5542 = ~n4891 | ~REG2_REG_29__SCAN_IN;
  assign n5548 = n5543 & n5542;
  assign n5546 = ~n6015 | ~REG1_REG_29__SCAN_IN;
  assign n5545 = n5544 | n5684;
  assign n5547 = n5546 & n5545;
  assign n6030 = ~n6020 | ~DATAI_29_;
  assign n6052 = n6023 ^ ~n6030;
  assign n5553 = n5550 ^ ~n5549;
  assign n5552 = ~n5267 | ~n6131;
  assign n5551 = n7516 | n5666;
  assign n7678 = ~n5552 | ~n5551;
  assign n5566 = ~n5553 | ~n7678;
  assign n5555 = ~n4359 | ~REG2_REG_30__SCAN_IN;
  assign n5554 = ~n6015 | ~REG1_REG_30__SCAN_IN;
  assign n5557 = n5555 & n5554;
  assign n5556 = ~n5188 | ~REG0_REG_30__SCAN_IN;
  assign n8001 = n5557 & n5556;
  assign n5559 = ~n7067 | ~B_REG_SCAN_IN;
  assign n6223 = ~n7709 | ~n5559;
  assign n5564 = ~n8001 & ~n6223;
  assign n7668 = n7069 | n5560;
  assign n7533 = ~n7668;
  assign n5562 = ~n7994 | ~n7533;
  assign n6022 = ~n6030;
  assign n5561 = ~n7714 | ~n6022;
  assign n5563 = ~n5562 | ~n5561;
  assign n5565 = ~n5564 & ~n5563;
  assign n5687 = ~n5566 | ~n5565;
  assign n5569 = n5568 & n5567;
  assign n7641 = ~n5569 | ~n7670;
  assign n7570 = ~n7598 | ~n7599;
  assign n5571 = n7379 & n6954;
  assign n6582 = ~n6611 | ~n6610;
  assign n6397 = n6419 & n6448;
  assign n5573 = n5815 & n6397;
  assign n6273 = ~n6258;
  assign n5779 = ~n5790;
  assign n6231 = ~n5574 | ~n6030;
  assign n5575 = n5574 | n6030;
  assign n5683 = ~n6231 | ~n5575;
  assign n5576 = ~n5683 & ~n7858;
  assign n5669 = ~n5687 & ~n5576;
  assign n5580 = ~n5577;
  assign n7683 = n6854 & n5578;
  assign n7685 = ~n7684 | ~n7683;
  assign n5579 = ~n5496 | ~n4729;
  assign n5582 = ~n5581 | ~n5567;
  assign n5583 = ~n7582 | ~n7629;
  assign n5585 = ~n7612 | ~n5583;
  assign n5584 = ~n7651 | ~n7618;
  assign n7591 = ~n5585 | ~n5584;
  assign n7592 = ~n4377 | ~n6147;
  assign n5587 = ~n7591 | ~n7592;
  assign n5586 = ~n7617 | ~n7584;
  assign n7556 = ~n5587 | ~n5586;
  assign n5589 = ~n5588 | ~n7563;
  assign n5591 = ~n7556 | ~n5589;
  assign n5590 = ~n7583 | ~n7571;
  assign n7526 = ~n5591 | ~n5590;
  assign n5592 = ~n7574 | ~n7529;
  assign n5594 = ~n7526 | ~n5592;
  assign n5593 = ~n7503 | ~n7534;
  assign n7511 = ~n5594 | ~n5593;
  assign n5597 = ~n7511 | ~n6152;
  assign n5596 = ~n7486 | ~n7504;
  assign n7478 = ~n5597 | ~n5596;
  assign n7502 = ~n7451;
  assign n5598 = ~n7502 | ~n7468;
  assign n5599 = ~n7451 | ~n7471;
  assign n5600 = ~n7470 | ~n6921;
  assign n5601 = ~n6840 | ~n7452;
  assign n5603 = ~n7450 | ~n5602;
  assign n5605 = ~n7415 | ~n5603;
  assign n5604 = ~n7393 | ~n4886;
  assign n7340 = ~n5606;
  assign n5608 = ~n5607 | ~n6954;
  assign n6587 = ~n7394 & ~n7368;
  assign n5636 = ~n7958 | ~n6598;
  assign n5620 = ~n5636;
  assign n5614 = ~n7316 | ~n5609;
  assign n5611 = n7316 | n5609;
  assign n6738 = ~n6725 | ~n5610;
  assign n5612 = ~n5611 | ~n6738;
  assign n5616 = ~n5614 | ~n5612;
  assign n6736 = ~n7314 | ~n7352;
  assign n5613 = ~n6736;
  assign n6735 = ~n7367 | ~n7330;
  assign n6590 = n6735 & n5616;
  assign n5617 = n6590 & n6595;
  assign n5634 = n6537 & n5902;
  assign n6458 = ~n5898 | ~n5972;
  assign n6460 = ~n5969 | ~n5826;
  assign n5644 = ~n6458 | ~n6460;
  assign n6462 = ~n7970 | ~n5621;
  assign n6459 = n5969 | n5826;
  assign n6367 = n6462 & n6459;
  assign n5626 = ~n6345 | ~n5815;
  assign n5624 = ~n5626;
  assign n5622 = ~n7979 | ~n6398;
  assign n6374 = ~n7976 | ~n6410;
  assign n5623 = n5622 & n6374;
  assign n5629 = ~n5630;
  assign n6428 = n6381 & n5625;
  assign n6373 = ~n6428;
  assign n5627 = n6373 & n5626;
  assign n6371 = ~n6466 | ~n6448;
  assign n5628 = n5627 & n6371;
  assign n5649 = n5629 | n5628;
  assign n5632 = ~n5649;
  assign n6370 = ~n7973 | ~n6437;
  assign n5631 = n6370 & n5630;
  assign n5648 = n5632 | n5631;
  assign n6334 = n6367 & n5648;
  assign n5647 = ~n7982 | ~n6356;
  assign n5645 = n6334 & n5647;
  assign n5641 = ~n5634;
  assign n6588 = ~n7394 | ~n7368;
  assign n5637 = n6588 & n5635;
  assign n5638 = n5637 & n5636;
  assign n5640 = ~n6562;
  assign n5643 = ~n5641 | ~n5640;
  assign n5642 = ~n7961 | ~n6583;
  assign n5656 = ~n6333 | ~n5646;
  assign n5652 = ~n5647;
  assign n5651 = ~n5648;
  assign n6461 = ~n6436 | ~n6489;
  assign n5650 = n6461 & n5649;
  assign n5654 = n5652 | n6335;
  assign n5653 = ~n6315 | ~n5920;
  assign n5655 = n5654 & n5653;
  assign n5658 = ~n7985 | ~n5657;
  assign n5917 = ~n7985;
  assign n5659 = ~n5722 | ~n6298;
  assign n6267 = ~n5660 | ~n5659;
  assign n5661 = ~n7991 | ~n6273;
  assign n6285 = ~n7991;
  assign n5662 = ~n6285 | ~n6258;
  assign n6014 = ~n5663;
  assign n6032 = ~n5664;
  assign n5723 = ~n7994;
  assign n5667 = n5688 ^ ~n5666;
  assign n7887 = ~n7707 | ~n7901;
  assign n5668 = ~n5689 | ~n7887;
  assign n5768 = ~n5669 | ~n5668;
  assign n5671 = ~n5670;
  assign n5673 = ~n5671 | ~n5680;
  assign n5675 = ~n5673 & ~n5672;
  assign n5767 = ~n5675 | ~n5674;
  assign n5676 = ~n5766;
  assign n7952 = n5767 | n5676;
  assign n7954 = ~n7952;
  assign n5678 = ~n5768 | ~n7954;
  assign n5677 = ~n7952 | ~REG1_REG_29__SCAN_IN;
  assign U3547 = ~n5678 | ~n5677;
  assign n5681 = ~n5680 | ~n5679;
  assign n7608 = ~n5682 | ~n7632;
  assign n7418 = ~n7572;
  assign n7642 = ~n7608 | ~n7418;
  assign n5685 = n5683 | n7642;
  assign n5686 = ~n7608 | ~n4596;
  assign n5691 = ~n4589 | ~n4597;
  assign n7698 = ~n7608;
  assign n7691 = n5688 | n7516;
  assign n6244 = n7707 & n7691;
  assign n6528 = ~n7698 & ~n6244;
  assign n5690 = ~n5689 | ~n6528;
  assign U3354 = ~n5691 | ~n5690;
  assign n5693 = ~n7988 | ~n4362;
  assign n5692 = n5774 | n6298;
  assign n5694 = ~n5693 | ~n5692;
  assign n5710 = n5694 ^ ~n4711;
  assign n5696 = ~n7988 | ~n5778;
  assign n5695 = ~n4934 | ~n6286;
  assign n5709 = ~n5696 | ~n5695;
  assign n5739 = n5710 | n5709;
  assign n5715 = n5697 & n5739;
  assign n5699 = ~n7991 | ~n4362;
  assign n5698 = n5774 | n6258;
  assign n5701 = ~n5699 | ~n5698;
  assign n5705 = n5701 ^ ~n5700;
  assign n5703 = ~n7991 | ~n5778;
  assign n5702 = ~n4362 | ~n6273;
  assign n5704 = n5703 & n5702;
  assign n5786 = n5705 | n5704;
  assign n5706 = ~n5705 | ~n5704;
  assign n5717 = ~n5786 | ~n5706;
  assign n5707 = ~n5717;
  assign n5708 = n5715 & n5707;
  assign n5714 = ~n5736 | ~n5708;
  assign n5712 = ~n5739;
  assign n5738 = n5710 & n5709;
  assign n5711 = ~n5738 & ~n5735;
  assign n5716 = n5712 | n5711;
  assign n5713 = n5717 | n5716;
  assign n5719 = ~n5736 | ~n5715;
  assign n5718 = n5717 & n5716;
  assign n5720 = ~n5719 | ~n5718;
  assign n5721 = ~n5720 | ~n6970;
  assign n5734 = ~n5804 & ~n5721;
  assign n5730 = ~n5722 & ~n6955;
  assign n5728 = ~n6990 | ~n6273;
  assign n5726 = ~n6951 & ~n5723;
  assign n5725 = ~n5724 & ~STATE_REG_SCAN_IN;
  assign n5727 = ~n5726 & ~n5725;
  assign n5729 = ~n5728 | ~n5727;
  assign n5732 = ~n5730 & ~n5729;
  assign n5731 = ~n6264 | ~n6798;
  assign n5733 = ~n5732 | ~n5731;
  assign U3211 = n5734 | n5733;
  assign n5740 = ~n5738;
  assign n5751 = ~n5741 | ~n6970;
  assign n5749 = ~n6285 & ~n6951;
  assign n5747 = ~n6301 | ~n6798;
  assign n5745 = ~n6974 & ~n6298;
  assign n5743 = n6955 | n5917;
  assign n5742 = ~REG3_REG_26__SCAN_IN | ~U3149;
  assign n5744 = ~n5743 | ~n5742;
  assign n5746 = ~n5745 & ~n5744;
  assign n5748 = ~n5747 | ~n5746;
  assign n5750 = ~n5749 & ~n5748;
  assign U3237 = ~n5751 | ~n5750;
  assign n5753 = n6102 ^ n5752;
  assign n5759 = ~n5753 | ~n7678;
  assign n5757 = ~n6285 & ~n7668;
  assign n7997 = ~n6023;
  assign n5755 = ~n7997 | ~n7709;
  assign n5754 = ~n7714 | ~n5779;
  assign n5756 = ~n5755 | ~n5754;
  assign n5758 = ~n5757 & ~n5756;
  assign n6243 = ~n5759 | ~n5758;
  assign n5760 = n6275 ^ ~n5779;
  assign n6240 = ~n5760 & ~n7858;
  assign n5763 = ~n6243 & ~n6240;
  assign n6245 = n6102 ^ n5761;
  assign n5762 = ~n6245 | ~n7887;
  assign n5771 = ~n5763 | ~n5762;
  assign n5765 = ~n5771 | ~n7954;
  assign n5764 = ~n7952 | ~REG1_REG_28__SCAN_IN;
  assign U3546 = ~n5765 | ~n5764;
  assign n7900 = n5767 | n5766;
  assign n7907 = ~n7900;
  assign n5770 = ~n5768 | ~n7907;
  assign n5769 = ~n7900 | ~REG0_REG_29__SCAN_IN;
  assign U3515 = ~n5770 | ~n5769;
  assign n5773 = ~n5771 | ~n7907;
  assign n5772 = ~n7900 | ~REG0_REG_28__SCAN_IN;
  assign U3514 = ~n5773 | ~n5772;
  assign n5776 = ~n7994 | ~n4934;
  assign n5775 = n5774 | n5790;
  assign n5777 = ~n5776 | ~n5775;
  assign n5783 = n5777 ^ ~n4711;
  assign n5781 = ~n5778 | ~n7994;
  assign n5780 = ~n4362 | ~n5779;
  assign n5782 = ~n5781 | ~n5780;
  assign n5787 = n5783 ^ ~n5782;
  assign n5784 = ~n5787 & ~n7007;
  assign n5785 = ~n5786 | ~n5784;
  assign n5788 = ~n5786;
  assign n5803 = n5787 & n6970;
  assign n5800 = ~n5788 | ~n5803;
  assign n5798 = ~n6285 & ~n6955;
  assign n6251 = ~n5789;
  assign n5796 = ~n6798 | ~n6251;
  assign n5794 = ~n6974 & ~n5790;
  assign n5792 = n6951 | n6023;
  assign n5791 = ~REG3_REG_28__SCAN_IN | ~U3149;
  assign n5793 = ~n5792 | ~n5791;
  assign n5795 = ~n5794 & ~n5793;
  assign n5797 = ~n5796 | ~n5795;
  assign n5799 = ~n5798 & ~n5797;
  assign n5801 = ~n5800 | ~n5799;
  assign n5806 = ~n5802 & ~n5801;
  assign n5805 = ~n5804 | ~n5803;
  assign U3217 = ~n5806 | ~n5805;
  assign n5809 = n5808 ^ ~n5807;
  assign n5821 = ~n5809 & ~n7007;
  assign n5810 = ~n6399;
  assign n5819 = ~n6798 | ~n5810;
  assign n5812 = n6955 | n6387;
  assign n5811 = ~REG3_REG_23__SCAN_IN | ~U3149;
  assign n5814 = ~n5812 | ~n5811;
  assign n5813 = ~n6951 & ~n6315;
  assign n5817 = ~n5814 & ~n5813;
  assign n5816 = n6974 | n5815;
  assign n5818 = n5817 & n5816;
  assign n5820 = ~n5819 | ~n5818;
  assign U3213 = n5821 | n5820;
  assign n5824 = n4380 & n5823;
  assign n5825 = ~n5822 & ~n5824;
  assign n5836 = ~n5825 & ~n7007;
  assign n5834 = ~n6798 | ~n6521;
  assign n5830 = ~n6955 & ~n5898;
  assign n5827 = ~n5826 & ~n6974;
  assign n5829 = n5828 | n5827;
  assign n5832 = ~n5830 & ~n5829;
  assign n5831 = ~n7970 | ~n6991;
  assign n5833 = n5832 & n5831;
  assign n5835 = ~n5834 | ~n5833;
  assign U3216 = n5836 | n5835;
  assign n5838 = ~n5929 | ~n5927;
  assign n5928 = ~n5837;
  assign n5842 = ~n5838 | ~n5928;
  assign n5841 = n5840 ^ ~n5839;
  assign n5843 = n5842 ^ ~n5841;
  assign n5854 = ~n5843 | ~n6970;
  assign n6449 = ~n5844;
  assign n5852 = n6798 & n6449;
  assign n5848 = ~n6974 & ~n6448;
  assign n5846 = n6951 | n6387;
  assign n5845 = ~REG3_REG_21__SCAN_IN | ~U3149;
  assign n5847 = ~n5846 | ~n5845;
  assign n5850 = ~n5848 & ~n5847;
  assign n5849 = ~n7970 | ~n6988;
  assign n5851 = ~n5850 | ~n5849;
  assign n5853 = ~n5852 & ~n5851;
  assign U3220 = ~n5854 | ~n5853;
  assign n5857 = ~n5855 | ~n6796;
  assign n6847 = ~n5857 | ~n5856;
  assign n5858 = ~n6847 | ~n6845;
  assign n6938 = ~n5858 | ~n6846;
  assign n5861 = n6938 | n5859;
  assign n6935 = ~n5861 | ~n5860;
  assign n6808 = ~n6935 & ~n6941;
  assign n6809 = ~n5862 | ~n5863;
  assign n5865 = ~n6808 & ~n6809;
  assign n5864 = ~n5863;
  assign n5866 = ~n5865 & ~n5864;
  assign n5870 = ~n5866 | ~n5867;
  assign n5869 = ~n5866;
  assign n5868 = ~n5867;
  assign n5871 = ~n5869 | ~n5868;
  assign n5979 = ~n5870 | ~n5871;
  assign n5873 = ~n5979 & ~n5980;
  assign n5872 = ~n5871;
  assign n5874 = ~n5873 & ~n5872;
  assign n5876 = n5875 ^ n5874;
  assign n5886 = ~n5876 & ~n7007;
  assign n6613 = ~n5877;
  assign n5884 = ~n6798 | ~n6613;
  assign n5878 = n6955 | n6597;
  assign n7245 = ~REG3_REG_16__SCAN_IN | ~U3149;
  assign n5880 = ~n5878 | ~n7245;
  assign n5879 = ~n6951 & ~n6537;
  assign n5882 = ~n5880 & ~n5879;
  assign n5881 = n6974 | n6610;
  assign n5883 = n5882 & n5881;
  assign n5885 = ~n5884 | ~n5883;
  assign U3223 = n5886 | n5885;
  assign n5888 = ~n5887;
  assign n5895 = ~n5888 & ~n5892;
  assign n5891 = ~n5890;
  assign n5893 = ~n5892 & ~n5891;
  assign n5894 = ~n5889 & ~n5893;
  assign n5896 = ~n5895 & ~n5894;
  assign n5908 = ~n5896 & ~n7007;
  assign n6574 = ~n5897;
  assign n5906 = ~n6798 | ~n6574;
  assign n5899 = n6951 | n5898;
  assign n7257 = ~REG3_REG_17__SCAN_IN | ~U3149;
  assign n5901 = ~n5899 | ~n7257;
  assign n6567 = ~n7958;
  assign n5900 = ~n6955 & ~n6567;
  assign n5904 = ~n5901 & ~n5900;
  assign n5903 = n6974 | n5902;
  assign n5905 = n5904 & n5903;
  assign n5907 = ~n5906 | ~n5905;
  assign U3225 = n5908 | n5907;
  assign n5912 = n5911 ^ ~n5910;
  assign n5913 = n5909 ^ ~n5912;
  assign n5926 = ~n5913 & ~n7007;
  assign n6360 = ~n5914;
  assign n5924 = ~n6798 | ~n6360;
  assign n5916 = n6955 | n6345;
  assign n5915 = ~REG3_REG_24__SCAN_IN | ~U3149;
  assign n5919 = ~n5916 | ~n5915;
  assign n5918 = ~n6951 & ~n5917;
  assign n5922 = ~n5919 & ~n5918;
  assign n5921 = n6974 | n5920;
  assign n5923 = n5922 & n5921;
  assign n5925 = ~n5924 | ~n5923;
  assign U3226 = n5926 | n5925;
  assign n5930 = ~n5928 | ~n5927;
  assign n5931 = n5930 ^ n5929;
  assign n5942 = ~n5931 & ~n7007;
  assign n5932 = ~n6495;
  assign n5940 = ~n6798 | ~n5932;
  assign n5934 = n6951 | n6466;
  assign n5933 = ~REG3_REG_20__SCAN_IN | ~U3149;
  assign n5936 = ~n5934 | ~n5933;
  assign n5935 = ~n6955 & ~n5969;
  assign n5938 = ~n5936 & ~n5935;
  assign n5937 = n6974 | n6489;
  assign n5939 = n5938 & n5937;
  assign n5941 = ~n5940 | ~n5939;
  assign U3230 = n5942 | n5941;
  assign n5946 = n5945 & n5944;
  assign n5947 = ~n5943 & ~n5946;
  assign n5958 = ~n5947 & ~n7007;
  assign n5948 = ~n6423;
  assign n5956 = ~n6798 | ~n5948;
  assign n5950 = n6951 | n6345;
  assign n5949 = ~U3149 | ~REG3_REG_22__SCAN_IN;
  assign n5952 = ~n5950 | ~n5949;
  assign n5951 = ~n6955 & ~n6466;
  assign n5954 = ~n5952 & ~n5951;
  assign n5953 = n6974 | n6419;
  assign n5955 = n5954 & n5953;
  assign n5957 = ~n5956 | ~n5955;
  assign U3232 = n5958 | n5957;
  assign n5965 = ~n4370 & ~n5960;
  assign n5963 = ~n5959;
  assign n5962 = ~n5961 & ~n5960;
  assign n5964 = ~n5963 & ~n5962;
  assign n5966 = ~n5965 & ~n5964;
  assign n5978 = ~n5966 & ~n7007;
  assign n6558 = ~n5967;
  assign n5976 = ~n6798 | ~n6558;
  assign n5968 = n6955 | n6537;
  assign n7272 = ~REG3_REG_18__SCAN_IN | ~U3149;
  assign n5971 = ~n5968 | ~n7272;
  assign n5970 = ~n6951 & ~n5969;
  assign n5974 = ~n5971 & ~n5970;
  assign n5973 = n6974 | n5972;
  assign n5975 = n5974 & n5973;
  assign n5977 = ~n5976 | ~n5975;
  assign U3235 = n5978 | n5977;
  assign n5981 = n5980 ^ n5979;
  assign n5991 = ~n5981 & ~n7007;
  assign n5982 = ~n7292;
  assign n5989 = ~n6798 | ~n5982;
  assign n5983 = n6955 | n6725;
  assign n7231 = ~REG3_REG_15__SCAN_IN | ~U3149;
  assign n5985 = ~n5983 | ~n7231;
  assign n5984 = ~n6951 & ~n6567;
  assign n5987 = ~n5985 & ~n5984;
  assign n5986 = n6974 | n6732;
  assign n5988 = n5987 & n5986;
  assign n5990 = ~n5989 | ~n5988;
  assign U3238 = n5991 | n5990;
  assign n5996 = ~n5993;
  assign n5995 = ~n5994 | ~n5999;
  assign n6124 = ~n5996 & ~n5995;
  assign n6000 = ~n5992 | ~n6124;
  assign n6127 = ~n5998 | ~n5997;
  assign n6125 = ~n6127 | ~n5999;
  assign n6001 = n6000 & n6125;
  assign n6004 = ~n6001 & ~n6179;
  assign n6169 = ~n6002 & ~n6502;
  assign n6003 = ~n6169 | ~n4410;
  assign n6006 = ~n6004 & ~n6003;
  assign n6173 = ~n6005 | ~n6478;
  assign n6007 = ~n6006 & ~n6173;
  assign n6009 = ~n6007 & ~n6168;
  assign n6011 = ~n6009 & ~n6008;
  assign n6012 = ~n6011 & ~n6010;
  assign n6013 = ~n6012 & ~n6187;
  assign n6029 = ~n6013 & ~n6188;
  assign n6035 = ~n6050 | ~n6014;
  assign n6027 = ~n6035;
  assign n6017 = ~n4359 | ~REG2_REG_31__SCAN_IN;
  assign n6016 = ~n6015 | ~REG1_REG_31__SCAN_IN;
  assign n6019 = n6017 & n6016;
  assign n6018 = ~n5188 | ~REG0_REG_31__SCAN_IN;
  assign n6224 = n6019 & n6018;
  assign n6225 = ~n6020 | ~DATAI_31_;
  assign n6043 = ~n6225;
  assign n6197 = ~n6224 & ~n6043;
  assign n6232 = n4771 & DATAI_30_;
  assign n6021 = n8001 & n6232;
  assign n6064 = ~n6197 & ~n6021;
  assign n6024 = ~n6023 | ~n6022;
  assign n6036 = n6064 & n6024;
  assign n6025 = ~n6036;
  assign n6026 = ~n6191 & ~n6025;
  assign n6028 = ~n6027 | ~n6026;
  assign n6040 = ~n6029 & ~n6028;
  assign n6031 = ~n7997 | ~n6030;
  assign n6110 = n6032 & n6031;
  assign n6033 = ~n6110;
  assign n6038 = ~n6034 & ~n6033;
  assign n6037 = ~n6035 | ~n6110;
  assign n6198 = ~n6037 | ~n6036;
  assign n6039 = ~n6038 & ~n6198;
  assign n6042 = ~n6040 & ~n6039;
  assign n8006 = ~n6224;
  assign n6233 = ~n6232;
  assign n6041 = ~n8006 & ~n6233;
  assign n6046 = ~n6042 & ~n6041;
  assign n6062 = ~n8001 & ~n6232;
  assign n6044 = ~n6062 | ~n6043;
  assign n6060 = ~n6224 | ~n6043;
  assign n6045 = ~n6044 | ~n6060;
  assign n6047 = ~n6046 & ~n6045;
  assign n6048 = n6047 ^ ~n7516;
  assign n6108 = ~n6048 | ~n6131;
  assign n6051 = ~n6049;
  assign n6268 = n6051 & n6050;
  assign n6101 = ~n6052 | ~n6268;
  assign n6282 = n7988 ^ ~n6298;
  assign n7426 = ~n6118 | ~n6120;
  assign n7448 = ~n6157 | ~n6159;
  assign n6058 = ~n7426 & ~n7448;
  assign n6312 = ~n6280 | ~n6053;
  assign n7479 = ~n6158 | ~n6113;
  assign n6055 = ~n7479;
  assign n6132 = ~n6854 | ~n5568;
  assign n6054 = ~n6132;
  assign n7787 = n7674 | n6054;
  assign n7703 = ~n7787;
  assign n6056 = ~n6055 | ~n7703;
  assign n6057 = ~n6312 & ~n6056;
  assign n6059 = ~n6058 | ~n6057;
  assign n6099 = ~n6282 & ~n6059;
  assign n6061 = ~n6060;
  assign n6196 = ~n6062 & ~n6061;
  assign n6342 = ~n6310 | ~n6063;
  assign n6065 = ~n6064;
  assign n6066 = ~n6342 & ~n6065;
  assign n6097 = ~n6196 | ~n6066;
  assign n6068 = ~n6152 & ~n7557;
  assign n7539 = ~n7496 | ~n7495;
  assign n6067 = ~n7539;
  assign n6072 = ~n6068 | ~n6067;
  assign n6340 = ~n6069;
  assign n6382 = ~n6070 & ~n6340;
  assign n6071 = ~n6428 | ~n6382;
  assign n6095 = ~n6072 & ~n6071;
  assign n6076 = ~n6073 | ~n7398;
  assign n6075 = ~n5577 | ~n6074;
  assign n6081 = ~n6076 & ~n6075;
  assign n6077 = ~n7592;
  assign n6079 = ~n6077 | ~n7309;
  assign n6078 = ~n6549 | ~n7558;
  assign n6080 = ~n6079 & ~n6078;
  assign n6093 = ~n6081 | ~n6080;
  assign n6082 = ~n6167;
  assign n6433 = n6082 & n6379;
  assign n6499 = ~n6461 | ~n6462;
  assign n6089 = ~n6433 | ~n6499;
  assign n6526 = ~n6084 | ~n6083;
  assign n6085 = ~n6502;
  assign n6565 = ~n6085 | ~n6531;
  assign n6087 = ~n6526 & ~n6565;
  assign n7347 = n7314 ^ ~n7330;
  assign n7375 = ~n7343 | ~n7344;
  assign n6086 = ~n7347 & ~n7375;
  assign n6088 = ~n6087 | ~n6086;
  assign n6091 = ~n6089 & ~n6088;
  assign n7614 = ~n7611;
  assign n6090 = ~n7614 & ~n6740;
  assign n6092 = ~n6091 | ~n6090;
  assign n6094 = ~n6093 & ~n6092;
  assign n6096 = ~n6095 | ~n6094;
  assign n6098 = ~n6097 & ~n6096;
  assign n6100 = ~n6099 | ~n6098;
  assign n6103 = ~n6101 & ~n6100;
  assign n6104 = ~n6103 | ~n6102;
  assign n6106 = n6104 ^ ~n7712;
  assign n6107 = ~n6106 | ~n6105;
  assign n6109 = ~n6108 | ~n6107;
  assign n6206 = ~n6109 | ~n5267;
  assign n6193 = ~n6110 | ~n6196;
  assign n6185 = ~n6111;
  assign n6115 = ~n6159;
  assign n6114 = ~n6113 | ~n6112;
  assign n6155 = ~n6115 & ~n6114;
  assign n6116 = ~n7495;
  assign n6117 = ~n6116 & ~n7558;
  assign n6119 = ~n6155 | ~n6117;
  assign n6122 = ~n6119 | ~n6118;
  assign n6128 = ~n7340 | ~n6120;
  assign n6121 = ~n6128 & ~n6129;
  assign n6123 = ~n6122 | ~n6121;
  assign n6126 = ~n6124 | ~n6123;
  assign n6166 = ~n6126 | ~n6125;
  assign n6130 = n6128 | n6127;
  assign n6164 = ~n6130 & ~n6129;
  assign n6135 = ~n7674 & ~n6131;
  assign n6134 = ~n6133 | ~n6132;
  assign n6139 = ~n6135 & ~n6134;
  assign n6138 = ~n6137 | ~n6136;
  assign n6143 = ~n6139 & ~n6138;
  assign n6142 = ~n6141 | ~n6140;
  assign n6146 = ~n6143 & ~n6142;
  assign n6145 = ~n4377 | ~n6144;
  assign n6150 = n6146 | n6145;
  assign n6148 = ~n7495 | ~n6147;
  assign n6149 = ~n6148 & ~n7557;
  assign n6154 = ~n6150 | ~n6149;
  assign n6151 = ~n7496;
  assign n6153 = ~n6152 & ~n6151;
  assign n6156 = ~n6154 | ~n6153;
  assign n6162 = ~n6156 | ~n6155;
  assign n6160 = ~n6158 | ~n6157;
  assign n6161 = ~n6160 | ~n6159;
  assign n6163 = ~n6162 | ~n6161;
  assign n6165 = ~n6164 | ~n6163;
  assign n6172 = ~n6166 | ~n6165;
  assign n6174 = ~n6168 & ~n6167;
  assign n6177 = ~n6169 | ~n6174;
  assign n6171 = ~n6170 & ~n6177;
  assign n6176 = ~n6172 | ~n6171;
  assign n6175 = ~n6174 | ~n6173;
  assign n6183 = ~n6176 | ~n6175;
  assign n6178 = ~n6177;
  assign n6180 = ~n6179 | ~n6178;
  assign n6182 = ~n6181 | ~n6180;
  assign n6184 = ~n6183 & ~n6182;
  assign n6186 = ~n6185 & ~n6184;
  assign n6189 = ~n6187 & ~n6186;
  assign n6190 = ~n6189 & ~n6188;
  assign n6192 = ~n6191 & ~n6190;
  assign n6194 = ~n6193 & ~n6192;
  assign n6201 = ~n6195 | ~n6194;
  assign n6199 = n6197 | n6196;
  assign n6200 = ~n6199 | ~n6198;
  assign n6202 = ~n6201 | ~n6200;
  assign n6204 = n6202 ^ ~n7516;
  assign n6205 = ~n6204 | ~n6203;
  assign n6208 = ~n6206 | ~n6205;
  assign n6207 = ~n6213;
  assign n6222 = ~n6208 | ~n6207;
  assign n6210 = ~n7058 & ~n6209;
  assign n6211 = ~n6210 | ~n7516;
  assign n6212 = ~n7069 & ~n6211;
  assign n6214 = ~n4934 | ~n6212;
  assign n6219 = ~n6214 | ~n6213;
  assign n6217 = ~n6215;
  assign n6218 = ~n6217 | ~n6216;
  assign n6220 = ~n6219 | ~n6218;
  assign n6221 = ~n6220 | ~B_REG_SCAN_IN;
  assign U3239 = ~n6222 | ~n6221;
  assign n7665 = ~n7642;
  assign n6230 = ~n6620 | ~n7665;
  assign n6235 = ~n6224 & ~n6223;
  assign n6226 = ~n7671 & ~n6225;
  assign n6621 = ~n6235 & ~n6226;
  assign n6228 = ~n6621 | ~n7608;
  assign n6227 = n7608 | REG2_REG_31__SCAN_IN;
  assign n6229 = ~n6228 | ~n6227;
  assign U3260 = ~n6230 | ~n6229;
  assign n6624 = n6232 ^ n6231;
  assign n6239 = ~n6624 | ~n7665;
  assign n6234 = ~n7671 & ~n6233;
  assign n6625 = ~n6235 & ~n6234;
  assign n6237 = ~n6625 | ~n7608;
  assign n6236 = n7608 | REG2_REG_30__SCAN_IN;
  assign n6238 = ~n6237 | ~n6236;
  assign U3261 = ~n6239 | ~n6238;
  assign n6241 = ~n6240 | ~n7516;
  assign n6242 = ~n6241 | ~n7608;
  assign n6247 = ~n6243 & ~n6242;
  assign n7513 = ~n6244;
  assign n6246 = ~n6245 | ~n7513;
  assign n6250 = ~n6247 | ~n6246;
  assign n6249 = ~n7698 | ~n6248;
  assign n6253 = ~n6250 | ~n6249;
  assign n7699 = ~n7632;
  assign n6252 = ~n7699 | ~n6251;
  assign U3262 = ~n6253 | ~n6252;
  assign n6257 = ~n6255 & ~n6268;
  assign n6262 = ~n7988 | ~n7533;
  assign n6260 = ~n7994 | ~n7709;
  assign n6259 = n7671 | n6258;
  assign n6261 = n6260 & n6259;
  assign n6263 = ~n6262 | ~n6261;
  assign n6265 = ~n6264 | ~n7699;
  assign n6266 = ~n6265 | ~n7608;
  assign n6270 = ~n6631 & ~n6266;
  assign n6632 = n6268 ^ n6267;
  assign n6269 = ~n6632 | ~n7513;
  assign n6272 = ~n6270 | ~n6269;
  assign n6271 = n7608 | REG2_REG_27__SCAN_IN;
  assign n6277 = ~n6272 | ~n6271;
  assign n6274 = ~n4366 | ~n6273;
  assign n6629 = ~n6275 | ~n6274;
  assign n6276 = n6629 | n7642;
  assign U3263 = ~n6277 | ~n6276;
  assign n6637 = n6282 ^ n6278;
  assign n6294 = ~n6637 & ~n7707;
  assign n6281 = ~n6280;
  assign n6283 = ~n6279 & ~n6281;
  assign n6284 = n6283 ^ ~n6282;
  assign n6292 = ~n6284 | ~n7678;
  assign n7573 = ~n7709;
  assign n6290 = ~n6285 & ~n7573;
  assign n6288 = ~n7985 | ~n7533;
  assign n6287 = ~n7714 | ~n6286;
  assign n6289 = ~n6288 | ~n6287;
  assign n6291 = ~n6290 & ~n6289;
  assign n6293 = ~n6292 | ~n6291;
  assign n6642 = ~n6294 & ~n6293;
  assign n6297 = ~n6642 | ~n7608;
  assign n6296 = ~n7698 | ~n6295;
  assign n6307 = ~n6297 | ~n6296;
  assign n7613 = ~n7691;
  assign n7702 = ~n7608 | ~n7613;
  assign n6305 = ~n6637 & ~n7702;
  assign n6300 = n6299 | n6298;
  assign n6638 = ~n6300 | ~n4366;
  assign n6303 = n6638 | n7642;
  assign n6302 = ~n6301 | ~n7699;
  assign n6304 = ~n6303 | ~n6302;
  assign n6306 = ~n6305 & ~n6304;
  assign U3264 = ~n6307 | ~n6306;
  assign n6645 = n6308 ^ ~n6312;
  assign n6326 = ~n6645 | ~n7513;
  assign n6311 = ~n6310;
  assign n6313 = ~n6309 & ~n6311;
  assign n6314 = n6313 ^ ~n6312;
  assign n6321 = ~n6314 & ~n7706;
  assign n6319 = ~n7988 | ~n7709;
  assign n6317 = ~n6315 & ~n7668;
  assign n6316 = ~n7671 & ~n6330;
  assign n6318 = ~n6317 & ~n6316;
  assign n6320 = ~n6319 | ~n6318;
  assign n6648 = n6321 | n6320;
  assign n6323 = ~n7699 | ~n6322;
  assign n6324 = ~n7608 | ~n6323;
  assign n6325 = ~n6648 & ~n6324;
  assign n6328 = ~n6326 | ~n6325;
  assign n6327 = n7608 | REG2_REG_25__SCAN_IN;
  assign n6332 = ~n6328 | ~n6327;
  assign n6646 = n6329 ^ ~n6330;
  assign n6331 = n6646 | n7642;
  assign U3265 = ~n6332 | ~n6331;
  assign n6336 = ~n6368 | ~n6334;
  assign n6337 = ~n6336 | ~n6335;
  assign n6653 = n6342 ^ n6337;
  assign n6353 = ~n6653 & ~n7707;
  assign n6341 = ~n6338 | ~n6339;
  assign n6343 = ~n6341 & ~n6340;
  assign n6344 = n6343 ^ ~n6342;
  assign n6351 = ~n6344 | ~n7678;
  assign n6349 = ~n6345 & ~n7668;
  assign n6347 = ~n7985 | ~n7709;
  assign n6346 = ~n7714 | ~n6356;
  assign n6348 = ~n6347 | ~n6346;
  assign n6350 = ~n6349 & ~n6348;
  assign n6352 = ~n6351 | ~n6350;
  assign n6658 = ~n6353 & ~n6352;
  assign n6355 = ~n6658 | ~n7608;
  assign n6354 = n7608 | REG2_REG_24__SCAN_IN;
  assign n6366 = ~n6355 | ~n6354;
  assign n6364 = ~n6653 & ~n7702;
  assign n6359 = ~n6329;
  assign n6358 = ~n6357 | ~n6356;
  assign n6654 = ~n6359 | ~n6358;
  assign n6362 = n6654 | n7642;
  assign n6361 = ~n7699 | ~n6360;
  assign n6363 = ~n6362 | ~n6361;
  assign n6365 = ~n6364 & ~n6363;
  assign U3266 = ~n6366 | ~n6365;
  assign n6369 = ~n6368 | ~n6367;
  assign n6432 = ~n6369 | ~n6461;
  assign n6372 = ~n6432 | ~n6370;
  assign n6393 = ~n6661 & ~n7707;
  assign n6378 = n6375 | n6376;
  assign n6434 = ~n6378 | ~n6377;
  assign n6380 = ~n6434 | ~n6433;
  assign n6406 = ~n6380 | ~n6379;
  assign n6408 = ~n6406 | ~n6428;
  assign n6383 = ~n6408 | ~n6381;
  assign n6384 = n6383 ^ ~n6382;
  assign n6391 = ~n6384 | ~n7678;
  assign n6386 = ~n7982 | ~n7709;
  assign n6385 = ~n7714 | ~n6398;
  assign n6389 = ~n6386 | ~n6385;
  assign n6388 = ~n6387 & ~n7668;
  assign n6390 = ~n6389 & ~n6388;
  assign n6392 = ~n6391 | ~n6390;
  assign n6666 = ~n6393 & ~n6392;
  assign n6395 = ~n6666 | ~n7608;
  assign n6394 = n7608 | REG2_REG_23__SCAN_IN;
  assign n6405 = ~n6395 | ~n6394;
  assign n6403 = n6661 | n7702;
  assign n6422 = ~n6396 | ~n6397;
  assign n6662 = n6422 ^ ~n6398;
  assign n6401 = n6662 | n7642;
  assign n6400 = n7632 | n6399;
  assign n6402 = n6401 & n6400;
  assign n6404 = n6403 & n6402;
  assign U3267 = ~n6405 | ~n6404;
  assign n6407 = n6406 | n6428;
  assign n6409 = ~n6408 | ~n6407;
  assign n6416 = ~n6409 | ~n7678;
  assign n6412 = ~n7979 | ~n7709;
  assign n6411 = ~n7714 | ~n6410;
  assign n6414 = ~n6412 | ~n6411;
  assign n6413 = ~n6466 & ~n7668;
  assign n6415 = ~n6414 & ~n6413;
  assign n6672 = ~n6416 | ~n6415;
  assign n6418 = ~n6672 & ~n7698;
  assign n6417 = ~n7608 & ~REG2_REG_22__SCAN_IN;
  assign n6427 = ~n6418 & ~n6417;
  assign n6420 = n6396 & n6448;
  assign n6421 = n6420 | n6419;
  assign n6670 = ~n6422 | ~n6421;
  assign n6425 = ~n6670 & ~n7642;
  assign n6424 = ~n7632 & ~n6423;
  assign n6426 = n6425 | n6424;
  assign n6431 = ~n6427 & ~n6426;
  assign n6669 = n6429 ^ ~n6428;
  assign n6430 = ~n6669 | ~n6528;
  assign U3268 = ~n6431 | ~n6430;
  assign n6677 = n6432 ^ ~n6433;
  assign n6445 = ~n6677 & ~n7707;
  assign n6435 = n6434 ^ ~n6433;
  assign n6443 = ~n6435 | ~n7678;
  assign n6441 = ~n6436 & ~n7668;
  assign n6439 = ~n7976 | ~n7709;
  assign n6438 = ~n7714 | ~n6437;
  assign n6440 = ~n6439 | ~n6438;
  assign n6442 = ~n6441 & ~n6440;
  assign n6444 = ~n6443 | ~n6442;
  assign n6682 = ~n6445 & ~n6444;
  assign n6447 = ~n6682 | ~n7608;
  assign n6446 = n7608 | REG2_REG_21__SCAN_IN;
  assign n6455 = ~n6447 | ~n6446;
  assign n6453 = ~n6677 & ~n7702;
  assign n6678 = n6396 ^ ~n6448;
  assign n6451 = n6678 | n7642;
  assign n6450 = ~n7699 | ~n6449;
  assign n6452 = ~n6451 | ~n6450;
  assign n6454 = ~n6453 & ~n6452;
  assign U3269 = ~n6455 | ~n6454;
  assign n6548 = n7376 | n6456;
  assign n6552 = ~n6548 | ~n6457;
  assign n6527 = ~n6552 | ~n6458;
  assign n6475 = ~n6527 | ~n6459;
  assign n6498 = ~n6475 | ~n6460;
  assign n6464 = ~n6461 | ~n6460;
  assign n6463 = ~n6462;
  assign n6473 = n6464 | n6463;
  assign n7648 = ~n7707;
  assign n6465 = ~n6473 | ~n7648;
  assign n6472 = ~n6498 & ~n6465;
  assign n6468 = ~n6466 & ~n7573;
  assign n6467 = ~n7671 & ~n6489;
  assign n6470 = ~n6468 & ~n6467;
  assign n6469 = ~n7967 | ~n7533;
  assign n6471 = ~n6470 | ~n6469;
  assign n6488 = ~n6472 & ~n6471;
  assign n6474 = ~n6473;
  assign n6476 = ~n6475 | ~n6474;
  assign n6482 = ~n6476 | ~n7648;
  assign n6479 = n6375 | n6477;
  assign n6483 = ~n6479 | ~n6478;
  assign n6480 = ~n6483 & ~n7706;
  assign n6481 = ~n6480 & ~n6499;
  assign n6486 = ~n6482 | ~n6481;
  assign n6484 = ~n6483 | ~n7678;
  assign n6485 = ~n6484 | ~n6499;
  assign n6487 = ~n6486 | ~n6485;
  assign n6686 = ~n6488 | ~n6487;
  assign n6490 = n6516 ^ ~n6489;
  assign n6685 = ~n6490 & ~n7858;
  assign n6491 = ~n6685 | ~n7516;
  assign n6492 = ~n6491 | ~n7608;
  assign n6494 = ~n6686 & ~n6492;
  assign n6493 = ~n7608 & ~REG2_REG_20__SCAN_IN;
  assign n6497 = ~n6494 & ~n6493;
  assign n6496 = ~n6495 & ~n7632;
  assign n6501 = ~n6497 & ~n6496;
  assign n6687 = n6499 ^ n6498;
  assign n7527 = ~n7702;
  assign n6500 = ~n6687 | ~n7527;
  assign U3270 = ~n6501 | ~n6500;
  assign n6505 = ~n6532 | ~n6503;
  assign n6506 = ~n6505 | ~n6504;
  assign n6507 = n6506 ^ ~n6526;
  assign n6513 = ~n6507 | ~n7678;
  assign n6511 = ~n7970 | ~n7709;
  assign n6509 = ~n7964 | ~n7533;
  assign n6508 = ~n7714 | ~n6517;
  assign n6510 = n6509 & n6508;
  assign n6512 = n6511 & n6510;
  assign n6695 = ~n6513 | ~n6512;
  assign n6515 = ~n6695 & ~n7698;
  assign n6514 = ~n7608 & ~REG2_REG_19__SCAN_IN;
  assign n6525 = ~n6515 & ~n6514;
  assign n6520 = ~n6516;
  assign n6519 = ~n6518 | ~n6517;
  assign n6693 = ~n6520 | ~n6519;
  assign n6523 = n6693 | n7642;
  assign n6522 = ~n7699 | ~n6521;
  assign n6524 = ~n6523 | ~n6522;
  assign n6530 = ~n6525 & ~n6524;
  assign n6692 = n6527 ^ ~n6526;
  assign n6529 = ~n6692 | ~n6528;
  assign U3271 = ~n6530 | ~n6529;
  assign n6533 = ~n6532 | ~n6531;
  assign n6534 = n6533 ^ ~n6549;
  assign n6541 = ~n6534 | ~n7678;
  assign n6536 = ~n7967 | ~n7709;
  assign n6535 = ~n7714 | ~n6543;
  assign n6539 = ~n6536 | ~n6535;
  assign n6538 = ~n6537 & ~n7668;
  assign n6540 = ~n6539 & ~n6538;
  assign n6701 = ~n6541 | ~n6540;
  assign n6544 = n6542 ^ ~n6543;
  assign n6700 = ~n6544 & ~n7858;
  assign n6545 = ~n6700 | ~n7516;
  assign n6546 = ~n6545 | ~n7608;
  assign n6554 = ~n6701 & ~n6546;
  assign n6550 = ~n6548 | ~n6547;
  assign n6551 = ~n6550 | ~n6549;
  assign n6702 = ~n6552 | ~n6551;
  assign n6553 = ~n6702 | ~n7513;
  assign n6557 = ~n6554 | ~n6553;
  assign n6555 = ~REG2_REG_18__SCAN_IN;
  assign n6556 = ~n7698 | ~n6555;
  assign n6560 = ~n6557 | ~n6556;
  assign n6559 = ~n7699 | ~n6558;
  assign U3272 = ~n6560 | ~n6559;
  assign n6563 = n7376 | n6561;
  assign n6564 = ~n6563 | ~n6562;
  assign n6707 = n6565 ^ n6564;
  assign n6578 = ~n6707 | ~n7513;
  assign n6566 = n6375 ^ ~n6565;
  assign n6573 = ~n6566 | ~n7678;
  assign n6571 = ~n6567 & ~n7668;
  assign n6569 = ~n7964 | ~n7709;
  assign n6568 = ~n7714 | ~n6583;
  assign n6570 = ~n6569 | ~n6568;
  assign n6572 = ~n6571 & ~n6570;
  assign n6710 = ~n6573 | ~n6572;
  assign n6575 = ~n7699 | ~n6574;
  assign n6576 = ~n7608 | ~n6575;
  assign n6577 = ~n6710 & ~n6576;
  assign n6581 = ~n6578 | ~n6577;
  assign n6579 = ~REG2_REG_17__SCAN_IN;
  assign n6580 = ~n7698 | ~n6579;
  assign n6586 = ~n6581 | ~n6580;
  assign n6584 = ~n6582 | ~n6583;
  assign n6708 = ~n6542 | ~n6584;
  assign n6585 = n6708 | n7642;
  assign U3273 = ~n6586 | ~n6585;
  assign n7329 = ~n6589 | ~n6588;
  assign n6592 = ~n7329 | ~n6590;
  assign n6593 = ~n6592 | ~n6591;
  assign n6715 = n6593 ^ ~n6595;
  assign n6606 = ~n6715 & ~n7707;
  assign n6596 = n6594 ^ ~n6595;
  assign n6604 = ~n6596 | ~n7678;
  assign n6602 = ~n6597 & ~n7668;
  assign n6600 = ~n7961 | ~n7709;
  assign n6599 = ~n7714 | ~n6598;
  assign n6601 = ~n6600 | ~n6599;
  assign n6603 = ~n6602 & ~n6601;
  assign n6605 = ~n6604 | ~n6603;
  assign n6720 = ~n6606 & ~n6605;
  assign n6609 = ~n6720 | ~n7608;
  assign n6607 = ~REG2_REG_16__SCAN_IN;
  assign n6608 = ~n7698 | ~n6607;
  assign n6619 = ~n6609 | ~n6608;
  assign n6617 = ~n6715 & ~n7702;
  assign n6612 = n6611 | n6610;
  assign n6716 = ~n6582 | ~n6612;
  assign n6615 = n6716 | n7642;
  assign n6614 = ~n7699 | ~n6613;
  assign n6616 = ~n6615 | ~n6614;
  assign n6618 = ~n6617 & ~n6616;
  assign U3274 = ~n6619 | ~n6618;
  assign n7883 = ~n7858;
  assign n6623 = ~n6746 | ~n7954;
  assign n6622 = ~n7952 | ~REG1_REG_31__SCAN_IN;
  assign U3549 = ~n6623 | ~n6622;
  assign n6626 = ~n6624 | ~n7883;
  assign n6749 = ~n6626 | ~n6625;
  assign n6628 = ~n6749 | ~n7954;
  assign n6627 = ~n7952 | ~REG1_REG_30__SCAN_IN;
  assign U3548 = ~n6628 | ~n6627;
  assign n6630 = ~n6629 & ~n7858;
  assign n6633 = ~n6632 | ~n7887;
  assign n6752 = ~n6634 | ~n6633;
  assign n6636 = ~n6752 | ~n7954;
  assign n6635 = ~n7952 | ~REG1_REG_27__SCAN_IN;
  assign U3545 = ~n6636 | ~n6635;
  assign n6640 = ~n6637 & ~n7901;
  assign n6639 = ~n6638 & ~n7858;
  assign n6641 = ~n6640 & ~n6639;
  assign n6755 = ~n6642 | ~n6641;
  assign n6644 = ~n6755 | ~n7954;
  assign n6643 = ~n7952 | ~REG1_REG_26__SCAN_IN;
  assign U3544 = ~n6644 | ~n6643;
  assign n6650 = ~n6645 | ~n7887;
  assign n6647 = ~n6646 & ~n7858;
  assign n6649 = ~n6648 & ~n6647;
  assign n6758 = ~n6650 | ~n6649;
  assign n6652 = ~n6758 | ~n7954;
  assign n6651 = ~n7952 | ~REG1_REG_25__SCAN_IN;
  assign U3543 = ~n6652 | ~n6651;
  assign n6656 = ~n6653 & ~n7901;
  assign n6655 = ~n6654 & ~n7858;
  assign n6657 = ~n6656 & ~n6655;
  assign n6761 = ~n6658 | ~n6657;
  assign n6660 = ~n6761 | ~n7954;
  assign n6659 = ~n7952 | ~REG1_REG_24__SCAN_IN;
  assign U3542 = ~n6660 | ~n6659;
  assign n6663 = n6662 | n7858;
  assign n6665 = n6664 & n6663;
  assign n6764 = ~n6666 | ~n6665;
  assign n6668 = ~n6764 | ~n7954;
  assign n6667 = ~n7952 | ~REG1_REG_23__SCAN_IN;
  assign U3541 = ~n6668 | ~n6667;
  assign n6674 = ~n6669 | ~n7887;
  assign n6671 = ~n6670 & ~n7858;
  assign n6673 = ~n6672 & ~n6671;
  assign n6767 = ~n6674 | ~n6673;
  assign n6676 = ~n6767 | ~n7954;
  assign n6675 = ~n7952 | ~REG1_REG_22__SCAN_IN;
  assign U3540 = ~n6676 | ~n6675;
  assign n6680 = ~n6677 & ~n7901;
  assign n6679 = ~n6678 & ~n7858;
  assign n6681 = ~n6680 & ~n6679;
  assign n6770 = ~n6682 | ~n6681;
  assign n6684 = ~n6770 | ~n7954;
  assign n6683 = ~n7952 | ~REG1_REG_21__SCAN_IN;
  assign U3539 = ~n6684 | ~n6683;
  assign n6689 = ~n6686 & ~n6685;
  assign n7852 = ~n7901;
  assign n6688 = ~n6687 | ~n7852;
  assign n6773 = ~n6689 | ~n6688;
  assign n6691 = ~n6773 | ~n7954;
  assign n6690 = ~n7952 | ~REG1_REG_20__SCAN_IN;
  assign U3538 = ~n6691 | ~n6690;
  assign n6697 = ~n6692 | ~n7887;
  assign n6694 = ~n6693 & ~n7858;
  assign n6696 = ~n6695 & ~n6694;
  assign n6776 = ~n6697 | ~n6696;
  assign n6699 = ~n6776 | ~n7954;
  assign n6698 = ~n7952 | ~REG1_REG_19__SCAN_IN;
  assign U3537 = ~n6699 | ~n6698;
  assign n6704 = ~n6701 & ~n6700;
  assign n6703 = ~n6702 | ~n7887;
  assign n6779 = ~n6704 | ~n6703;
  assign n6706 = ~n6779 | ~n7954;
  assign n6705 = ~n7952 | ~REG1_REG_18__SCAN_IN;
  assign U3536 = ~n6706 | ~n6705;
  assign n6712 = ~n6707 | ~n7887;
  assign n6709 = ~n6708 & ~n7858;
  assign n6711 = ~n6710 & ~n6709;
  assign n6782 = ~n6712 | ~n6711;
  assign n6714 = ~n6782 | ~n7954;
  assign n6713 = ~n7952 | ~REG1_REG_17__SCAN_IN;
  assign U3535 = ~n6714 | ~n6713;
  assign n6718 = ~n6715 & ~n7901;
  assign n6717 = ~n6716 & ~n7858;
  assign n6719 = ~n6718 & ~n6717;
  assign n6785 = ~n6720 | ~n6719;
  assign n6722 = ~n6785 | ~n7954;
  assign n6721 = ~n7952 | ~REG1_REG_16__SCAN_IN;
  assign U3534 = ~n6722 | ~n6721;
  assign n6724 = n6723 ^ ~n6740;
  assign n6731 = ~n6724 & ~n7706;
  assign n6727 = ~n6725 & ~n7668;
  assign n6726 = ~n7671 & ~n6732;
  assign n6729 = ~n6727 & ~n6726;
  assign n6728 = ~n7958 | ~n7709;
  assign n6730 = ~n6729 | ~n6728;
  assign n7295 = ~n6731 & ~n6730;
  assign n7289 = n6733 ^ ~n6732;
  assign n6734 = ~n7289 | ~n7883;
  assign n6743 = n7295 & n6734;
  assign n6737 = ~n7329 | ~n6735;
  assign n7300 = ~n6737 | ~n6736;
  assign n6739 = n7300 | n7309;
  assign n6741 = ~n6739 | ~n6738;
  assign n7288 = n6741 ^ ~n6740;
  assign n6742 = ~n7288 | ~n7887;
  assign n6788 = ~n6743 | ~n6742;
  assign n6745 = ~n6788 | ~n7954;
  assign n6744 = ~n7952 | ~REG1_REG_15__SCAN_IN;
  assign U3533 = ~n6745 | ~n6744;
  assign n6748 = ~n6746 | ~n7907;
  assign n6747 = ~n7900 | ~REG0_REG_31__SCAN_IN;
  assign U3517 = ~n6748 | ~n6747;
  assign n6751 = ~n6749 | ~n7907;
  assign n6750 = ~n7900 | ~REG0_REG_30__SCAN_IN;
  assign U3516 = ~n6751 | ~n6750;
  assign n6754 = ~n6752 | ~n7907;
  assign n6753 = ~n7900 | ~REG0_REG_27__SCAN_IN;
  assign U3513 = ~n6754 | ~n6753;
  assign n6757 = ~n6755 | ~n7907;
  assign n6756 = ~n7900 | ~REG0_REG_26__SCAN_IN;
  assign U3512 = ~n6757 | ~n6756;
  assign n6760 = ~n6758 | ~n7907;
  assign n6759 = ~n7900 | ~REG0_REG_25__SCAN_IN;
  assign U3511 = ~n6760 | ~n6759;
  assign n6763 = ~n6761 | ~n7907;
  assign n6762 = ~n7900 | ~REG0_REG_24__SCAN_IN;
  assign U3510 = ~n6763 | ~n6762;
  assign n6766 = ~n6764 | ~n7907;
  assign n6765 = ~n7900 | ~REG0_REG_23__SCAN_IN;
  assign U3509 = ~n6766 | ~n6765;
  assign n6769 = ~n6767 | ~n7907;
  assign n6768 = ~n7900 | ~REG0_REG_22__SCAN_IN;
  assign U3508 = ~n6769 | ~n6768;
  assign n6772 = ~n6770 | ~n7907;
  assign n6771 = ~n7900 | ~REG0_REG_21__SCAN_IN;
  assign U3507 = ~n6772 | ~n6771;
  assign n6775 = ~n6773 | ~n7907;
  assign n6774 = ~n7900 | ~REG0_REG_20__SCAN_IN;
  assign U3506 = ~n6775 | ~n6774;
  assign n6778 = ~n6776 | ~n7907;
  assign n6777 = ~n7900 | ~REG0_REG_19__SCAN_IN;
  assign U3505 = ~n6778 | ~n6777;
  assign n6781 = ~n6779 | ~n7907;
  assign n6780 = ~n7900 | ~REG0_REG_18__SCAN_IN;
  assign U3503 = ~n6781 | ~n6780;
  assign n6784 = ~n6782 | ~n7907;
  assign n6783 = ~n7900 | ~REG0_REG_17__SCAN_IN;
  assign U3501 = ~n6784 | ~n6783;
  assign n6787 = ~n6785 | ~n7907;
  assign n6786 = ~n7900 | ~REG0_REG_16__SCAN_IN;
  assign U3499 = ~n6787 | ~n6786;
  assign n6790 = ~n6788 | ~n7907;
  assign n6789 = ~n7900 | ~REG0_REG_15__SCAN_IN;
  assign U3497 = ~n6790 | ~n6789;
  assign n6791 = ~n6991 | ~n7451;
  assign n7118 = ~REG3_REG_7__SCAN_IN | ~U3149;
  assign n6795 = ~n6791 | ~n7118;
  assign n6793 = ~n6990 | ~n7504;
  assign n6792 = ~n6988 | ~n7503;
  assign n6794 = ~n6793 | ~n6792;
  assign n6802 = ~n6795 & ~n6794;
  assign n6797 = n5855 ^ ~n6796;
  assign n6800 = ~n6797 & ~n7007;
  assign n6799 = ~n7009 & ~n7521;
  assign n6801 = ~n6800 & ~n6799;
  assign U3210 = ~n6802 | ~n6801;
  assign n6803 = ~n6988 | ~n7314;
  assign n7219 = ~REG3_REG_14__SCAN_IN | ~U3149;
  assign n6807 = ~n6803 | ~n7219;
  assign n6805 = ~n6990 | ~n7315;
  assign n6804 = ~n6991 | ~n7316;
  assign n6806 = ~n6805 | ~n6804;
  assign n6814 = ~n6807 & ~n6806;
  assign n6810 = n6809 ^ n6808;
  assign n6812 = ~n6810 & ~n7007;
  assign n6811 = ~n7009 & ~n7305;
  assign n6813 = ~n6812 & ~n6811;
  assign U3212 = ~n6814 | ~n6813;
  assign n6815 = ~n6988 | ~n6840;
  assign n7163 = ~REG3_REG_10__SCAN_IN | ~U3149;
  assign n6819 = ~n6815 | ~n7163;
  assign n6817 = ~n6990 | ~n4886;
  assign n6816 = ~n6991 | ~n4906;
  assign n6818 = ~n6817 | ~n6816;
  assign n6825 = ~n6819 & ~n6818;
  assign n6821 = n6962 ^ ~n6963;
  assign n6823 = ~n6821 & ~n7007;
  assign n6822 = ~n7009 & ~n7435;
  assign n6824 = ~n6823 & ~n6822;
  assign U3214 = ~n6825 | ~n6824;
  assign n6827 = ~n6988 | ~n7680;
  assign n6831 = ~n6827 | ~n6826;
  assign n6829 = ~n6990 | ~n7618;
  assign n6828 = ~n6991 | ~n7617;
  assign n6830 = ~n6829 | ~n6828;
  assign n6838 = ~n6831 & ~n6830;
  assign n6834 = n6832 ^ n6833;
  assign n6836 = ~n6834 & ~n7007;
  assign n6835 = ~REG3_REG_3__SCAN_IN & ~n7009;
  assign n6837 = ~n6836 & ~n6835;
  assign U3215 = ~n6838 | ~n6837;
  assign n6839 = ~n6988 | ~n7486;
  assign n7136 = ~REG3_REG_8__SCAN_IN | ~U3149;
  assign n6844 = ~n6839 | ~n7136;
  assign n6842 = ~n6990 | ~n7471;
  assign n6841 = ~n6991 | ~n6840;
  assign n6843 = ~n6842 | ~n6841;
  assign n6853 = ~n6844 & ~n6843;
  assign n6848 = ~n6846 | ~n6845;
  assign n6849 = n6848 ^ n6847;
  assign n6851 = ~n6849 & ~n7007;
  assign n6850 = ~n7009 & ~n7465;
  assign n6852 = ~n6851 & ~n6850;
  assign U3218 = ~n6853 | ~n6852;
  assign n7669 = ~n6854;
  assign n6856 = ~n6955 & ~n7669;
  assign n6855 = ~n6951 & ~n5581;
  assign n6866 = ~n6856 & ~n6855;
  assign n6857 = ~REG3_REG_1__SCAN_IN;
  assign n6864 = ~n6983 & ~n6857;
  assign n6860 = n6858 ^ n6859;
  assign n6862 = ~n6860 | ~n6970;
  assign n6861 = ~n6990 | ~n4729;
  assign n6863 = ~n6862 | ~n6861;
  assign n6865 = ~n6864 & ~n6863;
  assign U3219 = ~n6866 | ~n6865;
  assign n6867 = ~n6991 | ~n7314;
  assign n7191 = ~REG3_REG_12__SCAN_IN | ~U3149;
  assign n6871 = ~n6867 | ~n7191;
  assign n6869 = ~n6990 | ~n7368;
  assign n6868 = ~n6988 | ~n4906;
  assign n6870 = ~n6869 | ~n6868;
  assign n6888 = ~n6871 & ~n6870;
  assign n6877 = ~n6963 | ~n6872;
  assign n6874 = ~n6877 | ~n6873;
  assign n6883 = ~n6874 & ~n6879;
  assign n6876 = ~n6875;
  assign n6881 = n6877 & n6876;
  assign n6880 = ~n6879 & ~n6878;
  assign n6882 = ~n6881 & ~n6880;
  assign n6884 = ~n6883 & ~n6882;
  assign n6886 = ~n6884 & ~n7007;
  assign n6885 = ~n7009 & ~n7387;
  assign n6887 = ~n6886 & ~n6885;
  assign U3221 = ~n6888 | ~n6887;
  assign n6889 = ~n6991 | ~n7503;
  assign n7092 = ~REG3_REG_5__SCAN_IN | ~U3149;
  assign n6893 = ~n6889 | ~n7092;
  assign n6891 = ~n6990 | ~n7571;
  assign n6890 = ~n6988 | ~n7617;
  assign n6892 = ~n6891 | ~n6890;
  assign n6903 = ~n6893 & ~n6892;
  assign n6896 = n6894 | n6909;
  assign n6897 = ~n6896 | ~n6895;
  assign n6899 = n6898 ^ ~n6897;
  assign n6901 = ~n6899 & ~n7007;
  assign n6900 = ~n7009 & ~n7553;
  assign n6902 = ~n6901 & ~n6900;
  assign U3224 = ~n6903 | ~n6902;
  assign n6904 = ~n6991 | ~n7583;
  assign n7075 = ~REG3_REG_4__SCAN_IN | ~U3149;
  assign n6908 = ~n6904 | ~n7075;
  assign n6906 = ~n6990 | ~n7584;
  assign n6905 = ~n6988 | ~n7651;
  assign n6907 = ~n6906 | ~n6905;
  assign n6914 = ~n6908 & ~n6907;
  assign n6910 = n6894 ^ ~n6909;
  assign n6912 = ~n6910 & ~n7007;
  assign n6911 = ~n7009 & ~n7602;
  assign n6913 = ~n6912 & ~n6911;
  assign U3227 = ~n6914 | ~n6913;
  assign n6916 = ~n6955 & ~n7502;
  assign n7147 = ~STATE_REG_SCAN_IN & ~n6915;
  assign n6929 = ~n6916 & ~n7147;
  assign n6918 = ~n6938 | ~n6917;
  assign n6920 = ~n6919 | ~n6918;
  assign n6925 = ~n6920 | ~n6970;
  assign n6923 = ~n6974 & ~n6921;
  assign n6922 = ~n6951 & ~n7450;
  assign n6924 = ~n6923 & ~n6922;
  assign n6927 = ~n6925 | ~n6924;
  assign n6926 = ~n7009 & ~n7440;
  assign n6928 = ~n6927 & ~n6926;
  assign U3228 = ~n6929 | ~n6928;
  assign n6930 = ~n6991 | ~n7351;
  assign n7203 = ~REG3_REG_13__SCAN_IN | ~U3149;
  assign n6934 = ~n6930 | ~n7203;
  assign n6932 = ~n6990 | ~n7352;
  assign n6931 = ~n6988 | ~n7394;
  assign n6933 = ~n6932 | ~n6931;
  assign n6950 = ~n6934 & ~n6933;
  assign n6936 = ~n6935;
  assign n6945 = ~n6936 & ~n6941;
  assign n6940 = n6938 | n6937;
  assign n6943 = ~n6940 | ~n6939;
  assign n6942 = ~n4386 & ~n6941;
  assign n6944 = ~n6943 & ~n6942;
  assign n6946 = ~n6945 & ~n6944;
  assign n6948 = ~n6946 & ~n7007;
  assign n6947 = ~n7009 & ~n7336;
  assign n6949 = ~n6948 & ~n6947;
  assign U3231 = ~n6950 | ~n6949;
  assign n6953 = ~n6951 & ~n7350;
  assign n7175 = ~STATE_REG_SCAN_IN & ~n6952;
  assign n6959 = ~n6953 & ~n7175;
  assign n6957 = ~n6974 & ~n6954;
  assign n6956 = ~n6955 & ~n7450;
  assign n6958 = ~n6957 & ~n6956;
  assign n6961 = ~n6959 | ~n6958;
  assign n6960 = ~n7009 & ~n7407;
  assign n6973 = ~n6961 & ~n6960;
  assign n6965 = ~n6963 | ~n6962;
  assign n6969 = ~n6965 | ~n6964;
  assign n6968 = ~n6967 | ~n6966;
  assign n6971 = n6969 ^ ~n6968;
  assign n6972 = ~n6971 | ~n6970;
  assign U3233 = ~n6973 | ~n6972;
  assign n6978 = ~n6974 & ~n5567;
  assign n6976 = ~n6988 | ~n5496;
  assign n6975 = ~n6991 | ~n7651;
  assign n6977 = ~n6976 | ~n6975;
  assign n6987 = ~n6978 & ~n6977;
  assign n6981 = n6980 ^ n6979;
  assign n6985 = ~n6981 & ~n7007;
  assign n6982 = ~REG3_REG_2__SCAN_IN;
  assign n6984 = ~n6983 & ~n6982;
  assign n6986 = ~n6985 & ~n6984;
  assign U3234 = ~n6987 | ~n6986;
  assign n6989 = ~n6988 | ~n7583;
  assign n7106 = ~REG3_REG_6__SCAN_IN | ~U3149;
  assign n6995 = ~n6989 | ~n7106;
  assign n6993 = ~n6990 | ~n7534;
  assign n6992 = ~n6991 | ~n7486;
  assign n6994 = ~n6993 | ~n6992;
  assign n7013 = ~n6995 & ~n6994;
  assign n6996 = ~n7002;
  assign n7006 = ~n6997 & ~n6996;
  assign n6999 = ~n6998;
  assign n7004 = ~n6999 & ~n7000;
  assign n7003 = n7002 & n7001;
  assign n7005 = ~n7004 & ~n7003;
  assign n7008 = ~n7006 & ~n7005;
  assign n7011 = ~n7008 & ~n7007;
  assign n7010 = ~n7009 & ~n7546;
  assign n7012 = ~n7011 & ~n7010;
  assign U3236 = ~n7013 | ~n7012;
  assign n7014 = ~n7058 & ~REG2_REG_0__SCAN_IN;
  assign n7062 = n7069 | n7014;
  assign n7015 = ~n7067 & ~REG1_REG_0__SCAN_IN;
  assign n7016 = n7062 | n7015;
  assign n7017 = IR_REG_0__SCAN_IN ^ n7016;
  assign n7021 = ~n7018 & ~n7017;
  assign n7020 = ~STATE_REG_SCAN_IN & ~n7019;
  assign n7023 = ~n7021 & ~n7020;
  assign n7022 = ~n7270 | ~ADDR_REG_0__SCAN_IN;
  assign U3240 = ~n7023 | ~n7022;
  assign n7025 = ~ADDR_REG_1__SCAN_IN | ~n7270;
  assign n7024 = ~REG3_REG_1__SCAN_IN | ~U3149;
  assign n7033 = ~n7025 | ~n7024;
  assign n7028 = n7027 ^ ~n7026;
  assign n7031 = ~n7275 | ~n7028;
  assign n7030 = ~n7277 | ~n7029;
  assign n7032 = ~n7031 | ~n7030;
  assign n7038 = ~n7033 & ~n7032;
  assign n7036 = n7035 ^ n7034;
  assign n7037 = ~n7284 | ~n7036;
  assign U3241 = ~n7038 | ~n7037;
  assign n7040 = ~ADDR_REG_2__SCAN_IN | ~n7270;
  assign n7039 = ~REG3_REG_2__SCAN_IN | ~U3149;
  assign n7057 = ~n7040 | ~n7039;
  assign n7045 = ~n7275 | ~n7041;
  assign n7044 = ~n7043 & ~n7042;
  assign n7052 = ~n7045 & ~n7044;
  assign n7050 = ~n7047 & ~n7046;
  assign n7049 = ~n7284 | ~n7048;
  assign n7051 = ~n7050 & ~n7049;
  assign n7055 = ~n7052 & ~n7051;
  assign n7054 = ~n7277 | ~n7053;
  assign n7056 = ~n7055 | ~n7054;
  assign n7073 = ~n7057 & ~n7056;
  assign n7060 = ~n7059 | ~n7058;
  assign n7065 = ~n7061 & ~n7060;
  assign n7063 = ~n7062;
  assign n7064 = ~n7063 & ~IR_REG_0__SCAN_IN;
  assign n7072 = ~n7065 & ~n7064;
  assign n7068 = ~n7067 | ~n7066;
  assign n7070 = ~n7069 & ~n7068;
  assign n7071 = ~n8000 & ~n7070;
  assign n7089 = ~n7072 | ~n7071;
  assign U3242 = ~n7073 | ~n7089;
  assign n7074 = ~n7270 | ~ADDR_REG_4__SCAN_IN;
  assign n7088 = ~n7075 | ~n7074;
  assign n7078 = n7076 ^ ~REG1_REG_4__SCAN_IN;
  assign n7082 = ~n7078 & ~n7077;
  assign n7081 = ~n7080 & ~n7079;
  assign n7086 = ~n7082 & ~n7081;
  assign n7084 = n7083 ^ ~REG2_REG_4__SCAN_IN;
  assign n7085 = ~n7275 | ~n7084;
  assign n7087 = ~n7086 | ~n7085;
  assign n7090 = ~n7088 & ~n7087;
  assign U3244 = ~n7090 | ~n7089;
  assign n7091 = ~n7270 | ~ADDR_REG_5__SCAN_IN;
  assign n7102 = ~n7092 | ~n7091;
  assign n7095 = n7094 ^ n7093;
  assign n7100 = ~n7095 | ~n7275;
  assign n7098 = n7097 ^ n7096;
  assign n7099 = ~n7098 | ~n7284;
  assign n7101 = ~n7100 | ~n7099;
  assign n7104 = ~n7102 & ~n7101;
  assign n7103 = ~n7277 | ~n7768;
  assign U3245 = ~n7104 | ~n7103;
  assign n7105 = ~n7270 | ~ADDR_REG_6__SCAN_IN;
  assign n7112 = ~n7106 | ~n7105;
  assign n7108 = n7107 ^ REG1_REG_6__SCAN_IN;
  assign n7110 = ~n7108 | ~n7284;
  assign n7109 = ~n7277 | ~n7765;
  assign n7111 = ~n7110 | ~n7109;
  assign n7116 = ~n7112 & ~n7111;
  assign n7114 = n7113 ^ REG2_REG_6__SCAN_IN;
  assign n7115 = ~n7275 | ~n7114;
  assign U3246 = ~n7116 | ~n7115;
  assign n7117 = ~n7270 | ~ADDR_REG_7__SCAN_IN;
  assign n7132 = ~n7118 | ~n7117;
  assign n7121 = ~n7120 | ~n7119;
  assign n7123 = n7122 ^ n7121;
  assign n7130 = ~n7123 | ~n7275;
  assign n7127 = ~n7125 & ~n7124;
  assign n7128 = n7127 ^ n7126;
  assign n7129 = ~n7128 | ~n7284;
  assign n7131 = ~n7130 | ~n7129;
  assign n7134 = ~n7132 & ~n7131;
  assign n7133 = ~n7277 | ~n7762;
  assign U3247 = ~n7134 | ~n7133;
  assign n7135 = ~n7270 | ~ADDR_REG_8__SCAN_IN;
  assign n7142 = ~n7136 | ~n7135;
  assign n7138 = n7137 ^ REG2_REG_8__SCAN_IN;
  assign n7140 = ~n7138 | ~n7275;
  assign n7139 = ~n7277 | ~n7759;
  assign n7141 = ~n7140 | ~n7139;
  assign n7146 = ~n7142 & ~n7141;
  assign n7144 = n7143 ^ REG1_REG_8__SCAN_IN;
  assign n7145 = ~n7144 | ~n7284;
  assign U3248 = ~n7146 | ~n7145;
  assign n7149 = ~n7147;
  assign n7148 = ~n7270 | ~ADDR_REG_9__SCAN_IN;
  assign n7159 = ~n7149 | ~n7148;
  assign n7152 = n7151 ^ n7150;
  assign n7157 = ~n7152 | ~n7275;
  assign n7155 = n7154 ^ n7153;
  assign n7156 = ~n7155 | ~n7284;
  assign n7158 = ~n7157 | ~n7156;
  assign n7161 = ~n7159 & ~n7158;
  assign n7160 = ~n7277 | ~n7756;
  assign U3249 = ~n7161 | ~n7160;
  assign n7162 = ~n7270 | ~ADDR_REG_10__SCAN_IN;
  assign n7171 = ~n7163 | ~n7162;
  assign n7165 = n7164 ^ REG2_REG_10__SCAN_IN;
  assign n7169 = ~n7165 | ~n7275;
  assign n7167 = REG1_REG_10__SCAN_IN ^ n7166;
  assign n7168 = ~n7167 | ~n7284;
  assign n7170 = ~n7169 | ~n7168;
  assign n7173 = ~n7171 & ~n7170;
  assign n7172 = ~n7277 | ~n7753;
  assign U3250 = ~n7173 | ~n7172;
  assign n7174 = n7270 & ADDR_REG_11__SCAN_IN;
  assign n7189 = ~n7175 & ~n7174;
  assign n7178 = n7177 ^ n7176;
  assign n7180 = ~n7178 | ~n7275;
  assign n7179 = ~n7277 | ~n7750;
  assign n7187 = ~n7180 | ~n7179;
  assign n7185 = ~n7182 & ~n7181;
  assign n7184 = ~n7183 | ~n7284;
  assign n7186 = ~n7185 & ~n7184;
  assign n7188 = ~n7187 & ~n7186;
  assign U3251 = ~n7189 | ~n7188;
  assign n7190 = ~n7270 | ~ADDR_REG_12__SCAN_IN;
  assign n7199 = ~n7191 | ~n7190;
  assign n7193 = REG2_REG_12__SCAN_IN ^ n7192;
  assign n7197 = ~n7193 | ~n7275;
  assign n7195 = REG1_REG_12__SCAN_IN ^ n7194;
  assign n7196 = ~n7195 | ~n7284;
  assign n7198 = ~n7197 | ~n7196;
  assign n7201 = ~n7199 & ~n7198;
  assign n7200 = ~n7277 | ~n7747;
  assign U3252 = ~n7201 | ~n7200;
  assign n7202 = ~n7270 | ~ADDR_REG_13__SCAN_IN;
  assign n7215 = ~n7203 | ~n7202;
  assign n7206 = ~n7205 | ~n7204;
  assign n7208 = n7207 ^ n7206;
  assign n7213 = ~n7208 | ~n7275;
  assign n7211 = n7210 ^ n7209;
  assign n7212 = ~n7211 | ~n7284;
  assign n7214 = ~n7213 | ~n7212;
  assign n7217 = ~n7215 & ~n7214;
  assign n7216 = ~n7277 | ~n7744;
  assign U3253 = ~n7217 | ~n7216;
  assign n7218 = ~n7270 | ~ADDR_REG_14__SCAN_IN;
  assign n7227 = ~n7219 | ~n7218;
  assign n7221 = REG2_REG_14__SCAN_IN ^ n7220;
  assign n7225 = ~n7221 | ~n7275;
  assign n7223 = REG1_REG_14__SCAN_IN ^ n7222;
  assign n7224 = ~n7223 | ~n7284;
  assign n7226 = ~n7225 | ~n7224;
  assign n7229 = ~n7227 & ~n7226;
  assign n7228 = ~n7277 | ~n7741;
  assign U3254 = ~n7229 | ~n7228;
  assign n7230 = ~n7270 | ~ADDR_REG_15__SCAN_IN;
  assign n7238 = ~n7231 | ~n7230;
  assign n7234 = n7233 ^ n7232;
  assign n7236 = ~n7234 | ~n7275;
  assign n7235 = ~n7277 | ~n7738;
  assign n7237 = ~n7236 | ~n7235;
  assign n7243 = ~n7238 & ~n7237;
  assign n7241 = n7240 ^ n7239;
  assign n7242 = ~n7241 | ~n7284;
  assign U3255 = ~n7243 | ~n7242;
  assign n7244 = ~n7270 | ~ADDR_REG_16__SCAN_IN;
  assign n7251 = ~n7245 | ~n7244;
  assign n7247 = n7246 ^ ~REG2_REG_16__SCAN_IN;
  assign n7249 = ~n7247 | ~n7275;
  assign n7248 = ~n7277 | ~n7735;
  assign n7250 = ~n7249 | ~n7248;
  assign n7255 = ~n7251 & ~n7250;
  assign n7253 = REG1_REG_16__SCAN_IN ^ ~n7252;
  assign n7254 = ~n7253 | ~n7284;
  assign U3256 = ~n7255 | ~n7254;
  assign n7256 = ~n7270 | ~ADDR_REG_17__SCAN_IN;
  assign n7264 = ~n7257 | ~n7256;
  assign n7262 = ~n7277 | ~n7732;
  assign n7260 = n7258 ^ ~n7259;
  assign n7261 = ~n7275 | ~n7260;
  assign n7263 = ~n7262 | ~n7261;
  assign n7269 = ~n7264 & ~n7263;
  assign n7267 = n7266 ^ ~n7265;
  assign n7268 = ~n7267 | ~n7284;
  assign U3257 = ~n7269 | ~n7268;
  assign n7271 = ~n7270 | ~ADDR_REG_18__SCAN_IN;
  assign n7281 = ~n7272 | ~n7271;
  assign n7276 = n7274 ^ n7273;
  assign n7279 = ~n7276 | ~n7275;
  assign n7278 = ~n7277 | ~n7729;
  assign n7280 = ~n7279 | ~n7278;
  assign n7287 = ~n7281 & ~n7280;
  assign n7285 = n7283 ^ n7282;
  assign n7286 = ~n7285 | ~n7284;
  assign U3258 = ~n7287 | ~n7286;
  assign n7291 = ~n7288 | ~n7513;
  assign n7290 = ~n7289 | ~n7418;
  assign n7294 = ~n7291 | ~n7290;
  assign n7293 = ~n7292 & ~n7632;
  assign n7296 = ~n7294 & ~n7293;
  assign n7297 = ~n7296 | ~n7295;
  assign n7299 = ~n7608 | ~n7297;
  assign n7298 = ~n7698 | ~REG2_REG_15__SCAN_IN;
  assign U3275 = ~n7299 | ~n7298;
  assign n7902 = n7309 ^ n7300;
  assign n7301 = ~n7902;
  assign n7304 = ~n7301 | ~n7613;
  assign n7302 = n7332 ^ ~n7315;
  assign n7904 = ~n7302 & ~n7858;
  assign n7303 = ~n7904 | ~n7516;
  assign n7307 = ~n7304 | ~n7303;
  assign n7306 = ~n7305 & ~n7632;
  assign n7325 = ~n7307 & ~n7306;
  assign n7312 = ~n7308;
  assign n7311 = ~n7310 & ~n7309;
  assign n7313 = ~n7312 & ~n7311;
  assign n7324 = ~n7313 & ~n7706;
  assign n7322 = ~n7314 | ~n7533;
  assign n7318 = ~n7714 | ~n7315;
  assign n7317 = ~n7709 | ~n7316;
  assign n7320 = ~n7318 | ~n7317;
  assign n7319 = ~n7707 & ~n7902;
  assign n7321 = ~n7320 & ~n7319;
  assign n7323 = ~n7322 | ~n7321;
  assign n7906 = ~n7324 & ~n7323;
  assign n7326 = ~n7325 | ~n7906;
  assign n7328 = ~n7608 | ~n7326;
  assign n7327 = ~n7698 | ~REG2_REG_14__SCAN_IN;
  assign U3276 = ~n7328 | ~n7327;
  assign n7893 = n7329 ^ ~n7347;
  assign n7349 = ~n7893;
  assign n7335 = ~n7349 | ~n7613;
  assign n7331 = ~n7381 & ~n7330;
  assign n7333 = ~n7331 & ~n7858;
  assign n7895 = n7333 & n7332;
  assign n7334 = ~n7895 | ~n7516;
  assign n7338 = ~n7335 | ~n7334;
  assign n7337 = ~n7336 & ~n7632;
  assign n7361 = ~n7338 & ~n7337;
  assign n7342 = ~n7339 | ~n7340;
  assign n7345 = ~n7365 | ~n7343;
  assign n7346 = ~n7345 | ~n7344;
  assign n7348 = n7347 ^ n7346;
  assign n7360 = ~n7706 & ~n7348;
  assign n7358 = ~n7349 | ~n7648;
  assign n7356 = ~n7350 & ~n7668;
  assign n7354 = ~n7351 | ~n7709;
  assign n7353 = ~n7714 | ~n7352;
  assign n7355 = ~n7354 | ~n7353;
  assign n7357 = ~n7356 & ~n7355;
  assign n7359 = ~n7358 | ~n7357;
  assign n7897 = ~n7360 & ~n7359;
  assign n7362 = ~n7361 | ~n7897;
  assign n7364 = ~n7608 | ~n7362;
  assign n7363 = ~n7698 | ~REG2_REG_13__SCAN_IN;
  assign U3277 = ~n7364 | ~n7363;
  assign n7366 = n7365 ^ ~n7375;
  assign n7374 = ~n7366 | ~n7678;
  assign n7372 = ~n7367 & ~n7573;
  assign n7370 = ~n4906 | ~n7533;
  assign n7369 = ~n7368 | ~n7714;
  assign n7371 = ~n7370 | ~n7369;
  assign n7373 = ~n7372 & ~n7371;
  assign n7886 = ~n7374 | ~n7373;
  assign n7888 = n7376 ^ ~n7375;
  assign n7384 = ~n7888 | ~n7513;
  assign n7378 = ~n7377;
  assign n7380 = ~n7378 & ~n7405;
  assign n7382 = ~n7380 & ~n7379;
  assign n7884 = ~n7382 & ~n7381;
  assign n7383 = ~n7884 | ~n7418;
  assign n7385 = ~n7384 | ~n7383;
  assign n7386 = ~n7886 & ~n7385;
  assign n7389 = ~n7698 & ~n7386;
  assign n7388 = ~n7387 & ~n7632;
  assign n7391 = ~n7389 & ~n7388;
  assign n7390 = ~REG2_REG_12__SCAN_IN | ~n7698;
  assign U3278 = ~n7391 | ~n7390;
  assign n7392 = n7339 ^ n7398;
  assign n7404 = ~n7392 & ~n7706;
  assign n7402 = ~n7393 | ~n7533;
  assign n7396 = ~n7714 | ~n7405;
  assign n7395 = ~n7709 | ~n7394;
  assign n7400 = ~n7396 | ~n7395;
  assign n7876 = n7398 ^ n7397;
  assign n7399 = ~n7707 & ~n7876;
  assign n7401 = ~n7400 & ~n7399;
  assign n7403 = ~n7402 | ~n7401;
  assign n7880 = ~n7404 & ~n7403;
  assign n7875 = n7377 ^ ~n7405;
  assign n7406 = ~n7875 | ~n7418;
  assign n7409 = ~n7880 | ~n7406;
  assign n7408 = ~n7407 & ~n7632;
  assign n7410 = ~n7409 & ~n7408;
  assign n7412 = ~n7698 & ~n7410;
  assign n7411 = ~n7876 & ~n7702;
  assign n7414 = ~n7412 & ~n7411;
  assign n7413 = ~REG2_REG_11__SCAN_IN | ~n7698;
  assign U3279 = ~n7414 | ~n7413;
  assign n7868 = n7415 ^ ~n7426;
  assign n7433 = ~n7868 & ~n7691;
  assign n7417 = n7416 & n4886;
  assign n7867 = ~n7377 & ~n7417;
  assign n7431 = ~n7867 | ~n7418;
  assign n7422 = ~n7470 & ~n7668;
  assign n7420 = ~n7709 | ~n4906;
  assign n7419 = ~n7714 | ~n4886;
  assign n7421 = ~n7420 | ~n7419;
  assign n7425 = ~n7422 & ~n7421;
  assign n7423 = ~n7868;
  assign n7424 = ~n7648 | ~n7423;
  assign n7430 = ~n7425 | ~n7424;
  assign n7428 = n7427 ^ ~n7426;
  assign n7429 = ~n7706 & ~n7428;
  assign n7872 = ~n7430 & ~n7429;
  assign n7432 = ~n7431 | ~n7872;
  assign n7434 = ~n7433 & ~n7432;
  assign n7437 = ~n7698 & ~n7434;
  assign n7436 = ~n7435 & ~n7632;
  assign n7439 = ~n7437 & ~n7436;
  assign n7438 = ~REG2_REG_10__SCAN_IN | ~n7698;
  assign U3280 = ~n7439 | ~n7438;
  assign n7442 = ~n7698 | ~REG2_REG_9__SCAN_IN;
  assign n7441 = n7632 | n7440;
  assign n7445 = ~n7442 | ~n7441;
  assign n7859 = n7443 ^ ~n7452;
  assign n7444 = ~n7859 & ~n7642;
  assign n7464 = ~n7445 & ~n7444;
  assign n7860 = n7446 ^ ~n7448;
  assign n7462 = ~n7860 & ~n7702;
  assign n7449 = n7447 ^ n7448;
  assign n7458 = ~n7449 | ~n7678;
  assign n7456 = ~n7450 & ~n7573;
  assign n7454 = ~n7451 | ~n7533;
  assign n7453 = ~n7714 | ~n7452;
  assign n7455 = ~n7454 | ~n7453;
  assign n7457 = ~n7456 & ~n7455;
  assign n7460 = ~n7458 | ~n7457;
  assign n7459 = ~n7860 & ~n7707;
  assign n7864 = ~n7460 & ~n7459;
  assign n7461 = ~n7698 & ~n7864;
  assign n7463 = ~n7462 & ~n7461;
  assign U3281 = ~n7464 | ~n7463;
  assign n7467 = ~n7465 & ~n7632;
  assign n7466 = n7698 & REG2_REG_8__SCAN_IN;
  assign n7494 = ~n7467 & ~n7466;
  assign n7469 = n4397 | n7468;
  assign n7848 = ~n7443 | ~n7469;
  assign n7489 = ~n7848 & ~n7572;
  assign n7485 = ~n7470 & ~n7573;
  assign n7483 = ~n7714 | ~n7471;
  assign n7540 = ~n7472 | ~n7558;
  assign n7475 = ~n7540 | ~n7473;
  assign n7476 = ~n7475 | ~n7474;
  assign n7477 = n7476 ^ ~n7479;
  assign n7481 = ~n7706 & ~n7477;
  assign n7851 = n7478 ^ ~n7479;
  assign n7480 = ~n7707 & ~n7851;
  assign n7482 = ~n7481 & ~n7480;
  assign n7484 = ~n7483 | ~n7482;
  assign n7488 = ~n7485 & ~n7484;
  assign n7487 = ~n7486 | ~n7533;
  assign n7850 = ~n7488 | ~n7487;
  assign n7490 = ~n7489 & ~n7850;
  assign n7492 = ~n7698 & ~n7490;
  assign n7491 = ~n7851 & ~n7702;
  assign n7493 = ~n7492 & ~n7491;
  assign U3282 = ~n7494 | ~n7493;
  assign n7497 = ~n7540 | ~n7495;
  assign n7498 = ~n7497 | ~n7496;
  assign n7500 = n7498 | n7512;
  assign n7499 = ~n7498 | ~n7512;
  assign n7501 = ~n7500 | ~n7499;
  assign n7510 = ~n7501 | ~n7678;
  assign n7508 = ~n7502 & ~n7573;
  assign n7506 = ~n7503 | ~n7533;
  assign n7505 = ~n7714 | ~n7504;
  assign n7507 = ~n7506 | ~n7505;
  assign n7509 = ~n7508 & ~n7507;
  assign n7841 = ~n7510 | ~n7509;
  assign n7843 = n7511 ^ ~n7512;
  assign n7518 = ~n7843 | ~n7513;
  assign n7515 = n4390 ^ ~n7514;
  assign n7842 = ~n7515 & ~n7858;
  assign n7517 = ~n7842 | ~n7516;
  assign n7519 = ~n7518 | ~n7517;
  assign n7520 = ~n7841 & ~n7519;
  assign n7523 = ~n7698 & ~n7520;
  assign n7522 = ~n7632 & ~n7521;
  assign n7525 = ~n7523 & ~n7522;
  assign n7524 = ~REG2_REG_7__SCAN_IN | ~n7698;
  assign U3283 = ~n7525 | ~n7524;
  assign n7833 = n7526 ^ ~n7539;
  assign n7528 = ~n7833;
  assign n7531 = ~n7528 | ~n7527;
  assign n7836 = n4587 ^ ~n7529;
  assign n7530 = ~n7836 | ~n7665;
  assign n7550 = ~n7531 | ~n7530;
  assign n7538 = ~n7532 & ~n7573;
  assign n7536 = ~n7583 | ~n7533;
  assign n7535 = ~n7714 | ~n7534;
  assign n7537 = ~n7536 | ~n7535;
  assign n7545 = ~n7538 & ~n7537;
  assign n7541 = n7540 ^ ~n7539;
  assign n7543 = ~n7541 & ~n7706;
  assign n7542 = ~n7833 & ~n7707;
  assign n7544 = ~n7543 & ~n7542;
  assign n7835 = ~n7545 | ~n7544;
  assign n7547 = ~n7546 & ~n7632;
  assign n7548 = ~n7835 & ~n7547;
  assign n7549 = ~n7698 & ~n7548;
  assign n7552 = ~n7550 & ~n7549;
  assign n7551 = ~REG2_REG_6__SCAN_IN | ~n7698;
  assign U3284 = ~n7552 | ~n7551;
  assign n7555 = REG2_REG_5__SCAN_IN & n7698;
  assign n7554 = ~n7632 & ~n7553;
  assign n7581 = ~n7555 & ~n7554;
  assign n7559 = ~n5498 | ~n7558;
  assign n7826 = n7556 ^ ~n7559;
  assign n7569 = ~n7826 & ~n7707;
  assign n7561 = n7560 ^ ~n7559;
  assign n7567 = ~n7561 | ~n7678;
  assign n7562 = ~n7617;
  assign n7565 = ~n7562 & ~n7668;
  assign n7564 = ~n7671 & ~n7563;
  assign n7566 = ~n7565 & ~n7564;
  assign n7568 = ~n7567 | ~n7566;
  assign n7830 = ~n7569 & ~n7568;
  assign n7823 = n7570 ^ ~n7571;
  assign n7575 = ~n7823 & ~n7572;
  assign n7824 = ~n7574 & ~n7573;
  assign n7576 = ~n7575 & ~n7824;
  assign n7577 = n7830 & n7576;
  assign n7579 = ~n7698 & ~n7577;
  assign n7578 = ~n7826 & ~n7702;
  assign n7580 = ~n7579 & ~n7578;
  assign U3285 = ~n7581 | ~n7580;
  assign n7588 = ~n7582 & ~n7668;
  assign n7586 = ~n7583 | ~n7709;
  assign n7585 = ~n7714 | ~n7584;
  assign n7587 = ~n7586 | ~n7585;
  assign n7596 = ~n7588 & ~n7587;
  assign n7590 = n7589 ^ ~n7592;
  assign n7594 = ~n7590 & ~n7706;
  assign n7816 = n7591 ^ ~n7592;
  assign n7593 = ~n7816 & ~n7707;
  assign n7595 = ~n7594 & ~n7593;
  assign n7818 = ~n7596 | ~n7595;
  assign n7597 = ~n7816 & ~n7691;
  assign n7606 = ~n7818 & ~n7597;
  assign n7600 = ~n7598 & ~n7599;
  assign n7601 = ~n7600 & ~n7858;
  assign n7819 = ~n7601 | ~n7570;
  assign n7604 = ~n7819 & ~n7712;
  assign n7603 = ~n7632 & ~n7602;
  assign n7605 = ~n7604 & ~n7603;
  assign n7607 = ~n7606 | ~n7605;
  assign n7610 = ~n7608 | ~n7607;
  assign n7609 = ~n7698 | ~REG2_REG_4__SCAN_IN;
  assign U3286 = ~n7610 | ~n7609;
  assign n7808 = n7612 ^ ~n7611;
  assign n7627 = ~n7808 | ~n7613;
  assign n7616 = n7615 ^ ~n7614;
  assign n7626 = ~n7616 & ~n7706;
  assign n7624 = ~n7808 | ~n7648;
  assign n7622 = ~n5581 & ~n7668;
  assign n7620 = ~n7617 | ~n7709;
  assign n7619 = ~n7714 | ~n7618;
  assign n7621 = ~n7620 | ~n7619;
  assign n7623 = ~n7622 & ~n7621;
  assign n7625 = ~n7624 | ~n7623;
  assign n7813 = ~n7626 & ~n7625;
  assign n7628 = ~n7627 | ~n7813;
  assign n7636 = ~n7628 | ~n7608;
  assign n7809 = n7641 ^ ~n7629;
  assign n7631 = ~n7665 | ~n7809;
  assign n7630 = ~n7698 | ~REG2_REG_3__SCAN_IN;
  assign n7634 = ~n7631 | ~n7630;
  assign n7633 = ~REG3_REG_3__SCAN_IN & ~n7632;
  assign n7635 = ~n7634 & ~n7633;
  assign U3287 = ~n7636 | ~n7635;
  assign n7638 = ~n7698 | ~REG2_REG_2__SCAN_IN;
  assign n7637 = ~n7699 | ~REG3_REG_2__SCAN_IN;
  assign n7644 = ~n7638 | ~n7637;
  assign n7639 = ~n7670 | ~n5568;
  assign n7640 = ~n7652 | ~n7639;
  assign n7800 = ~n7641 | ~n7640;
  assign n7643 = ~n7642 & ~n7800;
  assign n7664 = ~n7644 & ~n7643;
  assign n7801 = n5577 ^ n7645;
  assign n7662 = ~n7801 & ~n7702;
  assign n7647 = n7646 ^ n5577;
  assign n7660 = ~n7647 & ~n7706;
  assign n7649 = ~n7801;
  assign n7658 = ~n7649 | ~n7648;
  assign n7656 = ~n7650 & ~n7668;
  assign n7654 = ~n7651 | ~n7709;
  assign n7653 = ~n7714 | ~n7652;
  assign n7655 = ~n7654 | ~n7653;
  assign n7657 = ~n7656 & ~n7655;
  assign n7659 = ~n7658 | ~n7657;
  assign n7805 = ~n7660 & ~n7659;
  assign n7661 = ~n7698 & ~n7805;
  assign n7663 = ~n7662 & ~n7661;
  assign U3288 = ~n7664 | ~n7663;
  assign n7795 = n4729 ^ ~n5568;
  assign n7667 = ~n7665 | ~n7795;
  assign n7666 = ~n7699 | ~REG3_REG_1__SCAN_IN;
  assign n7695 = ~n7667 | ~n7666;
  assign n7673 = ~n7669 & ~n7668;
  assign n7672 = ~n7671 & ~n7670;
  assign n7690 = ~n7673 & ~n7672;
  assign n7675 = ~n7674;
  assign n7677 = ~n7684 | ~n7675;
  assign n7679 = ~n7677 | ~n7676;
  assign n7682 = ~n7679 | ~n7678;
  assign n7681 = ~n7680 | ~n7709;
  assign n7688 = ~n7682 | ~n7681;
  assign n7686 = n7684 | n7683;
  assign n7792 = ~n7686 | ~n7685;
  assign n7687 = ~n7792 & ~n7707;
  assign n7689 = ~n7688 & ~n7687;
  assign n7794 = ~n7690 | ~n7689;
  assign n7692 = ~n7792 & ~n7691;
  assign n7693 = ~n7794 & ~n7692;
  assign n7694 = ~n7698 & ~n7693;
  assign n7697 = ~n7695 & ~n7694;
  assign n7696 = ~REG2_REG_1__SCAN_IN | ~n7698;
  assign U3289 = ~n7697 | ~n7696;
  assign n7701 = ~n7698 | ~REG2_REG_0__SCAN_IN;
  assign n7700 = ~n7699 | ~REG3_REG_0__SCAN_IN;
  assign n7705 = ~n7701 | ~n7700;
  assign n7704 = ~n7703 & ~n7702;
  assign n7719 = ~n7705 & ~n7704;
  assign n7708 = ~n7707 | ~n7706;
  assign n7711 = ~n7787 | ~n7708;
  assign n7710 = ~n5496 | ~n7709;
  assign n7786 = ~n7711 | ~n7710;
  assign n7713 = ~n7712 & ~n7784;
  assign n7715 = ~n7714 & ~n7713;
  assign n7716 = ~n7715 & ~n5568;
  assign n7717 = n7786 | n7716;
  assign n7718 = ~n7717 | ~n7608;
  assign U3290 = ~n7719 | ~n7718;
  assign n7779 = ~n7721 | ~n7720;
  assign U3291 = D_REG_31__SCAN_IN & n7779;
  assign U3292 = D_REG_30__SCAN_IN & n7779;
  assign U3293 = D_REG_29__SCAN_IN & n7779;
  assign U3294 = D_REG_28__SCAN_IN & n7779;
  assign U3295 = D_REG_27__SCAN_IN & n7779;
  assign U3296 = D_REG_26__SCAN_IN & n7779;
  assign U3297 = D_REG_25__SCAN_IN & n7779;
  assign U3298 = D_REG_24__SCAN_IN & n7779;
  assign U3299 = D_REG_23__SCAN_IN & n7779;
  assign U3300 = D_REG_22__SCAN_IN & n7779;
  assign U3301 = D_REG_21__SCAN_IN & n7779;
  assign U3302 = D_REG_20__SCAN_IN & n7779;
  assign U3303 = D_REG_19__SCAN_IN & n7779;
  assign U3304 = D_REG_18__SCAN_IN & n7779;
  assign U3305 = D_REG_17__SCAN_IN & n7779;
  assign U3306 = D_REG_16__SCAN_IN & n7779;
  assign U3307 = D_REG_15__SCAN_IN & n7779;
  assign U3308 = D_REG_14__SCAN_IN & n7779;
  assign U3309 = D_REG_13__SCAN_IN & n7779;
  assign U3310 = D_REG_12__SCAN_IN & n7779;
  assign U3311 = D_REG_11__SCAN_IN & n7779;
  assign U3312 = D_REG_10__SCAN_IN & n7779;
  assign U3313 = D_REG_9__SCAN_IN & n7779;
  assign U3314 = D_REG_8__SCAN_IN & n7779;
  assign U3315 = D_REG_7__SCAN_IN & n7779;
  assign U3316 = D_REG_6__SCAN_IN & n7779;
  assign U3317 = D_REG_5__SCAN_IN & n7779;
  assign U3318 = D_REG_4__SCAN_IN & n7779;
  assign U3319 = D_REG_3__SCAN_IN & n7779;
  assign U3320 = D_REG_2__SCAN_IN & n7779;
  assign n7724 = ~n7723 | ~STATE_REG_SCAN_IN;
  assign n7725 = ~n7722 & ~n7724;
  assign n7727 = ~IR_REG_31__SCAN_IN | ~n7725;
  assign n7726 = ~DATAI_31_ | ~U3149;
  assign U3321 = ~n7727 | ~n7726;
  assign n7728 = ~STATE_REG_SCAN_IN & ~DATAI_23_;
  assign U3329 = ~n7774 & ~n7728;
  assign n7731 = ~STATE_REG_SCAN_IN | ~n7729;
  assign n7730 = ~DATAI_18_ | ~U3149;
  assign U3334 = ~n7731 | ~n7730;
  assign n7734 = ~STATE_REG_SCAN_IN | ~n7732;
  assign n7733 = ~DATAI_17_ | ~U3149;
  assign U3335 = ~n7734 | ~n7733;
  assign n7737 = ~STATE_REG_SCAN_IN | ~n7735;
  assign n7736 = ~DATAI_16_ | ~U3149;
  assign U3336 = ~n7737 | ~n7736;
  assign n7740 = ~STATE_REG_SCAN_IN | ~n7738;
  assign n7739 = ~DATAI_15_ | ~U3149;
  assign U3337 = ~n7740 | ~n7739;
  assign n7743 = ~STATE_REG_SCAN_IN | ~n7741;
  assign n7742 = ~DATAI_14_ | ~U3149;
  assign U3338 = ~n7743 | ~n7742;
  assign n7746 = ~STATE_REG_SCAN_IN | ~n7744;
  assign n7745 = ~DATAI_13_ | ~U3149;
  assign U3339 = ~n7746 | ~n7745;
  assign n7749 = ~STATE_REG_SCAN_IN | ~n7747;
  assign n7748 = ~DATAI_12_ | ~U3149;
  assign U3340 = ~n7749 | ~n7748;
  assign n7752 = ~STATE_REG_SCAN_IN | ~n7750;
  assign n7751 = ~DATAI_11_ | ~U3149;
  assign U3341 = ~n7752 | ~n7751;
  assign n7755 = ~STATE_REG_SCAN_IN | ~n7753;
  assign n7754 = ~DATAI_10_ | ~U3149;
  assign U3342 = ~n7755 | ~n7754;
  assign n7758 = ~STATE_REG_SCAN_IN | ~n7756;
  assign n7757 = ~DATAI_9_ | ~U3149;
  assign U3343 = ~n7758 | ~n7757;
  assign n7761 = ~STATE_REG_SCAN_IN | ~n7759;
  assign n7760 = ~DATAI_8_ | ~U3149;
  assign U3344 = ~n7761 | ~n7760;
  assign n7764 = ~STATE_REG_SCAN_IN | ~n7762;
  assign n7763 = ~DATAI_7_ | ~U3149;
  assign U3345 = ~n7764 | ~n7763;
  assign n7767 = ~STATE_REG_SCAN_IN | ~n7765;
  assign n7766 = ~DATAI_6_ | ~U3149;
  assign U3346 = ~n7767 | ~n7766;
  assign n7770 = ~STATE_REG_SCAN_IN | ~n7768;
  assign n7769 = ~DATAI_5_ | ~U3149;
  assign U3347 = ~n7770 | ~n7769;
  assign n7772 = ~IR_REG_0__SCAN_IN | ~STATE_REG_SCAN_IN;
  assign n7771 = ~DATAI_0_ | ~U3149;
  assign U3352 = ~n7772 | ~n7771;
  assign n7775 = ~n7774 | ~n7773;
  assign n7778 = ~n7776 & ~n7775;
  assign n7781 = ~n7779;
  assign n7777 = ~D_REG_0__SCAN_IN & ~n7781;
  assign U3458 = ~n7778 & ~n7777;
  assign n7783 = ~D_REG_1__SCAN_IN | ~n7779;
  assign n7782 = ~n7781 | ~n7780;
  assign U3459 = ~n7783 | ~n7782;
  assign n7791 = ~REG0_REG_0__SCAN_IN | ~n7900;
  assign n7785 = ~n5568 & ~n7784;
  assign n7789 = ~n7786 & ~n7785;
  assign n7788 = ~n7787 | ~n7852;
  assign n7910 = ~n7789 | ~n7788;
  assign n7790 = ~n7907 | ~n7910;
  assign U3467 = ~n7791 | ~n7790;
  assign n7799 = ~REG0_REG_1__SCAN_IN | ~n7900;
  assign n7793 = ~n7792 & ~n7901;
  assign n7797 = ~n7794 & ~n7793;
  assign n7796 = ~n7795 | ~n7883;
  assign n7913 = ~n7797 | ~n7796;
  assign n7798 = ~n7907 | ~n7913;
  assign U3469 = ~n7799 | ~n7798;
  assign n7807 = ~REG0_REG_2__SCAN_IN | ~n7900;
  assign n7803 = ~n7800 & ~n7858;
  assign n7802 = ~n7801 & ~n7901;
  assign n7804 = ~n7803 & ~n7802;
  assign n7916 = ~n7805 | ~n7804;
  assign n7806 = ~n7907 | ~n7916;
  assign U3471 = ~n7807 | ~n7806;
  assign n7815 = ~REG0_REG_3__SCAN_IN | ~n7900;
  assign n7811 = ~n7808 | ~n7852;
  assign n7810 = ~n7809 | ~n7883;
  assign n7812 = n7811 & n7810;
  assign n7919 = ~n7813 | ~n7812;
  assign n7814 = ~n7907 | ~n7919;
  assign U3473 = ~n7815 | ~n7814;
  assign n7822 = ~REG0_REG_4__SCAN_IN | ~n7900;
  assign n7817 = ~n7816 & ~n7901;
  assign n7820 = ~n7818 & ~n7817;
  assign n7922 = ~n7820 | ~n7819;
  assign n7821 = ~n7907 | ~n7922;
  assign U3475 = ~n7822 | ~n7821;
  assign n7832 = ~REG0_REG_5__SCAN_IN | ~n7900;
  assign n7825 = ~n7823 & ~n7858;
  assign n7828 = n7825 | n7824;
  assign n7827 = ~n7826 & ~n7901;
  assign n7829 = ~n7828 & ~n7827;
  assign n7925 = ~n7830 | ~n7829;
  assign n7831 = ~n7907 | ~n7925;
  assign U3477 = ~n7832 | ~n7831;
  assign n7840 = ~REG0_REG_6__SCAN_IN | ~n7900;
  assign n7834 = ~n7833 & ~n7901;
  assign n7838 = ~n7835 & ~n7834;
  assign n7837 = ~n7836 | ~n7883;
  assign n7928 = ~n7838 | ~n7837;
  assign n7839 = ~n7907 | ~n7928;
  assign U3479 = ~n7840 | ~n7839;
  assign n7847 = ~REG0_REG_7__SCAN_IN | ~n7900;
  assign n7845 = ~n7842 & ~n7841;
  assign n7844 = ~n7843 | ~n7887;
  assign n7931 = ~n7845 | ~n7844;
  assign n7846 = ~n7907 | ~n7931;
  assign U3481 = ~n7847 | ~n7846;
  assign n7857 = ~REG0_REG_8__SCAN_IN | ~n7900;
  assign n7849 = ~n7848 & ~n7858;
  assign n7855 = ~n7850 & ~n7849;
  assign n7853 = ~n7851;
  assign n7854 = ~n7853 | ~n7852;
  assign n7934 = ~n7855 | ~n7854;
  assign n7856 = ~n7907 | ~n7934;
  assign U3483 = ~n7857 | ~n7856;
  assign n7866 = ~REG0_REG_9__SCAN_IN | ~n7900;
  assign n7862 = ~n7859 & ~n7858;
  assign n7861 = ~n7860 & ~n7901;
  assign n7863 = ~n7862 & ~n7861;
  assign n7937 = ~n7864 | ~n7863;
  assign n7865 = ~n7907 | ~n7937;
  assign U3485 = ~n7866 | ~n7865;
  assign n7874 = ~REG0_REG_10__SCAN_IN | ~n7900;
  assign n7870 = n7867 & n7883;
  assign n7869 = ~n7868 & ~n7901;
  assign n7871 = ~n7870 & ~n7869;
  assign n7940 = ~n7872 | ~n7871;
  assign n7873 = ~n7907 | ~n7940;
  assign U3487 = ~n7874 | ~n7873;
  assign n7882 = ~REG0_REG_11__SCAN_IN | ~n7900;
  assign n7878 = n7875 & n7883;
  assign n7877 = ~n7876 & ~n7901;
  assign n7879 = ~n7878 & ~n7877;
  assign n7943 = ~n7880 | ~n7879;
  assign n7881 = ~n7907 | ~n7943;
  assign U3489 = ~n7882 | ~n7881;
  assign n7892 = ~REG0_REG_12__SCAN_IN | ~n7900;
  assign n7885 = n7884 & n7883;
  assign n7890 = ~n7886 & ~n7885;
  assign n7889 = ~n7888 | ~n7887;
  assign n7946 = ~n7890 | ~n7889;
  assign n7891 = ~n7907 | ~n7946;
  assign U3491 = ~n7892 | ~n7891;
  assign n7899 = ~REG0_REG_13__SCAN_IN | ~n7900;
  assign n7894 = ~n7893 & ~n7901;
  assign n7896 = ~n7895 & ~n7894;
  assign n7949 = ~n7897 | ~n7896;
  assign n7898 = ~n7907 | ~n7949;
  assign U3493 = ~n7899 | ~n7898;
  assign n7909 = ~REG0_REG_14__SCAN_IN | ~n7900;
  assign n7903 = ~n7902 & ~n7901;
  assign n7905 = ~n7904 & ~n7903;
  assign n7953 = ~n7906 | ~n7905;
  assign n7908 = ~n7907 | ~n7953;
  assign U3495 = ~n7909 | ~n7908;
  assign n7912 = ~REG1_REG_0__SCAN_IN | ~n7952;
  assign n7911 = ~n7954 | ~n7910;
  assign U3518 = ~n7912 | ~n7911;
  assign n7915 = ~REG1_REG_1__SCAN_IN | ~n7952;
  assign n7914 = ~n7954 | ~n7913;
  assign U3519 = ~n7915 | ~n7914;
  assign n7918 = ~REG1_REG_2__SCAN_IN | ~n7952;
  assign n7917 = ~n7954 | ~n7916;
  assign U3520 = ~n7918 | ~n7917;
  assign n7921 = ~REG1_REG_3__SCAN_IN | ~n7952;
  assign n7920 = ~n7954 | ~n7919;
  assign U3521 = ~n7921 | ~n7920;
  assign n7924 = ~REG1_REG_4__SCAN_IN | ~n7952;
  assign n7923 = ~n7954 | ~n7922;
  assign U3522 = ~n7924 | ~n7923;
  assign n7927 = ~REG1_REG_5__SCAN_IN | ~n7952;
  assign n7926 = ~n7954 | ~n7925;
  assign U3523 = ~n7927 | ~n7926;
  assign n7930 = ~REG1_REG_6__SCAN_IN | ~n7952;
  assign n7929 = ~n7954 | ~n7928;
  assign U3524 = ~n7930 | ~n7929;
  assign n7933 = ~REG1_REG_7__SCAN_IN | ~n7952;
  assign n7932 = ~n7954 | ~n7931;
  assign U3525 = ~n7933 | ~n7932;
  assign n7936 = ~REG1_REG_8__SCAN_IN | ~n7952;
  assign n7935 = ~n7954 | ~n7934;
  assign U3526 = ~n7936 | ~n7935;
  assign n7939 = ~REG1_REG_9__SCAN_IN | ~n7952;
  assign n7938 = ~n7954 | ~n7937;
  assign U3527 = ~n7939 | ~n7938;
  assign n7942 = ~REG1_REG_10__SCAN_IN | ~n7952;
  assign n7941 = ~n7954 | ~n7940;
  assign U3528 = ~n7942 | ~n7941;
  assign n7945 = ~REG1_REG_11__SCAN_IN | ~n7952;
  assign n7944 = ~n7954 | ~n7943;
  assign U3529 = ~n7945 | ~n7944;
  assign n7948 = ~REG1_REG_12__SCAN_IN | ~n7952;
  assign n7947 = ~n7954 | ~n7946;
  assign U3530 = ~n7948 | ~n7947;
  assign n7951 = ~REG1_REG_13__SCAN_IN | ~n7952;
  assign n7950 = ~n7954 | ~n7949;
  assign U3531 = ~n7951 | ~n7950;
  assign n7956 = ~REG1_REG_14__SCAN_IN | ~n7952;
  assign n7955 = ~n7954 | ~n7953;
  assign U3532 = ~n7956 | ~n7955;
  assign n7960 = ~n8000 | ~DATAO_REG_16__SCAN_IN;
  assign n7959 = ~n7958 | ~n7957;
  assign U3566 = ~n7960 | ~n7959;
  assign n7963 = ~n8000 | ~DATAO_REG_17__SCAN_IN;
  assign n7962 = ~n7961 | ~U4043;
  assign U3567 = ~n7963 | ~n7962;
  assign n7966 = ~n8000 | ~DATAO_REG_18__SCAN_IN;
  assign n7965 = ~n7964 | ~U4043;
  assign U3568 = ~n7966 | ~n7965;
  assign n7969 = ~n8000 | ~DATAO_REG_19__SCAN_IN;
  assign n7968 = ~n7967 | ~U4043;
  assign U3569 = ~n7969 | ~n7968;
  assign n7972 = ~n8000 | ~DATAO_REG_20__SCAN_IN;
  assign n7971 = ~n7970 | ~U4043;
  assign U3570 = ~n7972 | ~n7971;
  assign n7975 = ~n8000 | ~DATAO_REG_21__SCAN_IN;
  assign n7974 = ~n7973 | ~U4043;
  assign U3571 = ~n7975 | ~n7974;
  assign n7978 = ~n8000 | ~DATAO_REG_22__SCAN_IN;
  assign n7977 = ~n7976 | ~U4043;
  assign U3572 = ~n7978 | ~n7977;
  assign n7981 = ~n8000 | ~DATAO_REG_23__SCAN_IN;
  assign n7980 = ~n7979 | ~U4043;
  assign U3573 = ~n7981 | ~n7980;
  assign n7984 = ~n8000 | ~DATAO_REG_24__SCAN_IN;
  assign n7983 = ~n7982 | ~U4043;
  assign U3574 = ~n7984 | ~n7983;
  assign n7987 = ~n8000 | ~DATAO_REG_25__SCAN_IN;
  assign n7986 = ~n7985 | ~U4043;
  assign U3575 = ~n7987 | ~n7986;
  assign n7990 = ~n8005 | ~DATAO_REG_26__SCAN_IN;
  assign n7989 = ~n7988 | ~U4043;
  assign U3576 = ~n7990 | ~n7989;
  assign n7993 = ~n8000 | ~DATAO_REG_27__SCAN_IN;
  assign n7992 = ~n7991 | ~U4043;
  assign U3577 = ~n7993 | ~n7992;
  assign n7996 = ~n8000 | ~DATAO_REG_28__SCAN_IN;
  assign n7995 = ~n7994 | ~U4043;
  assign U3578 = ~n7996 | ~n7995;
  assign n7999 = ~n8000 | ~DATAO_REG_29__SCAN_IN;
  assign n7998 = ~n7997 | ~U4043;
  assign U3579 = ~n7999 | ~n7998;
  assign n8004 = ~n8000 | ~DATAO_REG_30__SCAN_IN;
  assign n8002 = ~n8001;
  assign n8003 = ~n8002 | ~U4043;
  assign U3580 = ~n8004 | ~n8003;
  assign n8008 = ~n8005 | ~DATAO_REG_31__SCAN_IN;
  assign n8007 = ~n8006 | ~U4043;
  assign U3581 = ~n8008 | ~n8007;
  assign n5752 = n4545 & n4544;
endmodule


