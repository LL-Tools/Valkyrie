

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput127, keyinput126, keyinput125, keyinput124, keyinput123, 
        keyinput122, keyinput121, keyinput120, keyinput119, keyinput118, 
        keyinput117, keyinput116, keyinput115, keyinput114, keyinput113, 
        keyinput112, keyinput111, keyinput110, keyinput109, keyinput108, 
        keyinput107, keyinput106, keyinput105, keyinput104, keyinput103, 
        keyinput102, keyinput101, keyinput100, keyinput99, keyinput98, 
        keyinput97, keyinput96, keyinput95, keyinput94, keyinput93, keyinput92, 
        keyinput91, keyinput90, keyinput89, keyinput88, keyinput87, keyinput86, 
        keyinput85, keyinput84, keyinput83, keyinput82, keyinput81, keyinput80, 
        keyinput79, keyinput78, keyinput77, keyinput76, keyinput75, keyinput74, 
        keyinput73, keyinput72, keyinput71, keyinput70, keyinput69, keyinput68, 
        keyinput67, keyinput66, keyinput65, keyinput64, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4401, n4403, n4404, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415;

  AND2_X1 U4907 ( .A1(n4892), .A2(n4437), .ZN(n8601) );
  NAND2_X1 U4908 ( .A1(n8164), .A2(n8163), .ZN(n8375) );
  OR2_X1 U4909 ( .A1(n8412), .A2(n4857), .ZN(n4856) );
  AND2_X1 U4910 ( .A1(n5944), .A2(n7363), .ZN(n5930) );
  CLKBUF_X2 U4911 ( .A(n7453), .Z(n8201) );
  CLKBUF_X2 U4912 ( .A(n5250), .Z(n5579) );
  INV_X2 U4913 ( .A(n6138), .ZN(n6370) );
  NAND3_X2 U4914 ( .A1(n6104), .A2(n6103), .A3(n6102), .ZN(n6893) );
  CLKBUF_X2 U4915 ( .A(n6114), .Z(n6299) );
  XNOR2_X1 U4916 ( .A(n5038), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7363) );
  CLKBUF_X2 U4917 ( .A(n6109), .Z(n6133) );
  CLKBUF_X3 U4918 ( .A(n6956), .Z(n9089) );
  INV_X1 U4919 ( .A(n9062), .ZN(n4409) );
  AOI21_X1 U4921 ( .B1(n8710), .B2(n8717), .A(n4640), .ZN(n8699) );
  INV_X1 U4922 ( .A(n5930), .ZN(n6617) );
  INV_X1 U4923 ( .A(n6959), .ZN(n9165) );
  CLKBUF_X2 U4924 ( .A(n7453), .Z(n4406) );
  OR2_X1 U4925 ( .A1(n5073), .A2(n5058), .ZN(n5070) );
  INV_X1 U4926 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5058) );
  NAND2_X1 U4927 ( .A1(n4819), .A2(n4817), .ZN(n5103) );
  INV_X1 U4928 ( .A(n8392), .ZN(n8702) );
  NAND2_X1 U4929 ( .A1(n6536), .A2(n6127), .ZN(n6974) );
  XNOR2_X1 U4930 ( .A(n6584), .B(P1_IR_REG_22__SCAN_IN), .ZN(n6745) );
  OAI211_X2 U4931 ( .C1(n7201), .C2(n4897), .A(n5105), .B(n4895), .ZN(n10317)
         );
  AND4_X1 U4932 ( .A1(n4521), .A2(n10013), .A3(n4570), .A4(n4569), .ZN(n4401)
         );
  NAND4_X2 U4933 ( .A1(n6132), .A2(n6131), .A3(n6130), .A4(n6129), .ZN(n9318)
         );
  AOI21_X2 U4935 ( .B1(n7083), .B2(n6538), .A(n6151), .ZN(n7242) );
  XNOR2_X2 U4936 ( .A(n5070), .B(n5069), .ZN(n7199) );
  XNOR2_X2 U4937 ( .A(n5059), .B(n4537), .ZN(n8153) );
  NAND2_X2 U4938 ( .A1(n4960), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5059) );
  CLKBUF_X1 U4939 ( .A(n6365), .Z(n4403) );
  BUF_X4 U4940 ( .A(n6365), .Z(n4404) );
  INV_X1 U4941 ( .A(n6097), .ZN(n6365) );
  AND2_X2 U4942 ( .A1(n7242), .A2(n7181), .ZN(n7165) );
  NAND2_X2 U4943 ( .A1(n5082), .A2(n5081), .ZN(n7285) );
  OAI21_X2 U4944 ( .B1(n4852), .B2(n4848), .A(n4845), .ZN(n4853) );
  OAI21_X2 U4945 ( .B1(n8125), .B2(n8035), .A(n8034), .ZN(n9006) );
  NOR2_X2 U4946 ( .A1(n8126), .A2(n8127), .ZN(n8125) );
  NAND2_X2 U4947 ( .A1(n7368), .A2(n7367), .ZN(n7453) );
  XNOR2_X2 U4949 ( .A(n4686), .B(P1_IR_REG_1__SCAN_IN), .ZN(n9324) );
  AOI21_X2 U4951 ( .B1(n9549), .B2(n9551), .A(n9467), .ZN(n9537) );
  AND2_X1 U4952 ( .A1(n4577), .A2(n4575), .ZN(n9704) );
  NAND2_X1 U4953 ( .A1(n8000), .A2(n6251), .ZN(n7998) );
  NOR2_X1 U4954 ( .A1(n7672), .A2(n5011), .ZN(n4418) );
  NAND2_X1 U4955 ( .A1(n7664), .A2(n8132), .ZN(n7388) );
  NAND2_X1 U4956 ( .A1(n6417), .A2(n6537), .ZN(n6999) );
  INV_X1 U4957 ( .A(n9314), .ZN(n7397) );
  INV_X1 U4958 ( .A(n8406), .ZN(n7656) );
  INV_X2 U4959 ( .A(n9319), .ZN(n7012) );
  CLKBUF_X2 U4960 ( .A(n6959), .Z(n4410) );
  NAND3_X1 U4961 ( .A1(n6755), .A2(n6786), .A3(n6724), .ZN(n6959) );
  AND3_X1 U4962 ( .A1(n5108), .A2(n5107), .A3(n5106), .ZN(n10344) );
  CLKBUF_X2 U4963 ( .A(n5104), .Z(n6619) );
  INV_X2 U4966 ( .A(n5103), .ZN(n6624) );
  AND2_X1 U4968 ( .A1(n4607), .A2(n4608), .ZN(n4598) );
  NAND2_X1 U4969 ( .A1(n4909), .A2(n4913), .ZN(n9565) );
  NAND2_X1 U4970 ( .A1(n9078), .A2(n9077), .ZN(n9142) );
  AND2_X1 U4971 ( .A1(n4773), .A2(n4772), .ZN(n5777) );
  NAND2_X1 U4972 ( .A1(n9460), .A2(n4806), .ZN(n9606) );
  NOR2_X1 U4973 ( .A1(n8692), .A2(n5903), .ZN(n8684) );
  AOI21_X1 U4974 ( .B1(n8982), .B2(n5733), .A(n5730), .ZN(n8929) );
  AND2_X1 U4975 ( .A1(n9027), .A2(n9028), .ZN(n9299) );
  NAND2_X1 U4976 ( .A1(n8723), .A2(n4642), .ZN(n8710) );
  NAND2_X1 U4977 ( .A1(n8724), .A2(n8728), .ZN(n8723) );
  AOI21_X1 U4978 ( .B1(n5008), .B2(n4438), .A(n4668), .ZN(n9132) );
  NOR2_X1 U4979 ( .A1(n8734), .A2(n8745), .ZN(n8737) );
  NAND2_X1 U4980 ( .A1(n9716), .A2(n6462), .ZN(n9702) );
  NOR2_X1 U4981 ( .A1(n9390), .A2(n4684), .ZN(n9410) );
  OR2_X1 U4982 ( .A1(n8499), .A2(n8498), .ZN(n8522) );
  NAND2_X1 U4983 ( .A1(n8023), .A2(n4663), .ZN(n8126) );
  NAND2_X1 U4984 ( .A1(n7998), .A2(n4812), .ZN(n9741) );
  AOI21_X1 U4985 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n8466), .A(n8458), .ZN(
        n8492) );
  OR2_X1 U4986 ( .A1(n8482), .A2(n8481), .ZN(n8507) );
  NAND2_X1 U4987 ( .A1(n7833), .A2(n7834), .ZN(n8000) );
  NAND2_X1 U4988 ( .A1(n8434), .A2(n4859), .ZN(n4858) );
  NAND2_X1 U4989 ( .A1(n7742), .A2(n7741), .ZN(n7896) );
  NAND2_X1 U4990 ( .A1(n5362), .A2(n5361), .ZN(n8877) );
  NAND2_X1 U4991 ( .A1(n4519), .A2(n4422), .ZN(n7868) );
  OAI21_X1 U4992 ( .B1(n7792), .B2(n7791), .A(n4861), .ZN(n4864) );
  NAND2_X1 U4993 ( .A1(n5954), .A2(n10345), .ZN(n10350) );
  NAND2_X1 U4994 ( .A1(n6164), .A2(n6163), .ZN(n7664) );
  NAND2_X1 U4995 ( .A1(n7878), .A2(n8085), .ZN(n8079) );
  NAND2_X1 U4996 ( .A1(n6174), .A2(n6173), .ZN(n7578) );
  OR2_X1 U4997 ( .A1(n4573), .A2(n4574), .ZN(n7014) );
  NAND2_X1 U4998 ( .A1(n4644), .A2(n4694), .ZN(n5233) );
  NAND2_X1 U4999 ( .A1(n6094), .A2(n6533), .ZN(n6926) );
  AOI21_X1 U5000 ( .B1(n7547), .B2(n7548), .A(n7549), .ZN(n7686) );
  INV_X1 U5001 ( .A(n5785), .ZN(n7484) );
  CLKBUF_X1 U5002 ( .A(n6748), .Z(n9320) );
  NAND4_X1 U5003 ( .A1(n5115), .A2(n5114), .A3(n5113), .A4(n5112), .ZN(n8406)
         );
  NAND4_X1 U5004 ( .A1(n5096), .A2(n5095), .A3(n5094), .A4(n5093), .ZN(n8407)
         );
  AND2_X1 U5005 ( .A1(n7799), .A2(n6755), .ZN(n4662) );
  OAI211_X1 U5006 ( .C1(n6138), .C2(n6635), .A(n6137), .B(n6136), .ZN(n7106)
         );
  NAND4_X1 U5007 ( .A1(n6083), .A2(n6082), .A3(n6081), .A4(n6080), .ZN(n6748)
         );
  NAND2_X1 U5008 ( .A1(n4595), .A2(n5162), .ZN(n5174) );
  OR2_X1 U5009 ( .A1(n6721), .A2(n6745), .ZN(n6722) );
  NAND2_X1 U5010 ( .A1(n7002), .A2(n6723), .ZN(n7799) );
  OR2_X1 U5011 ( .A1(n5663), .A2(n5662), .ZN(n5664) );
  INV_X1 U5012 ( .A(n6099), .ZN(n6114) );
  CLKBUF_X3 U5013 ( .A(n6095), .Z(n6364) );
  CLKBUF_X3 U5014 ( .A(n6115), .Z(n6366) );
  INV_X2 U5015 ( .A(n6133), .ZN(n6376) );
  AND2_X2 U5016 ( .A1(n5064), .A2(n8989), .ZN(n5128) );
  AND2_X1 U5017 ( .A1(n7751), .A2(n6607), .ZN(n6723) );
  OR2_X1 U5018 ( .A1(n6631), .A2(n6109), .ZN(n4823) );
  NAND2_X1 U5019 ( .A1(n4596), .A2(n5137), .ZN(n5160) );
  NAND2_X1 U5020 ( .A1(n6733), .A2(n6602), .ZN(n6755) );
  INV_X1 U5021 ( .A(n8106), .ZN(n6733) );
  NAND2_X1 U5022 ( .A1(n6532), .A2(n6531), .ZN(n7751) );
  OR2_X1 U5023 ( .A1(n5251), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5273) );
  XNOR2_X1 U5024 ( .A(n6318), .B(n6317), .ZN(n6603) );
  NAND2_X1 U5025 ( .A1(n10219), .A2(n5997), .ZN(n6097) );
  NAND2_X1 U5026 ( .A1(n6384), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6584) );
  NAND2_X1 U5027 ( .A1(n6593), .A2(n6594), .ZN(n8106) );
  NAND2_X1 U5028 ( .A1(n5990), .A2(n5995), .ZN(n10219) );
  XNOR2_X1 U5029 ( .A(n6385), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6607) );
  NAND3_X1 U5030 ( .A1(n4976), .A2(n4977), .A3(n4979), .ZN(n5997) );
  XNOR2_X1 U5031 ( .A(n5061), .B(n4536), .ZN(n8989) );
  OR2_X1 U5032 ( .A1(n6531), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n6384) );
  NAND2_X1 U5033 ( .A1(n5994), .A2(n5993), .ZN(n5995) );
  NAND2_X1 U5034 ( .A1(n6528), .A2(n10010), .ZN(n6531) );
  AND2_X1 U5035 ( .A1(n6383), .A2(n6382), .ZN(n6528) );
  AND2_X2 U5036 ( .A1(n5975), .A2(n5972), .ZN(n5991) );
  NAND2_X2 U5037 ( .A1(n5553), .A2(P1_U3086), .ZN(n10222) );
  NOR2_X1 U5038 ( .A1(n4803), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n4566) );
  NAND2_X1 U5039 ( .A1(n4804), .A2(n5056), .ZN(n4803) );
  INV_X2 U5040 ( .A(n6624), .ZN(n5553) );
  XNOR2_X1 U5041 ( .A(n5141), .B(n5153), .ZN(n7444) );
  AND2_X1 U5042 ( .A1(n4444), .A2(n5024), .ZN(n6382) );
  AND3_X1 U5043 ( .A1(n4954), .A2(n4932), .A3(n4759), .ZN(n4758) );
  CLKBUF_X1 U5044 ( .A(n6107), .Z(n6123) );
  AND4_X1 U5045 ( .A1(n5029), .A2(n9976), .A3(n5031), .A4(n5153), .ZN(n4425)
         );
  NAND2_X1 U5046 ( .A1(n5992), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5993) );
  AND3_X1 U5047 ( .A1(n5050), .A2(n5646), .A3(n5049), .ZN(n5054) );
  AND2_X1 U5048 ( .A1(n6105), .A2(n5968), .ZN(n6107) );
  NAND2_X1 U5049 ( .A1(n5058), .A2(n4896), .ZN(n4895) );
  INV_X1 U5050 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n9976) );
  NOR2_X1 U5051 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n6292) );
  INV_X4 U5052 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U5053 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n10010) );
  NOR2_X1 U5054 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n4521) );
  INV_X1 U5055 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5049) );
  INV_X1 U5056 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5153) );
  INV_X1 U5057 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5646) );
  INV_X1 U5058 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5031) );
  INV_X2 U5059 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U5060 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5229) );
  NOR2_X1 U5061 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5029) );
  NAND2_X1 U5062 ( .A1(n6959), .A2(n9168), .ZN(n4407) );
  NAND2_X1 U5063 ( .A1(n6959), .A2(n9168), .ZN(n6956) );
  AND2_X4 U5064 ( .A1(n8153), .A2(n8989), .ZN(n5110) );
  AND2_X1 U5065 ( .A1(n6755), .A2(n6723), .ZN(n6720) );
  INV_X1 U5066 ( .A(n6720), .ZN(n9062) );
  NAND2_X1 U5067 ( .A1(n4873), .A2(n4461), .ZN(n4871) );
  NAND2_X1 U5068 ( .A1(n9079), .A2(n9267), .ZN(n4963) );
  AND2_X1 U5069 ( .A1(n4921), .A2(n4911), .ZN(n4910) );
  NAND2_X1 U5070 ( .A1(n4913), .A2(n4915), .ZN(n4911) );
  NOR2_X1 U5071 ( .A1(n9502), .A2(n4922), .ZN(n4921) );
  INV_X1 U5072 ( .A(n9500), .ZN(n4922) );
  INV_X1 U5073 ( .A(n9737), .ZN(n9478) );
  NAND2_X1 U5074 ( .A1(n5924), .A2(n5742), .ZN(n5921) );
  OAI21_X1 U5075 ( .B1(n8653), .B2(n8388), .A(n5632), .ZN(n5694) );
  NAND2_X1 U5076 ( .A1(n7199), .A2(n5636), .ZN(n5104) );
  NOR2_X1 U5077 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5032) );
  NOR2_X1 U5078 ( .A1(n8823), .A2(n4561), .ZN(n4560) );
  NOR2_X1 U5079 ( .A1(n5844), .A2(n5760), .ZN(n4561) );
  NOR2_X1 U5080 ( .A1(n5904), .A2(n5903), .ZN(n4556) );
  NAND2_X1 U5081 ( .A1(n4549), .A2(n4548), .ZN(n4547) );
  INV_X1 U5082 ( .A(n4552), .ZN(n4548) );
  INV_X1 U5083 ( .A(n4550), .ZN(n4549) );
  NOR2_X1 U5084 ( .A1(n5921), .A2(n5919), .ZN(n4533) );
  AND2_X1 U5085 ( .A1(n5744), .A2(n5743), .ZN(n5748) );
  NOR2_X1 U5086 ( .A1(n5381), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n5043) );
  INV_X1 U5087 ( .A(n6084), .ZN(n6120) );
  AND2_X1 U5088 ( .A1(n5019), .A2(n5035), .ZN(n5037) );
  INV_X1 U5089 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5035) );
  NAND2_X1 U5090 ( .A1(n4849), .A2(n4855), .ZN(n4848) );
  NAND2_X1 U5091 ( .A1(n4871), .A2(n7534), .ZN(n4869) );
  OR3_X1 U5092 ( .A1(n7217), .A2(n4875), .A3(n7450), .ZN(n4870) );
  OAI21_X1 U5093 ( .B1(n4424), .B2(n4413), .A(n4466), .ZN(n4613) );
  OR2_X1 U5094 ( .A1(n8368), .A2(n8671), .ZN(n5912) );
  AND2_X1 U5095 ( .A1(n8368), .A2(n8671), .ZN(n5913) );
  OR2_X1 U5096 ( .A1(n8285), .A2(n8680), .ZN(n5909) );
  OR2_X1 U5097 ( .A1(n8729), .A2(n8713), .ZN(n5887) );
  OAI21_X1 U5098 ( .B1(n8754), .B2(n5629), .A(n5630), .ZN(n8734) );
  OR2_X1 U5099 ( .A1(n8772), .A2(n8757), .ZN(n5875) );
  NAND3_X1 U5100 ( .A1(n4535), .A2(n4763), .A3(n5068), .ZN(n5782) );
  INV_X1 U5101 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n4759) );
  NAND2_X1 U5102 ( .A1(n5996), .A2(n5997), .ZN(n6099) );
  INV_X1 U5103 ( .A(n4721), .ZN(n4717) );
  OR2_X1 U5104 ( .A1(n10052), .A2(n9528), .ZN(n6403) );
  OR2_X1 U5105 ( .A1(n9532), .A2(n10067), .ZN(n6509) );
  AOI21_X1 U5106 ( .B1(n4914), .B2(n9498), .A(n4454), .ZN(n4913) );
  NAND2_X1 U5107 ( .A1(n5987), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6019) );
  INV_X1 U5108 ( .A(n6056), .ZN(n5987) );
  NAND2_X1 U5109 ( .A1(n9719), .A2(n9725), .ZN(n4576) );
  INV_X1 U5110 ( .A(n5018), .ZN(n4590) );
  NAND2_X1 U5111 ( .A1(n6641), .A2(n5553), .ZN(n6109) );
  NAND2_X1 U5112 ( .A1(n5732), .A2(n4722), .ZN(n4720) );
  XNOR2_X1 U5113 ( .A(n5718), .B(n5717), .ZN(n5721) );
  AND2_X1 U5114 ( .A1(n5571), .A2(n5556), .ZN(n5570) );
  NAND2_X1 U5115 ( .A1(n5552), .A2(n5551), .ZN(n5569) );
  NAND2_X1 U5116 ( .A1(n5971), .A2(n4995), .ZN(n4994) );
  INV_X1 U5117 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4995) );
  AND2_X1 U5118 ( .A1(n5534), .A2(n5519), .ZN(n5532) );
  OAI21_X1 U5119 ( .B1(n5469), .B2(n5468), .A(n5467), .ZN(n5485) );
  AND2_X1 U5120 ( .A1(n5450), .A2(n5438), .ZN(n5448) );
  AOI21_X1 U5121 ( .B1(n4749), .B2(n4752), .A(n4748), .ZN(n4747) );
  INV_X1 U5122 ( .A(n5432), .ZN(n4748) );
  NOR2_X1 U5123 ( .A1(n4753), .A2(n5433), .ZN(n4749) );
  NAND2_X1 U5124 ( .A1(n4752), .A2(n4751), .ZN(n4750) );
  INV_X1 U5125 ( .A(n5433), .ZN(n4751) );
  AOI21_X1 U5126 ( .B1(n4411), .B2(n4738), .A(n4464), .ZN(n4731) );
  INV_X1 U5127 ( .A(n4737), .ZN(n4736) );
  OAI21_X1 U5128 ( .B1(n4740), .B2(n4738), .A(n5281), .ZN(n4737) );
  NAND2_X1 U5129 ( .A1(n4941), .A2(n8398), .ZN(n4940) );
  INV_X1 U5130 ( .A(n7458), .ZN(n4942) );
  AOI21_X1 U5131 ( .B1(n4940), .B2(n4941), .A(n8900), .ZN(n4938) );
  INV_X1 U5132 ( .A(n5128), .ZN(n5640) );
  INV_X1 U5133 ( .A(n5111), .ZN(n5582) );
  MUX2_X1 U5134 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5072), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5075) );
  NAND2_X1 U5135 ( .A1(n4852), .A2(n4851), .ZN(n4850) );
  INV_X1 U5136 ( .A(n8077), .ZN(n4882) );
  OAI22_X1 U5137 ( .A1(n8699), .A2(n8703), .B1(n8393), .B2(n8331), .ZN(n8689)
         );
  NOR2_X1 U5138 ( .A1(n8737), .A2(n4643), .ZN(n8724) );
  AND2_X1 U5139 ( .A1(n8744), .A2(n8725), .ZN(n4643) );
  INV_X1 U5140 ( .A(n5734), .ZN(n5418) );
  INV_X1 U5141 ( .A(n6619), .ZN(n5417) );
  INV_X1 U5142 ( .A(n5117), .ZN(n5733) );
  NAND2_X1 U5143 ( .A1(n5104), .A2(n6624), .ZN(n5117) );
  NAND2_X1 U5144 ( .A1(n5104), .A2(n5553), .ZN(n5139) );
  INV_X1 U5145 ( .A(n5055), .ZN(n4804) );
  NOR2_X1 U5146 ( .A1(n9275), .A2(n4657), .ZN(n4656) );
  INV_X1 U5147 ( .A(n9046), .ZN(n4657) );
  NAND2_X1 U5148 ( .A1(n9186), .A2(n4666), .ZN(n9079) );
  AND2_X1 U5149 ( .A1(n9076), .A2(n9073), .ZN(n4666) );
  NOR2_X1 U5150 ( .A1(n4837), .A2(n9571), .ZN(n9507) );
  OR2_X1 U5151 ( .A1(n10052), .A2(n4838), .ZN(n4837) );
  NOR2_X1 U5152 ( .A1(n9535), .A2(n9469), .ZN(n9520) );
  AND2_X1 U5153 ( .A1(n6509), .A2(n9470), .ZN(n9521) );
  OR2_X1 U5154 ( .A1(n9522), .A2(n9521), .ZN(n9524) );
  NOR2_X1 U5155 ( .A1(n9537), .A2(n9536), .ZN(n9535) );
  INV_X1 U5156 ( .A(n6299), .ZN(n6355) );
  OR2_X1 U5157 ( .A1(n10096), .A2(n9150), .ZN(n9465) );
  NAND2_X1 U5158 ( .A1(n9458), .A2(n9457), .ZN(n9460) );
  INV_X1 U5159 ( .A(n9489), .ZN(n4931) );
  NAND2_X1 U5160 ( .A1(n9741), .A2(n6550), .ZN(n9718) );
  NAND2_X1 U5161 ( .A1(n4904), .A2(n4906), .ZN(n4902) );
  OAI21_X1 U5162 ( .B1(n5975), .B2(n10213), .A(P1_IR_REG_28__SCAN_IN), .ZN(
        n4572) );
  NAND2_X1 U5163 ( .A1(n4746), .A2(n4752), .ZN(n5434) );
  NAND2_X1 U5164 ( .A1(n5396), .A2(n4753), .ZN(n4746) );
  NAND2_X1 U5165 ( .A1(n4777), .A2(n4779), .ZN(n5716) );
  OR2_X1 U5166 ( .A1(n5694), .A2(n4601), .ZN(n4597) );
  NAND2_X1 U5167 ( .A1(n4602), .A2(n8785), .ZN(n4601) );
  NAND2_X1 U5168 ( .A1(n4603), .A2(n4606), .ZN(n4602) );
  NAND2_X1 U5169 ( .A1(n5633), .A2(n4417), .ZN(n4606) );
  NAND2_X1 U5170 ( .A1(n5694), .A2(n4600), .ZN(n4599) );
  NOR2_X1 U5171 ( .A1(n4429), .A2(n8896), .ZN(n4600) );
  INV_X1 U5172 ( .A(n5644), .ZN(n4608) );
  AOI21_X1 U5173 ( .B1(n5698), .B2(n8785), .A(n5697), .ZN(n8647) );
  OR2_X1 U5174 ( .A1(n5696), .A2(n5695), .ZN(n5697) );
  OAI21_X1 U5175 ( .B1(n6526), .B2(n4726), .A(n4729), .ZN(n6591) );
  NAND2_X1 U5176 ( .A1(n4471), .A2(n7002), .ZN(n4726) );
  NAND2_X1 U5177 ( .A1(n6527), .A2(n4408), .ZN(n4729) );
  NAND2_X1 U5178 ( .A1(n4559), .A2(n5847), .ZN(n4558) );
  NAND2_X1 U5179 ( .A1(n4560), .A2(n4456), .ZN(n4559) );
  NAND2_X1 U5180 ( .A1(n6469), .A2(n4523), .ZN(n6470) );
  AOI21_X1 U5181 ( .B1(n6467), .B2(n6505), .A(n4426), .ZN(n4523) );
  AOI21_X1 U5182 ( .B1(n4470), .B2(n4556), .A(n4427), .ZN(n4550) );
  AND2_X1 U5183 ( .A1(n4555), .A2(n4553), .ZN(n4552) );
  NOR2_X1 U5184 ( .A1(n5904), .A2(n6617), .ZN(n4555) );
  NAND2_X1 U5185 ( .A1(n5902), .A2(n4554), .ZN(n4553) );
  INV_X1 U5186 ( .A(n5898), .ZN(n4554) );
  AOI21_X1 U5187 ( .B1(n5572), .B2(n5571), .A(n4704), .ZN(n4703) );
  INV_X1 U5188 ( .A(n5586), .ZN(n4704) );
  INV_X1 U5189 ( .A(n5571), .ZN(n4700) );
  INV_X1 U5190 ( .A(n4779), .ZN(n4776) );
  INV_X1 U5191 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n4982) );
  INV_X1 U5192 ( .A(n5448), .ZN(n4745) );
  NAND2_X1 U5193 ( .A1(n5265), .A2(n5264), .ZN(n5281) );
  AND2_X1 U5194 ( .A1(n8264), .A2(n8261), .ZN(n8234) );
  OR2_X1 U5195 ( .A1(n7362), .A2(n5013), .ZN(n7365) );
  OR2_X1 U5196 ( .A1(n5921), .A2(n5922), .ZN(n4531) );
  NAND2_X1 U5197 ( .A1(n4529), .A2(n8651), .ZN(n4528) );
  INV_X1 U5198 ( .A(n4531), .ZN(n4529) );
  NAND2_X1 U5199 ( .A1(n4534), .A2(n4533), .ZN(n4532) );
  NAND2_X1 U5200 ( .A1(n4534), .A2(n4530), .ZN(n5932) );
  AND2_X1 U5201 ( .A1(n4533), .A2(n5923), .ZN(n4530) );
  AOI21_X1 U5202 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n7687), .A(n7686), .ZN(
        n7688) );
  OR2_X1 U5203 ( .A1(n5688), .A2(n8211), .ZN(n5924) );
  OR2_X1 U5204 ( .A1(n8317), .A2(n8691), .ZN(n5901) );
  OR2_X1 U5205 ( .A1(n8868), .A2(n8769), .ZN(n5876) );
  INV_X1 U5206 ( .A(n4796), .ZN(n4795) );
  INV_X1 U5207 ( .A(n7932), .ZN(n4799) );
  NAND2_X1 U5208 ( .A1(n8342), .A2(n8249), .ZN(n5829) );
  OR2_X1 U5209 ( .A1(n8342), .A2(n8249), .ZN(n5828) );
  OR2_X1 U5210 ( .A1(n8401), .A2(n7956), .ZN(n5819) );
  OR2_X1 U5211 ( .A1(n8403), .A2(n7745), .ZN(n5808) );
  NOR2_X1 U5212 ( .A1(n7362), .A2(n8109), .ZN(n5661) );
  AND2_X1 U5213 ( .A1(n5043), .A2(n5009), .ZN(n5019) );
  NAND3_X1 U5214 ( .A1(n4818), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4817) );
  INV_X1 U5215 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4818) );
  INV_X1 U5216 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4820) );
  AOI21_X1 U5217 ( .B1(n9255), .B2(n9256), .A(n5006), .ZN(n5005) );
  INV_X1 U5218 ( .A(n9018), .ZN(n5006) );
  NOR2_X1 U5219 ( .A1(n9021), .A2(n9132), .ZN(n9026) );
  INV_X1 U5220 ( .A(n4724), .ZN(n4719) );
  OR2_X1 U5221 ( .A1(n9545), .A2(n9555), .ZN(n6508) );
  NOR2_X1 U5222 ( .A1(n9663), .A2(n9682), .ZN(n4830) );
  INV_X1 U5223 ( .A(n4925), .ZN(n4588) );
  INV_X1 U5224 ( .A(n9474), .ZN(n4587) );
  OR2_X1 U5225 ( .A1(n9012), .A2(n9000), .ZN(n4836) );
  AND2_X1 U5226 ( .A1(n4926), .A2(n4929), .ZN(n4925) );
  AND2_X1 U5227 ( .A1(n8003), .A2(n4930), .ZN(n4929) );
  NAND2_X1 U5228 ( .A1(n4431), .A2(n7800), .ZN(n4926) );
  OR2_X1 U5229 ( .A1(n9000), .A2(n10154), .ZN(n8003) );
  NAND2_X1 U5230 ( .A1(n7090), .A2(n7106), .ZN(n6417) );
  OR2_X1 U5231 ( .A1(n9570), .A2(n9574), .ZN(n9571) );
  OR2_X1 U5232 ( .A1(n4831), .A2(n9629), .ZN(n9627) );
  NAND2_X1 U5233 ( .A1(n4725), .A2(n5728), .ZN(n4724) );
  INV_X1 U5234 ( .A(n5731), .ZN(n4725) );
  AOI21_X1 U5235 ( .B1(n4722), .B2(n5731), .A(n4495), .ZN(n4721) );
  AND2_X1 U5236 ( .A1(n5992), .A2(P1_IR_REG_30__SCAN_IN), .ZN(n4980) );
  NAND2_X1 U5237 ( .A1(n4982), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4981) );
  OAI22_X1 U5238 ( .A1(n4981), .A2(n5992), .B1(P1_IR_REG_31__SCAN_IN), .B2(
        n4982), .ZN(n4978) );
  OAI21_X1 U5239 ( .B1(n5721), .B2(n5720), .A(n5719), .ZN(n5732) );
  OR2_X1 U5240 ( .A1(n5718), .A2(n5717), .ZN(n5719) );
  INV_X1 U5241 ( .A(n5570), .ZN(n5572) );
  INV_X1 U5242 ( .A(n4710), .ZN(n4709) );
  AND2_X1 U5243 ( .A1(n5551), .A2(n5538), .ZN(n5549) );
  AOI21_X1 U5244 ( .B1(n4753), .B2(n5395), .A(n4493), .ZN(n4752) );
  AOI21_X1 U5245 ( .B1(n5354), .B2(n4690), .A(n4492), .ZN(n4689) );
  NOR2_X1 U5246 ( .A1(n5261), .A2(n4741), .ZN(n4740) );
  INV_X1 U5247 ( .A(n5241), .ZN(n4741) );
  INV_X1 U5248 ( .A(n5257), .ZN(n5261) );
  OAI21_X1 U5249 ( .B1(n5233), .B2(n5232), .A(n5231), .ZN(n5240) );
  NOR2_X1 U5250 ( .A1(n4696), .A2(n4693), .ZN(n4692) );
  INV_X1 U5251 ( .A(n5205), .ZN(n4696) );
  INV_X1 U5252 ( .A(n5188), .ZN(n4693) );
  INV_X1 U5253 ( .A(n5192), .ZN(n4695) );
  INV_X1 U5254 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5968) );
  NAND2_X1 U5255 ( .A1(n8362), .A2(n8363), .ZN(n8200) );
  CLKBUF_X1 U5256 ( .A(n7453), .Z(n8206) );
  INV_X1 U5257 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5145) );
  NAND2_X1 U5258 ( .A1(n8375), .A2(n4950), .ZN(n8302) );
  NOR2_X1 U5259 ( .A1(n8290), .A2(n4951), .ZN(n4950) );
  INV_X1 U5260 ( .A(n8167), .ZN(n4951) );
  XNOR2_X1 U5261 ( .A(n7453), .B(n7826), .ZN(n7369) );
  AND2_X1 U5262 ( .A1(n5775), .A2(n5939), .ZN(n5776) );
  OR2_X1 U5263 ( .A1(n5774), .A2(n7363), .ZN(n5775) );
  AND2_X1 U5264 ( .A1(n5067), .A2(n5066), .ZN(n4535) );
  AND2_X1 U5265 ( .A1(n5063), .A2(n5062), .ZN(n5068) );
  NAND2_X1 U5266 ( .A1(n4866), .A2(n4867), .ZN(n4873) );
  NAND2_X1 U5267 ( .A1(n4874), .A2(n4876), .ZN(n4872) );
  INV_X1 U5268 ( .A(n4875), .ZN(n4874) );
  AOI21_X1 U5269 ( .B1(n4436), .B2(n7450), .A(n7539), .ZN(n7435) );
  INV_X1 U5270 ( .A(n4848), .ZN(n4847) );
  NAND2_X1 U5271 ( .A1(n4881), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8078) );
  AND2_X1 U5272 ( .A1(n4843), .A2(n4473), .ZN(n8451) );
  NAND2_X1 U5273 ( .A1(n5679), .A2(n5678), .ZN(n7221) );
  NOR2_X1 U5274 ( .A1(n5677), .A2(n8109), .ZN(n5678) );
  INV_X1 U5275 ( .A(n8103), .ZN(n5679) );
  INV_X1 U5276 ( .A(n4611), .ZN(n8649) );
  OR2_X1 U5277 ( .A1(n4617), .A2(n4413), .ZN(n4614) );
  INV_X1 U5278 ( .A(n4613), .ZN(n4612) );
  AND2_X1 U5279 ( .A1(n5548), .A2(n5547), .ZN(n8671) );
  NAND2_X1 U5280 ( .A1(n8948), .A2(n8691), .ZN(n4627) );
  INV_X1 U5281 ( .A(n4434), .ZN(n4621) );
  AND2_X1 U5282 ( .A1(n5530), .A2(n5529), .ZN(n8680) );
  AOI21_X1 U5283 ( .B1(n4784), .B2(n4790), .A(n5895), .ZN(n4783) );
  NOR2_X1 U5284 ( .A1(n8268), .A2(n4641), .ZN(n4640) );
  AND2_X1 U5285 ( .A1(n5894), .A2(n5897), .ZN(n8703) );
  NAND2_X1 U5286 ( .A1(n5889), .A2(n4788), .ZN(n4787) );
  INV_X1 U5287 ( .A(n5886), .ZN(n4788) );
  AND2_X1 U5288 ( .A1(n5431), .A2(n5860), .ZN(n8745) );
  NAND2_X1 U5289 ( .A1(n8766), .A2(n8767), .ZN(n4647) );
  AOI21_X1 U5290 ( .B1(n4767), .B2(n4770), .A(n4766), .ZN(n4765) );
  AOI21_X1 U5291 ( .B1(n4414), .B2(n4769), .A(n4768), .ZN(n4767) );
  INV_X1 U5292 ( .A(n5856), .ZN(n4768) );
  INV_X1 U5293 ( .A(n5352), .ZN(n4769) );
  INV_X1 U5294 ( .A(n4414), .ZN(n4770) );
  NAND2_X1 U5295 ( .A1(n8824), .A2(n5352), .ZN(n4771) );
  OR2_X1 U5296 ( .A1(n5363), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5387) );
  AOI21_X1 U5297 ( .B1(n4637), .B2(n4635), .A(n4455), .ZN(n4634) );
  INV_X1 U5298 ( .A(n4637), .ZN(n4636) );
  OR2_X1 U5299 ( .A1(n8885), .A2(n8898), .ZN(n8804) );
  NAND2_X1 U5300 ( .A1(n4639), .A2(n5845), .ZN(n8815) );
  NAND2_X1 U5301 ( .A1(n5289), .A2(n5288), .ZN(n5306) );
  INV_X1 U5302 ( .A(n5290), .ZN(n5289) );
  NOR2_X1 U5303 ( .A1(n5758), .A2(n4797), .ZN(n4796) );
  INV_X1 U5304 ( .A(n5813), .ZN(n4797) );
  NAND2_X1 U5305 ( .A1(n4800), .A2(n4799), .ZN(n4798) );
  INV_X1 U5306 ( .A(n7928), .ZN(n4800) );
  NAND2_X1 U5307 ( .A1(n5828), .A2(n5829), .ZN(n8137) );
  OR2_X1 U5308 ( .A1(n8405), .A2(n7650), .ZN(n7712) );
  OR2_X1 U5309 ( .A1(n6617), .A2(n7358), .ZN(n8901) );
  INV_X1 U5310 ( .A(n8780), .ZN(n8899) );
  AND2_X1 U5311 ( .A1(n8922), .A2(n7764), .ZN(n5952) );
  NOR3_X1 U5312 ( .A1(n7292), .A2(n5708), .A3(n6615), .ZN(n5951) );
  OR2_X1 U5313 ( .A1(n5946), .A2(n5704), .ZN(n5949) );
  OR2_X1 U5314 ( .A1(n5947), .A2(n5705), .ZN(n5950) );
  AND3_X1 U5315 ( .A1(n5198), .A2(n5197), .A3(n5196), .ZN(n7902) );
  NAND2_X1 U5316 ( .A1(n7923), .A2(n7764), .ZN(n8917) );
  INV_X1 U5317 ( .A(n5661), .ZN(n6987) );
  NAND2_X1 U5318 ( .A1(n7221), .A2(n7300), .ZN(n6986) );
  NAND2_X1 U5319 ( .A1(n4959), .A2(n5033), .ZN(n4568) );
  NAND2_X1 U5320 ( .A1(n5357), .A2(n5033), .ZN(n5381) );
  NAND2_X1 U5321 ( .A1(n5357), .A2(n4566), .ZN(n5650) );
  INV_X1 U5322 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5030) );
  NOR2_X1 U5323 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n4760) );
  INV_X1 U5324 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n9967) );
  INV_X1 U5325 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4896) );
  OR2_X1 U5326 ( .A1(n9111), .A2(n4443), .ZN(n4975) );
  AOI22_X1 U5327 ( .A1(n4419), .A2(n4443), .B1(n9124), .B2(n4973), .ZN(n4972)
         );
  INV_X1 U5328 ( .A(n9111), .ZN(n4973) );
  NAND2_X1 U5329 ( .A1(n9289), .A2(n9124), .ZN(n9175) );
  AND2_X1 U5330 ( .A1(n7557), .A2(n7556), .ZN(n7669) );
  NAND2_X1 U5331 ( .A1(n6030), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6043) );
  NAND2_X1 U5332 ( .A1(n9236), .A2(n9100), .ZN(n9207) );
  NAND2_X1 U5333 ( .A1(n5980), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6176) );
  OR2_X1 U5334 ( .A1(n6176), .A2(n6165), .ZN(n6205) );
  NAND2_X1 U5335 ( .A1(n4654), .A2(n4421), .ZN(n4651) );
  NAND2_X1 U5336 ( .A1(n4421), .A2(n9276), .ZN(n4652) );
  INV_X1 U5337 ( .A(n9197), .ZN(n5007) );
  NAND2_X1 U5338 ( .A1(n5982), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6243) );
  OR2_X1 U5339 ( .A1(n6243), .A2(n10016), .ZN(n6256) );
  INV_X1 U5340 ( .A(n4963), .ZN(n4962) );
  NAND2_X1 U5341 ( .A1(n4984), .A2(n4983), .ZN(n8035) );
  NAND2_X1 U5342 ( .A1(n4986), .A2(n4989), .ZN(n4983) );
  INV_X1 U5343 ( .A(n8022), .ZN(n4989) );
  OR2_X1 U5344 ( .A1(n6205), .A2(n6920), .ZN(n6218) );
  NAND2_X1 U5345 ( .A1(n6364), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6118) );
  NOR2_X1 U5346 ( .A1(n6097), .A2(n6096), .ZN(n6101) );
  NOR2_X1 U5347 ( .A1(n6099), .A2(n6098), .ZN(n6100) );
  OR2_X1 U5348 ( .A1(n6097), .A2(n6079), .ZN(n6082) );
  AND2_X1 U5349 ( .A1(n8216), .A2(n5996), .ZN(n6095) );
  AND2_X1 U5350 ( .A1(n9391), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4684) );
  NAND2_X1 U5351 ( .A1(n6354), .A2(n6353), .ZN(n10052) );
  NAND2_X1 U5352 ( .A1(n4910), .A2(n4582), .ZN(n4581) );
  AND2_X1 U5353 ( .A1(n4908), .A2(n4917), .ZN(n4907) );
  INV_X1 U5354 ( .A(n9494), .ZN(n4582) );
  INV_X1 U5355 ( .A(n4910), .ZN(n4583) );
  AND2_X1 U5356 ( .A1(n4811), .A2(n9465), .ZN(n4810) );
  NAND2_X1 U5357 ( .A1(n9591), .A2(n4914), .ZN(n4909) );
  INV_X1 U5358 ( .A(n6019), .ZN(n5988) );
  NAND2_X1 U5359 ( .A1(n9580), .A2(n9579), .ZN(n9578) );
  NAND2_X1 U5360 ( .A1(n9606), .A2(n4453), .ZN(n9596) );
  NOR2_X1 U5361 ( .A1(n10100), .A2(n9610), .ZN(n9592) );
  NAND2_X1 U5362 ( .A1(n6329), .A2(n6569), .ZN(n9458) );
  AND2_X1 U5363 ( .A1(n6304), .A2(n6559), .ZN(n4813) );
  NAND2_X1 U5364 ( .A1(n4512), .A2(n4511), .ZN(n9716) );
  INV_X1 U5365 ( .A(n9720), .ZN(n4511) );
  NAND2_X1 U5366 ( .A1(n9478), .A2(n10244), .ZN(n9479) );
  NAND2_X1 U5367 ( .A1(n8045), .A2(n9202), .ZN(n4930) );
  NAND2_X1 U5368 ( .A1(n4924), .A2(n4923), .ZN(n7832) );
  INV_X1 U5369 ( .A(n7800), .ZN(n4923) );
  NAND2_X1 U5370 ( .A1(n4814), .A2(n6448), .ZN(n7833) );
  NOR2_X1 U5371 ( .A1(n6453), .A2(n4816), .ZN(n4815) );
  NAND2_X1 U5372 ( .A1(n7498), .A2(n6452), .ZN(n7803) );
  INV_X1 U5373 ( .A(n4905), .ZN(n4904) );
  OAI21_X1 U5374 ( .B1(n7185), .B2(n4906), .A(n7334), .ZN(n4905) );
  INV_X1 U5375 ( .A(n7328), .ZN(n4906) );
  NAND2_X1 U5376 ( .A1(n7235), .A2(n7184), .ZN(n7186) );
  NAND2_X1 U5377 ( .A1(n7186), .A2(n7185), .ZN(n7329) );
  NAND2_X1 U5378 ( .A1(n5977), .A2(n5976), .ZN(n10096) );
  NAND2_X1 U5379 ( .A1(n6016), .A2(n6015), .ZN(n10106) );
  NAND2_X1 U5380 ( .A1(n6063), .A2(n6062), .ZN(n10116) );
  NAND2_X1 U5381 ( .A1(n6295), .A2(n6294), .ZN(n9695) );
  NAND2_X1 U5382 ( .A1(n6267), .A2(n6266), .ZN(n10247) );
  INV_X1 U5383 ( .A(n10241), .ZN(n10152) );
  INV_X1 U5384 ( .A(n4515), .ZN(n4514) );
  OAI21_X1 U5385 ( .B1(n6133), .B2(n6627), .A(n6126), .ZN(n4515) );
  INV_X1 U5386 ( .A(n10125), .ZN(n10250) );
  NAND2_X1 U5387 ( .A1(n7807), .A2(n6925), .ZN(n10302) );
  NOR2_X1 U5388 ( .A1(n4992), .A2(n10213), .ZN(n4525) );
  NOR2_X1 U5389 ( .A1(n4991), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4990) );
  NAND2_X1 U5390 ( .A1(n4993), .A2(n4992), .ZN(n4991) );
  INV_X1 U5391 ( .A(n4994), .ZN(n4993) );
  NAND2_X1 U5392 ( .A1(n4708), .A2(n5516), .ZN(n5533) );
  NAND2_X1 U5393 ( .A1(n5515), .A2(n5514), .ZN(n4708) );
  AND2_X1 U5394 ( .A1(n5499), .A2(n5490), .ZN(n5497) );
  AOI21_X1 U5395 ( .B1(P1_IR_REG_17__SCAN_IN), .B2(P1_IR_REG_31__SCAN_IN), .A(
        P1_IR_REG_18__SCAN_IN), .ZN(n4665) );
  NAND2_X1 U5396 ( .A1(n4755), .A2(n5394), .ZN(n5412) );
  OR2_X1 U5397 ( .A1(n5396), .A2(n5395), .ZN(n4755) );
  NAND2_X1 U5398 ( .A1(n4732), .A2(n4736), .ZN(n5300) );
  NAND2_X1 U5399 ( .A1(n4734), .A2(n4733), .ZN(n4732) );
  NAND2_X1 U5400 ( .A1(n5178), .A2(n5177), .ZN(n5189) );
  XNOR2_X1 U5401 ( .A(n5099), .B(SI_1_), .ZN(n5098) );
  NAND2_X1 U5402 ( .A1(n6091), .A2(n5090), .ZN(n5097) );
  INV_X1 U5403 ( .A(n8783), .ZN(n8818) );
  NAND2_X1 U5404 ( .A1(n7409), .A2(n7408), .ZN(n7407) );
  XNOR2_X1 U5405 ( .A(n7369), .B(n4513), .ZN(n7409) );
  AND4_X1 U5406 ( .A1(n5447), .A2(n5446), .A3(n5445), .A4(n5444), .ZN(n8713)
         );
  NAND2_X1 U5407 ( .A1(n8375), .A2(n8167), .ZN(n8289) );
  OR2_X1 U5408 ( .A1(n7639), .A2(n7638), .ZN(n4944) );
  NAND2_X1 U5409 ( .A1(n5440), .A2(n5439), .ZN(n8729) );
  NAND2_X1 U5410 ( .A1(n4938), .A2(n4939), .ZN(n4935) );
  NAND2_X1 U5411 ( .A1(n5304), .A2(n5303), .ZN(n8892) );
  INV_X1 U5412 ( .A(n8940), .ZN(n8368) );
  AND4_X1 U5413 ( .A1(n5368), .A2(n5367), .A3(n5366), .A4(n5365), .ZN(n8801)
         );
  AOI21_X1 U5414 ( .B1(n4543), .B2(n4507), .A(n7926), .ZN(n4538) );
  NAND2_X1 U5415 ( .A1(n4543), .A2(n4544), .ZN(n4542) );
  NAND2_X1 U5416 ( .A1(n5941), .A2(n8611), .ZN(n4544) );
  XNOR2_X1 U5417 ( .A(n5036), .B(P2_IR_REG_22__SCAN_IN), .ZN(n5944) );
  NAND4_X1 U5418 ( .A1(n5256), .A2(n5255), .A3(n5254), .A4(n5253), .ZN(n8399)
         );
  NAND2_X1 U5419 ( .A1(n4882), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4880) );
  NAND2_X1 U5420 ( .A1(n4879), .A2(n4882), .ZN(n4878) );
  INV_X1 U5421 ( .A(n8079), .ZN(n4879) );
  AND2_X1 U5422 ( .A1(n5325), .A2(n5339), .ZN(n8503) );
  NAND2_X1 U5423 ( .A1(n8594), .A2(n8628), .ZN(n4675) );
  INV_X1 U5424 ( .A(n8620), .ZN(n4671) );
  AOI21_X1 U5425 ( .B1(n10332), .B2(n8605), .A(n4673), .ZN(n4672) );
  OAI21_X1 U5426 ( .B1(n10330), .B2(n8595), .A(n4674), .ZN(n4673) );
  INV_X1 U5427 ( .A(n8593), .ZN(n4674) );
  AND2_X1 U5428 ( .A1(n7210), .A2(n8622), .ZN(n10327) );
  NOR2_X1 U5429 ( .A1(n8631), .A2(n4510), .ZN(n4509) );
  OAI21_X1 U5430 ( .B1(n10330), .B2(n4821), .A(n8630), .ZN(n4510) );
  NAND2_X1 U5431 ( .A1(n5420), .A2(n5419), .ZN(n8744) );
  OR2_X1 U5432 ( .A1(n5957), .A2(n8912), .ZN(n4607) );
  NAND2_X1 U5433 ( .A1(n8647), .A2(n5701), .ZN(n5714) );
  AND2_X1 U5434 ( .A1(n5559), .A2(n5558), .ZN(n8936) );
  OR2_X1 U5435 ( .A1(n10375), .A2(n8917), .ZN(n8980) );
  XNOR2_X1 U5436 ( .A(n6587), .B(n6586), .ZN(n6639) );
  INV_X1 U5437 ( .A(n9607), .ZN(n9496) );
  INV_X1 U5438 ( .A(n10076), .ZN(n9499) );
  MUX2_X1 U5439 ( .A(n6520), .B(n6519), .S(n6790), .Z(n6521) );
  NAND2_X1 U5440 ( .A1(n6037), .A2(n6036), .ZN(n10086) );
  NAND2_X1 U5441 ( .A1(n9446), .A2(n9746), .ZN(n9761) );
  XNOR2_X1 U5442 ( .A(n4805), .B(n9505), .ZN(n10057) );
  OAI21_X1 U5443 ( .B1(n9520), .B2(n9471), .A(n9470), .ZN(n4805) );
  AND2_X1 U5444 ( .A1(n6360), .A2(n6359), .ZN(n9528) );
  AND2_X1 U5445 ( .A1(n9524), .A2(n9523), .ZN(n10063) );
  CLKBUF_X1 U5446 ( .A(n6846), .Z(n8124) );
  AND2_X1 U5447 ( .A1(n5788), .A2(n6617), .ZN(n4565) );
  OAI21_X1 U5448 ( .B1(n7377), .B2(n4564), .A(n4562), .ZN(n5805) );
  INV_X1 U5449 ( .A(n4563), .ZN(n4562) );
  NAND2_X1 U5450 ( .A1(n5780), .A2(n4565), .ZN(n4564) );
  OAI21_X1 U5451 ( .B1(n5787), .B2(n6617), .A(n7654), .ZN(n4563) );
  AOI21_X1 U5452 ( .B1(n5846), .B2(n4560), .A(n4558), .ZN(n4557) );
  AOI22_X1 U5453 ( .A1(n4550), .A2(n4551), .B1(n4552), .B2(n5900), .ZN(n4546)
         );
  INV_X1 U5454 ( .A(n4556), .ZN(n4551) );
  AOI21_X1 U5455 ( .B1(n6489), .B2(n4524), .A(n4467), .ZN(n6492) );
  AND2_X1 U5456 ( .A1(n6488), .A2(n6487), .ZN(n4524) );
  INV_X1 U5457 ( .A(n5516), .ZN(n4711) );
  NAND2_X1 U5458 ( .A1(n4645), .A2(n5616), .ZN(n5613) );
  NAND2_X1 U5459 ( .A1(n7991), .A2(n8137), .ZN(n4645) );
  OR2_X1 U5460 ( .A1(n9033), .A2(n9222), .ZN(n9035) );
  NAND2_X1 U5461 ( .A1(n10176), .A2(n10180), .ZN(n4841) );
  INV_X1 U5462 ( .A(n5725), .ZN(n4723) );
  NOR2_X1 U5463 ( .A1(n5728), .A2(n4723), .ZN(n4722) );
  OAI21_X1 U5464 ( .B1(n5573), .B2(n4701), .A(n4699), .ZN(n5718) );
  AOI21_X1 U5465 ( .B1(n4703), .B2(n4700), .A(n4498), .ZN(n4699) );
  INV_X1 U5466 ( .A(n4703), .ZN(n4701) );
  NOR2_X1 U5467 ( .A1(n4707), .A2(n4711), .ZN(n4706) );
  INV_X1 U5468 ( .A(n5499), .ZN(n4707) );
  OAI21_X1 U5469 ( .B1(n5514), .B2(n4711), .A(n5532), .ZN(n4710) );
  NOR2_X1 U5470 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5965) );
  NOR2_X1 U5471 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5966) );
  NOR2_X1 U5472 ( .A1(n5353), .A2(n5334), .ZN(n4688) );
  INV_X1 U5473 ( .A(n5338), .ZN(n4690) );
  INV_X1 U5474 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5284) );
  INV_X1 U5475 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5263) );
  AOI21_X1 U5476 ( .B1(n5748), .B2(n4457), .A(n5747), .ZN(n4772) );
  INV_X1 U5477 ( .A(n5924), .ZN(n4778) );
  OAI21_X1 U5478 ( .B1(n5636), .B2(n7279), .A(n4676), .ZN(n7194) );
  NAND2_X1 U5479 ( .A1(n4866), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4875) );
  NAND2_X1 U5480 ( .A1(n8522), .A2(n8521), .ZN(n8546) );
  AOI21_X1 U5481 ( .B1(n8586), .B2(n8597), .A(n8585), .ZN(n8587) );
  AND2_X1 U5482 ( .A1(n8952), .A2(n8392), .ZN(n5903) );
  INV_X1 U5483 ( .A(n5875), .ZN(n4766) );
  AND2_X1 U5484 ( .A1(n5625), .A2(n4638), .ZN(n4637) );
  NAND2_X1 U5485 ( .A1(n5623), .A2(n5842), .ZN(n4638) );
  INV_X1 U5486 ( .A(n5623), .ZN(n4635) );
  AND2_X1 U5487 ( .A1(n7929), .A2(n5613), .ZN(n5612) );
  NAND2_X1 U5488 ( .A1(n5222), .A2(n5221), .ZN(n5251) );
  INV_X1 U5489 ( .A(n5223), .ZN(n5222) );
  NOR2_X1 U5490 ( .A1(n6987), .A2(n5676), .ZN(n5708) );
  OAI21_X1 U5491 ( .B1(n6987), .B2(P2_D_REG_0__SCAN_IN), .A(n6989), .ZN(n5946)
         );
  NAND2_X1 U5492 ( .A1(n6992), .A2(n5660), .ZN(n5947) );
  OR2_X1 U5493 ( .A1(n5709), .A2(n5708), .ZN(n7291) );
  AND2_X1 U5494 ( .A1(n4801), .A2(n5357), .ZN(n5073) );
  NOR2_X1 U5495 ( .A1(n4803), .A2(n4802), .ZN(n4801) );
  NAND2_X1 U5496 ( .A1(n5057), .A2(n5033), .ZN(n4802) );
  NAND2_X1 U5497 ( .A1(n5681), .A2(n5680), .ZN(n5652) );
  OAI21_X2 U5498 ( .B1(n5645), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5681) );
  INV_X1 U5499 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5680) );
  INV_X1 U5500 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5045) );
  AND2_X1 U5501 ( .A1(n4438), .A2(n9020), .ZN(n5002) );
  INV_X1 U5502 ( .A(n5005), .ZN(n5001) );
  NAND2_X1 U5503 ( .A1(n5002), .A2(n4998), .ZN(n4997) );
  INV_X1 U5504 ( .A(n9198), .ZN(n4998) );
  OR2_X1 U5505 ( .A1(n9072), .A2(n9071), .ZN(n9073) );
  AND2_X1 U5506 ( .A1(n9028), .A2(n9035), .ZN(n9034) );
  INV_X1 U5507 ( .A(n10219), .ZN(n5996) );
  NAND2_X1 U5508 ( .A1(n4679), .A2(n4678), .ZN(n7474) );
  NAND2_X1 U5509 ( .A1(n7263), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4678) );
  INV_X1 U5510 ( .A(n7257), .ZN(n4679) );
  NAND2_X1 U5511 ( .A1(n4840), .A2(n4839), .ZN(n4838) );
  INV_X1 U5512 ( .A(n4841), .ZN(n4840) );
  NAND2_X1 U5513 ( .A1(n4910), .A2(n4912), .ZN(n4908) );
  INV_X1 U5514 ( .A(n4913), .ZN(n4912) );
  AOI21_X1 U5515 ( .B1(n4920), .B2(n4919), .A(n4918), .ZN(n4917) );
  NOR2_X1 U5516 ( .A1(n10180), .A2(n10066), .ZN(n4918) );
  INV_X1 U5517 ( .A(n9502), .ZN(n4919) );
  AND2_X1 U5518 ( .A1(n9501), .A2(n9500), .ZN(n4920) );
  NAND2_X1 U5519 ( .A1(n9702), .A2(n9481), .ZN(n6288) );
  AND2_X1 U5520 ( .A1(n6464), .A2(n6559), .ZN(n9481) );
  NOR2_X1 U5521 ( .A1(n4835), .A2(n10247), .ZN(n4833) );
  OR2_X1 U5522 ( .A1(n9752), .A2(n4836), .ZN(n4835) );
  OR2_X1 U5523 ( .A1(n9752), .A2(n10244), .ZN(n6550) );
  NAND2_X1 U5524 ( .A1(n6196), .A2(n6195), .ZN(n6541) );
  AND2_X1 U5525 ( .A1(n7388), .A2(n7330), .ZN(n6434) );
  AND2_X1 U5526 ( .A1(n7045), .A2(n10269), .ZN(n4825) );
  NAND2_X1 U5527 ( .A1(n7012), .A2(n6977), .ZN(n6127) );
  NAND2_X1 U5528 ( .A1(n6846), .A2(n6748), .ZN(n6533) );
  NOR2_X1 U5529 ( .A1(n9571), .A2(n9561), .ZN(n9556) );
  NOR2_X1 U5530 ( .A1(n4829), .A2(n10116), .ZN(n4828) );
  INV_X1 U5531 ( .A(n4830), .ZN(n4829) );
  AND2_X1 U5532 ( .A1(n9693), .A2(n10201), .ZN(n9694) );
  INV_X1 U5533 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6161) );
  AOI21_X1 U5534 ( .B1(n4747), .B2(n4750), .A(n4745), .ZN(n4744) );
  NOR2_X1 U5535 ( .A1(n5411), .A2(n4754), .ZN(n4753) );
  INV_X1 U5536 ( .A(n5394), .ZN(n4754) );
  INV_X1 U5537 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6252) );
  INV_X1 U5538 ( .A(n5282), .ZN(n4739) );
  INV_X1 U5539 ( .A(n5242), .ZN(n4734) );
  XNOR2_X1 U5540 ( .A(n5258), .B(SI_10_), .ZN(n5257) );
  INV_X1 U5541 ( .A(SI_9_), .ZN(n5234) );
  OR2_X1 U5542 ( .A1(n6147), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n6158) );
  OAI21_X1 U5543 ( .B1(n6624), .B2(P2_DATAO_REG_3__SCAN_IN), .A(n4698), .ZN(
        n5135) );
  OAI211_X1 U5544 ( .C1(n4819), .C2(P2_DATAO_REG_1__SCAN_IN), .A(n4633), .B(
        n4631), .ZN(n5099) );
  NAND2_X1 U5545 ( .A1(n4632), .A2(n5076), .ZN(n4631) );
  INV_X1 U5546 ( .A(n4817), .ZN(n4632) );
  OR2_X1 U5547 ( .A1(n8179), .A2(n8325), .ZN(n8261) );
  INV_X1 U5548 ( .A(n7519), .ZN(n4948) );
  INV_X1 U5549 ( .A(n8189), .ZN(n8309) );
  AND2_X1 U5550 ( .A1(n7518), .A2(n8406), .ZN(n7519) );
  NAND2_X1 U5551 ( .A1(n4946), .A2(n4947), .ZN(n7640) );
  AND2_X1 U5552 ( .A1(n7522), .A2(n4948), .ZN(n4947) );
  NAND2_X1 U5553 ( .A1(n7896), .A2(n4956), .ZN(n7951) );
  NOR2_X1 U5554 ( .A1(n7899), .A2(n4957), .ZN(n4956) );
  INV_X1 U5555 ( .A(n7895), .ZN(n4957) );
  INV_X1 U5556 ( .A(n4940), .ZN(n4939) );
  AND2_X1 U5557 ( .A1(n5021), .A2(n8271), .ZN(n4934) );
  OR2_X1 U5558 ( .A1(n4476), .A2(n4937), .ZN(n4936) );
  AND2_X1 U5559 ( .A1(n8186), .A2(n8332), .ZN(n8235) );
  NAND2_X1 U5560 ( .A1(n5455), .A2(n5454), .ZN(n5478) );
  INV_X1 U5561 ( .A(n5456), .ZN(n5455) );
  OR3_X1 U5562 ( .A1(n7293), .A2(n5930), .A3(n8908), .ZN(n7286) );
  OR2_X1 U5563 ( .A1(n7302), .A2(n7769), .ZN(n7359) );
  NAND2_X1 U5564 ( .A1(n4532), .A2(n4531), .ZN(n5933) );
  AND2_X1 U5565 ( .A1(n5932), .A2(n4483), .ZN(n4526) );
  AND2_X1 U5566 ( .A1(n7274), .A2(n7273), .ZN(n7271) );
  OR2_X1 U5567 ( .A1(n7278), .A2(n7279), .ZN(n7276) );
  NAND2_X1 U5568 ( .A1(n7276), .A2(n7213), .ZN(n10319) );
  NAND2_X1 U5569 ( .A1(n10319), .A2(n10320), .ZN(n10318) );
  NAND2_X1 U5570 ( .A1(n4852), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7423) );
  NAND2_X1 U5571 ( .A1(n4876), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7428) );
  INV_X1 U5572 ( .A(n4871), .ZN(n4868) );
  AOI21_X1 U5573 ( .B1(n4846), .B2(n4849), .A(n7450), .ZN(n4845) );
  NOR2_X1 U5574 ( .A1(n4851), .A2(n4854), .ZN(n4846) );
  NAND2_X1 U5575 ( .A1(n7542), .A2(n4853), .ZN(n4887) );
  NAND2_X1 U5576 ( .A1(n4441), .A2(n4884), .ZN(n7785) );
  NAND2_X1 U5577 ( .A1(n7792), .A2(n7790), .ZN(n4860) );
  INV_X1 U5578 ( .A(n4862), .ZN(n4861) );
  OAI21_X1 U5579 ( .B1(n7790), .B2(n7791), .A(n4865), .ZN(n4862) );
  NAND2_X1 U5580 ( .A1(n7875), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4865) );
  NAND2_X1 U5581 ( .A1(n8410), .A2(n8409), .ZN(n8431) );
  INV_X1 U5582 ( .A(n8436), .ZN(n4859) );
  NAND2_X1 U5583 ( .A1(n8463), .A2(n8464), .ZN(n8485) );
  XNOR2_X1 U5584 ( .A(n8546), .B(n8523), .ZN(n8524) );
  NOR2_X1 U5585 ( .A1(n8509), .A2(n8524), .ZN(n8549) );
  NAND2_X1 U5586 ( .A1(n8572), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4893) );
  INV_X1 U5587 ( .A(n4677), .ZN(n8622) );
  NAND2_X1 U5588 ( .A1(n8591), .A2(n8605), .ZN(n8620) );
  NAND2_X1 U5589 ( .A1(n4781), .A2(n4780), .ZN(n4779) );
  OAI21_X1 U5590 ( .B1(n5633), .B2(n4605), .A(n4604), .ZN(n4603) );
  NOR2_X1 U5591 ( .A1(n4610), .A2(n4417), .ZN(n4605) );
  NAND2_X1 U5592 ( .A1(n5633), .A2(n4609), .ZN(n4604) );
  OR2_X1 U5593 ( .A1(n5577), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5592) );
  OR2_X1 U5594 ( .A1(n5541), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5562) );
  AOI21_X1 U5595 ( .B1(n8663), .B2(n5912), .A(n5913), .ZN(n8655) );
  NAND2_X1 U5596 ( .A1(n4623), .A2(n4629), .ZN(n4622) );
  NAND2_X1 U5597 ( .A1(n4616), .A2(n4618), .ZN(n4615) );
  INV_X1 U5598 ( .A(n8674), .ZN(n4623) );
  INV_X1 U5599 ( .A(n5631), .ZN(n4619) );
  NOR2_X1 U5600 ( .A1(n4626), .A2(n4625), .ZN(n4624) );
  INV_X1 U5601 ( .A(n4627), .ZN(n4625) );
  AND2_X1 U5602 ( .A1(n5749), .A2(n5912), .ZN(n8662) );
  OAI21_X1 U5603 ( .B1(n8684), .B2(n5900), .A(n5901), .ZN(n8675) );
  NAND2_X1 U5604 ( .A1(n5508), .A2(n5507), .ZN(n5524) );
  INV_X1 U5605 ( .A(n5509), .ZN(n5508) );
  AND3_X1 U5606 ( .A1(n5482), .A2(n5481), .A3(n5480), .ZN(n8712) );
  OR2_X1 U5607 ( .A1(n8729), .A2(n8739), .ZN(n4642) );
  NAND2_X1 U5608 ( .A1(n5423), .A2(n5422), .ZN(n5441) );
  INV_X1 U5609 ( .A(n5424), .ZN(n5423) );
  NAND2_X1 U5610 ( .A1(n5386), .A2(n5385), .ZN(n5400) );
  INV_X1 U5611 ( .A(n5387), .ZN(n5386) );
  NAND2_X1 U5612 ( .A1(n5344), .A2(n5343), .ZN(n5363) );
  INV_X1 U5613 ( .A(n5345), .ZN(n5344) );
  NAND2_X1 U5614 ( .A1(n5305), .A2(n8147), .ZN(n5328) );
  OAI21_X1 U5615 ( .B1(n7928), .B2(n4794), .A(n4791), .ZN(n8046) );
  AOI21_X1 U5616 ( .B1(n4793), .B2(n4795), .A(n4792), .ZN(n4791) );
  INV_X1 U5617 ( .A(n5828), .ZN(n4792) );
  NAND2_X1 U5618 ( .A1(n5615), .A2(n4646), .ZN(n7991) );
  NAND2_X1 U5619 ( .A1(n5611), .A2(n7972), .ZN(n4646) );
  OR2_X1 U5620 ( .A1(n8399), .A2(n8251), .ZN(n5611) );
  NAND2_X1 U5621 ( .A1(n4798), .A2(n5813), .ZN(n7970) );
  OR2_X1 U5622 ( .A1(n5199), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5223) );
  INV_X1 U5623 ( .A(n7816), .ZN(n4518) );
  OR2_X1 U5624 ( .A1(n5166), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5182) );
  NAND2_X1 U5625 ( .A1(n5181), .A2(n9823), .ZN(n5199) );
  INV_X1 U5626 ( .A(n5182), .ZN(n5181) );
  INV_X1 U5627 ( .A(n7654), .ZN(n5603) );
  AND2_X1 U5628 ( .A1(n7712), .A2(n5790), .ZN(n7654) );
  NAND2_X1 U5629 ( .A1(n7649), .A2(n7654), .ZN(n7713) );
  INV_X1 U5630 ( .A(n8901), .ZN(n8782) );
  CLKBUF_X1 U5631 ( .A(n5750), .Z(n7322) );
  AND2_X1 U5632 ( .A1(n5930), .A2(n7358), .ZN(n8780) );
  NAND2_X1 U5633 ( .A1(n5475), .A2(n5474), .ZN(n8331) );
  AND3_X1 U5634 ( .A1(n5219), .A2(n5218), .A3(n5217), .ZN(n7956) );
  AND3_X1 U5635 ( .A1(n5144), .A2(n5143), .A3(n5142), .ZN(n7650) );
  OR2_X1 U5636 ( .A1(n6617), .A2(n7367), .ZN(n7769) );
  AND2_X1 U5637 ( .A1(n7286), .A2(n10343), .ZN(n7295) );
  NOR2_X1 U5638 ( .A1(n7291), .A2(n6986), .ZN(n7305) );
  INV_X1 U5639 ( .A(n8917), .ZN(n8908) );
  NAND2_X1 U5640 ( .A1(n7219), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6615) );
  NAND2_X1 U5641 ( .A1(n5652), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5663) );
  XNOR2_X1 U5642 ( .A(n5681), .B(n5680), .ZN(n7219) );
  NAND2_X1 U5643 ( .A1(n5041), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5038) );
  AND2_X1 U5644 ( .A1(n5042), .A2(n5041), .ZN(n5939) );
  AND2_X1 U5645 ( .A1(n4954), .A2(n4953), .ZN(n4952) );
  INV_X1 U5646 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n4953) );
  OR2_X1 U5647 ( .A1(n5193), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5214) );
  INV_X1 U5648 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5194) );
  INV_X1 U5649 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6583) );
  OAI21_X1 U5650 ( .B1(n9006), .B2(n4999), .A(n4996), .ZN(n9131) );
  INV_X1 U5651 ( .A(n5002), .ZN(n4999) );
  AND2_X1 U5652 ( .A1(n4997), .A2(n5000), .ZN(n4996) );
  NAND2_X1 U5653 ( .A1(n5001), .A2(n9020), .ZN(n5000) );
  NAND2_X1 U5654 ( .A1(n5005), .A2(n4440), .ZN(n4668) );
  AND2_X1 U5655 ( .A1(n9232), .A2(n9088), .ZN(n9143) );
  NAND2_X1 U5656 ( .A1(n5984), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6297) );
  INV_X1 U5657 ( .A(n6282), .ZN(n5984) );
  NAND2_X1 U5658 ( .A1(n4967), .A2(n7061), .ZN(n7100) );
  AND2_X1 U5659 ( .A1(n7056), .A2(n7055), .ZN(n4967) );
  NAND2_X1 U5660 ( .A1(n4418), .A2(n4448), .ZN(n4988) );
  INV_X1 U5661 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6165) );
  NAND2_X1 U5662 ( .A1(n5986), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6325) );
  INV_X1 U5663 ( .A(n6323), .ZN(n5986) );
  OR2_X1 U5664 ( .A1(n6325), .A2(n9249), .ZN(n6065) );
  AOI21_X1 U5665 ( .B1(n4651), .B2(n4652), .A(n4649), .ZN(n4648) );
  INV_X1 U5666 ( .A(n9247), .ZN(n4649) );
  INV_X1 U5667 ( .A(n6218), .ZN(n5981) );
  NAND2_X1 U5668 ( .A1(n5985), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6323) );
  INV_X1 U5669 ( .A(n6308), .ZN(n5985) );
  OR2_X1 U5670 ( .A1(n9045), .A2(n9044), .ZN(n9046) );
  NAND2_X1 U5671 ( .A1(n4966), .A2(n7127), .ZN(n4965) );
  INV_X1 U5672 ( .A(n7066), .ZN(n4966) );
  NAND2_X1 U5673 ( .A1(n5983), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6268) );
  NOR2_X1 U5674 ( .A1(n4728), .A2(n6400), .ZN(n4727) );
  OR2_X1 U5675 ( .A1(n6573), .A2(n6578), .ZN(n4728) );
  NAND2_X1 U5676 ( .A1(n6578), .A2(n9449), .ZN(n6519) );
  NAND2_X1 U5677 ( .A1(n6859), .A2(n6860), .ZN(n6858) );
  AND2_X1 U5678 ( .A1(n6858), .A2(n4685), .ZN(n6662) );
  NAND2_X1 U5679 ( .A1(n6861), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4685) );
  NOR2_X1 U5680 ( .A1(n6662), .A2(n6661), .ZN(n6684) );
  NOR2_X1 U5681 ( .A1(n6880), .A2(n4488), .ZN(n6883) );
  NAND2_X1 U5682 ( .A1(n6883), .A2(n6882), .ZN(n6911) );
  INV_X1 U5683 ( .A(n7474), .ZN(n7473) );
  NOR2_X1 U5684 ( .A1(n7583), .A2(n4683), .ZN(n7587) );
  AND2_X1 U5685 ( .A1(n7584), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4683) );
  NOR2_X1 U5686 ( .A1(n7587), .A2(n7586), .ZN(n7845) );
  NOR2_X1 U5687 ( .A1(n7845), .A2(n4682), .ZN(n9369) );
  AND2_X1 U5688 ( .A1(n7846), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4682) );
  OAI21_X1 U5689 ( .B1(n9410), .B2(n9409), .A(n9408), .ZN(n9412) );
  OAI21_X1 U5690 ( .B1(n4720), .B2(n6133), .A(n4714), .ZN(n9450) );
  NAND2_X1 U5691 ( .A1(n4579), .A2(n4578), .ZN(n9522) );
  AOI21_X1 U5692 ( .B1(n4423), .B2(n4583), .A(n4468), .ZN(n4578) );
  AOI21_X1 U5693 ( .B1(n4810), .B2(n4808), .A(n6333), .ZN(n4807) );
  INV_X1 U5694 ( .A(n4810), .ZN(n4809) );
  AND2_X1 U5695 ( .A1(n6341), .A2(n6032), .ZN(n9552) );
  OR2_X1 U5696 ( .A1(n6009), .A2(n9241), .ZN(n6041) );
  AND2_X1 U5697 ( .A1(n6490), .A2(n9464), .ZN(n9597) );
  AND2_X1 U5698 ( .A1(n9462), .A2(n9459), .ZN(n4806) );
  NAND2_X1 U5699 ( .A1(n9694), .A2(n4830), .ZN(n9655) );
  NAND2_X1 U5700 ( .A1(n9694), .A2(n10197), .ZN(n9679) );
  OR2_X1 U5701 ( .A1(n9682), .A2(n10119), .ZN(n9484) );
  AND2_X1 U5702 ( .A1(n6563), .A2(n6569), .ZN(n9653) );
  AND2_X1 U5703 ( .A1(n9689), .A2(n6480), .ZN(n9669) );
  NAND2_X1 U5704 ( .A1(n9669), .A2(n9671), .ZN(n9668) );
  AND2_X1 U5705 ( .A1(n6562), .A2(n6481), .ZN(n9671) );
  NAND2_X1 U5706 ( .A1(n6288), .A2(n6559), .ZN(n9687) );
  NAND2_X1 U5707 ( .A1(n9480), .A2(n10247), .ZN(n4577) );
  NAND2_X1 U5708 ( .A1(n4576), .A2(n10144), .ZN(n4575) );
  NAND2_X1 U5709 ( .A1(n4832), .A2(n4834), .ZN(n9745) );
  INV_X1 U5710 ( .A(n4835), .ZN(n4834) );
  NAND2_X1 U5711 ( .A1(n7998), .A2(n6545), .ZN(n9739) );
  AND2_X1 U5712 ( .A1(n6262), .A2(n6545), .ZN(n4812) );
  INV_X1 U5713 ( .A(n4586), .ZN(n4584) );
  INV_X1 U5714 ( .A(n4927), .ZN(n4585) );
  AOI21_X1 U5715 ( .B1(n4589), .B2(n4588), .A(n4587), .ZN(n4586) );
  NOR2_X1 U5716 ( .A1(n7837), .A2(n4836), .ZN(n9747) );
  NAND2_X1 U5717 ( .A1(n6233), .A2(n6232), .ZN(n9000) );
  NOR2_X1 U5718 ( .A1(n7837), .A2(n9000), .ZN(n8012) );
  OR2_X1 U5719 ( .A1(n7664), .A2(n9313), .ZN(n7495) );
  NAND2_X1 U5720 ( .A1(n6212), .A2(n6211), .ZN(n7498) );
  AND2_X1 U5721 ( .A1(n4442), .A2(n7177), .ZN(n7237) );
  INV_X1 U5722 ( .A(n9746), .ZN(n9723) );
  NAND2_X1 U5723 ( .A1(n7017), .A2(n10269), .ZN(n7016) );
  AOI21_X1 U5724 ( .B1(n6111), .B2(n6112), .A(n6893), .ZN(n4574) );
  INV_X1 U5725 ( .A(n6535), .ZN(n4573) );
  NAND2_X1 U5726 ( .A1(n6093), .A2(n6928), .ZN(n6933) );
  NOR2_X1 U5727 ( .A1(n4901), .A2(n6928), .ZN(n7017) );
  AND2_X1 U5728 ( .A1(n6815), .A2(n7751), .ZN(n9746) );
  NAND2_X1 U5729 ( .A1(n6372), .A2(n6371), .ZN(n6386) );
  NAND2_X1 U5730 ( .A1(n6370), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n6371) );
  NAND2_X1 U5731 ( .A1(n8154), .A2(n6376), .ZN(n6372) );
  NAND2_X1 U5732 ( .A1(n6006), .A2(n6005), .ZN(n10100) );
  INV_X1 U5733 ( .A(n10153), .ZN(n10244) );
  NAND2_X1 U5734 ( .A1(n4720), .A2(n4712), .ZN(n8982) );
  INV_X1 U5735 ( .A(n4713), .ZN(n4712) );
  INV_X1 U5736 ( .A(n4978), .ZN(n4977) );
  XNOR2_X1 U5737 ( .A(n5732), .B(n5731), .ZN(n8154) );
  INV_X1 U5738 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5992) );
  XNOR2_X1 U5739 ( .A(n5721), .B(SI_29_), .ZN(n8986) );
  XNOR2_X1 U5740 ( .A(n5587), .B(n5586), .ZN(n8113) );
  NAND2_X1 U5741 ( .A1(n4702), .A2(n5571), .ZN(n5587) );
  XNOR2_X1 U5742 ( .A(n5569), .B(n5570), .ZN(n8110) );
  NAND2_X1 U5743 ( .A1(n4743), .A2(n4747), .ZN(n5449) );
  OR2_X1 U5744 ( .A1(n5396), .A2(n4750), .ZN(n4743) );
  OAI21_X1 U5745 ( .B1(n6293), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6315) );
  NAND2_X1 U5746 ( .A1(n6293), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6305) );
  NAND2_X1 U5747 ( .A1(n4691), .A2(n5338), .ZN(n5355) );
  NAND2_X1 U5748 ( .A1(n5336), .A2(n5335), .ZN(n4691) );
  AND2_X1 U5749 ( .A1(n6230), .A2(n10014), .ZN(n6253) );
  NAND2_X1 U5750 ( .A1(n4735), .A2(n5260), .ZN(n5283) );
  AND2_X1 U5751 ( .A1(n6202), .A2(n6213), .ZN(n7026) );
  AOI21_X1 U5752 ( .B1(n4695), .B2(n5205), .A(n4465), .ZN(n4694) );
  NAND2_X1 U5753 ( .A1(n5189), .A2(n4692), .ZN(n4644) );
  INV_X1 U5754 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n6122) );
  NAND2_X1 U5755 ( .A1(n7896), .A2(n7895), .ZN(n7898) );
  NAND2_X1 U5756 ( .A1(n8200), .A2(n8199), .ZN(n8219) );
  XNOR2_X1 U5757 ( .A(n8308), .B(n8309), .ZN(n8310) );
  NAND2_X1 U5758 ( .A1(n5492), .A2(n5491), .ZN(n8240) );
  OR2_X1 U5759 ( .A1(n7454), .A2(n8407), .ZN(n7455) );
  AND2_X1 U5760 ( .A1(n5741), .A2(n5596), .ZN(n8211) );
  NAND2_X1 U5761 ( .A1(n7951), .A2(n7950), .ZN(n8061) );
  INV_X1 U5762 ( .A(n8396), .ZN(n8819) );
  NAND2_X1 U5763 ( .A1(n8343), .A2(n4940), .ZN(n8273) );
  NAND2_X1 U5764 ( .A1(n5521), .A2(n5520), .ZN(n8285) );
  NAND2_X1 U5765 ( .A1(n5384), .A2(n5383), .ZN(n8772) );
  NAND2_X1 U5766 ( .A1(n8063), .A2(n8062), .ZN(n8065) );
  NAND2_X1 U5767 ( .A1(n7951), .A2(n4955), .ZN(n8063) );
  AND2_X1 U5768 ( .A1(n4502), .A2(n7950), .ZN(n4955) );
  AND4_X1 U5769 ( .A1(n5430), .A2(n5429), .A3(n5428), .A4(n5427), .ZN(n8758)
         );
  AOI21_X1 U5770 ( .B1(n8145), .B2(n8144), .A(n8143), .ZN(n8345) );
  NOR2_X1 U5771 ( .A1(n8142), .A2(n8399), .ZN(n8143) );
  NAND2_X1 U5772 ( .A1(n8345), .A2(n5021), .ZN(n8343) );
  NAND2_X1 U5773 ( .A1(n7407), .A2(n4435), .ZN(n7371) );
  AND4_X1 U5774 ( .A1(n5392), .A2(n5391), .A3(n5390), .A4(n5389), .ZN(n8757)
         );
  NOR2_X1 U5775 ( .A1(n7740), .A2(n5010), .ZN(n7742) );
  INV_X1 U5776 ( .A(n8379), .ZN(n8355) );
  XNOR2_X1 U5777 ( .A(n8197), .B(n8671), .ZN(n8363) );
  INV_X1 U5778 ( .A(n8374), .ZN(n8163) );
  NAND2_X1 U5779 ( .A1(n7452), .A2(n7926), .ZN(n8381) );
  INV_X1 U5780 ( .A(n8712), .ZN(n8393) );
  INV_X1 U5781 ( .A(n8758), .ZN(n8725) );
  INV_X1 U5782 ( .A(n8757), .ZN(n8781) );
  NAND4_X1 U5783 ( .A1(n5132), .A2(n5131), .A3(n5130), .A4(n5129), .ZN(n8405)
         );
  NAND2_X1 U5784 ( .A1(n4850), .A2(n4849), .ZN(n7434) );
  INV_X1 U5785 ( .A(n8078), .ZN(n8075) );
  NOR2_X1 U5786 ( .A1(n8412), .A2(n5275), .ZN(n8433) );
  INV_X1 U5787 ( .A(n8936), .ZN(n8653) );
  NAND2_X1 U5788 ( .A1(n4628), .A2(n4627), .ZN(n8669) );
  NAND2_X1 U5789 ( .A1(n4630), .A2(n4620), .ZN(n4628) );
  NAND2_X1 U5790 ( .A1(n4630), .A2(n4434), .ZN(n8678) );
  NAND2_X1 U5791 ( .A1(n4786), .A2(n4787), .ZN(n8704) );
  NAND2_X1 U5792 ( .A1(n4782), .A2(n4789), .ZN(n4786) );
  NAND2_X1 U5793 ( .A1(n4782), .A2(n4415), .ZN(n8715) );
  NOR2_X1 U5794 ( .A1(n8864), .A2(n5881), .ZN(n8727) );
  NAND2_X1 U5795 ( .A1(n5399), .A2(n5398), .ZN(n8868) );
  OAI21_X1 U5796 ( .B1(n8802), .B2(n4770), .A(n4767), .ZN(n8771) );
  AND2_X1 U5797 ( .A1(n4771), .A2(n4439), .ZN(n8789) );
  NAND2_X1 U5798 ( .A1(n8815), .A2(n5623), .ZN(n8798) );
  NAND2_X1 U5799 ( .A1(n5327), .A2(n5326), .ZN(n8885) );
  AND2_X1 U5800 ( .A1(n7731), .A2(n8611), .ZN(n10231) );
  NAND2_X1 U5801 ( .A1(n5287), .A2(n5286), .ZN(n8907) );
  NAND2_X1 U5802 ( .A1(n4798), .A2(n4796), .ZN(n7987) );
  INV_X1 U5803 ( .A(n8251), .ZN(n8918) );
  OR2_X1 U5804 ( .A1(n6619), .A2(n10317), .ZN(n5106) );
  OR2_X1 U5805 ( .A1(n6986), .A2(n5953), .ZN(n10345) );
  INV_X1 U5806 ( .A(n10345), .ZN(n8822) );
  NAND2_X1 U5807 ( .A1(n5714), .A2(n8925), .ZN(n5712) );
  OR2_X1 U5808 ( .A1(n5104), .A2(n7285), .ZN(n5083) );
  OR2_X1 U5809 ( .A1(n5139), .A2(n6629), .ZN(n4761) );
  OR2_X1 U5810 ( .A1(n5117), .A2(n6631), .ZN(n4762) );
  AND3_X2 U5811 ( .A1(n5710), .A2(n5951), .A3(n5709), .ZN(n8925) );
  INV_X1 U5812 ( .A(n5745), .ZN(n8932) );
  AND2_X1 U5813 ( .A1(n5540), .A2(n5539), .ZN(n8940) );
  INV_X1 U5814 ( .A(n8240), .ZN(n8952) );
  OR2_X1 U5815 ( .A1(n8867), .A2(n8866), .ZN(n8963) );
  CLKBUF_X1 U5816 ( .A(n7366), .Z(n6989) );
  NAND2_X1 U5817 ( .A1(n6988), .A2(n6987), .ZN(n7040) );
  AND2_X1 U5818 ( .A1(n4959), .A2(n4536), .ZN(n4958) );
  NOR2_X1 U5819 ( .A1(n4803), .A2(n4568), .ZN(n4567) );
  NOR2_X1 U5820 ( .A1(n4677), .A2(P2_U3151), .ZN(n8111) );
  NAND2_X1 U5821 ( .A1(n5650), .A2(n5649), .ZN(n8109) );
  XNOR2_X1 U5822 ( .A(n5647), .B(n5646), .ZN(n8103) );
  NAND2_X1 U5823 ( .A1(n5665), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5647) );
  INV_X1 U5824 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n9786) );
  INV_X1 U5825 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n9991) );
  INV_X1 U5826 ( .A(n5944), .ZN(n7923) );
  INV_X1 U5827 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n9990) );
  INV_X1 U5828 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7763) );
  INV_X1 U5829 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n9989) );
  INV_X1 U5830 ( .A(n5939), .ZN(n7731) );
  INV_X1 U5831 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7532) );
  INV_X1 U5832 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7357) );
  INV_X1 U5833 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7231) );
  AND2_X1 U5834 ( .A1(n4954), .A2(n4932), .ZN(n4757) );
  INV_X1 U5835 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9978) );
  AND2_X1 U5836 ( .A1(P2_U3151), .A2(n5553), .ZN(n8991) );
  INV_X1 U5837 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6783) );
  INV_X1 U5838 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6682) );
  INV_X1 U5839 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9977) );
  INV_X1 U5840 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6644) );
  XNOR2_X1 U5841 ( .A(n5172), .B(n9967), .ZN(n7687) );
  INV_X1 U5842 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5028) );
  NOR2_X1 U5843 ( .A1(n4419), .A2(n4970), .ZN(n4969) );
  INV_X1 U5844 ( .A(n4972), .ZN(n4970) );
  NAND2_X1 U5845 ( .A1(n4972), .A2(n4974), .ZN(n4971) );
  INV_X1 U5846 ( .A(n9124), .ZN(n4974) );
  AND2_X1 U5847 ( .A1(n4987), .A2(n4985), .ZN(n8021) );
  NAND2_X1 U5848 ( .A1(n9224), .A2(n4656), .ZN(n4653) );
  NAND2_X1 U5849 ( .A1(n6321), .A2(n6320), .ZN(n9663) );
  INV_X1 U5850 ( .A(n9318), .ZN(n7090) );
  NAND2_X1 U5851 ( .A1(n7100), .A2(n7066), .ZN(n7128) );
  NAND2_X1 U5852 ( .A1(n4987), .A2(n4988), .ZN(n8017) );
  OAI21_X1 U5853 ( .B1(n5008), .B2(n9256), .A(n5003), .ZN(n9254) );
  INV_X1 U5854 ( .A(n5004), .ZN(n5003) );
  OAI21_X1 U5855 ( .B1(n5007), .B2(n9256), .A(n9255), .ZN(n5004) );
  AND2_X1 U5856 ( .A1(n9079), .A2(n9142), .ZN(n9266) );
  INV_X1 U5857 ( .A(n9312), .ZN(n8040) );
  INV_X1 U5858 ( .A(n7020), .ZN(n10269) );
  AND2_X1 U5859 ( .A1(n4667), .A2(n4428), .ZN(n7150) );
  AND2_X1 U5860 ( .A1(n9111), .A2(n4659), .ZN(n4658) );
  AND2_X1 U5861 ( .A1(n6849), .A2(n6747), .ZN(n9300) );
  OR2_X1 U5862 ( .A1(n6955), .A2(n7915), .ZN(n9307) );
  NAND2_X1 U5863 ( .A1(n6049), .A2(n6048), .ZN(n10076) );
  NAND2_X1 U5864 ( .A1(n6014), .A2(n6013), .ZN(n9607) );
  OR2_X1 U5865 ( .A1(n9148), .A2(n6355), .ZN(n6014) );
  NAND2_X1 U5866 ( .A1(n6025), .A2(n6024), .ZN(n9624) );
  OR2_X1 U5867 ( .A1(n9269), .A2(n6355), .ZN(n6025) );
  NAND2_X1 U5868 ( .A1(n6061), .A2(n6060), .ZN(n9641) );
  NAND4_X1 U5869 ( .A1(n6180), .A2(n6179), .A3(n6178), .A4(n6177), .ZN(n9314)
         );
  NAND4_X2 U5870 ( .A1(n6119), .A2(n6118), .A3(n6117), .A4(n6116), .ZN(n9319)
         );
  NAND2_X1 U5871 ( .A1(n9330), .A2(n9331), .ZN(n9329) );
  NOR2_X1 U5872 ( .A1(n6765), .A2(n4681), .ZN(n6770) );
  AND2_X1 U5873 ( .A1(n6766), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4681) );
  NOR2_X1 U5874 ( .A1(n6770), .A2(n6769), .ZN(n6880) );
  NOR2_X1 U5875 ( .A1(n7025), .A2(n4680), .ZN(n7029) );
  AND2_X1 U5876 ( .A1(n7026), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4680) );
  NOR2_X1 U5877 ( .A1(n7029), .A2(n7028), .ZN(n7257) );
  XNOR2_X1 U5878 ( .A(n9369), .B(n9368), .ZN(n7847) );
  OR2_X1 U5879 ( .A1(n6664), .A2(n6935), .ZN(n9431) );
  INV_X1 U5880 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9444) );
  NAND2_X1 U5881 ( .A1(n4580), .A2(n4420), .ZN(n9539) );
  OR2_X1 U5882 ( .A1(n9495), .A2(n4583), .ZN(n4580) );
  OAI21_X1 U5883 ( .B1(n9565), .B2(n9501), .A(n9500), .ZN(n9550) );
  NAND2_X1 U5884 ( .A1(n9578), .A2(n9465), .ZN(n9564) );
  INV_X1 U5885 ( .A(n10086), .ZN(n10066) );
  NAND2_X1 U5886 ( .A1(n6039), .A2(n6038), .ZN(n9574) );
  NAND2_X1 U5887 ( .A1(n4916), .A2(n9497), .ZN(n9577) );
  OR2_X1 U5888 ( .A1(n9591), .A2(n9498), .ZN(n4916) );
  INV_X1 U5889 ( .A(n10100), .ZN(n9595) );
  NAND2_X1 U5891 ( .A1(n6280), .A2(n6279), .ZN(n9713) );
  INV_X1 U5892 ( .A(n9690), .ZN(n10242) );
  OAI21_X1 U5893 ( .B1(n7832), .B2(n4928), .A(n4431), .ZN(n8004) );
  INV_X1 U5894 ( .A(n4930), .ZN(n4928) );
  AND2_X1 U5895 ( .A1(n9757), .A2(n7004), .ZN(n9751) );
  OAI21_X1 U5896 ( .B1(n7186), .B2(n4906), .A(n4904), .ZN(n7399) );
  NAND2_X1 U5897 ( .A1(n7329), .A2(n7328), .ZN(n7331) );
  INV_X1 U5898 ( .A(n9673), .ZN(n9748) );
  INV_X1 U5899 ( .A(n9755), .ZN(n9733) );
  OR2_X1 U5900 ( .A1(n6795), .A2(n6798), .ZN(n9673) );
  AND2_X1 U5901 ( .A1(n7919), .A2(n7767), .ZN(n6815) );
  INV_X1 U5902 ( .A(n10316), .ZN(n10313) );
  INV_X1 U5903 ( .A(n6386), .ZN(n10168) );
  NAND2_X1 U5904 ( .A1(n4593), .A2(n4592), .ZN(n10169) );
  AOI21_X1 U5905 ( .B1(n10057), .B2(n10125), .A(n4472), .ZN(n4592) );
  NAND2_X1 U5906 ( .A1(n10051), .A2(n10302), .ZN(n4593) );
  AOI21_X1 U5907 ( .B1(n10063), .B2(n10302), .A(n10062), .ZN(n10170) );
  INV_X1 U5908 ( .A(n9574), .ZN(n10184) );
  INV_X1 U5909 ( .A(n9695), .ZN(n10201) );
  INV_X1 U5910 ( .A(n7089), .ZN(n7177) );
  AND2_X2 U5911 ( .A1(n6943), .A2(n6942), .ZN(n10306) );
  NAND2_X1 U5912 ( .A1(n4572), .A2(n4571), .ZN(n5974) );
  NAND2_X1 U5913 ( .A1(n5972), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4571) );
  NOR2_X1 U5914 ( .A1(n5975), .A2(n4899), .ZN(n4898) );
  NAND2_X1 U5915 ( .A1(n6594), .A2(n4525), .ZN(n4900) );
  NOR2_X1 U5916 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4899) );
  INV_X1 U5917 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7752) );
  INV_X1 U5918 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6317) );
  NAND2_X1 U5919 ( .A1(n6316), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6318) );
  INV_X1 U5920 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n9845) );
  INV_X1 U5921 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7230) );
  INV_X1 U5922 ( .A(n9362), .ZN(n9368) );
  INV_X1 U5923 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6804) );
  INV_X1 U5924 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6785) );
  INV_X1 U5925 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6653) );
  NAND2_X1 U5926 ( .A1(n4697), .A2(n5192), .ZN(n5206) );
  NAND2_X1 U5927 ( .A1(n5189), .A2(n5188), .ZN(n4697) );
  INV_X1 U5928 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6646) );
  NAND2_X1 U5929 ( .A1(n10226), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4686) );
  CLKBUF_X1 U5930 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n10226) );
  NAND2_X1 U5931 ( .A1(n4542), .A2(n5942), .ZN(n4541) );
  NAND2_X1 U5932 ( .A1(n4877), .A2(n4878), .ZN(n8423) );
  INV_X1 U5933 ( .A(n4894), .ZN(n8559) );
  NOR2_X1 U5934 ( .A1(n8604), .A2(n4669), .ZN(n8606) );
  AOI21_X1 U5935 ( .B1(n8632), .B2(n10327), .A(n4508), .ZN(n8633) );
  NAND2_X1 U5936 ( .A1(n8629), .A2(n4509), .ZN(n4508) );
  AOI21_X1 U5937 ( .B1(n5688), .B2(n8795), .A(n5956), .ZN(n5958) );
  MUX2_X1 U5938 ( .A(n9925), .B(n8933), .S(n8925), .Z(n8834) );
  NOR2_X1 U5939 ( .A1(n5689), .A2(n5691), .ZN(n5692) );
  OAI21_X1 U5940 ( .B1(n5714), .B2(n10375), .A(n5713), .ZN(n5715) );
  MUX2_X1 U5941 ( .A(n8934), .B(n8933), .S(n10372), .Z(n8935) );
  NAND2_X1 U5942 ( .A1(n4961), .A2(n6903), .ZN(n6844) );
  MUX2_X1 U5943 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n10164), .S(n10316), .Z(
        n10046) );
  AND2_X1 U5944 ( .A1(n4736), .A2(n5297), .ZN(n4411) );
  AND2_X1 U5945 ( .A1(n4760), .A2(n5080), .ZN(n4412) );
  AND2_X1 U5946 ( .A1(n8940), .A2(n8671), .ZN(n4413) );
  AND2_X1 U5947 ( .A1(n5370), .A2(n4439), .ZN(n4414) );
  AND2_X1 U5948 ( .A1(n5064), .A2(n5065), .ZN(n5250) );
  AND2_X1 U5949 ( .A1(n5431), .A2(n5887), .ZN(n4415) );
  AND4_X1 U5950 ( .A1(n4932), .A2(n7201), .A3(n5029), .A4(n4475), .ZN(n4416)
         );
  OR2_X1 U5951 ( .A1(n8213), .A2(n8387), .ZN(n4417) );
  NAND2_X1 U5952 ( .A1(n7444), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4855) );
  AND2_X1 U5953 ( .A1(n4975), .A2(n9123), .ZN(n4419) );
  AND2_X1 U5954 ( .A1(n4907), .A2(n4581), .ZN(n4420) );
  NAND2_X1 U5955 ( .A1(n9059), .A2(n9155), .ZN(n4421) );
  OR2_X1 U5956 ( .A1(n4864), .A2(n8085), .ZN(n4422) );
  AND2_X1 U5957 ( .A1(n4420), .A2(n9536), .ZN(n4423) );
  AND2_X1 U5958 ( .A1(n4615), .A2(n4622), .ZN(n4424) );
  NOR2_X1 U5959 ( .A1(n4621), .A2(n4460), .ZN(n4620) );
  INV_X1 U5960 ( .A(n4620), .ZN(n4618) );
  AND2_X1 U5961 ( .A1(n6468), .A2(n6790), .ZN(n4426) );
  OR2_X1 U5962 ( .A1(n5907), .A2(n5930), .ZN(n4427) );
  NAND2_X1 U5963 ( .A1(n4650), .A2(n4648), .ZN(n9246) );
  AND2_X1 U5964 ( .A1(n4469), .A2(n4965), .ZN(n4428) );
  AND3_X1 U5965 ( .A1(n5513), .A2(n5512), .A3(n5511), .ZN(n8691) );
  INV_X1 U5966 ( .A(n5353), .ZN(n5354) );
  AND2_X1 U5967 ( .A1(n9465), .A2(n6494), .ZN(n9579) );
  INV_X1 U5968 ( .A(n9579), .ZN(n4808) );
  AND2_X1 U5969 ( .A1(n4603), .A2(n4450), .ZN(n4429) );
  NAND2_X1 U5970 ( .A1(n5453), .A2(n5452), .ZN(n8268) );
  INV_X1 U5971 ( .A(n4738), .ZN(n4733) );
  NAND2_X1 U5972 ( .A1(n4739), .A2(n5260), .ZN(n4738) );
  INV_X1 U5973 ( .A(n7578), .ZN(n4826) );
  INV_X1 U5974 ( .A(n4790), .ZN(n4789) );
  NAND2_X1 U5975 ( .A1(n5889), .A2(n4415), .ZN(n4790) );
  NAND2_X1 U5976 ( .A1(n6073), .A2(n6072), .ZN(n9545) );
  INV_X1 U5977 ( .A(n9545), .ZN(n10176) );
  AND2_X1 U5978 ( .A1(n4878), .A2(n4491), .ZN(n4430) );
  INV_X1 U5979 ( .A(n8651), .ZN(n4780) );
  INV_X1 U5980 ( .A(n4946), .ZN(n7520) );
  OR2_X1 U5981 ( .A1(n8045), .A2(n9202), .ZN(n4431) );
  NAND2_X1 U5982 ( .A1(n5080), .A2(n4896), .ZN(n5105) );
  NAND2_X1 U5983 ( .A1(n4962), .A2(n9142), .ZN(n9141) );
  OR2_X1 U5984 ( .A1(n6595), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n4432) );
  INV_X1 U5985 ( .A(n4610), .ZN(n4609) );
  OR2_X1 U5986 ( .A1(n8082), .A2(n8081), .ZN(n4433) );
  OR2_X1 U5987 ( .A1(n8702), .A2(n8952), .ZN(n4434) );
  NAND2_X1 U5988 ( .A1(n6216), .A2(n6215), .ZN(n8028) );
  OR2_X1 U5989 ( .A1(n7369), .A2(n7304), .ZN(n4435) );
  AND2_X1 U5990 ( .A1(n6457), .A2(n6545), .ZN(n8007) );
  INV_X1 U5991 ( .A(n7684), .ZN(n4886) );
  INV_X1 U5992 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5033) );
  INV_X1 U5993 ( .A(n7791), .ZN(n4863) );
  AND2_X1 U5994 ( .A1(n4850), .A2(n4847), .ZN(n4436) );
  OR2_X1 U5995 ( .A1(n8268), .A2(n8701), .ZN(n5889) );
  INV_X1 U5996 ( .A(n4763), .ZN(n7826) );
  OR2_X1 U5997 ( .A1(n8597), .A2(n8596), .ZN(n4437) );
  AND2_X1 U5998 ( .A1(n9255), .A2(n5007), .ZN(n4438) );
  OR2_X1 U5999 ( .A1(n5351), .A2(n8804), .ZN(n4439) );
  NAND2_X1 U6000 ( .A1(n4653), .A2(n9276), .ZN(n9154) );
  XOR2_X1 U6001 ( .A(n9019), .B(n4410), .Z(n4440) );
  OR2_X1 U6002 ( .A1(n4888), .A2(n4886), .ZN(n4441) );
  INV_X1 U6003 ( .A(n6452), .ZN(n4816) );
  NAND2_X1 U6004 ( .A1(n6029), .A2(n6028), .ZN(n9561) );
  INV_X1 U6005 ( .A(n9561), .ZN(n10180) );
  INV_X1 U6006 ( .A(n7815), .ZN(n4517) );
  AND2_X1 U6007 ( .A1(n6403), .A2(n6575), .ZN(n9505) );
  AND3_X1 U6008 ( .A1(n4825), .A2(n10275), .A3(n7017), .ZN(n4442) );
  AND2_X1 U6009 ( .A1(n9122), .A2(n9121), .ZN(n4443) );
  AND2_X1 U6010 ( .A1(n4416), .A2(n5229), .ZN(n5243) );
  AND4_X1 U6011 ( .A1(n6289), .A2(n5966), .A3(n5965), .A4(n6252), .ZN(n4444)
         );
  NAND2_X1 U6012 ( .A1(n4932), .A2(n5080), .ZN(n5140) );
  NAND2_X1 U6013 ( .A1(n9187), .A2(n9188), .ZN(n9186) );
  INV_X1 U6014 ( .A(n7427), .ZN(n4866) );
  AND3_X1 U6015 ( .A1(n4597), .A2(n4608), .A3(n4599), .ZN(n4445) );
  NAND2_X1 U6016 ( .A1(n6204), .A2(n6203), .ZN(n8134) );
  OR2_X1 U6017 ( .A1(n9571), .A2(n4838), .ZN(n4446) );
  OR2_X1 U6018 ( .A1(n9571), .A2(n4841), .ZN(n4447) );
  AND2_X1 U6019 ( .A1(n7668), .A2(n7669), .ZN(n4448) );
  INV_X1 U6020 ( .A(n4617), .ZN(n4616) );
  OAI21_X1 U6021 ( .B1(n4619), .B2(n4618), .A(n4624), .ZN(n4617) );
  OR2_X1 U6022 ( .A1(n10096), .A2(n10085), .ZN(n4449) );
  NOR2_X1 U6023 ( .A1(n8007), .A2(n4590), .ZN(n4589) );
  OR2_X1 U6024 ( .A1(n5633), .A2(n4610), .ZN(n4450) );
  INV_X1 U6025 ( .A(n9629), .ZN(n10191) );
  NAND2_X1 U6026 ( .A1(n6054), .A2(n6053), .ZN(n9629) );
  AND2_X1 U6027 ( .A1(n7687), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4451) );
  INV_X1 U6028 ( .A(n9276), .ZN(n4655) );
  NOR2_X1 U6029 ( .A1(n8187), .A2(n8235), .ZN(n4452) );
  INV_X1 U6030 ( .A(n9682), .ZN(n10197) );
  NAND2_X1 U6031 ( .A1(n6307), .A2(n6306), .ZN(n9682) );
  AND2_X1 U6032 ( .A1(n9597), .A2(n9463), .ZN(n4453) );
  XNOR2_X1 U6033 ( .A(n5298), .B(SI_12_), .ZN(n5297) );
  AND2_X1 U6034 ( .A1(n10096), .A2(n10085), .ZN(n4454) );
  AND2_X1 U6035 ( .A1(n8371), .A2(n8783), .ZN(n4455) );
  AND2_X1 U6036 ( .A1(n6508), .A2(n9468), .ZN(n9538) );
  AND2_X1 U6037 ( .A1(n5845), .A2(n5844), .ZN(n4456) );
  OR2_X1 U6038 ( .A1(n4778), .A2(n4776), .ZN(n4457) );
  NAND2_X1 U6039 ( .A1(n8019), .A2(n8018), .ZN(n4458) );
  AND2_X1 U6040 ( .A1(n9578), .A2(n4810), .ZN(n4459) );
  INV_X1 U6041 ( .A(n4915), .ZN(n4914) );
  NAND2_X1 U6042 ( .A1(n4449), .A2(n9497), .ZN(n4915) );
  NOR2_X1 U6043 ( .A1(n8948), .A2(n8691), .ZN(n4460) );
  INV_X1 U6044 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4992) );
  OR2_X1 U6045 ( .A1(n8331), .A2(n8712), .ZN(n5894) );
  INV_X1 U6046 ( .A(n4629), .ZN(n4626) );
  NAND2_X1 U6047 ( .A1(n8944), .A2(n8680), .ZN(n4629) );
  NAND2_X1 U6048 ( .A1(n5576), .A2(n5575), .ZN(n8213) );
  INV_X1 U6049 ( .A(n8213), .ZN(n4781) );
  NAND2_X1 U6050 ( .A1(n7444), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4461) );
  NOR2_X1 U6051 ( .A1(n5931), .A2(n5930), .ZN(n4462) );
  INV_X1 U6052 ( .A(n4794), .ZN(n4793) );
  OAI21_X1 U6053 ( .B1(n4799), .B2(n4795), .A(n5280), .ZN(n4794) );
  OR2_X1 U6054 ( .A1(n5381), .A2(n5055), .ZN(n4463) );
  INV_X1 U6055 ( .A(n4855), .ZN(n4854) );
  INV_X1 U6056 ( .A(n6893), .ZN(n6976) );
  AND2_X1 U6057 ( .A1(n5299), .A2(SI_12_), .ZN(n4464) );
  AND2_X1 U6058 ( .A1(n5208), .A2(SI_7_), .ZN(n4465) );
  NAND2_X1 U6059 ( .A1(n8389), .A2(n8368), .ZN(n4466) );
  OR2_X1 U6060 ( .A1(n6408), .A2(n9461), .ZN(n4467) );
  INV_X1 U6061 ( .A(n7534), .ZN(n7450) );
  INV_X1 U6062 ( .A(n4785), .ZN(n4784) );
  NAND2_X1 U6063 ( .A1(n5897), .A2(n4787), .ZN(n4785) );
  INV_X1 U6064 ( .A(n8948), .ZN(n8317) );
  AND2_X1 U6065 ( .A1(n5506), .A2(n5505), .ZN(n8948) );
  AND2_X1 U6066 ( .A1(n9555), .A2(n10176), .ZN(n4468) );
  OR2_X1 U6067 ( .A1(n8744), .A2(n8758), .ZN(n5431) );
  NAND2_X1 U6068 ( .A1(n7126), .A2(n7125), .ZN(n4469) );
  NAND2_X1 U6069 ( .A1(n5898), .A2(n5905), .ZN(n4470) );
  NAND2_X1 U6070 ( .A1(n6522), .A2(n4727), .ZN(n4471) );
  OAI21_X1 U6071 ( .B1(n4656), .B2(n4655), .A(n9060), .ZN(n4654) );
  INV_X1 U6072 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6314) );
  OR2_X1 U6073 ( .A1(n10056), .A2(n10055), .ZN(n4472) );
  INV_X1 U6074 ( .A(n4986), .ZN(n4985) );
  NAND2_X1 U6075 ( .A1(n4988), .A2(n4458), .ZN(n4986) );
  OR2_X1 U6076 ( .A1(n8448), .A2(n8447), .ZN(n4473) );
  AND2_X1 U6077 ( .A1(n5057), .A2(n5069), .ZN(n4959) );
  INV_X1 U6078 ( .A(n8271), .ZN(n4937) );
  AND2_X1 U6079 ( .A1(n9474), .A2(n10153), .ZN(n4474) );
  NAND2_X1 U6080 ( .A1(n6125), .A2(n4514), .ZN(n6977) );
  INV_X1 U6081 ( .A(n6977), .ZN(n7045) );
  NAND2_X1 U6082 ( .A1(n6255), .A2(n6254), .ZN(n9752) );
  AND3_X1 U6083 ( .A1(n9976), .A2(n5194), .A3(n5153), .ZN(n4475) );
  INV_X1 U6084 ( .A(n9012), .ZN(n10210) );
  NAND2_X1 U6085 ( .A1(n6242), .A2(n6241), .ZN(n9012) );
  AND2_X1 U6086 ( .A1(n4940), .A2(n8900), .ZN(n4476) );
  OR2_X1 U6087 ( .A1(n4938), .A2(n4934), .ZN(n4477) );
  AND2_X1 U6088 ( .A1(n7127), .A2(n7055), .ZN(n4478) );
  AND2_X1 U6089 ( .A1(n6893), .A2(n6112), .ZN(n4479) );
  AND2_X1 U6090 ( .A1(n9460), .A2(n9459), .ZN(n4480) );
  AND2_X1 U6091 ( .A1(n9606), .A2(n9463), .ZN(n4481) );
  AND2_X1 U6092 ( .A1(n8203), .A2(n8199), .ZN(n4482) );
  AND2_X1 U6093 ( .A1(n4462), .A2(n4528), .ZN(n4483) );
  AND2_X1 U6094 ( .A1(n4936), .A2(n4935), .ZN(n4484) );
  OR2_X1 U6095 ( .A1(n7541), .A2(n4886), .ZN(n4485) );
  INV_X1 U6096 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4536) );
  INV_X1 U6097 ( .A(n6505), .ZN(n6790) );
  AND2_X1 U6098 ( .A1(n5008), .A2(n5007), .ZN(n4486) );
  NAND2_X1 U6099 ( .A1(n6338), .A2(n6337), .ZN(n9532) );
  INV_X1 U6100 ( .A(n9532), .ZN(n4839) );
  NAND2_X1 U6101 ( .A1(n4416), .A2(n4954), .ZN(n5245) );
  NAND2_X1 U6102 ( .A1(n4416), .A2(n4952), .ZN(n4487) );
  AND2_X1 U6103 ( .A1(n6881), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4488) );
  NAND2_X1 U6104 ( .A1(n4522), .A2(n9479), .ZN(n9719) );
  NAND2_X1 U6105 ( .A1(n4647), .A2(n5628), .ZN(n8754) );
  NAND2_X1 U6106 ( .A1(n9224), .A2(n9046), .ZN(n9274) );
  NAND2_X1 U6107 ( .A1(n5591), .A2(n5590), .ZN(n5688) );
  NOR2_X1 U6108 ( .A1(n10191), .A2(n9491), .ZN(n4489) );
  NAND2_X1 U6109 ( .A1(n4591), .A2(n5018), .ZN(n8005) );
  OR2_X1 U6110 ( .A1(n5247), .A2(n5246), .ZN(n8424) );
  AND4_X1 U6111 ( .A1(n5279), .A2(n5278), .A3(n5277), .A4(n5276), .ZN(n8249)
         );
  AND4_X1 U6112 ( .A1(n5463), .A2(n5462), .A3(n5461), .A4(n5460), .ZN(n8701)
         );
  INV_X1 U6113 ( .A(n8701), .ZN(n4641) );
  AND2_X1 U6114 ( .A1(n4771), .A2(n4414), .ZN(n4490) );
  OR2_X1 U6115 ( .A1(n8414), .A2(n8076), .ZN(n4491) );
  AND2_X1 U6116 ( .A1(n5356), .A2(SI_15_), .ZN(n4492) );
  INV_X1 U6117 ( .A(n8397), .ZN(n8900) );
  AND2_X1 U6118 ( .A1(n5410), .A2(SI_18_), .ZN(n4493) );
  NOR2_X1 U6119 ( .A1(n4489), .A2(n4931), .ZN(n4494) );
  NAND2_X1 U6120 ( .A1(n7566), .A2(n7565), .ZN(n7673) );
  NAND2_X1 U6121 ( .A1(n4518), .A2(n4517), .ZN(n7814) );
  AND2_X1 U6122 ( .A1(n5728), .A2(n4723), .ZN(n4495) );
  NOR2_X1 U6123 ( .A1(n8434), .A2(n8433), .ZN(n4496) );
  AND2_X1 U6124 ( .A1(n7497), .A2(n7501), .ZN(n7801) );
  INV_X1 U6125 ( .A(n7801), .ZN(n4924) );
  NOR2_X1 U6126 ( .A1(n7236), .A2(n7326), .ZN(n4827) );
  NAND2_X1 U6127 ( .A1(n4860), .A2(n4863), .ZN(n4497) );
  AND2_X1 U6128 ( .A1(n5589), .A2(n5588), .ZN(n4498) );
  AND2_X1 U6129 ( .A1(n6377), .A2(n4716), .ZN(n4499) );
  INV_X1 U6130 ( .A(n7208), .ZN(n4852) );
  INV_X1 U6131 ( .A(n8611), .ZN(n8617) );
  OR2_X1 U6132 ( .A1(n7421), .A2(n7422), .ZN(n4849) );
  AND2_X1 U6133 ( .A1(n8572), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4500) );
  AND2_X1 U6134 ( .A1(n4825), .A2(n7017), .ZN(n4501) );
  INV_X1 U6135 ( .A(n7217), .ZN(n4876) );
  OR2_X2 U6136 ( .A1(n7221), .A2(n6615), .ZN(n8592) );
  NAND2_X1 U6137 ( .A1(n5635), .A2(n5634), .ZN(n8785) );
  INV_X1 U6138 ( .A(n8785), .ZN(n8896) );
  OR2_X1 U6139 ( .A1(n7952), .A2(n8401), .ZN(n4502) );
  INV_X1 U6140 ( .A(n7304), .ZN(n4513) );
  AND2_X1 U6141 ( .A1(n4872), .A2(n4873), .ZN(n4503) );
  OR2_X1 U6142 ( .A1(n8617), .A2(n7731), .ZN(n4504) );
  AND2_X1 U6143 ( .A1(n4889), .A2(n4887), .ZN(n4505) );
  OR2_X1 U6144 ( .A1(n4500), .A2(n8561), .ZN(n4506) );
  XNOR2_X1 U6145 ( .A(n5047), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8611) );
  INV_X1 U6146 ( .A(n6603), .ZN(n7002) );
  NAND2_X1 U6147 ( .A1(n8617), .A2(n7731), .ZN(n4507) );
  NAND2_X1 U6148 ( .A1(n5991), .A2(n5992), .ZN(n5990) );
  INV_X1 U6149 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4821) );
  AOI21_X1 U6150 ( .B1(n7445), .B2(n7444), .A(n7443), .ZN(n7446) );
  AOI21_X1 U6151 ( .B1(n7195), .B2(n10317), .A(n10322), .ZN(n7197) );
  AOI21_X1 U6152 ( .B1(n7535), .B2(n7534), .A(n7533), .ZN(n7537) );
  OAI22_X1 U6153 ( .A1(n7871), .A2(n7870), .B1(n7869), .B2(n7875), .ZN(n7873)
         );
  AND2_X2 U6154 ( .A1(n6931), .A2(n6094), .ZN(n7010) );
  INV_X1 U6155 ( .A(n9718), .ZN(n4512) );
  NAND4_X2 U6156 ( .A1(n6085), .A2(n6086), .A3(n6088), .A4(n6087), .ZN(n9321)
         );
  AND3_X2 U6157 ( .A1(n4758), .A2(n4412), .A3(n4425), .ZN(n5321) );
  OAI21_X2 U6158 ( .B1(n6409), .B2(n6974), .A(n6127), .ZN(n6994) );
  NAND2_X1 U6159 ( .A1(n4943), .A2(n4942), .ZN(n4946) );
  NAND2_X1 U6160 ( .A1(n7456), .A2(n7455), .ZN(n7457) );
  AOI21_X1 U6161 ( .B1(n8255), .B2(n8176), .A(n5016), .ZN(n8262) );
  NOR2_X1 U6162 ( .A1(n8467), .A2(n8903), .ZN(n8477) );
  XNOR2_X1 U6163 ( .A(n8476), .B(n8493), .ZN(n8467) );
  NOR2_X1 U6164 ( .A1(n8560), .A2(n8875), .ZN(n8580) );
  NOR2_X1 U6166 ( .A1(n8508), .A2(n8883), .ZN(n8532) );
  XNOR2_X1 U6167 ( .A(n8530), .B(n8523), .ZN(n8508) );
  NOR2_X1 U6168 ( .A1(n7685), .A2(n7823), .ZN(n7783) );
  NAND3_X1 U6169 ( .A1(n4884), .A2(n4441), .A3(n4885), .ZN(n7685) );
  NAND3_X1 U6170 ( .A1(n4762), .A2(n4761), .A3(n5083), .ZN(n4763) );
  OAI211_X1 U6171 ( .C1(n4541), .C2(n5940), .A(n4516), .B(n5945), .ZN(P2_U3296) );
  NAND2_X1 U6172 ( .A1(n4538), .A2(n5940), .ZN(n4516) );
  NAND2_X1 U6173 ( .A1(n4756), .A2(n5109), .ZN(n7377) );
  OAI21_X2 U6174 ( .B1(n5777), .B2(n7764), .A(n5776), .ZN(n5941) );
  NAND2_X1 U6175 ( .A1(n4540), .A2(n4539), .ZN(n4543) );
  NAND2_X1 U6176 ( .A1(n4433), .A2(n8083), .ZN(n8410) );
  AOI21_X1 U6177 ( .B1(n7438), .B2(n7450), .A(n7545), .ZN(n7439) );
  NOR2_X1 U6178 ( .A1(n7868), .A2(n7937), .ZN(n8082) );
  INV_X1 U6179 ( .A(n8081), .ZN(n4519) );
  OAI21_X1 U6180 ( .B1(n10317), .B2(n10352), .A(n4520), .ZN(n10320) );
  NAND2_X1 U6181 ( .A1(n10317), .A2(n10352), .ZN(n4520) );
  NOR2_X1 U6182 ( .A1(n9131), .A2(n9134), .ZN(n9021) );
  NOR2_X1 U6183 ( .A1(n8477), .A2(n8478), .ZN(n8482) );
  INV_X1 U6184 ( .A(n7541), .ZN(n4889) );
  NOR2_X1 U6185 ( .A1(n4853), .A2(n7541), .ZN(n4883) );
  OAI211_X1 U6186 ( .C1(n7542), .C2(n7541), .A(n4888), .B(n4886), .ZN(n4885)
         );
  NOR2_X1 U6187 ( .A1(n8532), .A2(n8533), .ZN(n8536) );
  NOR2_X2 U6188 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4932) );
  NAND2_X1 U6189 ( .A1(n9477), .A2(n9476), .ZN(n4522) );
  NAND2_X1 U6190 ( .A1(n4591), .A2(n4589), .ZN(n9475) );
  OAI22_X1 U6191 ( .A1(n9704), .A2(n9481), .B1(n10205), .B2(n10242), .ZN(n9685) );
  NAND2_X1 U6192 ( .A1(n7014), .A2(n7015), .ZN(n7013) );
  NOR2_X1 U6193 ( .A1(n8494), .A2(n8495), .ZN(n8499) );
  NOR2_X1 U6194 ( .A1(n8552), .A2(n8551), .ZN(n8571) );
  AND3_X2 U6195 ( .A1(n6382), .A2(n6171), .A3(n5012), .ZN(n6598) );
  AND2_X2 U6196 ( .A1(n4401), .A2(n6107), .ZN(n6171) );
  NOR2_X2 U6197 ( .A1(n8601), .A2(n8600), .ZN(n8615) );
  NAND2_X1 U6198 ( .A1(n4858), .A2(n4856), .ZN(n8458) );
  NAND2_X1 U6199 ( .A1(n4870), .A2(n4869), .ZN(n7545) );
  NOR2_X1 U6200 ( .A1(n10238), .A2(n8459), .ZN(n8494) );
  OAI21_X1 U6201 ( .B1(n4532), .B2(n4780), .A(n4526), .ZN(n4527) );
  INV_X1 U6202 ( .A(n5920), .ZN(n4534) );
  NAND2_X1 U6203 ( .A1(n5779), .A2(n5782), .ZN(n5597) );
  NAND2_X2 U6204 ( .A1(n4535), .A2(n5068), .ZN(n7304) );
  NAND3_X1 U6205 ( .A1(n8153), .A2(P2_REG0_REG_1__SCAN_IN), .A3(n8989), .ZN(
        n5062) );
  INV_X1 U6206 ( .A(n8989), .ZN(n5065) );
  INV_X1 U6207 ( .A(n8153), .ZN(n5064) );
  INV_X1 U6208 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n4537) );
  OR2_X1 U6209 ( .A1(n5941), .A2(n8617), .ZN(n4539) );
  NAND2_X1 U6210 ( .A1(n5941), .A2(n4504), .ZN(n4540) );
  NAND2_X1 U6211 ( .A1(n4545), .A2(n4546), .ZN(n5911) );
  NAND2_X1 U6212 ( .A1(n5899), .A2(n4547), .ZN(n4545) );
  INV_X1 U6213 ( .A(n4557), .ZN(n5849) );
  NAND2_X1 U6214 ( .A1(n5357), .A2(n4567), .ZN(n5060) );
  INV_X1 U6215 ( .A(n5650), .ZN(n5071) );
  INV_X1 U6216 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n4570) );
  INV_X1 U6217 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4569) );
  INV_X1 U6218 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n10013) );
  AND2_X2 U6219 ( .A1(n6598), .A2(n4990), .ZN(n5975) );
  NAND2_X1 U6220 ( .A1(n7020), .A2(n6976), .ZN(n6388) );
  NAND2_X1 U6221 ( .A1(n6111), .A2(n6112), .ZN(n7020) );
  NAND2_X1 U6222 ( .A1(n6111), .A2(n4479), .ZN(n6535) );
  NAND2_X1 U6223 ( .A1(n9495), .A2(n4423), .ZN(n4579) );
  NAND2_X1 U6224 ( .A1(n9495), .A2(n9494), .ZN(n9591) );
  NAND2_X1 U6225 ( .A1(n4927), .A2(n4925), .ZN(n4591) );
  AOI21_X2 U6226 ( .B1(n4585), .B2(n4589), .A(n4584), .ZN(n9737) );
  INV_X1 U6227 ( .A(n6641), .ZN(n6319) );
  NAND2_X2 U6228 ( .A1(n6605), .A2(n10223), .ZN(n6641) );
  OAI21_X1 U6229 ( .B1(n6133), .B2(n6625), .A(n4594), .ZN(n6110) );
  NAND3_X1 U6230 ( .A1(n10223), .A2(n6605), .A3(n9337), .ZN(n4594) );
  NAND2_X1 U6231 ( .A1(n5160), .A2(n5159), .ZN(n4595) );
  NAND2_X1 U6232 ( .A1(n5134), .A2(n5133), .ZN(n4596) );
  NAND3_X1 U6233 ( .A1(n4597), .A2(n4598), .A3(n4599), .ZN(n5963) );
  NOR2_X1 U6234 ( .A1(n8651), .A2(n4781), .ZN(n4610) );
  OAI21_X1 U6235 ( .B1(n8689), .B2(n4617), .A(n4424), .ZN(n8659) );
  OAI21_X1 U6236 ( .B1(n8689), .B2(n4614), .A(n4612), .ZN(n4611) );
  OR2_X1 U6237 ( .A1(n8689), .A2(n5631), .ZN(n4630) );
  NAND2_X1 U6238 ( .A1(n5098), .A2(n5097), .ZN(n5102) );
  NAND3_X1 U6239 ( .A1(n4819), .A2(n4817), .A3(n5078), .ZN(n5090) );
  NAND3_X1 U6240 ( .A1(n4819), .A2(n4817), .A3(n6629), .ZN(n4633) );
  OAI21_X1 U6241 ( .B1(n8895), .B2(n4636), .A(n4634), .ZN(n8779) );
  INV_X1 U6242 ( .A(n8895), .ZN(n4639) );
  NAND2_X1 U6243 ( .A1(n9224), .A2(n4651), .ZN(n4650) );
  OAI21_X1 U6244 ( .B1(n9224), .B2(n4652), .A(n4651), .ZN(n9245) );
  OAI21_X1 U6245 ( .B1(n9236), .B2(n4661), .A(n4658), .ZN(n9289) );
  NAND2_X1 U6246 ( .A1(n9208), .A2(n4660), .ZN(n4659) );
  INV_X1 U6247 ( .A(n9100), .ZN(n4660) );
  INV_X1 U6248 ( .A(n9208), .ZN(n4661) );
  NAND2_X2 U6249 ( .A1(n9207), .A2(n9208), .ZN(n9288) );
  NAND2_X2 U6250 ( .A1(n6722), .A2(n4662), .ZN(n9168) );
  INV_X1 U6251 ( .A(n8035), .ZN(n4663) );
  NAND2_X1 U6252 ( .A1(n6293), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4664) );
  NAND2_X1 U6253 ( .A1(n4664), .A2(n4665), .ZN(n6316) );
  NAND2_X1 U6254 ( .A1(n9186), .A2(n9073), .ZN(n9078) );
  NAND3_X1 U6255 ( .A1(n7056), .A2(n4478), .A3(n7061), .ZN(n4667) );
  NAND3_X1 U6256 ( .A1(n4667), .A2(n4428), .A3(n7149), .ZN(n7152) );
  INV_X1 U6257 ( .A(n4967), .ZN(n7102) );
  NAND2_X1 U6258 ( .A1(n6171), .A2(n6161), .ZN(n6381) );
  NAND3_X1 U6259 ( .A1(n4675), .A2(n4672), .A3(n4670), .ZN(n4669) );
  NAND3_X1 U6260 ( .A1(n8619), .A2(n4671), .A3(P2_U3893), .ZN(n4670) );
  NAND2_X1 U6261 ( .A1(n5636), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4676) );
  CLKBUF_X1 U6262 ( .A(n5636), .Z(n4677) );
  MUX2_X1 U6263 ( .A(n7777), .B(n7193), .S(n5636), .Z(n7250) );
  MUX2_X1 U6264 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n5636), .Z(n7195) );
  MUX2_X1 U6265 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n5636), .Z(n7417) );
  MUX2_X1 U6266 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n5636), .Z(n7445) );
  MUX2_X1 U6267 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n4677), .Z(n7535) );
  MUX2_X1 U6268 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n4677), .Z(n7683) );
  MUX2_X1 U6269 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n4677), .Z(n7778) );
  MUX2_X1 U6270 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n4677), .Z(n7869) );
  MUX2_X1 U6271 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n4677), .Z(n8086) );
  MUX2_X1 U6272 ( .A(n9811), .B(n8076), .S(n4677), .Z(n8413) );
  MUX2_X1 U6273 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n4677), .Z(n8437) );
  MUX2_X1 U6274 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n4677), .Z(n8460) );
  MUX2_X1 U6275 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n4677), .Z(n8483) );
  MUX2_X1 U6276 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n4677), .Z(n8511) );
  MUX2_X1 U6277 ( .A(n8509), .B(n8883), .S(n4677), .Z(n8537) );
  MUX2_X1 U6278 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n4677), .Z(n8562) );
  MUX2_X1 U6279 ( .A(n8774), .B(n8875), .S(n4677), .Z(n8586) );
  MUX2_X1 U6280 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n4677), .Z(n8588) );
  NAND3_X1 U6281 ( .A1(n7298), .A2(n4677), .A3(n7198), .ZN(n5943) );
  MUX2_X1 U6282 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6079), .S(n9324), .Z(n9330)
         );
  NAND2_X1 U6283 ( .A1(n5336), .A2(n4688), .ZN(n4687) );
  NAND2_X1 U6284 ( .A1(n4687), .A2(n4689), .ZN(n5373) );
  NAND2_X1 U6285 ( .A1(n6624), .A2(n6628), .ZN(n4698) );
  MUX2_X1 U6286 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n6624), .Z(n5161) );
  MUX2_X1 U6287 ( .A(n6636), .B(n6637), .S(n6624), .Z(n5175) );
  MUX2_X1 U6288 ( .A(n6646), .B(n6644), .S(n6624), .Z(n5190) );
  MUX2_X1 U6289 ( .A(n6653), .B(n9977), .S(n6624), .Z(n5207) );
  MUX2_X1 U6290 ( .A(n9979), .B(n6682), .S(n6624), .Z(n5210) );
  MUX2_X1 U6291 ( .A(n6785), .B(n6783), .S(n6624), .Z(n5235) );
  MUX2_X1 U6292 ( .A(n6804), .B(n6802), .S(n6624), .Z(n5258) );
  MUX2_X1 U6293 ( .A(n6873), .B(n5263), .S(n6624), .Z(n5265) );
  MUX2_X1 U6294 ( .A(n5284), .B(n9978), .S(n6624), .Z(n5298) );
  MUX2_X1 U6295 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n6624), .Z(n5318) );
  OR2_X1 U6296 ( .A1(n5573), .A2(n5572), .ZN(n4702) );
  NAND2_X1 U6297 ( .A1(n5500), .A2(n4706), .ZN(n4705) );
  NAND2_X1 U6298 ( .A1(n5500), .A2(n5499), .ZN(n5515) );
  NAND2_X1 U6299 ( .A1(n4705), .A2(n4709), .ZN(n5535) );
  OAI21_X1 U6300 ( .B1(n5732), .B2(n4724), .A(n4721), .ZN(n4713) );
  INV_X1 U6301 ( .A(n4715), .ZN(n4714) );
  OAI21_X1 U6302 ( .B1(n5732), .B2(n4718), .A(n4499), .ZN(n4715) );
  NAND2_X1 U6303 ( .A1(n4717), .A2(n6376), .ZN(n4716) );
  NAND2_X1 U6304 ( .A1(n6376), .A2(n4719), .ZN(n4718) );
  NAND2_X1 U6305 ( .A1(n5242), .A2(n4411), .ZN(n4730) );
  NAND2_X1 U6306 ( .A1(n4730), .A2(n4731), .ZN(n5317) );
  NAND2_X1 U6307 ( .A1(n5242), .A2(n4740), .ZN(n4735) );
  NAND2_X1 U6308 ( .A1(n5242), .A2(n5241), .ZN(n5262) );
  NAND2_X1 U6309 ( .A1(n4742), .A2(n4744), .ZN(n5451) );
  NAND2_X1 U6310 ( .A1(n5396), .A2(n4747), .ZN(n4742) );
  OAI21_X1 U6311 ( .B1(n7483), .B2(n7484), .A(n4756), .ZN(n10348) );
  NAND2_X1 U6312 ( .A1(n7483), .A2(n7484), .ZN(n4756) );
  NAND3_X1 U6313 ( .A1(n4425), .A2(n4412), .A3(n4757), .ZN(n5301) );
  NAND2_X1 U6314 ( .A1(n8802), .A2(n4767), .ZN(n4764) );
  NAND2_X1 U6315 ( .A1(n4764), .A2(n4765), .ZN(n5393) );
  NAND2_X1 U6316 ( .A1(n5748), .A2(n4775), .ZN(n4774) );
  OR2_X1 U6317 ( .A1(n5699), .A2(n8205), .ZN(n4777) );
  OR2_X1 U6318 ( .A1(n5699), .A2(n4774), .ZN(n4773) );
  INV_X1 U6319 ( .A(n8205), .ZN(n4775) );
  CLKBUF_X1 U6320 ( .A(n8747), .Z(n4782) );
  OAI21_X2 U6321 ( .B1(n8747), .B2(n4785), .A(n4783), .ZN(n8692) );
  OAI21_X1 U6322 ( .B1(n7707), .B2(n7704), .A(n5808), .ZN(n7816) );
  INV_X1 U6323 ( .A(n5597), .ZN(n5750) );
  AOI21_X1 U6324 ( .B1(n8675), .B2(n5908), .A(n5531), .ZN(n8663) );
  AOI21_X1 U6325 ( .B1(n8655), .B2(n8648), .A(n5917), .ZN(n5699) );
  NAND2_X1 U6326 ( .A1(n5750), .A2(n7320), .ZN(n7319) );
  NAND2_X1 U6327 ( .A1(n8048), .A2(n5296), .ZN(n8891) );
  NAND2_X1 U6328 ( .A1(n5393), .A2(n5853), .ZN(n8751) );
  NAND2_X1 U6329 ( .A1(n8046), .A2(n8050), .ZN(n8048) );
  NAND2_X1 U6330 ( .A1(n7376), .A2(n5788), .ZN(n7649) );
  NAND2_X2 U6331 ( .A1(n5075), .A2(n5074), .ZN(n5636) );
  NAND2_X1 U6332 ( .A1(n5407), .A2(n5406), .ZN(n8753) );
  OAI21_X2 U6333 ( .B1(n9580), .B2(n4809), .A(n4807), .ZN(n9549) );
  INV_X1 U6334 ( .A(n9566), .ZN(n4811) );
  NAND2_X1 U6335 ( .A1(n6288), .A2(n4813), .ZN(n9689) );
  NAND2_X1 U6336 ( .A1(n7498), .A2(n4815), .ZN(n4814) );
  NAND3_X1 U6337 ( .A1(n9444), .A2(n4821), .A3(n4820), .ZN(n4819) );
  OAI211_X2 U6338 ( .C1(n6641), .C2(n4824), .A(n4823), .B(n4822), .ZN(n4901)
         );
  OR2_X1 U6339 ( .A1(n6084), .A2(n5076), .ZN(n4822) );
  NAND2_X1 U6340 ( .A1(n6641), .A2(n6624), .ZN(n6084) );
  INV_X1 U6341 ( .A(n9324), .ZN(n4824) );
  INV_X1 U6342 ( .A(n4827), .ZN(n7341) );
  NAND2_X1 U6343 ( .A1(n7504), .A2(n10287), .ZN(n7809) );
  NOR2_X1 U6344 ( .A1(n7503), .A2(n7664), .ZN(n7504) );
  NAND2_X1 U6345 ( .A1(n4827), .A2(n4826), .ZN(n7503) );
  NAND2_X1 U6346 ( .A1(n9694), .A2(n4828), .ZN(n4831) );
  INV_X1 U6347 ( .A(n4831), .ZN(n9644) );
  INV_X1 U6348 ( .A(n7837), .ZN(n4832) );
  NAND2_X1 U6349 ( .A1(n4833), .A2(n4832), .ZN(n9709) );
  AND2_X1 U6350 ( .A1(n4843), .A2(n4842), .ZN(n8426) );
  NAND2_X1 U6351 ( .A1(n8425), .A2(n5272), .ZN(n4842) );
  NAND2_X1 U6352 ( .A1(n4844), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4843) );
  INV_X1 U6353 ( .A(n8425), .ZN(n4844) );
  NOR2_X1 U6354 ( .A1(n7422), .A2(n7384), .ZN(n4851) );
  INV_X1 U6355 ( .A(n4853), .ZN(n7539) );
  XNOR2_X2 U6356 ( .A(n8431), .B(n8411), .ZN(n8412) );
  NAND2_X1 U6357 ( .A1(n4859), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4857) );
  AND2_X1 U6358 ( .A1(n4864), .A2(n8085), .ZN(n8081) );
  INV_X1 U6359 ( .A(n7426), .ZN(n4867) );
  AND2_X1 U6360 ( .A1(n4868), .A2(n4872), .ZN(n7438) );
  OR2_X2 U6362 ( .A1(n7879), .A2(n4880), .ZN(n4877) );
  INV_X1 U6363 ( .A(n7879), .ZN(n4881) );
  NOR2_X1 U6364 ( .A1(n4883), .A2(n4451), .ZN(n4888) );
  OR2_X2 U6365 ( .A1(n7542), .A2(n4485), .ZN(n4884) );
  NAND3_X1 U6366 ( .A1(n4890), .A2(n4891), .A3(P2_REG2_REG_17__SCAN_IN), .ZN(
        n4892) );
  NAND2_X1 U6367 ( .A1(n4890), .A2(n4891), .ZN(n8573) );
  NOR2_X1 U6368 ( .A1(n8571), .A2(n4500), .ZN(n8596) );
  OR2_X1 U6369 ( .A1(n8571), .A2(n4506), .ZN(n4890) );
  OAI21_X1 U6370 ( .B1(n8571), .B2(n4500), .A(n8561), .ZN(n4891) );
  INV_X1 U6371 ( .A(n4892), .ZN(n8598) );
  AND2_X2 U6372 ( .A1(n4894), .A2(n4893), .ZN(n8579) );
  NAND2_X1 U6374 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4897) );
  NOR2_X2 U6375 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6105) );
  NAND2_X2 U6376 ( .A1(n4900), .A2(n4898), .ZN(n10223) );
  INV_X1 U6377 ( .A(n4901), .ZN(n6846) );
  NAND2_X1 U6378 ( .A1(n7186), .A2(n4904), .ZN(n4903) );
  NAND3_X1 U6379 ( .A1(n4903), .A2(n7398), .A3(n4902), .ZN(n7401) );
  NAND2_X1 U6380 ( .A1(n7801), .A2(n4431), .ZN(n4927) );
  NAND2_X1 U6381 ( .A1(n9490), .A2(n4494), .ZN(n9602) );
  NAND2_X1 U6382 ( .A1(n9602), .A2(n9493), .ZN(n9495) );
  NAND2_X1 U6383 ( .A1(n9490), .A2(n9489), .ZN(n9618) );
  NAND2_X1 U6384 ( .A1(n9475), .A2(n4474), .ZN(n9477) );
  OR2_X2 U6385 ( .A1(n6595), .A2(n4994), .ZN(n6594) );
  NAND2_X2 U6386 ( .A1(n6598), .A2(n5970), .ZN(n6595) );
  NAND2_X1 U6387 ( .A1(n4933), .A2(n4484), .ZN(n8159) );
  NAND2_X1 U6388 ( .A1(n8345), .A2(n4477), .ZN(n4933) );
  INV_X1 U6389 ( .A(n5021), .ZN(n4941) );
  INV_X1 U6390 ( .A(n7457), .ZN(n4943) );
  NAND2_X1 U6391 ( .A1(n4945), .A2(n4944), .ZN(n7740) );
  NAND4_X1 U6392 ( .A1(n4946), .A2(n7522), .A3(n4948), .A4(n4949), .ZN(n4945)
         );
  NOR2_X1 U6393 ( .A1(n7520), .A2(n7519), .ZN(n7523) );
  INV_X1 U6394 ( .A(n7639), .ZN(n4949) );
  NAND2_X1 U6395 ( .A1(n8221), .A2(n8204), .ZN(n8208) );
  NAND2_X1 U6396 ( .A1(n8200), .A2(n4482), .ZN(n8221) );
  AND2_X2 U6397 ( .A1(n5229), .A2(n5030), .ZN(n4954) );
  NAND2_X1 U6398 ( .A1(n5071), .A2(n4958), .ZN(n4960) );
  NAND3_X1 U6399 ( .A1(n4961), .A2(n6842), .A3(n6903), .ZN(n6892) );
  NAND2_X1 U6400 ( .A1(n6841), .A2(n6840), .ZN(n6903) );
  NAND2_X1 U6401 ( .A1(n6839), .A2(n6838), .ZN(n4961) );
  NAND2_X1 U6402 ( .A1(n4963), .A2(n9142), .ZN(n4964) );
  NAND2_X1 U6403 ( .A1(n4964), .A2(n9143), .ZN(n9146) );
  NAND2_X1 U6404 ( .A1(n9288), .A2(n4969), .ZN(n4968) );
  OAI211_X1 U6405 ( .C1(n9288), .C2(n4971), .A(n9300), .B(n4968), .ZN(n9130)
         );
  INV_X1 U6406 ( .A(n9175), .ZN(n9172) );
  OR2_X1 U6407 ( .A1(n5991), .A2(n4981), .ZN(n4976) );
  NAND2_X1 U6408 ( .A1(n5991), .A2(n4980), .ZN(n4979) );
  NAND4_X1 U6409 ( .A1(n7566), .A2(n7565), .A3(n4989), .A4(n4418), .ZN(n4984)
         );
  NAND3_X1 U6410 ( .A1(n7566), .A2(n7565), .A3(n4418), .ZN(n4987) );
  NAND2_X1 U6411 ( .A1(n9006), .A2(n9198), .ZN(n5008) );
  CLKBUF_X1 U6412 ( .A(n6994), .Z(n6995) );
  NAND2_X1 U6413 ( .A1(n5025), .A2(n5700), .ZN(n5701) );
  NAND2_X1 U6414 ( .A1(n5092), .A2(n7768), .ZN(n7370) );
  INV_X1 U6415 ( .A(n8408), .ZN(n5092) );
  CLKBUF_X1 U6416 ( .A(n8802), .Z(n8824) );
  NAND2_X1 U6417 ( .A1(n5111), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5066) );
  NAND2_X1 U6418 ( .A1(n4403), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6088) );
  INV_X1 U6419 ( .A(n4404), .ZN(n6046) );
  NAND2_X1 U6420 ( .A1(n6114), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6080) );
  INV_X1 U6421 ( .A(n9475), .ZN(n8006) );
  NAND2_X2 U6422 ( .A1(n6113), .A2(n6535), .ZN(n6409) );
  XNOR2_X1 U6423 ( .A(n8142), .B(n8399), .ZN(n8244) );
  INV_X1 U6424 ( .A(n5110), .ZN(n5458) );
  NAND2_X1 U6425 ( .A1(n6964), .A2(n6965), .ZN(n7056) );
  AOI21_X1 U6426 ( .B1(n9320), .B2(n9115), .A(n6837), .ZN(n6840) );
  INV_X1 U6427 ( .A(n6748), .ZN(n6970) );
  INV_X1 U6428 ( .A(n7001), .ZN(n9757) );
  AND2_X1 U6429 ( .A1(n5045), .A2(n5034), .ZN(n5009) );
  AND2_X1 U6430 ( .A1(n7739), .A2(n7744), .ZN(n5010) );
  AND2_X1 U6431 ( .A1(n7671), .A2(n7670), .ZN(n5011) );
  AND4_X1 U6432 ( .A1(n5969), .A2(n10010), .A3(n6161), .A4(n6583), .ZN(n5012)
         );
  OAI21_X1 U6433 ( .B1(n7710), .B2(n5753), .A(n5751), .ZN(n7703) );
  INV_X1 U6434 ( .A(n7239), .ZN(n7183) );
  NAND2_X1 U6435 ( .A1(n5663), .A2(n5662), .ZN(n5665) );
  OR2_X1 U6436 ( .A1(n8109), .A2(P2_D_REG_0__SCAN_IN), .ZN(n5013) );
  AND2_X1 U6437 ( .A1(n6350), .A2(n6349), .ZN(n10067) );
  OR2_X1 U6438 ( .A1(n4781), .A2(n8890), .ZN(n5014) );
  OR2_X1 U6439 ( .A1(n10197), .A2(n9483), .ZN(n5015) );
  NOR2_X1 U6440 ( .A1(n8175), .A2(n8320), .ZN(n5016) );
  OR2_X1 U6441 ( .A1(n4781), .A2(n8980), .ZN(n5017) );
  OR2_X1 U6442 ( .A1(n10293), .A2(n9261), .ZN(n5018) );
  INV_X1 U6443 ( .A(n7363), .ZN(n7764) );
  NOR2_X2 U6444 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n6289) );
  INV_X1 U6445 ( .A(n8387), .ZN(n8651) );
  INV_X1 U6446 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n5959) );
  AND2_X1 U6447 ( .A1(n5241), .A2(n5237), .ZN(n5020) );
  INV_X1 U6448 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n10016) );
  NOR2_X1 U6449 ( .A1(n5961), .A2(n8980), .ZN(n5689) );
  INV_X1 U6450 ( .A(n8755), .ZN(n5406) );
  XOR2_X1 U6451 ( .A(n8137), .B(n4406), .Z(n5021) );
  OR2_X1 U6452 ( .A1(n6612), .A2(n6611), .ZN(n5022) );
  AND2_X1 U6453 ( .A1(n7979), .A2(n7964), .ZN(n8912) );
  INV_X1 U6454 ( .A(n8912), .ZN(n5700) );
  AND4_X1 U6455 ( .A1(n6292), .A2(n6289), .A3(n6291), .A4(n6290), .ZN(n5023)
         );
  AND3_X1 U6456 ( .A1(n6292), .A2(n6314), .A3(n5967), .ZN(n5024) );
  XOR2_X1 U6457 ( .A(n5699), .B(n8205), .Z(n5025) );
  AND2_X1 U6458 ( .A1(n5712), .A2(n5711), .ZN(n5026) );
  INV_X1 U6459 ( .A(n9686), .ZN(n6304) );
  OR2_X1 U6460 ( .A1(n5957), .A2(n8792), .ZN(n5027) );
  AND2_X1 U6461 ( .A1(n9100), .A2(n9098), .ZN(n9233) );
  INV_X1 U6462 ( .A(n9738), .ZN(n6262) );
  INV_X1 U6463 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5034) );
  INV_X1 U6464 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5967) );
  INV_X1 U6465 ( .A(n8546), .ZN(n8547) );
  INV_X1 U6466 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5057) );
  INV_X1 U6467 ( .A(n10067), .ZN(n9503) );
  NOR2_X1 U6468 ( .A1(n7688), .A2(n4886), .ZN(n7789) );
  NAND2_X1 U6469 ( .A1(n7731), .A2(n8617), .ZN(n7367) );
  INV_X1 U6470 ( .A(n5073), .ZN(n5074) );
  OR2_X1 U6471 ( .A1(n9040), .A2(n9039), .ZN(n9041) );
  INV_X1 U6472 ( .A(n7558), .ZN(n7559) );
  AND2_X1 U6473 ( .A1(n6962), .A2(n6900), .ZN(n6902) );
  INV_X1 U6474 ( .A(n6041), .ZN(n6030) );
  INV_X1 U6475 ( .A(n6256), .ZN(n5983) );
  INV_X1 U6476 ( .A(n9461), .ZN(n9462) );
  OR2_X1 U6477 ( .A1(n6745), .A2(n4408), .ZN(n6505) );
  INV_X1 U6478 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5970) );
  INV_X1 U6479 ( .A(n5371), .ZN(n5372) );
  OR2_X1 U6480 ( .A1(n6381), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n6228) );
  OR2_X1 U6481 ( .A1(n8139), .A2(n8138), .ZN(n8140) );
  INV_X1 U6482 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5126) );
  INV_X1 U6483 ( .A(n8431), .ZN(n8432) );
  INV_X1 U6484 ( .A(n5921), .ZN(n5633) );
  INV_X1 U6485 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9823) );
  AND2_X1 U6486 ( .A1(n5703), .A2(n6617), .ZN(n5705) );
  INV_X1 U6487 ( .A(n6234), .ZN(n5982) );
  INV_X1 U6488 ( .A(n7103), .ZN(n7061) );
  AND2_X1 U6489 ( .A1(n9290), .A2(n9287), .ZN(n9111) );
  OR2_X1 U6490 ( .A1(n6043), .A2(n6031), .ZN(n6341) );
  NAND2_X1 U6491 ( .A1(n5988), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6009) );
  INV_X1 U6492 ( .A(n6364), .ZN(n6347) );
  NAND2_X1 U6493 ( .A1(n8216), .A2(n10219), .ZN(n5998) );
  INV_X1 U6494 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6920) );
  INV_X1 U6495 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7854) );
  INV_X1 U6496 ( .A(n9719), .ZN(n9480) );
  NAND2_X1 U6497 ( .A1(n10210), .A2(n9473), .ZN(n9474) );
  INV_X1 U6498 ( .A(n6746), .ZN(n6934) );
  INV_X1 U6499 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5971) );
  NOR2_X1 U6500 ( .A1(n6228), .A2(n6227), .ZN(n6230) );
  OR2_X1 U6501 ( .A1(n7901), .A2(n7894), .ZN(n7895) );
  INV_X1 U6502 ( .A(n8377), .ZN(n8358) );
  NAND2_X1 U6503 ( .A1(n7303), .A2(n7358), .ZN(n8379) );
  INV_X1 U6504 ( .A(n5592), .ZN(n5955) );
  INV_X1 U6505 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5069) );
  INV_X1 U6506 ( .A(n8448), .ZN(n8411) );
  XNOR2_X1 U6507 ( .A(n8213), .B(n8651), .ZN(n8205) );
  AND2_X1 U6508 ( .A1(n5901), .A2(n5906), .ZN(n8686) );
  INV_X1 U6509 ( .A(n8738), .ZN(n8769) );
  OR2_X1 U6510 ( .A1(n8917), .A2(n10231), .ZN(n10343) );
  INV_X1 U6511 ( .A(n7370), .ZN(n7320) );
  INV_X1 U6512 ( .A(n8395), .ZN(n8898) );
  INV_X1 U6513 ( .A(n8407), .ZN(n7461) );
  OR2_X1 U6514 ( .A1(n7297), .A2(n6986), .ZN(n7302) );
  INV_X1 U6515 ( .A(n9742), .ZN(n9473) );
  NAND2_X1 U6516 ( .A1(n8021), .A2(n8022), .ZN(n8023) );
  OR2_X1 U6517 ( .A1(n6065), .A2(n9190), .ZN(n6056) );
  OR2_X1 U6518 ( .A1(n6297), .A2(n6296), .ZN(n6308) );
  INV_X1 U6519 ( .A(n10154), .ZN(n9261) );
  NAND2_X1 U6520 ( .A1(n5981), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6234) );
  INV_X1 U6521 ( .A(n9303), .ZN(n9293) );
  OR2_X1 U6522 ( .A1(n6268), .A2(n7854), .ZN(n6282) );
  OR2_X1 U6523 ( .A1(n9176), .A2(n6355), .ZN(n6350) );
  INV_X1 U6524 ( .A(n9450), .ZN(n9445) );
  INV_X1 U6525 ( .A(n9505), .ZN(n9472) );
  INV_X1 U6526 ( .A(n10077), .ZN(n9555) );
  INV_X1 U6527 ( .A(n10143), .ZN(n9708) );
  INV_X1 U6528 ( .A(n10243), .ZN(n10155) );
  AND2_X1 U6529 ( .A1(n7999), .A2(n6454), .ZN(n7834) );
  INV_X1 U6530 ( .A(n8134), .ZN(n10287) );
  NAND2_X1 U6531 ( .A1(n9321), .A2(n6928), .ZN(n6927) );
  AND2_X1 U6532 ( .A1(n5516), .A2(n5504), .ZN(n5514) );
  NAND2_X1 U6533 ( .A1(n5451), .A2(n5450), .ZN(n5469) );
  INV_X1 U6534 ( .A(n8373), .ZN(n8344) );
  NAND2_X1 U6535 ( .A1(n7306), .A2(n10345), .ZN(n8367) );
  INV_X1 U6536 ( .A(n8618), .ZN(n10332) );
  AND2_X1 U6537 ( .A1(n8753), .A2(n8752), .ZN(n8870) );
  INV_X1 U6538 ( .A(n8792), .ZN(n8825) );
  OAI21_X1 U6539 ( .B1(n5961), .B2(n8890), .A(n5960), .ZN(n5962) );
  OR2_X1 U6540 ( .A1(n5947), .A2(n5946), .ZN(n5709) );
  NOR2_X1 U6541 ( .A1(n10372), .A2(n5690), .ZN(n5691) );
  AND2_X1 U6542 ( .A1(n6849), .A2(n6848), .ZN(n9303) );
  INV_X1 U6543 ( .A(n9305), .ZN(n9295) );
  OR2_X1 U6544 ( .A1(n9567), .A2(n6355), .ZN(n6049) );
  OR2_X1 U6545 ( .A1(n6664), .A2(n6660), .ZN(n9415) );
  INV_X1 U6546 ( .A(n9432), .ZN(n9436) );
  XNOR2_X1 U6547 ( .A(n9453), .B(n9445), .ZN(n9446) );
  INV_X1 U6548 ( .A(n9538), .ZN(n9536) );
  INV_X1 U6549 ( .A(n9481), .ZN(n9703) );
  NAND2_X1 U6550 ( .A1(n6792), .A2(n6791), .ZN(n10125) );
  AND2_X1 U6551 ( .A1(n7003), .A2(n9673), .ZN(n7001) );
  INV_X1 U6552 ( .A(n10299), .ZN(n10248) );
  NAND2_X1 U6553 ( .A1(n6734), .A2(n6733), .ZN(n6805) );
  AND2_X1 U6554 ( .A1(n6762), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7915) );
  NOR2_X1 U6555 ( .A1(n6231), .A2(n6253), .ZN(n7475) );
  XNOR2_X1 U6556 ( .A(n5120), .B(SI_2_), .ZN(n5118) );
  INV_X1 U6557 ( .A(n8381), .ZN(n8298) );
  AND2_X1 U6558 ( .A1(n7290), .A2(n7289), .ZN(n8373) );
  NAND2_X1 U6559 ( .A1(n5585), .A2(n5584), .ZN(n8387) );
  INV_X1 U6560 ( .A(n8713), .ZN(n8739) );
  OR2_X1 U6561 ( .A1(P2_U3150), .A2(n7222), .ZN(n10330) );
  INV_X1 U6562 ( .A(n10327), .ZN(n8602) );
  OR2_X1 U6563 ( .A1(n7249), .A2(n8622), .ZN(n8634) );
  INV_X1 U6564 ( .A(n8795), .ZN(n8810) );
  NAND2_X1 U6565 ( .A1(n10350), .A2(n10235), .ZN(n8792) );
  INV_X2 U6566 ( .A(n10350), .ZN(n10353) );
  NAND2_X1 U6567 ( .A1(n8925), .A2(n8908), .ZN(n8890) );
  INV_X1 U6568 ( .A(n8925), .ZN(n8924) );
  INV_X1 U6569 ( .A(n8268), .ZN(n8958) );
  AND2_X1 U6570 ( .A1(n5687), .A2(n5686), .ZN(n10375) );
  INV_X2 U6571 ( .A(n10375), .ZN(n10372) );
  INV_X1 U6572 ( .A(n6615), .ZN(n7300) );
  INV_X1 U6573 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6802) );
  INV_X1 U6574 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6628) );
  INV_X1 U6575 ( .A(n9443), .ZN(n9420) );
  INV_X1 U6576 ( .A(n9000), .ZN(n10293) );
  INV_X1 U6577 ( .A(n9300), .ZN(n9285) );
  NAND2_X1 U6578 ( .A1(n6078), .A2(n6077), .ZN(n10077) );
  NAND2_X1 U6579 ( .A1(n6004), .A2(n6003), .ZN(n10085) );
  OR2_X1 U6580 ( .A1(n6664), .A2(n6663), .ZN(n9432) );
  OR2_X1 U6581 ( .A1(n7003), .A2(n7002), .ZN(n9755) );
  INV_X1 U6582 ( .A(n9721), .ZN(n9759) );
  INV_X1 U6583 ( .A(n9751), .ZN(n9724) );
  NAND2_X1 U6584 ( .A1(n10316), .A2(n10248), .ZN(n10163) );
  AND2_X2 U6585 ( .A1(n6943), .A2(n6799), .ZN(n10316) );
  INV_X1 U6586 ( .A(n9713), .ZN(n10205) );
  INV_X1 U6587 ( .A(n10306), .ZN(n10304) );
  NAND2_X1 U6588 ( .A1(n6807), .A2(n6805), .ZN(n10265) );
  INV_X1 U6589 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7765) );
  INV_X1 U6590 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8116) );
  INV_X1 U6591 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6873) );
  INV_X1 U6592 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9979) );
  INV_X1 U6593 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10379) );
  INV_X1 U6594 ( .A(n8592), .ZN(P2_U3893) );
  OAI211_X1 U6595 ( .C1(n4445), .C2(n10353), .A(n5958), .B(n5027), .ZN(
        P2_U3204) );
  AND2_X2 U6596 ( .A1(n5321), .A2(n5032), .ZN(n5357) );
  NAND2_X1 U6597 ( .A1(n5037), .A2(n5049), .ZN(n5645) );
  NAND2_X1 U6598 ( .A1(n5645), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5036) );
  INV_X1 U6599 ( .A(n5037), .ZN(n5041) );
  INV_X1 U6600 ( .A(n5019), .ZN(n5039) );
  NAND2_X1 U6601 ( .A1(n5039), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5040) );
  MUX2_X1 U6602 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5040), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n5042) );
  INV_X1 U6603 ( .A(n5043), .ZN(n5044) );
  NAND2_X1 U6604 ( .A1(n5044), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U6605 ( .A1(n5397), .A2(n5045), .ZN(n5046) );
  NAND2_X1 U6606 ( .A1(n5046), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5047) );
  NAND2_X1 U6607 ( .A1(n5944), .A2(n8617), .ZN(n5702) );
  NAND2_X1 U6608 ( .A1(n5702), .A2(n7367), .ZN(n5048) );
  NAND3_X1 U6609 ( .A1(n7769), .A2(n8917), .A3(n5048), .ZN(n7979) );
  NAND2_X1 U6610 ( .A1(n7923), .A2(n10231), .ZN(n7964) );
  INV_X1 U6611 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5050) );
  NOR2_X1 U6612 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5053) );
  NOR2_X1 U6613 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5052) );
  NOR2_X1 U6614 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5051) );
  NAND4_X1 U6615 ( .A1(n5054), .A2(n5053), .A3(n5052), .A4(n5051), .ZN(n5055)
         );
  INV_X1 U6616 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5056) );
  NAND2_X1 U6617 ( .A1(n5060), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5061) );
  NAND2_X1 U6618 ( .A1(n5250), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5063) );
  NAND2_X1 U6619 ( .A1(n5128), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5067) );
  AND2_X4 U6620 ( .A1(n8153), .A2(n5065), .ZN(n5111) );
  NAND2_X1 U6621 ( .A1(n5650), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5072) );
  INV_X1 U6622 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6629) );
  INV_X1 U6623 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5076) );
  AND2_X1 U6624 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5077) );
  NAND2_X1 U6625 ( .A1(n5103), .A2(n5077), .ZN(n6091) );
  AND2_X1 U6626 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5078) );
  XNOR2_X1 U6627 ( .A(n5098), .B(n5097), .ZN(n6631) );
  NAND2_X1 U6628 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5079) );
  MUX2_X1 U6629 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5079), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5082) );
  BUF_X1 U6630 ( .A(n5080), .Z(n7201) );
  INV_X1 U6631 ( .A(n5080), .ZN(n5081) );
  NAND2_X1 U6632 ( .A1(n7304), .A2(n7826), .ZN(n5779) );
  NAND2_X1 U6633 ( .A1(n5250), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5087) );
  NAND2_X1 U6634 ( .A1(n5110), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5086) );
  NAND2_X1 U6635 ( .A1(n5111), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5085) );
  NAND2_X1 U6636 ( .A1(n5128), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5084) );
  NAND4_X1 U6637 ( .A1(n5087), .A2(n5086), .A3(n5085), .A4(n5084), .ZN(n8408)
         );
  NAND2_X1 U6638 ( .A1(n6624), .A2(SI_0_), .ZN(n5089) );
  INV_X1 U6639 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5088) );
  NAND2_X1 U6640 ( .A1(n5089), .A2(n5088), .ZN(n5091) );
  AND2_X1 U6641 ( .A1(n5091), .A2(n5090), .ZN(n8995) );
  MUX2_X1 U6642 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8995), .S(n5104), .Z(n7768) );
  INV_X1 U6643 ( .A(n7768), .ZN(n5754) );
  NAND2_X1 U6644 ( .A1(n7319), .A2(n5782), .ZN(n7483) );
  NAND2_X1 U6645 ( .A1(n5250), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5096) );
  NAND2_X1 U6646 ( .A1(n5110), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5095) );
  NAND2_X1 U6647 ( .A1(n5128), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5094) );
  NAND2_X1 U6648 ( .A1(n5111), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5093) );
  INV_X1 U6649 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6626) );
  OR2_X1 U6650 ( .A1(n5139), .A2(n6626), .ZN(n5108) );
  INV_X1 U6651 ( .A(n5099), .ZN(n5100) );
  NAND2_X1 U6652 ( .A1(n5100), .A2(SI_1_), .ZN(n5101) );
  NAND2_X1 U6653 ( .A1(n5102), .A2(n5101), .ZN(n5119) );
  INV_X1 U6654 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6622) );
  MUX2_X1 U6655 ( .A(n6626), .B(n6622), .S(n5103), .Z(n5120) );
  XNOR2_X1 U6656 ( .A(n5119), .B(n5118), .ZN(n6625) );
  OR2_X1 U6657 ( .A1(n5117), .A2(n6625), .ZN(n5107) );
  XNOR2_X1 U6658 ( .A(n8407), .B(n10344), .ZN(n5785) );
  INV_X1 U6659 ( .A(n10344), .ZN(n7361) );
  NAND2_X1 U6660 ( .A1(n7461), .A2(n7361), .ZN(n5109) );
  INV_X1 U6661 ( .A(n5250), .ZN(n5426) );
  OR2_X1 U6662 ( .A1(n5426), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5115) );
  NAND2_X1 U6663 ( .A1(n5110), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5114) );
  NAND2_X1 U6664 ( .A1(n5128), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5113) );
  NAND2_X1 U6665 ( .A1(n5111), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5112) );
  NAND2_X1 U6666 ( .A1(n5105), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5116) );
  XNOR2_X1 U6667 ( .A(n5116), .B(n5028), .ZN(n7416) );
  OR2_X1 U6668 ( .A1(n5139), .A2(n6628), .ZN(n5125) );
  NAND2_X1 U6669 ( .A1(n5119), .A2(n5118), .ZN(n5123) );
  INV_X1 U6670 ( .A(n5120), .ZN(n5121) );
  NAND2_X1 U6671 ( .A1(n5121), .A2(SI_2_), .ZN(n5122) );
  NAND2_X1 U6672 ( .A1(n5123), .A2(n5122), .ZN(n5134) );
  XNOR2_X1 U6673 ( .A(n5135), .B(SI_3_), .ZN(n5133) );
  XNOR2_X1 U6674 ( .A(n5134), .B(n5133), .ZN(n6627) );
  OR2_X1 U6675 ( .A1(n5117), .A2(n6627), .ZN(n5124) );
  OAI211_X1 U6676 ( .C1(n6619), .C2(n7416), .A(n5125), .B(n5124), .ZN(n7381)
         );
  NAND2_X1 U6677 ( .A1(n7656), .A2(n7381), .ZN(n5788) );
  INV_X1 U6678 ( .A(n7381), .ZN(n7697) );
  NAND2_X1 U6679 ( .A1(n8406), .A2(n7697), .ZN(n5802) );
  AND2_X1 U6680 ( .A1(n5788), .A2(n5802), .ZN(n7378) );
  NAND2_X1 U6681 ( .A1(n7377), .A2(n7378), .ZN(n7376) );
  NAND2_X1 U6682 ( .A1(n5110), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5132) );
  NAND2_X1 U6683 ( .A1(n5111), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5131) );
  NAND2_X1 U6684 ( .A1(n9822), .A2(n5126), .ZN(n5147) );
  NAND2_X1 U6685 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5127) );
  NAND2_X1 U6686 ( .A1(n5147), .A2(n5127), .ZN(n7723) );
  NAND2_X1 U6687 ( .A1(n5579), .A2(n7723), .ZN(n5130) );
  NAND2_X1 U6688 ( .A1(n5128), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5129) );
  INV_X1 U6689 ( .A(n5135), .ZN(n5136) );
  NAND2_X1 U6690 ( .A1(n5136), .A2(SI_3_), .ZN(n5137) );
  INV_X1 U6691 ( .A(SI_4_), .ZN(n5138) );
  XNOR2_X1 U6692 ( .A(n5161), .B(n5138), .ZN(n5159) );
  XNOR2_X1 U6693 ( .A(n5160), .B(n5159), .ZN(n6634) );
  OR2_X1 U6694 ( .A1(n5117), .A2(n6634), .ZN(n5144) );
  INV_X1 U6695 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6632) );
  OR2_X1 U6696 ( .A1(n5734), .A2(n6632), .ZN(n5143) );
  NAND2_X1 U6697 ( .A1(n5140), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5141) );
  OR2_X1 U6698 ( .A1(n6619), .A2(n7444), .ZN(n5142) );
  NAND2_X1 U6699 ( .A1(n8405), .A2(n7650), .ZN(n5790) );
  NAND2_X1 U6700 ( .A1(n5110), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5152) );
  NAND2_X1 U6701 ( .A1(n5111), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5151) );
  INV_X1 U6702 ( .A(n5147), .ZN(n5146) );
  NAND2_X1 U6703 ( .A1(n5146), .A2(n5145), .ZN(n5166) );
  NAND2_X1 U6704 ( .A1(n5147), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5148) );
  NAND2_X1 U6705 ( .A1(n5166), .A2(n5148), .ZN(n7716) );
  NAND2_X1 U6706 ( .A1(n5579), .A2(n7716), .ZN(n5150) );
  NAND2_X1 U6707 ( .A1(n5128), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5149) );
  NAND4_X1 U6708 ( .A1(n5152), .A2(n5151), .A3(n5150), .A4(n5149), .ZN(n8404)
         );
  INV_X1 U6709 ( .A(n5140), .ZN(n5154) );
  NAND2_X1 U6710 ( .A1(n5154), .A2(n5153), .ZN(n5156) );
  NAND2_X1 U6711 ( .A1(n5156), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5155) );
  MUX2_X1 U6712 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5155), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n5158) );
  INV_X1 U6713 ( .A(n5156), .ZN(n5157) );
  NAND2_X1 U6714 ( .A1(n5157), .A2(n9976), .ZN(n5193) );
  NAND2_X1 U6715 ( .A1(n5158), .A2(n5193), .ZN(n7534) );
  NAND2_X1 U6716 ( .A1(n5161), .A2(SI_4_), .ZN(n5162) );
  INV_X1 U6717 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6637) );
  INV_X1 U6718 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6636) );
  XNOR2_X1 U6719 ( .A(n5175), .B(SI_5_), .ZN(n5173) );
  XNOR2_X1 U6720 ( .A(n5174), .B(n5173), .ZN(n6638) );
  OR2_X1 U6721 ( .A1(n5117), .A2(n6638), .ZN(n5164) );
  OR2_X1 U6722 ( .A1(n5734), .A2(n6637), .ZN(n5163) );
  OAI211_X1 U6723 ( .C1(n6619), .C2(n7534), .A(n5164), .B(n5163), .ZN(n7717)
         );
  INV_X1 U6724 ( .A(n7717), .ZN(n7733) );
  OR2_X1 U6725 ( .A1(n8404), .A2(n7733), .ZN(n5792) );
  AND2_X1 U6726 ( .A1(n7712), .A2(n5792), .ZN(n5803) );
  NAND2_X1 U6727 ( .A1(n7713), .A2(n5803), .ZN(n5165) );
  NAND2_X1 U6728 ( .A1(n8404), .A2(n7733), .ZN(n5789) );
  NAND2_X1 U6729 ( .A1(n5165), .A2(n5789), .ZN(n7707) );
  NAND2_X1 U6730 ( .A1(n5111), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5171) );
  NAND2_X1 U6731 ( .A1(n5110), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5170) );
  NAND2_X1 U6732 ( .A1(n5166), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5167) );
  NAND2_X1 U6733 ( .A1(n5182), .A2(n5167), .ZN(n7737) );
  NAND2_X1 U6734 ( .A1(n5579), .A2(n7737), .ZN(n5169) );
  NAND2_X1 U6735 ( .A1(n5128), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5168) );
  NAND4_X1 U6736 ( .A1(n5171), .A2(n5170), .A3(n5169), .A4(n5168), .ZN(n8403)
         );
  NAND2_X1 U6737 ( .A1(n5193), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5172) );
  NAND2_X1 U6738 ( .A1(n5174), .A2(n5173), .ZN(n5178) );
  INV_X1 U6739 ( .A(n5175), .ZN(n5176) );
  NAND2_X1 U6740 ( .A1(n5176), .A2(SI_5_), .ZN(n5177) );
  XNOR2_X1 U6741 ( .A(n5190), .B(SI_6_), .ZN(n5188) );
  XNOR2_X1 U6742 ( .A(n5189), .B(n5188), .ZN(n6645) );
  OR2_X1 U6743 ( .A1(n5117), .A2(n6645), .ZN(n5180) );
  OR2_X1 U6744 ( .A1(n5734), .A2(n6644), .ZN(n5179) );
  OAI211_X1 U6745 ( .C1(n6619), .C2(n7687), .A(n5180), .B(n5179), .ZN(n7754)
         );
  INV_X1 U6746 ( .A(n7754), .ZN(n7745) );
  NAND2_X1 U6747 ( .A1(n8403), .A2(n7745), .ZN(n5793) );
  NAND2_X1 U6748 ( .A1(n5808), .A2(n5793), .ZN(n7704) );
  NAND2_X1 U6749 ( .A1(n5110), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5187) );
  NAND2_X1 U6750 ( .A1(n5111), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5186) );
  NAND2_X1 U6751 ( .A1(n5182), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5183) );
  NAND2_X1 U6752 ( .A1(n5199), .A2(n5183), .ZN(n7905) );
  NAND2_X1 U6753 ( .A1(n5579), .A2(n7905), .ZN(n5185) );
  NAND2_X1 U6754 ( .A1(n5128), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5184) );
  NAND4_X1 U6755 ( .A1(n5187), .A2(n5186), .A3(n5185), .A4(n5184), .ZN(n8402)
         );
  INV_X1 U6756 ( .A(n5190), .ZN(n5191) );
  NAND2_X1 U6757 ( .A1(n5191), .A2(SI_6_), .ZN(n5192) );
  XNOR2_X1 U6758 ( .A(n5207), .B(SI_7_), .ZN(n5205) );
  XNOR2_X1 U6759 ( .A(n5206), .B(n5205), .ZN(n6652) );
  OR2_X1 U6760 ( .A1(n5117), .A2(n6652), .ZN(n5198) );
  OR2_X1 U6761 ( .A1(n5734), .A2(n9977), .ZN(n5197) );
  NAND2_X1 U6762 ( .A1(n5214), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5195) );
  XNOR2_X1 U6763 ( .A(n5195), .B(n5194), .ZN(n7684) );
  OR2_X1 U6764 ( .A1(n6619), .A2(n7684), .ZN(n5196) );
  OR2_X1 U6765 ( .A1(n8402), .A2(n7902), .ZN(n5818) );
  NAND2_X1 U6766 ( .A1(n8402), .A2(n7902), .ZN(n7909) );
  NAND2_X1 U6767 ( .A1(n5818), .A2(n7909), .ZN(n7815) );
  NAND2_X1 U6768 ( .A1(n5111), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5204) );
  NAND2_X1 U6769 ( .A1(n5110), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5203) );
  NAND2_X1 U6770 ( .A1(n5199), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5200) );
  NAND2_X1 U6771 ( .A1(n5223), .A2(n5200), .ZN(n7959) );
  NAND2_X1 U6772 ( .A1(n5579), .A2(n7959), .ZN(n5202) );
  NAND2_X1 U6773 ( .A1(n5128), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5201) );
  NAND4_X1 U6774 ( .A1(n5204), .A2(n5203), .A3(n5202), .A4(n5201), .ZN(n8401)
         );
  INV_X1 U6775 ( .A(n5207), .ZN(n5208) );
  INV_X1 U6776 ( .A(SI_8_), .ZN(n5209) );
  NAND2_X1 U6777 ( .A1(n5210), .A2(n5209), .ZN(n5231) );
  INV_X1 U6778 ( .A(n5210), .ZN(n5211) );
  NAND2_X1 U6779 ( .A1(n5211), .A2(SI_8_), .ZN(n5212) );
  NAND2_X1 U6780 ( .A1(n5231), .A2(n5212), .ZN(n5232) );
  INV_X1 U6781 ( .A(n5232), .ZN(n5213) );
  XNOR2_X1 U6782 ( .A(n5233), .B(n5213), .ZN(n6683) );
  OR2_X1 U6783 ( .A1(n5117), .A2(n6683), .ZN(n5219) );
  OR2_X1 U6784 ( .A1(n5734), .A2(n6682), .ZN(n5218) );
  OAI21_X1 U6785 ( .B1(n5214), .B2(P2_IR_REG_7__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5216) );
  INV_X1 U6786 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5215) );
  XNOR2_X1 U6787 ( .A(n5216), .B(n5215), .ZN(n7875) );
  OR2_X1 U6788 ( .A1(n6619), .A2(n7875), .ZN(n5217) );
  NAND2_X1 U6789 ( .A1(n8401), .A2(n7956), .ZN(n5797) );
  AND2_X1 U6790 ( .A1(n5797), .A2(n7909), .ZN(n5811) );
  NAND2_X1 U6791 ( .A1(n7814), .A2(n5811), .ZN(n5220) );
  NAND2_X1 U6792 ( .A1(n5220), .A2(n5819), .ZN(n7928) );
  NAND2_X1 U6793 ( .A1(n5110), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5228) );
  NAND2_X1 U6794 ( .A1(n5111), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5227) );
  INV_X1 U6795 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5221) );
  NAND2_X1 U6796 ( .A1(n5223), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5224) );
  NAND2_X1 U6797 ( .A1(n5251), .A2(n5224), .ZN(n7936) );
  NAND2_X1 U6798 ( .A1(n5579), .A2(n7936), .ZN(n5226) );
  NAND2_X1 U6799 ( .A1(n5128), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5225) );
  NAND4_X1 U6800 ( .A1(n5228), .A2(n5227), .A3(n5226), .A4(n5225), .ZN(n8400)
         );
  OR2_X1 U6801 ( .A1(n4416), .A2(n5058), .ZN(n5230) );
  XNOR2_X1 U6802 ( .A(n5230), .B(n5229), .ZN(n8085) );
  NAND2_X1 U6803 ( .A1(n5235), .A2(n5234), .ZN(n5241) );
  INV_X1 U6804 ( .A(n5235), .ZN(n5236) );
  NAND2_X1 U6805 ( .A1(n5236), .A2(SI_9_), .ZN(n5237) );
  XNOR2_X1 U6806 ( .A(n5240), .B(n5020), .ZN(n6782) );
  NAND2_X1 U6807 ( .A1(n6782), .A2(n5733), .ZN(n5239) );
  OR2_X1 U6808 ( .A1(n5734), .A2(n6783), .ZN(n5238) );
  OAI211_X1 U6809 ( .C1(n6619), .C2(n8085), .A(n5239), .B(n5238), .ZN(n8072)
         );
  INV_X1 U6810 ( .A(n8072), .ZN(n7963) );
  OR2_X1 U6811 ( .A1(n8400), .A2(n7963), .ZN(n5820) );
  NAND2_X1 U6812 ( .A1(n8400), .A2(n7963), .ZN(n5813) );
  NAND2_X1 U6813 ( .A1(n5820), .A2(n5813), .ZN(n7932) );
  NAND2_X1 U6814 ( .A1(n5240), .A2(n5020), .ZN(n5242) );
  XNOR2_X1 U6815 ( .A(n5262), .B(n5257), .ZN(n6801) );
  NAND2_X1 U6816 ( .A1(n6801), .A2(n5733), .ZN(n5249) );
  NOR2_X1 U6817 ( .A1(n5243), .A2(n5058), .ZN(n5244) );
  MUX2_X1 U6818 ( .A(n5058), .B(n5244), .S(P2_IR_REG_10__SCAN_IN), .Z(n5247)
         );
  INV_X1 U6819 ( .A(n5245), .ZN(n5246) );
  INV_X1 U6820 ( .A(n8424), .ZN(n8414) );
  AOI22_X1 U6821 ( .A1(n5418), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5417), .B2(
        n8414), .ZN(n5248) );
  NAND2_X1 U6822 ( .A1(n5249), .A2(n5248), .ZN(n8251) );
  NAND2_X1 U6823 ( .A1(n5111), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5256) );
  NAND2_X1 U6824 ( .A1(n5110), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5255) );
  NAND2_X1 U6825 ( .A1(n5251), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5252) );
  NAND2_X1 U6826 ( .A1(n5273), .A2(n5252), .ZN(n8245) );
  NAND2_X1 U6827 ( .A1(n5579), .A2(n8245), .ZN(n5254) );
  NAND2_X1 U6828 ( .A1(n5128), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5253) );
  AND2_X1 U6829 ( .A1(n8918), .A2(n8399), .ZN(n5758) );
  INV_X1 U6830 ( .A(n5258), .ZN(n5259) );
  NAND2_X1 U6831 ( .A1(n5259), .A2(SI_10_), .ZN(n5260) );
  INV_X1 U6832 ( .A(SI_11_), .ZN(n5264) );
  INV_X1 U6833 ( .A(n5265), .ZN(n5266) );
  NAND2_X1 U6834 ( .A1(n5266), .A2(SI_11_), .ZN(n5267) );
  NAND2_X1 U6835 ( .A1(n5281), .A2(n5267), .ZN(n5282) );
  XNOR2_X1 U6836 ( .A(n5283), .B(n5282), .ZN(n6827) );
  NAND2_X1 U6837 ( .A1(n6827), .A2(n5733), .ZN(n5271) );
  NAND2_X1 U6838 ( .A1(n5245), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5268) );
  MUX2_X1 U6839 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5268), .S(
        P2_IR_REG_11__SCAN_IN), .Z(n5269) );
  AND2_X1 U6840 ( .A1(n5269), .A2(n4487), .ZN(n8448) );
  AOI22_X1 U6841 ( .A1(n5418), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5417), .B2(
        n8448), .ZN(n5270) );
  NAND2_X1 U6842 ( .A1(n5271), .A2(n5270), .ZN(n8342) );
  NAND2_X1 U6843 ( .A1(n5110), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5279) );
  INV_X1 U6844 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5272) );
  OR2_X1 U6845 ( .A1(n5582), .A2(n5272), .ZN(n5278) );
  OR2_X2 U6846 ( .A1(n5273), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5290) );
  NAND2_X1 U6847 ( .A1(n5273), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5274) );
  AND2_X1 U6848 ( .A1(n5290), .A2(n5274), .ZN(n8346) );
  OR2_X1 U6849 ( .A1(n5426), .A2(n8346), .ZN(n5277) );
  INV_X1 U6850 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n5275) );
  OR2_X1 U6851 ( .A1(n5640), .A2(n5275), .ZN(n5276) );
  OR2_X1 U6852 ( .A1(n8399), .A2(n8918), .ZN(n7986) );
  AND2_X1 U6853 ( .A1(n5829), .A2(n7986), .ZN(n5280) );
  XNOR2_X1 U6854 ( .A(n5300), .B(n5297), .ZN(n6889) );
  NAND2_X1 U6855 ( .A1(n6889), .A2(n5733), .ZN(n5287) );
  NAND2_X1 U6856 ( .A1(n4487), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5285) );
  XNOR2_X1 U6857 ( .A(n5285), .B(n5031), .ZN(n8466) );
  INV_X1 U6858 ( .A(n8466), .ZN(n8455) );
  AOI22_X1 U6859 ( .A1(n5418), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5417), .B2(
        n8455), .ZN(n5286) );
  NAND2_X1 U6860 ( .A1(n5110), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5295) );
  NAND2_X1 U6861 ( .A1(n5128), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5294) );
  INV_X1 U6862 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5288) );
  NAND2_X1 U6863 ( .A1(n5290), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5291) );
  NAND2_X1 U6864 ( .A1(n5306), .A2(n5291), .ZN(n8274) );
  NAND2_X1 U6865 ( .A1(n5579), .A2(n8274), .ZN(n5293) );
  NAND2_X1 U6866 ( .A1(n5111), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5292) );
  NAND4_X1 U6867 ( .A1(n5295), .A2(n5294), .A3(n5293), .A4(n5292), .ZN(n8397)
         );
  XNOR2_X1 U6868 ( .A(n8907), .B(n8397), .ZN(n8050) );
  OR2_X1 U6869 ( .A1(n8907), .A2(n8900), .ZN(n5296) );
  INV_X1 U6870 ( .A(n5298), .ZN(n5299) );
  XNOR2_X1 U6871 ( .A(n5318), .B(SI_13_), .ZN(n5315) );
  XNOR2_X1 U6872 ( .A(n5317), .B(n5315), .ZN(n6951) );
  NAND2_X1 U6873 ( .A1(n6951), .A2(n5733), .ZN(n5304) );
  NAND2_X1 U6874 ( .A1(n5301), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5302) );
  XNOR2_X1 U6875 ( .A(n5302), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8493) );
  AOI22_X1 U6876 ( .A1(n5418), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5417), .B2(
        n8493), .ZN(n5303) );
  NAND2_X1 U6877 ( .A1(n5111), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5311) );
  NAND2_X1 U6878 ( .A1(n5110), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5310) );
  INV_X1 U6879 ( .A(n5306), .ZN(n5305) );
  INV_X1 U6880 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8147) );
  NAND2_X1 U6881 ( .A1(n5306), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5307) );
  NAND2_X1 U6882 ( .A1(n5328), .A2(n5307), .ZN(n10229) );
  NAND2_X1 U6883 ( .A1(n5579), .A2(n10229), .ZN(n5309) );
  NAND2_X1 U6884 ( .A1(n5128), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5308) );
  NAND4_X1 U6885 ( .A1(n5311), .A2(n5310), .A3(n5309), .A4(n5308), .ZN(n8396)
         );
  NAND2_X1 U6886 ( .A1(n8892), .A2(n8819), .ZN(n5312) );
  NAND2_X1 U6887 ( .A1(n8891), .A2(n5312), .ZN(n5314) );
  OR2_X1 U6888 ( .A1(n8892), .A2(n8819), .ZN(n5313) );
  NAND2_X1 U6889 ( .A1(n5314), .A2(n5313), .ZN(n8802) );
  INV_X1 U6890 ( .A(n5315), .ZN(n5316) );
  NAND2_X1 U6891 ( .A1(n5317), .A2(n5316), .ZN(n5320) );
  NAND2_X1 U6892 ( .A1(n5318), .A2(SI_13_), .ZN(n5319) );
  NAND2_X1 U6893 ( .A1(n5320), .A2(n5319), .ZN(n5336) );
  MUX2_X1 U6894 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n5553), .Z(n5337) );
  XNOR2_X1 U6895 ( .A(n5337), .B(SI_14_), .ZN(n5334) );
  XNOR2_X1 U6896 ( .A(n5336), .B(n5334), .ZN(n7079) );
  NAND2_X1 U6897 ( .A1(n7079), .A2(n5733), .ZN(n5327) );
  OR2_X1 U6898 ( .A1(n5321), .A2(n5058), .ZN(n5324) );
  INV_X1 U6899 ( .A(n5324), .ZN(n5322) );
  NAND2_X1 U6900 ( .A1(n5322), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n5325) );
  INV_X1 U6901 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5323) );
  NAND2_X1 U6902 ( .A1(n5324), .A2(n5323), .ZN(n5339) );
  AOI22_X1 U6903 ( .A1(n5418), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5417), .B2(
        n8503), .ZN(n5326) );
  NAND2_X1 U6904 ( .A1(n5111), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5333) );
  NAND2_X1 U6905 ( .A1(n5110), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5332) );
  OR2_X2 U6906 ( .A1(n5328), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5345) );
  NAND2_X1 U6907 ( .A1(n5328), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5329) );
  NAND2_X1 U6908 ( .A1(n5345), .A2(n5329), .ZN(n8821) );
  NAND2_X1 U6909 ( .A1(n5579), .A2(n8821), .ZN(n5331) );
  NAND2_X1 U6910 ( .A1(n5128), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5330) );
  NAND4_X1 U6911 ( .A1(n5333), .A2(n5332), .A3(n5331), .A4(n5330), .ZN(n8395)
         );
  NAND2_X1 U6912 ( .A1(n8885), .A2(n8898), .ZN(n8803) );
  INV_X1 U6913 ( .A(n5334), .ZN(n5335) );
  NAND2_X1 U6914 ( .A1(n5337), .A2(SI_14_), .ZN(n5338) );
  MUX2_X1 U6915 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n5553), .Z(n5356) );
  XNOR2_X1 U6916 ( .A(n5356), .B(SI_15_), .ZN(n5353) );
  XNOR2_X1 U6917 ( .A(n5355), .B(n5353), .ZN(n7145) );
  NAND2_X1 U6918 ( .A1(n7145), .A2(n5733), .ZN(n5342) );
  NAND2_X1 U6919 ( .A1(n5339), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5340) );
  XNOR2_X1 U6920 ( .A(n5340), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8548) );
  AOI22_X1 U6921 ( .A1(n5418), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5417), .B2(
        n8548), .ZN(n5341) );
  NAND2_X1 U6922 ( .A1(n5342), .A2(n5341), .ZN(n8371) );
  NAND2_X1 U6923 ( .A1(n5111), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5350) );
  NAND2_X1 U6924 ( .A1(n5110), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5349) );
  INV_X1 U6925 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5343) );
  NAND2_X1 U6926 ( .A1(n5345), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5346) );
  NAND2_X1 U6927 ( .A1(n5363), .A2(n5346), .ZN(n8808) );
  NAND2_X1 U6928 ( .A1(n5579), .A2(n8808), .ZN(n5348) );
  NAND2_X1 U6929 ( .A1(n5128), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5347) );
  NAND4_X1 U6930 ( .A1(n5350), .A2(n5349), .A3(n5348), .A4(n5347), .ZN(n8783)
         );
  NAND2_X1 U6931 ( .A1(n8371), .A2(n8818), .ZN(n5871) );
  AND2_X1 U6932 ( .A1(n8803), .A2(n5871), .ZN(n5352) );
  INV_X1 U6933 ( .A(n5871), .ZN(n5351) );
  OR2_X1 U6934 ( .A1(n8371), .A2(n8818), .ZN(n8788) );
  MUX2_X1 U6935 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n5553), .Z(n5374) );
  XNOR2_X1 U6936 ( .A(n5374), .B(SI_16_), .ZN(n5371) );
  XNOR2_X1 U6937 ( .A(n5373), .B(n5371), .ZN(n7147) );
  NAND2_X1 U6938 ( .A1(n7147), .A2(n5733), .ZN(n5362) );
  NOR2_X1 U6939 ( .A1(n5357), .A2(n5058), .ZN(n5358) );
  MUX2_X1 U6940 ( .A(n5058), .B(n5358), .S(P2_IR_REG_16__SCAN_IN), .Z(n5359)
         );
  INV_X1 U6941 ( .A(n5359), .ZN(n5360) );
  AND2_X1 U6942 ( .A1(n5360), .A2(n5381), .ZN(n8556) );
  AOI22_X1 U6943 ( .A1(n5418), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5417), .B2(
        n8556), .ZN(n5361) );
  NAND2_X1 U6944 ( .A1(n5110), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5368) );
  INV_X1 U6945 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8534) );
  OR2_X1 U6946 ( .A1(n5582), .A2(n8534), .ZN(n5367) );
  NAND2_X1 U6947 ( .A1(n5363), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5364) );
  AND2_X1 U6948 ( .A1(n5387), .A2(n5364), .ZN(n8786) );
  OR2_X1 U6949 ( .A1(n5426), .A2(n8786), .ZN(n5366) );
  INV_X1 U6950 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8787) );
  OR2_X1 U6951 ( .A1(n5640), .A2(n8787), .ZN(n5365) );
  OR2_X1 U6952 ( .A1(n8877), .A2(n8801), .ZN(n5873) );
  NAND2_X1 U6953 ( .A1(n8877), .A2(n8801), .ZN(n5856) );
  NAND2_X1 U6954 ( .A1(n5873), .A2(n5856), .ZN(n8791) );
  INV_X1 U6955 ( .A(n8791), .ZN(n5369) );
  AND2_X1 U6956 ( .A1(n8788), .A2(n5369), .ZN(n5370) );
  NAND2_X1 U6957 ( .A1(n5373), .A2(n5372), .ZN(n5376) );
  NAND2_X1 U6958 ( .A1(n5374), .A2(SI_16_), .ZN(n5375) );
  NAND2_X1 U6959 ( .A1(n5376), .A2(n5375), .ZN(n5396) );
  MUX2_X1 U6960 ( .A(n7231), .B(n7230), .S(n5553), .Z(n5378) );
  INV_X1 U6961 ( .A(SI_17_), .ZN(n5377) );
  NAND2_X1 U6962 ( .A1(n5378), .A2(n5377), .ZN(n5394) );
  INV_X1 U6963 ( .A(n5378), .ZN(n5379) );
  NAND2_X1 U6964 ( .A1(n5379), .A2(SI_17_), .ZN(n5380) );
  NAND2_X1 U6965 ( .A1(n5394), .A2(n5380), .ZN(n5395) );
  XNOR2_X1 U6966 ( .A(n5396), .B(n5395), .ZN(n7229) );
  NAND2_X1 U6967 ( .A1(n7229), .A2(n5733), .ZN(n5384) );
  NAND2_X1 U6968 ( .A1(n5381), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5382) );
  XNOR2_X1 U6969 ( .A(n5382), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8597) );
  AOI22_X1 U6970 ( .A1(n5418), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5417), .B2(
        n8597), .ZN(n5383) );
  NAND2_X1 U6971 ( .A1(n5110), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5392) );
  INV_X1 U6972 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8875) );
  OR2_X1 U6973 ( .A1(n5582), .A2(n8875), .ZN(n5391) );
  INV_X1 U6974 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5385) );
  NAND2_X1 U6975 ( .A1(n5387), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5388) );
  AND2_X1 U6976 ( .A1(n5400), .A2(n5388), .ZN(n8773) );
  OR2_X1 U6977 ( .A1(n5426), .A2(n8773), .ZN(n5390) );
  INV_X1 U6978 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8774) );
  OR2_X1 U6979 ( .A1(n5640), .A2(n8774), .ZN(n5389) );
  NAND2_X1 U6980 ( .A1(n8772), .A2(n8757), .ZN(n5853) );
  INV_X1 U6981 ( .A(n8751), .ZN(n5407) );
  MUX2_X1 U6982 ( .A(n7357), .B(n9845), .S(n5553), .Z(n5409) );
  XNOR2_X1 U6983 ( .A(n5409), .B(SI_18_), .ZN(n5408) );
  XNOR2_X1 U6984 ( .A(n5412), .B(n5408), .ZN(n7355) );
  NAND2_X1 U6985 ( .A1(n7355), .A2(n5733), .ZN(n5399) );
  XNOR2_X1 U6986 ( .A(n5397), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8605) );
  AOI22_X1 U6987 ( .A1(n5418), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5417), .B2(
        n8605), .ZN(n5398) );
  NAND2_X1 U6988 ( .A1(n5110), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U6989 ( .A1(n5128), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5404) );
  OR2_X2 U6990 ( .A1(n5400), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5424) );
  NAND2_X1 U6991 ( .A1(n5400), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5401) );
  NAND2_X1 U6992 ( .A1(n5424), .A2(n5401), .ZN(n8759) );
  NAND2_X1 U6993 ( .A1(n5579), .A2(n8759), .ZN(n5403) );
  NAND2_X1 U6994 ( .A1(n5111), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5402) );
  NAND4_X1 U6995 ( .A1(n5405), .A2(n5404), .A3(n5403), .A4(n5402), .ZN(n8738)
         );
  NAND2_X1 U6996 ( .A1(n8868), .A2(n8769), .ZN(n5852) );
  NAND2_X1 U6997 ( .A1(n5876), .A2(n5852), .ZN(n8755) );
  NAND2_X1 U6998 ( .A1(n8753), .A2(n5876), .ZN(n8746) );
  INV_X1 U6999 ( .A(n5408), .ZN(n5411) );
  INV_X1 U7000 ( .A(n5409), .ZN(n5410) );
  MUX2_X1 U7001 ( .A(n7532), .B(n8116), .S(n5553), .Z(n5414) );
  INV_X1 U7002 ( .A(SI_19_), .ZN(n5413) );
  NAND2_X1 U7003 ( .A1(n5414), .A2(n5413), .ZN(n5432) );
  INV_X1 U7004 ( .A(n5414), .ZN(n5415) );
  NAND2_X1 U7005 ( .A1(n5415), .A2(SI_19_), .ZN(n5416) );
  NAND2_X1 U7006 ( .A1(n5432), .A2(n5416), .ZN(n5433) );
  XNOR2_X1 U7007 ( .A(n5434), .B(n5433), .ZN(n7531) );
  NAND2_X1 U7008 ( .A1(n7531), .A2(n5733), .ZN(n5420) );
  AOI22_X1 U7009 ( .A1(n5418), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8611), .B2(
        n5417), .ZN(n5419) );
  NAND2_X1 U7010 ( .A1(n5110), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5430) );
  INV_X1 U7011 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n5421) );
  OR2_X1 U7012 ( .A1(n5582), .A2(n5421), .ZN(n5429) );
  INV_X1 U7013 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5422) );
  NAND2_X1 U7014 ( .A1(n5424), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5425) );
  AND2_X1 U7015 ( .A1(n5441), .A2(n5425), .ZN(n8742) );
  OR2_X1 U7016 ( .A1(n5426), .A2(n8742), .ZN(n5428) );
  INV_X1 U7017 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n9980) );
  OR2_X1 U7018 ( .A1(n5640), .A2(n9980), .ZN(n5427) );
  NAND2_X1 U7019 ( .A1(n8744), .A2(n8758), .ZN(n5860) );
  AND2_X2 U7020 ( .A1(n8746), .A2(n8745), .ZN(n8864) );
  INV_X1 U7021 ( .A(n5431), .ZN(n5881) );
  MUX2_X1 U7022 ( .A(n9989), .B(n7752), .S(n5553), .Z(n5436) );
  INV_X1 U7023 ( .A(SI_20_), .ZN(n5435) );
  NAND2_X1 U7024 ( .A1(n5436), .A2(n5435), .ZN(n5450) );
  INV_X1 U7025 ( .A(n5436), .ZN(n5437) );
  NAND2_X1 U7026 ( .A1(n5437), .A2(SI_20_), .ZN(n5438) );
  XNOR2_X1 U7027 ( .A(n5449), .B(n5448), .ZN(n7730) );
  NAND2_X1 U7028 ( .A1(n7730), .A2(n5733), .ZN(n5440) );
  OR2_X1 U7029 ( .A1(n5734), .A2(n9989), .ZN(n5439) );
  OR2_X2 U7030 ( .A1(n5441), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5456) );
  NAND2_X1 U7031 ( .A1(n5441), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5442) );
  NAND2_X1 U7032 ( .A1(n5456), .A2(n5442), .ZN(n8730) );
  NAND2_X1 U7033 ( .A1(n5579), .A2(n8730), .ZN(n5447) );
  INV_X1 U7034 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8860) );
  OR2_X1 U7035 ( .A1(n5582), .A2(n8860), .ZN(n5446) );
  INV_X1 U7036 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8960) );
  OR2_X1 U7037 ( .A1(n5458), .A2(n8960), .ZN(n5445) );
  INV_X1 U7038 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n5443) );
  OR2_X1 U7039 ( .A1(n5640), .A2(n5443), .ZN(n5444) );
  MUX2_X1 U7040 ( .A(n7763), .B(n7765), .S(n5553), .Z(n5465) );
  XNOR2_X1 U7041 ( .A(n5465), .B(SI_21_), .ZN(n5464) );
  XNOR2_X1 U7042 ( .A(n5469), .B(n5464), .ZN(n7762) );
  NAND2_X1 U7043 ( .A1(n7762), .A2(n5733), .ZN(n5453) );
  OR2_X1 U7044 ( .A1(n5734), .A2(n7763), .ZN(n5452) );
  INV_X1 U7045 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5454) );
  NAND2_X1 U7046 ( .A1(n5456), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5457) );
  NAND2_X1 U7047 ( .A1(n5478), .A2(n5457), .ZN(n8718) );
  NAND2_X1 U7048 ( .A1(n5579), .A2(n8718), .ZN(n5463) );
  INV_X1 U7049 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n10033) );
  OR2_X1 U7050 ( .A1(n5582), .A2(n10033), .ZN(n5462) );
  INV_X1 U7051 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9972) );
  OR2_X1 U7052 ( .A1(n5458), .A2(n9972), .ZN(n5461) );
  INV_X1 U7053 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n5459) );
  OR2_X1 U7054 ( .A1(n5640), .A2(n5459), .ZN(n5460) );
  NAND2_X1 U7055 ( .A1(n8268), .A2(n8701), .ZN(n5891) );
  NAND2_X1 U7056 ( .A1(n8729), .A2(n8713), .ZN(n8714) );
  AND2_X1 U7057 ( .A1(n5891), .A2(n8714), .ZN(n5886) );
  INV_X1 U7058 ( .A(n5464), .ZN(n5468) );
  INV_X1 U7059 ( .A(n5465), .ZN(n5466) );
  NAND2_X1 U7060 ( .A1(n5466), .A2(SI_21_), .ZN(n5467) );
  INV_X1 U7061 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7920) );
  MUX2_X1 U7062 ( .A(n9990), .B(n7920), .S(n5553), .Z(n5471) );
  INV_X1 U7063 ( .A(SI_22_), .ZN(n5470) );
  NAND2_X1 U7064 ( .A1(n5471), .A2(n5470), .ZN(n5483) );
  INV_X1 U7065 ( .A(n5471), .ZN(n5472) );
  NAND2_X1 U7066 ( .A1(n5472), .A2(SI_22_), .ZN(n5473) );
  NAND2_X1 U7067 ( .A1(n5483), .A2(n5473), .ZN(n5484) );
  XNOR2_X1 U7068 ( .A(n5485), .B(n5484), .ZN(n7918) );
  NAND2_X1 U7069 ( .A1(n7918), .A2(n5733), .ZN(n5475) );
  OR2_X1 U7070 ( .A1(n5734), .A2(n9990), .ZN(n5474) );
  NAND2_X1 U7071 ( .A1(n5111), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5477) );
  NAND2_X1 U7072 ( .A1(n5110), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5476) );
  AND2_X1 U7073 ( .A1(n5477), .A2(n5476), .ZN(n5482) );
  OR2_X2 U7074 ( .A1(n5478), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5493) );
  NAND2_X1 U7075 ( .A1(n5478), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5479) );
  NAND2_X1 U7076 ( .A1(n5493), .A2(n5479), .ZN(n8705) );
  NAND2_X1 U7077 ( .A1(n8705), .A2(n5579), .ZN(n5481) );
  NAND2_X1 U7078 ( .A1(n5128), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5480) );
  NAND2_X1 U7079 ( .A1(n8331), .A2(n8712), .ZN(n5897) );
  OAI21_X1 U7080 ( .B1(n5485), .B2(n5484), .A(n5483), .ZN(n5498) );
  INV_X1 U7081 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5486) );
  MUX2_X1 U7082 ( .A(n9991), .B(n5486), .S(n5553), .Z(n5488) );
  INV_X1 U7083 ( .A(SI_23_), .ZN(n5487) );
  NAND2_X1 U7084 ( .A1(n5488), .A2(n5487), .ZN(n5499) );
  INV_X1 U7085 ( .A(n5488), .ZN(n5489) );
  NAND2_X1 U7086 ( .A1(n5489), .A2(SI_23_), .ZN(n5490) );
  XNOR2_X1 U7087 ( .A(n5498), .B(n5497), .ZN(n7925) );
  NAND2_X1 U7088 ( .A1(n7925), .A2(n5733), .ZN(n5492) );
  OR2_X1 U7089 ( .A1(n5734), .A2(n9991), .ZN(n5491) );
  INV_X1 U7090 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8848) );
  OR2_X2 U7091 ( .A1(n5493), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5509) );
  NAND2_X1 U7092 ( .A1(n5493), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5494) );
  NAND2_X1 U7093 ( .A1(n5509), .A2(n5494), .ZN(n8694) );
  NAND2_X1 U7094 ( .A1(n8694), .A2(n5579), .ZN(n5496) );
  AOI22_X1 U7095 ( .A1(n5128), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n5110), .B2(
        P2_REG0_REG_23__SCAN_IN), .ZN(n5495) );
  OAI211_X1 U7096 ( .C1(n5582), .C2(n8848), .A(n5496), .B(n5495), .ZN(n8392)
         );
  NAND2_X1 U7097 ( .A1(n5498), .A2(n5497), .ZN(n5500) );
  INV_X1 U7098 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8058) );
  MUX2_X1 U7099 ( .A(n9786), .B(n8058), .S(n5553), .Z(n5502) );
  INV_X1 U7100 ( .A(SI_24_), .ZN(n5501) );
  NAND2_X1 U7101 ( .A1(n5502), .A2(n5501), .ZN(n5516) );
  INV_X1 U7102 ( .A(n5502), .ZN(n5503) );
  NAND2_X1 U7103 ( .A1(n5503), .A2(SI_24_), .ZN(n5504) );
  XNOR2_X1 U7104 ( .A(n5515), .B(n5514), .ZN(n8057) );
  NAND2_X1 U7105 ( .A1(n8057), .A2(n5733), .ZN(n5506) );
  OR2_X1 U7106 ( .A1(n5734), .A2(n9786), .ZN(n5505) );
  INV_X1 U7107 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5507) );
  NAND2_X1 U7108 ( .A1(n5509), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5510) );
  NAND2_X1 U7109 ( .A1(n5524), .A2(n5510), .ZN(n8682) );
  NAND2_X1 U7110 ( .A1(n8682), .A2(n5579), .ZN(n5513) );
  AOI22_X1 U7111 ( .A1(n5111), .A2(P2_REG1_REG_24__SCAN_IN), .B1(n5110), .B2(
        P2_REG0_REG_24__SCAN_IN), .ZN(n5512) );
  NAND2_X1 U7112 ( .A1(n5128), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5511) );
  NAND2_X1 U7113 ( .A1(n8317), .A2(n8691), .ZN(n5906) );
  NAND2_X1 U7114 ( .A1(n8240), .A2(n8702), .ZN(n5905) );
  NAND2_X1 U7115 ( .A1(n5906), .A2(n5905), .ZN(n5900) );
  INV_X1 U7116 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8101) );
  INV_X1 U7117 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8099) );
  MUX2_X1 U7118 ( .A(n8101), .B(n8099), .S(n5553), .Z(n5517) );
  INV_X1 U7119 ( .A(SI_25_), .ZN(n9988) );
  NAND2_X1 U7120 ( .A1(n5517), .A2(n9988), .ZN(n5534) );
  INV_X1 U7121 ( .A(n5517), .ZN(n5518) );
  NAND2_X1 U7122 ( .A1(n5518), .A2(SI_25_), .ZN(n5519) );
  XNOR2_X1 U7123 ( .A(n5533), .B(n5532), .ZN(n8098) );
  NAND2_X1 U7124 ( .A1(n8098), .A2(n5733), .ZN(n5521) );
  OR2_X1 U7125 ( .A1(n5734), .A2(n8101), .ZN(n5520) );
  INV_X1 U7126 ( .A(n5524), .ZN(n5523) );
  INV_X1 U7127 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5522) );
  NAND2_X1 U7128 ( .A1(n5523), .A2(n5522), .ZN(n5541) );
  NAND2_X1 U7129 ( .A1(n5524), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5525) );
  NAND2_X1 U7130 ( .A1(n5541), .A2(n5525), .ZN(n8673) );
  NAND2_X1 U7131 ( .A1(n8673), .A2(n5579), .ZN(n5530) );
  INV_X1 U7132 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n10028) );
  NAND2_X1 U7133 ( .A1(n5110), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5527) );
  NAND2_X1 U7134 ( .A1(n5128), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5526) );
  OAI211_X1 U7135 ( .C1(n5582), .C2(n10028), .A(n5527), .B(n5526), .ZN(n5528)
         );
  INV_X1 U7136 ( .A(n5528), .ZN(n5529) );
  NAND2_X1 U7137 ( .A1(n8285), .A2(n8680), .ZN(n5908) );
  INV_X1 U7138 ( .A(n5909), .ZN(n5531) );
  NAND2_X1 U7139 ( .A1(n5535), .A2(n5534), .ZN(n5550) );
  INV_X1 U7140 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8107) );
  INV_X1 U7141 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8105) );
  MUX2_X1 U7142 ( .A(n8107), .B(n8105), .S(n5553), .Z(n5536) );
  INV_X1 U7143 ( .A(SI_26_), .ZN(n9818) );
  NAND2_X1 U7144 ( .A1(n5536), .A2(n9818), .ZN(n5551) );
  INV_X1 U7145 ( .A(n5536), .ZN(n5537) );
  NAND2_X1 U7146 ( .A1(n5537), .A2(SI_26_), .ZN(n5538) );
  XNOR2_X1 U7147 ( .A(n5550), .B(n5549), .ZN(n8104) );
  NAND2_X1 U7148 ( .A1(n8104), .A2(n5733), .ZN(n5540) );
  OR2_X1 U7149 ( .A1(n5734), .A2(n8107), .ZN(n5539) );
  NAND2_X1 U7150 ( .A1(n5541), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5542) );
  NAND2_X1 U7151 ( .A1(n5562), .A2(n5542), .ZN(n8664) );
  NAND2_X1 U7152 ( .A1(n8664), .A2(n5579), .ZN(n5548) );
  INV_X1 U7153 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n5545) );
  NAND2_X1 U7154 ( .A1(n5111), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5544) );
  NAND2_X1 U7155 ( .A1(n5110), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5543) );
  OAI211_X1 U7156 ( .C1(n5545), .C2(n5640), .A(n5544), .B(n5543), .ZN(n5546)
         );
  INV_X1 U7157 ( .A(n5546), .ZN(n5547) );
  NAND2_X1 U7158 ( .A1(n5550), .A2(n5549), .ZN(n5552) );
  INV_X1 U7159 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5557) );
  INV_X1 U7160 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10224) );
  MUX2_X1 U7161 ( .A(n5557), .B(n10224), .S(n5553), .Z(n5554) );
  INV_X1 U7162 ( .A(SI_27_), .ZN(n9820) );
  NAND2_X1 U7163 ( .A1(n5554), .A2(n9820), .ZN(n5571) );
  INV_X1 U7164 ( .A(n5554), .ZN(n5555) );
  NAND2_X1 U7165 ( .A1(n5555), .A2(SI_27_), .ZN(n5556) );
  NAND2_X1 U7166 ( .A1(n8110), .A2(n5733), .ZN(n5559) );
  OR2_X1 U7167 ( .A1(n5734), .A2(n5557), .ZN(n5558) );
  INV_X1 U7168 ( .A(n5562), .ZN(n5561) );
  INV_X1 U7169 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5560) );
  NAND2_X1 U7170 ( .A1(n5561), .A2(n5560), .ZN(n5577) );
  NAND2_X1 U7171 ( .A1(n5562), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5563) );
  NAND2_X1 U7172 ( .A1(n5577), .A2(n5563), .ZN(n8652) );
  NAND2_X1 U7173 ( .A1(n8652), .A2(n5579), .ZN(n5568) );
  INV_X1 U7174 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9925) );
  NAND2_X1 U7175 ( .A1(n5110), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5565) );
  NAND2_X1 U7176 ( .A1(n5128), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5564) );
  OAI211_X1 U7177 ( .C1(n9925), .C2(n5582), .A(n5565), .B(n5564), .ZN(n5566)
         );
  INV_X1 U7178 ( .A(n5566), .ZN(n5567) );
  AND2_X2 U7179 ( .A1(n5568), .A2(n5567), .ZN(n8661) );
  INV_X2 U7180 ( .A(n8661), .ZN(n8388) );
  XNOR2_X1 U7181 ( .A(n8653), .B(n8388), .ZN(n8648) );
  NOR2_X1 U7182 ( .A1(n8653), .A2(n8661), .ZN(n5917) );
  INV_X1 U7183 ( .A(n5569), .ZN(n5573) );
  INV_X1 U7184 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5574) );
  INV_X1 U7185 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8114) );
  MUX2_X1 U7186 ( .A(n5574), .B(n8114), .S(n5553), .Z(n5589) );
  XNOR2_X1 U7187 ( .A(n5589), .B(SI_28_), .ZN(n5586) );
  NAND2_X1 U7188 ( .A1(n8113), .A2(n5733), .ZN(n5576) );
  OR2_X1 U7189 ( .A1(n5734), .A2(n5574), .ZN(n5575) );
  NAND2_X1 U7190 ( .A1(n5577), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U7191 ( .A1(n5592), .A2(n5578), .ZN(n8643) );
  NAND2_X1 U7192 ( .A1(n8643), .A2(n5579), .ZN(n5585) );
  INV_X1 U7193 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9937) );
  NAND2_X1 U7194 ( .A1(n5128), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5581) );
  NAND2_X1 U7195 ( .A1(n5110), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5580) );
  OAI211_X1 U7196 ( .C1(n5582), .C2(n9937), .A(n5581), .B(n5580), .ZN(n5583)
         );
  INV_X1 U7197 ( .A(n5583), .ZN(n5584) );
  INV_X1 U7198 ( .A(SI_28_), .ZN(n5588) );
  INV_X1 U7199 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8988) );
  INV_X1 U7200 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10220) );
  MUX2_X1 U7201 ( .A(n8988), .B(n10220), .S(n5553), .Z(n5717) );
  NAND2_X1 U7202 ( .A1(n8986), .A2(n5733), .ZN(n5591) );
  OR2_X1 U7203 ( .A1(n5734), .A2(n8988), .ZN(n5590) );
  NAND2_X1 U7204 ( .A1(n5955), .A2(n5579), .ZN(n5741) );
  INV_X1 U7205 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n9856) );
  NAND2_X1 U7206 ( .A1(n5111), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U7207 ( .A1(n5110), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5593) );
  OAI211_X1 U7208 ( .C1(n9856), .C2(n5640), .A(n5594), .B(n5593), .ZN(n5595)
         );
  INV_X1 U7209 ( .A(n5595), .ZN(n5596) );
  NAND2_X1 U7210 ( .A1(n5688), .A2(n8211), .ZN(n5742) );
  XOR2_X1 U7211 ( .A(n5716), .B(n5921), .Z(n5957) );
  NAND2_X1 U7212 ( .A1(n8408), .A2(n7768), .ZN(n7321) );
  NAND2_X1 U7213 ( .A1(n5597), .A2(n7321), .ZN(n5599) );
  OR2_X1 U7214 ( .A1(n7304), .A2(n4763), .ZN(n5598) );
  NAND2_X1 U7215 ( .A1(n5599), .A2(n5598), .ZN(n7485) );
  NAND2_X1 U7216 ( .A1(n7485), .A2(n5785), .ZN(n5601) );
  OR2_X1 U7217 ( .A1(n8407), .A2(n7361), .ZN(n5600) );
  NAND2_X1 U7218 ( .A1(n5601), .A2(n5600), .ZN(n7379) );
  NOR2_X1 U7219 ( .A1(n8406), .A2(n7381), .ZN(n5602) );
  OAI22_X1 U7220 ( .A1(n7379), .A2(n5602), .B1(n7656), .B2(n7697), .ZN(n7653)
         );
  INV_X1 U7221 ( .A(n7653), .ZN(n5604) );
  NAND2_X1 U7222 ( .A1(n5604), .A2(n5603), .ZN(n7651) );
  INV_X1 U7223 ( .A(n7650), .ZN(n7724) );
  OR2_X1 U7224 ( .A1(n8405), .A2(n7724), .ZN(n5605) );
  NAND2_X1 U7225 ( .A1(n7651), .A2(n5605), .ZN(n7710) );
  NOR2_X1 U7226 ( .A1(n8404), .A2(n7717), .ZN(n5753) );
  NAND2_X1 U7227 ( .A1(n8404), .A2(n7717), .ZN(n5751) );
  OR2_X1 U7228 ( .A1(n8403), .A2(n7754), .ZN(n5606) );
  NAND2_X1 U7229 ( .A1(n7703), .A2(n5606), .ZN(n5608) );
  NAND2_X1 U7230 ( .A1(n8403), .A2(n7754), .ZN(n5607) );
  NAND2_X1 U7231 ( .A1(n5608), .A2(n5607), .ZN(n7818) );
  NAND2_X1 U7232 ( .A1(n7818), .A2(n7815), .ZN(n5610) );
  INV_X1 U7233 ( .A(n7902), .ZN(n7890) );
  NAND2_X1 U7234 ( .A1(n8402), .A2(n7890), .ZN(n5609) );
  NAND2_X1 U7235 ( .A1(n5610), .A2(n5609), .ZN(n7911) );
  NAND2_X1 U7236 ( .A1(n5819), .A2(n5797), .ZN(n7929) );
  INV_X1 U7237 ( .A(n8249), .ZN(n8398) );
  NAND2_X1 U7238 ( .A1(n8342), .A2(n8398), .ZN(n5616) );
  NAND2_X1 U7239 ( .A1(n8399), .A2(n8251), .ZN(n5615) );
  OR2_X1 U7240 ( .A1(n8400), .A2(n8072), .ZN(n7972) );
  NAND2_X1 U7241 ( .A1(n7911), .A2(n5612), .ZN(n5620) );
  INV_X1 U7242 ( .A(n5613), .ZN(n5618) );
  INV_X1 U7243 ( .A(n7956), .ZN(n7945) );
  NAND2_X1 U7244 ( .A1(n8401), .A2(n7945), .ZN(n7930) );
  NAND2_X1 U7245 ( .A1(n8400), .A2(n8072), .ZN(n5614) );
  AND2_X1 U7246 ( .A1(n7930), .A2(n5614), .ZN(n7971) );
  AND2_X1 U7247 ( .A1(n7971), .A2(n5615), .ZN(n7989) );
  AND2_X1 U7248 ( .A1(n7989), .A2(n5616), .ZN(n5617) );
  OR2_X1 U7249 ( .A1(n5618), .A2(n5617), .ZN(n5619) );
  NAND2_X1 U7250 ( .A1(n5620), .A2(n5619), .ZN(n8049) );
  AND2_X1 U7251 ( .A1(n8907), .A2(n8397), .ZN(n5621) );
  OAI22_X1 U7252 ( .A1(n8049), .A2(n5621), .B1(n8397), .B2(n8907), .ZN(n8895)
         );
  NOR2_X1 U7253 ( .A1(n8892), .A2(n8396), .ZN(n5842) );
  NAND2_X1 U7254 ( .A1(n8892), .A2(n8396), .ZN(n8814) );
  NAND2_X1 U7255 ( .A1(n8885), .A2(n8395), .ZN(n5622) );
  AND2_X1 U7256 ( .A1(n8814), .A2(n5622), .ZN(n5623) );
  OR2_X1 U7257 ( .A1(n8371), .A2(n8783), .ZN(n5624) );
  OR2_X1 U7258 ( .A1(n8885), .A2(n8395), .ZN(n8797) );
  AND2_X1 U7259 ( .A1(n5624), .A2(n8797), .ZN(n5625) );
  NAND2_X1 U7260 ( .A1(n8779), .A2(n8791), .ZN(n5627) );
  INV_X1 U7261 ( .A(n8801), .ZN(n8394) );
  NAND2_X1 U7262 ( .A1(n8877), .A2(n8394), .ZN(n5626) );
  NAND2_X1 U7263 ( .A1(n5627), .A2(n5626), .ZN(n8766) );
  NAND2_X1 U7264 ( .A1(n5875), .A2(n5853), .ZN(n8767) );
  NAND2_X1 U7265 ( .A1(n8772), .A2(n8781), .ZN(n5628) );
  AND2_X1 U7266 ( .A1(n8868), .A2(n8738), .ZN(n5629) );
  OR2_X1 U7267 ( .A1(n8868), .A2(n8738), .ZN(n5630) );
  NAND2_X1 U7268 ( .A1(n5887), .A2(n8714), .ZN(n8728) );
  NAND2_X1 U7269 ( .A1(n5889), .A2(n5891), .ZN(n8717) );
  NOR2_X1 U7270 ( .A1(n8240), .A2(n8392), .ZN(n5631) );
  INV_X1 U7271 ( .A(n8691), .ZN(n8391) );
  NAND2_X1 U7272 ( .A1(n5909), .A2(n5908), .ZN(n8674) );
  INV_X1 U7273 ( .A(n8285), .ZN(n8944) );
  INV_X1 U7274 ( .A(n8671), .ZN(n8389) );
  OAI21_X1 U7275 ( .B1(n8661), .B2(n8936), .A(n8649), .ZN(n5632) );
  NAND2_X1 U7276 ( .A1(n5944), .A2(n8611), .ZN(n5635) );
  NAND2_X1 U7277 ( .A1(n7363), .A2(n5939), .ZN(n5634) );
  INV_X1 U7278 ( .A(n7199), .ZN(n7198) );
  NAND2_X1 U7279 ( .A1(n7198), .A2(n8622), .ZN(n5637) );
  NAND2_X1 U7280 ( .A1(n6619), .A2(n5637), .ZN(n7358) );
  INV_X1 U7281 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n10031) );
  NAND2_X1 U7282 ( .A1(n5111), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5639) );
  NAND2_X1 U7283 ( .A1(n5110), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5638) );
  OAI211_X1 U7284 ( .C1(n10031), .C2(n5640), .A(n5639), .B(n5638), .ZN(n5641)
         );
  INV_X1 U7285 ( .A(n5641), .ZN(n5642) );
  AND2_X1 U7286 ( .A1(n5741), .A2(n5642), .ZN(n5746) );
  NAND2_X1 U7287 ( .A1(n6619), .A2(P2_B_REG_SCAN_IN), .ZN(n5643) );
  NAND2_X1 U7288 ( .A1(n8780), .A2(n5643), .ZN(n8636) );
  OAI22_X1 U7289 ( .A1(n8651), .A2(n8901), .B1(n5746), .B2(n8636), .ZN(n5644)
         );
  INV_X1 U7290 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5662) );
  NAND2_X1 U7291 ( .A1(n4463), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5648) );
  MUX2_X1 U7292 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5648), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5649) );
  NAND2_X1 U7293 ( .A1(n8103), .A2(n8109), .ZN(n6992) );
  XNOR2_X1 U7294 ( .A(P2_IR_REG_24__SCAN_IN), .B(P2_B_REG_SCAN_IN), .ZN(n5651)
         );
  NAND3_X1 U7295 ( .A1(n5652), .A2(P2_IR_REG_25__SCAN_IN), .A3(n5651), .ZN(
        n5659) );
  INV_X1 U7296 ( .A(n5652), .ZN(n5657) );
  NOR2_X1 U7297 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5654) );
  INV_X1 U7298 ( .A(P2_B_REG_SCAN_IN), .ZN(n5653) );
  AOI22_X1 U7299 ( .A1(n5654), .A2(P2_B_REG_SCAN_IN), .B1(n5653), .B2(
        P2_IR_REG_24__SCAN_IN), .ZN(n5655) );
  INV_X1 U7300 ( .A(n5655), .ZN(n5656) );
  NAND2_X1 U7301 ( .A1(n5657), .A2(n5656), .ZN(n5658) );
  NAND2_X1 U7302 ( .A1(n5659), .A2(n5658), .ZN(n7362) );
  INV_X1 U7303 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9996) );
  NAND2_X1 U7304 ( .A1(n5661), .A2(n9996), .ZN(n5660) );
  NAND2_X1 U7305 ( .A1(n5665), .A2(n5664), .ZN(n5677) );
  NAND2_X1 U7306 ( .A1(n5677), .A2(n8109), .ZN(n7366) );
  NOR2_X1 U7307 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .ZN(
        n5669) );
  NOR4_X1 U7308 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n5668) );
  NOR4_X1 U7309 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5667) );
  NOR4_X1 U7310 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n5666) );
  NAND4_X1 U7311 ( .A1(n5669), .A2(n5668), .A3(n5667), .A4(n5666), .ZN(n5675)
         );
  NOR4_X1 U7312 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5673) );
  NOR4_X1 U7313 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n5672) );
  NOR4_X1 U7314 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5671) );
  NOR4_X1 U7315 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n5670) );
  NAND4_X1 U7316 ( .A1(n5673), .A2(n5672), .A3(n5671), .A4(n5670), .ZN(n5674)
         );
  NOR2_X1 U7317 ( .A1(n5675), .A2(n5674), .ZN(n5676) );
  NAND2_X1 U7318 ( .A1(n5939), .A2(n8611), .ZN(n5682) );
  NOR2_X1 U7319 ( .A1(n5682), .A2(n7363), .ZN(n5683) );
  NAND2_X1 U7320 ( .A1(n5683), .A2(n5944), .ZN(n7288) );
  NAND2_X1 U7321 ( .A1(n7769), .A2(n7288), .ZN(n5684) );
  NAND2_X1 U7322 ( .A1(n7305), .A2(n5684), .ZN(n5687) );
  INV_X1 U7323 ( .A(n5708), .ZN(n5685) );
  NAND3_X1 U7324 ( .A1(n5947), .A2(n5685), .A3(n5946), .ZN(n7297) );
  INV_X1 U7325 ( .A(n7288), .ZN(n7293) );
  OR2_X1 U7326 ( .A1(n7302), .A2(n7295), .ZN(n5686) );
  NAND2_X1 U7327 ( .A1(n5963), .A2(n10372), .ZN(n5693) );
  INV_X1 U7328 ( .A(n5688), .ZN(n5961) );
  INV_X1 U7329 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5690) );
  NAND2_X1 U7330 ( .A1(n5693), .A2(n5692), .ZN(P2_U3456) );
  XNOR2_X1 U7331 ( .A(n5694), .B(n8205), .ZN(n5698) );
  INV_X1 U7332 ( .A(n8211), .ZN(n8386) );
  AND2_X1 U7333 ( .A1(n8386), .A2(n8780), .ZN(n5696) );
  AND2_X1 U7334 ( .A1(n8388), .A2(n8782), .ZN(n5695) );
  INV_X1 U7335 ( .A(n7964), .ZN(n8922) );
  OR2_X1 U7336 ( .A1(n5702), .A2(n7731), .ZN(n5703) );
  INV_X1 U7337 ( .A(n5705), .ZN(n5704) );
  OAI21_X1 U7338 ( .B1(n5952), .B2(n5949), .A(n5950), .ZN(n5710) );
  INV_X1 U7339 ( .A(n7367), .ZN(n5706) );
  OR2_X1 U7340 ( .A1(n6617), .A2(n5706), .ZN(n5707) );
  NAND2_X1 U7341 ( .A1(n7221), .A2(n5707), .ZN(n7292) );
  OR2_X1 U7342 ( .A1(n8925), .A2(n9937), .ZN(n5711) );
  NAND2_X1 U7343 ( .A1(n5026), .A2(n5014), .ZN(P2_U3487) );
  OR2_X1 U7344 ( .A1(n10372), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5713) );
  NAND2_X1 U7345 ( .A1(n5715), .A2(n5017), .ZN(P2_U3455) );
  INV_X1 U7346 ( .A(SI_29_), .ZN(n5720) );
  INV_X1 U7347 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8155) );
  INV_X1 U7348 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8218) );
  MUX2_X1 U7349 ( .A(n8155), .B(n8218), .S(n5553), .Z(n5722) );
  INV_X1 U7350 ( .A(SI_30_), .ZN(n9987) );
  NAND2_X1 U7351 ( .A1(n5722), .A2(n9987), .ZN(n5725) );
  INV_X1 U7352 ( .A(n5722), .ZN(n5723) );
  NAND2_X1 U7353 ( .A1(n5723), .A2(SI_30_), .ZN(n5724) );
  NAND2_X1 U7354 ( .A1(n5725), .A2(n5724), .ZN(n5731) );
  INV_X1 U7355 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n5729) );
  INV_X1 U7356 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n5726) );
  MUX2_X1 U7357 ( .A(n5729), .B(n5726), .S(n5553), .Z(n5727) );
  XNOR2_X1 U7358 ( .A(n5727), .B(SI_31_), .ZN(n5728) );
  NOR2_X1 U7359 ( .A1(n5734), .A2(n5729), .ZN(n5730) );
  NAND2_X1 U7360 ( .A1(n8154), .A2(n5733), .ZN(n5736) );
  OR2_X1 U7361 ( .A1(n5734), .A2(n8155), .ZN(n5735) );
  NAND2_X1 U7362 ( .A1(n5736), .A2(n5735), .ZN(n5745) );
  NAND2_X1 U7363 ( .A1(n5128), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n5739) );
  NAND2_X1 U7364 ( .A1(n5111), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n5738) );
  NAND2_X1 U7365 ( .A1(n5110), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5737) );
  AND3_X1 U7366 ( .A1(n5739), .A2(n5738), .A3(n5737), .ZN(n5740) );
  NAND2_X1 U7367 ( .A1(n5741), .A2(n5740), .ZN(n8638) );
  AND2_X1 U7368 ( .A1(n8929), .A2(n8638), .ZN(n5936) );
  AOI21_X1 U7369 ( .B1(n8929), .B2(n5745), .A(n5936), .ZN(n5744) );
  NAND2_X1 U7370 ( .A1(n5745), .A2(n5746), .ZN(n5929) );
  NAND2_X1 U7371 ( .A1(n5929), .A2(n5742), .ZN(n5931) );
  INV_X1 U7372 ( .A(n5931), .ZN(n5743) );
  INV_X1 U7373 ( .A(n5746), .ZN(n8385) );
  NAND2_X1 U7374 ( .A1(n8932), .A2(n8385), .ZN(n5926) );
  AOI21_X1 U7375 ( .B1(n8638), .B2(n5926), .A(n8929), .ZN(n5747) );
  NOR2_X1 U7376 ( .A1(n8929), .A2(n8638), .ZN(n5927) );
  INV_X1 U7377 ( .A(n5913), .ZN(n5749) );
  INV_X1 U7378 ( .A(n5905), .ZN(n8683) );
  NOR2_X1 U7379 ( .A1(n5903), .A2(n8683), .ZN(n8693) );
  INV_X1 U7380 ( .A(n8767), .ZN(n8770) );
  INV_X1 U7381 ( .A(n5751), .ZN(n5752) );
  OR2_X1 U7382 ( .A1(n5753), .A2(n5752), .ZN(n7714) );
  NAND3_X1 U7383 ( .A1(n7322), .A2(n7714), .A3(n7654), .ZN(n5756) );
  NAND2_X1 U7384 ( .A1(n8408), .A2(n5754), .ZN(n5778) );
  AND2_X1 U7385 ( .A1(n7370), .A2(n5778), .ZN(n7771) );
  NAND2_X1 U7386 ( .A1(n7378), .A2(n7771), .ZN(n5755) );
  NOR2_X1 U7387 ( .A1(n5756), .A2(n5755), .ZN(n5757) );
  INV_X1 U7388 ( .A(n7704), .ZN(n7706) );
  NAND4_X1 U7389 ( .A1(n5757), .A2(n4517), .A3(n7706), .A4(n7484), .ZN(n5759)
         );
  INV_X1 U7390 ( .A(n5758), .ZN(n5812) );
  NAND2_X1 U7391 ( .A1(n5812), .A2(n7986), .ZN(n7975) );
  NOR4_X1 U7392 ( .A1(n5759), .A2(n7975), .A3(n7932), .A4(n7929), .ZN(n5762)
         );
  INV_X1 U7393 ( .A(n8137), .ZN(n5761) );
  INV_X1 U7394 ( .A(n8814), .ZN(n5760) );
  OR2_X1 U7395 ( .A1(n5842), .A2(n5760), .ZN(n8894) );
  NAND4_X1 U7396 ( .A1(n5762), .A2(n5761), .A3(n8050), .A4(n8894), .ZN(n5763)
         );
  NAND2_X1 U7397 ( .A1(n8788), .A2(n5871), .ZN(n8806) );
  NAND2_X1 U7398 ( .A1(n8804), .A2(n8803), .ZN(n8823) );
  OR3_X1 U7399 ( .A1(n5763), .A2(n8806), .A3(n8823), .ZN(n5764) );
  NOR2_X1 U7400 ( .A1(n8791), .A2(n5764), .ZN(n5765) );
  NAND4_X1 U7401 ( .A1(n8745), .A2(n8770), .A3(n5406), .A4(n5765), .ZN(n5766)
         );
  OR2_X1 U7402 ( .A1(n8728), .A2(n5766), .ZN(n5767) );
  NOR2_X1 U7403 ( .A1(n8717), .A2(n5767), .ZN(n5768) );
  NAND4_X1 U7404 ( .A1(n8686), .A2(n8693), .A3(n8703), .A4(n5768), .ZN(n5769)
         );
  NOR2_X1 U7405 ( .A1(n8674), .A2(n5769), .ZN(n5770) );
  NAND3_X1 U7406 ( .A1(n8662), .A2(n8648), .A3(n5770), .ZN(n5771) );
  NOR2_X1 U7407 ( .A1(n8205), .A2(n5771), .ZN(n5772) );
  NAND4_X1 U7408 ( .A1(n5926), .A2(n5633), .A3(n5772), .A4(n5929), .ZN(n5773)
         );
  NOR3_X1 U7409 ( .A1(n5927), .A2(n5936), .A3(n5773), .ZN(n5774) );
  MUX2_X1 U7410 ( .A(n8387), .B(n8213), .S(n6617), .Z(n5923) );
  INV_X1 U7411 ( .A(n5923), .ZN(n5922) );
  AND2_X1 U7412 ( .A1(n5779), .A2(n5778), .ZN(n5781) );
  NAND3_X1 U7413 ( .A1(n7484), .A2(n7363), .A3(n5781), .ZN(n5780) );
  INV_X1 U7414 ( .A(n5781), .ZN(n5783) );
  NAND2_X1 U7415 ( .A1(n5783), .A2(n5782), .ZN(n5786) );
  NAND2_X1 U7416 ( .A1(n8407), .A2(n10344), .ZN(n5784) );
  OAI211_X1 U7417 ( .C1(n5786), .C2(n5785), .A(n5784), .B(n5802), .ZN(n5787)
         );
  INV_X1 U7418 ( .A(n5788), .ZN(n5791) );
  AND2_X1 U7419 ( .A1(n5793), .A2(n5789), .ZN(n5806) );
  OAI211_X1 U7420 ( .C1(n5805), .C2(n5791), .A(n5806), .B(n5790), .ZN(n5796)
         );
  INV_X1 U7421 ( .A(n5792), .ZN(n5794) );
  NAND2_X1 U7422 ( .A1(n5794), .A2(n5793), .ZN(n5795) );
  NAND4_X1 U7423 ( .A1(n5796), .A2(n5930), .A3(n5795), .A4(n5808), .ZN(n5801)
         );
  NAND2_X1 U7424 ( .A1(n5819), .A2(n5820), .ZN(n5799) );
  NAND2_X1 U7425 ( .A1(n5813), .A2(n5797), .ZN(n5798) );
  MUX2_X1 U7426 ( .A(n5799), .B(n5798), .S(n5930), .Z(n5810) );
  NOR2_X1 U7427 ( .A1(n5810), .A2(n7815), .ZN(n5800) );
  NAND2_X1 U7428 ( .A1(n5801), .A2(n5800), .ZN(n5835) );
  INV_X1 U7429 ( .A(n5802), .ZN(n5804) );
  OAI21_X1 U7430 ( .B1(n5805), .B2(n5804), .A(n5803), .ZN(n5807) );
  NAND2_X1 U7431 ( .A1(n5807), .A2(n5806), .ZN(n5809) );
  NAND2_X1 U7432 ( .A1(n5809), .A2(n5808), .ZN(n5817) );
  INV_X1 U7433 ( .A(n5810), .ZN(n5823) );
  INV_X1 U7434 ( .A(n5811), .ZN(n5815) );
  NAND4_X1 U7435 ( .A1(n5828), .A2(n6617), .A3(n5813), .A4(n5812), .ZN(n5814)
         );
  AOI21_X1 U7436 ( .B1(n5823), .B2(n5815), .A(n5814), .ZN(n5816) );
  OAI21_X1 U7437 ( .B1(n5835), .B2(n5817), .A(n5816), .ZN(n5837) );
  NAND2_X1 U7438 ( .A1(n5819), .A2(n5818), .ZN(n5822) );
  NAND4_X1 U7439 ( .A1(n5829), .A2(n5930), .A3(n5820), .A4(n7986), .ZN(n5821)
         );
  AOI21_X1 U7440 ( .B1(n5823), .B2(n5822), .A(n5821), .ZN(n5834) );
  NOR2_X1 U7441 ( .A1(n8249), .A2(n6617), .ZN(n5826) );
  NAND2_X1 U7442 ( .A1(n8249), .A2(n6617), .ZN(n5824) );
  NAND2_X1 U7443 ( .A1(n8342), .A2(n5824), .ZN(n5825) );
  OAI21_X1 U7444 ( .B1(n5826), .B2(n8342), .A(n5825), .ZN(n5832) );
  NOR2_X1 U7445 ( .A1(n8399), .A2(n5930), .ZN(n5827) );
  NAND3_X1 U7446 ( .A1(n5828), .A2(n5827), .A3(n8251), .ZN(n5831) );
  NAND4_X1 U7447 ( .A1(n5829), .A2(n5930), .A3(n8918), .A4(n8399), .ZN(n5830)
         );
  NAND3_X1 U7448 ( .A1(n5832), .A2(n5831), .A3(n5830), .ZN(n5833) );
  AOI21_X1 U7449 ( .B1(n5835), .B2(n5834), .A(n5833), .ZN(n5836) );
  NAND2_X1 U7450 ( .A1(n5837), .A2(n5836), .ZN(n5838) );
  NAND2_X1 U7451 ( .A1(n5838), .A2(n8050), .ZN(n5841) );
  MUX2_X1 U7452 ( .A(n5930), .B(n8900), .S(n8907), .Z(n5839) );
  OAI21_X1 U7453 ( .B1(n8397), .B2(n6617), .A(n5839), .ZN(n5840) );
  NAND2_X1 U7454 ( .A1(n5841), .A2(n5840), .ZN(n5846) );
  INV_X1 U7455 ( .A(n5842), .ZN(n5845) );
  MUX2_X1 U7456 ( .A(n8396), .B(n8892), .S(n5930), .Z(n5843) );
  INV_X1 U7457 ( .A(n5843), .ZN(n5844) );
  MUX2_X1 U7458 ( .A(n8803), .B(n8804), .S(n5930), .Z(n5847) );
  INV_X1 U7459 ( .A(n8806), .ZN(n5848) );
  NAND2_X1 U7460 ( .A1(n5849), .A2(n5848), .ZN(n5872) );
  NAND3_X1 U7461 ( .A1(n5872), .A2(n8788), .A3(n5873), .ZN(n5851) );
  AND2_X1 U7462 ( .A1(n5856), .A2(n5930), .ZN(n5850) );
  NAND2_X1 U7463 ( .A1(n5851), .A2(n5850), .ZN(n5857) );
  NAND2_X1 U7464 ( .A1(n5857), .A2(n8770), .ZN(n5854) );
  NAND3_X1 U7465 ( .A1(n5854), .A2(n5853), .A3(n5852), .ZN(n5855) );
  NAND2_X1 U7466 ( .A1(n5855), .A2(n5930), .ZN(n5859) );
  NAND3_X1 U7467 ( .A1(n5857), .A2(n8770), .A3(n5856), .ZN(n5858) );
  NAND2_X1 U7468 ( .A1(n5859), .A2(n5858), .ZN(n5879) );
  NAND2_X1 U7469 ( .A1(n5860), .A2(n5930), .ZN(n5870) );
  INV_X1 U7470 ( .A(n8744), .ZN(n8863) );
  NAND2_X1 U7471 ( .A1(n8738), .A2(n5930), .ZN(n5861) );
  NAND2_X1 U7472 ( .A1(n8725), .A2(n5930), .ZN(n5862) );
  OAI21_X1 U7473 ( .B1(n8868), .B2(n5861), .A(n5862), .ZN(n5867) );
  OAI21_X1 U7474 ( .B1(n5930), .B2(n8738), .A(n8868), .ZN(n5866) );
  INV_X1 U7475 ( .A(n5862), .ZN(n5863) );
  AND2_X1 U7476 ( .A1(n5863), .A2(n8738), .ZN(n5864) );
  OR2_X1 U7477 ( .A1(n8868), .A2(n5864), .ZN(n5865) );
  AOI22_X1 U7478 ( .A1(n8863), .A2(n5867), .B1(n5866), .B2(n5865), .ZN(n5869)
         );
  NAND3_X1 U7479 ( .A1(n8744), .A2(n8758), .A3(n6617), .ZN(n5868) );
  OAI211_X1 U7480 ( .C1(n5879), .C2(n5870), .A(n5869), .B(n5868), .ZN(n5884)
         );
  NAND2_X1 U7481 ( .A1(n5872), .A2(n5871), .ZN(n5874) );
  NAND2_X1 U7482 ( .A1(n5874), .A2(n5873), .ZN(n5878) );
  NAND3_X1 U7483 ( .A1(n5876), .A2(n6617), .A3(n5875), .ZN(n5877) );
  AOI21_X1 U7484 ( .B1(n5879), .B2(n5878), .A(n5877), .ZN(n5883) );
  NAND2_X1 U7485 ( .A1(n8714), .A2(n5930), .ZN(n5880) );
  OAI21_X1 U7486 ( .B1(n8728), .B2(n5881), .A(n5880), .ZN(n5882) );
  OAI21_X1 U7487 ( .B1(n5884), .B2(n5883), .A(n5882), .ZN(n5885) );
  OAI21_X1 U7488 ( .B1(n5930), .B2(n5886), .A(n5885), .ZN(n5890) );
  AOI21_X1 U7489 ( .B1(n5889), .B2(n5887), .A(n6617), .ZN(n5888) );
  AOI21_X1 U7490 ( .B1(n5890), .B2(n5889), .A(n5888), .ZN(n5893) );
  OAI21_X1 U7491 ( .B1(n6617), .B2(n5891), .A(n8703), .ZN(n5892) );
  OR2_X1 U7492 ( .A1(n5893), .A2(n5892), .ZN(n5899) );
  INV_X1 U7493 ( .A(n5894), .ZN(n5895) );
  NOR2_X1 U7494 ( .A1(n5903), .A2(n5895), .ZN(n5896) );
  MUX2_X1 U7495 ( .A(n5897), .B(n5896), .S(n5930), .Z(n5898) );
  INV_X1 U7496 ( .A(n5900), .ZN(n5902) );
  INV_X1 U7497 ( .A(n5901), .ZN(n5904) );
  INV_X1 U7498 ( .A(n5906), .ZN(n5907) );
  MUX2_X1 U7499 ( .A(n5909), .B(n5908), .S(n6617), .Z(n5910) );
  OAI21_X1 U7500 ( .B1(n5911), .B2(n8674), .A(n5910), .ZN(n5916) );
  INV_X1 U7501 ( .A(n8648), .ZN(n8654) );
  INV_X1 U7502 ( .A(n5912), .ZN(n5914) );
  MUX2_X1 U7503 ( .A(n5914), .B(n5913), .S(n6617), .Z(n5915) );
  AOI211_X1 U7504 ( .C1(n5916), .C2(n8662), .A(n8654), .B(n5915), .ZN(n5920)
         );
  NOR2_X1 U7505 ( .A1(n8936), .A2(n8388), .ZN(n5918) );
  MUX2_X1 U7506 ( .A(n5918), .B(n5917), .S(n6617), .Z(n5919) );
  NAND3_X1 U7507 ( .A1(n5932), .A2(n5926), .A3(n5924), .ZN(n5925) );
  AOI211_X1 U7508 ( .C1(n4781), .C2(n5933), .A(n5927), .B(n5925), .ZN(n5935)
         );
  INV_X1 U7509 ( .A(n5926), .ZN(n5928) );
  AOI211_X1 U7510 ( .C1(n5930), .C2(n5929), .A(n5928), .B(n5927), .ZN(n5934)
         );
  OAI21_X1 U7511 ( .B1(n5935), .B2(n5934), .A(n4527), .ZN(n5938) );
  INV_X1 U7512 ( .A(n5936), .ZN(n5937) );
  NAND2_X1 U7513 ( .A1(n5938), .A2(n5937), .ZN(n5940) );
  OR2_X1 U7514 ( .A1(n7219), .A2(P2_U3151), .ZN(n7926) );
  INV_X1 U7515 ( .A(n7926), .ZN(n5942) );
  NOR2_X1 U7516 ( .A1(n6986), .A2(n7769), .ZN(n7298) );
  OAI211_X1 U7517 ( .C1(n5944), .C2(n7926), .A(n5943), .B(P2_B_REG_SCAN_IN), 
        .ZN(n5945) );
  NAND2_X1 U7518 ( .A1(n5947), .A2(n5946), .ZN(n5948) );
  NAND4_X1 U7519 ( .A1(n5951), .A2(n5950), .A3(n5949), .A4(n5948), .ZN(n5954)
         );
  INV_X1 U7520 ( .A(n5952), .ZN(n5953) );
  NOR2_X2 U7521 ( .A1(n5954), .A2(n10343), .ZN(n8795) );
  NAND2_X1 U7522 ( .A1(n5955), .A2(n8822), .ZN(n8639) );
  OAI21_X1 U7523 ( .B1(n10350), .B2(n9856), .A(n8639), .ZN(n5956) );
  NAND2_X1 U7524 ( .A1(n10231), .A2(n7363), .ZN(n10342) );
  NAND2_X1 U7525 ( .A1(n7979), .A2(n10342), .ZN(n10235) );
  OR2_X1 U7526 ( .A1(n8925), .A2(n5959), .ZN(n5960) );
  AOI21_X1 U7527 ( .B1(n5963), .B2(n8925), .A(n5962), .ZN(n5964) );
  INV_X1 U7528 ( .A(n5964), .ZN(P2_U3488) );
  NOR2_X1 U7529 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5969) );
  INV_X1 U7530 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5972) );
  INV_X1 U7531 ( .A(n5991), .ZN(n5973) );
  NAND2_X2 U7532 ( .A1(n5974), .A2(n5973), .ZN(n6605) );
  NAND2_X1 U7533 ( .A1(n8057), .A2(n6376), .ZN(n5977) );
  NAND2_X1 U7534 ( .A1(n6370), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5976) );
  NAND3_X1 U7535 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n6152) );
  INV_X1 U7536 ( .A(n6152), .ZN(n5978) );
  NAND2_X1 U7537 ( .A1(n5978), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6187) );
  INV_X1 U7538 ( .A(n6187), .ZN(n5979) );
  NAND2_X1 U7539 ( .A1(n5979), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6189) );
  INV_X1 U7540 ( .A(n6189), .ZN(n5980) );
  INV_X1 U7541 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6296) );
  INV_X1 U7542 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9249) );
  INV_X1 U7543 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9190) );
  INV_X1 U7544 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9241) );
  NAND2_X1 U7545 ( .A1(n6009), .A2(n9241), .ZN(n5989) );
  AND2_X1 U7546 ( .A1(n6041), .A2(n5989), .ZN(n9585) );
  OAI21_X1 U7547 ( .B1(n5991), .B2(n10213), .A(P1_IR_REG_29__SCAN_IN), .ZN(
        n5994) );
  NAND2_X1 U7548 ( .A1(n9585), .A2(n6299), .ZN(n6004) );
  INV_X1 U7549 ( .A(n5997), .ZN(n8216) );
  INV_X1 U7550 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n6001) );
  NAND2_X1 U7551 ( .A1(n4404), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6000) );
  NAND2_X1 U7552 ( .A1(n6366), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5999) );
  OAI211_X1 U7553 ( .C1(n6347), .C2(n6001), .A(n6000), .B(n5999), .ZN(n6002)
         );
  INV_X1 U7554 ( .A(n6002), .ZN(n6003) );
  INV_X1 U7555 ( .A(n10085), .ZN(n9150) );
  NAND2_X1 U7556 ( .A1(n10096), .A2(n9150), .ZN(n6494) );
  NAND2_X1 U7557 ( .A1(n7925), .A2(n6376), .ZN(n6006) );
  INV_X1 U7558 ( .A(n6120), .ZN(n6138) );
  NAND2_X1 U7559 ( .A1(n6370), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6005) );
  INV_X1 U7560 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U7561 ( .A1(n6019), .A2(n6007), .ZN(n6008) );
  NAND2_X1 U7562 ( .A1(n6009), .A2(n6008), .ZN(n9148) );
  INV_X1 U7563 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9802) );
  NAND2_X1 U7564 ( .A1(n4404), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6011) );
  NAND2_X1 U7565 ( .A1(n6366), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6010) );
  OAI211_X1 U7566 ( .C1(n6347), .C2(n9802), .A(n6011), .B(n6010), .ZN(n6012)
         );
  INV_X1 U7567 ( .A(n6012), .ZN(n6013) );
  OR2_X1 U7568 ( .A1(n10100), .A2(n9496), .ZN(n6490) );
  NAND2_X1 U7569 ( .A1(n7918), .A2(n6376), .ZN(n6016) );
  NAND2_X1 U7570 ( .A1(n6370), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6015) );
  INV_X1 U7571 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6017) );
  NAND2_X1 U7572 ( .A1(n6056), .A2(n6017), .ZN(n6018) );
  NAND2_X1 U7573 ( .A1(n6019), .A2(n6018), .ZN(n9269) );
  INV_X1 U7574 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n6022) );
  NAND2_X1 U7575 ( .A1(n4404), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6021) );
  NAND2_X1 U7576 ( .A1(n6366), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6020) );
  OAI211_X1 U7577 ( .C1(n6347), .C2(n6022), .A(n6021), .B(n6020), .ZN(n6023)
         );
  INV_X1 U7578 ( .A(n6023), .ZN(n6024) );
  INV_X1 U7579 ( .A(n9624), .ZN(n9193) );
  OR2_X1 U7580 ( .A1(n10106), .A2(n9193), .ZN(n9463) );
  NAND2_X1 U7581 ( .A1(n6490), .A2(n9463), .ZN(n6406) );
  INV_X1 U7582 ( .A(n6406), .ZN(n6027) );
  NAND2_X1 U7583 ( .A1(n10100), .A2(n9496), .ZN(n9464) );
  INV_X1 U7584 ( .A(n9464), .ZN(n6026) );
  OAI21_X1 U7585 ( .B1(n6027), .B2(n6026), .A(n9465), .ZN(n6052) );
  NAND2_X1 U7586 ( .A1(n8104), .A2(n6376), .ZN(n6029) );
  NAND2_X1 U7587 ( .A1(n6370), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6028) );
  INV_X1 U7588 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U7589 ( .A1(n6043), .A2(n6031), .ZN(n6032) );
  NAND2_X1 U7590 ( .A1(n9552), .A2(n6299), .ZN(n6037) );
  INV_X1 U7591 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n10178) );
  NAND2_X1 U7592 ( .A1(n6364), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U7593 ( .A1(n4404), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6033) );
  OAI211_X1 U7594 ( .C1(n10178), .C2(n5998), .A(n6034), .B(n6033), .ZN(n6035)
         );
  INV_X1 U7595 ( .A(n6035), .ZN(n6036) );
  NOR2_X1 U7596 ( .A1(n9561), .A2(n10066), .ZN(n6500) );
  NAND2_X1 U7597 ( .A1(n8098), .A2(n6376), .ZN(n6039) );
  NAND2_X1 U7598 ( .A1(n6370), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6038) );
  INV_X1 U7599 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6040) );
  NAND2_X1 U7600 ( .A1(n6041), .A2(n6040), .ZN(n6042) );
  NAND2_X1 U7601 ( .A1(n6043), .A2(n6042), .ZN(n9567) );
  INV_X1 U7602 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9986) );
  NAND2_X1 U7603 ( .A1(n6364), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6045) );
  NAND2_X1 U7604 ( .A1(n6366), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6044) );
  OAI211_X1 U7605 ( .C1(n6046), .C2(n9986), .A(n6045), .B(n6044), .ZN(n6047)
         );
  INV_X1 U7606 ( .A(n6047), .ZN(n6048) );
  OR2_X1 U7607 ( .A1(n9574), .A2(n9499), .ZN(n6497) );
  INV_X1 U7608 ( .A(n6497), .ZN(n6050) );
  NOR2_X1 U7609 ( .A1(n6500), .A2(n6050), .ZN(n6504) );
  INV_X1 U7610 ( .A(n6504), .ZN(n6051) );
  AOI21_X1 U7611 ( .B1(n6494), .B2(n6052), .A(n6051), .ZN(n6336) );
  NAND2_X1 U7612 ( .A1(n7762), .A2(n6376), .ZN(n6054) );
  NAND2_X1 U7613 ( .A1(n6370), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U7614 ( .A1(n6065), .A2(n9190), .ZN(n6055) );
  AND2_X1 U7615 ( .A1(n6056), .A2(n6055), .ZN(n9630) );
  NAND2_X1 U7616 ( .A1(n9630), .A2(n6299), .ZN(n6061) );
  INV_X1 U7617 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n10189) );
  NAND2_X1 U7618 ( .A1(n6364), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6058) );
  NAND2_X1 U7619 ( .A1(n4404), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6057) );
  OAI211_X1 U7620 ( .C1(n5998), .C2(n10189), .A(n6058), .B(n6057), .ZN(n6059)
         );
  INV_X1 U7621 ( .A(n6059), .ZN(n6060) );
  INV_X1 U7622 ( .A(n9641), .ZN(n9491) );
  OR2_X1 U7623 ( .A1(n9629), .A2(n9491), .ZN(n6484) );
  NAND2_X1 U7624 ( .A1(n7730), .A2(n6376), .ZN(n6063) );
  NAND2_X1 U7625 ( .A1(n6370), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U7626 ( .A1(n6325), .A2(n9249), .ZN(n6064) );
  NAND2_X1 U7627 ( .A1(n6065), .A2(n6064), .ZN(n9645) );
  OR2_X1 U7628 ( .A1(n9645), .A2(n6355), .ZN(n6071) );
  INV_X1 U7629 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U7630 ( .A1(n4404), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6067) );
  NAND2_X1 U7631 ( .A1(n6366), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6066) );
  OAI211_X1 U7632 ( .C1(n6347), .C2(n6068), .A(n6067), .B(n6066), .ZN(n6069)
         );
  INV_X1 U7633 ( .A(n6069), .ZN(n6070) );
  NAND2_X1 U7634 ( .A1(n6071), .A2(n6070), .ZN(n10120) );
  INV_X1 U7635 ( .A(n10120), .ZN(n9661) );
  OR2_X1 U7636 ( .A1(n10116), .A2(n9661), .ZN(n9619) );
  AND2_X1 U7637 ( .A1(n6484), .A2(n9619), .ZN(n9457) );
  NAND2_X1 U7638 ( .A1(n8110), .A2(n6376), .ZN(n6073) );
  NAND2_X1 U7639 ( .A1(n6370), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6072) );
  XNOR2_X1 U7640 ( .A(n6341), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9540) );
  NAND2_X1 U7641 ( .A1(n9540), .A2(n6299), .ZN(n6078) );
  INV_X1 U7642 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n10074) );
  NAND2_X1 U7643 ( .A1(n4404), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U7644 ( .A1(n6366), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6074) );
  OAI211_X1 U7645 ( .C1(n6347), .C2(n10074), .A(n6075), .B(n6074), .ZN(n6076)
         );
  INV_X1 U7646 ( .A(n6076), .ZN(n6077) );
  AND3_X1 U7647 ( .A1(n6336), .A2(n9457), .A3(n6508), .ZN(n6566) );
  NAND2_X1 U7648 ( .A1(n6115), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6083) );
  INV_X1 U7649 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6079) );
  NAND2_X1 U7650 ( .A1(n6095), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6081) );
  NAND2_X1 U7651 ( .A1(n6970), .A2(n4901), .ZN(n6094) );
  NAND2_X1 U7652 ( .A1(n6095), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6087) );
  NAND2_X1 U7653 ( .A1(n6115), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7654 ( .A1(n6114), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6085) );
  INV_X1 U7655 ( .A(n9321), .ZN(n6093) );
  NAND2_X1 U7656 ( .A1(n5553), .A2(SI_0_), .ZN(n6090) );
  INV_X1 U7657 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6089) );
  NAND2_X1 U7658 ( .A1(n6090), .A2(n6089), .ZN(n6092) );
  AND2_X1 U7659 ( .A1(n6092), .A2(n6091), .ZN(n10227) );
  MUX2_X1 U7660 ( .A(n10226), .B(n10227), .S(n6641), .Z(n6928) );
  OR2_X2 U7661 ( .A1(n6926), .A2(n6933), .ZN(n6931) );
  NAND2_X1 U7662 ( .A1(n6095), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6104) );
  NAND2_X1 U7663 ( .A1(n6115), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6103) );
  INV_X1 U7664 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6096) );
  INV_X1 U7665 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6098) );
  NOR2_X1 U7666 ( .A1(n6101), .A2(n6100), .ZN(n6102) );
  NAND2_X1 U7667 ( .A1(n6120), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n6112) );
  INV_X2 U7668 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10213) );
  NOR2_X1 U7669 ( .A1(n6105), .A2(n10213), .ZN(n6106) );
  MUX2_X1 U7670 ( .A(n10213), .B(n6106), .S(P1_IR_REG_2__SCAN_IN), .Z(n6108)
         );
  NOR2_X1 U7671 ( .A1(n6108), .A2(n6123), .ZN(n9337) );
  INV_X1 U7672 ( .A(n6110), .ZN(n6111) );
  NAND2_X1 U7673 ( .A1(n7010), .A2(n6388), .ZN(n6113) );
  INV_X1 U7674 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7042) );
  NAND2_X1 U7675 ( .A1(n6114), .A2(n7042), .ZN(n6119) );
  NAND2_X1 U7676 ( .A1(n6115), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6117) );
  NAND2_X1 U7677 ( .A1(n4404), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6116) );
  NAND2_X1 U7678 ( .A1(n6120), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n6126) );
  NOR2_X1 U7679 ( .A1(n6123), .A2(n10213), .ZN(n6121) );
  MUX2_X1 U7680 ( .A(n10213), .B(n6121), .S(P1_IR_REG_3__SCAN_IN), .Z(n6124)
         );
  AND2_X1 U7681 ( .A1(n6123), .A2(n6122), .ZN(n6134) );
  NOR2_X1 U7682 ( .A1(n6124), .A2(n6134), .ZN(n9351) );
  NAND2_X1 U7683 ( .A1(n6319), .A2(n9351), .ZN(n6125) );
  NAND2_X1 U7684 ( .A1(n9319), .A2(n7045), .ZN(n6536) );
  NAND2_X1 U7685 ( .A1(n6364), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6132) );
  INV_X1 U7686 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n6128) );
  XNOR2_X1 U7687 ( .A(n6128), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n7104) );
  NAND2_X1 U7688 ( .A1(n6299), .A2(n7104), .ZN(n6131) );
  NAND2_X1 U7689 ( .A1(n6366), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6130) );
  NAND2_X1 U7690 ( .A1(n4404), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6129) );
  INV_X1 U7691 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6635) );
  OR2_X1 U7692 ( .A1(n6133), .A2(n6634), .ZN(n6137) );
  INV_X1 U7693 ( .A(n6134), .ZN(n6147) );
  NAND2_X1 U7694 ( .A1(n6147), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6135) );
  XNOR2_X1 U7695 ( .A(n6135), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6861) );
  NAND2_X1 U7696 ( .A1(n6319), .A2(n6861), .ZN(n6136) );
  INV_X1 U7697 ( .A(n7106), .ZN(n10275) );
  NAND2_X1 U7698 ( .A1(n9318), .A2(n10275), .ZN(n6537) );
  NAND2_X1 U7699 ( .A1(n6994), .A2(n6537), .ZN(n6139) );
  NAND2_X1 U7700 ( .A1(n6139), .A2(n6417), .ZN(n7083) );
  NAND2_X1 U7701 ( .A1(n6364), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6146) );
  INV_X1 U7702 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6141) );
  NAND2_X1 U7703 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6140) );
  NAND2_X1 U7704 ( .A1(n6141), .A2(n6140), .ZN(n6142) );
  AND2_X1 U7705 ( .A1(n6152), .A2(n6142), .ZN(n7113) );
  NAND2_X1 U7706 ( .A1(n6299), .A2(n7113), .ZN(n6145) );
  NAND2_X1 U7707 ( .A1(n4404), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6144) );
  NAND2_X1 U7708 ( .A1(n6366), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6143) );
  NAND4_X1 U7709 ( .A1(n6146), .A2(n6145), .A3(n6144), .A4(n6143), .ZN(n9317)
         );
  NAND2_X1 U7710 ( .A1(n6158), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6148) );
  XNOR2_X1 U7711 ( .A(n6148), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6685) );
  AOI22_X1 U7712 ( .A1(n6370), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6319), .B2(
        n6685), .ZN(n6150) );
  OR2_X1 U7713 ( .A1(n6638), .A2(n6133), .ZN(n6149) );
  NAND2_X1 U7714 ( .A1(n6150), .A2(n6149), .ZN(n7089) );
  NAND2_X1 U7715 ( .A1(n9317), .A2(n7177), .ZN(n6538) );
  INV_X1 U7716 ( .A(n9317), .ZN(n7178) );
  NAND2_X1 U7717 ( .A1(n7178), .A2(n7089), .ZN(n6418) );
  INV_X1 U7718 ( .A(n6418), .ZN(n6151) );
  NAND2_X1 U7719 ( .A1(n6364), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6157) );
  INV_X1 U7720 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6714) );
  NAND2_X1 U7721 ( .A1(n6152), .A2(n6714), .ZN(n6153) );
  AND2_X1 U7722 ( .A1(n6187), .A2(n6153), .ZN(n7238) );
  NAND2_X1 U7723 ( .A1(n6299), .A2(n7238), .ZN(n6156) );
  NAND2_X1 U7724 ( .A1(n4404), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6155) );
  NAND2_X1 U7725 ( .A1(n6366), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6154) );
  NAND4_X1 U7726 ( .A1(n6157), .A2(n6156), .A3(n6155), .A4(n6154), .ZN(n9316)
         );
  INV_X1 U7727 ( .A(n9316), .ZN(n7160) );
  OR2_X1 U7728 ( .A1(n6645), .A2(n6133), .ZN(n6160) );
  OAI21_X1 U7729 ( .B1(n6158), .B2(P1_IR_REG_5__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6181) );
  XNOR2_X1 U7730 ( .A(n6181), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6707) );
  AOI22_X1 U7731 ( .A1(n6370), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6319), .B2(
        n6707), .ZN(n6159) );
  NAND2_X1 U7732 ( .A1(n6160), .A2(n6159), .ZN(n7239) );
  NAND2_X1 U7733 ( .A1(n7160), .A2(n7239), .ZN(n7181) );
  NAND2_X1 U7734 ( .A1(n6782), .A2(n6376), .ZN(n6164) );
  NAND2_X1 U7735 ( .A1(n6381), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6162) );
  XNOR2_X1 U7736 ( .A(n6162), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6912) );
  AOI22_X1 U7737 ( .A1(n6370), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6319), .B2(
        n6912), .ZN(n6163) );
  NAND2_X1 U7738 ( .A1(n6364), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6170) );
  NAND2_X1 U7739 ( .A1(n6176), .A2(n6165), .ZN(n6166) );
  AND2_X1 U7740 ( .A1(n6205), .A2(n6166), .ZN(n7678) );
  NAND2_X1 U7741 ( .A1(n6299), .A2(n7678), .ZN(n6169) );
  NAND2_X1 U7742 ( .A1(n4404), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6168) );
  NAND2_X1 U7743 ( .A1(n6366), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6167) );
  NAND4_X1 U7744 ( .A1(n6170), .A2(n6169), .A3(n6168), .A4(n6167), .ZN(n9313)
         );
  INV_X1 U7745 ( .A(n9313), .ZN(n8132) );
  OR2_X1 U7746 ( .A1(n6683), .A2(n6133), .ZN(n6174) );
  OR2_X1 U7747 ( .A1(n6171), .A2(n10213), .ZN(n6172) );
  XNOR2_X1 U7748 ( .A(n6172), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6881) );
  AOI22_X1 U7749 ( .A1(n6370), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6319), .B2(
        n6881), .ZN(n6173) );
  NAND2_X1 U7750 ( .A1(n6364), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6180) );
  INV_X1 U7751 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n9804) );
  NAND2_X1 U7752 ( .A1(n6189), .A2(n9804), .ZN(n6175) );
  AND2_X1 U7753 ( .A1(n6176), .A2(n6175), .ZN(n7572) );
  NAND2_X1 U7754 ( .A1(n6299), .A2(n7572), .ZN(n6179) );
  NAND2_X1 U7755 ( .A1(n4404), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6178) );
  NAND2_X1 U7756 ( .A1(n6366), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6177) );
  NAND2_X1 U7757 ( .A1(n7578), .A2(n7397), .ZN(n7330) );
  OR2_X1 U7758 ( .A1(n6652), .A2(n6133), .ZN(n6185) );
  NAND2_X1 U7759 ( .A1(n6181), .A2(n4570), .ZN(n6182) );
  NAND2_X1 U7760 ( .A1(n6182), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6183) );
  XNOR2_X1 U7761 ( .A(n6183), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6766) );
  AOI22_X1 U7762 ( .A1(n6370), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6319), .B2(
        n6766), .ZN(n6184) );
  NAND2_X1 U7763 ( .A1(n6185), .A2(n6184), .ZN(n7326) );
  NAND2_X1 U7764 ( .A1(n6364), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6193) );
  INV_X1 U7765 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6186) );
  NAND2_X1 U7766 ( .A1(n6187), .A2(n6186), .ZN(n6188) );
  AND2_X1 U7767 ( .A1(n6189), .A2(n6188), .ZN(n7170) );
  NAND2_X1 U7768 ( .A1(n6299), .A2(n7170), .ZN(n6192) );
  NAND2_X1 U7769 ( .A1(n6366), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6191) );
  NAND2_X1 U7770 ( .A1(n4404), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6190) );
  NAND4_X1 U7771 ( .A1(n6193), .A2(n6192), .A3(n6191), .A4(n6190), .ZN(n9315)
         );
  INV_X1 U7772 ( .A(n9315), .ZN(n7576) );
  NAND2_X1 U7773 ( .A1(n7326), .A2(n7576), .ZN(n7335) );
  NAND3_X1 U7774 ( .A1(n7165), .A2(n6434), .A3(n7335), .ZN(n6199) );
  INV_X1 U7775 ( .A(n6434), .ZN(n6194) );
  INV_X1 U7776 ( .A(n7335), .ZN(n7332) );
  OR2_X1 U7777 ( .A1(n6194), .A2(n7332), .ZN(n6196) );
  OR2_X1 U7778 ( .A1(n7664), .A2(n8132), .ZN(n7389) );
  OR2_X1 U7779 ( .A1(n7578), .A2(n7397), .ZN(n7390) );
  NAND2_X1 U7780 ( .A1(n7389), .A2(n7390), .ZN(n6432) );
  NAND2_X1 U7781 ( .A1(n6432), .A2(n7388), .ZN(n6195) );
  OR2_X1 U7782 ( .A1(n7576), .A2(n7326), .ZN(n6426) );
  NAND2_X1 U7783 ( .A1(n7183), .A2(n9316), .ZN(n7182) );
  NAND2_X1 U7784 ( .A1(n6426), .A2(n7182), .ZN(n6197) );
  OR2_X1 U7785 ( .A1(n6432), .A2(n6197), .ZN(n6542) );
  NAND2_X1 U7786 ( .A1(n6541), .A2(n6542), .ZN(n6198) );
  NAND2_X1 U7787 ( .A1(n6199), .A2(n6198), .ZN(n7500) );
  INV_X1 U7788 ( .A(n7500), .ZN(n6212) );
  NAND2_X1 U7789 ( .A1(n6801), .A2(n6376), .ZN(n6204) );
  NAND2_X1 U7790 ( .A1(n6228), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6201) );
  INV_X1 U7791 ( .A(n6201), .ZN(n6200) );
  NAND2_X1 U7792 ( .A1(n6200), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6202) );
  INV_X1 U7793 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6226) );
  NAND2_X1 U7794 ( .A1(n6201), .A2(n6226), .ZN(n6213) );
  AOI22_X1 U7795 ( .A1(n6370), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6319), .B2(
        n7026), .ZN(n6203) );
  NAND2_X1 U7796 ( .A1(n6364), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6210) );
  NAND2_X1 U7797 ( .A1(n6205), .A2(n6920), .ZN(n6206) );
  AND2_X1 U7798 ( .A1(n6218), .A2(n6206), .ZN(n8128) );
  NAND2_X1 U7799 ( .A1(n6299), .A2(n8128), .ZN(n6209) );
  NAND2_X1 U7800 ( .A1(n4404), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6208) );
  NAND2_X1 U7801 ( .A1(n6366), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6207) );
  NAND4_X1 U7802 ( .A1(n6210), .A2(n6209), .A3(n6208), .A4(n6207), .ZN(n9312)
         );
  OR2_X1 U7803 ( .A1(n8134), .A2(n8040), .ZN(n6449) );
  NAND2_X1 U7804 ( .A1(n8134), .A2(n8040), .ZN(n6452) );
  NAND2_X1 U7805 ( .A1(n6449), .A2(n6452), .ZN(n7501) );
  INV_X1 U7806 ( .A(n7501), .ZN(n6211) );
  NAND2_X1 U7807 ( .A1(n6827), .A2(n6376), .ZN(n6216) );
  NAND2_X1 U7808 ( .A1(n6213), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6214) );
  XNOR2_X1 U7809 ( .A(n6214), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7263) );
  AOI22_X1 U7810 ( .A1(n6370), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6319), .B2(
        n7263), .ZN(n6215) );
  NAND2_X1 U7811 ( .A1(n6364), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6223) );
  INV_X1 U7812 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6217) );
  NAND2_X1 U7813 ( .A1(n6218), .A2(n6217), .ZN(n6219) );
  AND2_X1 U7814 ( .A1(n6234), .A2(n6219), .ZN(n8042) );
  NAND2_X1 U7815 ( .A1(n6299), .A2(n8042), .ZN(n6222) );
  NAND2_X1 U7816 ( .A1(n6366), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6221) );
  NAND2_X1 U7817 ( .A1(n4404), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6220) );
  NAND4_X1 U7818 ( .A1(n6223), .A2(n6222), .A3(n6221), .A4(n6220), .ZN(n9311)
         );
  INV_X1 U7819 ( .A(n9311), .ZN(n9202) );
  AND2_X1 U7820 ( .A1(n8028), .A2(n9202), .ZN(n6453) );
  INV_X1 U7821 ( .A(n6453), .ZN(n6224) );
  OR2_X1 U7822 ( .A1(n8028), .A2(n9202), .ZN(n6448) );
  NAND2_X1 U7823 ( .A1(n6889), .A2(n6376), .ZN(n6233) );
  INV_X1 U7824 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n6225) );
  NAND2_X1 U7825 ( .A1(n6226), .A2(n6225), .ZN(n6227) );
  NOR2_X1 U7826 ( .A1(n6230), .A2(n10213), .ZN(n6229) );
  MUX2_X1 U7827 ( .A(n10213), .B(n6229), .S(P1_IR_REG_12__SCAN_IN), .Z(n6231)
         );
  INV_X1 U7828 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n10014) );
  AOI22_X1 U7829 ( .A1(n6370), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6319), .B2(
        n7475), .ZN(n6232) );
  NAND2_X1 U7830 ( .A1(n6364), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6239) );
  INV_X1 U7831 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7256) );
  NAND2_X1 U7832 ( .A1(n6234), .A2(n7256), .ZN(n6235) );
  AND2_X1 U7833 ( .A1(n6243), .A2(n6235), .ZN(n9204) );
  NAND2_X1 U7834 ( .A1(n6299), .A2(n9204), .ZN(n6238) );
  NAND2_X1 U7835 ( .A1(n4404), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6237) );
  NAND2_X1 U7836 ( .A1(n6366), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6236) );
  NAND4_X1 U7837 ( .A1(n6239), .A2(n6238), .A3(n6237), .A4(n6236), .ZN(n10154)
         );
  OR2_X1 U7838 ( .A1(n9000), .A2(n9261), .ZN(n7999) );
  NAND2_X1 U7839 ( .A1(n9000), .A2(n9261), .ZN(n6454) );
  NAND2_X1 U7840 ( .A1(n6951), .A2(n6376), .ZN(n6242) );
  OR2_X1 U7841 ( .A1(n6253), .A2(n10213), .ZN(n6240) );
  XNOR2_X1 U7842 ( .A(n6240), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7584) );
  AOI22_X1 U7843 ( .A1(n6370), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6319), .B2(
        n7584), .ZN(n6241) );
  NAND2_X1 U7844 ( .A1(n6364), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6248) );
  NAND2_X1 U7845 ( .A1(n6243), .A2(n10016), .ZN(n6244) );
  AND2_X1 U7846 ( .A1(n6256), .A2(n6244), .ZN(n9263) );
  NAND2_X1 U7847 ( .A1(n6299), .A2(n9263), .ZN(n6247) );
  NAND2_X1 U7848 ( .A1(n6366), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6246) );
  NAND2_X1 U7849 ( .A1(n4404), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6245) );
  NAND4_X1 U7850 ( .A1(n6248), .A2(n6247), .A3(n6246), .A4(n6245), .ZN(n9742)
         );
  OR2_X1 U7851 ( .A1(n9012), .A2(n9473), .ZN(n6457) );
  NAND2_X1 U7852 ( .A1(n9012), .A2(n9473), .ZN(n6545) );
  INV_X1 U7853 ( .A(n8007), .ZN(n6250) );
  INV_X1 U7854 ( .A(n7999), .ZN(n6249) );
  NOR2_X1 U7855 ( .A1(n6250), .A2(n6249), .ZN(n6251) );
  NAND2_X1 U7856 ( .A1(n7079), .A2(n6376), .ZN(n6255) );
  NAND2_X1 U7857 ( .A1(n6253), .A2(n6252), .ZN(n6277) );
  NAND2_X1 U7858 ( .A1(n6277), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6263) );
  XNOR2_X1 U7859 ( .A(n6263), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7846) );
  AOI22_X1 U7860 ( .A1(n6370), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6319), .B2(
        n7846), .ZN(n6254) );
  NAND2_X1 U7861 ( .A1(n6364), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6261) );
  INV_X1 U7862 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9936) );
  NAND2_X1 U7863 ( .A1(n6256), .A2(n9936), .ZN(n6257) );
  AND2_X1 U7864 ( .A1(n6268), .A2(n6257), .ZN(n9749) );
  NAND2_X1 U7865 ( .A1(n6299), .A2(n9749), .ZN(n6260) );
  NAND2_X1 U7866 ( .A1(n4404), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6259) );
  NAND2_X1 U7867 ( .A1(n6366), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6258) );
  NAND4_X1 U7868 ( .A1(n6261), .A2(n6260), .A3(n6259), .A4(n6258), .ZN(n10153)
         );
  NAND2_X1 U7869 ( .A1(n9752), .A2(n10244), .ZN(n6443) );
  NAND2_X1 U7870 ( .A1(n6550), .A2(n6443), .ZN(n9738) );
  NAND2_X1 U7871 ( .A1(n7145), .A2(n6376), .ZN(n6267) );
  INV_X1 U7872 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6275) );
  NAND2_X1 U7873 ( .A1(n6263), .A2(n6275), .ZN(n6264) );
  NAND2_X1 U7874 ( .A1(n6264), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6265) );
  XNOR2_X1 U7875 ( .A(n6265), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9362) );
  AOI22_X1 U7876 ( .A1(n6370), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6319), .B2(
        n9362), .ZN(n6266) );
  NAND2_X1 U7877 ( .A1(n6364), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6273) );
  NAND2_X1 U7878 ( .A1(n6268), .A2(n7854), .ZN(n6269) );
  AND2_X1 U7879 ( .A1(n6282), .A2(n6269), .ZN(n9727) );
  NAND2_X1 U7880 ( .A1(n6299), .A2(n9727), .ZN(n6272) );
  NAND2_X1 U7881 ( .A1(n4404), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6271) );
  NAND2_X1 U7882 ( .A1(n6366), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6270) );
  NAND4_X1 U7883 ( .A1(n6273), .A2(n6272), .A3(n6271), .A4(n6270), .ZN(n10144)
         );
  INV_X1 U7884 ( .A(n10144), .ZN(n6446) );
  XNOR2_X1 U7885 ( .A(n10247), .B(n6446), .ZN(n9720) );
  NAND2_X1 U7886 ( .A1(n10247), .A2(n6446), .ZN(n6462) );
  NAND2_X1 U7887 ( .A1(n7147), .A2(n6376), .ZN(n6280) );
  INV_X1 U7888 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6274) );
  NAND2_X1 U7889 ( .A1(n6275), .A2(n6274), .ZN(n6276) );
  OAI21_X1 U7890 ( .B1(n6277), .B2(n6276), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6278) );
  XNOR2_X1 U7891 ( .A(n6278), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9391) );
  AOI22_X1 U7892 ( .A1(n6370), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6319), .B2(
        n9391), .ZN(n6279) );
  NAND2_X1 U7893 ( .A1(n6364), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6287) );
  INV_X1 U7894 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6281) );
  NAND2_X1 U7895 ( .A1(n6282), .A2(n6281), .ZN(n6283) );
  AND2_X1 U7896 ( .A1(n6297), .A2(n6283), .ZN(n9705) );
  NAND2_X1 U7897 ( .A1(n6299), .A2(n9705), .ZN(n6286) );
  NAND2_X1 U7898 ( .A1(n4404), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6285) );
  NAND2_X1 U7899 ( .A1(n6366), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6284) );
  NAND4_X1 U7900 ( .A1(n6287), .A2(n6286), .A3(n6285), .A4(n6284), .ZN(n9690)
         );
  OR2_X1 U7901 ( .A1(n9713), .A2(n10242), .ZN(n6464) );
  NAND2_X1 U7902 ( .A1(n9713), .A2(n10242), .ZN(n6559) );
  NAND2_X1 U7903 ( .A1(n7229), .A2(n6376), .ZN(n6295) );
  NOR2_X1 U7904 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n6291) );
  NOR2_X1 U7905 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n6290) );
  NAND2_X1 U7906 ( .A1(n6383), .A2(n5023), .ZN(n6293) );
  XNOR2_X1 U7907 ( .A(n6305), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9401) );
  AOI22_X1 U7908 ( .A1(n6370), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6319), .B2(
        n9401), .ZN(n6294) );
  NAND2_X1 U7909 ( .A1(n6297), .A2(n6296), .ZN(n6298) );
  AND2_X1 U7910 ( .A1(n6308), .A2(n6298), .ZN(n9696) );
  NAND2_X1 U7911 ( .A1(n9696), .A2(n6299), .ZN(n6303) );
  NAND2_X1 U7912 ( .A1(n6364), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6302) );
  NAND2_X1 U7913 ( .A1(n4404), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6301) );
  NAND2_X1 U7914 ( .A1(n6366), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6300) );
  NAND4_X1 U7915 ( .A1(n6303), .A2(n6302), .A3(n6301), .A4(n6300), .ZN(n10143)
         );
  OR2_X1 U7916 ( .A1(n9695), .A2(n9708), .ZN(n6480) );
  NAND2_X1 U7917 ( .A1(n9695), .A2(n9708), .ZN(n6471) );
  NAND2_X1 U7918 ( .A1(n6480), .A2(n6471), .ZN(n9686) );
  NAND2_X1 U7919 ( .A1(n7355), .A2(n6376), .ZN(n6307) );
  XNOR2_X1 U7920 ( .A(n6315), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9429) );
  AOI22_X1 U7921 ( .A1(n6370), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6319), .B2(
        n9429), .ZN(n6306) );
  INV_X1 U7922 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10195) );
  INV_X1 U7923 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9934) );
  NAND2_X1 U7924 ( .A1(n6308), .A2(n9934), .ZN(n6309) );
  NAND2_X1 U7925 ( .A1(n6323), .A2(n6309), .ZN(n9674) );
  OR2_X1 U7926 ( .A1(n9674), .A2(n6355), .ZN(n6313) );
  NAND2_X1 U7927 ( .A1(n6364), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6311) );
  NAND2_X1 U7928 ( .A1(n4404), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6310) );
  AND2_X1 U7929 ( .A1(n6311), .A2(n6310), .ZN(n6312) );
  OAI211_X1 U7930 ( .C1(n5998), .C2(n10195), .A(n6313), .B(n6312), .ZN(n10119)
         );
  INV_X1 U7931 ( .A(n10119), .ZN(n9483) );
  OR2_X1 U7932 ( .A1(n9682), .A2(n9483), .ZN(n6562) );
  NAND2_X1 U7933 ( .A1(n9682), .A2(n9483), .ZN(n6481) );
  NAND2_X1 U7934 ( .A1(n9668), .A2(n6481), .ZN(n9654) );
  NAND2_X1 U7935 ( .A1(n7531), .A2(n6376), .ZN(n6321) );
  AOI22_X1 U7936 ( .A1(n6370), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n6319), .B2(
        n7002), .ZN(n6320) );
  INV_X1 U7937 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n6328) );
  INV_X1 U7938 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6322) );
  NAND2_X1 U7939 ( .A1(n6323), .A2(n6322), .ZN(n6324) );
  NAND2_X1 U7940 ( .A1(n6325), .A2(n6324), .ZN(n9657) );
  OR2_X1 U7941 ( .A1(n9657), .A2(n6355), .ZN(n6327) );
  AOI22_X1 U7942 ( .A1(n6364), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n4404), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n6326) );
  OAI211_X1 U7943 ( .C1(n5998), .C2(n6328), .A(n6327), .B(n6326), .ZN(n10130)
         );
  INV_X1 U7944 ( .A(n10130), .ZN(n9678) );
  OR2_X1 U7945 ( .A1(n9663), .A2(n9678), .ZN(n6563) );
  NAND2_X1 U7946 ( .A1(n9663), .A2(n9678), .ZN(n6569) );
  NAND2_X1 U7947 ( .A1(n9654), .A2(n9653), .ZN(n6329) );
  INV_X1 U7948 ( .A(n6508), .ZN(n6351) );
  AND2_X1 U7949 ( .A1(n9561), .A2(n10066), .ZN(n9467) );
  INV_X1 U7950 ( .A(n9467), .ZN(n6330) );
  NOR2_X1 U7951 ( .A1(n6351), .A2(n6330), .ZN(n6570) );
  NAND2_X1 U7952 ( .A1(n10106), .A2(n9193), .ZN(n6387) );
  NAND2_X1 U7953 ( .A1(n9464), .A2(n6387), .ZN(n6407) );
  INV_X1 U7954 ( .A(n6407), .ZN(n6332) );
  NAND2_X1 U7955 ( .A1(n9629), .A2(n9491), .ZN(n6487) );
  NAND2_X1 U7956 ( .A1(n10116), .A2(n9661), .ZN(n6473) );
  NAND2_X1 U7957 ( .A1(n6487), .A2(n6473), .ZN(n6331) );
  NAND2_X1 U7958 ( .A1(n6331), .A2(n6484), .ZN(n9459) );
  NAND3_X1 U7959 ( .A1(n6494), .A2(n6332), .A3(n9459), .ZN(n6335) );
  INV_X1 U7960 ( .A(n6500), .ZN(n6334) );
  NAND2_X1 U7961 ( .A1(n9574), .A2(n9499), .ZN(n9466) );
  INV_X1 U7962 ( .A(n9466), .ZN(n6333) );
  AND2_X1 U7963 ( .A1(n6334), .A2(n6333), .ZN(n6502) );
  AOI21_X1 U7964 ( .B1(n6336), .B2(n6335), .A(n6502), .ZN(n6352) );
  NAND2_X1 U7965 ( .A1(n8113), .A2(n6376), .ZN(n6338) );
  NAND2_X1 U7966 ( .A1(n6370), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6337) );
  INV_X1 U7967 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6340) );
  INV_X1 U7968 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6339) );
  OAI21_X1 U7969 ( .B1(n6341), .B2(n6340), .A(n6339), .ZN(n6344) );
  INV_X1 U7970 ( .A(n6341), .ZN(n6343) );
  AND2_X1 U7971 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n6342) );
  NAND2_X1 U7972 ( .A1(n6343), .A2(n6342), .ZN(n9510) );
  NAND2_X1 U7973 ( .A1(n6344), .A2(n9510), .ZN(n9176) );
  INV_X1 U7974 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n10064) );
  NAND2_X1 U7975 ( .A1(n4404), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6346) );
  NAND2_X1 U7976 ( .A1(n6366), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6345) );
  OAI211_X1 U7977 ( .C1(n6347), .C2(n10064), .A(n6346), .B(n6345), .ZN(n6348)
         );
  INV_X1 U7978 ( .A(n6348), .ZN(n6349) );
  NAND2_X1 U7979 ( .A1(n9532), .A2(n10067), .ZN(n9470) );
  NAND2_X1 U7980 ( .A1(n9545), .A2(n9555), .ZN(n9468) );
  NAND2_X1 U7981 ( .A1(n9470), .A2(n9468), .ZN(n6514) );
  INV_X1 U7982 ( .A(n6514), .ZN(n6512) );
  OAI21_X1 U7983 ( .B1(n6352), .B2(n6351), .A(n6512), .ZN(n6572) );
  AOI211_X1 U7984 ( .C1(n6566), .C2(n9458), .A(n6570), .B(n6572), .ZN(n6374)
         );
  NAND2_X1 U7985 ( .A1(n8986), .A2(n6376), .ZN(n6354) );
  NAND2_X1 U7986 ( .A1(n6370), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6353) );
  OR2_X1 U7987 ( .A1(n9510), .A2(n6355), .ZN(n6360) );
  NAND2_X1 U7988 ( .A1(n6364), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6358) );
  NAND2_X1 U7989 ( .A1(n4404), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6357) );
  NAND2_X1 U7990 ( .A1(n6366), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6356) );
  AND3_X1 U7991 ( .A1(n6358), .A2(n6357), .A3(n6356), .ZN(n6359) );
  NAND2_X1 U7992 ( .A1(n6403), .A2(n6509), .ZN(n6576) );
  NAND2_X1 U7993 ( .A1(n6364), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6363) );
  NAND2_X1 U7994 ( .A1(n4404), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6362) );
  NAND2_X1 U7995 ( .A1(n6366), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6361) );
  NAND3_X1 U7996 ( .A1(n6363), .A2(n6362), .A3(n6361), .ZN(n9449) );
  INV_X1 U7997 ( .A(n9449), .ZN(n6380) );
  NAND2_X1 U7998 ( .A1(n6364), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6369) );
  NAND2_X1 U7999 ( .A1(n4404), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6368) );
  NAND2_X1 U8000 ( .A1(n6366), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6367) );
  NAND3_X1 U8001 ( .A1(n6369), .A2(n6368), .A3(n6367), .ZN(n9509) );
  INV_X1 U8002 ( .A(n9509), .ZN(n6375) );
  OAI21_X1 U8003 ( .B1(n6380), .B2(n6375), .A(n6386), .ZN(n6520) );
  NAND2_X1 U8004 ( .A1(n10052), .A2(n9528), .ZN(n6575) );
  NAND2_X1 U8005 ( .A1(n6520), .A2(n6575), .ZN(n6405) );
  INV_X1 U8006 ( .A(n6405), .ZN(n6373) );
  OAI21_X1 U8007 ( .B1(n6374), .B2(n6576), .A(n6373), .ZN(n6379) );
  NOR2_X1 U8008 ( .A1(n6386), .A2(n6375), .ZN(n6578) );
  NAND2_X1 U8009 ( .A1(n6370), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n6377) );
  OR2_X1 U8010 ( .A1(n9450), .A2(n6380), .ZN(n6610) );
  INV_X1 U8011 ( .A(n6610), .ZN(n6378) );
  AOI21_X1 U8012 ( .B1(n6379), .B2(n6519), .A(n6378), .ZN(n6402) );
  NAND2_X1 U8013 ( .A1(n9450), .A2(n6380), .ZN(n6580) );
  INV_X1 U8014 ( .A(n6381), .ZN(n6383) );
  NAND2_X1 U8015 ( .A1(n6531), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6385) );
  NAND2_X1 U8016 ( .A1(n6745), .A2(n6607), .ZN(n6746) );
  NAND2_X1 U8017 ( .A1(n6580), .A2(n6934), .ZN(n6401) );
  AND2_X1 U8018 ( .A1(n6610), .A2(n6580), .ZN(n6522) );
  NOR2_X1 U8019 ( .A1(n10168), .A2(n9509), .ZN(n6573) );
  NAND2_X1 U8020 ( .A1(n6497), .A2(n9466), .ZN(n9566) );
  NAND2_X1 U8021 ( .A1(n9463), .A2(n6387), .ZN(n9461) );
  OR2_X1 U8022 ( .A1(n10116), .A2(n10120), .ZN(n9488) );
  NAND2_X1 U8023 ( .A1(n10116), .A2(n10120), .ZN(n9489) );
  NAND2_X1 U8024 ( .A1(n9488), .A2(n9489), .ZN(n9639) );
  INV_X1 U8025 ( .A(n7834), .ZN(n6393) );
  INV_X1 U8026 ( .A(n6928), .ZN(n6389) );
  NAND2_X1 U8027 ( .A1(n9321), .A2(n6389), .ZN(n6534) );
  NAND2_X1 U8028 ( .A1(n6933), .A2(n6534), .ZN(n6814) );
  OR4_X1 U8029 ( .A1(n7014), .A2(n6926), .A3(n6814), .A4(n6607), .ZN(n6390) );
  NAND2_X1 U8030 ( .A1(n6418), .A2(n6538), .ZN(n7086) );
  NOR4_X1 U8031 ( .A1(n6390), .A2(n7086), .A3(n6999), .A4(n6974), .ZN(n6391)
         );
  NAND4_X1 U8032 ( .A1(n6391), .A2(n6434), .A3(n7181), .A4(n7335), .ZN(n6392)
         );
  NOR4_X1 U8033 ( .A1(n6393), .A2(n7501), .A3(n6542), .A4(n6392), .ZN(n6394)
         );
  XNOR2_X1 U8034 ( .A(n8028), .B(n9311), .ZN(n7802) );
  NAND4_X1 U8035 ( .A1(n6262), .A2(n8007), .A3(n6394), .A4(n7802), .ZN(n6395)
         );
  NOR4_X1 U8036 ( .A1(n9703), .A2(n9720), .A3(n9686), .A4(n6395), .ZN(n6396)
         );
  AND4_X1 U8037 ( .A1(n9639), .A2(n9653), .A3(n9671), .A4(n6396), .ZN(n6397)
         );
  XNOR2_X1 U8038 ( .A(n9629), .B(n9641), .ZN(n9620) );
  NAND4_X1 U8039 ( .A1(n9597), .A2(n9462), .A3(n6397), .A4(n9620), .ZN(n6398)
         );
  NOR4_X1 U8040 ( .A1(n9536), .A2(n9566), .A3(n4808), .A4(n6398), .ZN(n6399)
         );
  XNOR2_X1 U8041 ( .A(n9561), .B(n10086), .ZN(n9551) );
  NAND4_X1 U8042 ( .A1(n9505), .A2(n9521), .A3(n6399), .A4(n9551), .ZN(n6400)
         );
  OAI21_X1 U8043 ( .B1(n6402), .B2(n6401), .A(n4471), .ZN(n6527) );
  NAND2_X1 U8044 ( .A1(n6519), .A2(n6403), .ZN(n6404) );
  MUX2_X1 U8045 ( .A(n6405), .B(n6404), .S(n6505), .Z(n6524) );
  MUX2_X1 U8046 ( .A(n6407), .B(n6406), .S(n6790), .Z(n6493) );
  NOR2_X1 U8047 ( .A1(n9459), .A2(n6505), .ZN(n6408) );
  NAND2_X1 U8048 ( .A1(n6537), .A2(n6536), .ZN(n6410) );
  AOI21_X1 U8049 ( .B1(n6409), .B2(n6127), .A(n6410), .ZN(n6414) );
  INV_X1 U8050 ( .A(n6536), .ZN(n6411) );
  OAI211_X1 U8051 ( .C1(n6409), .C2(n6411), .A(n6417), .B(n6127), .ZN(n6412)
         );
  NAND2_X1 U8052 ( .A1(n6412), .A2(n6537), .ZN(n6413) );
  MUX2_X1 U8053 ( .A(n6414), .B(n6413), .S(n6790), .Z(n6421) );
  NAND2_X1 U8054 ( .A1(n6421), .A2(n6418), .ZN(n6416) );
  AND2_X1 U8055 ( .A1(n7182), .A2(n6538), .ZN(n6419) );
  INV_X1 U8056 ( .A(n7181), .ZN(n6415) );
  AOI21_X1 U8057 ( .B1(n6416), .B2(n6419), .A(n6415), .ZN(n6424) );
  NAND2_X1 U8058 ( .A1(n6418), .A2(n6417), .ZN(n6420) );
  OAI21_X1 U8059 ( .B1(n6421), .B2(n6420), .A(n6419), .ZN(n6422) );
  NAND2_X1 U8060 ( .A1(n6422), .A2(n7181), .ZN(n6423) );
  MUX2_X1 U8061 ( .A(n6424), .B(n6423), .S(n6505), .Z(n6425) );
  NAND2_X1 U8062 ( .A1(n6426), .A2(n7335), .ZN(n7185) );
  INV_X1 U8063 ( .A(n7185), .ZN(n7167) );
  NAND2_X1 U8064 ( .A1(n6425), .A2(n7167), .ZN(n6431) );
  NAND2_X1 U8065 ( .A1(n7390), .A2(n6426), .ZN(n6428) );
  NAND2_X1 U8066 ( .A1(n7330), .A2(n7335), .ZN(n6427) );
  MUX2_X1 U8067 ( .A(n6428), .B(n6427), .S(n6505), .Z(n6429) );
  INV_X1 U8068 ( .A(n6429), .ZN(n6430) );
  NAND2_X1 U8069 ( .A1(n6431), .A2(n6430), .ZN(n6436) );
  INV_X1 U8070 ( .A(n6432), .ZN(n6433) );
  MUX2_X1 U8071 ( .A(n6434), .B(n6433), .S(n6505), .Z(n6435) );
  NAND2_X1 U8072 ( .A1(n6436), .A2(n6435), .ZN(n6450) );
  NAND2_X1 U8073 ( .A1(n6450), .A2(n7389), .ZN(n6437) );
  NAND2_X1 U8074 ( .A1(n6437), .A2(n6452), .ZN(n6438) );
  NAND3_X1 U8075 ( .A1(n6438), .A2(n6449), .A3(n6448), .ZN(n6439) );
  NAND3_X1 U8076 ( .A1(n6439), .A2(n6454), .A3(n6224), .ZN(n6440) );
  NAND2_X1 U8077 ( .A1(n6440), .A2(n7999), .ZN(n6442) );
  INV_X1 U8078 ( .A(n6457), .ZN(n6551) );
  OR2_X1 U8079 ( .A1(n9738), .A2(n6551), .ZN(n6441) );
  AOI21_X1 U8080 ( .B1(n6442), .B2(n6545), .A(n6441), .ZN(n6444) );
  NAND2_X1 U8081 ( .A1(n6462), .A2(n6443), .ZN(n6555) );
  OAI21_X1 U8082 ( .B1(n6444), .B2(n6555), .A(n6464), .ZN(n6445) );
  NAND3_X1 U8083 ( .A1(n6445), .A2(n6790), .A3(n6559), .ZN(n6469) );
  OR2_X1 U8084 ( .A1(n10247), .A2(n6446), .ZN(n6460) );
  INV_X1 U8085 ( .A(n6460), .ZN(n6447) );
  AND2_X1 U8086 ( .A1(n6559), .A2(n6447), .ZN(n6468) );
  AND2_X1 U8087 ( .A1(n7999), .A2(n6448), .ZN(n6451) );
  NAND2_X1 U8088 ( .A1(n6451), .A2(n6449), .ZN(n6544) );
  AOI21_X1 U8089 ( .B1(n6450), .B2(n7388), .A(n6544), .ZN(n6458) );
  INV_X1 U8090 ( .A(n6451), .ZN(n6456) );
  NOR2_X1 U8091 ( .A1(n6453), .A2(n4816), .ZN(n6455) );
  OAI21_X1 U8092 ( .B1(n6456), .B2(n6455), .A(n6454), .ZN(n6546) );
  OAI21_X1 U8093 ( .B1(n6458), .B2(n6546), .A(n6457), .ZN(n6459) );
  NAND3_X1 U8094 ( .A1(n6459), .A2(n6262), .A3(n6545), .ZN(n6461) );
  AND2_X1 U8095 ( .A1(n6464), .A2(n6460), .ZN(n6554) );
  NAND3_X1 U8096 ( .A1(n6461), .A2(n6554), .A3(n6550), .ZN(n6466) );
  INV_X1 U8097 ( .A(n6462), .ZN(n6463) );
  NAND2_X1 U8098 ( .A1(n6464), .A2(n6463), .ZN(n6465) );
  NAND3_X1 U8099 ( .A1(n6466), .A2(n6559), .A3(n6465), .ZN(n6467) );
  NAND2_X1 U8100 ( .A1(n6470), .A2(n6304), .ZN(n6483) );
  AND2_X1 U8101 ( .A1(n6481), .A2(n6471), .ZN(n6561) );
  NAND2_X1 U8102 ( .A1(n6483), .A2(n6561), .ZN(n6472) );
  NAND4_X1 U8103 ( .A1(n6472), .A2(n6563), .A3(n6562), .A4(n6505), .ZN(n6478)
         );
  INV_X1 U8104 ( .A(n9663), .ZN(n10123) );
  AOI21_X1 U8105 ( .B1(n6473), .B2(n10123), .A(n6790), .ZN(n6476) );
  NAND2_X1 U8106 ( .A1(n9619), .A2(n6563), .ZN(n6475) );
  NAND3_X1 U8107 ( .A1(n6473), .A2(n10130), .A3(n6505), .ZN(n6474) );
  OAI21_X1 U8108 ( .B1(n6476), .B2(n6475), .A(n6474), .ZN(n6477) );
  NAND2_X1 U8109 ( .A1(n6478), .A2(n6477), .ZN(n6479) );
  OAI21_X1 U8110 ( .B1(n9457), .B2(n6790), .A(n6479), .ZN(n6489) );
  AND2_X1 U8111 ( .A1(n6562), .A2(n6480), .ZN(n6557) );
  NAND2_X1 U8112 ( .A1(n6569), .A2(n6481), .ZN(n6482) );
  AOI21_X1 U8113 ( .B1(n6483), .B2(n6557), .A(n6482), .ZN(n6486) );
  INV_X1 U8114 ( .A(n6484), .ZN(n6485) );
  OAI21_X1 U8115 ( .B1(n6486), .B2(n6485), .A(n6790), .ZN(n6488) );
  MUX2_X1 U8116 ( .A(n6490), .B(n9464), .S(n6790), .Z(n6491) );
  OAI211_X1 U8117 ( .C1(n6493), .C2(n6492), .A(n9579), .B(n6491), .ZN(n6496)
         );
  MUX2_X1 U8118 ( .A(n6494), .B(n9465), .S(n6790), .Z(n6495) );
  NAND2_X1 U8119 ( .A1(n6496), .A2(n6495), .ZN(n6503) );
  INV_X1 U8120 ( .A(n6503), .ZN(n6498) );
  AOI21_X1 U8121 ( .B1(n6498), .B2(n6497), .A(n9467), .ZN(n6501) );
  INV_X1 U8122 ( .A(n6502), .ZN(n6499) );
  OAI21_X1 U8123 ( .B1(n6501), .B2(n6500), .A(n6499), .ZN(n6507) );
  AOI211_X1 U8124 ( .C1(n6504), .C2(n6503), .A(n9467), .B(n6502), .ZN(n6506)
         );
  MUX2_X1 U8125 ( .A(n6507), .B(n6506), .S(n6505), .Z(n6515) );
  OR2_X1 U8126 ( .A1(n6514), .A2(n6508), .ZN(n6510) );
  AND2_X1 U8127 ( .A1(n6510), .A2(n6509), .ZN(n6513) );
  INV_X1 U8128 ( .A(n6513), .ZN(n6511) );
  AOI21_X1 U8129 ( .B1(n6515), .B2(n6512), .A(n6511), .ZN(n6517) );
  OAI21_X1 U8130 ( .B1(n6515), .B2(n6514), .A(n6513), .ZN(n6516) );
  MUX2_X1 U8131 ( .A(n6517), .B(n6516), .S(n6790), .Z(n6518) );
  NOR2_X1 U8132 ( .A1(n6518), .A2(n9472), .ZN(n6523) );
  OAI211_X1 U8133 ( .C1(n6524), .C2(n6523), .A(n6522), .B(n6521), .ZN(n6525)
         );
  OAI21_X1 U8134 ( .B1(n6790), .B2(n6580), .A(n6525), .ZN(n6612) );
  INV_X1 U8135 ( .A(n6607), .ZN(n7767) );
  AOI21_X1 U8136 ( .B1(n6612), .B2(n6745), .A(n7767), .ZN(n6526) );
  INV_X1 U8137 ( .A(n6528), .ZN(n6529) );
  NAND2_X1 U8138 ( .A1(n6529), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6530) );
  MUX2_X1 U8139 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6530), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n6532) );
  INV_X1 U8140 ( .A(n7751), .ZN(n6750) );
  NOR2_X1 U8141 ( .A1(n4408), .A2(n6750), .ZN(n6818) );
  AND4_X1 U8142 ( .A1(n6535), .A2(n6534), .A3(n6533), .A4(n6607), .ZN(n6539)
         );
  NAND4_X1 U8143 ( .A1(n6539), .A2(n6538), .A3(n6537), .A4(n6536), .ZN(n6540)
         );
  AND2_X1 U8144 ( .A1(n7165), .A2(n6540), .ZN(n6543) );
  OAI21_X1 U8145 ( .B1(n6543), .B2(n6542), .A(n6541), .ZN(n6549) );
  INV_X1 U8146 ( .A(n6544), .ZN(n6548) );
  INV_X1 U8147 ( .A(n6545), .ZN(n6547) );
  AOI211_X1 U8148 ( .C1(n6549), .C2(n6548), .A(n6547), .B(n6546), .ZN(n6553)
         );
  INV_X1 U8149 ( .A(n6550), .ZN(n6552) );
  NOR3_X1 U8150 ( .A1(n6553), .A2(n6552), .A3(n6551), .ZN(n6556) );
  OAI21_X1 U8151 ( .B1(n6556), .B2(n6555), .A(n6554), .ZN(n6560) );
  INV_X1 U8152 ( .A(n6557), .ZN(n6558) );
  AOI21_X1 U8153 ( .B1(n6560), .B2(n6559), .A(n6558), .ZN(n6565) );
  INV_X1 U8154 ( .A(n6561), .ZN(n6564) );
  OAI211_X1 U8155 ( .C1(n6565), .C2(n6564), .A(n6563), .B(n6562), .ZN(n6568)
         );
  INV_X1 U8156 ( .A(n6566), .ZN(n6567) );
  AOI21_X1 U8157 ( .B1(n6569), .B2(n6568), .A(n6567), .ZN(n6571) );
  NOR3_X1 U8158 ( .A1(n6572), .A2(n6571), .A3(n6570), .ZN(n6577) );
  INV_X1 U8159 ( .A(n6573), .ZN(n6574) );
  OAI211_X1 U8160 ( .C1(n6577), .C2(n6576), .A(n6575), .B(n6574), .ZN(n6581)
         );
  INV_X1 U8161 ( .A(n6578), .ZN(n6579) );
  NAND3_X1 U8162 ( .A1(n6581), .A2(n6580), .A3(n6579), .ZN(n6582) );
  NAND2_X1 U8163 ( .A1(n6582), .A2(n6610), .ZN(n6589) );
  NAND2_X1 U8164 ( .A1(n6584), .A2(n6583), .ZN(n6585) );
  NAND2_X1 U8165 ( .A1(n6585), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6587) );
  INV_X1 U8166 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6586) );
  INV_X1 U8167 ( .A(n6639), .ZN(n6762) );
  INV_X1 U8168 ( .A(n7915), .ZN(n6642) );
  NAND2_X1 U8169 ( .A1(n4408), .A2(n7751), .ZN(n6721) );
  NOR2_X1 U8170 ( .A1(n6589), .A2(n6721), .ZN(n6588) );
  AOI211_X1 U8171 ( .C1(n6818), .C2(n6589), .A(n6642), .B(n6588), .ZN(n6590)
         );
  OAI21_X1 U8172 ( .B1(n6591), .B2(n7751), .A(n6590), .ZN(n6614) );
  NAND2_X1 U8173 ( .A1(n4432), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6592) );
  MUX2_X1 U8174 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6592), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n6593) );
  NAND2_X1 U8175 ( .A1(n6595), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6596) );
  MUX2_X1 U8176 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6596), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n6597) );
  NAND2_X1 U8177 ( .A1(n6597), .A2(n4432), .ZN(n8100) );
  INV_X1 U8178 ( .A(n6598), .ZN(n6599) );
  NAND2_X1 U8179 ( .A1(n6599), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6600) );
  MUX2_X1 U8180 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6600), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n6601) );
  NAND2_X1 U8181 ( .A1(n6601), .A2(n6595), .ZN(n8060) );
  NOR2_X1 U8182 ( .A1(n8100), .A2(n8060), .ZN(n6602) );
  NAND3_X1 U8183 ( .A1(n6755), .A2(n6639), .A3(P1_STATE_REG_SCAN_IN), .ZN(
        n6798) );
  INV_X1 U8184 ( .A(n6798), .ZN(n6807) );
  NAND2_X1 U8185 ( .A1(n4408), .A2(n6745), .ZN(n6786) );
  INV_X1 U8186 ( .A(n6786), .ZN(n6604) );
  AND2_X1 U8187 ( .A1(n6604), .A2(n6723), .ZN(n6816) );
  NAND2_X1 U8188 ( .A1(n6807), .A2(n6816), .ZN(n6847) );
  INV_X1 U8189 ( .A(n6605), .ZN(n6935) );
  INV_X1 U8190 ( .A(n10223), .ZN(n6663) );
  NAND2_X1 U8191 ( .A1(n6935), .A2(n6663), .ZN(n6660) );
  NOR2_X1 U8192 ( .A1(n6642), .A2(n6745), .ZN(n6609) );
  INV_X1 U8193 ( .A(n6609), .ZN(n6606) );
  OAI211_X1 U8194 ( .C1(n6847), .C2(n6660), .A(P1_B_REG_SCAN_IN), .B(n6606), 
        .ZN(n6613) );
  NAND2_X1 U8195 ( .A1(n6607), .A2(n6750), .ZN(n6791) );
  INV_X1 U8196 ( .A(n6791), .ZN(n6608) );
  OAI211_X1 U8197 ( .C1(n6610), .C2(n4408), .A(n6609), .B(n6608), .ZN(n6611)
         );
  NAND3_X1 U8198 ( .A1(n6614), .A2(n6613), .A3(n5022), .ZN(P1_U3242) );
  NOR2_X1 U8199 ( .A1(n6755), .A2(P1_U3086), .ZN(n6616) );
  AND2_X2 U8200 ( .A1(n6616), .A2(n6639), .ZN(P1_U3973) );
  NAND2_X1 U8201 ( .A1(n7221), .A2(n6617), .ZN(n6618) );
  NAND2_X1 U8202 ( .A1(n6618), .A2(n7219), .ZN(n7200) );
  NAND2_X1 U8203 ( .A1(n7200), .A2(n6619), .ZN(n6620) );
  NAND2_X1 U8204 ( .A1(n6620), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  NOR2_X1 U8205 ( .A1(n5553), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10215) );
  INV_X1 U8206 ( .A(n10215), .ZN(n10225) );
  INV_X1 U8207 ( .A(n9337), .ZN(n6621) );
  OAI222_X1 U8208 ( .A1(n10225), .A2(n6622), .B1(n10222), .B2(n6625), .C1(
        P1_U3086), .C2(n6621), .ZN(P1_U3353) );
  AOI22_X1 U8209 ( .A1(n9351), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n10215), .ZN(n6623) );
  OAI21_X1 U8210 ( .B1(n6627), .B2(n10222), .A(n6623), .ZN(P1_U3352) );
  INV_X2 U8211 ( .A(n8991), .ZN(n8987) );
  NAND2_X1 U8212 ( .A1(n6624), .A2(P2_U3151), .ZN(n8993) );
  OAI222_X1 U8213 ( .A1(n8987), .A2(n6626), .B1(n8993), .B2(n6625), .C1(n10317), .C2(P2_U3151), .ZN(P2_U3293) );
  OAI222_X1 U8214 ( .A1(n8987), .A2(n6628), .B1(n8993), .B2(n6627), .C1(n7416), 
        .C2(P2_U3151), .ZN(P2_U3292) );
  INV_X1 U8215 ( .A(n8993), .ZN(n7924) );
  INV_X1 U8216 ( .A(n7924), .ZN(n7922) );
  OAI222_X1 U8217 ( .A1(n8987), .A2(n6629), .B1(n7922), .B2(n6631), .C1(n7285), 
        .C2(P2_U3151), .ZN(P2_U3294) );
  AOI22_X1 U8218 ( .A1(n10215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(n9324), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6630) );
  OAI21_X1 U8219 ( .B1(n6631), .B2(n10222), .A(n6630), .ZN(P1_U3354) );
  OAI222_X1 U8220 ( .A1(n7444), .A2(P2_U3151), .B1(n8993), .B2(n6634), .C1(
        n6632), .C2(n8987), .ZN(P2_U3291) );
  INV_X1 U8221 ( .A(n6861), .ZN(n6633) );
  OAI222_X1 U8222 ( .A1(n10225), .A2(n6635), .B1(n10222), .B2(n6634), .C1(
        P1_U3086), .C2(n6633), .ZN(P1_U3351) );
  INV_X1 U8223 ( .A(n6685), .ZN(n6691) );
  OAI222_X1 U8224 ( .A1(n10225), .A2(n6636), .B1(n10222), .B2(n6638), .C1(
        P1_U3086), .C2(n6691), .ZN(P1_U3350) );
  OAI222_X1 U8225 ( .A1(n7534), .A2(P2_U3151), .B1(n8993), .B2(n6638), .C1(
        n6637), .C2(n8987), .ZN(P2_U3290) );
  NAND2_X1 U8226 ( .A1(n6934), .A2(n6639), .ZN(n6640) );
  AND2_X1 U8227 ( .A1(n6641), .A2(n6640), .ZN(n6649) );
  INV_X1 U8228 ( .A(n6649), .ZN(n6643) );
  NAND2_X1 U8229 ( .A1(n6642), .A2(n6798), .ZN(n6648) );
  NAND2_X1 U8230 ( .A1(n6643), .A2(n6648), .ZN(n9443) );
  NOR2_X1 U8231 ( .A1(n9420), .A2(P1_U3973), .ZN(P1_U3085) );
  OAI222_X1 U8232 ( .A1(n7687), .A2(P2_U3151), .B1(n8993), .B2(n6645), .C1(
        n6644), .C2(n8987), .ZN(P2_U3289) );
  INV_X1 U8233 ( .A(n6707), .ZN(n6717) );
  OAI222_X1 U8234 ( .A1(n10225), .A2(n6646), .B1(n10222), .B2(n6645), .C1(
        P1_U3086), .C2(n6717), .ZN(P1_U3349) );
  INV_X1 U8235 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6826) );
  AOI21_X1 U8236 ( .B1(n6663), .B2(n6826), .A(n6605), .ZN(n6857) );
  OAI21_X1 U8237 ( .B1(n6663), .B2(P1_REG1_REG_0__SCAN_IN), .A(n6857), .ZN(
        n6647) );
  XOR2_X1 U8238 ( .A(n10226), .B(n6647), .Z(n6651) );
  NAND2_X1 U8239 ( .A1(n6649), .A2(n6648), .ZN(n6664) );
  AOI22_X1 U8240 ( .A1(n9420), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n6650) );
  OAI21_X1 U8241 ( .B1(n6651), .B2(n6664), .A(n6650), .ZN(P1_U3243) );
  OAI222_X1 U8242 ( .A1(n7684), .A2(P2_U3151), .B1(n7922), .B2(n6652), .C1(
        n9977), .C2(n8987), .ZN(P2_U3288) );
  INV_X1 U8243 ( .A(n6766), .ZN(n6771) );
  OAI222_X1 U8244 ( .A1(n10225), .A2(n6653), .B1(n10222), .B2(n6652), .C1(
        P1_U3086), .C2(n6771), .ZN(P1_U3348) );
  XNOR2_X1 U8245 ( .A(n9337), .B(n6096), .ZN(n9342) );
  AND2_X1 U8246 ( .A1(n10226), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9331) );
  NAND2_X1 U8247 ( .A1(n9324), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6654) );
  NAND2_X1 U8248 ( .A1(n9329), .A2(n6654), .ZN(n9341) );
  NAND2_X1 U8249 ( .A1(n9342), .A2(n9341), .ZN(n9340) );
  NAND2_X1 U8250 ( .A1(n9337), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6655) );
  NAND2_X1 U8251 ( .A1(n9340), .A2(n6655), .ZN(n9348) );
  INV_X1 U8252 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6656) );
  XNOR2_X1 U8253 ( .A(n9351), .B(n6656), .ZN(n9349) );
  NAND2_X1 U8254 ( .A1(n9348), .A2(n9349), .ZN(n9347) );
  NAND2_X1 U8255 ( .A1(n9351), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6657) );
  NAND2_X1 U8256 ( .A1(n9347), .A2(n6657), .ZN(n6859) );
  INV_X1 U8257 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6658) );
  XNOR2_X1 U8258 ( .A(n6861), .B(n6658), .ZN(n6860) );
  INV_X1 U8259 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6659) );
  MUX2_X1 U8260 ( .A(n6659), .B(P1_REG2_REG_5__SCAN_IN), .S(n6685), .Z(n6661)
         );
  AOI211_X1 U8261 ( .C1(n6662), .C2(n6661), .A(n6684), .B(n9415), .ZN(n6679)
         );
  INV_X1 U8262 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6665) );
  MUX2_X1 U8263 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6665), .S(n9337), .Z(n9339)
         );
  INV_X1 U8264 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6666) );
  MUX2_X1 U8265 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6666), .S(n9324), .Z(n6667)
         );
  AND2_X1 U8266 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(n10226), .ZN(n9328) );
  NAND2_X1 U8267 ( .A1(n6667), .A2(n9328), .ZN(n9326) );
  NAND2_X1 U8268 ( .A1(n9324), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6668) );
  NAND2_X1 U8269 ( .A1(n9326), .A2(n6668), .ZN(n9338) );
  NAND2_X1 U8270 ( .A1(n9339), .A2(n9338), .ZN(n9353) );
  NAND2_X1 U8271 ( .A1(n9337), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9352) );
  NAND2_X1 U8272 ( .A1(n9353), .A2(n9352), .ZN(n6671) );
  INV_X1 U8273 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6669) );
  MUX2_X1 U8274 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6669), .S(n9351), .Z(n6670)
         );
  NAND2_X1 U8275 ( .A1(n6671), .A2(n6670), .ZN(n9356) );
  NAND2_X1 U8276 ( .A1(n9351), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6863) );
  NAND2_X1 U8277 ( .A1(n9356), .A2(n6863), .ZN(n6674) );
  INV_X1 U8278 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6672) );
  MUX2_X1 U8279 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6672), .S(n6861), .Z(n6673)
         );
  NAND2_X1 U8280 ( .A1(n6674), .A2(n6673), .ZN(n6865) );
  NAND2_X1 U8281 ( .A1(n6861), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6676) );
  INV_X1 U8282 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7093) );
  MUX2_X1 U8283 ( .A(n7093), .B(P1_REG1_REG_5__SCAN_IN), .S(n6685), .Z(n6675)
         );
  AOI21_X1 U8284 ( .B1(n6865), .B2(n6676), .A(n6675), .ZN(n6713) );
  AND3_X1 U8285 ( .A1(n6865), .A2(n6676), .A3(n6675), .ZN(n6677) );
  NOR3_X1 U8286 ( .A1(n9432), .A2(n6713), .A3(n6677), .ZN(n6678) );
  NOR2_X1 U8287 ( .A1(n6679), .A2(n6678), .ZN(n6681) );
  NOR2_X1 U8288 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6141), .ZN(n7073) );
  AOI21_X1 U8289 ( .B1(n9420), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n7073), .ZN(
        n6680) );
  OAI211_X1 U8290 ( .C1(n6691), .C2(n9431), .A(n6681), .B(n6680), .ZN(P1_U3248) );
  OAI222_X1 U8291 ( .A1(n7875), .A2(P2_U3151), .B1(n8993), .B2(n6683), .C1(
        n6682), .C2(n8987), .ZN(P2_U3287) );
  INV_X1 U8292 ( .A(n6881), .ZN(n6875) );
  OAI222_X1 U8293 ( .A1(n10225), .A2(n9979), .B1(n10222), .B2(n6683), .C1(
        P1_U3086), .C2(n6875), .ZN(P1_U3347) );
  AOI21_X1 U8294 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n6685), .A(n6684), .ZN(
        n6706) );
  INV_X1 U8295 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6686) );
  MUX2_X1 U8296 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6686), .S(n6707), .Z(n6687)
         );
  INV_X1 U8297 ( .A(n6687), .ZN(n6705) );
  NOR2_X1 U8298 ( .A1(n6706), .A2(n6705), .ZN(n6704) );
  AOI21_X1 U8299 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n6707), .A(n6704), .ZN(
        n6690) );
  INV_X1 U8300 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6688) );
  MUX2_X1 U8301 ( .A(n6688), .B(P1_REG2_REG_7__SCAN_IN), .S(n6766), .Z(n6689)
         );
  NOR2_X1 U8302 ( .A1(n6690), .A2(n6689), .ZN(n6765) );
  AOI211_X1 U8303 ( .C1(n6690), .C2(n6689), .A(n9415), .B(n6765), .ZN(n6702)
         );
  NOR2_X1 U8304 ( .A1(n6691), .A2(n7093), .ZN(n6708) );
  INV_X1 U8305 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6692) );
  MUX2_X1 U8306 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6692), .S(n6707), .Z(n6693)
         );
  OAI21_X1 U8307 ( .B1(n6713), .B2(n6708), .A(n6693), .ZN(n6711) );
  NAND2_X1 U8308 ( .A1(n6707), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6696) );
  INV_X1 U8309 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6694) );
  MUX2_X1 U8310 ( .A(n6694), .B(P1_REG1_REG_7__SCAN_IN), .S(n6766), .Z(n6695)
         );
  AOI21_X1 U8311 ( .B1(n6711), .B2(n6696), .A(n6695), .ZN(n6777) );
  INV_X1 U8312 ( .A(n6777), .ZN(n6698) );
  NAND3_X1 U8313 ( .A1(n6711), .A2(n6696), .A3(n6695), .ZN(n6697) );
  NAND3_X1 U8314 ( .A1(n6698), .A2(n9436), .A3(n6697), .ZN(n6700) );
  AND2_X1 U8315 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7157) );
  AOI21_X1 U8316 ( .B1(n9420), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n7157), .ZN(
        n6699) );
  OAI211_X1 U8317 ( .C1(n9431), .C2(n6771), .A(n6700), .B(n6699), .ZN(n6701)
         );
  OR2_X1 U8318 ( .A1(n6702), .A2(n6701), .ZN(P1_U3250) );
  NAND2_X1 U8319 ( .A1(n9449), .A2(P1_U3973), .ZN(n6703) );
  OAI21_X1 U8320 ( .B1(P1_U3973), .B2(n5729), .A(n6703), .ZN(P1_U3585) );
  AOI211_X1 U8321 ( .C1(n6706), .C2(n6705), .A(n9415), .B(n6704), .ZN(n6719)
         );
  MUX2_X1 U8322 ( .A(n6692), .B(P1_REG1_REG_6__SCAN_IN), .S(n6707), .Z(n6710)
         );
  INV_X1 U8323 ( .A(n6708), .ZN(n6709) );
  NAND2_X1 U8324 ( .A1(n6710), .A2(n6709), .ZN(n6712) );
  OAI211_X1 U8325 ( .C1(n6713), .C2(n6712), .A(n9436), .B(n6711), .ZN(n6716)
         );
  NOR2_X1 U8326 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6714), .ZN(n7139) );
  AOI21_X1 U8327 ( .B1(n9420), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n7139), .ZN(
        n6715) );
  OAI211_X1 U8328 ( .C1(n9431), .C2(n6717), .A(n6716), .B(n6715), .ZN(n6718)
         );
  OR2_X1 U8329 ( .A1(n6719), .A2(n6718), .ZN(P1_U3249) );
  NAND2_X1 U8330 ( .A1(n9321), .A2(n6720), .ZN(n6727) );
  INV_X1 U8331 ( .A(n6723), .ZN(n6724) );
  NAND2_X1 U8332 ( .A1(n6928), .A2(n4407), .ZN(n6831) );
  INV_X1 U8333 ( .A(n6755), .ZN(n6728) );
  NAND2_X1 U8334 ( .A1(n6728), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6725) );
  AND2_X1 U8335 ( .A1(n6831), .A2(n6725), .ZN(n6726) );
  NAND2_X1 U8336 ( .A1(n6727), .A2(n6726), .ZN(n6829) );
  INV_X2 U8337 ( .A(n9168), .ZN(n9115) );
  NAND2_X1 U8338 ( .A1(n9321), .A2(n9115), .ZN(n6730) );
  AOI22_X1 U8339 ( .A1(n6928), .A2(n6720), .B1(n10226), .B2(n6728), .ZN(n6729)
         );
  NAND2_X1 U8340 ( .A1(n6730), .A2(n6729), .ZN(n6830) );
  XNOR2_X1 U8341 ( .A(n6829), .B(n6830), .ZN(n6854) );
  NAND2_X1 U8342 ( .A1(n8100), .A2(P1_B_REG_SCAN_IN), .ZN(n6732) );
  INV_X1 U8343 ( .A(n8060), .ZN(n6731) );
  MUX2_X1 U8344 ( .A(n6732), .B(P1_B_REG_SCAN_IN), .S(n6731), .Z(n6734) );
  NAND2_X1 U8345 ( .A1(n8106), .A2(n8100), .ZN(n10211) );
  OAI21_X1 U8346 ( .B1(n6805), .B2(P1_D_REG_1__SCAN_IN), .A(n10211), .ZN(n6810) );
  NOR2_X1 U8347 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .ZN(
        n10023) );
  NOR4_X1 U8348 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6737) );
  NOR4_X1 U8349 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n6736) );
  NOR4_X1 U8350 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_31__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6735) );
  AND4_X1 U8351 ( .A1(n10023), .A2(n6737), .A3(n6736), .A4(n6735), .ZN(n6743)
         );
  NOR4_X1 U8352 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n6741) );
  NOR4_X1 U8353 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n6740) );
  NOR4_X1 U8354 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_27__SCAN_IN), .ZN(n6739) );
  NOR4_X1 U8355 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n6738) );
  AND4_X1 U8356 ( .A1(n6741), .A2(n6740), .A3(n6739), .A4(n6738), .ZN(n6742)
         );
  AND2_X1 U8357 ( .A1(n6743), .A2(n6742), .ZN(n6806) );
  NOR2_X1 U8358 ( .A1(n6805), .A2(n6806), .ZN(n6794) );
  NOR2_X1 U8359 ( .A1(n6810), .A2(n6794), .ZN(n6744) );
  NAND2_X1 U8360 ( .A1(n8106), .A2(n8060), .ZN(n10212) );
  OAI21_X1 U8361 ( .B1(n6805), .B2(P1_D_REG_0__SCAN_IN), .A(n10212), .ZN(n6811) );
  INV_X1 U8362 ( .A(n6811), .ZN(n6941) );
  AND2_X1 U8363 ( .A1(n6744), .A2(n6941), .ZN(n6849) );
  INV_X1 U8364 ( .A(n6745), .ZN(n7919) );
  NAND2_X1 U8365 ( .A1(n6815), .A2(n6721), .ZN(n10299) );
  NAND2_X1 U8366 ( .A1(n10299), .A2(n6746), .ZN(n6753) );
  NOR2_X1 U8367 ( .A1(n6753), .A2(n6798), .ZN(n6747) );
  NOR2_X1 U8368 ( .A1(n6847), .A2(n6935), .ZN(n6749) );
  NAND2_X1 U8369 ( .A1(n6849), .A2(n6749), .ZN(n9305) );
  INV_X1 U8370 ( .A(n6849), .ZN(n6759) );
  AND2_X1 U8371 ( .A1(n6815), .A2(n6750), .ZN(n7004) );
  NAND2_X1 U8372 ( .A1(n6807), .A2(n7004), .ZN(n6751) );
  OR2_X1 U8373 ( .A1(n6759), .A2(n6751), .ZN(n6752) );
  NAND2_X1 U8374 ( .A1(n9746), .A2(n7002), .ZN(n6795) );
  NAND2_X1 U8375 ( .A1(n6752), .A2(n9673), .ZN(n9283) );
  AOI22_X1 U8376 ( .A1(n9320), .A2(n9295), .B1(n6928), .B2(n9283), .ZN(n6764)
         );
  NAND2_X1 U8377 ( .A1(n6753), .A2(n7751), .ZN(n6754) );
  NAND2_X1 U8378 ( .A1(n6759), .A2(n6754), .ZN(n6756) );
  NAND2_X1 U8379 ( .A1(n6934), .A2(n6721), .ZN(n6797) );
  NAND3_X1 U8380 ( .A1(n6756), .A2(n6755), .A3(n6797), .ZN(n6757) );
  NAND2_X1 U8381 ( .A1(n6757), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6761) );
  INV_X1 U8382 ( .A(n6847), .ZN(n6758) );
  NAND2_X1 U8383 ( .A1(n6759), .A2(n6758), .ZN(n6760) );
  NAND2_X1 U8384 ( .A1(n6761), .A2(n6760), .ZN(n6955) );
  OR3_X1 U8385 ( .A1(n6955), .A2(n6762), .A3(P1_U3086), .ZN(n6908) );
  NAND2_X1 U8386 ( .A1(n6908), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6763) );
  OAI211_X1 U8387 ( .C1(n6854), .C2(n9285), .A(n6764), .B(n6763), .ZN(P1_U3232) );
  INV_X1 U8388 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6767) );
  MUX2_X1 U8389 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n6767), .S(n6881), .Z(n6768)
         );
  INV_X1 U8390 ( .A(n6768), .ZN(n6769) );
  AOI211_X1 U8391 ( .C1(n6770), .C2(n6769), .A(n9415), .B(n6880), .ZN(n6781)
         );
  NOR2_X1 U8392 ( .A1(n6771), .A2(n6694), .ZN(n6775) );
  INV_X1 U8393 ( .A(n6775), .ZN(n6773) );
  INV_X1 U8394 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6876) );
  MUX2_X1 U8395 ( .A(n6876), .B(P1_REG1_REG_8__SCAN_IN), .S(n6881), .Z(n6772)
         );
  NAND2_X1 U8396 ( .A1(n6773), .A2(n6772), .ZN(n6776) );
  MUX2_X1 U8397 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n6876), .S(n6881), .Z(n6774)
         );
  OAI21_X1 U8398 ( .B1(n6777), .B2(n6775), .A(n6774), .ZN(n6874) );
  OAI211_X1 U8399 ( .C1(n6777), .C2(n6776), .A(n6874), .B(n9436), .ZN(n6779)
         );
  NOR2_X1 U8400 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9804), .ZN(n7573) );
  AOI21_X1 U8401 ( .B1(n9420), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n7573), .ZN(
        n6778) );
  OAI211_X1 U8402 ( .C1(n9431), .C2(n6875), .A(n6779), .B(n6778), .ZN(n6780)
         );
  OR2_X1 U8403 ( .A1(n6781), .A2(n6780), .ZN(P1_U3251) );
  INV_X1 U8404 ( .A(n6782), .ZN(n6784) );
  OAI222_X1 U8405 ( .A1(P2_U3151), .A2(n8085), .B1(n7922), .B2(n6784), .C1(
        n6783), .C2(n8987), .ZN(P2_U3286) );
  INV_X1 U8406 ( .A(n6912), .ZN(n6916) );
  OAI222_X1 U8407 ( .A1(n10225), .A2(n6785), .B1(n10222), .B2(n6784), .C1(
        n6916), .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U8408 ( .A(n6815), .ZN(n6788) );
  NAND2_X1 U8409 ( .A1(n6721), .A2(n6786), .ZN(n6787) );
  NAND2_X1 U8410 ( .A1(n6788), .A2(n6787), .ZN(n6789) );
  OR2_X1 U8411 ( .A1(n6816), .A2(n6789), .ZN(n7807) );
  NAND2_X1 U8412 ( .A1(n6790), .A2(n7751), .ZN(n6925) );
  OR2_X1 U8413 ( .A1(n7919), .A2(n4408), .ZN(n6792) );
  OAI21_X1 U8414 ( .B1(n10302), .B2(n10125), .A(n6814), .ZN(n6793) );
  NAND2_X1 U8415 ( .A1(n6928), .A2(n6815), .ZN(n6819) );
  NAND2_X1 U8416 ( .A1(n6605), .A2(n6934), .ZN(n10241) );
  NAND2_X1 U8417 ( .A1(n9320), .A2(n10152), .ZN(n6821) );
  AND3_X1 U8418 ( .A1(n6793), .A2(n6819), .A3(n6821), .ZN(n10267) );
  INV_X1 U8419 ( .A(n6794), .ZN(n6796) );
  AND3_X1 U8420 ( .A1(n6796), .A2(n6810), .A3(n6795), .ZN(n6943) );
  INV_X1 U8421 ( .A(n6797), .ZN(n6809) );
  OR2_X1 U8422 ( .A1(n6798), .A2(n6809), .ZN(n6940) );
  NOR2_X1 U8423 ( .A1(n6940), .A2(n6811), .ZN(n6799) );
  NAND2_X1 U8424 ( .A1(n10313), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6800) );
  OAI21_X1 U8425 ( .B1(n10267), .B2(n10313), .A(n6800), .ZN(P1_U3522) );
  INV_X1 U8426 ( .A(n6801), .ZN(n6803) );
  OAI222_X1 U8427 ( .A1(P2_U3151), .A2(n8424), .B1(n7922), .B2(n6803), .C1(
        n6802), .C2(n8987), .ZN(P2_U3285) );
  INV_X1 U8428 ( .A(n7026), .ZN(n7031) );
  OAI222_X1 U8429 ( .A1(n10225), .A2(n6804), .B1(n10222), .B2(n6803), .C1(
        n7031), .C2(P1_U3086), .ZN(P1_U3345) );
  NAND2_X1 U8430 ( .A1(n6807), .A2(n6806), .ZN(n6808) );
  NAND2_X1 U8431 ( .A1(n10265), .A2(n6808), .ZN(n6813) );
  NOR2_X1 U8432 ( .A1(n6810), .A2(n6809), .ZN(n6812) );
  NAND3_X1 U8433 ( .A1(n6813), .A2(n6812), .A3(n6811), .ZN(n7003) );
  INV_X1 U8434 ( .A(n6814), .ZN(n6817) );
  NOR3_X1 U8435 ( .A1(n6817), .A2(n6816), .A3(n6815), .ZN(n6824) );
  INV_X1 U8436 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6822) );
  OR2_X1 U8437 ( .A1(n6819), .A2(n6818), .ZN(n6820) );
  OAI211_X1 U8438 ( .C1(n6822), .C2(n9673), .A(n6821), .B(n6820), .ZN(n6823)
         );
  OAI21_X1 U8439 ( .B1(n6824), .B2(n6823), .A(n9757), .ZN(n6825) );
  OAI21_X1 U8440 ( .B1(n6826), .B2(n9757), .A(n6825), .ZN(P1_U3293) );
  INV_X1 U8441 ( .A(n6827), .ZN(n6872) );
  AOI22_X1 U8442 ( .A1(n8448), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n8991), .ZN(n6828) );
  OAI21_X1 U8443 ( .B1(n6872), .B2(n8993), .A(n6828), .ZN(P2_U3284) );
  NAND2_X1 U8444 ( .A1(n6830), .A2(n6829), .ZN(n6833) );
  NAND2_X1 U8445 ( .A1(n6831), .A2(n9165), .ZN(n6832) );
  NAND2_X1 U8446 ( .A1(n6833), .A2(n6832), .ZN(n6845) );
  NAND2_X1 U8447 ( .A1(n9320), .A2(n6720), .ZN(n6835) );
  NAND2_X1 U8448 ( .A1(n4901), .A2(n6956), .ZN(n6834) );
  NAND2_X1 U8449 ( .A1(n6835), .A2(n6834), .ZN(n6836) );
  XNOR2_X1 U8450 ( .A(n6836), .B(n9165), .ZN(n6841) );
  INV_X1 U8451 ( .A(n6841), .ZN(n6839) );
  INV_X2 U8452 ( .A(n9062), .ZN(n9074) );
  AND2_X1 U8453 ( .A1(n4901), .A2(n6720), .ZN(n6837) );
  INV_X1 U8454 ( .A(n6840), .ZN(n6838) );
  INV_X1 U8455 ( .A(n6845), .ZN(n6842) );
  INV_X1 U8456 ( .A(n6892), .ZN(n6843) );
  AOI21_X1 U8457 ( .B1(n6845), .B2(n6844), .A(n6843), .ZN(n6853) );
  INV_X1 U8458 ( .A(n9283), .ZN(n9310) );
  NOR2_X1 U8459 ( .A1(n6847), .A2(n6605), .ZN(n6848) );
  AOI22_X1 U8460 ( .A1(n9295), .A2(n6893), .B1(n9321), .B2(n9303), .ZN(n6850)
         );
  OAI21_X1 U8461 ( .B1(n8124), .B2(n9310), .A(n6850), .ZN(n6851) );
  AOI21_X1 U8462 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n6908), .A(n6851), .ZN(
        n6852) );
  OAI21_X1 U8463 ( .B1(n6853), .B2(n9285), .A(n6852), .ZN(P1_U3222) );
  MUX2_X1 U8464 ( .A(n9331), .B(n6854), .S(n10223), .Z(n6855) );
  NAND2_X1 U8465 ( .A1(n6855), .A2(n6935), .ZN(n6856) );
  OAI211_X1 U8466 ( .C1(n10226), .C2(n6857), .A(n6856), .B(P1_U3973), .ZN(
        n9346) );
  INV_X1 U8467 ( .A(n9346), .ZN(n6871) );
  INV_X1 U8468 ( .A(n9415), .ZN(n9437) );
  OAI211_X1 U8469 ( .C1(n6860), .C2(n6859), .A(n9437), .B(n6858), .ZN(n6869)
         );
  AND2_X1 U8470 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n7105) );
  AOI21_X1 U8471 ( .B1(n9420), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n7105), .ZN(
        n6868) );
  INV_X1 U8472 ( .A(n9431), .ZN(n9379) );
  NAND2_X1 U8473 ( .A1(n9379), .A2(n6861), .ZN(n6867) );
  MUX2_X1 U8474 ( .A(n6672), .B(P1_REG1_REG_4__SCAN_IN), .S(n6861), .Z(n6862)
         );
  NAND3_X1 U8475 ( .A1(n9356), .A2(n6863), .A3(n6862), .ZN(n6864) );
  NAND3_X1 U8476 ( .A1(n9436), .A2(n6865), .A3(n6864), .ZN(n6866) );
  NAND4_X1 U8477 ( .A1(n6869), .A2(n6868), .A3(n6867), .A4(n6866), .ZN(n6870)
         );
  OR2_X1 U8478 ( .A1(n6871), .A2(n6870), .ZN(P1_U3247) );
  INV_X1 U8479 ( .A(n7263), .ZN(n7037) );
  OAI222_X1 U8480 ( .A1(n10225), .A2(n6873), .B1(n10222), .B2(n6872), .C1(
        P1_U3086), .C2(n7037), .ZN(P1_U3344) );
  OAI21_X1 U8481 ( .B1(n6876), .B2(n6875), .A(n6874), .ZN(n6879) );
  INV_X1 U8482 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6877) );
  MUX2_X1 U8483 ( .A(n6877), .B(P1_REG1_REG_9__SCAN_IN), .S(n6912), .Z(n6878)
         );
  NOR2_X1 U8484 ( .A1(n6878), .A2(n6879), .ZN(n6915) );
  AOI21_X1 U8485 ( .B1(n6879), .B2(n6878), .A(n6915), .ZN(n6888) );
  INV_X1 U8486 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9784) );
  AOI22_X1 U8487 ( .A1(n6912), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n9784), .B2(
        n6916), .ZN(n6882) );
  AOI221_X1 U8488 ( .B1(n6883), .B2(n6911), .C1(n6882), .C2(n6911), .A(n9415), 
        .ZN(n6884) );
  INV_X1 U8489 ( .A(n6884), .ZN(n6887) );
  AND2_X1 U8490 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7675) );
  INV_X1 U8491 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10003) );
  NOR2_X1 U8492 ( .A1(n9443), .A2(n10003), .ZN(n6885) );
  AOI211_X1 U8493 ( .C1(n9379), .C2(n6912), .A(n7675), .B(n6885), .ZN(n6886)
         );
  OAI211_X1 U8494 ( .C1(n6888), .C2(n9432), .A(n6887), .B(n6886), .ZN(P1_U3252) );
  INV_X1 U8495 ( .A(n6889), .ZN(n6950) );
  AOI22_X1 U8496 ( .A1(n7475), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n10215), .ZN(n6890) );
  OAI21_X1 U8497 ( .B1(n6950), .B2(n10222), .A(n6890), .ZN(P1_U3343) );
  AOI22_X1 U8498 ( .A1(n9303), .A2(n9320), .B1(n9319), .B2(n9295), .ZN(n6891)
         );
  OAI21_X1 U8499 ( .B1(n10269), .B2(n9310), .A(n6891), .ZN(n6907) );
  NAND2_X1 U8500 ( .A1(n6892), .A2(n6903), .ZN(n6901) );
  NAND2_X1 U8501 ( .A1(n6893), .A2(n6720), .ZN(n6895) );
  NAND2_X1 U8502 ( .A1(n7020), .A2(n6956), .ZN(n6894) );
  NAND2_X1 U8503 ( .A1(n6895), .A2(n6894), .ZN(n6896) );
  XNOR2_X1 U8504 ( .A(n6896), .B(n9165), .ZN(n6899) );
  AND2_X1 U8505 ( .A1(n7020), .A2(n6720), .ZN(n6897) );
  AOI21_X1 U8506 ( .B1(n6893), .B2(n9115), .A(n6897), .ZN(n6898) );
  NAND2_X1 U8507 ( .A1(n6899), .A2(n6898), .ZN(n6962) );
  OR2_X1 U8508 ( .A1(n6899), .A2(n6898), .ZN(n6900) );
  NAND2_X1 U8509 ( .A1(n6901), .A2(n6902), .ZN(n6963) );
  INV_X1 U8510 ( .A(n6902), .ZN(n6904) );
  NAND3_X1 U8511 ( .A1(n6904), .A2(n6892), .A3(n6903), .ZN(n6905) );
  AOI21_X1 U8512 ( .B1(n6963), .B2(n6905), .A(n9285), .ZN(n6906) );
  AOI211_X1 U8513 ( .C1(P1_REG3_REG_2__SCAN_IN), .C2(n6908), .A(n6907), .B(
        n6906), .ZN(n6909) );
  INV_X1 U8514 ( .A(n6909), .ZN(P1_U3237) );
  NAND2_X1 U8515 ( .A1(n7026), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6910) );
  OAI21_X1 U8516 ( .B1(n7026), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6910), .ZN(
        n6914) );
  OAI21_X1 U8517 ( .B1(n6912), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6911), .ZN(
        n6913) );
  NOR2_X1 U8518 ( .A1(n6914), .A2(n6913), .ZN(n7025) );
  AOI211_X1 U8519 ( .C1(n6914), .C2(n6913), .A(n7025), .B(n9415), .ZN(n6924)
         );
  AOI21_X1 U8520 ( .B1(n6916), .B2(n6877), .A(n6915), .ZN(n6919) );
  INV_X1 U8521 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6917) );
  MUX2_X1 U8522 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6917), .S(n7026), .Z(n6918)
         );
  NAND2_X1 U8523 ( .A1(n6918), .A2(n6919), .ZN(n7030) );
  OAI211_X1 U8524 ( .C1(n6919), .C2(n6918), .A(n9436), .B(n7030), .ZN(n6922)
         );
  NOR2_X1 U8525 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6920), .ZN(n8129) );
  AOI21_X1 U8526 ( .B1(n9420), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n8129), .ZN(
        n6921) );
  OAI211_X1 U8527 ( .C1(n9431), .C2(n7031), .A(n6922), .B(n6921), .ZN(n6923)
         );
  OR2_X1 U8528 ( .A1(n6924), .A2(n6923), .ZN(P1_U3253) );
  INV_X1 U8529 ( .A(n6925), .ZN(n7861) );
  NAND2_X1 U8530 ( .A1(n6926), .A2(n6927), .ZN(n6972) );
  OAI21_X1 U8531 ( .B1(n6926), .B2(n6927), .A(n6972), .ZN(n8118) );
  NAND2_X1 U8532 ( .A1(n4901), .A2(n6928), .ZN(n6929) );
  NAND2_X1 U8533 ( .A1(n6929), .A2(n9746), .ZN(n6930) );
  NOR2_X1 U8534 ( .A1(n7017), .A2(n6930), .ZN(n8121) );
  INV_X1 U8535 ( .A(n6931), .ZN(n6932) );
  AOI21_X1 U8536 ( .B1(n6933), .B2(n6926), .A(n6932), .ZN(n6939) );
  NAND2_X1 U8537 ( .A1(n6935), .A2(n6934), .ZN(n10243) );
  AOI22_X1 U8538 ( .A1(n10152), .A2(n6893), .B1(n9321), .B2(n10155), .ZN(n6938) );
  INV_X1 U8539 ( .A(n7807), .ZN(n6936) );
  NAND2_X1 U8540 ( .A1(n8118), .A2(n6936), .ZN(n6937) );
  OAI211_X1 U8541 ( .C1(n6939), .C2(n10250), .A(n6938), .B(n6937), .ZN(n8117)
         );
  AOI211_X1 U8542 ( .C1(n7861), .C2(n8118), .A(n8121), .B(n8117), .ZN(n6949)
         );
  NOR2_X1 U8543 ( .A1(n6941), .A2(n6940), .ZN(n6942) );
  NAND2_X1 U8544 ( .A1(n10306), .A2(n10248), .ZN(n10209) );
  INV_X1 U8545 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6944) );
  OAI22_X1 U8546 ( .A1(n10209), .A2(n8124), .B1(n10306), .B2(n6944), .ZN(n6945) );
  INV_X1 U8547 ( .A(n6945), .ZN(n6946) );
  OAI21_X1 U8548 ( .B1(n6949), .B2(n10304), .A(n6946), .ZN(P1_U3456) );
  OAI22_X1 U8549 ( .A1(n10163), .A2(n8124), .B1(n10316), .B2(n6666), .ZN(n6947) );
  INV_X1 U8550 ( .A(n6947), .ZN(n6948) );
  OAI21_X1 U8551 ( .B1(n6949), .B2(n10313), .A(n6948), .ZN(P1_U3523) );
  OAI222_X1 U8552 ( .A1(P2_U3151), .A2(n8466), .B1(n7922), .B2(n6950), .C1(
        n9978), .C2(n8987), .ZN(P2_U3283) );
  INV_X1 U8553 ( .A(n6951), .ZN(n6954) );
  AOI22_X1 U8554 ( .A1(n7584), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n10215), .ZN(n6952) );
  OAI21_X1 U8555 ( .B1(n6954), .B2(n10222), .A(n6952), .ZN(P1_U3342) );
  AOI22_X1 U8556 ( .A1(n8493), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n8991), .ZN(n6953) );
  OAI21_X1 U8557 ( .B1(n6954), .B2(n7922), .A(n6953), .ZN(P2_U3282) );
  INV_X1 U8558 ( .A(n9307), .ZN(n9281) );
  NAND2_X1 U8559 ( .A1(n9319), .A2(n6720), .ZN(n6958) );
  NAND2_X1 U8560 ( .A1(n6977), .A2(n9089), .ZN(n6957) );
  NAND2_X1 U8561 ( .A1(n6958), .A2(n6957), .ZN(n6960) );
  XNOR2_X1 U8562 ( .A(n6960), .B(n4410), .ZN(n7052) );
  AND2_X1 U8563 ( .A1(n6977), .A2(n6720), .ZN(n6961) );
  AOI21_X1 U8564 ( .B1(n9319), .B2(n9115), .A(n6961), .ZN(n7053) );
  XNOR2_X1 U8565 ( .A(n7052), .B(n7053), .ZN(n6965) );
  NAND2_X1 U8566 ( .A1(n6963), .A2(n6962), .ZN(n6964) );
  OAI21_X1 U8567 ( .B1(n6965), .B2(n6964), .A(n7056), .ZN(n6966) );
  NAND2_X1 U8568 ( .A1(n6966), .A2(n9300), .ZN(n6969) );
  NOR2_X1 U8569 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7042), .ZN(n9350) );
  OAI22_X1 U8570 ( .A1(n6976), .A2(n9293), .B1(n9310), .B2(n7045), .ZN(n6967)
         );
  AOI211_X1 U8571 ( .C1(n9295), .C2(n9318), .A(n9350), .B(n6967), .ZN(n6968)
         );
  OAI211_X1 U8572 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9281), .A(n6969), .B(
        n6968), .ZN(P1_U3218) );
  XOR2_X1 U8573 ( .A(n6409), .B(n6974), .Z(n7051) );
  NAND2_X1 U8574 ( .A1(n6970), .A2(n8124), .ZN(n6971) );
  NAND2_X1 U8575 ( .A1(n6972), .A2(n6971), .ZN(n7015) );
  NAND2_X1 U8576 ( .A1(n6976), .A2(n10269), .ZN(n6973) );
  NAND2_X1 U8577 ( .A1(n7013), .A2(n6973), .ZN(n6975) );
  NAND2_X1 U8578 ( .A1(n6975), .A2(n6974), .ZN(n6998) );
  OAI21_X1 U8579 ( .B1(n6975), .B2(n6974), .A(n6998), .ZN(n7048) );
  OAI22_X1 U8580 ( .A1(n6976), .A2(n10243), .B1(n7090), .B2(n10241), .ZN(n6978) );
  AOI211_X1 U8581 ( .C1(n6977), .C2(n7016), .A(n9723), .B(n4501), .ZN(n7047)
         );
  AOI211_X1 U8582 ( .C1(n10302), .C2(n7048), .A(n6978), .B(n7047), .ZN(n6979)
         );
  OAI21_X1 U8583 ( .B1(n7051), .B2(n10250), .A(n6979), .ZN(n6984) );
  INV_X1 U8584 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6980) );
  OAI22_X1 U8585 ( .A1(n10209), .A2(n7045), .B1(n10306), .B2(n6980), .ZN(n6981) );
  AOI21_X1 U8586 ( .B1(n6984), .B2(n10306), .A(n6981), .ZN(n6982) );
  INV_X1 U8587 ( .A(n6982), .ZN(P1_U3462) );
  OAI22_X1 U8588 ( .A1(n10163), .A2(n7045), .B1(n10316), .B2(n6669), .ZN(n6983) );
  AOI21_X1 U8589 ( .B1(n6984), .B2(n10316), .A(n6983), .ZN(n6985) );
  INV_X1 U8590 ( .A(n6985), .ZN(P1_U3525) );
  INV_X1 U8591 ( .A(n6986), .ZN(n6988) );
  INV_X1 U8592 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6991) );
  INV_X1 U8593 ( .A(n6989), .ZN(n6990) );
  AOI22_X1 U8594 ( .A1(n7040), .A2(n6991), .B1(n7300), .B2(n6990), .ZN(
        P2_U3376) );
  INV_X1 U8595 ( .A(n6992), .ZN(n6993) );
  AOI22_X1 U8596 ( .A1(n7040), .A2(n9996), .B1(n7300), .B2(n6993), .ZN(
        P2_U3377) );
  AND2_X1 U8597 ( .A1(n7040), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8598 ( .A1(n7040), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8599 ( .A1(n7040), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8600 ( .A1(n7040), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8601 ( .A1(n7040), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8602 ( .A1(n7040), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8603 ( .A1(n7040), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8604 ( .A1(n7040), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8605 ( .A1(n7040), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8606 ( .A1(n7040), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8607 ( .A1(n7040), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8608 ( .A1(n7040), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8609 ( .A1(n7040), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8610 ( .A1(n7040), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8611 ( .A1(n7040), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8612 ( .A1(n7040), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8613 ( .A1(n7040), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8614 ( .A1(n7040), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8615 ( .A1(n7040), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8616 ( .A1(n7040), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8617 ( .A1(n7040), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8618 ( .A1(n7040), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8619 ( .A1(n7040), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8620 ( .A1(n7040), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8621 ( .A1(n7040), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8622 ( .A1(n7040), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8623 ( .A1(n7040), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  XNOR2_X1 U8624 ( .A(n6995), .B(n6999), .ZN(n6996) );
  OAI222_X1 U8625 ( .A1(n10241), .A2(n7178), .B1(n10243), .B2(n7012), .C1(
        n6996), .C2(n10250), .ZN(n10276) );
  INV_X1 U8626 ( .A(n10276), .ZN(n7009) );
  NAND2_X1 U8627 ( .A1(n7012), .A2(n7045), .ZN(n6997) );
  NAND2_X1 U8628 ( .A1(n6998), .A2(n6997), .ZN(n7000) );
  NAND2_X1 U8629 ( .A1(n7000), .A2(n6999), .ZN(n7085) );
  OAI21_X1 U8630 ( .B1(n7000), .B2(n6999), .A(n7085), .ZN(n10278) );
  AOI21_X2 U8631 ( .B1(n7799), .B2(n7807), .A(n7001), .ZN(n9721) );
  INV_X1 U8632 ( .A(n4442), .ZN(n7088) );
  OAI211_X1 U8633 ( .C1(n10275), .C2(n4501), .A(n7088), .B(n9746), .ZN(n10274)
         );
  INV_X1 U8634 ( .A(n9757), .ZN(n9750) );
  AOI22_X1 U8635 ( .A1(n9750), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7104), .B2(
        n9748), .ZN(n7006) );
  NAND2_X1 U8636 ( .A1(n9751), .A2(n7106), .ZN(n7005) );
  OAI211_X1 U8637 ( .C1(n10274), .C2(n9755), .A(n7006), .B(n7005), .ZN(n7007)
         );
  AOI21_X1 U8638 ( .B1(n10278), .B2(n9721), .A(n7007), .ZN(n7008) );
  OAI21_X1 U8639 ( .B1(n7009), .B2(n7001), .A(n7008), .ZN(P1_U3289) );
  XOR2_X1 U8640 ( .A(n7014), .B(n7010), .Z(n7011) );
  OAI222_X1 U8641 ( .A1(n10241), .A2(n7012), .B1(n10243), .B2(n6970), .C1(
        n7011), .C2(n10250), .ZN(n10270) );
  INV_X1 U8642 ( .A(n10270), .ZN(n7024) );
  OAI21_X1 U8643 ( .B1(n7015), .B2(n7014), .A(n7013), .ZN(n10272) );
  OAI211_X1 U8644 ( .C1(n7017), .C2(n10269), .A(n7016), .B(n9746), .ZN(n10268)
         );
  NAND2_X1 U8645 ( .A1(n7001), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7018) );
  OAI21_X1 U8646 ( .B1(n9673), .B2(n6098), .A(n7018), .ZN(n7019) );
  AOI21_X1 U8647 ( .B1(n9751), .B2(n7020), .A(n7019), .ZN(n7021) );
  OAI21_X1 U8648 ( .B1(n9755), .B2(n10268), .A(n7021), .ZN(n7022) );
  AOI21_X1 U8649 ( .B1(n10272), .B2(n9721), .A(n7022), .ZN(n7023) );
  OAI21_X1 U8650 ( .B1(n7024), .B2(n7001), .A(n7023), .ZN(P1_U3291) );
  NAND2_X1 U8651 ( .A1(n7263), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7027) );
  OAI21_X1 U8652 ( .B1(n7263), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7027), .ZN(
        n7028) );
  AOI211_X1 U8653 ( .C1(n7029), .C2(n7028), .A(n7257), .B(n9415), .ZN(n7039)
         );
  OAI21_X1 U8654 ( .B1(n7031), .B2(n6917), .A(n7030), .ZN(n7034) );
  INV_X1 U8655 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7032) );
  MUX2_X1 U8656 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n7032), .S(n7263), .Z(n7033)
         );
  NAND2_X1 U8657 ( .A1(n7033), .A2(n7034), .ZN(n7261) );
  OAI211_X1 U8658 ( .C1(n7034), .C2(n7033), .A(n9436), .B(n7261), .ZN(n7036)
         );
  AND2_X1 U8659 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8038) );
  AOI21_X1 U8660 ( .B1(n9420), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n8038), .ZN(
        n7035) );
  OAI211_X1 U8661 ( .C1(n9431), .C2(n7037), .A(n7036), .B(n7035), .ZN(n7038)
         );
  OR2_X1 U8662 ( .A1(n7039), .A2(n7038), .ZN(P1_U3254) );
  INV_X1 U8663 ( .A(n7040), .ZN(n7041) );
  INV_X1 U8664 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n9949) );
  NOR2_X1 U8665 ( .A1(n7041), .A2(n9949), .ZN(P2_U3234) );
  INV_X1 U8666 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n10030) );
  NOR2_X1 U8667 ( .A1(n7041), .A2(n10030), .ZN(P2_U3262) );
  INV_X1 U8668 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n9847) );
  NOR2_X1 U8669 ( .A1(n7041), .A2(n9847), .ZN(P2_U3257) );
  NAND2_X1 U8670 ( .A1(n9757), .A2(n10125), .ZN(n9736) );
  OR2_X1 U8671 ( .A1(n7001), .A2(n10241), .ZN(n9730) );
  INV_X1 U8672 ( .A(n9730), .ZN(n7339) );
  NAND2_X1 U8673 ( .A1(n9757), .A2(n10155), .ZN(n9515) );
  INV_X1 U8674 ( .A(n9515), .ZN(n9726) );
  AOI22_X1 U8675 ( .A1(n7339), .A2(n9318), .B1(n9726), .B2(n6893), .ZN(n7044)
         );
  AOI22_X1 U8676 ( .A1(n9750), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9748), .B2(
        n7042), .ZN(n7043) );
  OAI211_X1 U8677 ( .C1(n7045), .C2(n9724), .A(n7044), .B(n7043), .ZN(n7046)
         );
  AOI21_X1 U8678 ( .B1(n7047), .B2(n9733), .A(n7046), .ZN(n7050) );
  NAND2_X1 U8679 ( .A1(n7048), .A2(n9721), .ZN(n7049) );
  OAI211_X1 U8680 ( .C1(n7051), .C2(n9736), .A(n7050), .B(n7049), .ZN(P1_U3290) );
  INV_X1 U8681 ( .A(n7052), .ZN(n7054) );
  NAND2_X1 U8682 ( .A1(n7054), .A2(n7053), .ZN(n7055) );
  NAND2_X1 U8683 ( .A1(n9318), .A2(n6720), .ZN(n7058) );
  NAND2_X1 U8684 ( .A1(n7106), .A2(n9089), .ZN(n7057) );
  NAND2_X1 U8685 ( .A1(n7058), .A2(n7057), .ZN(n7059) );
  XNOR2_X1 U8686 ( .A(n7059), .B(n9165), .ZN(n7062) );
  AND2_X1 U8687 ( .A1(n7106), .A2(n6720), .ZN(n7060) );
  AOI21_X1 U8688 ( .B1(n9318), .B2(n9115), .A(n7060), .ZN(n7063) );
  XNOR2_X1 U8689 ( .A(n7062), .B(n7063), .ZN(n7103) );
  INV_X1 U8690 ( .A(n7062), .ZN(n7065) );
  INV_X1 U8691 ( .A(n7063), .ZN(n7064) );
  NAND2_X1 U8692 ( .A1(n7065), .A2(n7064), .ZN(n7066) );
  NAND2_X1 U8693 ( .A1(n9317), .A2(n4409), .ZN(n7068) );
  NAND2_X1 U8694 ( .A1(n7089), .A2(n9089), .ZN(n7067) );
  NAND2_X1 U8695 ( .A1(n7068), .A2(n7067), .ZN(n7069) );
  XNOR2_X1 U8696 ( .A(n7069), .B(n4410), .ZN(n7126) );
  NAND2_X1 U8697 ( .A1(n9317), .A2(n9115), .ZN(n7071) );
  NAND2_X1 U8698 ( .A1(n7089), .A2(n4409), .ZN(n7070) );
  NAND2_X1 U8699 ( .A1(n7071), .A2(n7070), .ZN(n7125) );
  INV_X1 U8700 ( .A(n7125), .ZN(n7123) );
  XNOR2_X1 U8701 ( .A(n7126), .B(n7123), .ZN(n7072) );
  XNOR2_X1 U8702 ( .A(n7128), .B(n7072), .ZN(n7078) );
  NAND2_X1 U8703 ( .A1(n9307), .A2(n7113), .ZN(n7075) );
  AOI21_X1 U8704 ( .B1(n9316), .B2(n9295), .A(n7073), .ZN(n7074) );
  OAI211_X1 U8705 ( .C1(n7090), .C2(n9293), .A(n7075), .B(n7074), .ZN(n7076)
         );
  AOI21_X1 U8706 ( .B1(n7089), .B2(n9283), .A(n7076), .ZN(n7077) );
  OAI21_X1 U8707 ( .B1(n7078), .B2(n9285), .A(n7077), .ZN(P1_U3227) );
  INV_X1 U8708 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7080) );
  INV_X1 U8709 ( .A(n7079), .ZN(n7082) );
  INV_X1 U8710 ( .A(n7846), .ZN(n7852) );
  OAI222_X1 U8711 ( .A1(n10225), .A2(n7080), .B1(n10222), .B2(n7082), .C1(
        P1_U3086), .C2(n7852), .ZN(P1_U3341) );
  INV_X1 U8712 ( .A(n8503), .ZN(n8510) );
  INV_X1 U8713 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7081) );
  OAI222_X1 U8714 ( .A1(n8510), .A2(P2_U3151), .B1(n7922), .B2(n7082), .C1(
        n7081), .C2(n8987), .ZN(P2_U3281) );
  XNOR2_X1 U8715 ( .A(n7083), .B(n7086), .ZN(n7122) );
  NAND2_X1 U8716 ( .A1(n7090), .A2(n10275), .ZN(n7084) );
  NAND2_X1 U8717 ( .A1(n7085), .A2(n7084), .ZN(n7087) );
  NAND2_X1 U8718 ( .A1(n7087), .A2(n7086), .ZN(n7180) );
  OAI21_X1 U8719 ( .B1(n7087), .B2(n7086), .A(n7180), .ZN(n7119) );
  AOI211_X1 U8720 ( .C1(n7089), .C2(n7088), .A(n9723), .B(n7237), .ZN(n7118)
         );
  OAI22_X1 U8721 ( .A1(n7090), .A2(n10243), .B1(n7160), .B2(n10241), .ZN(n7091) );
  AOI211_X1 U8722 ( .C1(n7119), .C2(n10302), .A(n7118), .B(n7091), .ZN(n7092)
         );
  OAI21_X1 U8723 ( .B1(n10250), .B2(n7122), .A(n7092), .ZN(n7098) );
  OAI22_X1 U8724 ( .A1(n10163), .A2(n7177), .B1(n10316), .B2(n7093), .ZN(n7094) );
  AOI21_X1 U8725 ( .B1(n7098), .B2(n10316), .A(n7094), .ZN(n7095) );
  INV_X1 U8726 ( .A(n7095), .ZN(P1_U3527) );
  INV_X1 U8727 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7096) );
  OAI22_X1 U8728 ( .A1(n10209), .A2(n7177), .B1(n10306), .B2(n7096), .ZN(n7097) );
  AOI21_X1 U8729 ( .B1(n7098), .B2(n10306), .A(n7097), .ZN(n7099) );
  INV_X1 U8730 ( .A(n7099), .ZN(P1_U3468) );
  INV_X1 U8731 ( .A(n7100), .ZN(n7101) );
  AOI211_X1 U8732 ( .C1(n7103), .C2(n7102), .A(n9285), .B(n7101), .ZN(n7112)
         );
  NAND2_X1 U8733 ( .A1(n9307), .A2(n7104), .ZN(n7110) );
  AOI21_X1 U8734 ( .B1(n9317), .B2(n9295), .A(n7105), .ZN(n7109) );
  NAND2_X1 U8735 ( .A1(n9283), .A2(n7106), .ZN(n7108) );
  NAND2_X1 U8736 ( .A1(n9319), .A2(n9303), .ZN(n7107) );
  NAND4_X1 U8737 ( .A1(n7110), .A2(n7109), .A3(n7108), .A4(n7107), .ZN(n7111)
         );
  OR2_X1 U8738 ( .A1(n7112), .A2(n7111), .ZN(P1_U3230) );
  NOR2_X1 U8739 ( .A1(n9724), .A2(n7177), .ZN(n7117) );
  NAND2_X1 U8740 ( .A1(n9726), .A2(n9318), .ZN(n7115) );
  AOI22_X1 U8741 ( .A1(n9750), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7113), .B2(
        n9748), .ZN(n7114) );
  OAI211_X1 U8742 ( .C1(n7160), .C2(n9730), .A(n7115), .B(n7114), .ZN(n7116)
         );
  AOI211_X1 U8743 ( .C1(n7118), .C2(n9733), .A(n7117), .B(n7116), .ZN(n7121)
         );
  NAND2_X1 U8744 ( .A1(n7119), .A2(n9721), .ZN(n7120) );
  OAI211_X1 U8745 ( .C1(n7122), .C2(n9736), .A(n7121), .B(n7120), .ZN(P1_U3288) );
  INV_X1 U8746 ( .A(n7126), .ZN(n7124) );
  NAND2_X1 U8747 ( .A1(n7124), .A2(n7123), .ZN(n7127) );
  NAND2_X1 U8748 ( .A1(n7239), .A2(n9089), .ZN(n7130) );
  NAND2_X1 U8749 ( .A1(n9316), .A2(n4409), .ZN(n7129) );
  NAND2_X1 U8750 ( .A1(n7130), .A2(n7129), .ZN(n7131) );
  XNOR2_X1 U8751 ( .A(n7131), .B(n4410), .ZN(n7134) );
  NAND2_X1 U8752 ( .A1(n7239), .A2(n4409), .ZN(n7133) );
  NAND2_X1 U8753 ( .A1(n9316), .A2(n9115), .ZN(n7132) );
  NAND2_X1 U8754 ( .A1(n7133), .A2(n7132), .ZN(n7135) );
  NAND2_X1 U8755 ( .A1(n7134), .A2(n7135), .ZN(n7149) );
  INV_X1 U8756 ( .A(n7134), .ZN(n7137) );
  INV_X1 U8757 ( .A(n7135), .ZN(n7136) );
  NAND2_X1 U8758 ( .A1(n7137), .A2(n7136), .ZN(n7151) );
  NAND2_X1 U8759 ( .A1(n7149), .A2(n7151), .ZN(n7138) );
  XNOR2_X1 U8760 ( .A(n7150), .B(n7138), .ZN(n7144) );
  NAND2_X1 U8761 ( .A1(n9307), .A2(n7238), .ZN(n7141) );
  AOI21_X1 U8762 ( .B1(n9315), .B2(n9295), .A(n7139), .ZN(n7140) );
  OAI211_X1 U8763 ( .C1(n7178), .C2(n9293), .A(n7141), .B(n7140), .ZN(n7142)
         );
  AOI21_X1 U8764 ( .B1(n7239), .B2(n9283), .A(n7142), .ZN(n7143) );
  OAI21_X1 U8765 ( .B1(n7144), .B2(n9285), .A(n7143), .ZN(P1_U3239) );
  INV_X1 U8766 ( .A(n8548), .ZN(n8523) );
  INV_X1 U8767 ( .A(n7145), .ZN(n7146) );
  INV_X1 U8768 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n9816) );
  OAI222_X1 U8769 ( .A1(n8523), .A2(P2_U3151), .B1(n7922), .B2(n7146), .C1(
        n9816), .C2(n8987), .ZN(P2_U3280) );
  INV_X1 U8770 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n9997) );
  OAI222_X1 U8771 ( .A1(n10225), .A2(n9997), .B1(n10222), .B2(n7146), .C1(
        P1_U3086), .C2(n9368), .ZN(P1_U3340) );
  INV_X1 U8772 ( .A(n7147), .ZN(n7190) );
  AOI22_X1 U8773 ( .A1(n9391), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n10215), .ZN(n7148) );
  OAI21_X1 U8774 ( .B1(n7190), .B2(n10222), .A(n7148), .ZN(P1_U3339) );
  NAND2_X1 U8775 ( .A1(n7152), .A2(n7151), .ZN(n7561) );
  AOI22_X1 U8776 ( .A1(n7326), .A2(n9089), .B1(n4409), .B2(n9315), .ZN(n7153)
         );
  XNOR2_X1 U8777 ( .A(n7153), .B(n4410), .ZN(n7558) );
  NAND2_X1 U8778 ( .A1(n7326), .A2(n4409), .ZN(n7155) );
  NAND2_X1 U8779 ( .A1(n9315), .A2(n9115), .ZN(n7154) );
  AND2_X1 U8780 ( .A1(n7155), .A2(n7154), .ZN(n7562) );
  XNOR2_X1 U8781 ( .A(n7558), .B(n7562), .ZN(n7156) );
  XNOR2_X1 U8782 ( .A(n7561), .B(n7156), .ZN(n7163) );
  NAND2_X1 U8783 ( .A1(n9307), .A2(n7170), .ZN(n7159) );
  AOI21_X1 U8784 ( .B1(n9314), .B2(n9295), .A(n7157), .ZN(n7158) );
  OAI211_X1 U8785 ( .C1(n7160), .C2(n9293), .A(n7159), .B(n7158), .ZN(n7161)
         );
  AOI21_X1 U8786 ( .B1(n7326), .B2(n9283), .A(n7161), .ZN(n7162) );
  OAI21_X1 U8787 ( .B1(n7163), .B2(n9285), .A(n7162), .ZN(P1_U3213) );
  INV_X1 U8788 ( .A(n7182), .ZN(n7164) );
  NOR2_X1 U8789 ( .A1(n7165), .A2(n7164), .ZN(n7166) );
  NAND2_X1 U8790 ( .A1(n7166), .A2(n7167), .ZN(n7337) );
  OAI21_X1 U8791 ( .B1(n7167), .B2(n7166), .A(n7337), .ZN(n7168) );
  NAND2_X1 U8792 ( .A1(n7168), .A2(n10125), .ZN(n7311) );
  NAND2_X1 U8793 ( .A1(n7237), .A2(n7183), .ZN(n7236) );
  AOI21_X1 U8794 ( .B1(n7236), .B2(n7326), .A(n9723), .ZN(n7169) );
  NAND2_X1 U8795 ( .A1(n7169), .A2(n7341), .ZN(n7309) );
  INV_X1 U8796 ( .A(n7309), .ZN(n7176) );
  NAND2_X1 U8797 ( .A1(n7326), .A2(n9751), .ZN(n7174) );
  NAND2_X1 U8798 ( .A1(n7339), .A2(n9314), .ZN(n7173) );
  AOI22_X1 U8799 ( .A1(n9750), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7170), .B2(
        n9748), .ZN(n7172) );
  NAND2_X1 U8800 ( .A1(n9726), .A2(n9316), .ZN(n7171) );
  NAND4_X1 U8801 ( .A1(n7174), .A2(n7173), .A3(n7172), .A4(n7171), .ZN(n7175)
         );
  AOI21_X1 U8802 ( .B1(n7176), .B2(n9733), .A(n7175), .ZN(n7188) );
  NAND2_X1 U8803 ( .A1(n7178), .A2(n7177), .ZN(n7179) );
  NAND2_X1 U8804 ( .A1(n7180), .A2(n7179), .ZN(n7233) );
  NAND2_X1 U8805 ( .A1(n7182), .A2(n7181), .ZN(n7241) );
  NAND2_X1 U8806 ( .A1(n7233), .A2(n7241), .ZN(n7235) );
  NAND2_X1 U8807 ( .A1(n7183), .A2(n7160), .ZN(n7184) );
  OAI21_X1 U8808 ( .B1(n7186), .B2(n7185), .A(n7329), .ZN(n7313) );
  NAND2_X1 U8809 ( .A1(n7313), .A2(n9721), .ZN(n7187) );
  OAI211_X1 U8810 ( .C1(n7311), .C2(n7001), .A(n7188), .B(n7187), .ZN(P1_U3286) );
  INV_X1 U8811 ( .A(n8556), .ZN(n8572) );
  INV_X1 U8812 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7189) );
  OAI222_X1 U8813 ( .A1(n8572), .A2(P2_U3151), .B1(n7922), .B2(n7190), .C1(
        n7189), .C2(n8987), .ZN(P2_U3279) );
  NAND2_X1 U8814 ( .A1(n7200), .A2(n8111), .ZN(n7191) );
  MUX2_X1 U8815 ( .A(n8592), .B(n7191), .S(n7199), .Z(n8618) );
  INV_X1 U8816 ( .A(n7285), .ZN(n7192) );
  XNOR2_X1 U8817 ( .A(n7194), .B(n7192), .ZN(n7274) );
  INV_X1 U8818 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7777) );
  INV_X1 U8819 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7193) );
  NAND2_X1 U8820 ( .A1(n7250), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7273) );
  AOI21_X1 U8821 ( .B1(n7194), .B2(n7285), .A(n7271), .ZN(n10323) );
  XNOR2_X1 U8822 ( .A(n7195), .B(n10317), .ZN(n10324) );
  NOR2_X1 U8823 ( .A1(n10323), .A2(n10324), .ZN(n10322) );
  XOR2_X1 U8824 ( .A(n7416), .B(n7417), .Z(n7196) );
  NAND2_X1 U8825 ( .A1(n7197), .A2(n7196), .ZN(n7415) );
  OAI21_X1 U8826 ( .B1(n7197), .B2(n7196), .A(n7415), .ZN(n7227) );
  NOR2_X2 U8827 ( .A1(n8592), .A2(n7198), .ZN(n8628) );
  NOR2_X1 U8828 ( .A1(n7199), .A2(P2_U3151), .ZN(n8990) );
  AND2_X1 U8829 ( .A1(n7200), .A2(n8990), .ZN(n7210) );
  INV_X1 U8830 ( .A(n7210), .ZN(n7249) );
  INV_X1 U8831 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7384) );
  INV_X1 U8832 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7492) );
  MUX2_X1 U8833 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n7492), .S(n10317), .Z(n10336) );
  INV_X1 U8834 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7211) );
  AND2_X1 U8835 ( .A1(n7211), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7202) );
  NAND2_X1 U8836 ( .A1(n7201), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7203) );
  OAI21_X1 U8837 ( .B1(n7285), .B2(n7202), .A(n7203), .ZN(n7270) );
  INV_X1 U8838 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9965) );
  OR2_X1 U8839 ( .A1(n7270), .A2(n9965), .ZN(n7204) );
  NAND2_X1 U8840 ( .A1(n7204), .A2(n7203), .ZN(n10335) );
  NAND2_X1 U8841 ( .A1(n10336), .A2(n10335), .ZN(n10334) );
  NAND2_X1 U8842 ( .A1(n10317), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7205) );
  NAND2_X1 U8843 ( .A1(n10334), .A2(n7205), .ZN(n7206) );
  NAND2_X1 U8844 ( .A1(n7206), .A2(n7416), .ZN(n7421) );
  OAI21_X1 U8845 ( .B1(n7206), .B2(n7416), .A(n7421), .ZN(n7208) );
  INV_X1 U8846 ( .A(n7423), .ZN(n7207) );
  AOI21_X1 U8847 ( .B1(n7384), .B2(n7208), .A(n7207), .ZN(n7209) );
  NAND2_X1 U8848 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7460) );
  OAI21_X1 U8849 ( .B1(n8634), .B2(n7209), .A(n7460), .ZN(n7226) );
  INV_X1 U8850 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7218) );
  INV_X1 U8851 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10352) );
  AND2_X1 U8852 ( .A1(n7211), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7212) );
  NAND2_X1 U8853 ( .A1(n7201), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7213) );
  OAI21_X1 U8854 ( .B1(n7285), .B2(n7212), .A(n7213), .ZN(n7278) );
  INV_X1 U8855 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7279) );
  NAND2_X1 U8856 ( .A1(n10317), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7214) );
  NAND2_X1 U8857 ( .A1(n10318), .A2(n7214), .ZN(n7215) );
  NAND2_X1 U8858 ( .A1(n7215), .A2(n7416), .ZN(n7426) );
  OAI21_X1 U8859 ( .B1(n7215), .B2(n7416), .A(n7426), .ZN(n7217) );
  INV_X1 U8860 ( .A(n7428), .ZN(n7216) );
  AOI21_X1 U8861 ( .B1(n7218), .B2(n7217), .A(n7216), .ZN(n7224) );
  INV_X1 U8862 ( .A(n7219), .ZN(n7220) );
  NOR2_X1 U8863 ( .A1(n7221), .A2(n7220), .ZN(n7222) );
  INV_X1 U8864 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n7223) );
  OAI22_X1 U8865 ( .A1(n8602), .A2(n7224), .B1(n10330), .B2(n7223), .ZN(n7225)
         );
  AOI211_X1 U8866 ( .C1(n7227), .C2(n8628), .A(n7226), .B(n7225), .ZN(n7228)
         );
  OAI21_X1 U8867 ( .B1(n7416), .B2(n8618), .A(n7228), .ZN(P2_U3185) );
  INV_X1 U8868 ( .A(n7229), .ZN(n7232) );
  INV_X1 U8869 ( .A(n9401), .ZN(n9408) );
  OAI222_X1 U8870 ( .A1(n10225), .A2(n7230), .B1(n10222), .B2(n7232), .C1(
        P1_U3086), .C2(n9408), .ZN(P1_U3338) );
  INV_X1 U8871 ( .A(n8597), .ZN(n8561) );
  OAI222_X1 U8872 ( .A1(n8561), .A2(P2_U3151), .B1(n7922), .B2(n7232), .C1(
        n7231), .C2(n8987), .ZN(P2_U3278) );
  OR2_X1 U8873 ( .A1(n7233), .A2(n7241), .ZN(n7234) );
  NAND2_X1 U8874 ( .A1(n7235), .A2(n7234), .ZN(n10280) );
  OAI211_X1 U8875 ( .C1(n7237), .C2(n7183), .A(n9746), .B(n7236), .ZN(n10281)
         );
  AOI22_X1 U8876 ( .A1(n9751), .A2(n7239), .B1(n9748), .B2(n7238), .ZN(n7240)
         );
  OAI21_X1 U8877 ( .B1(n10281), .B2(n9755), .A(n7240), .ZN(n7247) );
  XNOR2_X1 U8878 ( .A(n7242), .B(n7241), .ZN(n7243) );
  NAND2_X1 U8879 ( .A1(n7243), .A2(n10125), .ZN(n7245) );
  AOI22_X1 U8880 ( .A1(n10155), .A2(n9317), .B1(n9315), .B2(n10152), .ZN(n7244) );
  NAND2_X1 U8881 ( .A1(n7245), .A2(n7244), .ZN(n10284) );
  MUX2_X1 U8882 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10284), .S(n9757), .Z(n7246)
         );
  AOI211_X1 U8883 ( .C1(n9721), .C2(n10280), .A(n7247), .B(n7246), .ZN(n7248)
         );
  INV_X1 U8884 ( .A(n7248), .ZN(P1_U3287) );
  INV_X1 U8885 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n7255) );
  INV_X1 U8886 ( .A(n8628), .ZN(n10321) );
  NAND2_X1 U8887 ( .A1(n10321), .A2(n7249), .ZN(n7252) );
  OAI21_X1 U8888 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n7250), .A(n7273), .ZN(n7251) );
  AOI22_X1 U8889 ( .A1(n7252), .A2(n7251), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        P2_U3151), .ZN(n7254) );
  NAND2_X1 U8890 ( .A1(n10332), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7253) );
  OAI211_X1 U8891 ( .C1(n10330), .C2(n7255), .A(n7254), .B(n7253), .ZN(
        P2_U3182) );
  INV_X1 U8892 ( .A(n7475), .ZN(n7269) );
  NOR2_X1 U8893 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7256), .ZN(n9200) );
  INV_X1 U8894 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7472) );
  MUX2_X1 U8895 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n7472), .S(n7475), .Z(n7258)
         );
  NAND2_X1 U8896 ( .A1(n7473), .A2(n7258), .ZN(n7259) );
  AOI221_X1 U8897 ( .B1(n7473), .B2(n7259), .C1(n7258), .C2(n7259), .A(n9415), 
        .ZN(n7260) );
  AOI211_X1 U8898 ( .C1(n9420), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n9200), .B(
        n7260), .ZN(n7268) );
  INV_X1 U8899 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10311) );
  MUX2_X1 U8900 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10311), .S(n7475), .Z(n7265) );
  INV_X1 U8901 ( .A(n7261), .ZN(n7262) );
  AOI21_X1 U8902 ( .B1(n7263), .B2(P1_REG1_REG_11__SCAN_IN), .A(n7262), .ZN(
        n7264) );
  NAND2_X1 U8903 ( .A1(n7265), .A2(n7264), .ZN(n7466) );
  OAI21_X1 U8904 ( .B1(n7265), .B2(n7264), .A(n7466), .ZN(n7266) );
  NAND2_X1 U8905 ( .A1(n9436), .A2(n7266), .ZN(n7267) );
  OAI211_X1 U8906 ( .C1(n9431), .C2(n7269), .A(n7268), .B(n7267), .ZN(P1_U3255) );
  INV_X1 U8907 ( .A(n8634), .ZN(n10338) );
  XNOR2_X1 U8908 ( .A(n7270), .B(n9965), .ZN(n7283) );
  INV_X1 U8909 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7825) );
  INV_X1 U8910 ( .A(n7271), .ZN(n7272) );
  OAI211_X1 U8911 ( .C1(n7274), .C2(n7273), .A(n8628), .B(n7272), .ZN(n7275)
         );
  OAI21_X1 U8912 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n7825), .A(n7275), .ZN(n7282) );
  INV_X1 U8913 ( .A(n7276), .ZN(n7277) );
  AOI21_X1 U8914 ( .B1(n7279), .B2(n7278), .A(n7277), .ZN(n7280) );
  OAI22_X1 U8915 ( .A1(n8602), .A2(n7280), .B1(n10379), .B2(n10330), .ZN(n7281) );
  AOI211_X1 U8916 ( .C1(n10338), .C2(n7283), .A(n7282), .B(n7281), .ZN(n7284)
         );
  OAI21_X1 U8917 ( .B1(n7285), .B2(n8618), .A(n7284), .ZN(P2_U3183) );
  INV_X1 U8918 ( .A(n7286), .ZN(n7287) );
  NAND2_X1 U8919 ( .A1(n7305), .A2(n7287), .ZN(n7290) );
  OR2_X1 U8920 ( .A1(n7302), .A2(n7288), .ZN(n7289) );
  INV_X1 U8921 ( .A(n7291), .ZN(n7296) );
  AOI21_X1 U8922 ( .B1(n7297), .B2(n7293), .A(n7292), .ZN(n7294) );
  OAI21_X1 U8923 ( .B1(n7296), .B2(n7295), .A(n7294), .ZN(n7299) );
  AOI22_X1 U8924 ( .A1(n7299), .A2(P2_STATE_REG_SCAN_IN), .B1(n7298), .B2(
        n7297), .ZN(n7452) );
  AND2_X1 U8925 ( .A1(n7452), .A2(n7300), .ZN(n7414) );
  INV_X1 U8926 ( .A(n7414), .ZN(n7301) );
  NAND2_X1 U8927 ( .A1(n7301), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7308) );
  INV_X1 U8928 ( .A(n7359), .ZN(n7303) );
  NAND2_X1 U8929 ( .A1(n7305), .A2(n8908), .ZN(n7306) );
  AOI22_X1 U8930 ( .A1(n8355), .A2(n7304), .B1(n8367), .B2(n7768), .ZN(n7307)
         );
  OAI211_X1 U8931 ( .C1(n7771), .C2(n8373), .A(n7308), .B(n7307), .ZN(P2_U3172) );
  AOI22_X1 U8932 ( .A1(n10155), .A2(n9316), .B1(n9314), .B2(n10152), .ZN(n7310) );
  NAND3_X1 U8933 ( .A1(n7311), .A2(n7310), .A3(n7309), .ZN(n7312) );
  AOI21_X1 U8934 ( .B1(n10302), .B2(n7313), .A(n7312), .ZN(n7318) );
  INV_X1 U8935 ( .A(n10163), .ZN(n7863) );
  AOI22_X1 U8936 ( .A1(n7326), .A2(n7863), .B1(n10313), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n7314) );
  OAI21_X1 U8937 ( .B1(n7318), .B2(n10313), .A(n7314), .ZN(P1_U3529) );
  INV_X1 U8938 ( .A(n10209), .ZN(n7865) );
  INV_X1 U8939 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7315) );
  NOR2_X1 U8940 ( .A1(n10306), .A2(n7315), .ZN(n7316) );
  AOI21_X1 U8941 ( .B1(n7326), .B2(n7865), .A(n7316), .ZN(n7317) );
  OAI21_X1 U8942 ( .B1(n7318), .B2(n10304), .A(n7317), .ZN(P1_U3474) );
  OAI21_X1 U8943 ( .B1(n7322), .B2(n7320), .A(n7319), .ZN(n7830) );
  XNOR2_X1 U8944 ( .A(n7322), .B(n7321), .ZN(n7323) );
  OAI222_X1 U8945 ( .A1(n8899), .A2(n7461), .B1(n8901), .B2(n5092), .C1(n8896), 
        .C2(n7323), .ZN(n7827) );
  AOI21_X1 U8946 ( .B1(n5700), .B2(n7830), .A(n7827), .ZN(n7493) );
  INV_X1 U8947 ( .A(n8890), .ZN(n7324) );
  AOI22_X1 U8948 ( .A1(n7324), .A2(n4763), .B1(n8924), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n7325) );
  OAI21_X1 U8949 ( .B1(n7493), .B2(n8924), .A(n7325), .ZN(P2_U3460) );
  INV_X1 U8950 ( .A(n7326), .ZN(n7327) );
  NAND2_X1 U8951 ( .A1(n7327), .A2(n7576), .ZN(n7328) );
  NAND2_X1 U8952 ( .A1(n7390), .A2(n7330), .ZN(n7334) );
  OAI21_X1 U8953 ( .B1(n7331), .B2(n7334), .A(n7399), .ZN(n7351) );
  INV_X1 U8954 ( .A(n7351), .ZN(n7346) );
  INV_X1 U8955 ( .A(n7337), .ZN(n7333) );
  OAI21_X1 U8956 ( .B1(n7333), .B2(n7332), .A(n7334), .ZN(n7338) );
  INV_X1 U8957 ( .A(n7334), .ZN(n7336) );
  NAND3_X1 U8958 ( .A1(n7337), .A2(n7336), .A3(n7335), .ZN(n7391) );
  NAND3_X1 U8959 ( .A1(n7338), .A2(n10125), .A3(n7391), .ZN(n7349) );
  MUX2_X1 U8960 ( .A(n6767), .B(n7349), .S(n9757), .Z(n7345) );
  AOI22_X1 U8961 ( .A1(n7339), .A2(n9313), .B1(n9748), .B2(n7572), .ZN(n7340)
         );
  OAI21_X1 U8962 ( .B1(n7576), .B2(n9515), .A(n7340), .ZN(n7343) );
  OAI211_X1 U8963 ( .C1(n4827), .C2(n4826), .A(n9746), .B(n7503), .ZN(n7347)
         );
  NOR2_X1 U8964 ( .A1(n7347), .A2(n9755), .ZN(n7342) );
  AOI211_X1 U8965 ( .C1(n9751), .C2(n7578), .A(n7343), .B(n7342), .ZN(n7344)
         );
  OAI211_X1 U8966 ( .C1(n7346), .C2(n9759), .A(n7345), .B(n7344), .ZN(P1_U3285) );
  AOI22_X1 U8967 ( .A1(n10155), .A2(n9315), .B1(n9313), .B2(n10152), .ZN(n7348) );
  NAND3_X1 U8968 ( .A1(n7349), .A2(n7348), .A3(n7347), .ZN(n7350) );
  AOI21_X1 U8969 ( .B1(n10302), .B2(n7351), .A(n7350), .ZN(n7354) );
  AOI22_X1 U8970 ( .A1(n7578), .A2(n7863), .B1(n10313), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n7352) );
  OAI21_X1 U8971 ( .B1(n7354), .B2(n10313), .A(n7352), .ZN(P1_U3530) );
  AOI22_X1 U8972 ( .A1(n7578), .A2(n7865), .B1(n10304), .B2(
        P1_REG0_REG_8__SCAN_IN), .ZN(n7353) );
  OAI21_X1 U8973 ( .B1(n7354), .B2(n10304), .A(n7353), .ZN(P1_U3477) );
  INV_X1 U8974 ( .A(n9429), .ZN(n9423) );
  INV_X1 U8975 ( .A(n7355), .ZN(n7356) );
  OAI222_X1 U8976 ( .A1(P1_U3086), .A2(n9423), .B1(n10222), .B2(n7356), .C1(
        n9845), .C2(n10225), .ZN(P1_U3337) );
  INV_X1 U8977 ( .A(n8605), .ZN(n8599) );
  OAI222_X1 U8978 ( .A1(n8987), .A2(n7357), .B1(n7922), .B2(n7356), .C1(
        P2_U3151), .C2(n8599), .ZN(P2_U3277) );
  NOR2_X2 U8979 ( .A1(n7359), .A2(n7358), .ZN(n8377) );
  OAI22_X1 U8980 ( .A1(n8358), .A2(n4513), .B1(n7656), .B2(n8379), .ZN(n7360)
         );
  AOI21_X1 U8981 ( .B1(n7361), .B2(n8367), .A(n7360), .ZN(n7375) );
  XNOR2_X1 U8982 ( .A(n7731), .B(n7363), .ZN(n7364) );
  NAND3_X1 U8983 ( .A1(n7366), .A2(n7365), .A3(n7364), .ZN(n7368) );
  XNOR2_X1 U8984 ( .A(n8206), .B(n10344), .ZN(n7454) );
  XNOR2_X1 U8985 ( .A(n7454), .B(n7461), .ZN(n7372) );
  OAI21_X1 U8986 ( .B1(n7768), .B2(n8206), .A(n7370), .ZN(n7408) );
  NAND2_X1 U8987 ( .A1(n7371), .A2(n7372), .ZN(n7456) );
  OAI21_X1 U8988 ( .B1(n7372), .B2(n7371), .A(n7456), .ZN(n7373) );
  NAND2_X1 U8989 ( .A1(n7373), .A2(n8344), .ZN(n7374) );
  OAI211_X1 U8990 ( .C1(n7414), .C2(n10341), .A(n7375), .B(n7374), .ZN(
        P2_U3177) );
  OAI21_X1 U8991 ( .B1(n7377), .B2(n7378), .A(n7376), .ZN(n7701) );
  INV_X1 U8992 ( .A(n8405), .ZN(n7643) );
  XNOR2_X1 U8993 ( .A(n7379), .B(n7378), .ZN(n7380) );
  OAI222_X1 U8994 ( .A1(n8901), .A2(n7461), .B1(n8899), .B2(n7643), .C1(n8896), 
        .C2(n7380), .ZN(n7698) );
  AOI21_X1 U8995 ( .B1(n5700), .B2(n7701), .A(n7698), .ZN(n7387) );
  INV_X1 U8996 ( .A(n8980), .ZN(n7382) );
  AOI22_X1 U8997 ( .A1(n7382), .A2(n7381), .B1(n10375), .B2(
        P2_REG0_REG_3__SCAN_IN), .ZN(n7383) );
  OAI21_X1 U8998 ( .B1(n7387), .B2(n10375), .A(n7383), .ZN(P2_U3399) );
  OAI22_X1 U8999 ( .A1(n8890), .A2(n7697), .B1(n8925), .B2(n7384), .ZN(n7385)
         );
  INV_X1 U9000 ( .A(n7385), .ZN(n7386) );
  OAI21_X1 U9001 ( .B1(n7387), .B2(n8924), .A(n7386), .ZN(P2_U3462) );
  NAND2_X1 U9002 ( .A1(n7389), .A2(n7388), .ZN(n7400) );
  NAND2_X1 U9003 ( .A1(n7391), .A2(n7390), .ZN(n7392) );
  XOR2_X1 U9004 ( .A(n7400), .B(n7392), .Z(n7512) );
  XNOR2_X1 U9005 ( .A(n7503), .B(n7664), .ZN(n7393) );
  OAI22_X1 U9006 ( .A1(n7393), .A2(n9723), .B1(n8040), .B2(n10241), .ZN(n7510)
         );
  NAND2_X1 U9007 ( .A1(n7664), .A2(n9751), .ZN(n7395) );
  AOI22_X1 U9008 ( .A1(n9750), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7678), .B2(
        n9748), .ZN(n7394) );
  OAI211_X1 U9009 ( .C1(n7397), .C2(n9515), .A(n7395), .B(n7394), .ZN(n7396)
         );
  AOI21_X1 U9010 ( .B1(n7510), .B2(n9733), .A(n7396), .ZN(n7403) );
  NAND2_X1 U9011 ( .A1(n4826), .A2(n7397), .ZN(n7398) );
  NAND2_X1 U9012 ( .A1(n7401), .A2(n7400), .ZN(n7496) );
  OAI21_X1 U9013 ( .B1(n7401), .B2(n7400), .A(n7496), .ZN(n7514) );
  NAND2_X1 U9014 ( .A1(n7514), .A2(n9721), .ZN(n7402) );
  OAI211_X1 U9015 ( .C1(n7512), .C2(n9736), .A(n7403), .B(n7402), .ZN(P1_U3284) );
  INV_X1 U9016 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9834) );
  AND2_X1 U9017 ( .A1(n8912), .A2(n8896), .ZN(n7405) );
  NAND2_X1 U9018 ( .A1(n7768), .A2(n8908), .ZN(n7404) );
  NAND2_X1 U9019 ( .A1(n7304), .A2(n8780), .ZN(n7772) );
  OAI211_X1 U9020 ( .C1(n7771), .C2(n7405), .A(n7404), .B(n7772), .ZN(n8926)
         );
  NAND2_X1 U9021 ( .A1(n10372), .A2(n8926), .ZN(n7406) );
  OAI21_X1 U9022 ( .B1(n10372), .B2(n9834), .A(n7406), .ZN(P2_U3390) );
  OAI21_X1 U9023 ( .B1(n7409), .B2(n7408), .A(n7407), .ZN(n7412) );
  INV_X1 U9024 ( .A(n8367), .ZN(n8384) );
  AOI22_X1 U9025 ( .A1(n8355), .A2(n8407), .B1(n8377), .B2(n8408), .ZN(n7410)
         );
  OAI21_X1 U9026 ( .B1(n7826), .B2(n8384), .A(n7410), .ZN(n7411) );
  AOI21_X1 U9027 ( .B1(n8344), .B2(n7412), .A(n7411), .ZN(n7413) );
  OAI21_X1 U9028 ( .B1(n7414), .B2(n7825), .A(n7413), .ZN(P2_U3162) );
  XNOR2_X1 U9029 ( .A(n7445), .B(n7444), .ZN(n7419) );
  OAI21_X1 U9030 ( .B1(n7417), .B2(n7416), .A(n7415), .ZN(n7418) );
  NOR2_X1 U9031 ( .A1(n7418), .A2(n7419), .ZN(n7443) );
  AOI211_X1 U9032 ( .C1(n7419), .C2(n7418), .A(n10321), .B(n7443), .ZN(n7420)
         );
  INV_X1 U9033 ( .A(n7420), .ZN(n7433) );
  INV_X1 U9034 ( .A(n10330), .ZN(n7796) );
  XNOR2_X1 U9035 ( .A(n7444), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n7422) );
  AND3_X1 U9036 ( .A1(n7423), .A2(n7422), .A3(n7421), .ZN(n7424) );
  NOR2_X1 U9037 ( .A1(n7434), .A2(n7424), .ZN(n7425) );
  NAND2_X1 U9038 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7525) );
  OAI21_X1 U9039 ( .B1(n8634), .B2(n7425), .A(n7525), .ZN(n7431) );
  INV_X1 U9040 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10009) );
  MUX2_X1 U9041 ( .A(n10009), .B(P2_REG2_REG_4__SCAN_IN), .S(n7444), .Z(n7427)
         );
  NAND3_X1 U9042 ( .A1(n7428), .A2(n7427), .A3(n7426), .ZN(n7429) );
  AOI21_X1 U9043 ( .B1(n4503), .B2(n7429), .A(n8602), .ZN(n7430) );
  AOI211_X1 U9044 ( .C1(n7796), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n7431), .B(
        n7430), .ZN(n7432) );
  OAI211_X1 U9045 ( .C1(n8618), .C2(n7444), .A(n7433), .B(n7432), .ZN(P2_U3186) );
  INV_X1 U9046 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9981) );
  INV_X1 U9047 ( .A(n7435), .ZN(n7437) );
  NAND2_X1 U9048 ( .A1(n7435), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7542) );
  INV_X1 U9049 ( .A(n7542), .ZN(n7436) );
  AOI21_X1 U9050 ( .B1(n9981), .B2(n7437), .A(n7436), .ZN(n7442) );
  OAI21_X1 U9051 ( .B1(n7439), .B2(P2_REG2_REG_5__SCAN_IN), .A(n7547), .ZN(
        n7440) );
  AOI22_X1 U9052 ( .A1(n7796), .A2(P2_ADDR_REG_5__SCAN_IN), .B1(n10327), .B2(
        n7440), .ZN(n7441) );
  NAND2_X1 U9053 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7642) );
  OAI211_X1 U9054 ( .C1(n7442), .C2(n8634), .A(n7441), .B(n7642), .ZN(n7449)
         );
  XNOR2_X1 U9055 ( .A(n7535), .B(n7534), .ZN(n7447) );
  NOR2_X1 U9056 ( .A1(n7446), .A2(n7447), .ZN(n7533) );
  AOI211_X1 U9057 ( .C1(n7447), .C2(n7446), .A(n10321), .B(n7533), .ZN(n7448)
         );
  AOI211_X1 U9058 ( .C1(n10332), .C2(n7450), .A(n7449), .B(n7448), .ZN(n7451)
         );
  INV_X1 U9059 ( .A(n7451), .ZN(P2_U3187) );
  XNOR2_X1 U9060 ( .A(n8201), .B(n7697), .ZN(n7518) );
  XNOR2_X1 U9061 ( .A(n7518), .B(n8406), .ZN(n7458) );
  AOI211_X1 U9062 ( .C1(n7458), .C2(n7457), .A(n8373), .B(n7520), .ZN(n7459)
         );
  INV_X1 U9063 ( .A(n7459), .ZN(n7465) );
  INV_X1 U9064 ( .A(n7460), .ZN(n7463) );
  OAI22_X1 U9065 ( .A1(n7697), .A2(n8384), .B1(n8358), .B2(n7461), .ZN(n7462)
         );
  AOI211_X1 U9066 ( .C1(n8355), .C2(n8405), .A(n7463), .B(n7462), .ZN(n7464)
         );
  OAI211_X1 U9067 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8298), .A(n7465), .B(
        n7464), .ZN(P2_U3158) );
  INV_X1 U9068 ( .A(n7584), .ZN(n7482) );
  OAI21_X1 U9069 ( .B1(n7475), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7466), .ZN(
        n7468) );
  INV_X1 U9070 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10161) );
  MUX2_X1 U9071 ( .A(n10161), .B(P1_REG1_REG_13__SCAN_IN), .S(n7584), .Z(n7467) );
  NOR2_X1 U9072 ( .A1(n7468), .A2(n7467), .ZN(n7581) );
  AOI211_X1 U9073 ( .C1(n7468), .C2(n7467), .A(n9432), .B(n7581), .ZN(n7469)
         );
  INV_X1 U9074 ( .A(n7469), .ZN(n7481) );
  NOR2_X1 U9075 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10016), .ZN(n9259) );
  INV_X1 U9076 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7470) );
  MUX2_X1 U9077 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n7470), .S(n7584), .Z(n7471)
         );
  INV_X1 U9078 ( .A(n7471), .ZN(n7478) );
  NOR2_X1 U9079 ( .A1(n7473), .A2(n7472), .ZN(n7476) );
  OAI22_X1 U9080 ( .A1(n7476), .A2(n7475), .B1(n7474), .B2(
        P1_REG2_REG_12__SCAN_IN), .ZN(n7477) );
  NOR2_X1 U9081 ( .A1(n7477), .A2(n7478), .ZN(n7583) );
  AOI211_X1 U9082 ( .C1(n7478), .C2(n7477), .A(n7583), .B(n9415), .ZN(n7479)
         );
  AOI211_X1 U9083 ( .C1(n9420), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n9259), .B(
        n7479), .ZN(n7480) );
  OAI211_X1 U9084 ( .C1(n9431), .C2(n7482), .A(n7481), .B(n7480), .ZN(P1_U3256) );
  NOR2_X1 U9085 ( .A1(n10344), .A2(n8917), .ZN(n7490) );
  XNOR2_X1 U9086 ( .A(n7485), .B(n7484), .ZN(n7489) );
  INV_X1 U9087 ( .A(n7979), .ZN(n7486) );
  NAND2_X1 U9088 ( .A1(n10348), .A2(n7486), .ZN(n7488) );
  AOI22_X1 U9089 ( .A1(n8782), .A2(n7304), .B1(n8406), .B2(n8780), .ZN(n7487)
         );
  OAI211_X1 U9090 ( .C1(n8896), .C2(n7489), .A(n7488), .B(n7487), .ZN(n10346)
         );
  AOI211_X1 U9091 ( .C1(n8922), .C2(n10348), .A(n7490), .B(n10346), .ZN(n10354) );
  OR2_X1 U9092 ( .A1(n10354), .A2(n8924), .ZN(n7491) );
  OAI21_X1 U9093 ( .B1(n8925), .B2(n7492), .A(n7491), .ZN(P2_U3461) );
  INV_X1 U9094 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9764) );
  MUX2_X1 U9095 ( .A(n9764), .B(n7493), .S(n10372), .Z(n7494) );
  OAI21_X1 U9096 ( .B1(n7826), .B2(n8980), .A(n7494), .ZN(P2_U3393) );
  NAND2_X1 U9097 ( .A1(n7496), .A2(n7495), .ZN(n7497) );
  OAI21_X1 U9098 ( .B1(n7497), .B2(n7501), .A(n4924), .ZN(n10290) );
  INV_X1 U9099 ( .A(n10290), .ZN(n7509) );
  INV_X1 U9100 ( .A(n7498), .ZN(n7499) );
  AOI21_X1 U9101 ( .B1(n7501), .B2(n7500), .A(n7499), .ZN(n7502) );
  OAI222_X1 U9102 ( .A1(n10241), .A2(n9202), .B1(n10243), .B2(n8132), .C1(
        n10250), .C2(n7502), .ZN(n10288) );
  OAI211_X1 U9103 ( .C1(n7504), .C2(n10287), .A(n7809), .B(n9746), .ZN(n10286)
         );
  AOI22_X1 U9104 ( .A1(n7001), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n8128), .B2(
        n9748), .ZN(n7506) );
  NAND2_X1 U9105 ( .A1(n8134), .A2(n9751), .ZN(n7505) );
  OAI211_X1 U9106 ( .C1(n10286), .C2(n9755), .A(n7506), .B(n7505), .ZN(n7507)
         );
  AOI21_X1 U9107 ( .B1(n10288), .B2(n9757), .A(n7507), .ZN(n7508) );
  OAI21_X1 U9108 ( .B1(n7509), .B2(n9759), .A(n7508), .ZN(P1_U3283) );
  AOI21_X1 U9109 ( .B1(n10155), .B2(n9314), .A(n7510), .ZN(n7511) );
  OAI21_X1 U9110 ( .B1(n7512), .B2(n10250), .A(n7511), .ZN(n7513) );
  AOI21_X1 U9111 ( .B1(n10302), .B2(n7514), .A(n7513), .ZN(n7517) );
  AOI22_X1 U9112 ( .A1(n7664), .A2(n7863), .B1(n10313), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n7515) );
  OAI21_X1 U9113 ( .B1(n7517), .B2(n10313), .A(n7515), .ZN(P1_U3531) );
  AOI22_X1 U9114 ( .A1(n7664), .A2(n7865), .B1(n10304), .B2(
        P1_REG0_REG_9__SCAN_IN), .ZN(n7516) );
  OAI21_X1 U9115 ( .B1(n7517), .B2(n10304), .A(n7516), .ZN(P1_U3480) );
  INV_X1 U9116 ( .A(n7723), .ZN(n7530) );
  XNOR2_X1 U9117 ( .A(n4406), .B(n7650), .ZN(n7521) );
  NOR2_X1 U9118 ( .A1(n7521), .A2(n8405), .ZN(n7637) );
  AOI21_X1 U9119 ( .B1(n7521), .B2(n8405), .A(n7637), .ZN(n7522) );
  OAI21_X1 U9120 ( .B1(n7523), .B2(n7522), .A(n7640), .ZN(n7524) );
  NAND2_X1 U9121 ( .A1(n7524), .A2(n8344), .ZN(n7529) );
  INV_X1 U9122 ( .A(n7525), .ZN(n7527) );
  OAI22_X1 U9123 ( .A1(n7650), .A2(n8384), .B1(n8358), .B2(n7656), .ZN(n7526)
         );
  AOI211_X1 U9124 ( .C1(n8355), .C2(n8404), .A(n7527), .B(n7526), .ZN(n7528)
         );
  OAI211_X1 U9125 ( .C1(n7530), .C2(n8298), .A(n7529), .B(n7528), .ZN(P2_U3170) );
  INV_X1 U9126 ( .A(n7531), .ZN(n8115) );
  OAI222_X1 U9127 ( .A1(n8617), .A2(P2_U3151), .B1(n7922), .B2(n8115), .C1(
        n7532), .C2(n8987), .ZN(P2_U3276) );
  XOR2_X1 U9128 ( .A(n7687), .B(n7683), .Z(n7536) );
  NAND2_X1 U9129 ( .A1(n7537), .A2(n7536), .ZN(n7682) );
  OAI21_X1 U9130 ( .B1(n7537), .B2(n7536), .A(n7682), .ZN(n7538) );
  NAND2_X1 U9131 ( .A1(n7538), .A2(n8628), .ZN(n7555) );
  INV_X1 U9132 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7540) );
  MUX2_X1 U9133 ( .A(n7540), .B(P2_REG1_REG_6__SCAN_IN), .S(n7687), .Z(n7541)
         );
  AND3_X1 U9134 ( .A1(n7542), .A2(n7541), .A3(n4853), .ZN(n7543) );
  NOR2_X1 U9135 ( .A1(n4505), .A2(n7543), .ZN(n7544) );
  NAND2_X1 U9136 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7743) );
  OAI21_X1 U9137 ( .B1(n8634), .B2(n7544), .A(n7743), .ZN(n7553) );
  INV_X1 U9138 ( .A(n7545), .ZN(n7548) );
  INV_X1 U9139 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7546) );
  MUX2_X1 U9140 ( .A(n7546), .B(P2_REG2_REG_6__SCAN_IN), .S(n7687), .Z(n7549)
         );
  INV_X1 U9141 ( .A(n7686), .ZN(n7551) );
  NAND3_X1 U9142 ( .A1(n7547), .A2(n7549), .A3(n7548), .ZN(n7550) );
  AOI21_X1 U9143 ( .B1(n7551), .B2(n7550), .A(n8602), .ZN(n7552) );
  AOI211_X1 U9144 ( .C1(n7796), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n7553), .B(
        n7552), .ZN(n7554) );
  OAI211_X1 U9145 ( .C1(n8618), .C2(n7687), .A(n7555), .B(n7554), .ZN(P2_U3188) );
  NAND2_X1 U9146 ( .A1(n7578), .A2(n4409), .ZN(n7557) );
  NAND2_X1 U9147 ( .A1(n9314), .A2(n9115), .ZN(n7556) );
  NAND2_X1 U9148 ( .A1(n7561), .A2(n7562), .ZN(n7560) );
  NAND2_X1 U9149 ( .A1(n7560), .A2(n7559), .ZN(n7566) );
  INV_X1 U9150 ( .A(n7561), .ZN(n7564) );
  INV_X1 U9151 ( .A(n7562), .ZN(n7563) );
  NAND2_X1 U9152 ( .A1(n7564), .A2(n7563), .ZN(n7565) );
  NAND2_X1 U9153 ( .A1(n7578), .A2(n9089), .ZN(n7568) );
  NAND2_X1 U9154 ( .A1(n9314), .A2(n4409), .ZN(n7567) );
  NAND2_X1 U9155 ( .A1(n7568), .A2(n7567), .ZN(n7569) );
  XNOR2_X1 U9156 ( .A(n7569), .B(n9165), .ZN(n7668) );
  INV_X1 U9157 ( .A(n7668), .ZN(n7671) );
  NOR2_X1 U9158 ( .A1(n7673), .A2(n7671), .ZN(n7665) );
  AOI21_X1 U9159 ( .B1(n7673), .B2(n7671), .A(n7665), .ZN(n7570) );
  NAND2_X1 U9160 ( .A1(n7570), .A2(n7669), .ZN(n7667) );
  OAI21_X1 U9161 ( .B1(n7669), .B2(n7570), .A(n7667), .ZN(n7571) );
  NAND2_X1 U9162 ( .A1(n7571), .A2(n9300), .ZN(n7580) );
  NAND2_X1 U9163 ( .A1(n9307), .A2(n7572), .ZN(n7575) );
  AOI21_X1 U9164 ( .B1(n9313), .B2(n9295), .A(n7573), .ZN(n7574) );
  OAI211_X1 U9165 ( .C1(n7576), .C2(n9293), .A(n7575), .B(n7574), .ZN(n7577)
         );
  AOI21_X1 U9166 ( .B1(n7578), .B2(n9283), .A(n7577), .ZN(n7579) );
  NAND2_X1 U9167 ( .A1(n7580), .A2(n7579), .ZN(P1_U3221) );
  INV_X1 U9168 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10314) );
  MUX2_X1 U9169 ( .A(n10314), .B(P1_REG1_REG_14__SCAN_IN), .S(n7846), .Z(n7850) );
  AOI21_X1 U9170 ( .B1(n7584), .B2(P1_REG1_REG_13__SCAN_IN), .A(n7581), .ZN(
        n7849) );
  XOR2_X1 U9171 ( .A(n7850), .B(n7849), .Z(n7590) );
  NOR2_X1 U9172 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9936), .ZN(n9135) );
  AOI21_X1 U9173 ( .B1(n9420), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n9135), .ZN(
        n7582) );
  OAI21_X1 U9174 ( .B1(n7852), .B2(n9431), .A(n7582), .ZN(n7589) );
  INV_X1 U9175 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7585) );
  AOI22_X1 U9176 ( .A1(n7846), .A2(n7585), .B1(P1_REG2_REG_14__SCAN_IN), .B2(
        n7852), .ZN(n7586) );
  AOI211_X1 U9177 ( .C1(n7587), .C2(n7586), .A(n7845), .B(n9415), .ZN(n7588)
         );
  AOI211_X1 U9178 ( .C1(n9436), .C2(n7590), .A(n7589), .B(n7588), .ZN(n7591)
         );
  INV_X1 U9179 ( .A(n7591), .ZN(P1_U3257) );
  NOR2_X1 U9180 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(P2_ADDR_REG_17__SCAN_IN), 
        .ZN(n7632) );
  NOR2_X1 U9181 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7630) );
  INV_X1 U9182 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9831) );
  INV_X1 U9183 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8520) );
  NOR2_X1 U9184 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7627) );
  NOR2_X1 U9185 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7624) );
  NOR2_X1 U9186 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7621) );
  NOR2_X1 U9187 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7618) );
  NOR2_X1 U9188 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7615) );
  NOR2_X1 U9189 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(P2_ADDR_REG_9__SCAN_IN), 
        .ZN(n7612) );
  NOR2_X1 U9190 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7609) );
  NOR2_X1 U9191 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7606) );
  NOR2_X1 U9192 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7604) );
  NOR2_X1 U9193 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7602) );
  NOR2_X1 U9194 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7600) );
  NAND2_X1 U9195 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n7597) );
  INV_X1 U9196 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n7592) );
  AOI22_X1 U9197 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .B1(n7592), .B2(n7223), .ZN(n10413) );
  NAND2_X1 U9198 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7595) );
  XOR2_X1 U9199 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10411) );
  INV_X1 U9200 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10380) );
  INV_X1 U9201 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9853) );
  OAI21_X1 U9202 ( .B1(n7255), .B2(n10380), .A(n9853), .ZN(n10376) );
  INV_X1 U9203 ( .A(n10376), .ZN(n7593) );
  NAND3_X1 U9204 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10377) );
  OAI21_X1 U9205 ( .B1(n7593), .B2(n10379), .A(n10377), .ZN(n10410) );
  NAND2_X1 U9206 ( .A1(n10411), .A2(n10410), .ZN(n7594) );
  NAND2_X1 U9207 ( .A1(n7595), .A2(n7594), .ZN(n10412) );
  NAND2_X1 U9208 ( .A1(n10413), .A2(n10412), .ZN(n7596) );
  NAND2_X1 U9209 ( .A1(n7597), .A2(n7596), .ZN(n10415) );
  INV_X1 U9210 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7598) );
  INV_X1 U9211 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9940) );
  AOI22_X1 U9212 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n7598), .B1(
        P2_ADDR_REG_4__SCAN_IN), .B2(n9940), .ZN(n10414) );
  NOR2_X1 U9213 ( .A1(n10415), .A2(n10414), .ZN(n7599) );
  NOR2_X1 U9214 ( .A1(n7600), .A2(n7599), .ZN(n10403) );
  XNOR2_X1 U9215 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10402) );
  NOR2_X1 U9216 ( .A1(n10403), .A2(n10402), .ZN(n7601) );
  NOR2_X1 U9217 ( .A1(n7602), .A2(n7601), .ZN(n10401) );
  XNOR2_X1 U9218 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n10400) );
  NOR2_X1 U9219 ( .A1(n10401), .A2(n10400), .ZN(n7603) );
  NOR2_X1 U9220 ( .A1(n7604), .A2(n7603), .ZN(n10407) );
  XNOR2_X1 U9221 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10406) );
  NOR2_X1 U9222 ( .A1(n10407), .A2(n10406), .ZN(n7605) );
  NOR2_X1 U9223 ( .A1(n7606), .A2(n7605), .ZN(n10409) );
  INV_X1 U9224 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n7607) );
  INV_X1 U9225 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n9773) );
  AOI22_X1 U9226 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n7607), .B1(
        P1_ADDR_REG_8__SCAN_IN), .B2(n9773), .ZN(n10408) );
  NOR2_X1 U9227 ( .A1(n10409), .A2(n10408), .ZN(n7608) );
  NOR2_X1 U9228 ( .A1(n7609), .A2(n7608), .ZN(n10405) );
  INV_X1 U9229 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7610) );
  AOI22_X1 U9230 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n7610), .B1(
        P2_ADDR_REG_9__SCAN_IN), .B2(n10003), .ZN(n10404) );
  NOR2_X1 U9231 ( .A1(n10405), .A2(n10404), .ZN(n7611) );
  NOR2_X1 U9232 ( .A1(n7612), .A2(n7611), .ZN(n10399) );
  INV_X1 U9233 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7613) );
  INV_X1 U9234 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n8094) );
  AOI22_X1 U9235 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n7613), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n8094), .ZN(n10398) );
  NOR2_X1 U9236 ( .A1(n10399), .A2(n10398), .ZN(n7614) );
  NOR2_X1 U9237 ( .A1(n7615), .A2(n7614), .ZN(n10397) );
  INV_X1 U9238 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7616) );
  INV_X1 U9239 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n8422) );
  AOI22_X1 U9240 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n7616), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n8422), .ZN(n10396) );
  NOR2_X1 U9241 ( .A1(n10397), .A2(n10396), .ZN(n7617) );
  NOR2_X1 U9242 ( .A1(n7618), .A2(n7617), .ZN(n10395) );
  INV_X1 U9243 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7619) );
  INV_X1 U9244 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n8446) );
  AOI22_X1 U9245 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n7619), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n8446), .ZN(n10394) );
  NOR2_X1 U9246 ( .A1(n10395), .A2(n10394), .ZN(n7620) );
  NOR2_X1 U9247 ( .A1(n7621), .A2(n7620), .ZN(n10393) );
  INV_X1 U9248 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7622) );
  INV_X1 U9249 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n9951) );
  AOI22_X1 U9250 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(n7622), .B1(
        P1_ADDR_REG_13__SCAN_IN), .B2(n9951), .ZN(n10392) );
  NOR2_X1 U9251 ( .A1(n10393), .A2(n10392), .ZN(n7623) );
  NOR2_X1 U9252 ( .A1(n7624), .A2(n7623), .ZN(n10391) );
  INV_X1 U9253 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7625) );
  INV_X1 U9254 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n9772) );
  AOI22_X1 U9255 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n7625), .B1(
        P1_ADDR_REG_14__SCAN_IN), .B2(n9772), .ZN(n10390) );
  NOR2_X1 U9256 ( .A1(n10391), .A2(n10390), .ZN(n7626) );
  NOR2_X1 U9257 ( .A1(n7627), .A2(n7626), .ZN(n10389) );
  AOI22_X1 U9258 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n8520), .B1(
        P2_ADDR_REG_15__SCAN_IN), .B2(n9831), .ZN(n10388) );
  NOR2_X1 U9259 ( .A1(n10389), .A2(n10388), .ZN(n7628) );
  AOI21_X1 U9260 ( .B1(n9831), .B2(n8520), .A(n7628), .ZN(n10387) );
  XNOR2_X1 U9261 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10386) );
  NOR2_X1 U9262 ( .A1(n10387), .A2(n10386), .ZN(n7629) );
  NOR2_X1 U9263 ( .A1(n7630), .A2(n7629), .ZN(n10385) );
  XNOR2_X1 U9264 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(P2_ADDR_REG_17__SCAN_IN), 
        .ZN(n10384) );
  NOR2_X1 U9265 ( .A1(n10385), .A2(n10384), .ZN(n7631) );
  NOR2_X1 U9266 ( .A1(n7632), .A2(n7631), .ZN(n7633) );
  AND2_X1 U9267 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n7633), .ZN(n10381) );
  NOR2_X1 U9268 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10381), .ZN(n7634) );
  NOR2_X1 U9269 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n7633), .ZN(n10382) );
  NOR2_X1 U9270 ( .A1(n7634), .A2(n10382), .ZN(n7636) );
  XNOR2_X1 U9271 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7635) );
  XNOR2_X1 U9272 ( .A(n7636), .B(n7635), .ZN(ADD_1068_U4) );
  INV_X1 U9273 ( .A(n7716), .ZN(n7648) );
  INV_X1 U9274 ( .A(n7637), .ZN(n7638) );
  XNOR2_X1 U9275 ( .A(n8201), .B(n7733), .ZN(n7738) );
  XNOR2_X1 U9276 ( .A(n7738), .B(n8404), .ZN(n7639) );
  AND3_X1 U9277 ( .A1(n7640), .A2(n7639), .A3(n7638), .ZN(n7641) );
  OAI21_X1 U9278 ( .B1(n7740), .B2(n7641), .A(n8344), .ZN(n7647) );
  INV_X1 U9279 ( .A(n7642), .ZN(n7645) );
  OAI22_X1 U9280 ( .A1(n7733), .A2(n8384), .B1(n8358), .B2(n7643), .ZN(n7644)
         );
  AOI211_X1 U9281 ( .C1(n8355), .C2(n8403), .A(n7645), .B(n7644), .ZN(n7646)
         );
  OAI211_X1 U9282 ( .C1(n7648), .C2(n8298), .A(n7647), .B(n7646), .ZN(P2_U3167) );
  INV_X1 U9283 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7659) );
  OAI21_X1 U9284 ( .B1(n7649), .B2(n7654), .A(n7713), .ZN(n7727) );
  NOR2_X1 U9285 ( .A1(n7650), .A2(n8917), .ZN(n7657) );
  INV_X1 U9286 ( .A(n8404), .ZN(n7744) );
  INV_X1 U9287 ( .A(n7651), .ZN(n7652) );
  AOI21_X1 U9288 ( .B1(n7654), .B2(n7653), .A(n7652), .ZN(n7655) );
  OAI222_X1 U9289 ( .A1(n8901), .A2(n7656), .B1(n8899), .B2(n7744), .C1(n8896), 
        .C2(n7655), .ZN(n7722) );
  AOI211_X1 U9290 ( .C1(n5700), .C2(n7727), .A(n7657), .B(n7722), .ZN(n10356)
         );
  OR2_X1 U9291 ( .A1(n10356), .A2(n8924), .ZN(n7658) );
  OAI21_X1 U9292 ( .B1(n8925), .B2(n7659), .A(n7658), .ZN(P2_U3463) );
  INV_X1 U9293 ( .A(n7664), .ZN(n7681) );
  NAND2_X1 U9294 ( .A1(n7664), .A2(n9089), .ZN(n7661) );
  NAND2_X1 U9295 ( .A1(n9313), .A2(n4409), .ZN(n7660) );
  NAND2_X1 U9296 ( .A1(n7661), .A2(n7660), .ZN(n7662) );
  XNOR2_X1 U9297 ( .A(n7662), .B(n9165), .ZN(n8019) );
  AND2_X1 U9298 ( .A1(n9313), .A2(n9115), .ZN(n7663) );
  AOI21_X1 U9299 ( .B1(n7664), .B2(n4409), .A(n7663), .ZN(n8018) );
  XNOR2_X1 U9300 ( .A(n8019), .B(n8018), .ZN(n7672) );
  INV_X1 U9301 ( .A(n7665), .ZN(n7666) );
  AND3_X1 U9302 ( .A1(n7667), .A2(n7672), .A3(n7666), .ZN(n7674) );
  INV_X1 U9303 ( .A(n7669), .ZN(n7670) );
  OAI21_X1 U9304 ( .B1(n7674), .B2(n8017), .A(n9300), .ZN(n7680) );
  AOI21_X1 U9305 ( .B1(n9312), .B2(n9295), .A(n7675), .ZN(n7676) );
  OAI21_X1 U9306 ( .B1(n7397), .B2(n9293), .A(n7676), .ZN(n7677) );
  AOI21_X1 U9307 ( .B1(n7678), .B2(n9307), .A(n7677), .ZN(n7679) );
  OAI211_X1 U9308 ( .C1(n7681), .C2(n9310), .A(n7680), .B(n7679), .ZN(P1_U3231) );
  XNOR2_X1 U9309 ( .A(n7778), .B(n4886), .ZN(n7780) );
  OAI21_X1 U9310 ( .B1(n7683), .B2(n7687), .A(n7682), .ZN(n7781) );
  XOR2_X1 U9311 ( .A(n7780), .B(n7781), .Z(n7696) );
  INV_X1 U9312 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7823) );
  AOI21_X1 U9313 ( .B1(n7823), .B2(n7685), .A(n7783), .ZN(n7693) );
  AND2_X1 U9314 ( .A1(n7688), .A2(n4886), .ZN(n7689) );
  NOR2_X1 U9315 ( .A1(n7789), .A2(n7689), .ZN(n7690) );
  NAND2_X1 U9316 ( .A1(n7690), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7792) );
  OAI21_X1 U9317 ( .B1(n7690), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7792), .ZN(
        n7691) );
  AOI22_X1 U9318 ( .A1(n7691), .A2(n10327), .B1(n7796), .B2(
        P2_ADDR_REG_7__SCAN_IN), .ZN(n7692) );
  NAND2_X1 U9319 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7900) );
  OAI211_X1 U9320 ( .C1(n7693), .C2(n8634), .A(n7692), .B(n7900), .ZN(n7694)
         );
  AOI21_X1 U9321 ( .B1(n4886), .B2(n10332), .A(n7694), .ZN(n7695) );
  OAI21_X1 U9322 ( .B1(n7696), .B2(n10321), .A(n7695), .ZN(P2_U3189) );
  OAI22_X1 U9323 ( .A1(n8810), .A2(n7697), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n10345), .ZN(n7700) );
  MUX2_X1 U9324 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n7698), .S(n10350), .Z(n7699)
         );
  AOI211_X1 U9325 ( .C1(n8825), .C2(n7701), .A(n7700), .B(n7699), .ZN(n7702)
         );
  INV_X1 U9326 ( .A(n7702), .ZN(P2_U3230) );
  INV_X1 U9327 ( .A(n8402), .ZN(n7955) );
  XNOR2_X1 U9328 ( .A(n7703), .B(n7704), .ZN(n7705) );
  OAI222_X1 U9329 ( .A1(n8901), .A2(n7744), .B1(n8899), .B2(n7955), .C1(n7705), 
        .C2(n8896), .ZN(n7760) );
  XNOR2_X1 U9330 ( .A(n7707), .B(n7706), .ZN(n7753) );
  OAI22_X1 U9331 ( .A1(n7753), .A2(n8912), .B1(n7745), .B2(n8917), .ZN(n7708)
         );
  NOR2_X1 U9332 ( .A1(n7760), .A2(n7708), .ZN(n10360) );
  OR2_X1 U9333 ( .A1(n8925), .A2(n7540), .ZN(n7709) );
  OAI21_X1 U9334 ( .B1(n10360), .B2(n8924), .A(n7709), .ZN(P2_U3465) );
  XOR2_X1 U9335 ( .A(n7710), .B(n7714), .Z(n7711) );
  AOI222_X1 U9336 ( .A1(n8785), .A2(n7711), .B1(n8405), .B2(n8782), .C1(n8403), 
        .C2(n8780), .ZN(n7732) );
  NAND2_X1 U9337 ( .A1(n7713), .A2(n7712), .ZN(n7715) );
  XNOR2_X1 U9338 ( .A(n7715), .B(n7714), .ZN(n7735) );
  INV_X1 U9339 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7719) );
  AOI22_X1 U9340 ( .A1(n8795), .A2(n7717), .B1(n8822), .B2(n7716), .ZN(n7718)
         );
  OAI21_X1 U9341 ( .B1(n7719), .B2(n10350), .A(n7718), .ZN(n7720) );
  AOI21_X1 U9342 ( .B1(n7735), .B2(n8825), .A(n7720), .ZN(n7721) );
  OAI21_X1 U9343 ( .B1(n7732), .B2(n10353), .A(n7721), .ZN(P2_U3228) );
  INV_X1 U9344 ( .A(n7722), .ZN(n7729) );
  AOI22_X1 U9345 ( .A1(n8795), .A2(n7724), .B1(n8822), .B2(n7723), .ZN(n7725)
         );
  OAI21_X1 U9346 ( .B1(n10009), .B2(n10350), .A(n7725), .ZN(n7726) );
  AOI21_X1 U9347 ( .B1(n7727), .B2(n8825), .A(n7726), .ZN(n7728) );
  OAI21_X1 U9348 ( .B1(n7729), .B2(n10353), .A(n7728), .ZN(P2_U3229) );
  INV_X1 U9349 ( .A(n7730), .ZN(n7750) );
  OAI222_X1 U9350 ( .A1(P2_U3151), .A2(n7731), .B1(n7922), .B2(n7750), .C1(
        n9989), .C2(n8987), .ZN(P2_U3275) );
  OAI21_X1 U9351 ( .B1(n7733), .B2(n8917), .A(n7732), .ZN(n7734) );
  AOI21_X1 U9352 ( .B1(n5700), .B2(n7735), .A(n7734), .ZN(n10358) );
  OR2_X1 U9353 ( .A1(n8925), .A2(n9981), .ZN(n7736) );
  OAI21_X1 U9354 ( .B1(n10358), .B2(n8924), .A(n7736), .ZN(P2_U3464) );
  INV_X1 U9355 ( .A(n7737), .ZN(n7755) );
  INV_X1 U9356 ( .A(n7738), .ZN(n7739) );
  XNOR2_X1 U9357 ( .A(n8201), .B(n7754), .ZN(n7894) );
  XNOR2_X1 U9358 ( .A(n7894), .B(n8403), .ZN(n7741) );
  OAI211_X1 U9359 ( .C1(n7742), .C2(n7741), .A(n7896), .B(n8344), .ZN(n7749)
         );
  INV_X1 U9360 ( .A(n7743), .ZN(n7747) );
  OAI22_X1 U9361 ( .A1(n7745), .A2(n8384), .B1(n8358), .B2(n7744), .ZN(n7746)
         );
  AOI211_X1 U9362 ( .C1(n8355), .C2(n8402), .A(n7747), .B(n7746), .ZN(n7748)
         );
  OAI211_X1 U9363 ( .C1(n7755), .C2(n8298), .A(n7749), .B(n7748), .ZN(P2_U3179) );
  OAI222_X1 U9364 ( .A1(n10225), .A2(n7752), .B1(P1_U3086), .B2(n7751), .C1(
        n10222), .C2(n7750), .ZN(P1_U3335) );
  NOR2_X1 U9365 ( .A1(n7753), .A2(n8792), .ZN(n7759) );
  NAND2_X1 U9366 ( .A1(n8795), .A2(n7754), .ZN(n7757) );
  OR2_X1 U9367 ( .A1(n10345), .A2(n7755), .ZN(n7756) );
  OAI211_X1 U9368 ( .C1(n7546), .C2(n10350), .A(n7757), .B(n7756), .ZN(n7758)
         );
  AOI211_X1 U9369 ( .C1(n7760), .C2(n10350), .A(n7759), .B(n7758), .ZN(n7761)
         );
  INV_X1 U9370 ( .A(n7761), .ZN(P2_U3227) );
  INV_X1 U9371 ( .A(n7762), .ZN(n7766) );
  OAI222_X1 U9372 ( .A1(P2_U3151), .A2(n7764), .B1(n7922), .B2(n7766), .C1(
        n7763), .C2(n8987), .ZN(P2_U3274) );
  OAI222_X1 U9373 ( .A1(P1_U3086), .A2(n7767), .B1(n10222), .B2(n7766), .C1(
        n7765), .C2(n10225), .ZN(P1_U3334) );
  AOI22_X1 U9374 ( .A1(n8795), .A2(n7768), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n8822), .ZN(n7776) );
  INV_X1 U9375 ( .A(n7769), .ZN(n7770) );
  NOR3_X1 U9376 ( .A1(n7771), .A2(n7770), .A3(n8908), .ZN(n7774) );
  INV_X1 U9377 ( .A(n7772), .ZN(n7773) );
  OAI21_X1 U9378 ( .B1(n7774), .B2(n7773), .A(n10350), .ZN(n7775) );
  OAI211_X1 U9379 ( .C1(n7777), .C2(n10350), .A(n7776), .B(n7775), .ZN(
        P2_U3233) );
  INV_X1 U9380 ( .A(n7778), .ZN(n7779) );
  AOI22_X1 U9381 ( .A1(n7781), .A2(n7780), .B1(n4886), .B2(n7779), .ZN(n7871)
         );
  XNOR2_X1 U9382 ( .A(n7869), .B(n7875), .ZN(n7870) );
  XNOR2_X1 U9383 ( .A(n7871), .B(n7870), .ZN(n7782) );
  NAND2_X1 U9384 ( .A1(n7782), .A2(n8628), .ZN(n7798) );
  INV_X1 U9385 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9968) );
  MUX2_X1 U9386 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9968), .S(n7875), .Z(n7784)
         );
  OAI21_X1 U9387 ( .B1(n7785), .B2(n7783), .A(n7784), .ZN(n7876) );
  INV_X1 U9388 ( .A(n7876), .ZN(n7787) );
  NOR3_X1 U9389 ( .A1(n7785), .A2(n7784), .A3(n7783), .ZN(n7786) );
  NOR2_X1 U9390 ( .A1(n7787), .A2(n7786), .ZN(n7788) );
  NAND2_X1 U9391 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7954) );
  OAI21_X1 U9392 ( .B1(n7788), .B2(n8634), .A(n7954), .ZN(n7795) );
  INV_X1 U9393 ( .A(n7789), .ZN(n7790) );
  XNOR2_X1 U9394 ( .A(n7875), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n7791) );
  NAND3_X1 U9395 ( .A1(n7792), .A2(n7791), .A3(n7790), .ZN(n7793) );
  AOI21_X1 U9396 ( .B1(n4497), .B2(n7793), .A(n8602), .ZN(n7794) );
  AOI211_X1 U9397 ( .C1(n7796), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n7795), .B(
        n7794), .ZN(n7797) );
  OAI211_X1 U9398 ( .C1(n8618), .C2(n7875), .A(n7798), .B(n7797), .ZN(P2_U3190) );
  INV_X1 U9399 ( .A(n7799), .ZN(n8119) );
  NOR2_X1 U9400 ( .A1(n8134), .A2(n9312), .ZN(n7800) );
  XNOR2_X1 U9401 ( .A(n7832), .B(n7802), .ZN(n7808) );
  INV_X1 U9402 ( .A(n7808), .ZN(n7862) );
  XNOR2_X1 U9403 ( .A(n7803), .B(n7802), .ZN(n7805) );
  OAI22_X1 U9404 ( .A1(n8040), .A2(n10243), .B1(n9261), .B2(n10241), .ZN(n7804) );
  AOI21_X1 U9405 ( .B1(n7805), .B2(n10125), .A(n7804), .ZN(n7806) );
  OAI21_X1 U9406 ( .B1(n7808), .B2(n7807), .A(n7806), .ZN(n7859) );
  AOI21_X1 U9407 ( .B1(n8119), .B2(n7862), .A(n7859), .ZN(n7813) );
  OR2_X1 U9408 ( .A1(n7809), .A2(n8028), .ZN(n7837) );
  AOI211_X1 U9409 ( .C1(n8028), .C2(n7809), .A(n9723), .B(n4832), .ZN(n7860)
         );
  INV_X1 U9410 ( .A(n8028), .ZN(n8045) );
  AOI22_X1 U9411 ( .A1(n9750), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n8042), .B2(
        n9748), .ZN(n7810) );
  OAI21_X1 U9412 ( .B1(n8045), .B2(n9724), .A(n7810), .ZN(n7811) );
  AOI21_X1 U9413 ( .B1(n7860), .B2(n9733), .A(n7811), .ZN(n7812) );
  OAI21_X1 U9414 ( .B1(n7813), .B2(n9750), .A(n7812), .ZN(P1_U3282) );
  NAND2_X1 U9415 ( .A1(n7816), .A2(n7815), .ZN(n7817) );
  NAND2_X1 U9416 ( .A1(n7814), .A2(n7817), .ZN(n7893) );
  AOI22_X1 U9417 ( .A1(n8780), .A2(n8401), .B1(n8403), .B2(n8782), .ZN(n7821)
         );
  XNOR2_X1 U9418 ( .A(n7818), .B(n4517), .ZN(n7819) );
  NAND2_X1 U9419 ( .A1(n7819), .A2(n8785), .ZN(n7820) );
  OAI211_X1 U9420 ( .C1(n7893), .C2(n7979), .A(n7821), .B(n7820), .ZN(n7887)
         );
  OAI22_X1 U9421 ( .A1(n7893), .A2(n7964), .B1(n7902), .B2(n8917), .ZN(n7822)
         );
  NOR2_X1 U9422 ( .A1(n7887), .A2(n7822), .ZN(n10362) );
  OR2_X1 U9423 ( .A1(n8925), .A2(n7823), .ZN(n7824) );
  OAI21_X1 U9424 ( .B1(n10362), .B2(n8924), .A(n7824), .ZN(P2_U3466) );
  OAI22_X1 U9425 ( .A1(n8810), .A2(n7826), .B1(n7825), .B2(n10345), .ZN(n7829)
         );
  MUX2_X1 U9426 ( .A(n7827), .B(P2_REG2_REG_1__SCAN_IN), .S(n10353), .Z(n7828)
         );
  AOI211_X1 U9427 ( .C1(n8825), .C2(n7830), .A(n7829), .B(n7828), .ZN(n7831)
         );
  INV_X1 U9428 ( .A(n7831), .ZN(P2_U3232) );
  XNOR2_X1 U9429 ( .A(n8004), .B(n7834), .ZN(n10296) );
  INV_X1 U9430 ( .A(n10296), .ZN(n7844) );
  OAI211_X1 U9431 ( .C1(n7834), .C2(n7833), .A(n8000), .B(n10125), .ZN(n7836)
         );
  AOI22_X1 U9432 ( .A1(n10155), .A2(n9311), .B1(n9742), .B2(n10152), .ZN(n7835) );
  NAND2_X1 U9433 ( .A1(n7836), .A2(n7835), .ZN(n10295) );
  INV_X1 U9434 ( .A(n8012), .ZN(n7838) );
  OAI211_X1 U9435 ( .C1(n10293), .C2(n4832), .A(n7838), .B(n9746), .ZN(n10292)
         );
  INV_X1 U9436 ( .A(n9204), .ZN(n7839) );
  OAI22_X1 U9437 ( .A1(n9757), .A2(n7472), .B1(n7839), .B2(n9673), .ZN(n7840)
         );
  AOI21_X1 U9438 ( .B1(n9000), .B2(n9751), .A(n7840), .ZN(n7841) );
  OAI21_X1 U9439 ( .B1(n10292), .B2(n9755), .A(n7841), .ZN(n7842) );
  AOI21_X1 U9440 ( .B1(n10295), .B2(n9757), .A(n7842), .ZN(n7843) );
  OAI21_X1 U9441 ( .B1(n7844), .B2(n9759), .A(n7843), .ZN(P1_U3281) );
  INV_X1 U9442 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7848) );
  NOR2_X1 U9443 ( .A1(n7848), .A2(n7847), .ZN(n9370) );
  AOI211_X1 U9444 ( .C1(n7848), .C2(n7847), .A(n9370), .B(n9415), .ZN(n7858)
         );
  OR2_X1 U9445 ( .A1(n7850), .A2(n7849), .ZN(n7851) );
  OAI21_X1 U9446 ( .B1(n10314), .B2(n7852), .A(n7851), .ZN(n9361) );
  XNOR2_X1 U9447 ( .A(n9368), .B(n9361), .ZN(n7853) );
  NAND2_X1 U9448 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n7853), .ZN(n9363) );
  OAI211_X1 U9449 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n7853), .A(n9436), .B(
        n9363), .ZN(n7856) );
  NOR2_X1 U9450 ( .A1(n7854), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9302) );
  AOI21_X1 U9451 ( .B1(n9420), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n9302), .ZN(
        n7855) );
  OAI211_X1 U9452 ( .C1(n9431), .C2(n9368), .A(n7856), .B(n7855), .ZN(n7857)
         );
  OR2_X1 U9453 ( .A1(n7858), .A2(n7857), .ZN(P1_U3258) );
  AOI211_X1 U9454 ( .C1(n7862), .C2(n7861), .A(n7860), .B(n7859), .ZN(n7867)
         );
  AOI22_X1 U9455 ( .A1(n8028), .A2(n7863), .B1(n10313), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n7864) );
  OAI21_X1 U9456 ( .B1(n7867), .B2(n10313), .A(n7864), .ZN(P1_U3533) );
  AOI22_X1 U9457 ( .A1(n8028), .A2(n7865), .B1(n10304), .B2(
        P1_REG0_REG_11__SCAN_IN), .ZN(n7866) );
  OAI21_X1 U9458 ( .B1(n7867), .B2(n10304), .A(n7866), .ZN(P1_U3486) );
  INV_X1 U9459 ( .A(n8085), .ZN(n7883) );
  INV_X1 U9460 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7937) );
  AOI21_X1 U9461 ( .B1(n7868), .B2(n7937), .A(n8082), .ZN(n7886) );
  XOR2_X1 U9462 ( .A(n8085), .B(n8086), .Z(n7872) );
  NAND2_X1 U9463 ( .A1(n7873), .A2(n7872), .ZN(n8087) );
  OAI21_X1 U9464 ( .B1(n7873), .B2(n7872), .A(n8087), .ZN(n7874) );
  NAND2_X1 U9465 ( .A1(n7874), .A2(n8628), .ZN(n7885) );
  NAND2_X1 U9466 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8066) );
  OAI21_X1 U9467 ( .B1(n10330), .B2(n7610), .A(n8066), .ZN(n7882) );
  INV_X1 U9468 ( .A(n7875), .ZN(n7877) );
  OAI21_X1 U9469 ( .B1(n7877), .B2(n9968), .A(n7876), .ZN(n7878) );
  OAI21_X1 U9470 ( .B1(n7878), .B2(n8085), .A(n8079), .ZN(n7879) );
  INV_X1 U9471 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9855) );
  AOI21_X1 U9472 ( .B1(n7879), .B2(n9855), .A(n8075), .ZN(n7880) );
  NOR2_X1 U9473 ( .A1(n7880), .A2(n8634), .ZN(n7881) );
  AOI211_X1 U9474 ( .C1(n10332), .C2(n7883), .A(n7882), .B(n7881), .ZN(n7884)
         );
  OAI211_X1 U9475 ( .C1(n7886), .C2(n8602), .A(n7885), .B(n7884), .ZN(P2_U3191) );
  NOR2_X1 U9476 ( .A1(n10353), .A2(n10342), .ZN(n7983) );
  INV_X1 U9477 ( .A(n7983), .ZN(n7941) );
  INV_X1 U9478 ( .A(n7887), .ZN(n7889) );
  INV_X1 U9479 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7888) );
  MUX2_X1 U9480 ( .A(n7889), .B(n7888), .S(n10353), .Z(n7892) );
  AOI22_X1 U9481 ( .A1(n8795), .A2(n7890), .B1(n8822), .B2(n7905), .ZN(n7891)
         );
  OAI211_X1 U9482 ( .C1(n7893), .C2(n7941), .A(n7892), .B(n7891), .ZN(P2_U3226) );
  XNOR2_X1 U9483 ( .A(n4406), .B(n7902), .ZN(n7949) );
  XNOR2_X1 U9484 ( .A(n7949), .B(n8402), .ZN(n7899) );
  INV_X1 U9485 ( .A(n8403), .ZN(n7901) );
  INV_X1 U9486 ( .A(n7951), .ZN(n7897) );
  AOI21_X1 U9487 ( .B1(n7899), .B2(n7898), .A(n7897), .ZN(n7908) );
  INV_X1 U9488 ( .A(n7900), .ZN(n7904) );
  OAI22_X1 U9489 ( .A1(n7902), .A2(n8384), .B1(n8358), .B2(n7901), .ZN(n7903)
         );
  AOI211_X1 U9490 ( .C1(n8355), .C2(n8401), .A(n7904), .B(n7903), .ZN(n7907)
         );
  NAND2_X1 U9491 ( .A1(n8381), .A2(n7905), .ZN(n7906) );
  OAI211_X1 U9492 ( .C1(n7908), .C2(n8373), .A(n7907), .B(n7906), .ZN(P2_U3153) );
  NAND2_X1 U9493 ( .A1(n7814), .A2(n7909), .ZN(n7910) );
  XOR2_X1 U9494 ( .A(n7929), .B(n7910), .Z(n7948) );
  OAI22_X1 U9495 ( .A1(n7948), .A2(n8912), .B1(n7956), .B2(n8917), .ZN(n7913)
         );
  INV_X1 U9496 ( .A(n8400), .ZN(n8138) );
  XNOR2_X1 U9497 ( .A(n7911), .B(n7929), .ZN(n7912) );
  OAI222_X1 U9498 ( .A1(n8899), .A2(n8138), .B1(n8901), .B2(n7955), .C1(n7912), 
        .C2(n8896), .ZN(n7942) );
  NOR2_X1 U9499 ( .A1(n7913), .A2(n7942), .ZN(n10364) );
  NAND2_X1 U9500 ( .A1(n8924), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7914) );
  OAI21_X1 U9501 ( .B1(n10364), .B2(n8924), .A(n7914), .ZN(P2_U3467) );
  INV_X1 U9502 ( .A(n7925), .ZN(n7917) );
  AOI21_X1 U9503 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n10215), .A(n7915), .ZN(
        n7916) );
  OAI21_X1 U9504 ( .B1(n7917), .B2(n10222), .A(n7916), .ZN(P1_U3332) );
  INV_X1 U9505 ( .A(n7918), .ZN(n7921) );
  OAI222_X1 U9506 ( .A1(n10225), .A2(n7920), .B1(n10222), .B2(n7921), .C1(
        P1_U3086), .C2(n7919), .ZN(P1_U3333) );
  OAI222_X1 U9507 ( .A1(n7923), .A2(P2_U3151), .B1(n7922), .B2(n7921), .C1(
        n9990), .C2(n8987), .ZN(P2_U3273) );
  NAND2_X1 U9508 ( .A1(n7925), .A2(n7924), .ZN(n7927) );
  OAI211_X1 U9509 ( .C1(n9991), .C2(n8987), .A(n7927), .B(n7926), .ZN(P2_U3272) );
  XNOR2_X1 U9510 ( .A(n7928), .B(n7932), .ZN(n7965) );
  NAND2_X1 U9511 ( .A1(n7911), .A2(n7929), .ZN(n7990) );
  NAND2_X1 U9512 ( .A1(n7990), .A2(n7930), .ZN(n7931) );
  XOR2_X1 U9513 ( .A(n7932), .B(n7931), .Z(n7933) );
  NAND2_X1 U9514 ( .A1(n7933), .A2(n8785), .ZN(n7935) );
  AOI22_X1 U9515 ( .A1(n8780), .A2(n8399), .B1(n8401), .B2(n8782), .ZN(n7934)
         );
  OAI211_X1 U9516 ( .C1(n7979), .C2(n7965), .A(n7935), .B(n7934), .ZN(n7967)
         );
  NAND2_X1 U9517 ( .A1(n7967), .A2(n10350), .ZN(n7940) );
  INV_X1 U9518 ( .A(n7936), .ZN(n8069) );
  OAI22_X1 U9519 ( .A1(n10350), .A2(n7937), .B1(n8069), .B2(n10345), .ZN(n7938) );
  AOI21_X1 U9520 ( .B1(n8795), .B2(n8072), .A(n7938), .ZN(n7939) );
  OAI211_X1 U9521 ( .C1(n7965), .C2(n7941), .A(n7940), .B(n7939), .ZN(P2_U3224) );
  INV_X1 U9522 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7944) );
  INV_X1 U9523 ( .A(n7942), .ZN(n7943) );
  MUX2_X1 U9524 ( .A(n7944), .B(n7943), .S(n10350), .Z(n7947) );
  AOI22_X1 U9525 ( .A1(n8795), .A2(n7945), .B1(n8822), .B2(n7959), .ZN(n7946)
         );
  OAI211_X1 U9526 ( .C1(n7948), .C2(n8792), .A(n7947), .B(n7946), .ZN(P2_U3225) );
  OR2_X1 U9527 ( .A1(n7949), .A2(n8402), .ZN(n7950) );
  XNOR2_X1 U9528 ( .A(n4406), .B(n7956), .ZN(n7952) );
  NAND2_X1 U9529 ( .A1(n7952), .A2(n8401), .ZN(n8062) );
  NAND2_X1 U9530 ( .A1(n4502), .A2(n8062), .ZN(n7953) );
  XNOR2_X1 U9531 ( .A(n8061), .B(n7953), .ZN(n7962) );
  INV_X1 U9532 ( .A(n7954), .ZN(n7958) );
  OAI22_X1 U9533 ( .A1(n7956), .A2(n8384), .B1(n8358), .B2(n7955), .ZN(n7957)
         );
  AOI211_X1 U9534 ( .C1(n8355), .C2(n8400), .A(n7958), .B(n7957), .ZN(n7961)
         );
  NAND2_X1 U9535 ( .A1(n8381), .A2(n7959), .ZN(n7960) );
  OAI211_X1 U9536 ( .C1(n7962), .C2(n8373), .A(n7961), .B(n7960), .ZN(P2_U3161) );
  OAI22_X1 U9537 ( .A1(n7965), .A2(n7964), .B1(n7963), .B2(n8917), .ZN(n7966)
         );
  NOR2_X1 U9538 ( .A1(n7967), .A2(n7966), .ZN(n10366) );
  OR2_X1 U9539 ( .A1(n8925), .A2(n9855), .ZN(n7968) );
  OAI21_X1 U9540 ( .B1(n10366), .B2(n8924), .A(n7968), .ZN(P2_U3468) );
  INV_X1 U9541 ( .A(n7975), .ZN(n7969) );
  XNOR2_X1 U9542 ( .A(n7970), .B(n7969), .ZN(n7980) );
  NAND2_X1 U9543 ( .A1(n7990), .A2(n7971), .ZN(n7973) );
  AND2_X1 U9544 ( .A1(n7973), .A2(n7972), .ZN(n7974) );
  XOR2_X1 U9545 ( .A(n7975), .B(n7974), .Z(n7976) );
  NAND2_X1 U9546 ( .A1(n7976), .A2(n8785), .ZN(n7978) );
  AOI22_X1 U9547 ( .A1(n8398), .A2(n8780), .B1(n8782), .B2(n8400), .ZN(n7977)
         );
  OAI211_X1 U9548 ( .C1(n7980), .C2(n7979), .A(n7978), .B(n7977), .ZN(n8919)
         );
  INV_X1 U9549 ( .A(n8919), .ZN(n7985) );
  INV_X1 U9550 ( .A(n7980), .ZN(n8921) );
  AOI22_X1 U9551 ( .A1(n10353), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n8822), .B2(
        n8245), .ZN(n7981) );
  OAI21_X1 U9552 ( .B1(n8918), .B2(n8810), .A(n7981), .ZN(n7982) );
  AOI21_X1 U9553 ( .B1(n8921), .B2(n7983), .A(n7982), .ZN(n7984) );
  OAI21_X1 U9554 ( .B1(n7985), .B2(n10353), .A(n7984), .ZN(P2_U3223) );
  NAND2_X1 U9555 ( .A1(n7987), .A2(n7986), .ZN(n7988) );
  XNOR2_X1 U9556 ( .A(n7988), .B(n8137), .ZN(n8913) );
  INV_X1 U9557 ( .A(n8399), .ZN(n8068) );
  NAND2_X1 U9558 ( .A1(n7990), .A2(n7989), .ZN(n7992) );
  AND2_X1 U9559 ( .A1(n7992), .A2(n7991), .ZN(n7993) );
  XNOR2_X1 U9560 ( .A(n7993), .B(n8137), .ZN(n7994) );
  OAI222_X1 U9561 ( .A1(n8901), .A2(n8068), .B1(n8899), .B2(n8900), .C1(n7994), 
        .C2(n8896), .ZN(n8915) );
  NAND2_X1 U9562 ( .A1(n8915), .A2(n10350), .ZN(n7997) );
  OAI22_X1 U9563 ( .A1(n10350), .A2(n5275), .B1(n8346), .B2(n10345), .ZN(n7995) );
  AOI21_X1 U9564 ( .B1(n8795), .B2(n8342), .A(n7995), .ZN(n7996) );
  OAI211_X1 U9565 ( .C1(n8913), .C2(n8792), .A(n7997), .B(n7996), .ZN(P2_U3222) );
  INV_X1 U9566 ( .A(n7998), .ZN(n8002) );
  AOI21_X1 U9567 ( .B1(n8000), .B2(n7999), .A(n8007), .ZN(n8001) );
  NOR2_X1 U9568 ( .A1(n8002), .A2(n8001), .ZN(n10158) );
  AOI21_X1 U9569 ( .B1(n8007), .B2(n8005), .A(n8006), .ZN(n8008) );
  INV_X1 U9570 ( .A(n8008), .ZN(n10160) );
  NAND2_X1 U9571 ( .A1(n10160), .A2(n9721), .ZN(n8016) );
  NAND2_X1 U9572 ( .A1(n9726), .A2(n10154), .ZN(n8010) );
  AOI22_X1 U9573 ( .A1(n9750), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9263), .B2(
        n9748), .ZN(n8009) );
  OAI211_X1 U9574 ( .C1(n10244), .C2(n9730), .A(n8010), .B(n8009), .ZN(n8014)
         );
  INV_X1 U9575 ( .A(n9747), .ZN(n8011) );
  OAI211_X1 U9576 ( .C1(n10210), .C2(n8012), .A(n8011), .B(n9746), .ZN(n10156)
         );
  NOR2_X1 U9577 ( .A1(n10156), .A2(n9755), .ZN(n8013) );
  AOI211_X1 U9578 ( .C1(n9751), .C2(n9012), .A(n8014), .B(n8013), .ZN(n8015)
         );
  OAI211_X1 U9579 ( .C1(n10158), .C2(n9736), .A(n8016), .B(n8015), .ZN(
        P1_U3280) );
  AOI22_X1 U9580 ( .A1(n8134), .A2(n9089), .B1(n4409), .B2(n9312), .ZN(n8020)
         );
  XOR2_X1 U9581 ( .A(n4410), .B(n8020), .Z(n8022) );
  OAI22_X1 U9582 ( .A1(n10287), .A2(n9062), .B1(n8040), .B2(n9168), .ZN(n8127)
         );
  NAND2_X1 U9583 ( .A1(n8028), .A2(n9089), .ZN(n8025) );
  NAND2_X1 U9584 ( .A1(n9311), .A2(n4409), .ZN(n8024) );
  NAND2_X1 U9585 ( .A1(n8025), .A2(n8024), .ZN(n8026) );
  XNOR2_X1 U9586 ( .A(n8026), .B(n9165), .ZN(n8029) );
  AND2_X1 U9587 ( .A1(n9311), .A2(n9115), .ZN(n8027) );
  AOI21_X1 U9588 ( .B1(n8028), .B2(n9074), .A(n8027), .ZN(n8030) );
  NAND2_X1 U9589 ( .A1(n8029), .A2(n8030), .ZN(n9198) );
  INV_X1 U9590 ( .A(n8029), .ZN(n8032) );
  INV_X1 U9591 ( .A(n8030), .ZN(n8031) );
  NAND2_X1 U9592 ( .A1(n8032), .A2(n8031), .ZN(n8033) );
  AND2_X1 U9593 ( .A1(n9198), .A2(n8033), .ZN(n8034) );
  INV_X1 U9594 ( .A(n9006), .ZN(n8037) );
  NOR3_X1 U9595 ( .A1(n8035), .A2(n8125), .A3(n8034), .ZN(n8036) );
  OAI21_X1 U9596 ( .B1(n8037), .B2(n8036), .A(n9300), .ZN(n8044) );
  AOI21_X1 U9597 ( .B1(n10154), .B2(n9295), .A(n8038), .ZN(n8039) );
  OAI21_X1 U9598 ( .B1(n8040), .B2(n9293), .A(n8039), .ZN(n8041) );
  AOI21_X1 U9599 ( .B1(n8042), .B2(n9307), .A(n8041), .ZN(n8043) );
  OAI211_X1 U9600 ( .C1(n8045), .C2(n9310), .A(n8044), .B(n8043), .ZN(P1_U3236) );
  OR2_X1 U9601 ( .A1(n8046), .A2(n8050), .ZN(n8047) );
  NAND2_X1 U9602 ( .A1(n8048), .A2(n8047), .ZN(n8904) );
  XOR2_X1 U9603 ( .A(n8050), .B(n8049), .Z(n8051) );
  OAI222_X1 U9604 ( .A1(n8901), .A2(n8249), .B1(n8899), .B2(n8819), .C1(n8896), 
        .C2(n8051), .ZN(n8905) );
  NAND2_X1 U9605 ( .A1(n8905), .A2(n10350), .ZN(n8056) );
  INV_X1 U9606 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8053) );
  INV_X1 U9607 ( .A(n8274), .ZN(n8052) );
  OAI22_X1 U9608 ( .A1(n10350), .A2(n8053), .B1(n8052), .B2(n10345), .ZN(n8054) );
  AOI21_X1 U9609 ( .B1(n8795), .B2(n8907), .A(n8054), .ZN(n8055) );
  OAI211_X1 U9610 ( .C1(n8904), .C2(n8792), .A(n8056), .B(n8055), .ZN(P2_U3221) );
  INV_X1 U9611 ( .A(n8057), .ZN(n8059) );
  OAI222_X1 U9612 ( .A1(n5677), .A2(P2_U3151), .B1(n8993), .B2(n8059), .C1(
        n9786), .C2(n8987), .ZN(P2_U3271) );
  OAI222_X1 U9613 ( .A1(n8060), .A2(P1_U3086), .B1(n10222), .B2(n8059), .C1(
        n8058), .C2(n10225), .ZN(P1_U3331) );
  XNOR2_X1 U9614 ( .A(n8201), .B(n8072), .ZN(n8139) );
  XNOR2_X1 U9615 ( .A(n8139), .B(n8400), .ZN(n8064) );
  NAND2_X1 U9616 ( .A1(n8065), .A2(n8064), .ZN(n8141) );
  OAI211_X1 U9617 ( .C1(n8065), .C2(n8064), .A(n8141), .B(n8344), .ZN(n8074)
         );
  NAND2_X1 U9618 ( .A1(n8377), .A2(n8401), .ZN(n8067) );
  OAI211_X1 U9619 ( .C1(n8379), .C2(n8068), .A(n8067), .B(n8066), .ZN(n8071)
         );
  NOR2_X1 U9620 ( .A1(n8298), .A2(n8069), .ZN(n8070) );
  AOI211_X1 U9621 ( .C1(n8072), .C2(n8367), .A(n8071), .B(n8070), .ZN(n8073)
         );
  NAND2_X1 U9622 ( .A1(n8074), .A2(n8073), .ZN(P2_U3171) );
  INV_X1 U9623 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8076) );
  MUX2_X1 U9624 ( .A(n8076), .B(P2_REG1_REG_10__SCAN_IN), .S(n8424), .Z(n8077)
         );
  AND3_X1 U9625 ( .A1(n8079), .A2(n8078), .A3(n8077), .ZN(n8080) );
  NOR2_X1 U9626 ( .A1(n8423), .A2(n8080), .ZN(n8097) );
  INV_X1 U9627 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n9811) );
  MUX2_X1 U9628 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n9811), .S(n8424), .Z(n8083)
         );
  OAI21_X1 U9629 ( .B1(n8083), .B2(n4433), .A(n8410), .ZN(n8084) );
  NAND2_X1 U9630 ( .A1(n10327), .A2(n8084), .ZN(n8093) );
  XNOR2_X1 U9631 ( .A(n8413), .B(n8424), .ZN(n8090) );
  OR2_X1 U9632 ( .A1(n8086), .A2(n8085), .ZN(n8088) );
  NAND2_X1 U9633 ( .A1(n8088), .A2(n8087), .ZN(n8089) );
  NAND2_X1 U9634 ( .A1(n8090), .A2(n8089), .ZN(n8415) );
  OAI21_X1 U9635 ( .B1(n8090), .B2(n8089), .A(n8415), .ZN(n8091) );
  AND2_X1 U9636 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8246) );
  AOI21_X1 U9637 ( .B1(n8628), .B2(n8091), .A(n8246), .ZN(n8092) );
  OAI211_X1 U9638 ( .C1(n10330), .C2(n8094), .A(n8093), .B(n8092), .ZN(n8095)
         );
  AOI21_X1 U9639 ( .B1(n8414), .B2(n10332), .A(n8095), .ZN(n8096) );
  OAI21_X1 U9640 ( .B1(n8097), .B2(n8634), .A(n8096), .ZN(P2_U3192) );
  INV_X1 U9641 ( .A(n8098), .ZN(n8102) );
  OAI222_X1 U9642 ( .A1(n8100), .A2(P1_U3086), .B1(n10222), .B2(n8102), .C1(
        n8099), .C2(n10225), .ZN(P1_U3330) );
  OAI222_X1 U9643 ( .A1(n8103), .A2(P2_U3151), .B1(n8993), .B2(n8102), .C1(
        n8101), .C2(n8987), .ZN(P2_U3270) );
  INV_X1 U9644 ( .A(n8104), .ZN(n8108) );
  OAI222_X1 U9645 ( .A1(n8106), .A2(P1_U3086), .B1(n10222), .B2(n8108), .C1(
        n8105), .C2(n10225), .ZN(P1_U3329) );
  OAI222_X1 U9646 ( .A1(n8109), .A2(P2_U3151), .B1(n8993), .B2(n8108), .C1(
        n8107), .C2(n8987), .ZN(P2_U3269) );
  INV_X1 U9647 ( .A(n8110), .ZN(n10221) );
  AOI21_X1 U9648 ( .B1(n8991), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n8111), .ZN(
        n8112) );
  OAI21_X1 U9649 ( .B1(n10221), .B2(n8993), .A(n8112), .ZN(P2_U3268) );
  INV_X1 U9650 ( .A(n8113), .ZN(n8994) );
  OAI222_X1 U9651 ( .A1(n10225), .A2(n8114), .B1(P1_U3086), .B2(n6605), .C1(
        n10222), .C2(n8994), .ZN(P1_U3327) );
  OAI222_X1 U9652 ( .A1(n10225), .A2(n8116), .B1(n10222), .B2(n8115), .C1(
        P1_U3086), .C2(n4408), .ZN(P1_U3336) );
  AOI21_X1 U9653 ( .B1(n8119), .B2(n8118), .A(n8117), .ZN(n8120) );
  MUX2_X1 U9654 ( .A(n6079), .B(n8120), .S(n9757), .Z(n8123) );
  AOI22_X1 U9655 ( .A1(n8121), .A2(n9733), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n9748), .ZN(n8122) );
  OAI211_X1 U9656 ( .C1(n8124), .C2(n9724), .A(n8123), .B(n8122), .ZN(P1_U3292) );
  AOI21_X1 U9657 ( .B1(n8127), .B2(n8126), .A(n8125), .ZN(n8136) );
  NAND2_X1 U9658 ( .A1(n9307), .A2(n8128), .ZN(n8131) );
  AOI21_X1 U9659 ( .B1(n9311), .B2(n9295), .A(n8129), .ZN(n8130) );
  OAI211_X1 U9660 ( .C1(n8132), .C2(n9293), .A(n8131), .B(n8130), .ZN(n8133)
         );
  AOI21_X1 U9661 ( .B1(n8134), .B2(n9283), .A(n8133), .ZN(n8135) );
  OAI21_X1 U9662 ( .B1(n8136), .B2(n9285), .A(n8135), .ZN(P1_U3217) );
  NAND2_X1 U9663 ( .A1(n8141), .A2(n8140), .ZN(n8142) );
  INV_X1 U9664 ( .A(n8244), .ZN(n8145) );
  XNOR2_X1 U9665 ( .A(n8918), .B(n4406), .ZN(n8243) );
  INV_X1 U9666 ( .A(n8243), .ZN(n8144) );
  XOR2_X1 U9667 ( .A(n8201), .B(n8907), .Z(n8271) );
  XNOR2_X1 U9668 ( .A(n8892), .B(n8201), .ZN(n8156) );
  XNOR2_X1 U9669 ( .A(n8156), .B(n8396), .ZN(n8146) );
  XNOR2_X1 U9670 ( .A(n8159), .B(n8146), .ZN(n8152) );
  NAND2_X1 U9671 ( .A1(n8381), .A2(n10229), .ZN(n8149) );
  NOR2_X1 U9672 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8147), .ZN(n8470) );
  AOI21_X1 U9673 ( .B1(n8377), .B2(n8397), .A(n8470), .ZN(n8148) );
  OAI211_X1 U9674 ( .C1(n8898), .C2(n8379), .A(n8149), .B(n8148), .ZN(n8150)
         );
  AOI21_X1 U9675 ( .B1(n8892), .B2(n8367), .A(n8150), .ZN(n8151) );
  OAI21_X1 U9676 ( .B1(n8152), .B2(n8373), .A(n8151), .ZN(P2_U3174) );
  INV_X1 U9677 ( .A(n8154), .ZN(n8217) );
  OAI222_X1 U9678 ( .A1(n8153), .A2(P2_U3151), .B1(n8993), .B2(n8217), .C1(
        n8155), .C2(n8987), .ZN(P2_U3265) );
  NOR2_X1 U9679 ( .A1(n8156), .A2(n8819), .ZN(n8158) );
  INV_X1 U9680 ( .A(n8156), .ZN(n8157) );
  OAI22_X1 U9681 ( .A1(n8159), .A2(n8158), .B1(n8157), .B2(n8396), .ZN(n8227)
         );
  XNOR2_X1 U9682 ( .A(n8885), .B(n4406), .ZN(n8160) );
  XNOR2_X1 U9683 ( .A(n8160), .B(n8395), .ZN(n8228) );
  NAND2_X1 U9684 ( .A1(n8227), .A2(n8228), .ZN(n8162) );
  NAND2_X1 U9685 ( .A1(n8160), .A2(n8898), .ZN(n8161) );
  NAND2_X1 U9686 ( .A1(n8162), .A2(n8161), .ZN(n8372) );
  INV_X1 U9687 ( .A(n8372), .ZN(n8164) );
  XNOR2_X1 U9688 ( .A(n8371), .B(n8201), .ZN(n8165) );
  XNOR2_X1 U9689 ( .A(n8165), .B(n8818), .ZN(n8374) );
  INV_X1 U9690 ( .A(n8165), .ZN(n8166) );
  NAND2_X1 U9691 ( .A1(n8166), .A2(n8783), .ZN(n8167) );
  XNOR2_X1 U9692 ( .A(n8877), .B(n4406), .ZN(n8168) );
  XNOR2_X1 U9693 ( .A(n8168), .B(n8801), .ZN(n8290) );
  NAND2_X1 U9694 ( .A1(n8168), .A2(n8801), .ZN(n8300) );
  NAND2_X1 U9695 ( .A1(n8302), .A2(n8300), .ZN(n8169) );
  XNOR2_X1 U9696 ( .A(n8772), .B(n8201), .ZN(n8170) );
  XNOR2_X1 U9697 ( .A(n8170), .B(n8781), .ZN(n8299) );
  NAND2_X1 U9698 ( .A1(n8169), .A2(n8299), .ZN(n8304) );
  NAND2_X1 U9699 ( .A1(n8170), .A2(n8757), .ZN(n8171) );
  NAND2_X1 U9700 ( .A1(n8304), .A2(n8171), .ZN(n8353) );
  XNOR2_X1 U9701 ( .A(n8868), .B(n4406), .ZN(n8172) );
  XNOR2_X1 U9702 ( .A(n8172), .B(n8738), .ZN(n8354) );
  NAND2_X1 U9703 ( .A1(n8353), .A2(n8354), .ZN(n8255) );
  NAND2_X1 U9704 ( .A1(n8172), .A2(n8769), .ZN(n8254) );
  XNOR2_X1 U9705 ( .A(n8744), .B(n8201), .ZN(n8174) );
  NAND2_X1 U9706 ( .A1(n8174), .A2(n8758), .ZN(n8322) );
  XNOR2_X1 U9707 ( .A(n8729), .B(n4406), .ZN(n8178) );
  NAND2_X1 U9708 ( .A1(n8178), .A2(n8713), .ZN(n8177) );
  AND2_X1 U9709 ( .A1(n8322), .A2(n8177), .ZN(n8173) );
  AND2_X1 U9710 ( .A1(n8254), .A2(n8173), .ZN(n8176) );
  INV_X1 U9711 ( .A(n8173), .ZN(n8175) );
  XNOR2_X1 U9712 ( .A(n8174), .B(n8725), .ZN(n8320) );
  XNOR2_X1 U9713 ( .A(n8268), .B(n8201), .ZN(n8185) );
  XOR2_X1 U9714 ( .A(n8701), .B(n8185), .Z(n8264) );
  INV_X1 U9715 ( .A(n8177), .ZN(n8179) );
  XNOR2_X1 U9716 ( .A(n8178), .B(n8739), .ZN(n8325) );
  XNOR2_X1 U9717 ( .A(n8317), .B(n4406), .ZN(n8311) );
  XNOR2_X1 U9718 ( .A(n8240), .B(n8201), .ZN(n8189) );
  OAI22_X1 U9719 ( .A1(n8311), .A2(n8691), .B1(n8702), .B2(n8189), .ZN(n8182)
         );
  XNOR2_X1 U9720 ( .A(n8331), .B(n4406), .ZN(n8184) );
  INV_X1 U9721 ( .A(n8184), .ZN(n8180) );
  NAND2_X1 U9722 ( .A1(n8180), .A2(n8393), .ZN(n8236) );
  INV_X1 U9723 ( .A(n8236), .ZN(n8181) );
  NOR2_X1 U9724 ( .A1(n8182), .A2(n8181), .ZN(n8183) );
  AND2_X1 U9725 ( .A1(n8234), .A2(n8183), .ZN(n8188) );
  INV_X1 U9726 ( .A(n8183), .ZN(n8187) );
  XNOR2_X1 U9727 ( .A(n8184), .B(n8712), .ZN(n8334) );
  INV_X1 U9728 ( .A(n8334), .ZN(n8186) );
  NAND2_X1 U9729 ( .A1(n8185), .A2(n8701), .ZN(n8332) );
  AOI21_X1 U9730 ( .B1(n8262), .B2(n8188), .A(n4452), .ZN(n8193) );
  OAI21_X1 U9731 ( .B1(n8309), .B2(n8392), .A(n8391), .ZN(n8191) );
  NOR2_X1 U9732 ( .A1(n8391), .A2(n8392), .ZN(n8190) );
  AOI22_X1 U9733 ( .A1(n8311), .A2(n8191), .B1(n8190), .B2(n8189), .ZN(n8192)
         );
  NAND2_X1 U9734 ( .A1(n8193), .A2(n8192), .ZN(n8280) );
  XNOR2_X1 U9735 ( .A(n8285), .B(n8201), .ZN(n8194) );
  XOR2_X1 U9736 ( .A(n8680), .B(n8194), .Z(n8281) );
  NAND2_X1 U9737 ( .A1(n8280), .A2(n8281), .ZN(n8196) );
  NAND2_X1 U9738 ( .A1(n8194), .A2(n8680), .ZN(n8195) );
  NAND2_X1 U9739 ( .A1(n8196), .A2(n8195), .ZN(n8362) );
  XNOR2_X1 U9740 ( .A(n8940), .B(n4406), .ZN(n8197) );
  INV_X1 U9741 ( .A(n8197), .ZN(n8198) );
  NAND2_X1 U9742 ( .A1(n8198), .A2(n8671), .ZN(n8199) );
  XNOR2_X1 U9743 ( .A(n8936), .B(n4406), .ZN(n8202) );
  NAND2_X1 U9744 ( .A1(n8202), .A2(n8388), .ZN(n8204) );
  OAI21_X1 U9745 ( .B1(n8202), .B2(n8388), .A(n8204), .ZN(n8220) );
  INV_X1 U9746 ( .A(n8220), .ZN(n8203) );
  XOR2_X1 U9747 ( .A(n8201), .B(n8205), .Z(n8207) );
  XNOR2_X1 U9748 ( .A(n8208), .B(n8207), .ZN(n8215) );
  AOI22_X1 U9749 ( .A1(n8388), .A2(n8377), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8210) );
  NAND2_X1 U9750 ( .A1(n8381), .A2(n8643), .ZN(n8209) );
  OAI211_X1 U9751 ( .C1(n8211), .C2(n8379), .A(n8210), .B(n8209), .ZN(n8212)
         );
  AOI21_X1 U9752 ( .B1(n8213), .B2(n8367), .A(n8212), .ZN(n8214) );
  OAI21_X1 U9753 ( .B1(n8215), .B2(n8373), .A(n8214), .ZN(P2_U3160) );
  OAI222_X1 U9754 ( .A1(n10225), .A2(n8218), .B1(n10222), .B2(n8217), .C1(
        n8216), .C2(P1_U3086), .ZN(P1_U3325) );
  AOI21_X1 U9755 ( .B1(n8219), .B2(n8220), .A(n8373), .ZN(n8222) );
  NAND2_X1 U9756 ( .A1(n8222), .A2(n8221), .ZN(n8226) );
  AOI22_X1 U9757 ( .A1(n8377), .A2(n8389), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8223) );
  OAI21_X1 U9758 ( .B1(n8651), .B2(n8379), .A(n8223), .ZN(n8224) );
  AOI21_X1 U9759 ( .B1(n8652), .B2(n8381), .A(n8224), .ZN(n8225) );
  OAI211_X1 U9760 ( .C1(n8936), .C2(n8384), .A(n8226), .B(n8225), .ZN(P2_U3154) );
  XOR2_X1 U9761 ( .A(n8227), .B(n8228), .Z(n8233) );
  NAND2_X1 U9762 ( .A1(n8381), .A2(n8821), .ZN(n8230) );
  AOI22_X1 U9763 ( .A1(n8377), .A2(n8396), .B1(P2_REG3_REG_14__SCAN_IN), .B2(
        P2_U3151), .ZN(n8229) );
  OAI211_X1 U9764 ( .C1(n8818), .C2(n8379), .A(n8230), .B(n8229), .ZN(n8231)
         );
  AOI21_X1 U9765 ( .B1(n8885), .B2(n8367), .A(n8231), .ZN(n8232) );
  OAI21_X1 U9766 ( .B1(n8233), .B2(n8373), .A(n8232), .ZN(P2_U3155) );
  NAND2_X1 U9767 ( .A1(n8262), .A2(n8234), .ZN(n8333) );
  NAND2_X1 U9768 ( .A1(n8333), .A2(n8235), .ZN(n8336) );
  NAND2_X1 U9769 ( .A1(n8336), .A2(n8236), .ZN(n8308) );
  XNOR2_X1 U9770 ( .A(n8310), .B(n8702), .ZN(n8242) );
  NAND2_X1 U9771 ( .A1(n8381), .A2(n8694), .ZN(n8238) );
  AOI22_X1 U9772 ( .A1(n8377), .A2(n8393), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8237) );
  OAI211_X1 U9773 ( .C1(n8691), .C2(n8379), .A(n8238), .B(n8237), .ZN(n8239)
         );
  AOI21_X1 U9774 ( .B1(n8240), .B2(n8367), .A(n8239), .ZN(n8241) );
  OAI21_X1 U9775 ( .B1(n8242), .B2(n8373), .A(n8241), .ZN(P2_U3156) );
  XOR2_X1 U9776 ( .A(n8244), .B(n8243), .Z(n8253) );
  NAND2_X1 U9777 ( .A1(n8381), .A2(n8245), .ZN(n8248) );
  AOI21_X1 U9778 ( .B1(n8377), .B2(n8400), .A(n8246), .ZN(n8247) );
  OAI211_X1 U9779 ( .C1(n8249), .C2(n8379), .A(n8248), .B(n8247), .ZN(n8250)
         );
  AOI21_X1 U9780 ( .B1(n8251), .B2(n8367), .A(n8250), .ZN(n8252) );
  OAI21_X1 U9781 ( .B1(n8253), .B2(n8373), .A(n8252), .ZN(P2_U3157) );
  NAND2_X1 U9782 ( .A1(n8255), .A2(n8254), .ZN(n8321) );
  XOR2_X1 U9783 ( .A(n8320), .B(n8321), .Z(n8260) );
  AOI22_X1 U9784 ( .A1(n8355), .A2(n8739), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3151), .ZN(n8257) );
  NAND2_X1 U9785 ( .A1(n8377), .A2(n8738), .ZN(n8256) );
  OAI211_X1 U9786 ( .C1(n8298), .C2(n8742), .A(n8257), .B(n8256), .ZN(n8258)
         );
  AOI21_X1 U9787 ( .B1(n8744), .B2(n8367), .A(n8258), .ZN(n8259) );
  OAI21_X1 U9788 ( .B1(n8260), .B2(n8373), .A(n8259), .ZN(P2_U3159) );
  AND2_X1 U9789 ( .A1(n8262), .A2(n8261), .ZN(n8263) );
  XOR2_X1 U9790 ( .A(n8264), .B(n8263), .Z(n8270) );
  NAND2_X1 U9791 ( .A1(n8381), .A2(n8718), .ZN(n8266) );
  AOI22_X1 U9792 ( .A1(n8355), .A2(n8393), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8265) );
  OAI211_X1 U9793 ( .C1(n8713), .C2(n8358), .A(n8266), .B(n8265), .ZN(n8267)
         );
  AOI21_X1 U9794 ( .B1(n8268), .B2(n8367), .A(n8267), .ZN(n8269) );
  OAI21_X1 U9795 ( .B1(n8270), .B2(n8373), .A(n8269), .ZN(P2_U3163) );
  XNOR2_X1 U9796 ( .A(n8271), .B(n8900), .ZN(n8272) );
  XNOR2_X1 U9797 ( .A(n8273), .B(n8272), .ZN(n8279) );
  NAND2_X1 U9798 ( .A1(n8381), .A2(n8274), .ZN(n8276) );
  AND2_X1 U9799 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8443) );
  AOI21_X1 U9800 ( .B1(n8377), .B2(n8398), .A(n8443), .ZN(n8275) );
  OAI211_X1 U9801 ( .C1(n8819), .C2(n8379), .A(n8276), .B(n8275), .ZN(n8277)
         );
  AOI21_X1 U9802 ( .B1(n8907), .B2(n8367), .A(n8277), .ZN(n8278) );
  OAI21_X1 U9803 ( .B1(n8279), .B2(n8373), .A(n8278), .ZN(P2_U3164) );
  XOR2_X1 U9804 ( .A(n8281), .B(n8280), .Z(n8287) );
  NAND2_X1 U9805 ( .A1(n8381), .A2(n8673), .ZN(n8283) );
  AOI22_X1 U9806 ( .A1(n8355), .A2(n8389), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8282) );
  OAI211_X1 U9807 ( .C1(n8691), .C2(n8358), .A(n8283), .B(n8282), .ZN(n8284)
         );
  AOI21_X1 U9808 ( .B1(n8285), .B2(n8367), .A(n8284), .ZN(n8286) );
  OAI21_X1 U9809 ( .B1(n8287), .B2(n8373), .A(n8286), .ZN(P2_U3165) );
  INV_X1 U9810 ( .A(n8302), .ZN(n8288) );
  AOI21_X1 U9811 ( .B1(n8290), .B2(n8289), .A(n8288), .ZN(n8295) );
  AOI22_X1 U9812 ( .A1(n8355), .A2(n8781), .B1(P2_REG3_REG_16__SCAN_IN), .B2(
        P2_U3151), .ZN(n8292) );
  NAND2_X1 U9813 ( .A1(n8377), .A2(n8783), .ZN(n8291) );
  OAI211_X1 U9814 ( .C1(n8298), .C2(n8786), .A(n8292), .B(n8291), .ZN(n8293)
         );
  AOI21_X1 U9815 ( .B1(n8877), .B2(n8367), .A(n8293), .ZN(n8294) );
  OAI21_X1 U9816 ( .B1(n8295), .B2(n8373), .A(n8294), .ZN(P2_U3166) );
  AND2_X1 U9817 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8567) );
  NOR2_X1 U9818 ( .A1(n8379), .A2(n8769), .ZN(n8296) );
  AOI211_X1 U9819 ( .C1(n8377), .C2(n8394), .A(n8567), .B(n8296), .ZN(n8297)
         );
  OAI21_X1 U9820 ( .B1(n8773), .B2(n8298), .A(n8297), .ZN(n8306) );
  INV_X1 U9821 ( .A(n8299), .ZN(n8301) );
  NAND3_X1 U9822 ( .A1(n8302), .A2(n8301), .A3(n8300), .ZN(n8303) );
  AOI21_X1 U9823 ( .B1(n8304), .B2(n8303), .A(n8373), .ZN(n8305) );
  AOI211_X1 U9824 ( .C1(n8772), .C2(n8367), .A(n8306), .B(n8305), .ZN(n8307)
         );
  INV_X1 U9825 ( .A(n8307), .ZN(P2_U3168) );
  OAI22_X1 U9826 ( .A1(n8310), .A2(n8392), .B1(n8309), .B2(n8308), .ZN(n8313)
         );
  XNOR2_X1 U9827 ( .A(n8311), .B(n8691), .ZN(n8312) );
  XNOR2_X1 U9828 ( .A(n8313), .B(n8312), .ZN(n8319) );
  NAND2_X1 U9829 ( .A1(n8381), .A2(n8682), .ZN(n8315) );
  INV_X1 U9830 ( .A(n8680), .ZN(n8390) );
  AOI22_X1 U9831 ( .A1(n8355), .A2(n8390), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8314) );
  OAI211_X1 U9832 ( .C1(n8702), .C2(n8358), .A(n8315), .B(n8314), .ZN(n8316)
         );
  AOI21_X1 U9833 ( .B1(n8317), .B2(n8367), .A(n8316), .ZN(n8318) );
  OAI21_X1 U9834 ( .B1(n8319), .B2(n8373), .A(n8318), .ZN(P2_U3169) );
  NAND2_X1 U9835 ( .A1(n8321), .A2(n8320), .ZN(n8323) );
  NAND2_X1 U9836 ( .A1(n8323), .A2(n8322), .ZN(n8324) );
  XOR2_X1 U9837 ( .A(n8325), .B(n8324), .Z(n8330) );
  NAND2_X1 U9838 ( .A1(n8381), .A2(n8730), .ZN(n8327) );
  AOI22_X1 U9839 ( .A1(n8355), .A2(n4641), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8326) );
  OAI211_X1 U9840 ( .C1(n8758), .C2(n8358), .A(n8327), .B(n8326), .ZN(n8328)
         );
  AOI21_X1 U9841 ( .B1(n8729), .B2(n8367), .A(n8328), .ZN(n8329) );
  OAI21_X1 U9842 ( .B1(n8330), .B2(n8373), .A(n8329), .ZN(P2_U3173) );
  INV_X1 U9843 ( .A(n8331), .ZN(n8955) );
  NAND2_X1 U9844 ( .A1(n8333), .A2(n8332), .ZN(n8335) );
  AOI21_X1 U9845 ( .B1(n8335), .B2(n8334), .A(n8373), .ZN(n8337) );
  NAND2_X1 U9846 ( .A1(n8337), .A2(n8336), .ZN(n8341) );
  AOI22_X1 U9847 ( .A1(n8377), .A2(n4641), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8338) );
  OAI21_X1 U9848 ( .B1(n8702), .B2(n8379), .A(n8338), .ZN(n8339) );
  AOI21_X1 U9849 ( .B1(n8705), .B2(n8381), .A(n8339), .ZN(n8340) );
  OAI211_X1 U9850 ( .C1(n8955), .C2(n8384), .A(n8341), .B(n8340), .ZN(P2_U3175) );
  INV_X1 U9851 ( .A(n8342), .ZN(n8911) );
  OAI211_X1 U9852 ( .C1(n8345), .C2(n5021), .A(n8344), .B(n8343), .ZN(n8352)
         );
  INV_X1 U9853 ( .A(n8346), .ZN(n8350) );
  INV_X1 U9854 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8347) );
  NOR2_X1 U9855 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8347), .ZN(n8419) );
  AOI21_X1 U9856 ( .B1(n8377), .B2(n8399), .A(n8419), .ZN(n8348) );
  OAI21_X1 U9857 ( .B1(n8900), .B2(n8379), .A(n8348), .ZN(n8349) );
  AOI21_X1 U9858 ( .B1(n8350), .B2(n8381), .A(n8349), .ZN(n8351) );
  OAI211_X1 U9859 ( .C1(n8911), .C2(n8384), .A(n8352), .B(n8351), .ZN(P2_U3176) );
  XOR2_X1 U9860 ( .A(n8354), .B(n8353), .Z(n8361) );
  NAND2_X1 U9861 ( .A1(n8381), .A2(n8759), .ZN(n8357) );
  AND2_X1 U9862 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8593) );
  AOI21_X1 U9863 ( .B1(n8355), .B2(n8725), .A(n8593), .ZN(n8356) );
  OAI211_X1 U9864 ( .C1(n8757), .C2(n8358), .A(n8357), .B(n8356), .ZN(n8359)
         );
  AOI21_X1 U9865 ( .B1(n8868), .B2(n8367), .A(n8359), .ZN(n8360) );
  OAI21_X1 U9866 ( .B1(n8361), .B2(n8373), .A(n8360), .ZN(P2_U3178) );
  XOR2_X1 U9867 ( .A(n8363), .B(n8362), .Z(n8370) );
  NAND2_X1 U9868 ( .A1(n8381), .A2(n8664), .ZN(n8365) );
  AOI22_X1 U9869 ( .A1(n8377), .A2(n8390), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8364) );
  OAI211_X1 U9870 ( .C1(n8661), .C2(n8379), .A(n8365), .B(n8364), .ZN(n8366)
         );
  AOI21_X1 U9871 ( .B1(n8368), .B2(n8367), .A(n8366), .ZN(n8369) );
  OAI21_X1 U9872 ( .B1(n8370), .B2(n8373), .A(n8369), .ZN(P2_U3180) );
  INV_X1 U9873 ( .A(n8371), .ZN(n8976) );
  AOI21_X1 U9874 ( .B1(n8372), .B2(n8374), .A(n8373), .ZN(n8376) );
  NAND2_X1 U9875 ( .A1(n8376), .A2(n8375), .ZN(n8383) );
  NAND2_X1 U9876 ( .A1(n8377), .A2(n8395), .ZN(n8378) );
  NAND2_X1 U9877 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8516) );
  OAI211_X1 U9878 ( .C1(n8379), .C2(n8801), .A(n8378), .B(n8516), .ZN(n8380)
         );
  AOI21_X1 U9879 ( .B1(n8381), .B2(n8808), .A(n8380), .ZN(n8382) );
  OAI211_X1 U9880 ( .C1(n8976), .C2(n8384), .A(n8383), .B(n8382), .ZN(P2_U3181) );
  MUX2_X1 U9881 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8638), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U9882 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8385), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U9883 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8386), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U9884 ( .A(n8387), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8592), .Z(
        P2_U3519) );
  MUX2_X1 U9885 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8388), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9886 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8389), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U9887 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8390), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9888 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8391), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9889 ( .A(n8392), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8592), .Z(
        P2_U3514) );
  MUX2_X1 U9890 ( .A(n8393), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8592), .Z(
        P2_U3513) );
  MUX2_X1 U9891 ( .A(n4641), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8592), .Z(
        P2_U3512) );
  MUX2_X1 U9892 ( .A(n8739), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8592), .Z(
        P2_U3511) );
  MUX2_X1 U9893 ( .A(n8725), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8592), .Z(
        P2_U3510) );
  MUX2_X1 U9894 ( .A(n8738), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8592), .Z(
        P2_U3509) );
  MUX2_X1 U9895 ( .A(n8781), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8592), .Z(
        P2_U3508) );
  MUX2_X1 U9896 ( .A(n8394), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8592), .Z(
        P2_U3507) );
  MUX2_X1 U9897 ( .A(n8783), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8592), .Z(
        P2_U3506) );
  MUX2_X1 U9898 ( .A(n8395), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8592), .Z(
        P2_U3505) );
  MUX2_X1 U9899 ( .A(n8396), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8592), .Z(
        P2_U3504) );
  MUX2_X1 U9900 ( .A(n8397), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8592), .Z(
        P2_U3503) );
  MUX2_X1 U9901 ( .A(n8398), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8592), .Z(
        P2_U3502) );
  MUX2_X1 U9902 ( .A(n8399), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8592), .Z(
        P2_U3501) );
  MUX2_X1 U9903 ( .A(n8400), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8592), .Z(
        P2_U3500) );
  MUX2_X1 U9904 ( .A(n8401), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8592), .Z(
        P2_U3499) );
  MUX2_X1 U9905 ( .A(n8402), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8592), .Z(
        P2_U3498) );
  MUX2_X1 U9906 ( .A(n8403), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8592), .Z(
        P2_U3497) );
  MUX2_X1 U9907 ( .A(n8404), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8592), .Z(
        P2_U3496) );
  MUX2_X1 U9908 ( .A(n8405), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8592), .Z(
        P2_U3495) );
  MUX2_X1 U9909 ( .A(n8406), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8592), .Z(
        P2_U3494) );
  MUX2_X1 U9910 ( .A(n8407), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8592), .Z(
        P2_U3493) );
  MUX2_X1 U9911 ( .A(n7304), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8592), .Z(
        P2_U3492) );
  MUX2_X1 U9912 ( .A(n8408), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8592), .Z(
        P2_U3491) );
  NAND2_X1 U9913 ( .A1(n8424), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n8409) );
  AOI21_X1 U9914 ( .B1(n5275), .B2(n8412), .A(n8433), .ZN(n8430) );
  XNOR2_X1 U9915 ( .A(n8437), .B(n8448), .ZN(n8418) );
  NAND2_X1 U9916 ( .A1(n8414), .A2(n8413), .ZN(n8416) );
  NAND2_X1 U9917 ( .A1(n8416), .A2(n8415), .ZN(n8417) );
  NAND2_X1 U9918 ( .A1(n8418), .A2(n8417), .ZN(n8439) );
  OAI21_X1 U9919 ( .B1(n8418), .B2(n8417), .A(n8439), .ZN(n8420) );
  AOI21_X1 U9920 ( .B1(n8628), .B2(n8420), .A(n8419), .ZN(n8421) );
  OAI21_X1 U9921 ( .B1(n10330), .B2(n8422), .A(n8421), .ZN(n8428) );
  XNOR2_X1 U9922 ( .A(n8447), .B(n8448), .ZN(n8425) );
  NOR2_X1 U9923 ( .A1(n8426), .A2(n8634), .ZN(n8427) );
  AOI211_X1 U9924 ( .C1(n10332), .C2(n8448), .A(n8428), .B(n8427), .ZN(n8429)
         );
  OAI21_X1 U9925 ( .B1(n8430), .B2(n8602), .A(n8429), .ZN(P2_U3193) );
  NOR2_X1 U9926 ( .A1(n8448), .A2(n8432), .ZN(n8434) );
  NAND2_X1 U9927 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n8466), .ZN(n8435) );
  OAI21_X1 U9928 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n8466), .A(n8435), .ZN(
        n8436) );
  AOI21_X1 U9929 ( .B1(n4496), .B2(n8436), .A(n8458), .ZN(n8457) );
  XNOR2_X1 U9930 ( .A(n8460), .B(n8455), .ZN(n8442) );
  INV_X1 U9931 ( .A(n8437), .ZN(n8438) );
  NAND2_X1 U9932 ( .A1(n8448), .A2(n8438), .ZN(n8440) );
  NAND2_X1 U9933 ( .A1(n8440), .A2(n8439), .ZN(n8441) );
  NAND2_X1 U9934 ( .A1(n8442), .A2(n8441), .ZN(n8461) );
  OAI21_X1 U9935 ( .B1(n8442), .B2(n8441), .A(n8461), .ZN(n8444) );
  AOI21_X1 U9936 ( .B1(n8628), .B2(n8444), .A(n8443), .ZN(n8445) );
  OAI21_X1 U9937 ( .B1(n10330), .B2(n8446), .A(n8445), .ZN(n8454) );
  NAND2_X1 U9938 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n8466), .ZN(n8449) );
  OAI21_X1 U9939 ( .B1(n8466), .B2(P2_REG1_REG_12__SCAN_IN), .A(n8449), .ZN(
        n8450) );
  NOR2_X1 U9940 ( .A1(n8451), .A2(n8450), .ZN(n8465) );
  AOI21_X1 U9941 ( .B1(n8451), .B2(n8450), .A(n8465), .ZN(n8452) );
  NOR2_X1 U9942 ( .A1(n8452), .A2(n8634), .ZN(n8453) );
  AOI211_X1 U9943 ( .C1(n10332), .C2(n8455), .A(n8454), .B(n8453), .ZN(n8456)
         );
  OAI21_X1 U9944 ( .B1(n8457), .B2(n8602), .A(n8456), .ZN(P2_U3194) );
  INV_X1 U9945 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10238) );
  XNOR2_X1 U9946 ( .A(n8492), .B(n8493), .ZN(n8459) );
  AOI21_X1 U9947 ( .B1(n10238), .B2(n8459), .A(n8494), .ZN(n8475) );
  XNOR2_X1 U9948 ( .A(n8483), .B(n8493), .ZN(n8464) );
  OR2_X1 U9949 ( .A1(n8460), .A2(n8466), .ZN(n8462) );
  NAND2_X1 U9950 ( .A1(n8462), .A2(n8461), .ZN(n8463) );
  OAI21_X1 U9951 ( .B1(n8464), .B2(n8463), .A(n8485), .ZN(n8471) );
  AOI21_X1 U9952 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n8466), .A(n8465), .ZN(
        n8476) );
  INV_X1 U9953 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8903) );
  AOI21_X1 U9954 ( .B1(n8467), .B2(n8903), .A(n8477), .ZN(n8468) );
  NOR2_X1 U9955 ( .A1(n8634), .A2(n8468), .ZN(n8469) );
  AOI211_X1 U9956 ( .C1(n8628), .C2(n8471), .A(n8470), .B(n8469), .ZN(n8472)
         );
  OAI21_X1 U9957 ( .B1(n9951), .B2(n10330), .A(n8472), .ZN(n8473) );
  AOI21_X1 U9958 ( .B1(n8493), .B2(n10332), .A(n8473), .ZN(n8474) );
  OAI21_X1 U9959 ( .B1(n8475), .B2(n8602), .A(n8474), .ZN(P2_U3195) );
  NOR2_X1 U9960 ( .A1(n8493), .A2(n8476), .ZN(n8478) );
  NAND2_X1 U9961 ( .A1(n8510), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8506) );
  INV_X1 U9962 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8888) );
  NAND2_X1 U9963 ( .A1(n8503), .A2(n8888), .ZN(n8479) );
  NAND2_X1 U9964 ( .A1(n8506), .A2(n8479), .ZN(n8481) );
  INV_X1 U9965 ( .A(n8507), .ZN(n8480) );
  AOI21_X1 U9966 ( .B1(n8482), .B2(n8481), .A(n8480), .ZN(n8505) );
  XNOR2_X1 U9967 ( .A(n8511), .B(n8503), .ZN(n8488) );
  INV_X1 U9968 ( .A(n8483), .ZN(n8484) );
  NAND2_X1 U9969 ( .A1(n8493), .A2(n8484), .ZN(n8486) );
  NAND2_X1 U9970 ( .A1(n8486), .A2(n8485), .ZN(n8487) );
  NAND2_X1 U9971 ( .A1(n8488), .A2(n8487), .ZN(n8512) );
  OAI21_X1 U9972 ( .B1(n8488), .B2(n8487), .A(n8512), .ZN(n8490) );
  AND2_X1 U9973 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8489) );
  AOI21_X1 U9974 ( .B1(n8628), .B2(n8490), .A(n8489), .ZN(n8491) );
  OAI21_X1 U9975 ( .B1(n10330), .B2(n9772), .A(n8491), .ZN(n8502) );
  NOR2_X1 U9976 ( .A1(n8493), .A2(n8492), .ZN(n8495) );
  NAND2_X1 U9977 ( .A1(n8510), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8521) );
  INV_X1 U9978 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8496) );
  NAND2_X1 U9979 ( .A1(n8503), .A2(n8496), .ZN(n8497) );
  NAND2_X1 U9980 ( .A1(n8521), .A2(n8497), .ZN(n8498) );
  NAND2_X1 U9981 ( .A1(n8499), .A2(n8498), .ZN(n8500) );
  AOI21_X1 U9982 ( .B1(n8522), .B2(n8500), .A(n8602), .ZN(n8501) );
  AOI211_X1 U9983 ( .C1(n10332), .C2(n8503), .A(n8502), .B(n8501), .ZN(n8504)
         );
  OAI21_X1 U9984 ( .B1(n8505), .B2(n8634), .A(n8504), .ZN(P2_U3196) );
  NAND2_X1 U9985 ( .A1(n8507), .A2(n8506), .ZN(n8530) );
  INV_X1 U9986 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8883) );
  AOI21_X1 U9987 ( .B1(n8508), .B2(n8883), .A(n8532), .ZN(n8529) );
  INV_X1 U9988 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8509) );
  XNOR2_X1 U9989 ( .A(n8537), .B(n8523), .ZN(n8515) );
  OR2_X1 U9990 ( .A1(n8511), .A2(n8510), .ZN(n8513) );
  NAND2_X1 U9991 ( .A1(n8513), .A2(n8512), .ZN(n8514) );
  NAND2_X1 U9992 ( .A1(n8515), .A2(n8514), .ZN(n8538) );
  OAI21_X1 U9993 ( .B1(n8515), .B2(n8514), .A(n8538), .ZN(n8518) );
  INV_X1 U9994 ( .A(n8516), .ZN(n8517) );
  AOI21_X1 U9995 ( .B1(n8628), .B2(n8518), .A(n8517), .ZN(n8519) );
  OAI21_X1 U9996 ( .B1(n10330), .B2(n8520), .A(n8519), .ZN(n8527) );
  AOI21_X1 U9997 ( .B1(n8509), .B2(n8524), .A(n8549), .ZN(n8525) );
  NOR2_X1 U9998 ( .A1(n8525), .A2(n8602), .ZN(n8526) );
  AOI211_X1 U9999 ( .C1(n10332), .C2(n8548), .A(n8527), .B(n8526), .ZN(n8528)
         );
  OAI21_X1 U10000 ( .B1(n8529), .B2(n8634), .A(n8528), .ZN(P2_U3197) );
  INV_X1 U10001 ( .A(n8530), .ZN(n8531) );
  NOR2_X1 U10002 ( .A1(n8548), .A2(n8531), .ZN(n8533) );
  XNOR2_X1 U10003 ( .A(n8556), .B(n8534), .ZN(n8535) );
  AOI21_X1 U10004 ( .B1(n8536), .B2(n8535), .A(n8559), .ZN(n8558) );
  INV_X1 U10005 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8545) );
  NAND2_X1 U10006 ( .A1(n8537), .A2(n8548), .ZN(n8539) );
  NAND2_X1 U10007 ( .A1(n8539), .A2(n8538), .ZN(n8541) );
  XNOR2_X1 U10008 ( .A(n8562), .B(n8556), .ZN(n8540) );
  NAND2_X1 U10009 ( .A1(n8540), .A2(n8541), .ZN(n8563) );
  OAI21_X1 U10010 ( .B1(n8541), .B2(n8540), .A(n8563), .ZN(n8543) );
  INV_X1 U10011 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10032) );
  NOR2_X1 U10012 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10032), .ZN(n8542) );
  AOI21_X1 U10013 ( .B1(n8628), .B2(n8543), .A(n8542), .ZN(n8544) );
  OAI21_X1 U10014 ( .B1(n10330), .B2(n8545), .A(n8544), .ZN(n8555) );
  NOR2_X1 U10015 ( .A1(n8548), .A2(n8547), .ZN(n8550) );
  NOR2_X1 U10016 ( .A1(n8550), .A2(n8549), .ZN(n8552) );
  AOI22_X1 U10017 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8556), .B1(n8572), .B2(
        n8787), .ZN(n8551) );
  AOI21_X1 U10018 ( .B1(n8552), .B2(n8551), .A(n8571), .ZN(n8553) );
  NOR2_X1 U10019 ( .A1(n8553), .A2(n8602), .ZN(n8554) );
  AOI211_X1 U10020 ( .C1(n10332), .C2(n8556), .A(n8555), .B(n8554), .ZN(n8557)
         );
  OAI21_X1 U10021 ( .B1(n8558), .B2(n8634), .A(n8557), .ZN(P2_U3198) );
  AOI21_X1 U10022 ( .B1(n8875), .B2(n8560), .A(n8580), .ZN(n8578) );
  INV_X1 U10023 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8570) );
  XNOR2_X1 U10024 ( .A(n8586), .B(n8561), .ZN(n8566) );
  OR2_X1 U10025 ( .A1(n8562), .A2(n8572), .ZN(n8564) );
  NAND2_X1 U10026 ( .A1(n8564), .A2(n8563), .ZN(n8565) );
  NAND2_X1 U10027 ( .A1(n8566), .A2(n8565), .ZN(n8584) );
  OAI21_X1 U10028 ( .B1(n8566), .B2(n8565), .A(n8584), .ZN(n8568) );
  AOI21_X1 U10029 ( .B1(n8628), .B2(n8568), .A(n8567), .ZN(n8569) );
  OAI21_X1 U10030 ( .B1(n10330), .B2(n8570), .A(n8569), .ZN(n8576) );
  AOI21_X1 U10031 ( .B1(n8774), .B2(n8573), .A(n8598), .ZN(n8574) );
  NOR2_X1 U10032 ( .A1(n8574), .A2(n8602), .ZN(n8575) );
  OAI21_X1 U10033 ( .B1(n8578), .B2(n8634), .A(n8577), .ZN(P2_U3199) );
  NOR2_X1 U10034 ( .A1(n8597), .A2(n8579), .ZN(n8581) );
  NOR2_X1 U10035 ( .A1(n8581), .A2(n8580), .ZN(n8583) );
  NAND2_X1 U10036 ( .A1(n8599), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8608) );
  OAI21_X1 U10037 ( .B1(n8599), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8608), .ZN(
        n8582) );
  NOR2_X1 U10038 ( .A1(n8583), .A2(n8582), .ZN(n8610) );
  AOI21_X1 U10039 ( .B1(n8583), .B2(n8582), .A(n8610), .ZN(n8607) );
  INV_X1 U10040 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8595) );
  INV_X1 U10041 ( .A(n8584), .ZN(n8585) );
  NAND2_X1 U10042 ( .A1(n8587), .A2(n8588), .ZN(n8591) );
  INV_X1 U10043 ( .A(n8587), .ZN(n8590) );
  INV_X1 U10044 ( .A(n8588), .ZN(n8589) );
  NAND2_X1 U10045 ( .A1(n8590), .A2(n8589), .ZN(n8619) );
  AOI21_X1 U10046 ( .B1(n8591), .B2(n8619), .A(n8605), .ZN(n8594) );
  NAND2_X1 U10047 ( .A1(n8599), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8613) );
  OAI21_X1 U10048 ( .B1(n8599), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8613), .ZN(
        n8600) );
  AOI21_X1 U10049 ( .B1(n8601), .B2(n8600), .A(n8615), .ZN(n8603) );
  NOR2_X1 U10050 ( .A1(n8603), .A2(n8602), .ZN(n8604) );
  OAI21_X1 U10051 ( .B1(n8607), .B2(n8634), .A(n8606), .ZN(P2_U3200) );
  INV_X1 U10052 ( .A(n8608), .ZN(n8609) );
  NOR2_X1 U10053 ( .A1(n8610), .A2(n8609), .ZN(n8612) );
  XNOR2_X1 U10054 ( .A(n8611), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8624) );
  XNOR2_X1 U10055 ( .A(n8612), .B(n8624), .ZN(n8635) );
  INV_X1 U10056 ( .A(n8613), .ZN(n8614) );
  NOR2_X1 U10057 ( .A1(n8615), .A2(n8614), .ZN(n8616) );
  XNOR2_X1 U10058 ( .A(n8617), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8621) );
  XNOR2_X1 U10059 ( .A(n8616), .B(n8621), .ZN(n8632) );
  NOR2_X1 U10060 ( .A1(n8618), .A2(n8617), .ZN(n8631) );
  NAND2_X1 U10061 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3151), .ZN(n8630) );
  NAND2_X1 U10062 ( .A1(n8620), .A2(n8619), .ZN(n8626) );
  INV_X1 U10063 ( .A(n8621), .ZN(n8623) );
  MUX2_X1 U10064 ( .A(n8624), .B(n8623), .S(n8622), .Z(n8625) );
  XNOR2_X1 U10065 ( .A(n8626), .B(n8625), .ZN(n8627) );
  NAND2_X1 U10066 ( .A1(n8628), .A2(n8627), .ZN(n8629) );
  OAI21_X1 U10067 ( .B1(n8635), .B2(n8634), .A(n8633), .ZN(P2_U3201) );
  INV_X1 U10068 ( .A(n8636), .ZN(n8637) );
  NAND2_X1 U10069 ( .A1(n8638), .A2(n8637), .ZN(n8927) );
  AOI21_X1 U10070 ( .B1(n8639), .B2(n8927), .A(n10353), .ZN(n8641) );
  AOI21_X1 U10071 ( .B1(n10353), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8641), .ZN(
        n8640) );
  OAI21_X1 U10072 ( .B1(n8929), .B2(n8810), .A(n8640), .ZN(P2_U3202) );
  AOI21_X1 U10073 ( .B1(n10353), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8641), .ZN(
        n8642) );
  OAI21_X1 U10074 ( .B1(n8932), .B2(n8810), .A(n8642), .ZN(P2_U3203) );
  AOI22_X1 U10075 ( .A1(n10353), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8643), 
        .B2(n8822), .ZN(n8644) );
  OAI21_X1 U10076 ( .B1(n4781), .B2(n8810), .A(n8644), .ZN(n8645) );
  AOI21_X1 U10077 ( .B1(n5025), .B2(n8825), .A(n8645), .ZN(n8646) );
  OAI21_X1 U10078 ( .B1(n8647), .B2(n10353), .A(n8646), .ZN(P2_U3205) );
  XNOR2_X1 U10079 ( .A(n8649), .B(n8648), .ZN(n8650) );
  OAI222_X1 U10080 ( .A1(n8901), .A2(n8671), .B1(n8899), .B2(n8651), .C1(n8896), .C2(n8650), .ZN(n8832) );
  AOI21_X1 U10081 ( .B1(n8822), .B2(n8652), .A(n8832), .ZN(n8658) );
  AOI22_X1 U10082 ( .A1(n8653), .A2(n8795), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n10353), .ZN(n8657) );
  XNOR2_X1 U10083 ( .A(n8655), .B(n8654), .ZN(n8833) );
  NAND2_X1 U10084 ( .A1(n8833), .A2(n8825), .ZN(n8656) );
  OAI211_X1 U10085 ( .C1(n8658), .C2(n10353), .A(n8657), .B(n8656), .ZN(
        P2_U3206) );
  XOR2_X1 U10086 ( .A(n8662), .B(n8659), .Z(n8660) );
  OAI222_X1 U10087 ( .A1(n8901), .A2(n8680), .B1(n8899), .B2(n8661), .C1(n8896), .C2(n8660), .ZN(n8835) );
  INV_X1 U10088 ( .A(n8835), .ZN(n8668) );
  XNOR2_X1 U10089 ( .A(n8663), .B(n8662), .ZN(n8836) );
  AOI22_X1 U10090 ( .A1(n10353), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n8822), 
        .B2(n8664), .ZN(n8665) );
  OAI21_X1 U10091 ( .B1(n8940), .B2(n8810), .A(n8665), .ZN(n8666) );
  AOI21_X1 U10092 ( .B1(n8836), .B2(n8825), .A(n8666), .ZN(n8667) );
  OAI21_X1 U10093 ( .B1(n8668), .B2(n10353), .A(n8667), .ZN(P2_U3207) );
  NOR2_X1 U10094 ( .A1(n8944), .A2(n10343), .ZN(n8672) );
  XOR2_X1 U10095 ( .A(n8674), .B(n8669), .Z(n8670) );
  OAI222_X1 U10096 ( .A1(n8901), .A2(n8691), .B1(n8899), .B2(n8671), .C1(n8896), .C2(n8670), .ZN(n8839) );
  AOI211_X1 U10097 ( .C1(n8822), .C2(n8673), .A(n8672), .B(n8839), .ZN(n8677)
         );
  XNOR2_X1 U10098 ( .A(n8675), .B(n8674), .ZN(n8840) );
  AOI22_X1 U10099 ( .A1(n8840), .A2(n8825), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n10353), .ZN(n8676) );
  OAI21_X1 U10100 ( .B1(n8677), .B2(n10353), .A(n8676), .ZN(P2_U3208) );
  NOR2_X1 U10101 ( .A1(n8948), .A2(n10343), .ZN(n8681) );
  XOR2_X1 U10102 ( .A(n8686), .B(n8678), .Z(n8679) );
  OAI222_X1 U10103 ( .A1(n8901), .A2(n8702), .B1(n8899), .B2(n8680), .C1(n8679), .C2(n8896), .ZN(n8842) );
  AOI211_X1 U10104 ( .C1(n8822), .C2(n8682), .A(n8681), .B(n8842), .ZN(n8688)
         );
  NOR2_X1 U10105 ( .A1(n8684), .A2(n8683), .ZN(n8685) );
  XOR2_X1 U10106 ( .A(n8686), .B(n8685), .Z(n8843) );
  AOI22_X1 U10107 ( .A1(n8843), .A2(n8825), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n10353), .ZN(n8687) );
  OAI21_X1 U10108 ( .B1(n8688), .B2(n10353), .A(n8687), .ZN(P2_U3209) );
  XNOR2_X1 U10109 ( .A(n8689), .B(n8693), .ZN(n8690) );
  OAI222_X1 U10110 ( .A1(n8899), .A2(n8691), .B1(n8901), .B2(n8712), .C1(n8896), .C2(n8690), .ZN(n8846) );
  INV_X1 U10111 ( .A(n8846), .ZN(n8698) );
  XOR2_X1 U10112 ( .A(n8693), .B(n8692), .Z(n8847) );
  AOI22_X1 U10113 ( .A1(n10353), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8822), 
        .B2(n8694), .ZN(n8695) );
  OAI21_X1 U10114 ( .B1(n8952), .B2(n8810), .A(n8695), .ZN(n8696) );
  AOI21_X1 U10115 ( .B1(n8847), .B2(n8825), .A(n8696), .ZN(n8697) );
  OAI21_X1 U10116 ( .B1(n8698), .B2(n10353), .A(n8697), .ZN(P2_U3210) );
  XOR2_X1 U10117 ( .A(n8703), .B(n8699), .Z(n8700) );
  OAI222_X1 U10118 ( .A1(n8899), .A2(n8702), .B1(n8901), .B2(n8701), .C1(n8896), .C2(n8700), .ZN(n8850) );
  INV_X1 U10119 ( .A(n8850), .ZN(n8709) );
  XNOR2_X1 U10120 ( .A(n8704), .B(n8703), .ZN(n8851) );
  AOI22_X1 U10121 ( .A1(n10353), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8822), 
        .B2(n8705), .ZN(n8706) );
  OAI21_X1 U10122 ( .B1(n8955), .B2(n8810), .A(n8706), .ZN(n8707) );
  AOI21_X1 U10123 ( .B1(n8851), .B2(n8825), .A(n8707), .ZN(n8708) );
  OAI21_X1 U10124 ( .B1(n8709), .B2(n10353), .A(n8708), .ZN(P2_U3211) );
  XOR2_X1 U10125 ( .A(n8717), .B(n8710), .Z(n8711) );
  OAI222_X1 U10126 ( .A1(n8901), .A2(n8713), .B1(n8899), .B2(n8712), .C1(n8896), .C2(n8711), .ZN(n8854) );
  INV_X1 U10127 ( .A(n8854), .ZN(n8722) );
  NAND2_X1 U10128 ( .A1(n8715), .A2(n8714), .ZN(n8716) );
  XOR2_X1 U10129 ( .A(n8717), .B(n8716), .Z(n8855) );
  AOI22_X1 U10130 ( .A1(n10353), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8822), 
        .B2(n8718), .ZN(n8719) );
  OAI21_X1 U10131 ( .B1(n8958), .B2(n8810), .A(n8719), .ZN(n8720) );
  AOI21_X1 U10132 ( .B1(n8855), .B2(n8825), .A(n8720), .ZN(n8721) );
  OAI21_X1 U10133 ( .B1(n8722), .B2(n10353), .A(n8721), .ZN(P2_U3212) );
  OAI21_X1 U10134 ( .B1(n8724), .B2(n8728), .A(n8723), .ZN(n8726) );
  AOI222_X1 U10135 ( .A1(n8785), .A2(n8726), .B1(n4641), .B2(n8780), .C1(n8725), .C2(n8782), .ZN(n8857) );
  XOR2_X1 U10136 ( .A(n8728), .B(n8727), .Z(n8859) );
  INV_X1 U10137 ( .A(n8729), .ZN(n8962) );
  AOI22_X1 U10138 ( .A1(n10353), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8822), 
        .B2(n8730), .ZN(n8731) );
  OAI21_X1 U10139 ( .B1(n8962), .B2(n8810), .A(n8731), .ZN(n8732) );
  AOI21_X1 U10140 ( .B1(n8859), .B2(n8825), .A(n8732), .ZN(n8733) );
  OAI21_X1 U10141 ( .B1(n8857), .B2(n10353), .A(n8733), .ZN(P2_U3213) );
  NAND2_X1 U10142 ( .A1(n8734), .A2(n8745), .ZN(n8735) );
  NAND2_X1 U10143 ( .A1(n8735), .A2(n8785), .ZN(n8736) );
  OR2_X1 U10144 ( .A1(n8737), .A2(n8736), .ZN(n8741) );
  AOI22_X1 U10145 ( .A1(n8739), .A2(n8780), .B1(n8782), .B2(n8738), .ZN(n8740)
         );
  NAND2_X1 U10146 ( .A1(n8741), .A2(n8740), .ZN(n8867) );
  INV_X1 U10147 ( .A(n8867), .ZN(n8750) );
  OAI22_X1 U10148 ( .A1(n10350), .A2(n9980), .B1(n8742), .B2(n10345), .ZN(
        n8743) );
  AOI21_X1 U10149 ( .B1(n8744), .B2(n8795), .A(n8743), .ZN(n8749) );
  INV_X1 U10150 ( .A(n8864), .ZN(n8747) );
  OR2_X1 U10151 ( .A1(n8746), .A2(n8745), .ZN(n8862) );
  NAND3_X1 U10152 ( .A1(n8747), .A2(n8825), .A3(n8862), .ZN(n8748) );
  OAI211_X1 U10153 ( .C1(n8750), .C2(n10353), .A(n8749), .B(n8748), .ZN(
        P2_U3214) );
  NAND2_X1 U10154 ( .A1(n8751), .A2(n8755), .ZN(n8752) );
  INV_X1 U10155 ( .A(n8870), .ZN(n8765) );
  XNOR2_X1 U10156 ( .A(n8754), .B(n8755), .ZN(n8756) );
  OAI222_X1 U10157 ( .A1(n8899), .A2(n8758), .B1(n8901), .B2(n8757), .C1(n8756), .C2(n8896), .ZN(n8869) );
  NAND2_X1 U10158 ( .A1(n8869), .A2(n10350), .ZN(n8764) );
  INV_X1 U10159 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8761) );
  INV_X1 U10160 ( .A(n8759), .ZN(n8760) );
  OAI22_X1 U10161 ( .A1(n10350), .A2(n8761), .B1(n8760), .B2(n10345), .ZN(
        n8762) );
  AOI21_X1 U10162 ( .B1(n8868), .B2(n8795), .A(n8762), .ZN(n8763) );
  OAI211_X1 U10163 ( .C1(n8765), .C2(n8792), .A(n8764), .B(n8763), .ZN(
        P2_U3215) );
  XNOR2_X1 U10164 ( .A(n8766), .B(n8767), .ZN(n8768) );
  OAI222_X1 U10165 ( .A1(n8901), .A2(n8801), .B1(n8899), .B2(n8769), .C1(n8768), .C2(n8896), .ZN(n8873) );
  INV_X1 U10166 ( .A(n8873), .ZN(n8778) );
  XNOR2_X1 U10167 ( .A(n8771), .B(n8770), .ZN(n8874) );
  INV_X1 U10168 ( .A(n8772), .ZN(n8971) );
  NOR2_X1 U10169 ( .A1(n8971), .A2(n8810), .ZN(n8776) );
  OAI22_X1 U10170 ( .A1(n10350), .A2(n8774), .B1(n8773), .B2(n10345), .ZN(
        n8775) );
  AOI211_X1 U10171 ( .C1(n8874), .C2(n8825), .A(n8776), .B(n8775), .ZN(n8777)
         );
  OAI21_X1 U10172 ( .B1(n8778), .B2(n10353), .A(n8777), .ZN(P2_U3216) );
  XOR2_X1 U10173 ( .A(n8779), .B(n8791), .Z(n8784) );
  AOI222_X1 U10174 ( .A1(n8785), .A2(n8784), .B1(n8783), .B2(n8782), .C1(n8781), .C2(n8780), .ZN(n8879) );
  OAI22_X1 U10175 ( .A1(n10350), .A2(n8787), .B1(n8786), .B2(n10345), .ZN(
        n8794) );
  NAND2_X1 U10176 ( .A1(n8789), .A2(n8788), .ZN(n8790) );
  AOI21_X1 U10177 ( .B1(n8791), .B2(n8790), .A(n4490), .ZN(n8880) );
  NOR2_X1 U10178 ( .A1(n8880), .A2(n8792), .ZN(n8793) );
  AOI211_X1 U10179 ( .C1(n8795), .C2(n8877), .A(n8794), .B(n8793), .ZN(n8796)
         );
  OAI21_X1 U10180 ( .B1(n10353), .B2(n8879), .A(n8796), .ZN(P2_U3217) );
  AND2_X1 U10181 ( .A1(n8798), .A2(n8797), .ZN(n8799) );
  XNOR2_X1 U10182 ( .A(n8799), .B(n8806), .ZN(n8800) );
  OAI222_X1 U10183 ( .A1(n8901), .A2(n8898), .B1(n8899), .B2(n8801), .C1(n8800), .C2(n8896), .ZN(n8881) );
  INV_X1 U10184 ( .A(n8881), .ZN(n8813) );
  NAND2_X1 U10185 ( .A1(n8824), .A2(n8803), .ZN(n8805) );
  NAND2_X1 U10186 ( .A1(n8805), .A2(n8804), .ZN(n8807) );
  XNOR2_X1 U10187 ( .A(n8807), .B(n8806), .ZN(n8882) );
  AOI22_X1 U10188 ( .A1(n10353), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8822), 
        .B2(n8808), .ZN(n8809) );
  OAI21_X1 U10189 ( .B1(n8976), .B2(n8810), .A(n8809), .ZN(n8811) );
  AOI21_X1 U10190 ( .B1(n8882), .B2(n8825), .A(n8811), .ZN(n8812) );
  OAI21_X1 U10191 ( .B1(n8813), .B2(n10353), .A(n8812), .ZN(P2_U3218) );
  INV_X1 U10192 ( .A(n10343), .ZN(n8820) );
  NAND2_X1 U10193 ( .A1(n8815), .A2(n8814), .ZN(n8816) );
  XNOR2_X1 U10194 ( .A(n8816), .B(n8823), .ZN(n8817) );
  OAI222_X1 U10195 ( .A1(n8901), .A2(n8819), .B1(n8899), .B2(n8818), .C1(n8817), .C2(n8896), .ZN(n8886) );
  AOI21_X1 U10196 ( .B1(n8820), .B2(n8885), .A(n8886), .ZN(n8828) );
  AOI22_X1 U10197 ( .A1(n10353), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8822), 
        .B2(n8821), .ZN(n8827) );
  XNOR2_X1 U10198 ( .A(n8824), .B(n8823), .ZN(n8887) );
  NAND2_X1 U10199 ( .A1(n8887), .A2(n8825), .ZN(n8826) );
  OAI211_X1 U10200 ( .C1(n8828), .C2(n10353), .A(n8827), .B(n8826), .ZN(
        P2_U3219) );
  NOR2_X1 U10201 ( .A1(n8927), .A2(n8924), .ZN(n8830) );
  AOI21_X1 U10202 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n8924), .A(n8830), .ZN(
        n8829) );
  OAI21_X1 U10203 ( .B1(n8929), .B2(n8890), .A(n8829), .ZN(P2_U3490) );
  AOI21_X1 U10204 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n8924), .A(n8830), .ZN(
        n8831) );
  OAI21_X1 U10205 ( .B1(n8932), .B2(n8890), .A(n8831), .ZN(P2_U3489) );
  AOI21_X1 U10206 ( .B1(n5700), .B2(n8833), .A(n8832), .ZN(n8933) );
  OAI21_X1 U10207 ( .B1(n8936), .B2(n8890), .A(n8834), .ZN(P2_U3486) );
  INV_X1 U10208 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8837) );
  AOI21_X1 U10209 ( .B1(n5700), .B2(n8836), .A(n8835), .ZN(n8937) );
  MUX2_X1 U10210 ( .A(n8837), .B(n8937), .S(n8925), .Z(n8838) );
  OAI21_X1 U10211 ( .B1(n8940), .B2(n8890), .A(n8838), .ZN(P2_U3485) );
  AOI21_X1 U10212 ( .B1(n5700), .B2(n8840), .A(n8839), .ZN(n8941) );
  MUX2_X1 U10213 ( .A(n10028), .B(n8941), .S(n8925), .Z(n8841) );
  OAI21_X1 U10214 ( .B1(n8944), .B2(n8890), .A(n8841), .ZN(P2_U3484) );
  INV_X1 U10215 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8844) );
  AOI21_X1 U10216 ( .B1(n8843), .B2(n5700), .A(n8842), .ZN(n8945) );
  MUX2_X1 U10217 ( .A(n8844), .B(n8945), .S(n8925), .Z(n8845) );
  OAI21_X1 U10218 ( .B1(n8948), .B2(n8890), .A(n8845), .ZN(P2_U3483) );
  AOI21_X1 U10219 ( .B1(n5700), .B2(n8847), .A(n8846), .ZN(n8949) );
  MUX2_X1 U10220 ( .A(n8848), .B(n8949), .S(n8925), .Z(n8849) );
  OAI21_X1 U10221 ( .B1(n8952), .B2(n8890), .A(n8849), .ZN(P2_U3482) );
  INV_X1 U10222 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8852) );
  AOI21_X1 U10223 ( .B1(n5700), .B2(n8851), .A(n8850), .ZN(n8953) );
  MUX2_X1 U10224 ( .A(n8852), .B(n8953), .S(n8925), .Z(n8853) );
  OAI21_X1 U10225 ( .B1(n8955), .B2(n8890), .A(n8853), .ZN(P2_U3481) );
  AOI21_X1 U10226 ( .B1(n8855), .B2(n5700), .A(n8854), .ZN(n8956) );
  MUX2_X1 U10227 ( .A(n10033), .B(n8956), .S(n8925), .Z(n8856) );
  OAI21_X1 U10228 ( .B1(n8958), .B2(n8890), .A(n8856), .ZN(P2_U3480) );
  INV_X1 U10229 ( .A(n8857), .ZN(n8858) );
  AOI21_X1 U10230 ( .B1(n5700), .B2(n8859), .A(n8858), .ZN(n8959) );
  MUX2_X1 U10231 ( .A(n8860), .B(n8959), .S(n8925), .Z(n8861) );
  OAI21_X1 U10232 ( .B1(n8962), .B2(n8890), .A(n8861), .ZN(P2_U3479) );
  NAND2_X1 U10233 ( .A1(n8862), .A2(n5700), .ZN(n8865) );
  OAI22_X1 U10234 ( .A1(n8865), .A2(n8864), .B1(n8863), .B2(n8917), .ZN(n8866)
         );
  MUX2_X1 U10235 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8963), .S(n8925), .Z(
        P2_U3478) );
  INV_X1 U10236 ( .A(n8868), .ZN(n8967) );
  INV_X1 U10237 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8871) );
  AOI21_X1 U10238 ( .B1(n8870), .B2(n5700), .A(n8869), .ZN(n8964) );
  MUX2_X1 U10239 ( .A(n8871), .B(n8964), .S(n8925), .Z(n8872) );
  OAI21_X1 U10240 ( .B1(n8967), .B2(n8890), .A(n8872), .ZN(P2_U3477) );
  AOI21_X1 U10241 ( .B1(n8874), .B2(n5700), .A(n8873), .ZN(n8968) );
  MUX2_X1 U10242 ( .A(n8875), .B(n8968), .S(n8925), .Z(n8876) );
  OAI21_X1 U10243 ( .B1(n8971), .B2(n8890), .A(n8876), .ZN(P2_U3476) );
  NAND2_X1 U10244 ( .A1(n8877), .A2(n8908), .ZN(n8878) );
  OAI211_X1 U10245 ( .C1(n8912), .C2(n8880), .A(n8879), .B(n8878), .ZN(n8972)
         );
  MUX2_X1 U10246 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8972), .S(n8925), .Z(
        P2_U3475) );
  AOI21_X1 U10247 ( .B1(n5700), .B2(n8882), .A(n8881), .ZN(n8973) );
  MUX2_X1 U10248 ( .A(n8883), .B(n8973), .S(n8925), .Z(n8884) );
  OAI21_X1 U10249 ( .B1(n8976), .B2(n8890), .A(n8884), .ZN(P2_U3474) );
  INV_X1 U10250 ( .A(n8885), .ZN(n8981) );
  AOI21_X1 U10251 ( .B1(n5700), .B2(n8887), .A(n8886), .ZN(n8977) );
  MUX2_X1 U10252 ( .A(n8888), .B(n8977), .S(n8925), .Z(n8889) );
  OAI21_X1 U10253 ( .B1(n8981), .B2(n8890), .A(n8889), .ZN(P2_U3473) );
  XOR2_X1 U10254 ( .A(n8891), .B(n8894), .Z(n10236) );
  INV_X1 U10255 ( .A(n8892), .ZN(n8893) );
  NOR2_X1 U10256 ( .A1(n8893), .A2(n8917), .ZN(n10228) );
  XNOR2_X1 U10257 ( .A(n8895), .B(n8894), .ZN(n8897) );
  OAI222_X1 U10258 ( .A1(n8901), .A2(n8900), .B1(n8899), .B2(n8898), .C1(n8897), .C2(n8896), .ZN(n10233) );
  AOI211_X1 U10259 ( .C1(n10236), .C2(n5700), .A(n10228), .B(n10233), .ZN(
        n10239) );
  OR2_X1 U10260 ( .A1(n10239), .A2(n8924), .ZN(n8902) );
  OAI21_X1 U10261 ( .B1(n8925), .B2(n8903), .A(n8902), .ZN(P2_U3472) );
  INV_X1 U10262 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8910) );
  NOR2_X1 U10263 ( .A1(n8904), .A2(n8912), .ZN(n8906) );
  AOI211_X1 U10264 ( .C1(n8908), .C2(n8907), .A(n8906), .B(n8905), .ZN(n10373)
         );
  OR2_X1 U10265 ( .A1(n10373), .A2(n8924), .ZN(n8909) );
  OAI21_X1 U10266 ( .B1(n8925), .B2(n8910), .A(n8909), .ZN(P2_U3471) );
  OAI22_X1 U10267 ( .A1(n8913), .A2(n8912), .B1(n8911), .B2(n8917), .ZN(n8914)
         );
  NOR2_X1 U10268 ( .A1(n8915), .A2(n8914), .ZN(n10370) );
  OR2_X1 U10269 ( .A1(n8925), .A2(n5272), .ZN(n8916) );
  OAI21_X1 U10270 ( .B1(n10370), .B2(n8924), .A(n8916), .ZN(P2_U3470) );
  NOR2_X1 U10271 ( .A1(n8918), .A2(n8917), .ZN(n8920) );
  AOI211_X1 U10272 ( .C1(n8922), .C2(n8921), .A(n8920), .B(n8919), .ZN(n10368)
         );
  NAND2_X1 U10273 ( .A1(n8924), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8923) );
  OAI21_X1 U10274 ( .B1(n10368), .B2(n8924), .A(n8923), .ZN(P2_U3469) );
  MUX2_X1 U10275 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n8926), .S(n8925), .Z(
        P2_U3459) );
  NOR2_X1 U10276 ( .A1(n8927), .A2(n10375), .ZN(n8930) );
  AOI21_X1 U10277 ( .B1(n10375), .B2(P2_REG0_REG_31__SCAN_IN), .A(n8930), .ZN(
        n8928) );
  OAI21_X1 U10278 ( .B1(n8929), .B2(n8980), .A(n8928), .ZN(P2_U3458) );
  AOI21_X1 U10279 ( .B1(n10375), .B2(P2_REG0_REG_30__SCAN_IN), .A(n8930), .ZN(
        n8931) );
  OAI21_X1 U10280 ( .B1(n8932), .B2(n8980), .A(n8931), .ZN(P2_U3457) );
  INV_X1 U10281 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8934) );
  OAI21_X1 U10282 ( .B1(n8936), .B2(n8980), .A(n8935), .ZN(P2_U3454) );
  INV_X1 U10283 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8938) );
  MUX2_X1 U10284 ( .A(n8938), .B(n8937), .S(n10372), .Z(n8939) );
  OAI21_X1 U10285 ( .B1(n8940), .B2(n8980), .A(n8939), .ZN(P2_U3453) );
  INV_X1 U10286 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8942) );
  MUX2_X1 U10287 ( .A(n8942), .B(n8941), .S(n10372), .Z(n8943) );
  OAI21_X1 U10288 ( .B1(n8944), .B2(n8980), .A(n8943), .ZN(P2_U3452) );
  INV_X1 U10289 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8946) );
  MUX2_X1 U10290 ( .A(n8946), .B(n8945), .S(n10372), .Z(n8947) );
  OAI21_X1 U10291 ( .B1(n8948), .B2(n8980), .A(n8947), .ZN(P2_U3451) );
  INV_X1 U10292 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8950) );
  MUX2_X1 U10293 ( .A(n8950), .B(n8949), .S(n10372), .Z(n8951) );
  OAI21_X1 U10294 ( .B1(n8952), .B2(n8980), .A(n8951), .ZN(P2_U3450) );
  INV_X1 U10295 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9793) );
  MUX2_X1 U10296 ( .A(n9793), .B(n8953), .S(n10372), .Z(n8954) );
  OAI21_X1 U10297 ( .B1(n8955), .B2(n8980), .A(n8954), .ZN(P2_U3449) );
  MUX2_X1 U10298 ( .A(n9972), .B(n8956), .S(n10372), .Z(n8957) );
  OAI21_X1 U10299 ( .B1(n8958), .B2(n8980), .A(n8957), .ZN(P2_U3448) );
  MUX2_X1 U10300 ( .A(n8960), .B(n8959), .S(n10372), .Z(n8961) );
  OAI21_X1 U10301 ( .B1(n8962), .B2(n8980), .A(n8961), .ZN(P2_U3447) );
  MUX2_X1 U10302 ( .A(n8963), .B(P2_REG0_REG_19__SCAN_IN), .S(n10375), .Z(
        P2_U3446) );
  INV_X1 U10303 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8965) );
  MUX2_X1 U10304 ( .A(n8965), .B(n8964), .S(n10372), .Z(n8966) );
  OAI21_X1 U10305 ( .B1(n8967), .B2(n8980), .A(n8966), .ZN(P2_U3444) );
  INV_X1 U10306 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8969) );
  MUX2_X1 U10307 ( .A(n8969), .B(n8968), .S(n10372), .Z(n8970) );
  OAI21_X1 U10308 ( .B1(n8971), .B2(n8980), .A(n8970), .ZN(P2_U3441) );
  MUX2_X1 U10309 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8972), .S(n10372), .Z(
        P2_U3438) );
  INV_X1 U10310 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8974) );
  MUX2_X1 U10311 ( .A(n8974), .B(n8973), .S(n10372), .Z(n8975) );
  OAI21_X1 U10312 ( .B1(n8976), .B2(n8980), .A(n8975), .ZN(P2_U3435) );
  INV_X1 U10313 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8978) );
  MUX2_X1 U10314 ( .A(n8978), .B(n8977), .S(n10372), .Z(n8979) );
  OAI21_X1 U10315 ( .B1(n8981), .B2(n8980), .A(n8979), .ZN(P2_U3432) );
  INV_X1 U10316 ( .A(n8982), .ZN(n10217) );
  NOR4_X1 U10317 ( .A1(n4960), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n5058), .ZN(n8984) );
  AOI21_X1 U10318 ( .B1(n8991), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8984), .ZN(
        n8985) );
  OAI21_X1 U10319 ( .B1(n10217), .B2(n8993), .A(n8985), .ZN(P2_U3264) );
  INV_X1 U10320 ( .A(n8986), .ZN(n10218) );
  OAI222_X1 U10321 ( .A1(P2_U3151), .A2(n8989), .B1(n8993), .B2(n10218), .C1(
        n8988), .C2(n8987), .ZN(P2_U3266) );
  AOI21_X1 U10322 ( .B1(n8991), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n8990), .ZN(
        n8992) );
  OAI21_X1 U10323 ( .B1(n8994), .B2(n8993), .A(n8992), .ZN(P2_U3267) );
  MUX2_X1 U10324 ( .A(n8995), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  NAND2_X1 U10325 ( .A1(n9000), .A2(n9089), .ZN(n8997) );
  NAND2_X1 U10326 ( .A1(n10154), .A2(n9074), .ZN(n8996) );
  NAND2_X1 U10327 ( .A1(n8997), .A2(n8996), .ZN(n8998) );
  XNOR2_X1 U10328 ( .A(n8998), .B(n9165), .ZN(n9001) );
  AND2_X1 U10329 ( .A1(n10154), .A2(n9115), .ZN(n8999) );
  AOI21_X1 U10330 ( .B1(n9000), .B2(n4409), .A(n8999), .ZN(n9002) );
  NAND2_X1 U10331 ( .A1(n9001), .A2(n9002), .ZN(n9007) );
  INV_X1 U10332 ( .A(n9001), .ZN(n9004) );
  INV_X1 U10333 ( .A(n9002), .ZN(n9003) );
  NAND2_X1 U10334 ( .A1(n9004), .A2(n9003), .ZN(n9005) );
  NAND2_X1 U10335 ( .A1(n9007), .A2(n9005), .ZN(n9197) );
  INV_X1 U10336 ( .A(n9007), .ZN(n9256) );
  NAND2_X1 U10337 ( .A1(n9012), .A2(n9089), .ZN(n9009) );
  NAND2_X1 U10338 ( .A1(n9742), .A2(n4409), .ZN(n9008) );
  NAND2_X1 U10339 ( .A1(n9009), .A2(n9008), .ZN(n9010) );
  XNOR2_X1 U10340 ( .A(n9010), .B(n9165), .ZN(n9013) );
  AND2_X1 U10341 ( .A1(n9742), .A2(n9115), .ZN(n9011) );
  AOI21_X1 U10342 ( .B1(n9012), .B2(n9074), .A(n9011), .ZN(n9014) );
  NAND2_X1 U10343 ( .A1(n9013), .A2(n9014), .ZN(n9018) );
  INV_X1 U10344 ( .A(n9013), .ZN(n9016) );
  INV_X1 U10345 ( .A(n9014), .ZN(n9015) );
  NAND2_X1 U10346 ( .A1(n9016), .A2(n9015), .ZN(n9017) );
  AND2_X1 U10347 ( .A1(n9018), .A2(n9017), .ZN(n9255) );
  AOI22_X1 U10348 ( .A1(n9752), .A2(n9089), .B1(n4409), .B2(n10153), .ZN(n9019) );
  INV_X1 U10349 ( .A(n4440), .ZN(n9020) );
  AOI22_X1 U10350 ( .A1(n9752), .A2(n9074), .B1(n9115), .B2(n10153), .ZN(n9134) );
  INV_X1 U10351 ( .A(n9026), .ZN(n9024) );
  AOI22_X1 U10352 ( .A1(n10247), .A2(n9089), .B1(n9074), .B2(n10144), .ZN(
        n9022) );
  XNOR2_X1 U10353 ( .A(n9022), .B(n4410), .ZN(n9025) );
  INV_X1 U10354 ( .A(n9025), .ZN(n9023) );
  NAND2_X1 U10355 ( .A1(n9024), .A2(n9023), .ZN(n9027) );
  NAND2_X1 U10356 ( .A1(n9026), .A2(n9025), .ZN(n9028) );
  AOI22_X1 U10357 ( .A1(n10247), .A2(n9074), .B1(n9115), .B2(n10144), .ZN(
        n9298) );
  NAND2_X1 U10358 ( .A1(n9299), .A2(n9298), .ZN(n9214) );
  NAND2_X1 U10359 ( .A1(n9695), .A2(n9089), .ZN(n9030) );
  NAND2_X1 U10360 ( .A1(n10143), .A2(n9074), .ZN(n9029) );
  NAND2_X1 U10361 ( .A1(n9030), .A2(n9029), .ZN(n9031) );
  XNOR2_X1 U10362 ( .A(n9031), .B(n4410), .ZN(n9045) );
  AOI22_X1 U10363 ( .A1(n9695), .A2(n9074), .B1(n9115), .B2(n10143), .ZN(n9043) );
  XNOR2_X1 U10364 ( .A(n9045), .B(n9043), .ZN(n9226) );
  INV_X1 U10365 ( .A(n9226), .ZN(n9033) );
  AOI22_X1 U10366 ( .A1(n9713), .A2(n9089), .B1(n9074), .B2(n9690), .ZN(n9032)
         );
  XOR2_X1 U10367 ( .A(n4410), .B(n9032), .Z(n9038) );
  OAI22_X1 U10368 ( .A1(n10205), .A2(n9062), .B1(n10242), .B2(n9168), .ZN(
        n9037) );
  NOR2_X1 U10369 ( .A1(n9038), .A2(n9037), .ZN(n9036) );
  INV_X1 U10370 ( .A(n9036), .ZN(n9222) );
  NAND2_X1 U10371 ( .A1(n9214), .A2(n9034), .ZN(n9042) );
  INV_X1 U10372 ( .A(n9035), .ZN(n9040) );
  AOI21_X1 U10373 ( .B1(n9038), .B2(n9037), .A(n9036), .ZN(n9216) );
  AND2_X1 U10374 ( .A1(n9216), .A2(n9226), .ZN(n9039) );
  NAND2_X1 U10375 ( .A1(n9042), .A2(n9041), .ZN(n9224) );
  INV_X1 U10376 ( .A(n9043), .ZN(n9044) );
  NAND2_X1 U10377 ( .A1(n9682), .A2(n9089), .ZN(n9048) );
  NAND2_X1 U10378 ( .A1(n10119), .A2(n9074), .ZN(n9047) );
  NAND2_X1 U10379 ( .A1(n9048), .A2(n9047), .ZN(n9049) );
  XNOR2_X1 U10380 ( .A(n9049), .B(n4410), .ZN(n9053) );
  NAND2_X1 U10381 ( .A1(n9682), .A2(n9074), .ZN(n9051) );
  NAND2_X1 U10382 ( .A1(n10119), .A2(n9115), .ZN(n9050) );
  NAND2_X1 U10383 ( .A1(n9051), .A2(n9050), .ZN(n9052) );
  NOR2_X1 U10384 ( .A1(n9053), .A2(n9052), .ZN(n9275) );
  NAND2_X1 U10385 ( .A1(n9053), .A2(n9052), .ZN(n9276) );
  NAND2_X1 U10386 ( .A1(n9663), .A2(n9089), .ZN(n9055) );
  NAND2_X1 U10387 ( .A1(n10130), .A2(n9074), .ZN(n9054) );
  NAND2_X1 U10388 ( .A1(n9055), .A2(n9054), .ZN(n9056) );
  XNOR2_X1 U10389 ( .A(n9056), .B(n9165), .ZN(n9156) );
  AND2_X1 U10390 ( .A1(n10130), .A2(n9115), .ZN(n9057) );
  AOI21_X1 U10391 ( .B1(n9663), .B2(n9074), .A(n9057), .ZN(n9058) );
  NAND2_X1 U10392 ( .A1(n9156), .A2(n9058), .ZN(n9060) );
  INV_X1 U10393 ( .A(n9156), .ZN(n9059) );
  INV_X1 U10394 ( .A(n9058), .ZN(n9155) );
  AOI22_X1 U10395 ( .A1(n10116), .A2(n9089), .B1(n9074), .B2(n10120), .ZN(
        n9061) );
  XOR2_X1 U10396 ( .A(n4410), .B(n9061), .Z(n9064) );
  INV_X1 U10397 ( .A(n10116), .ZN(n9649) );
  OAI22_X1 U10398 ( .A1(n9649), .A2(n9062), .B1(n9661), .B2(n9168), .ZN(n9063)
         );
  NOR2_X1 U10399 ( .A1(n9064), .A2(n9063), .ZN(n9065) );
  AOI21_X1 U10400 ( .B1(n9064), .B2(n9063), .A(n9065), .ZN(n9247) );
  INV_X1 U10401 ( .A(n9065), .ZN(n9066) );
  NAND2_X1 U10402 ( .A1(n9246), .A2(n9066), .ZN(n9187) );
  NAND2_X1 U10403 ( .A1(n9629), .A2(n9089), .ZN(n9068) );
  NAND2_X1 U10404 ( .A1(n9641), .A2(n9074), .ZN(n9067) );
  NAND2_X1 U10405 ( .A1(n9068), .A2(n9067), .ZN(n9069) );
  XNOR2_X1 U10406 ( .A(n9069), .B(n4410), .ZN(n9072) );
  AOI22_X1 U10407 ( .A1(n9629), .A2(n9074), .B1(n9115), .B2(n9641), .ZN(n9070)
         );
  XNOR2_X1 U10408 ( .A(n9072), .B(n9070), .ZN(n9188) );
  INV_X1 U10409 ( .A(n9070), .ZN(n9071) );
  AOI22_X1 U10410 ( .A1(n10106), .A2(n9089), .B1(n9074), .B2(n9624), .ZN(n9075) );
  XNOR2_X1 U10411 ( .A(n9075), .B(n4410), .ZN(n9077) );
  INV_X1 U10412 ( .A(n9077), .ZN(n9076) );
  AOI22_X1 U10413 ( .A1(n10106), .A2(n9074), .B1(n9115), .B2(n9624), .ZN(n9267) );
  NAND2_X1 U10414 ( .A1(n10100), .A2(n9089), .ZN(n9081) );
  NAND2_X1 U10415 ( .A1(n9607), .A2(n9074), .ZN(n9080) );
  NAND2_X1 U10416 ( .A1(n9081), .A2(n9080), .ZN(n9082) );
  XNOR2_X1 U10417 ( .A(n9082), .B(n9165), .ZN(n9084) );
  AND2_X1 U10418 ( .A1(n9607), .A2(n9115), .ZN(n9083) );
  AOI21_X1 U10419 ( .B1(n10100), .B2(n9074), .A(n9083), .ZN(n9085) );
  NAND2_X1 U10420 ( .A1(n9084), .A2(n9085), .ZN(n9232) );
  INV_X1 U10421 ( .A(n9084), .ZN(n9087) );
  INV_X1 U10422 ( .A(n9085), .ZN(n9086) );
  NAND2_X1 U10423 ( .A1(n9087), .A2(n9086), .ZN(n9088) );
  NAND2_X1 U10424 ( .A1(n9146), .A2(n9232), .ZN(n9099) );
  NAND2_X1 U10425 ( .A1(n10096), .A2(n4407), .ZN(n9091) );
  NAND2_X1 U10426 ( .A1(n10085), .A2(n9074), .ZN(n9090) );
  NAND2_X1 U10427 ( .A1(n9091), .A2(n9090), .ZN(n9092) );
  XNOR2_X1 U10428 ( .A(n9092), .B(n9165), .ZN(n9094) );
  AND2_X1 U10429 ( .A1(n10085), .A2(n9115), .ZN(n9093) );
  AOI21_X1 U10430 ( .B1(n10096), .B2(n9074), .A(n9093), .ZN(n9095) );
  NAND2_X1 U10431 ( .A1(n9094), .A2(n9095), .ZN(n9100) );
  INV_X1 U10432 ( .A(n9094), .ZN(n9097) );
  INV_X1 U10433 ( .A(n9095), .ZN(n9096) );
  NAND2_X1 U10434 ( .A1(n9097), .A2(n9096), .ZN(n9098) );
  NAND2_X1 U10435 ( .A1(n9099), .A2(n9233), .ZN(n9236) );
  NAND2_X1 U10436 ( .A1(n9574), .A2(n9089), .ZN(n9102) );
  NAND2_X1 U10437 ( .A1(n10076), .A2(n9074), .ZN(n9101) );
  NAND2_X1 U10438 ( .A1(n9102), .A2(n9101), .ZN(n9103) );
  XNOR2_X1 U10439 ( .A(n9103), .B(n4410), .ZN(n9108) );
  AOI22_X1 U10440 ( .A1(n9574), .A2(n9074), .B1(n9115), .B2(n10076), .ZN(n9109) );
  XNOR2_X1 U10441 ( .A(n9108), .B(n9109), .ZN(n9208) );
  NAND2_X1 U10442 ( .A1(n9561), .A2(n9089), .ZN(n9105) );
  NAND2_X1 U10443 ( .A1(n10086), .A2(n9074), .ZN(n9104) );
  NAND2_X1 U10444 ( .A1(n9105), .A2(n9104), .ZN(n9106) );
  XNOR2_X1 U10445 ( .A(n9106), .B(n4410), .ZN(n9122) );
  AND2_X1 U10446 ( .A1(n10086), .A2(n9115), .ZN(n9107) );
  AOI21_X1 U10447 ( .B1(n9561), .B2(n9074), .A(n9107), .ZN(n9120) );
  XNOR2_X1 U10448 ( .A(n9122), .B(n9120), .ZN(n9290) );
  INV_X1 U10449 ( .A(n9108), .ZN(n9110) );
  NAND2_X1 U10450 ( .A1(n9110), .A2(n9109), .ZN(n9287) );
  NAND2_X1 U10451 ( .A1(n9545), .A2(n9089), .ZN(n9113) );
  NAND2_X1 U10452 ( .A1(n10077), .A2(n9074), .ZN(n9112) );
  NAND2_X1 U10453 ( .A1(n9113), .A2(n9112), .ZN(n9114) );
  XNOR2_X1 U10454 ( .A(n9114), .B(n4410), .ZN(n9119) );
  NAND2_X1 U10455 ( .A1(n9545), .A2(n9074), .ZN(n9117) );
  NAND2_X1 U10456 ( .A1(n10077), .A2(n9115), .ZN(n9116) );
  NAND2_X1 U10457 ( .A1(n9117), .A2(n9116), .ZN(n9118) );
  NOR2_X1 U10458 ( .A1(n9119), .A2(n9118), .ZN(n9180) );
  AOI21_X1 U10459 ( .B1(n9119), .B2(n9118), .A(n9180), .ZN(n9125) );
  INV_X1 U10460 ( .A(n9125), .ZN(n9123) );
  INV_X1 U10461 ( .A(n9120), .ZN(n9121) );
  NOR2_X1 U10462 ( .A1(n9123), .A2(n4443), .ZN(n9124) );
  AOI22_X1 U10463 ( .A1(n10086), .A2(n9303), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9127) );
  NAND2_X1 U10464 ( .A1(n9540), .A2(n9307), .ZN(n9126) );
  OAI211_X1 U10465 ( .C1(n10067), .C2(n9305), .A(n9127), .B(n9126), .ZN(n9128)
         );
  AOI21_X1 U10466 ( .B1(n9545), .B2(n9283), .A(n9128), .ZN(n9129) );
  NAND2_X1 U10467 ( .A1(n9130), .A2(n9129), .ZN(P1_U3214) );
  NOR2_X1 U10468 ( .A1(n9132), .A2(n9131), .ZN(n9133) );
  XOR2_X1 U10469 ( .A(n9134), .B(n9133), .Z(n9140) );
  NAND2_X1 U10470 ( .A1(n9307), .A2(n9749), .ZN(n9137) );
  AOI21_X1 U10471 ( .B1(n10144), .B2(n9295), .A(n9135), .ZN(n9136) );
  OAI211_X1 U10472 ( .C1(n9473), .C2(n9293), .A(n9137), .B(n9136), .ZN(n9138)
         );
  AOI21_X1 U10473 ( .B1(n9752), .B2(n9283), .A(n9138), .ZN(n9139) );
  OAI21_X1 U10474 ( .B1(n9140), .B2(n9285), .A(n9139), .ZN(P1_U3215) );
  INV_X1 U10475 ( .A(n9141), .ZN(n9145) );
  INV_X1 U10476 ( .A(n9142), .ZN(n9144) );
  NOR3_X1 U10477 ( .A1(n9145), .A2(n9144), .A3(n9143), .ZN(n9147) );
  INV_X1 U10478 ( .A(n9146), .ZN(n9235) );
  OAI21_X1 U10479 ( .B1(n9147), .B2(n9235), .A(n9300), .ZN(n9153) );
  INV_X1 U10480 ( .A(n9148), .ZN(n9593) );
  AOI22_X1 U10481 ( .A1(n9624), .A2(n9303), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n9149) );
  OAI21_X1 U10482 ( .B1(n9150), .B2(n9305), .A(n9149), .ZN(n9151) );
  AOI21_X1 U10483 ( .B1(n9593), .B2(n9307), .A(n9151), .ZN(n9152) );
  OAI211_X1 U10484 ( .C1(n9595), .C2(n9310), .A(n9153), .B(n9152), .ZN(
        P1_U3216) );
  XNOR2_X1 U10485 ( .A(n9156), .B(n9155), .ZN(n9157) );
  XNOR2_X1 U10486 ( .A(n9154), .B(n9157), .ZN(n9162) );
  NAND2_X1 U10487 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9441) );
  OAI21_X1 U10488 ( .B1(n9661), .B2(n9305), .A(n9441), .ZN(n9158) );
  AOI21_X1 U10489 ( .B1(n9303), .B2(n10119), .A(n9158), .ZN(n9159) );
  OAI21_X1 U10490 ( .B1(n9281), .B2(n9657), .A(n9159), .ZN(n9160) );
  AOI21_X1 U10491 ( .B1(n9663), .B2(n9283), .A(n9160), .ZN(n9161) );
  OAI21_X1 U10492 ( .B1(n9162), .B2(n9285), .A(n9161), .ZN(P1_U3219) );
  NAND2_X1 U10493 ( .A1(n9532), .A2(n9089), .ZN(n9164) );
  NAND2_X1 U10494 ( .A1(n9503), .A2(n9074), .ZN(n9163) );
  NAND2_X1 U10495 ( .A1(n9164), .A2(n9163), .ZN(n9166) );
  XNOR2_X1 U10496 ( .A(n9166), .B(n9165), .ZN(n9170) );
  NAND2_X1 U10497 ( .A1(n9532), .A2(n9074), .ZN(n9167) );
  OAI21_X1 U10498 ( .B1(n10067), .B2(n9168), .A(n9167), .ZN(n9169) );
  XNOR2_X1 U10499 ( .A(n9170), .B(n9169), .ZN(n9181) );
  AND2_X1 U10500 ( .A1(n9181), .A2(n9300), .ZN(n9171) );
  NAND2_X1 U10501 ( .A1(n9172), .A2(n9171), .ZN(n9185) );
  INV_X1 U10502 ( .A(n9180), .ZN(n9174) );
  INV_X1 U10503 ( .A(n9181), .ZN(n9173) );
  NAND4_X1 U10504 ( .A1(n9175), .A2(n9174), .A3(n9173), .A4(n9300), .ZN(n9184)
         );
  INV_X1 U10505 ( .A(n9176), .ZN(n9525) );
  AOI22_X1 U10506 ( .A1(n9525), .A2(n9307), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n9178) );
  NAND2_X1 U10507 ( .A1(n10077), .A2(n9303), .ZN(n9177) );
  OAI211_X1 U10508 ( .C1(n9528), .C2(n9305), .A(n9178), .B(n9177), .ZN(n9179)
         );
  AOI21_X1 U10509 ( .B1(n9532), .B2(n9283), .A(n9179), .ZN(n9183) );
  NAND3_X1 U10510 ( .A1(n9181), .A2(n9300), .A3(n9180), .ZN(n9182) );
  NAND4_X1 U10511 ( .A1(n9185), .A2(n9184), .A3(n9183), .A4(n9182), .ZN(
        P1_U3220) );
  OAI21_X1 U10512 ( .B1(n9188), .B2(n9187), .A(n9186), .ZN(n9189) );
  NAND2_X1 U10513 ( .A1(n9189), .A2(n9300), .ZN(n9196) );
  NOR2_X1 U10514 ( .A1(n9190), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9191) );
  AOI21_X1 U10515 ( .B1(n10120), .B2(n9303), .A(n9191), .ZN(n9192) );
  OAI21_X1 U10516 ( .B1(n9193), .B2(n9305), .A(n9192), .ZN(n9194) );
  AOI21_X1 U10517 ( .B1(n9630), .B2(n9307), .A(n9194), .ZN(n9195) );
  OAI211_X1 U10518 ( .C1(n10191), .C2(n9310), .A(n9196), .B(n9195), .ZN(
        P1_U3223) );
  AND3_X1 U10519 ( .A1(n9006), .A2(n9198), .A3(n9197), .ZN(n9199) );
  OAI21_X1 U10520 ( .B1(n4486), .B2(n9199), .A(n9300), .ZN(n9206) );
  AOI21_X1 U10521 ( .B1(n9742), .B2(n9295), .A(n9200), .ZN(n9201) );
  OAI21_X1 U10522 ( .B1(n9202), .B2(n9293), .A(n9201), .ZN(n9203) );
  AOI21_X1 U10523 ( .B1(n9204), .B2(n9307), .A(n9203), .ZN(n9205) );
  OAI211_X1 U10524 ( .C1(n10293), .C2(n9310), .A(n9206), .B(n9205), .ZN(
        P1_U3224) );
  OAI21_X1 U10525 ( .B1(n9208), .B2(n9207), .A(n9288), .ZN(n9209) );
  NAND2_X1 U10526 ( .A1(n9209), .A2(n9300), .ZN(n9213) );
  AOI22_X1 U10527 ( .A1(n10085), .A2(n9303), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9210) );
  OAI21_X1 U10528 ( .B1(n9281), .B2(n9567), .A(n9210), .ZN(n9211) );
  AOI21_X1 U10529 ( .B1(n9295), .B2(n10086), .A(n9211), .ZN(n9212) );
  OAI211_X1 U10530 ( .C1(n10184), .C2(n9310), .A(n9213), .B(n9212), .ZN(
        P1_U3225) );
  NAND2_X1 U10531 ( .A1(n9028), .A2(n9214), .ZN(n9215) );
  NAND2_X1 U10532 ( .A1(n9215), .A2(n9216), .ZN(n9223) );
  OAI21_X1 U10533 ( .B1(n9216), .B2(n9215), .A(n9223), .ZN(n9217) );
  NAND2_X1 U10534 ( .A1(n9217), .A2(n9300), .ZN(n9221) );
  NAND2_X1 U10535 ( .A1(n10144), .A2(n9303), .ZN(n9218) );
  NAND2_X1 U10536 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9376) );
  OAI211_X1 U10537 ( .C1(n9708), .C2(n9305), .A(n9218), .B(n9376), .ZN(n9219)
         );
  AOI21_X1 U10538 ( .B1(n9705), .B2(n9307), .A(n9219), .ZN(n9220) );
  OAI211_X1 U10539 ( .C1(n10205), .C2(n9310), .A(n9221), .B(n9220), .ZN(
        P1_U3226) );
  NAND2_X1 U10540 ( .A1(n9223), .A2(n9222), .ZN(n9225) );
  OAI21_X1 U10541 ( .B1(n9226), .B2(n9225), .A(n9224), .ZN(n9227) );
  NAND2_X1 U10542 ( .A1(n9227), .A2(n9300), .ZN(n9231) );
  NAND2_X1 U10543 ( .A1(n10119), .A2(n9295), .ZN(n9228) );
  NAND2_X1 U10544 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9388) );
  OAI211_X1 U10545 ( .C1(n10242), .C2(n9293), .A(n9228), .B(n9388), .ZN(n9229)
         );
  AOI21_X1 U10546 ( .B1(n9696), .B2(n9307), .A(n9229), .ZN(n9230) );
  OAI211_X1 U10547 ( .C1(n10201), .C2(n9310), .A(n9231), .B(n9230), .ZN(
        P1_U3228) );
  INV_X1 U10548 ( .A(n10096), .ZN(n9588) );
  INV_X1 U10549 ( .A(n9232), .ZN(n9234) );
  NOR3_X1 U10550 ( .A1(n9235), .A2(n9234), .A3(n9233), .ZN(n9238) );
  INV_X1 U10551 ( .A(n9236), .ZN(n9237) );
  OAI21_X1 U10552 ( .B1(n9238), .B2(n9237), .A(n9300), .ZN(n9244) );
  NAND2_X1 U10553 ( .A1(n9607), .A2(n9303), .ZN(n9240) );
  NAND2_X1 U10554 ( .A1(n9585), .A2(n9307), .ZN(n9239) );
  OAI211_X1 U10555 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n9241), .A(n9240), .B(
        n9239), .ZN(n9242) );
  AOI21_X1 U10556 ( .B1(n10076), .B2(n9295), .A(n9242), .ZN(n9243) );
  OAI211_X1 U10557 ( .C1(n9588), .C2(n9310), .A(n9244), .B(n9243), .ZN(
        P1_U3229) );
  OAI21_X1 U10558 ( .B1(n9247), .B2(n9245), .A(n9246), .ZN(n9248) );
  NAND2_X1 U10559 ( .A1(n9248), .A2(n9300), .ZN(n9253) );
  NOR2_X1 U10560 ( .A1(n9281), .A2(n9645), .ZN(n9251) );
  OAI22_X1 U10561 ( .A1(n9491), .A2(n9305), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9249), .ZN(n9250) );
  AOI211_X1 U10562 ( .C1(n9303), .C2(n10130), .A(n9251), .B(n9250), .ZN(n9252)
         );
  OAI211_X1 U10563 ( .C1(n9649), .C2(n9310), .A(n9253), .B(n9252), .ZN(
        P1_U3233) );
  INV_X1 U10564 ( .A(n9254), .ZN(n9258) );
  NOR3_X1 U10565 ( .A1(n4486), .A2(n9256), .A3(n9255), .ZN(n9257) );
  OAI21_X1 U10566 ( .B1(n9258), .B2(n9257), .A(n9300), .ZN(n9265) );
  AOI21_X1 U10567 ( .B1(n10153), .B2(n9295), .A(n9259), .ZN(n9260) );
  OAI21_X1 U10568 ( .B1(n9261), .B2(n9293), .A(n9260), .ZN(n9262) );
  AOI21_X1 U10569 ( .B1(n9263), .B2(n9307), .A(n9262), .ZN(n9264) );
  OAI211_X1 U10570 ( .C1(n10210), .C2(n9310), .A(n9265), .B(n9264), .ZN(
        P1_U3234) );
  INV_X1 U10571 ( .A(n10106), .ZN(n9615) );
  OAI21_X1 U10572 ( .B1(n9267), .B2(n9266), .A(n9141), .ZN(n9268) );
  NAND2_X1 U10573 ( .A1(n9268), .A2(n9300), .ZN(n9273) );
  INV_X1 U10574 ( .A(n9269), .ZN(n9612) );
  AOI22_X1 U10575 ( .A1(n9641), .A2(n9303), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9270) );
  OAI21_X1 U10576 ( .B1(n9496), .B2(n9305), .A(n9270), .ZN(n9271) );
  AOI21_X1 U10577 ( .B1(n9612), .B2(n9307), .A(n9271), .ZN(n9272) );
  OAI211_X1 U10578 ( .C1(n9615), .C2(n9310), .A(n9273), .B(n9272), .ZN(
        P1_U3235) );
  INV_X1 U10579 ( .A(n9275), .ZN(n9277) );
  NAND2_X1 U10580 ( .A1(n9277), .A2(n9276), .ZN(n9278) );
  XNOR2_X1 U10581 ( .A(n9274), .B(n9278), .ZN(n9286) );
  NAND2_X1 U10582 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9407) );
  OAI21_X1 U10583 ( .B1(n9708), .B2(n9293), .A(n9407), .ZN(n9279) );
  AOI21_X1 U10584 ( .B1(n9295), .B2(n10130), .A(n9279), .ZN(n9280) );
  OAI21_X1 U10585 ( .B1(n9281), .B2(n9674), .A(n9280), .ZN(n9282) );
  AOI21_X1 U10586 ( .B1(n9682), .B2(n9283), .A(n9282), .ZN(n9284) );
  OAI21_X1 U10587 ( .B1(n9286), .B2(n9285), .A(n9284), .ZN(P1_U3238) );
  AND2_X1 U10588 ( .A1(n9288), .A2(n9287), .ZN(n9291) );
  OAI211_X1 U10589 ( .C1(n9291), .C2(n9290), .A(n9300), .B(n9289), .ZN(n9297)
         );
  AOI22_X1 U10590 ( .A1(n9552), .A2(n9307), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9292) );
  OAI21_X1 U10591 ( .B1(n9499), .B2(n9293), .A(n9292), .ZN(n9294) );
  AOI21_X1 U10592 ( .B1(n9295), .B2(n10077), .A(n9294), .ZN(n9296) );
  OAI211_X1 U10593 ( .C1(n10180), .C2(n9310), .A(n9297), .B(n9296), .ZN(
        P1_U3240) );
  INV_X1 U10594 ( .A(n10247), .ZN(n9725) );
  OAI21_X1 U10595 ( .B1(n9299), .B2(n9298), .A(n9214), .ZN(n9301) );
  NAND2_X1 U10596 ( .A1(n9301), .A2(n9300), .ZN(n9309) );
  AOI21_X1 U10597 ( .B1(n10153), .B2(n9303), .A(n9302), .ZN(n9304) );
  OAI21_X1 U10598 ( .B1(n10242), .B2(n9305), .A(n9304), .ZN(n9306) );
  AOI21_X1 U10599 ( .B1(n9727), .B2(n9307), .A(n9306), .ZN(n9308) );
  OAI211_X1 U10600 ( .C1(n9725), .C2(n9310), .A(n9309), .B(n9308), .ZN(
        P1_U3241) );
  MUX2_X1 U10601 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9509), .S(P1_U3973), .Z(
        P1_U3584) );
  INV_X1 U10602 ( .A(n9528), .ZN(n10058) );
  MUX2_X1 U10603 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n10058), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10604 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9503), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10605 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n10077), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10606 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n10086), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10607 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n10076), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10608 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n10085), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10609 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9607), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10610 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9624), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10611 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9641), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10612 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n10120), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10613 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n10130), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10614 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n10119), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10615 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n10143), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10616 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9690), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10617 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n10144), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10618 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n10153), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10619 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9742), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10620 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n10154), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10621 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9311), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10622 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9312), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10623 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9313), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10624 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9314), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10625 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9315), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10626 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9316), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10627 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9317), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10628 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9318), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10629 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9319), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10630 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n6893), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10631 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9320), .S(P1_U3973), .Z(
        P1_U3555) );
  MUX2_X1 U10632 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9321), .S(P1_U3973), .Z(
        P1_U3554) );
  INV_X1 U10633 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9322) );
  OAI22_X1 U10634 ( .A1(n9443), .A2(n9853), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9322), .ZN(n9323) );
  AOI21_X1 U10635 ( .B1(n9324), .B2(n9379), .A(n9323), .ZN(n9334) );
  MUX2_X1 U10636 ( .A(n6666), .B(P1_REG1_REG_1__SCAN_IN), .S(n9324), .Z(n9325)
         );
  INV_X1 U10637 ( .A(n9325), .ZN(n9327) );
  OAI211_X1 U10638 ( .C1(n9328), .C2(n9327), .A(n9436), .B(n9326), .ZN(n9333)
         );
  OAI211_X1 U10639 ( .C1(n9331), .C2(n9330), .A(n9437), .B(n9329), .ZN(n9332)
         );
  NAND3_X1 U10640 ( .A1(n9334), .A2(n9333), .A3(n9332), .ZN(P1_U3244) );
  INV_X1 U10641 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9335) );
  OAI22_X1 U10642 ( .A1(n9443), .A2(n9335), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6098), .ZN(n9336) );
  AOI21_X1 U10643 ( .B1(n9337), .B2(n9379), .A(n9336), .ZN(n9345) );
  OAI211_X1 U10644 ( .C1(n9339), .C2(n9338), .A(n9436), .B(n9353), .ZN(n9344)
         );
  OAI211_X1 U10645 ( .C1(n9342), .C2(n9341), .A(n9437), .B(n9340), .ZN(n9343)
         );
  NAND4_X1 U10646 ( .A1(n9346), .A2(n9345), .A3(n9344), .A4(n9343), .ZN(
        P1_U3245) );
  OAI211_X1 U10647 ( .C1(n9349), .C2(n9348), .A(n9437), .B(n9347), .ZN(n9360)
         );
  AOI21_X1 U10648 ( .B1(n9420), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n9350), .ZN(
        n9359) );
  NAND2_X1 U10649 ( .A1(n9379), .A2(n9351), .ZN(n9358) );
  MUX2_X1 U10650 ( .A(n6669), .B(P1_REG1_REG_3__SCAN_IN), .S(n9351), .Z(n9354)
         );
  NAND3_X1 U10651 ( .A1(n9354), .A2(n9353), .A3(n9352), .ZN(n9355) );
  NAND3_X1 U10652 ( .A1(n9436), .A2(n9356), .A3(n9355), .ZN(n9357) );
  NAND4_X1 U10653 ( .A1(n9360), .A2(n9359), .A3(n9358), .A4(n9357), .ZN(
        P1_U3246) );
  NAND2_X1 U10654 ( .A1(n9362), .A2(n9361), .ZN(n9364) );
  NAND2_X1 U10655 ( .A1(n9364), .A2(n9363), .ZN(n9367) );
  NOR2_X1 U10656 ( .A1(n9391), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9384) );
  AOI21_X1 U10657 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(n9391), .A(n9384), .ZN(
        n9365) );
  INV_X1 U10658 ( .A(n9365), .ZN(n9366) );
  NOR2_X1 U10659 ( .A1(n9366), .A2(n9367), .ZN(n9383) );
  AOI21_X1 U10660 ( .B1(n9367), .B2(n9366), .A(n9383), .ZN(n9382) );
  NOR2_X1 U10661 ( .A1(n9369), .A2(n9368), .ZN(n9371) );
  NOR2_X1 U10662 ( .A1(n9371), .A2(n9370), .ZN(n9374) );
  NAND2_X1 U10663 ( .A1(n9391), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9372) );
  OAI21_X1 U10664 ( .B1(n9391), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9372), .ZN(
        n9373) );
  NOR2_X1 U10665 ( .A1(n9374), .A2(n9373), .ZN(n9390) );
  AOI211_X1 U10666 ( .C1(n9374), .C2(n9373), .A(n9390), .B(n9415), .ZN(n9375)
         );
  INV_X1 U10667 ( .A(n9375), .ZN(n9381) );
  INV_X1 U10668 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9377) );
  OAI21_X1 U10669 ( .B1(n9443), .B2(n9377), .A(n9376), .ZN(n9378) );
  AOI21_X1 U10670 ( .B1(n9391), .B2(n9379), .A(n9378), .ZN(n9380) );
  OAI211_X1 U10671 ( .C1(n9382), .C2(n9432), .A(n9381), .B(n9380), .ZN(
        P1_U3259) );
  NOR2_X1 U10672 ( .A1(n9384), .A2(n9383), .ZN(n9386) );
  XNOR2_X1 U10673 ( .A(n9401), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9385) );
  NOR2_X1 U10674 ( .A1(n9386), .A2(n9385), .ZN(n9404) );
  AOI21_X1 U10675 ( .B1(n9386), .B2(n9385), .A(n9404), .ZN(n9387) );
  NOR2_X1 U10676 ( .A1(n9387), .A2(n9432), .ZN(n9399) );
  INV_X1 U10677 ( .A(n9388), .ZN(n9398) );
  INV_X1 U10678 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9389) );
  NOR2_X1 U10679 ( .A1(n9443), .A2(n9389), .ZN(n9397) );
  OR2_X1 U10680 ( .A1(n9401), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9393) );
  NAND2_X1 U10681 ( .A1(n9401), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9392) );
  AND2_X1 U10682 ( .A1(n9393), .A2(n9392), .ZN(n9394) );
  NAND2_X1 U10683 ( .A1(n9410), .A2(n9394), .ZN(n9395) );
  AOI221_X1 U10684 ( .B1(n9410), .B2(n9395), .C1(n9394), .C2(n9395), .A(n9415), 
        .ZN(n9396) );
  NOR4_X1 U10685 ( .A1(n9399), .A2(n9398), .A3(n9397), .A4(n9396), .ZN(n9400)
         );
  OAI21_X1 U10686 ( .B1(n9408), .B2(n9431), .A(n9400), .ZN(P1_U3260) );
  NOR2_X1 U10687 ( .A1(n9401), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9403) );
  XNOR2_X1 U10688 ( .A(n9429), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9402) );
  NOR3_X1 U10689 ( .A1(n9404), .A2(n9403), .A3(n9402), .ZN(n9428) );
  INV_X1 U10690 ( .A(n9428), .ZN(n9406) );
  OAI21_X1 U10691 ( .B1(n9404), .B2(n9403), .A(n9402), .ZN(n9405) );
  NAND3_X1 U10692 ( .A1(n9406), .A2(n9436), .A3(n9405), .ZN(n9422) );
  INV_X1 U10693 ( .A(n9407), .ZN(n9419) );
  INV_X1 U10694 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9409) );
  NAND2_X1 U10695 ( .A1(n9410), .A2(n9409), .ZN(n9411) );
  NAND2_X1 U10696 ( .A1(n9412), .A2(n9411), .ZN(n9417) );
  INV_X1 U10697 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9675) );
  OR2_X1 U10698 ( .A1(n9429), .A2(n9675), .ZN(n9414) );
  NAND2_X1 U10699 ( .A1(n9429), .A2(n9675), .ZN(n9413) );
  AND2_X1 U10700 ( .A1(n9414), .A2(n9413), .ZN(n9416) );
  NOR2_X1 U10701 ( .A1(n9417), .A2(n9416), .ZN(n9425) );
  AOI211_X1 U10702 ( .C1(n9417), .C2(n9416), .A(n9425), .B(n9415), .ZN(n9418)
         );
  AOI211_X1 U10703 ( .C1(n9420), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n9419), .B(
        n9418), .ZN(n9421) );
  OAI211_X1 U10704 ( .C1(n9431), .C2(n9423), .A(n9422), .B(n9421), .ZN(
        P1_U3261) );
  AND2_X1 U10705 ( .A1(n9429), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9424) );
  OR2_X1 U10706 ( .A1(n9425), .A2(n9424), .ZN(n9427) );
  INV_X1 U10707 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9426) );
  XNOR2_X1 U10708 ( .A(n9427), .B(n9426), .ZN(n9438) );
  INV_X1 U10709 ( .A(n9438), .ZN(n9434) );
  AOI21_X1 U10710 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n9429), .A(n9428), .ZN(
        n9430) );
  XNOR2_X1 U10711 ( .A(n9430), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9435) );
  OAI21_X1 U10712 ( .B1(n9435), .B2(n9432), .A(n9431), .ZN(n9433) );
  AOI21_X1 U10713 ( .B1(n9434), .B2(n9437), .A(n9433), .ZN(n9440) );
  AOI22_X1 U10714 ( .A1(n9438), .A2(n9437), .B1(n9436), .B2(n9435), .ZN(n9439)
         );
  MUX2_X1 U10715 ( .A(n9440), .B(n9439), .S(n4408), .Z(n9442) );
  OAI211_X1 U10716 ( .C1(n9444), .C2(n9443), .A(n9442), .B(n9441), .ZN(
        P1_U3262) );
  NOR2_X1 U10717 ( .A1(n9709), .A2(n9713), .ZN(n9693) );
  OR2_X1 U10718 ( .A1(n10106), .A2(n9627), .ZN(n9610) );
  NAND2_X1 U10719 ( .A1(n9588), .A2(n9592), .ZN(n9570) );
  NAND2_X1 U10720 ( .A1(n10168), .A2(n9507), .ZN(n9453) );
  INV_X1 U10721 ( .A(P1_B_REG_SCAN_IN), .ZN(n9447) );
  NOR2_X1 U10722 ( .A1(n10223), .A2(n9447), .ZN(n9448) );
  NOR2_X1 U10723 ( .A1(n10241), .A2(n9448), .ZN(n9508) );
  NAND2_X1 U10724 ( .A1(n9449), .A2(n9508), .ZN(n10047) );
  NOR2_X1 U10725 ( .A1(n10047), .A2(n7001), .ZN(n9455) );
  NOR2_X1 U10726 ( .A1(n9445), .A2(n9724), .ZN(n9451) );
  AOI211_X1 U10727 ( .C1(n7001), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9455), .B(
        n9451), .ZN(n9452) );
  OAI21_X1 U10728 ( .B1(n9761), .B2(n9755), .A(n9452), .ZN(P1_U3263) );
  OAI211_X1 U10729 ( .C1(n10168), .C2(n9507), .A(n9746), .B(n9453), .ZN(n10048) );
  NOR2_X1 U10730 ( .A1(n10168), .A2(n9724), .ZN(n9454) );
  AOI211_X1 U10731 ( .C1(n7001), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9455), .B(
        n9454), .ZN(n9456) );
  OAI21_X1 U10732 ( .B1(n9755), .B2(n10048), .A(n9456), .ZN(P1_U3264) );
  AND2_X2 U10733 ( .A1(n9596), .A2(n9464), .ZN(n9580) );
  INV_X1 U10734 ( .A(n9468), .ZN(n9469) );
  INV_X1 U10735 ( .A(n9521), .ZN(n9471) );
  INV_X1 U10736 ( .A(n10057), .ZN(n9519) );
  INV_X1 U10737 ( .A(n9752), .ZN(n9476) );
  NAND2_X1 U10738 ( .A1(n10201), .A2(n9708), .ZN(n9482) );
  AOI22_X1 U10739 ( .A1(n9685), .A2(n9482), .B1(n9695), .B2(n10143), .ZN(n9672) );
  NAND2_X1 U10740 ( .A1(n9672), .A2(n5015), .ZN(n9485) );
  NAND2_X1 U10741 ( .A1(n9485), .A2(n9484), .ZN(n9652) );
  NAND2_X1 U10742 ( .A1(n9663), .A2(n10130), .ZN(n9487) );
  NOR2_X1 U10743 ( .A1(n9663), .A2(n10130), .ZN(n9486) );
  AOI21_X1 U10744 ( .B1(n9652), .B2(n9487), .A(n9486), .ZN(n9636) );
  NAND2_X1 U10745 ( .A1(n9636), .A2(n9488), .ZN(n9490) );
  OR2_X1 U10746 ( .A1(n10106), .A2(n9624), .ZN(n9492) );
  NAND2_X1 U10747 ( .A1(n10191), .A2(n9491), .ZN(n9604) );
  AND2_X1 U10748 ( .A1(n9492), .A2(n9604), .ZN(n9493) );
  NAND2_X1 U10749 ( .A1(n10106), .A2(n9624), .ZN(n9494) );
  NOR2_X1 U10750 ( .A1(n9595), .A2(n9496), .ZN(n9498) );
  NAND2_X1 U10751 ( .A1(n9595), .A2(n9496), .ZN(n9497) );
  NOR2_X1 U10752 ( .A1(n10184), .A2(n9499), .ZN(n9501) );
  NAND2_X1 U10753 ( .A1(n10184), .A2(n9499), .ZN(n9500) );
  NOR2_X1 U10754 ( .A1(n9561), .A2(n10086), .ZN(n9502) );
  NAND2_X1 U10755 ( .A1(n9532), .A2(n9503), .ZN(n9504) );
  NAND2_X1 U10756 ( .A1(n9524), .A2(n9504), .ZN(n9506) );
  XNOR2_X1 U10757 ( .A(n9506), .B(n9505), .ZN(n10051) );
  NAND2_X1 U10758 ( .A1(n10051), .A2(n9721), .ZN(n9518) );
  AOI211_X1 U10759 ( .C1(n10052), .C2(n4446), .A(n9723), .B(n9507), .ZN(n10056) );
  NAND2_X1 U10760 ( .A1(n10052), .A2(n9751), .ZN(n9514) );
  NAND2_X1 U10761 ( .A1(n9509), .A2(n9508), .ZN(n10053) );
  NOR2_X1 U10762 ( .A1(n10053), .A2(n7001), .ZN(n9512) );
  NOR2_X1 U10763 ( .A1(n9510), .A2(n9673), .ZN(n9511) );
  AOI211_X1 U10764 ( .C1(n7001), .C2(P1_REG2_REG_29__SCAN_IN), .A(n9512), .B(
        n9511), .ZN(n9513) );
  OAI211_X1 U10765 ( .C1(n10067), .C2(n9515), .A(n9514), .B(n9513), .ZN(n9516)
         );
  AOI21_X1 U10766 ( .B1(n10056), .B2(n9733), .A(n9516), .ZN(n9517) );
  OAI211_X1 U10767 ( .C1(n9519), .C2(n9736), .A(n9518), .B(n9517), .ZN(
        P1_U3356) );
  XNOR2_X1 U10768 ( .A(n9520), .B(n9521), .ZN(n10061) );
  NAND2_X1 U10769 ( .A1(n9522), .A2(n9521), .ZN(n9523) );
  NAND2_X1 U10770 ( .A1(n10063), .A2(n9721), .ZN(n9534) );
  AOI22_X1 U10771 ( .A1(n9525), .A2(n9748), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9750), .ZN(n9527) );
  NAND2_X1 U10772 ( .A1(n10077), .A2(n9726), .ZN(n9526) );
  OAI211_X1 U10773 ( .C1(n9528), .C2(n9730), .A(n9527), .B(n9526), .ZN(n9531)
         );
  AOI21_X1 U10774 ( .B1(n4447), .B2(n9532), .A(n9723), .ZN(n9529) );
  NAND2_X1 U10775 ( .A1(n9529), .A2(n4446), .ZN(n10059) );
  NOR2_X1 U10776 ( .A1(n10059), .A2(n9755), .ZN(n9530) );
  AOI211_X1 U10777 ( .C1(n9751), .C2(n9532), .A(n9531), .B(n9530), .ZN(n9533)
         );
  OAI211_X1 U10778 ( .C1(n9736), .C2(n10061), .A(n9534), .B(n9533), .ZN(
        P1_U3265) );
  AOI21_X1 U10779 ( .B1(n9537), .B2(n9536), .A(n9535), .ZN(n10071) );
  XNOR2_X1 U10780 ( .A(n9539), .B(n9538), .ZN(n10073) );
  NAND2_X1 U10781 ( .A1(n10073), .A2(n9721), .ZN(n9547) );
  AOI22_X1 U10782 ( .A1(n10086), .A2(n9726), .B1(n7001), .B2(
        P1_REG2_REG_27__SCAN_IN), .ZN(n9542) );
  NAND2_X1 U10783 ( .A1(n9540), .A2(n9748), .ZN(n9541) );
  OAI211_X1 U10784 ( .C1(n10067), .C2(n9730), .A(n9542), .B(n9541), .ZN(n9544)
         );
  OAI211_X1 U10785 ( .C1(n10176), .C2(n9556), .A(n9746), .B(n4447), .ZN(n10069) );
  NOR2_X1 U10786 ( .A1(n10069), .A2(n9755), .ZN(n9543) );
  AOI211_X1 U10787 ( .C1(n9751), .C2(n9545), .A(n9544), .B(n9543), .ZN(n9546)
         );
  OAI211_X1 U10788 ( .C1(n10071), .C2(n9736), .A(n9547), .B(n9546), .ZN(
        P1_U3266) );
  INV_X1 U10789 ( .A(n9551), .ZN(n9548) );
  XNOR2_X1 U10790 ( .A(n9549), .B(n9548), .ZN(n10080) );
  XOR2_X1 U10791 ( .A(n9551), .B(n9550), .Z(n10082) );
  NAND2_X1 U10792 ( .A1(n10082), .A2(n9721), .ZN(n9563) );
  AOI22_X1 U10793 ( .A1(n9552), .A2(n9748), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9750), .ZN(n9554) );
  NAND2_X1 U10794 ( .A1(n10076), .A2(n9726), .ZN(n9553) );
  OAI211_X1 U10795 ( .C1(n9555), .C2(n9730), .A(n9554), .B(n9553), .ZN(n9560)
         );
  INV_X1 U10796 ( .A(n9571), .ZN(n9558) );
  INV_X1 U10797 ( .A(n9556), .ZN(n9557) );
  OAI211_X1 U10798 ( .C1(n10180), .C2(n9558), .A(n9557), .B(n9746), .ZN(n10078) );
  NOR2_X1 U10799 ( .A1(n10078), .A2(n9755), .ZN(n9559) );
  AOI211_X1 U10800 ( .C1(n9751), .C2(n9561), .A(n9560), .B(n9559), .ZN(n9562)
         );
  OAI211_X1 U10801 ( .C1(n10080), .C2(n9736), .A(n9563), .B(n9562), .ZN(
        P1_U3267) );
  AOI21_X1 U10802 ( .B1(n9566), .B2(n9564), .A(n4459), .ZN(n10089) );
  XOR2_X1 U10803 ( .A(n9566), .B(n9565), .Z(n10091) );
  NAND2_X1 U10804 ( .A1(n10091), .A2(n9721), .ZN(n9576) );
  OAI22_X1 U10805 ( .A1(n9567), .A2(n9673), .B1(n9986), .B2(n9757), .ZN(n9568)
         );
  AOI21_X1 U10806 ( .B1(n9726), .B2(n10085), .A(n9568), .ZN(n9569) );
  OAI21_X1 U10807 ( .B1(n10066), .B2(n9730), .A(n9569), .ZN(n9573) );
  INV_X1 U10808 ( .A(n9570), .ZN(n9583) );
  OAI211_X1 U10809 ( .C1(n9583), .C2(n10184), .A(n9746), .B(n9571), .ZN(n10087) );
  NOR2_X1 U10810 ( .A1(n10087), .A2(n9755), .ZN(n9572) );
  AOI211_X1 U10811 ( .C1(n9751), .C2(n9574), .A(n9573), .B(n9572), .ZN(n9575)
         );
  OAI211_X1 U10812 ( .C1(n10089), .C2(n9736), .A(n9576), .B(n9575), .ZN(
        P1_U3268) );
  XNOR2_X1 U10813 ( .A(n9577), .B(n9579), .ZN(n10098) );
  OAI211_X1 U10814 ( .C1(n9580), .C2(n9579), .A(n9578), .B(n10125), .ZN(n9582)
         );
  AOI22_X1 U10815 ( .A1(n10076), .A2(n10152), .B1(n10155), .B2(n9607), .ZN(
        n9581) );
  NAND2_X1 U10816 ( .A1(n9582), .A2(n9581), .ZN(n10094) );
  INV_X1 U10817 ( .A(n9592), .ZN(n9584) );
  AOI211_X1 U10818 ( .C1(n10096), .C2(n9584), .A(n9723), .B(n9583), .ZN(n10095) );
  NAND2_X1 U10819 ( .A1(n10095), .A2(n9733), .ZN(n9587) );
  AOI22_X1 U10820 ( .A1(n9585), .A2(n9748), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9750), .ZN(n9586) );
  OAI211_X1 U10821 ( .C1(n9588), .C2(n9724), .A(n9587), .B(n9586), .ZN(n9589)
         );
  AOI21_X1 U10822 ( .B1(n10094), .B2(n9757), .A(n9589), .ZN(n9590) );
  OAI21_X1 U10823 ( .B1(n10098), .B2(n9759), .A(n9590), .ZN(P1_U3269) );
  XOR2_X1 U10824 ( .A(n9591), .B(n9597), .Z(n10103) );
  AOI211_X1 U10825 ( .C1(n10100), .C2(n9610), .A(n9723), .B(n9592), .ZN(n10099) );
  AOI22_X1 U10826 ( .A1(n9593), .A2(n9748), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n7001), .ZN(n9594) );
  OAI21_X1 U10827 ( .B1(n9595), .B2(n9724), .A(n9594), .ZN(n9600) );
  OAI21_X1 U10828 ( .B1(n9597), .B2(n4481), .A(n9596), .ZN(n9598) );
  AOI222_X1 U10829 ( .A1(n10125), .A2(n9598), .B1(n10085), .B2(n10152), .C1(
        n9624), .C2(n10155), .ZN(n10102) );
  NOR2_X1 U10830 ( .A1(n10102), .A2(n7001), .ZN(n9599) );
  AOI211_X1 U10831 ( .C1(n10099), .C2(n9733), .A(n9600), .B(n9599), .ZN(n9601)
         );
  OAI21_X1 U10832 ( .B1(n10103), .B2(n9759), .A(n9601), .ZN(P1_U3270) );
  NAND2_X1 U10833 ( .A1(n9602), .A2(n9604), .ZN(n9605) );
  XNOR2_X1 U10834 ( .A(n9605), .B(n9462), .ZN(n10108) );
  OAI211_X1 U10835 ( .C1(n4480), .C2(n9462), .A(n9606), .B(n10125), .ZN(n9609)
         );
  AOI22_X1 U10836 ( .A1(n9607), .A2(n10152), .B1(n10155), .B2(n9641), .ZN(
        n9608) );
  NAND2_X1 U10837 ( .A1(n9609), .A2(n9608), .ZN(n10104) );
  INV_X1 U10838 ( .A(n9610), .ZN(n9611) );
  AOI211_X1 U10839 ( .C1(n10106), .C2(n9627), .A(n9723), .B(n9611), .ZN(n10105) );
  NAND2_X1 U10840 ( .A1(n10105), .A2(n9733), .ZN(n9614) );
  AOI22_X1 U10841 ( .A1(n9612), .A2(n9748), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n7001), .ZN(n9613) );
  OAI211_X1 U10842 ( .C1(n9615), .C2(n9724), .A(n9614), .B(n9613), .ZN(n9616)
         );
  AOI21_X1 U10843 ( .B1(n10104), .B2(n9757), .A(n9616), .ZN(n9617) );
  OAI21_X1 U10844 ( .B1(n10108), .B2(n9759), .A(n9617), .ZN(P1_U3271) );
  XNOR2_X1 U10845 ( .A(n9618), .B(n9620), .ZN(n10111) );
  INV_X1 U10846 ( .A(n10111), .ZN(n9635) );
  INV_X1 U10847 ( .A(n9639), .ZN(n9637) );
  OR2_X1 U10848 ( .A1(n9458), .A2(n9637), .ZN(n9638) );
  NAND2_X1 U10849 ( .A1(n9638), .A2(n9619), .ZN(n9622) );
  INV_X1 U10850 ( .A(n9620), .ZN(n9621) );
  XNOR2_X1 U10851 ( .A(n9622), .B(n9621), .ZN(n9623) );
  NAND2_X1 U10852 ( .A1(n9623), .A2(n10125), .ZN(n9626) );
  AOI22_X1 U10853 ( .A1(n9624), .A2(n10152), .B1(n10155), .B2(n10120), .ZN(
        n9625) );
  NAND2_X1 U10854 ( .A1(n9626), .A2(n9625), .ZN(n10109) );
  INV_X1 U10855 ( .A(n9627), .ZN(n9628) );
  AOI211_X1 U10856 ( .C1(n9629), .C2(n4831), .A(n9723), .B(n9628), .ZN(n10110)
         );
  NAND2_X1 U10857 ( .A1(n10110), .A2(n9733), .ZN(n9632) );
  AOI22_X1 U10858 ( .A1(n9630), .A2(n9748), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9750), .ZN(n9631) );
  OAI211_X1 U10859 ( .C1(n10191), .C2(n9724), .A(n9632), .B(n9631), .ZN(n9633)
         );
  AOI21_X1 U10860 ( .B1(n10109), .B2(n9757), .A(n9633), .ZN(n9634) );
  OAI21_X1 U10861 ( .B1(n9635), .B2(n9759), .A(n9634), .ZN(P1_U3272) );
  XNOR2_X1 U10862 ( .A(n9636), .B(n9637), .ZN(n10118) );
  INV_X1 U10863 ( .A(n9458), .ZN(n9640) );
  OAI211_X1 U10864 ( .C1(n9640), .C2(n9639), .A(n10125), .B(n9638), .ZN(n9643)
         );
  AOI22_X1 U10865 ( .A1(n9641), .A2(n10152), .B1(n10155), .B2(n10130), .ZN(
        n9642) );
  NAND2_X1 U10866 ( .A1(n9643), .A2(n9642), .ZN(n10114) );
  AOI211_X1 U10867 ( .C1(n10116), .C2(n9655), .A(n9723), .B(n9644), .ZN(n10115) );
  NAND2_X1 U10868 ( .A1(n10115), .A2(n9733), .ZN(n9648) );
  INV_X1 U10869 ( .A(n9645), .ZN(n9646) );
  AOI22_X1 U10870 ( .A1(n9646), .A2(n9748), .B1(P1_REG2_REG_20__SCAN_IN), .B2(
        n7001), .ZN(n9647) );
  OAI211_X1 U10871 ( .C1(n9649), .C2(n9724), .A(n9648), .B(n9647), .ZN(n9650)
         );
  AOI21_X1 U10872 ( .B1(n10114), .B2(n9757), .A(n9650), .ZN(n9651) );
  OAI21_X1 U10873 ( .B1(n10118), .B2(n9759), .A(n9651), .ZN(P1_U3273) );
  XNOR2_X1 U10874 ( .A(n9652), .B(n9653), .ZN(n10129) );
  XNOR2_X1 U10875 ( .A(n9654), .B(n9653), .ZN(n10126) );
  INV_X1 U10876 ( .A(n9736), .ZN(n9666) );
  INV_X1 U10877 ( .A(n9679), .ZN(n9656) );
  OAI211_X1 U10878 ( .C1(n9656), .C2(n10123), .A(n9746), .B(n9655), .ZN(n10122) );
  INV_X1 U10879 ( .A(n9657), .ZN(n9658) );
  AOI22_X1 U10880 ( .A1(n9658), .A2(n9748), .B1(P1_REG2_REG_19__SCAN_IN), .B2(
        n9750), .ZN(n9660) );
  NAND2_X1 U10881 ( .A1(n10119), .A2(n9726), .ZN(n9659) );
  OAI211_X1 U10882 ( .C1(n9661), .C2(n9730), .A(n9660), .B(n9659), .ZN(n9662)
         );
  AOI21_X1 U10883 ( .B1(n9663), .B2(n9751), .A(n9662), .ZN(n9664) );
  OAI21_X1 U10884 ( .B1(n10122), .B2(n9755), .A(n9664), .ZN(n9665) );
  AOI21_X1 U10885 ( .B1(n10126), .B2(n9666), .A(n9665), .ZN(n9667) );
  OAI21_X1 U10886 ( .B1(n10129), .B2(n9759), .A(n9667), .ZN(P1_U3274) );
  OAI21_X1 U10887 ( .B1(n9669), .B2(n9671), .A(n9668), .ZN(n9670) );
  INV_X1 U10888 ( .A(n9670), .ZN(n10133) );
  XOR2_X1 U10889 ( .A(n9672), .B(n9671), .Z(n10135) );
  NAND2_X1 U10890 ( .A1(n10135), .A2(n9721), .ZN(n9684) );
  OAI22_X1 U10891 ( .A1(n9757), .A2(n9675), .B1(n9674), .B2(n9673), .ZN(n9676)
         );
  AOI21_X1 U10892 ( .B1(n9726), .B2(n10143), .A(n9676), .ZN(n9677) );
  OAI21_X1 U10893 ( .B1(n9678), .B2(n9730), .A(n9677), .ZN(n9681) );
  OAI211_X1 U10894 ( .C1(n9694), .C2(n10197), .A(n9746), .B(n9679), .ZN(n10131) );
  NOR2_X1 U10895 ( .A1(n10131), .A2(n9755), .ZN(n9680) );
  AOI211_X1 U10896 ( .C1(n9751), .C2(n9682), .A(n9681), .B(n9680), .ZN(n9683)
         );
  OAI211_X1 U10897 ( .C1(n10133), .C2(n9736), .A(n9684), .B(n9683), .ZN(
        P1_U3275) );
  XNOR2_X1 U10898 ( .A(n9685), .B(n6304), .ZN(n10140) );
  INV_X1 U10899 ( .A(n10140), .ZN(n9701) );
  NAND2_X1 U10900 ( .A1(n9687), .A2(n9686), .ZN(n9688) );
  NAND3_X1 U10901 ( .A1(n9689), .A2(n10125), .A3(n9688), .ZN(n9692) );
  AOI22_X1 U10902 ( .A1(n10119), .A2(n10152), .B1(n10155), .B2(n9690), .ZN(
        n9691) );
  NAND2_X1 U10903 ( .A1(n9692), .A2(n9691), .ZN(n10138) );
  INV_X1 U10904 ( .A(n9693), .ZN(n9710) );
  AOI211_X1 U10905 ( .C1(n9695), .C2(n9710), .A(n9723), .B(n9694), .ZN(n10139)
         );
  NAND2_X1 U10906 ( .A1(n10139), .A2(n9733), .ZN(n9698) );
  AOI22_X1 U10907 ( .A1(n7001), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9696), .B2(
        n9748), .ZN(n9697) );
  OAI211_X1 U10908 ( .C1(n10201), .C2(n9724), .A(n9698), .B(n9697), .ZN(n9699)
         );
  AOI21_X1 U10909 ( .B1(n10138), .B2(n9757), .A(n9699), .ZN(n9700) );
  OAI21_X1 U10910 ( .B1(n9701), .B2(n9759), .A(n9700), .ZN(P1_U3276) );
  XNOR2_X1 U10911 ( .A(n9702), .B(n9703), .ZN(n10147) );
  XNOR2_X1 U10912 ( .A(n9704), .B(n9703), .ZN(n10149) );
  NAND2_X1 U10913 ( .A1(n10149), .A2(n9721), .ZN(n9715) );
  NAND2_X1 U10914 ( .A1(n9726), .A2(n10144), .ZN(n9707) );
  AOI22_X1 U10915 ( .A1(n9750), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9705), .B2(
        n9748), .ZN(n9706) );
  OAI211_X1 U10916 ( .C1(n9708), .C2(n9730), .A(n9707), .B(n9706), .ZN(n9712)
         );
  INV_X1 U10917 ( .A(n9709), .ZN(n9722) );
  OAI211_X1 U10918 ( .C1(n10205), .C2(n9722), .A(n9710), .B(n9746), .ZN(n10145) );
  NOR2_X1 U10919 ( .A1(n10145), .A2(n9755), .ZN(n9711) );
  AOI211_X1 U10920 ( .C1(n9751), .C2(n9713), .A(n9712), .B(n9711), .ZN(n9714)
         );
  OAI211_X1 U10921 ( .C1(n10147), .C2(n9736), .A(n9715), .B(n9714), .ZN(
        P1_U3277) );
  INV_X1 U10922 ( .A(n9716), .ZN(n9717) );
  AOI21_X1 U10923 ( .B1(n9720), .B2(n9718), .A(n9717), .ZN(n10251) );
  XNOR2_X1 U10924 ( .A(n9719), .B(n9720), .ZN(n10253) );
  NAND2_X1 U10925 ( .A1(n10253), .A2(n9721), .ZN(n9735) );
  AOI211_X1 U10926 ( .C1(n10247), .C2(n9745), .A(n9723), .B(n9722), .ZN(n10245) );
  NOR2_X1 U10927 ( .A1(n9725), .A2(n9724), .ZN(n9732) );
  NAND2_X1 U10928 ( .A1(n9726), .A2(n10153), .ZN(n9729) );
  AOI22_X1 U10929 ( .A1(n9750), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9727), .B2(
        n9748), .ZN(n9728) );
  OAI211_X1 U10930 ( .C1(n10242), .C2(n9730), .A(n9729), .B(n9728), .ZN(n9731)
         );
  AOI211_X1 U10931 ( .C1(n10245), .C2(n9733), .A(n9732), .B(n9731), .ZN(n9734)
         );
  OAI211_X1 U10932 ( .C1(n10251), .C2(n9736), .A(n9735), .B(n9734), .ZN(
        P1_U3278) );
  XNOR2_X1 U10933 ( .A(n9737), .B(n6262), .ZN(n10303) );
  INV_X1 U10934 ( .A(n10303), .ZN(n9760) );
  NAND2_X1 U10935 ( .A1(n9739), .A2(n9738), .ZN(n9740) );
  NAND3_X1 U10936 ( .A1(n9741), .A2(n10125), .A3(n9740), .ZN(n9744) );
  AOI22_X1 U10937 ( .A1(n10155), .A2(n9742), .B1(n10144), .B2(n10152), .ZN(
        n9743) );
  NAND2_X1 U10938 ( .A1(n9744), .A2(n9743), .ZN(n10301) );
  OAI211_X1 U10939 ( .C1(n9747), .C2(n9476), .A(n9746), .B(n9745), .ZN(n10298)
         );
  AOI22_X1 U10940 ( .A1(n9750), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9749), .B2(
        n9748), .ZN(n9754) );
  NAND2_X1 U10941 ( .A1(n9752), .A2(n9751), .ZN(n9753) );
  OAI211_X1 U10942 ( .C1(n10298), .C2(n9755), .A(n9754), .B(n9753), .ZN(n9756)
         );
  AOI21_X1 U10943 ( .B1(n10301), .B2(n9757), .A(n9756), .ZN(n9758) );
  OAI21_X1 U10944 ( .B1(n9760), .B2(n9759), .A(n9758), .ZN(P1_U3279) );
  OAI211_X1 U10945 ( .C1(n9445), .C2(n10299), .A(n9761), .B(n10047), .ZN(
        n10164) );
  INV_X1 U10946 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10257) );
  AOI22_X1 U10947 ( .A1(n10257), .A2(keyinput53), .B1(n5653), .B2(keyinput71), 
        .ZN(n9762) );
  OAI221_X1 U10948 ( .B1(n10257), .B2(keyinput53), .C1(n5653), .C2(keyinput71), 
        .A(n9762), .ZN(n9770) );
  INV_X1 U10949 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9961) );
  AOI22_X1 U10950 ( .A1(n9961), .A2(keyinput38), .B1(n9764), .B2(keyinput10), 
        .ZN(n9763) );
  OAI221_X1 U10951 ( .B1(n9961), .B2(keyinput38), .C1(n9764), .C2(keyinput10), 
        .A(n9763), .ZN(n9769) );
  INV_X1 U10952 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10262) );
  AOI22_X1 U10953 ( .A1(n9987), .A2(keyinput79), .B1(n10262), .B2(keyinput25), 
        .ZN(n9765) );
  OAI221_X1 U10954 ( .B1(n9987), .B2(keyinput79), .C1(n10262), .C2(keyinput25), 
        .A(n9765), .ZN(n9768) );
  AOI22_X1 U10955 ( .A1(n7042), .A2(keyinput59), .B1(n9967), .B2(keyinput95), 
        .ZN(n9766) );
  OAI221_X1 U10956 ( .B1(n7042), .B2(keyinput59), .C1(n9967), .C2(keyinput95), 
        .A(n9766), .ZN(n9767) );
  OR4_X1 U10957 ( .A1(n9770), .A2(n9769), .A3(n9768), .A4(n9767), .ZN(n9782)
         );
  INV_X1 U10958 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10260) );
  AOI22_X1 U10959 ( .A1(n10260), .A2(keyinput107), .B1(n5959), .B2(keyinput123), .ZN(n9771) );
  OAI221_X1 U10960 ( .B1(n10260), .B2(keyinput107), .C1(n5959), .C2(
        keyinput123), .A(n9771), .ZN(n9781) );
  XNOR2_X1 U10961 ( .A(n9772), .B(keyinput115), .ZN(n9780) );
  XOR2_X1 U10962 ( .A(n9773), .B(keyinput90), .Z(n9778) );
  XOR2_X1 U10963 ( .A(n10009), .B(keyinput45), .Z(n9777) );
  INV_X1 U10964 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10369) );
  XOR2_X1 U10965 ( .A(n10369), .B(keyinput54), .Z(n9776) );
  INV_X1 U10966 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9774) );
  XOR2_X1 U10967 ( .A(n9774), .B(keyinput69), .Z(n9775) );
  NAND4_X1 U10968 ( .A1(n9778), .A2(n9777), .A3(n9776), .A4(n9775), .ZN(n9779)
         );
  OR4_X1 U10969 ( .A1(n9782), .A2(n9781), .A3(n9780), .A4(n9779), .ZN(n9921)
         );
  INV_X1 U10970 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10255) );
  AOI22_X1 U10971 ( .A1(n10255), .A2(keyinput78), .B1(n9784), .B2(keyinput106), 
        .ZN(n9783) );
  OAI221_X1 U10972 ( .B1(n10255), .B2(keyinput78), .C1(n9784), .C2(keyinput106), .A(n9783), .ZN(n9790) );
  AOI22_X1 U10973 ( .A1(n9786), .A2(keyinput48), .B1(n9988), .B2(keyinput1), 
        .ZN(n9785) );
  OAI221_X1 U10974 ( .B1(n9786), .B2(keyinput48), .C1(n9988), .C2(keyinput1), 
        .A(n9785), .ZN(n9789) );
  XNOR2_X1 U10975 ( .A(keyinput98), .B(n10161), .ZN(n9788) );
  XNOR2_X1 U10976 ( .A(keyinput86), .B(n9965), .ZN(n9787) );
  OR4_X1 U10977 ( .A1(n9790), .A2(n9789), .A3(n9788), .A4(n9787), .ZN(n9798)
         );
  INV_X1 U10978 ( .A(keyinput24), .ZN(n9792) );
  AOI22_X1 U10979 ( .A1(n9793), .A2(keyinput117), .B1(P2_ADDR_REG_10__SCAN_IN), 
        .B2(n9792), .ZN(n9791) );
  OAI221_X1 U10980 ( .B1(n9793), .B2(keyinput117), .C1(n9792), .C2(
        P2_ADDR_REG_10__SCAN_IN), .A(n9791), .ZN(n9797) );
  INV_X1 U10981 ( .A(keyinput15), .ZN(n9795) );
  AOI22_X1 U10982 ( .A1(n9409), .A2(keyinput43), .B1(P2_ADDR_REG_18__SCAN_IN), 
        .B2(n9795), .ZN(n9794) );
  OAI221_X1 U10983 ( .B1(n9409), .B2(keyinput43), .C1(n9795), .C2(
        P2_ADDR_REG_18__SCAN_IN), .A(n9794), .ZN(n9796) );
  NOR3_X1 U10984 ( .A1(n9798), .A2(n9797), .A3(n9796), .ZN(n9842) );
  INV_X1 U10985 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9800) );
  INV_X1 U10986 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10357) );
  AOI22_X1 U10987 ( .A1(n9800), .A2(keyinput119), .B1(n10357), .B2(keyinput104), .ZN(n9799) );
  OAI221_X1 U10988 ( .B1(n9800), .B2(keyinput119), .C1(n10357), .C2(
        keyinput104), .A(n9799), .ZN(n9807) );
  AOI22_X1 U10989 ( .A1(n9802), .A2(keyinput105), .B1(n9972), .B2(keyinput85), 
        .ZN(n9801) );
  OAI221_X1 U10990 ( .B1(n9802), .B2(keyinput105), .C1(n9972), .C2(keyinput85), 
        .A(n9801), .ZN(n9806) );
  AOI22_X1 U10991 ( .A1(n9804), .A2(keyinput63), .B1(n9997), .B2(keyinput29), 
        .ZN(n9803) );
  OAI221_X1 U10992 ( .B1(n9804), .B2(keyinput63), .C1(n9997), .C2(keyinput29), 
        .A(n9803), .ZN(n9805) );
  OR3_X1 U10993 ( .A1(n9807), .A2(n9806), .A3(n9805), .ZN(n9814) );
  INV_X1 U10994 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n9809) );
  AOI22_X1 U10995 ( .A1(n9809), .A2(keyinput39), .B1(n10030), .B2(keyinput116), 
        .ZN(n9808) );
  OAI221_X1 U10996 ( .B1(n9809), .B2(keyinput39), .C1(n10030), .C2(keyinput116), .A(n9808), .ZN(n9813) );
  AOI22_X1 U10997 ( .A1(n10003), .A2(keyinput18), .B1(n9811), .B2(keyinput126), 
        .ZN(n9810) );
  OAI221_X1 U10998 ( .B1(n10003), .B2(keyinput18), .C1(n9811), .C2(keyinput126), .A(n9810), .ZN(n9812) );
  NOR3_X1 U10999 ( .A1(n9814), .A2(n9813), .A3(n9812), .ZN(n9841) );
  INV_X1 U11000 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10259) );
  AOI22_X1 U11001 ( .A1(n9816), .A2(keyinput49), .B1(keyinput23), .B2(n10259), 
        .ZN(n9815) );
  OAI221_X1 U11002 ( .B1(n9816), .B2(keyinput49), .C1(n10259), .C2(keyinput23), 
        .A(n9815), .ZN(n9827) );
  INV_X1 U11003 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10341) );
  AOI22_X1 U11004 ( .A1(n9818), .A2(keyinput80), .B1(keyinput41), .B2(n10341), 
        .ZN(n9817) );
  OAI221_X1 U11005 ( .B1(n9818), .B2(keyinput80), .C1(n10341), .C2(keyinput41), 
        .A(n9817), .ZN(n9826) );
  AOI22_X1 U11006 ( .A1(n9820), .A2(keyinput65), .B1(keyinput94), .B2(n6141), 
        .ZN(n9819) );
  OAI221_X1 U11007 ( .B1(n9820), .B2(keyinput65), .C1(n6141), .C2(keyinput94), 
        .A(n9819), .ZN(n9825) );
  INV_X1 U11008 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9822) );
  AOI22_X1 U11009 ( .A1(n9823), .A2(keyinput113), .B1(keyinput83), .B2(n9822), 
        .ZN(n9821) );
  OAI221_X1 U11010 ( .B1(n9823), .B2(keyinput113), .C1(n9822), .C2(keyinput83), 
        .A(n9821), .ZN(n9824) );
  NOR4_X1 U11011 ( .A1(n9827), .A2(n9826), .A3(n9825), .A4(n9824), .ZN(n9840)
         );
  INV_X1 U11012 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9829) );
  AOI22_X1 U11013 ( .A1(n9829), .A2(keyinput76), .B1(n9981), .B2(keyinput4), 
        .ZN(n9828) );
  OAI221_X1 U11014 ( .B1(n9829), .B2(keyinput76), .C1(n9981), .C2(keyinput4), 
        .A(n9828), .ZN(n9838) );
  AOI22_X1 U11015 ( .A1(n10016), .A2(keyinput93), .B1(keyinput16), .B2(n9831), 
        .ZN(n9830) );
  OAI221_X1 U11016 ( .B1(n10016), .B2(keyinput93), .C1(n9831), .C2(keyinput16), 
        .A(n9830), .ZN(n9837) );
  INV_X1 U11017 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10261) );
  AOI22_X1 U11018 ( .A1(n10261), .A2(keyinput9), .B1(keyinput6), .B2(n7223), 
        .ZN(n9832) );
  OAI221_X1 U11019 ( .B1(n10261), .B2(keyinput9), .C1(n7223), .C2(keyinput6), 
        .A(n9832), .ZN(n9836) );
  AOI22_X1 U11020 ( .A1(n9834), .A2(keyinput97), .B1(keyinput32), .B2(n6688), 
        .ZN(n9833) );
  OAI221_X1 U11021 ( .B1(n9834), .B2(keyinput97), .C1(n6688), .C2(keyinput32), 
        .A(n9833), .ZN(n9835) );
  NOR4_X1 U11022 ( .A1(n9838), .A2(n9837), .A3(n9836), .A4(n9835), .ZN(n9839)
         );
  NAND4_X1 U11023 ( .A1(n9842), .A2(n9841), .A3(n9840), .A4(n9839), .ZN(n9920)
         );
  AOI22_X1 U11024 ( .A1(n5545), .A2(keyinput37), .B1(keyinput44), .B2(n9968), 
        .ZN(n9843) );
  OAI221_X1 U11025 ( .B1(n5545), .B2(keyinput37), .C1(n9968), .C2(keyinput44), 
        .A(n9843), .ZN(n9851) );
  AOI22_X1 U11026 ( .A1(n9845), .A2(keyinput12), .B1(keyinput3), .B2(n8076), 
        .ZN(n9844) );
  OAI221_X1 U11027 ( .B1(n9845), .B2(keyinput12), .C1(n8076), .C2(keyinput3), 
        .A(n9844), .ZN(n9850) );
  INV_X1 U11028 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10374) );
  AOI22_X1 U11029 ( .A1(n10374), .A2(keyinput60), .B1(keyinput19), .B2(n7255), 
        .ZN(n9846) );
  OAI221_X1 U11030 ( .B1(n10374), .B2(keyinput60), .C1(n7255), .C2(keyinput19), 
        .A(n9846), .ZN(n9849) );
  XNOR2_X1 U11031 ( .A(n9847), .B(keyinput91), .ZN(n9848) );
  NOR4_X1 U11032 ( .A1(n9851), .A2(n9850), .A3(n9849), .A4(n9848), .ZN(n9873)
         );
  AOI22_X1 U11033 ( .A1(n9853), .A2(keyinput111), .B1(keyinput8), .B2(n10379), 
        .ZN(n9852) );
  OAI221_X1 U11034 ( .B1(n9853), .B2(keyinput111), .C1(n10379), .C2(keyinput8), 
        .A(n9852), .ZN(n9858) );
  AOI22_X1 U11035 ( .A1(n9856), .A2(keyinput82), .B1(keyinput58), .B2(n9855), 
        .ZN(n9854) );
  OAI221_X1 U11036 ( .B1(n9856), .B2(keyinput82), .C1(n9855), .C2(keyinput58), 
        .A(n9854), .ZN(n9857) );
  NOR2_X1 U11037 ( .A1(n9858), .A2(n9857), .ZN(n9872) );
  INV_X1 U11038 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n9960) );
  AOI22_X1 U11039 ( .A1(n9960), .A2(keyinput55), .B1(n9980), .B2(keyinput40), 
        .ZN(n9859) );
  OAI221_X1 U11040 ( .B1(n9960), .B2(keyinput55), .C1(n9980), .C2(keyinput40), 
        .A(n9859), .ZN(n9870) );
  INV_X1 U11041 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10258) );
  AOI22_X1 U11042 ( .A1(n10258), .A2(keyinput62), .B1(n9991), .B2(keyinput47), 
        .ZN(n9860) );
  OAI221_X1 U11043 ( .B1(n10258), .B2(keyinput62), .C1(n9991), .C2(keyinput47), 
        .A(n9860), .ZN(n9869) );
  INV_X1 U11044 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9862) );
  AOI22_X1 U11045 ( .A1(n9862), .A2(keyinput36), .B1(n9986), .B2(keyinput22), 
        .ZN(n9861) );
  OAI221_X1 U11046 ( .B1(n9862), .B2(keyinput36), .C1(n9986), .C2(keyinput22), 
        .A(n9861), .ZN(n9868) );
  XNOR2_X1 U11047 ( .A(SI_29_), .B(keyinput110), .ZN(n9866) );
  XNOR2_X1 U11048 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput99), .ZN(n9865) );
  XNOR2_X1 U11049 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput66), .ZN(n9864) );
  XNOR2_X1 U11050 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput27), .ZN(n9863) );
  NAND4_X1 U11051 ( .A1(n9866), .A2(n9865), .A3(n9864), .A4(n9863), .ZN(n9867)
         );
  NOR4_X1 U11052 ( .A1(n9870), .A2(n9869), .A3(n9868), .A4(n9867), .ZN(n9871)
         );
  NAND3_X1 U11053 ( .A1(n9873), .A2(n9872), .A3(n9871), .ZN(n9919) );
  XNOR2_X1 U11054 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(keyinput68), .ZN(n9877)
         );
  XNOR2_X1 U11055 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(keyinput0), .ZN(n9876) );
  XNOR2_X1 U11056 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(keyinput21), .ZN(n9875) );
  XNOR2_X1 U11057 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput87), .ZN(n9874) );
  NAND4_X1 U11058 ( .A1(n9877), .A2(n9876), .A3(n9875), .A4(n9874), .ZN(n9883)
         );
  XNOR2_X1 U11059 ( .A(P1_REG2_REG_2__SCAN_IN), .B(keyinput31), .ZN(n9881) );
  XNOR2_X1 U11060 ( .A(P1_REG0_REG_16__SCAN_IN), .B(keyinput2), .ZN(n9880) );
  XNOR2_X1 U11061 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(keyinput108), .ZN(n9879)
         );
  XNOR2_X1 U11062 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput81), .ZN(n9878) );
  NAND4_X1 U11063 ( .A1(n9881), .A2(n9880), .A3(n9879), .A4(n9878), .ZN(n9882)
         );
  NOR2_X1 U11064 ( .A1(n9883), .A2(n9882), .ZN(n9917) );
  XNOR2_X1 U11065 ( .A(P2_IR_REG_10__SCAN_IN), .B(keyinput109), .ZN(n9887) );
  XNOR2_X1 U11066 ( .A(P2_IR_REG_24__SCAN_IN), .B(keyinput72), .ZN(n9886) );
  XNOR2_X1 U11067 ( .A(P2_REG1_REG_18__SCAN_IN), .B(keyinput84), .ZN(n9885) );
  XNOR2_X1 U11068 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput75), .ZN(n9884) );
  NAND4_X1 U11069 ( .A1(n9887), .A2(n9886), .A3(n9885), .A4(n9884), .ZN(n9893)
         );
  XNOR2_X1 U11070 ( .A(P2_IR_REG_29__SCAN_IN), .B(keyinput34), .ZN(n9891) );
  XNOR2_X1 U11071 ( .A(P2_IR_REG_22__SCAN_IN), .B(keyinput33), .ZN(n9890) );
  XNOR2_X1 U11072 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput57), .ZN(n9889) );
  XNOR2_X1 U11073 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput92), .ZN(n9888) );
  NAND4_X1 U11074 ( .A1(n9891), .A2(n9890), .A3(n9889), .A4(n9888), .ZN(n9892)
         );
  NOR2_X1 U11075 ( .A1(n9893), .A2(n9892), .ZN(n9916) );
  XNOR2_X1 U11076 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(keyinput89), .ZN(n9897)
         );
  XNOR2_X1 U11077 ( .A(P1_REG0_REG_26__SCAN_IN), .B(keyinput112), .ZN(n9896)
         );
  XNOR2_X1 U11078 ( .A(P2_IR_REG_0__SCAN_IN), .B(keyinput67), .ZN(n9895) );
  XNOR2_X1 U11079 ( .A(P2_IR_REG_20__SCAN_IN), .B(keyinput88), .ZN(n9894) );
  NAND4_X1 U11080 ( .A1(n9897), .A2(n9896), .A3(n9895), .A4(n9894), .ZN(n9903)
         );
  XNOR2_X1 U11081 ( .A(P2_IR_REG_5__SCAN_IN), .B(keyinput46), .ZN(n9901) );
  XNOR2_X1 U11082 ( .A(P2_IR_REG_3__SCAN_IN), .B(keyinput17), .ZN(n9900) );
  XNOR2_X1 U11083 ( .A(SI_4_), .B(keyinput28), .ZN(n9899) );
  XNOR2_X1 U11084 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput52), .ZN(n9898) );
  NAND4_X1 U11085 ( .A1(n9901), .A2(n9900), .A3(n9899), .A4(n9898), .ZN(n9902)
         );
  NOR2_X1 U11086 ( .A1(n9903), .A2(n9902), .ZN(n9915) );
  XNOR2_X1 U11087 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput61), .ZN(n9907) );
  XNOR2_X1 U11088 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput125), .ZN(n9906) );
  XNOR2_X1 U11089 ( .A(P2_D_REG_0__SCAN_IN), .B(keyinput114), .ZN(n9905) );
  XNOR2_X1 U11090 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput122), .ZN(n9904) );
  NAND4_X1 U11091 ( .A1(n9907), .A2(n9906), .A3(n9905), .A4(n9904), .ZN(n9913)
         );
  XNOR2_X1 U11092 ( .A(P2_IR_REG_14__SCAN_IN), .B(keyinput127), .ZN(n9911) );
  XNOR2_X1 U11093 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput30), .ZN(n9910) );
  XNOR2_X1 U11094 ( .A(P2_IR_REG_28__SCAN_IN), .B(keyinput96), .ZN(n9909) );
  XNOR2_X1 U11095 ( .A(keyinput124), .B(P2_REG2_REG_7__SCAN_IN), .ZN(n9908) );
  NAND4_X1 U11096 ( .A1(n9911), .A2(n9910), .A3(n9909), .A4(n9908), .ZN(n9912)
         );
  NOR2_X1 U11097 ( .A1(n9913), .A2(n9912), .ZN(n9914) );
  NAND4_X1 U11098 ( .A1(n9917), .A2(n9916), .A3(n9915), .A4(n9914), .ZN(n9918)
         );
  NOR4_X1 U11099 ( .A1(n9921), .A2(n9920), .A3(n9919), .A4(n9918), .ZN(n9959)
         );
  INV_X1 U11100 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10263) );
  AOI22_X1 U11101 ( .A1(n10263), .A2(keyinput20), .B1(n9996), .B2(keyinput42), 
        .ZN(n9922) );
  OAI221_X1 U11102 ( .B1(n10263), .B2(keyinput20), .C1(n9996), .C2(keyinput42), 
        .A(n9922), .ZN(n9932) );
  INV_X1 U11103 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n9995) );
  INV_X1 U11104 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n10199) );
  AOI22_X1 U11105 ( .A1(n9995), .A2(keyinput74), .B1(n10199), .B2(keyinput13), 
        .ZN(n9923) );
  OAI221_X1 U11106 ( .B1(n9995), .B2(keyinput74), .C1(n10199), .C2(keyinput13), 
        .A(n9923), .ZN(n9931) );
  AOI22_X1 U11107 ( .A1(n9925), .A2(keyinput56), .B1(P2_U3151), .B2(
        keyinput120), .ZN(n9924) );
  OAI221_X1 U11108 ( .B1(n9925), .B2(keyinput56), .C1(P2_U3151), .C2(
        keyinput120), .A(n9924), .ZN(n9930) );
  INV_X1 U11109 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9928) );
  INV_X1 U11110 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9927) );
  AOI22_X1 U11111 ( .A1(n9928), .A2(keyinput101), .B1(n9927), .B2(keyinput51), 
        .ZN(n9926) );
  OAI221_X1 U11112 ( .B1(n9928), .B2(keyinput101), .C1(n9927), .C2(keyinput51), 
        .A(n9926), .ZN(n9929) );
  NOR4_X1 U11113 ( .A1(n9932), .A2(n9931), .A3(n9930), .A4(n9929), .ZN(n9958)
         );
  INV_X1 U11114 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10207) );
  AOI22_X1 U11115 ( .A1(n9934), .A2(keyinput50), .B1(keyinput26), .B2(n10207), 
        .ZN(n9933) );
  OAI221_X1 U11116 ( .B1(n9934), .B2(keyinput50), .C1(n10207), .C2(keyinput26), 
        .A(n9933), .ZN(n9944) );
  AOI22_X1 U11117 ( .A1(n9937), .A2(keyinput100), .B1(keyinput77), .B2(n9936), 
        .ZN(n9935) );
  OAI221_X1 U11118 ( .B1(n9937), .B2(keyinput100), .C1(n9936), .C2(keyinput77), 
        .A(n9935), .ZN(n9943) );
  AOI22_X1 U11119 ( .A1(n10033), .A2(keyinput11), .B1(n10031), .B2(keyinput5), 
        .ZN(n9938) );
  OAI221_X1 U11120 ( .B1(n10033), .B2(keyinput11), .C1(n10031), .C2(keyinput5), 
        .A(n9938), .ZN(n9942) );
  AOI22_X1 U11121 ( .A1(n9940), .A2(keyinput35), .B1(n10032), .B2(keyinput70), 
        .ZN(n9939) );
  OAI221_X1 U11122 ( .B1(n9940), .B2(keyinput35), .C1(n10032), .C2(keyinput70), 
        .A(n9939), .ZN(n9941) );
  NOR4_X1 U11123 ( .A1(n9944), .A2(n9943), .A3(n9942), .A4(n9941), .ZN(n9957)
         );
  INV_X1 U11124 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10355) );
  AOI22_X1 U11125 ( .A1(n10028), .A2(keyinput118), .B1(keyinput7), .B2(n10355), 
        .ZN(n9945) );
  OAI221_X1 U11126 ( .B1(n10028), .B2(keyinput118), .C1(n10355), .C2(keyinput7), .A(n9945), .ZN(n9955) );
  AOI22_X1 U11127 ( .A1(n9990), .A2(keyinput103), .B1(keyinput14), .B2(n10189), 
        .ZN(n9946) );
  OAI221_X1 U11128 ( .B1(n9990), .B2(keyinput103), .C1(n10189), .C2(keyinput14), .A(n9946), .ZN(n9954) );
  INV_X1 U11129 ( .A(keyinput64), .ZN(n9948) );
  AOI22_X1 U11130 ( .A1(n9949), .A2(keyinput102), .B1(P1_ADDR_REG_17__SCAN_IN), 
        .B2(n9948), .ZN(n9947) );
  OAI221_X1 U11131 ( .B1(n9949), .B2(keyinput102), .C1(n9948), .C2(
        P1_ADDR_REG_17__SCAN_IN), .A(n9947), .ZN(n9953) );
  AOI22_X1 U11132 ( .A1(n7825), .A2(keyinput121), .B1(keyinput73), .B2(n9951), 
        .ZN(n9950) );
  OAI221_X1 U11133 ( .B1(n7825), .B2(keyinput121), .C1(n9951), .C2(keyinput73), 
        .A(n9950), .ZN(n9952) );
  NOR4_X1 U11134 ( .A1(n9955), .A2(n9954), .A3(n9953), .A4(n9952), .ZN(n9956)
         );
  NAND4_X1 U11135 ( .A1(n9959), .A2(n9958), .A3(n9957), .A4(n9956), .ZN(n10044) );
  NOR4_X1 U11136 ( .A1(P2_B_REG_SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), .A3(
        n6141), .A4(n9960), .ZN(n9964) );
  INV_X1 U11137 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9962) );
  NOR4_X1 U11138 ( .A1(P2_REG0_REG_1__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), 
        .A3(n9962), .A4(n9961), .ZN(n9963) );
  NAND2_X1 U11139 ( .A1(n9964), .A2(n9963), .ZN(n10027) );
  NAND4_X1 U11140 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        n9965), .A4(n10161), .ZN(n9966) );
  NOR3_X1 U11141 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(P2_ADDR_REG_14__SCAN_IN), 
        .A3(n9966), .ZN(n9975) );
  NAND4_X1 U11142 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_REG0_REG_3__SCAN_IN), 
        .A3(P2_REG1_REG_10__SCAN_IN), .A4(n5959), .ZN(n9971) );
  NAND4_X1 U11143 ( .A1(P2_REG2_REG_29__SCAN_IN), .A2(P2_REG1_REG_9__SCAN_IN), 
        .A3(P1_REG3_REG_3__SCAN_IN), .A4(n9967), .ZN(n9970) );
  NAND4_X1 U11144 ( .A1(P2_REG2_REG_26__SCAN_IN), .A2(P2_REG2_REG_10__SCAN_IN), 
        .A3(P1_REG0_REG_26__SCAN_IN), .A4(n9968), .ZN(n9969) );
  NOR4_X1 U11145 ( .A1(n9972), .A2(n9971), .A3(n9970), .A4(n9969), .ZN(n9973)
         );
  AND4_X1 U11146 ( .A1(n9973), .A2(P1_REG0_REG_16__SCAN_IN), .A3(
        P1_REG1_REG_23__SCAN_IN), .A4(n6096), .ZN(n9974) );
  AND4_X1 U11147 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_REG1_REG_18__SCAN_IN), 
        .A3(n9975), .A4(n9974), .ZN(n10025) );
  NOR4_X1 U11148 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P1_REG2_REG_9__SCAN_IN), 
        .A3(P2_ADDR_REG_18__SCAN_IN), .A4(n10255), .ZN(n10024) );
  AND2_X1 U11149 ( .A1(n9976), .A2(SI_4_), .ZN(n10005) );
  NOR4_X1 U11150 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_4__SCAN_IN), 
        .A3(P2_ADDR_REG_8__SCAN_IN), .A4(n10379), .ZN(n9985) );
  NOR4_X1 U11151 ( .A1(P2_STATE_REG_SCAN_IN), .A2(P2_REG1_REG_27__SCAN_IN), 
        .A3(P1_REG2_REG_23__SCAN_IN), .A4(P1_REG0_REG_8__SCAN_IN), .ZN(n9984)
         );
  NOR4_X1 U11152 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n9979), .A3(n9978), .A4(
        n9977), .ZN(n9983) );
  NOR4_X1 U11153 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(P1_REG0_REG_9__SCAN_IN), 
        .A3(n9981), .A4(n9980), .ZN(n9982) );
  AND4_X1 U11154 ( .A1(n9985), .A2(n9984), .A3(n9983), .A4(n9982), .ZN(n10001)
         );
  NOR4_X1 U11155 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P1_REG0_REG_11__SCAN_IN), .A4(n9986), .ZN(n9994) );
  NOR4_X1 U11156 ( .A1(SI_27_), .A2(SI_26_), .A3(n9988), .A4(n9987), .ZN(n9993) );
  NOR4_X1 U11157 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n9991), .A3(n9990), .A4(
        n9989), .ZN(n9992) );
  AND3_X1 U11158 ( .A1(n9994), .A2(n9993), .A3(n9992), .ZN(n10000) );
  NOR4_X1 U11159 ( .A1(P1_REG0_REG_17__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .A3(n9996), .A4(n9995), .ZN(n9999) );
  NOR4_X1 U11160 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(P1_DATAO_REG_15__SCAN_IN), .A3(P1_DATAO_REG_13__SCAN_IN), .A4(n9997), .ZN(n9998) );
  NAND4_X1 U11161 ( .A1(n10001), .A2(n10000), .A3(n9999), .A4(n9998), .ZN(
        n10002) );
  NOR2_X1 U11162 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(n10002), .ZN(n10004) );
  NAND4_X1 U11163 ( .A1(n10005), .A2(P1_D_REG_28__SCAN_IN), .A3(n10004), .A4(
        n10003), .ZN(n10007) );
  NAND4_X1 U11164 ( .A1(P1_D_REG_0__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n10006) );
  NOR2_X1 U11165 ( .A1(n10007), .A2(n10006), .ZN(n10021) );
  INV_X1 U11166 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n10008) );
  NAND4_X1 U11167 ( .A1(n10010), .A2(n10009), .A3(n10008), .A4(
        P1_IR_REG_24__SCAN_IN), .ZN(n10012) );
  NAND4_X1 U11168 ( .A1(SI_29_), .A2(P1_DATAO_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .A4(P2_REG0_REG_0__SCAN_IN), .ZN(n10011) );
  NOR2_X1 U11169 ( .A1(n10012), .A2(n10011), .ZN(n10020) );
  INV_X1 U11170 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n10015) );
  NAND4_X1 U11171 ( .A1(n10015), .A2(n10014), .A3(n10013), .A4(
        P1_IR_REG_13__SCAN_IN), .ZN(n10018) );
  NAND4_X1 U11172 ( .A1(n10016), .A2(n9831), .A3(P1_REG2_REG_7__SCAN_IN), .A4(
        P2_DATAO_REG_2__SCAN_IN), .ZN(n10017) );
  NOR2_X1 U11173 ( .A1(n10018), .A2(n10017), .ZN(n10019) );
  AND4_X1 U11174 ( .A1(n10021), .A2(n10020), .A3(n10019), .A4(n10260), .ZN(
        n10022) );
  NAND4_X1 U11175 ( .A1(n10025), .A2(n10024), .A3(n10023), .A4(n10022), .ZN(
        n10026) );
  NOR2_X1 U11176 ( .A1(n10027), .A2(n10026), .ZN(n10042) );
  NOR4_X1 U11177 ( .A1(P2_IR_REG_29__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .A4(n7223), .ZN(n10041) );
  NAND4_X1 U11178 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(P2_REG0_REG_10__SCAN_IN), 
        .A3(P2_ADDR_REG_13__SCAN_IN), .A4(n10028), .ZN(n10029) );
  NOR3_X1 U11179 ( .A1(P2_REG0_REG_2__SCAN_IN), .A2(P1_REG0_REG_21__SCAN_IN), 
        .A3(n10029), .ZN(n10039) );
  NAND4_X1 U11180 ( .A1(P2_REG0_REG_22__SCAN_IN), .A2(P2_REG2_REG_7__SCAN_IN), 
        .A3(P1_REG3_REG_18__SCAN_IN), .A4(P2_ADDR_REG_10__SCAN_IN), .ZN(n10037) );
  NAND4_X1 U11181 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_REG2_REG_27__SCAN_IN), 
        .A3(n10030), .A4(n10357), .ZN(n10036) );
  NAND4_X1 U11182 ( .A1(P2_D_REG_0__SCAN_IN), .A2(P2_REG0_REG_12__SCAN_IN), 
        .A3(n10032), .A4(n10031), .ZN(n10035) );
  NAND4_X1 U11183 ( .A1(P2_REG1_REG_28__SCAN_IN), .A2(P1_REG3_REG_14__SCAN_IN), 
        .A3(P1_REG0_REG_13__SCAN_IN), .A4(n10033), .ZN(n10034) );
  NOR4_X1 U11184 ( .A1(n10037), .A2(n10036), .A3(n10035), .A4(n10034), .ZN(
        n10038) );
  AND4_X1 U11185 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .A3(n10039), .A4(n10038), .ZN(n10040) );
  NAND3_X1 U11186 ( .A1(n10042), .A2(n10041), .A3(n10040), .ZN(n10043) );
  XNOR2_X1 U11187 ( .A(n10044), .B(n10043), .ZN(n10045) );
  XNOR2_X1 U11188 ( .A(n10046), .B(n10045), .ZN(P1_U3553) );
  INV_X1 U11189 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10049) );
  AND2_X1 U11190 ( .A1(n10048), .A2(n10047), .ZN(n10165) );
  MUX2_X1 U11191 ( .A(n10049), .B(n10165), .S(n10316), .Z(n10050) );
  OAI21_X1 U11192 ( .B1(n10168), .B2(n10163), .A(n10050), .ZN(P1_U3552) );
  NAND2_X1 U11193 ( .A1(n10052), .A2(n10248), .ZN(n10054) );
  OAI211_X1 U11194 ( .C1(n10067), .C2(n10243), .A(n10054), .B(n10053), .ZN(
        n10055) );
  MUX2_X1 U11195 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n10169), .S(n10316), .Z(
        P1_U3551) );
  AOI22_X1 U11196 ( .A1(n10058), .A2(n10152), .B1(n10077), .B2(n10155), .ZN(
        n10060) );
  OAI211_X1 U11197 ( .C1(n10061), .C2(n10250), .A(n10060), .B(n10059), .ZN(
        n10062) );
  MUX2_X1 U11198 ( .A(n10064), .B(n10170), .S(n10316), .Z(n10065) );
  OAI21_X1 U11199 ( .B1(n4839), .B2(n10163), .A(n10065), .ZN(P1_U3550) );
  OAI22_X1 U11200 ( .A1(n10067), .A2(n10241), .B1(n10066), .B2(n10243), .ZN(
        n10068) );
  INV_X1 U11201 ( .A(n10068), .ZN(n10070) );
  OAI211_X1 U11202 ( .C1(n10071), .C2(n10250), .A(n10070), .B(n10069), .ZN(
        n10072) );
  AOI21_X1 U11203 ( .B1(n10073), .B2(n10302), .A(n10072), .ZN(n10173) );
  MUX2_X1 U11204 ( .A(n10074), .B(n10173), .S(n10316), .Z(n10075) );
  OAI21_X1 U11205 ( .B1(n10176), .B2(n10163), .A(n10075), .ZN(P1_U3549) );
  INV_X1 U11206 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n10083) );
  AOI22_X1 U11207 ( .A1(n10077), .A2(n10152), .B1(n10155), .B2(n10076), .ZN(
        n10079) );
  OAI211_X1 U11208 ( .C1(n10080), .C2(n10250), .A(n10079), .B(n10078), .ZN(
        n10081) );
  AOI21_X1 U11209 ( .B1(n10082), .B2(n10302), .A(n10081), .ZN(n10177) );
  MUX2_X1 U11210 ( .A(n10083), .B(n10177), .S(n10316), .Z(n10084) );
  OAI21_X1 U11211 ( .B1(n10180), .B2(n10163), .A(n10084), .ZN(P1_U3548) );
  INV_X1 U11212 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n10092) );
  AOI22_X1 U11213 ( .A1(n10086), .A2(n10152), .B1(n10155), .B2(n10085), .ZN(
        n10088) );
  OAI211_X1 U11214 ( .C1(n10089), .C2(n10250), .A(n10088), .B(n10087), .ZN(
        n10090) );
  AOI21_X1 U11215 ( .B1(n10091), .B2(n10302), .A(n10090), .ZN(n10181) );
  MUX2_X1 U11216 ( .A(n10092), .B(n10181), .S(n10316), .Z(n10093) );
  OAI21_X1 U11217 ( .B1(n10184), .B2(n10163), .A(n10093), .ZN(P1_U3547) );
  INV_X1 U11218 ( .A(n10302), .ZN(n10128) );
  AOI211_X1 U11219 ( .C1(n10248), .C2(n10096), .A(n10095), .B(n10094), .ZN(
        n10097) );
  OAI21_X1 U11220 ( .B1(n10098), .B2(n10128), .A(n10097), .ZN(n10185) );
  MUX2_X1 U11221 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10185), .S(n10316), .Z(
        P1_U3546) );
  AOI21_X1 U11222 ( .B1(n10248), .B2(n10100), .A(n10099), .ZN(n10101) );
  OAI211_X1 U11223 ( .C1(n10103), .C2(n10128), .A(n10102), .B(n10101), .ZN(
        n10186) );
  MUX2_X1 U11224 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10186), .S(n10316), .Z(
        P1_U3545) );
  AOI211_X1 U11225 ( .C1(n10248), .C2(n10106), .A(n10105), .B(n10104), .ZN(
        n10107) );
  OAI21_X1 U11226 ( .B1(n10108), .B2(n10128), .A(n10107), .ZN(n10187) );
  MUX2_X1 U11227 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10187), .S(n10316), .Z(
        P1_U3544) );
  INV_X1 U11228 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n10112) );
  AOI211_X1 U11229 ( .C1(n10111), .C2(n10302), .A(n10110), .B(n10109), .ZN(
        n10188) );
  MUX2_X1 U11230 ( .A(n10112), .B(n10188), .S(n10316), .Z(n10113) );
  OAI21_X1 U11231 ( .B1(n10191), .B2(n10163), .A(n10113), .ZN(P1_U3543) );
  AOI211_X1 U11232 ( .C1(n10248), .C2(n10116), .A(n10115), .B(n10114), .ZN(
        n10117) );
  OAI21_X1 U11233 ( .B1(n10118), .B2(n10128), .A(n10117), .ZN(n10192) );
  MUX2_X1 U11234 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10192), .S(n10316), .Z(
        P1_U3542) );
  AOI22_X1 U11235 ( .A1(n10120), .A2(n10152), .B1(n10155), .B2(n10119), .ZN(
        n10121) );
  OAI211_X1 U11236 ( .C1(n10123), .C2(n10299), .A(n10122), .B(n10121), .ZN(
        n10124) );
  AOI21_X1 U11237 ( .B1(n10126), .B2(n10125), .A(n10124), .ZN(n10127) );
  OAI21_X1 U11238 ( .B1(n10129), .B2(n10128), .A(n10127), .ZN(n10193) );
  MUX2_X1 U11239 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10193), .S(n10316), .Z(
        P1_U3541) );
  INV_X1 U11240 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10136) );
  AOI22_X1 U11241 ( .A1(n10130), .A2(n10152), .B1(n10155), .B2(n10143), .ZN(
        n10132) );
  OAI211_X1 U11242 ( .C1(n10133), .C2(n10250), .A(n10132), .B(n10131), .ZN(
        n10134) );
  AOI21_X1 U11243 ( .B1(n10135), .B2(n10302), .A(n10134), .ZN(n10194) );
  MUX2_X1 U11244 ( .A(n10136), .B(n10194), .S(n10316), .Z(n10137) );
  OAI21_X1 U11245 ( .B1(n10197), .B2(n10163), .A(n10137), .ZN(P1_U3540) );
  INV_X1 U11246 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10141) );
  AOI211_X1 U11247 ( .C1(n10140), .C2(n10302), .A(n10139), .B(n10138), .ZN(
        n10198) );
  MUX2_X1 U11248 ( .A(n10141), .B(n10198), .S(n10316), .Z(n10142) );
  OAI21_X1 U11249 ( .B1(n10201), .B2(n10163), .A(n10142), .ZN(P1_U3539) );
  INV_X1 U11250 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n10150) );
  AOI22_X1 U11251 ( .A1(n10155), .A2(n10144), .B1(n10143), .B2(n10152), .ZN(
        n10146) );
  OAI211_X1 U11252 ( .C1(n10147), .C2(n10250), .A(n10146), .B(n10145), .ZN(
        n10148) );
  AOI21_X1 U11253 ( .B1(n10149), .B2(n10302), .A(n10148), .ZN(n10202) );
  MUX2_X1 U11254 ( .A(n10150), .B(n10202), .S(n10316), .Z(n10151) );
  OAI21_X1 U11255 ( .B1(n10205), .B2(n10163), .A(n10151), .ZN(P1_U3538) );
  AOI22_X1 U11256 ( .A1(n10155), .A2(n10154), .B1(n10153), .B2(n10152), .ZN(
        n10157) );
  OAI211_X1 U11257 ( .C1(n10158), .C2(n10250), .A(n10157), .B(n10156), .ZN(
        n10159) );
  AOI21_X1 U11258 ( .B1(n10160), .B2(n10302), .A(n10159), .ZN(n10206) );
  MUX2_X1 U11259 ( .A(n10161), .B(n10206), .S(n10316), .Z(n10162) );
  OAI21_X1 U11260 ( .B1(n10210), .B2(n10163), .A(n10162), .ZN(P1_U3535) );
  MUX2_X1 U11261 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n10164), .S(n10306), .Z(
        P1_U3521) );
  INV_X1 U11262 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10166) );
  MUX2_X1 U11263 ( .A(n10166), .B(n10165), .S(n10306), .Z(n10167) );
  OAI21_X1 U11264 ( .B1(n10168), .B2(n10209), .A(n10167), .ZN(P1_U3520) );
  MUX2_X1 U11265 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n10169), .S(n10306), .Z(
        P1_U3519) );
  INV_X1 U11266 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n10171) );
  MUX2_X1 U11267 ( .A(n10171), .B(n10170), .S(n10306), .Z(n10172) );
  OAI21_X1 U11268 ( .B1(n4839), .B2(n10209), .A(n10172), .ZN(P1_U3518) );
  INV_X1 U11269 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n10174) );
  MUX2_X1 U11270 ( .A(n10174), .B(n10173), .S(n10306), .Z(n10175) );
  OAI21_X1 U11271 ( .B1(n10176), .B2(n10209), .A(n10175), .ZN(P1_U3517) );
  MUX2_X1 U11272 ( .A(n10178), .B(n10177), .S(n10306), .Z(n10179) );
  OAI21_X1 U11273 ( .B1(n10180), .B2(n10209), .A(n10179), .ZN(P1_U3516) );
  INV_X1 U11274 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n10182) );
  MUX2_X1 U11275 ( .A(n10182), .B(n10181), .S(n10306), .Z(n10183) );
  OAI21_X1 U11276 ( .B1(n10184), .B2(n10209), .A(n10183), .ZN(P1_U3515) );
  MUX2_X1 U11277 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10185), .S(n10306), .Z(
        P1_U3514) );
  MUX2_X1 U11278 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10186), .S(n10306), .Z(
        P1_U3513) );
  MUX2_X1 U11279 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10187), .S(n10306), .Z(
        P1_U3512) );
  MUX2_X1 U11280 ( .A(n10189), .B(n10188), .S(n10306), .Z(n10190) );
  OAI21_X1 U11281 ( .B1(n10191), .B2(n10209), .A(n10190), .ZN(P1_U3511) );
  MUX2_X1 U11282 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10192), .S(n10306), .Z(
        P1_U3510) );
  MUX2_X1 U11283 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10193), .S(n10306), .Z(
        P1_U3509) );
  MUX2_X1 U11284 ( .A(n10195), .B(n10194), .S(n10306), .Z(n10196) );
  OAI21_X1 U11285 ( .B1(n10197), .B2(n10209), .A(n10196), .ZN(P1_U3507) );
  MUX2_X1 U11286 ( .A(n10199), .B(n10198), .S(n10306), .Z(n10200) );
  OAI21_X1 U11287 ( .B1(n10201), .B2(n10209), .A(n10200), .ZN(P1_U3504) );
  INV_X1 U11288 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10203) );
  MUX2_X1 U11289 ( .A(n10203), .B(n10202), .S(n10306), .Z(n10204) );
  OAI21_X1 U11290 ( .B1(n10205), .B2(n10209), .A(n10204), .ZN(P1_U3501) );
  MUX2_X1 U11291 ( .A(n10207), .B(n10206), .S(n10306), .Z(n10208) );
  OAI21_X1 U11292 ( .B1(n10210), .B2(n10209), .A(n10208), .ZN(P1_U3492) );
  MUX2_X1 U11293 ( .A(n10211), .B(P1_D_REG_1__SCAN_IN), .S(n10265), .Z(
        P1_U3440) );
  MUX2_X1 U11294 ( .A(n10212), .B(P1_D_REG_0__SCAN_IN), .S(n10265), .Z(
        P1_U3439) );
  NOR4_X1 U11295 ( .A1(n5990), .A2(P1_IR_REG_30__SCAN_IN), .A3(n10213), .A4(
        P1_U3086), .ZN(n10214) );
  AOI21_X1 U11296 ( .B1(n10215), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n10214), 
        .ZN(n10216) );
  OAI21_X1 U11297 ( .B1(n10217), .B2(n10222), .A(n10216), .ZN(P1_U3324) );
  OAI222_X1 U11298 ( .A1(n10225), .A2(n10220), .B1(P1_U3086), .B2(n10219), 
        .C1(n10222), .C2(n10218), .ZN(P1_U3326) );
  OAI222_X1 U11299 ( .A1(n10225), .A2(n10224), .B1(P1_U3086), .B2(n10223), 
        .C1(n10222), .C2(n10221), .ZN(P1_U3328) );
  MUX2_X1 U11300 ( .A(n10227), .B(n10226), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3355) );
  INV_X1 U11301 ( .A(n10228), .ZN(n10232) );
  INV_X1 U11302 ( .A(n10229), .ZN(n10230) );
  OAI22_X1 U11303 ( .A1(n10232), .A2(n10231), .B1(n10230), .B2(n10345), .ZN(
        n10234) );
  AOI211_X1 U11304 ( .C1(n10236), .C2(n10235), .A(n10234), .B(n10233), .ZN(
        n10237) );
  AOI22_X1 U11305 ( .A1(n10353), .A2(n10238), .B1(n10237), .B2(n10350), .ZN(
        P2_U3220) );
  INV_X1 U11306 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10240) );
  AOI22_X1 U11307 ( .A1(n10375), .A2(n10240), .B1(n10239), .B2(n10372), .ZN(
        P2_U3429) );
  OAI22_X1 U11308 ( .A1(n10244), .A2(n10243), .B1(n10242), .B2(n10241), .ZN(
        n10246) );
  AOI211_X1 U11309 ( .C1(n10248), .C2(n10247), .A(n10246), .B(n10245), .ZN(
        n10249) );
  OAI21_X1 U11310 ( .B1(n10251), .B2(n10250), .A(n10249), .ZN(n10252) );
  AOI21_X1 U11311 ( .B1(n10253), .B2(n10302), .A(n10252), .ZN(n10256) );
  INV_X1 U11312 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10254) );
  AOI22_X1 U11313 ( .A1(n10316), .A2(n10256), .B1(n10254), .B2(n10313), .ZN(
        P1_U3537) );
  AOI22_X1 U11314 ( .A1(n10306), .A2(n10256), .B1(n10255), .B2(n10304), .ZN(
        P1_U3498) );
  XNOR2_X1 U11315 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11316 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U11317 ( .A(n10265), .ZN(n10264) );
  NOR2_X1 U11318 ( .A1(n10264), .A2(n10257), .ZN(P1_U3294) );
  AND2_X1 U11319 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10265), .ZN(P1_U3295) );
  AND2_X1 U11320 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10265), .ZN(P1_U3296) );
  NOR2_X1 U11321 ( .A1(n10264), .A2(n10258), .ZN(P1_U3297) );
  AND2_X1 U11322 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10265), .ZN(P1_U3298) );
  AND2_X1 U11323 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10265), .ZN(P1_U3299) );
  AND2_X1 U11324 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10265), .ZN(P1_U3300) );
  AND2_X1 U11325 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10265), .ZN(P1_U3301) );
  AND2_X1 U11326 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10265), .ZN(P1_U3302) );
  AND2_X1 U11327 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10265), .ZN(P1_U3303) );
  AND2_X1 U11328 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10265), .ZN(P1_U3304) );
  AND2_X1 U11329 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10265), .ZN(P1_U3305) );
  AND2_X1 U11330 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10265), .ZN(P1_U3306) );
  NOR2_X1 U11331 ( .A1(n10264), .A2(n10259), .ZN(P1_U3307) );
  AND2_X1 U11332 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10265), .ZN(P1_U3308) );
  AND2_X1 U11333 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10265), .ZN(P1_U3309) );
  AND2_X1 U11334 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10265), .ZN(P1_U3310) );
  AND2_X1 U11335 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10265), .ZN(P1_U3311) );
  NOR2_X1 U11336 ( .A1(n10264), .A2(n10260), .ZN(P1_U3312) );
  NOR2_X1 U11337 ( .A1(n10264), .A2(n10261), .ZN(P1_U3313) );
  AND2_X1 U11338 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10265), .ZN(P1_U3314) );
  AND2_X1 U11339 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10265), .ZN(P1_U3315) );
  AND2_X1 U11340 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10265), .ZN(P1_U3316) );
  NOR2_X1 U11341 ( .A1(n10264), .A2(n10262), .ZN(P1_U3317) );
  AND2_X1 U11342 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10265), .ZN(P1_U3318) );
  AND2_X1 U11343 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10265), .ZN(P1_U3319) );
  AND2_X1 U11344 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10265), .ZN(P1_U3320) );
  NOR2_X1 U11345 ( .A1(n10264), .A2(n10263), .ZN(P1_U3321) );
  AND2_X1 U11346 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10265), .ZN(P1_U3322) );
  AND2_X1 U11347 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10265), .ZN(P1_U3323) );
  INV_X1 U11348 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10266) );
  AOI22_X1 U11349 ( .A1(n10306), .A2(n10267), .B1(n10266), .B2(n10304), .ZN(
        P1_U3453) );
  OAI21_X1 U11350 ( .B1(n10269), .B2(n10299), .A(n10268), .ZN(n10271) );
  AOI211_X1 U11351 ( .C1(n10302), .C2(n10272), .A(n10271), .B(n10270), .ZN(
        n10307) );
  INV_X1 U11352 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10273) );
  AOI22_X1 U11353 ( .A1(n10306), .A2(n10307), .B1(n10273), .B2(n10304), .ZN(
        P1_U3459) );
  OAI21_X1 U11354 ( .B1(n10275), .B2(n10299), .A(n10274), .ZN(n10277) );
  AOI211_X1 U11355 ( .C1(n10302), .C2(n10278), .A(n10277), .B(n10276), .ZN(
        n10308) );
  INV_X1 U11356 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10279) );
  AOI22_X1 U11357 ( .A1(n10306), .A2(n10308), .B1(n10279), .B2(n10304), .ZN(
        P1_U3465) );
  NAND2_X1 U11358 ( .A1(n10280), .A2(n10302), .ZN(n10282) );
  OAI211_X1 U11359 ( .C1(n7183), .C2(n10299), .A(n10282), .B(n10281), .ZN(
        n10283) );
  NOR2_X1 U11360 ( .A1(n10284), .A2(n10283), .ZN(n10309) );
  INV_X1 U11361 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10285) );
  AOI22_X1 U11362 ( .A1(n10306), .A2(n10309), .B1(n10285), .B2(n10304), .ZN(
        P1_U3471) );
  OAI21_X1 U11363 ( .B1(n10287), .B2(n10299), .A(n10286), .ZN(n10289) );
  AOI211_X1 U11364 ( .C1(n10302), .C2(n10290), .A(n10289), .B(n10288), .ZN(
        n10310) );
  INV_X1 U11365 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10291) );
  AOI22_X1 U11366 ( .A1(n10306), .A2(n10310), .B1(n10291), .B2(n10304), .ZN(
        P1_U3483) );
  OAI21_X1 U11367 ( .B1(n10293), .B2(n10299), .A(n10292), .ZN(n10294) );
  AOI211_X1 U11368 ( .C1(n10296), .C2(n10302), .A(n10295), .B(n10294), .ZN(
        n10312) );
  INV_X1 U11369 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10297) );
  AOI22_X1 U11370 ( .A1(n10306), .A2(n10312), .B1(n10297), .B2(n10304), .ZN(
        P1_U3489) );
  OAI21_X1 U11371 ( .B1(n9476), .B2(n10299), .A(n10298), .ZN(n10300) );
  AOI211_X1 U11372 ( .C1(n10303), .C2(n10302), .A(n10301), .B(n10300), .ZN(
        n10315) );
  INV_X1 U11373 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10305) );
  AOI22_X1 U11374 ( .A1(n10306), .A2(n10315), .B1(n10305), .B2(n10304), .ZN(
        P1_U3495) );
  AOI22_X1 U11375 ( .A1(n10316), .A2(n10307), .B1(n6665), .B2(n10313), .ZN(
        P1_U3524) );
  AOI22_X1 U11376 ( .A1(n10316), .A2(n10308), .B1(n6672), .B2(n10313), .ZN(
        P1_U3526) );
  AOI22_X1 U11377 ( .A1(n10316), .A2(n10309), .B1(n6692), .B2(n10313), .ZN(
        P1_U3528) );
  AOI22_X1 U11378 ( .A1(n10316), .A2(n10310), .B1(n6917), .B2(n10313), .ZN(
        P1_U3532) );
  AOI22_X1 U11379 ( .A1(n10316), .A2(n10312), .B1(n10311), .B2(n10313), .ZN(
        P1_U3534) );
  AOI22_X1 U11380 ( .A1(n10316), .A2(n10315), .B1(n10314), .B2(n10313), .ZN(
        P1_U3536) );
  INV_X1 U11381 ( .A(n10317), .ZN(n10333) );
  INV_X1 U11382 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n10329) );
  OAI21_X1 U11383 ( .B1(n10320), .B2(n10319), .A(n10318), .ZN(n10326) );
  AOI211_X1 U11384 ( .C1(n10324), .C2(n10323), .A(n10322), .B(n10321), .ZN(
        n10325) );
  AOI21_X1 U11385 ( .B1(n10327), .B2(n10326), .A(n10325), .ZN(n10328) );
  OAI21_X1 U11386 ( .B1(n10330), .B2(n10329), .A(n10328), .ZN(n10331) );
  AOI21_X1 U11387 ( .B1(n10333), .B2(n10332), .A(n10331), .ZN(n10340) );
  OAI21_X1 U11388 ( .B1(n10336), .B2(n10335), .A(n10334), .ZN(n10337) );
  NAND2_X1 U11389 ( .A1(n10338), .A2(n10337), .ZN(n10339) );
  OAI211_X1 U11390 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10341), .A(n10340), .B(
        n10339), .ZN(P2_U3184) );
  INV_X1 U11391 ( .A(n10342), .ZN(n10349) );
  OAI22_X1 U11392 ( .A1(n10345), .A2(n10341), .B1(n10344), .B2(n10343), .ZN(
        n10347) );
  AOI211_X1 U11393 ( .C1(n10349), .C2(n10348), .A(n10347), .B(n10346), .ZN(
        n10351) );
  AOI22_X1 U11394 ( .A1(n10353), .A2(n10352), .B1(n10351), .B2(n10350), .ZN(
        P2_U3231) );
  AOI22_X1 U11395 ( .A1(n10375), .A2(n10355), .B1(n10354), .B2(n10372), .ZN(
        P2_U3396) );
  AOI22_X1 U11396 ( .A1(n10375), .A2(n10357), .B1(n10356), .B2(n10372), .ZN(
        P2_U3402) );
  INV_X1 U11397 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10359) );
  AOI22_X1 U11398 ( .A1(n10375), .A2(n10359), .B1(n10358), .B2(n10372), .ZN(
        P2_U3405) );
  INV_X1 U11399 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10361) );
  AOI22_X1 U11400 ( .A1(n10375), .A2(n10361), .B1(n10360), .B2(n10372), .ZN(
        P2_U3408) );
  INV_X1 U11401 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10363) );
  AOI22_X1 U11402 ( .A1(n10375), .A2(n10363), .B1(n10362), .B2(n10372), .ZN(
        P2_U3411) );
  INV_X1 U11403 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10365) );
  AOI22_X1 U11404 ( .A1(n10375), .A2(n10365), .B1(n10364), .B2(n10372), .ZN(
        P2_U3414) );
  INV_X1 U11405 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10367) );
  AOI22_X1 U11406 ( .A1(n10375), .A2(n10367), .B1(n10366), .B2(n10372), .ZN(
        P2_U3417) );
  AOI22_X1 U11407 ( .A1(n10375), .A2(n10369), .B1(n10368), .B2(n10372), .ZN(
        P2_U3420) );
  INV_X1 U11408 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10371) );
  AOI22_X1 U11409 ( .A1(n10375), .A2(n10371), .B1(n10370), .B2(n10372), .ZN(
        P2_U3423) );
  AOI22_X1 U11410 ( .A1(n10375), .A2(n10374), .B1(n10373), .B2(n10372), .ZN(
        P2_U3426) );
  NAND2_X1 U11411 ( .A1(n10377), .A2(n10376), .ZN(n10378) );
  XOR2_X1 U11412 ( .A(n10379), .B(n10378), .Z(ADD_1068_U5) );
  AOI22_X1 U11413 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .B1(n10380), .B2(n7255), .ZN(ADD_1068_U46) );
  NOR2_X1 U11414 ( .A1(n10382), .A2(n10381), .ZN(n10383) );
  XOR2_X1 U11415 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n10383), .Z(ADD_1068_U55)
         );
  XNOR2_X1 U11416 ( .A(n10385), .B(n10384), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11417 ( .A(n10387), .B(n10386), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11418 ( .A(n10389), .B(n10388), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11419 ( .A(n10391), .B(n10390), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11420 ( .A(n10393), .B(n10392), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11421 ( .A(n10395), .B(n10394), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11422 ( .A(n10397), .B(n10396), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11423 ( .A(n10399), .B(n10398), .ZN(ADD_1068_U63) );
  XNOR2_X1 U11424 ( .A(n10401), .B(n10400), .ZN(ADD_1068_U50) );
  XNOR2_X1 U11425 ( .A(n10403), .B(n10402), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11426 ( .A(n10405), .B(n10404), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11427 ( .A(n10407), .B(n10406), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11428 ( .A(n10409), .B(n10408), .ZN(ADD_1068_U48) );
  XOR2_X1 U11429 ( .A(n10411), .B(n10410), .Z(ADD_1068_U54) );
  XOR2_X1 U11430 ( .A(n10413), .B(n10412), .Z(ADD_1068_U53) );
  XNOR2_X1 U11431 ( .A(n10415), .B(n10414), .ZN(ADD_1068_U52) );
  AND2_X1 U4920 ( .A1(n4877), .A2(n4430), .ZN(n8447) );
  NAND2_X1 U4934 ( .A1(n7439), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7547) );
  OR2_X1 U4948 ( .A1(n8536), .A2(n8535), .ZN(n4894) );
  CLKBUF_X2 U4950 ( .A(n5139), .Z(n5734) );
  NOR2_X2 U4964 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5080) );
  INV_X1 U4965 ( .A(n5998), .ZN(n6115) );
  XNOR2_X1 U4967 ( .A(n8579), .B(n8597), .ZN(n8560) );
  AOI211_X1 U5890 ( .C1(n10332), .C2(n8597), .A(n8576), .B(n8575), .ZN(n8577)
         );
  CLKBUF_X2 U6165 ( .A(n6603), .Z(n4408) );
endmodule

