

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput127, keyinput126, keyinput125, keyinput124, keyinput123, 
        keyinput122, keyinput121, keyinput120, keyinput119, keyinput118, 
        keyinput117, keyinput116, keyinput115, keyinput114, keyinput113, 
        keyinput112, keyinput111, keyinput110, keyinput109, keyinput108, 
        keyinput107, keyinput106, keyinput105, keyinput104, keyinput103, 
        keyinput102, keyinput101, keyinput100, keyinput99, keyinput98, 
        keyinput97, keyinput96, keyinput95, keyinput94, keyinput93, keyinput92, 
        keyinput91, keyinput90, keyinput89, keyinput88, keyinput87, keyinput86, 
        keyinput85, keyinput84, keyinput83, keyinput82, keyinput81, keyinput80, 
        keyinput79, keyinput78, keyinput77, keyinput76, keyinput75, keyinput74, 
        keyinput73, keyinput72, keyinput71, keyinput70, keyinput69, keyinput68, 
        keyinput67, keyinput66, keyinput65, keyinput64, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855;

  INV_X2 U2370 ( .A(n3416), .ZN(n3373) );
  INV_X2 U2371 ( .A(n2649), .ZN(n3416) );
  NAND2_X1 U2372 ( .A1(n3703), .A2(n3767), .ZN(n2652) );
  NAND4_X2 U2373 ( .A1(n2795), .A2(n2792), .A3(n2790), .A4(n2791), .ZN(n2800)
         );
  CLKBUF_X2 U2374 ( .A(n2537), .Z(n3634) );
  XNOR2_X1 U2375 ( .A(n2332), .B(n2331), .ZN(n2334) );
  INV_X1 U2376 ( .A(n3448), .ZN(n3417) );
  INV_X1 U2377 ( .A(n3445), .ZN(n3422) );
  OAI21_X1 U2378 ( .B1(n3148), .B2(n2237), .A(n3149), .ZN(n3188) );
  CLKBUF_X3 U2379 ( .A(n2538), .Z(n3297) );
  AND4_X1 U2380 ( .A1(n2381), .A2(n2380), .A3(n2379), .A4(n2378), .ZN(n2764)
         );
  AOI21_X2 U2381 ( .B1(n4165), .B2(n3859), .A(n3858), .ZN(n4145) );
  XNOR2_X2 U2382 ( .A(n2329), .B(IR_REG_30__SCAN_IN), .ZN(n2434) );
  NAND2_X2 U2383 ( .A1(n2288), .A2(IR_REG_31__SCAN_IN), .ZN(n2329) );
  AND2_X1 U2384 ( .A1(n2667), .A2(n3767), .ZN(n4536) );
  XNOR2_X2 U2385 ( .A(n2371), .B(n2370), .ZN(n3767) );
  AND2_X1 U2386 ( .A1(n4145), .A2(n3860), .ZN(n4103) );
  AND2_X2 U2387 ( .A1(n2413), .A2(n4196), .ZN(n4477) );
  NAND2_X1 U2388 ( .A1(n2576), .A2(n2575), .ZN(n2649) );
  INV_X1 U2389 ( .A(n2577), .ZN(n2668) );
  INV_X2 U2390 ( .A(n3434), .ZN(n3446) );
  INV_X1 U2391 ( .A(n2760), .ZN(n2655) );
  NAND2_X2 U2392 ( .A1(n2576), .A2(n2652), .ZN(n3448) );
  INV_X2 U2393 ( .A(n3783), .ZN(U4043) );
  AND2_X1 U2394 ( .A1(n2336), .A2(n4344), .ZN(n2538) );
  NAND2_X1 U2395 ( .A1(n2342), .A2(IR_REG_31__SCAN_IN), .ZN(n2467) );
  AND2_X2 U2396 ( .A1(n2422), .A2(n2312), .ZN(n3327) );
  AND2_X1 U2397 ( .A1(n3328), .A2(n2314), .ZN(n2315) );
  NOR2_X1 U2398 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2302)
         );
  CLKBUF_X1 U2399 ( .A(IR_REG_0__SCAN_IN), .Z(n4357) );
  NOR2_X2 U2400 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2349)
         );
  NOR2_X1 U2401 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n4804)
         );
  NOR2_X2 U2402 ( .A1(n2868), .A2(n2887), .ZN(n2894) );
  NAND2_X1 U2403 ( .A1(n3295), .A2(n2216), .ZN(n2215) );
  NAND2_X1 U2404 ( .A1(n2336), .A2(n2334), .ZN(n2537) );
  AND2_X1 U2405 ( .A1(n2129), .A2(n2153), .ZN(n2197) );
  INV_X1 U2406 ( .A(IR_REG_25__SCAN_IN), .ZN(n2198) );
  OR2_X1 U2407 ( .A1(n4382), .A2(n2173), .ZN(n2240) );
  INV_X1 U2408 ( .A(n3897), .ZN(n2297) );
  NAND2_X1 U2409 ( .A1(n4129), .A2(n4116), .ZN(n2298) );
  AND2_X1 U2410 ( .A1(n2791), .A2(n2790), .ZN(n2794) );
  INV_X1 U2411 ( .A(n3248), .ZN(n2276) );
  INV_X1 U2412 ( .A(IR_REG_21__SCAN_IN), .ZN(n2300) );
  INV_X1 U2413 ( .A(IR_REG_11__SCAN_IN), .ZN(n3152) );
  INV_X1 U2414 ( .A(n3561), .ZN(n2223) );
  INV_X1 U2415 ( .A(n2139), .ZN(n2214) );
  AOI21_X1 U2416 ( .B1(n3291), .B2(n3290), .A(n3289), .ZN(n3296) );
  INV_X1 U2417 ( .A(n3288), .ZN(n3289) );
  AND2_X1 U2418 ( .A1(n3287), .A2(n3286), .ZN(n3291) );
  AOI21_X1 U2419 ( .B1(n2139), .B2(n2213), .A(n2164), .ZN(n2212) );
  NOR2_X1 U2420 ( .A1(n3295), .A2(n2216), .ZN(n2213) );
  NAND2_X1 U2421 ( .A1(n2369), .A2(IR_REG_31__SCAN_IN), .ZN(n2374) );
  INV_X1 U2422 ( .A(IR_REG_19__SCAN_IN), .ZN(n2373) );
  NAND2_X1 U2423 ( .A1(n2374), .A2(n2373), .ZN(n2372) );
  INV_X1 U2424 ( .A(n3439), .ZN(n3459) );
  AND2_X1 U2425 ( .A1(n3444), .A2(n3443), .ZN(n3946) );
  AOI21_X1 U2426 ( .B1(n4144), .B2(n3894), .A(n2156), .ZN(n4123) );
  NAND2_X1 U2427 ( .A1(n2283), .A2(n2282), .ZN(n3227) );
  AOI21_X1 U2428 ( .B1(n2284), .B2(n3139), .A(n2163), .ZN(n2282) );
  OR2_X1 U2429 ( .A1(n2861), .A2(n2860), .ZN(n2863) );
  NAND2_X1 U2430 ( .A1(n2330), .A2(IR_REG_31__SCAN_IN), .ZN(n2332) );
  NOR2_X1 U2431 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2316)
         );
  AND4_X1 U2432 ( .A1(n4804), .A2(n2311), .A3(n2310), .A4(n2309), .ZN(n2312)
         );
  NOR2_X1 U2433 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2311)
         );
  NOR2_X1 U2434 ( .A1(IR_REG_13__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2310)
         );
  OAI21_X1 U2435 ( .B1(n2374), .B2(n2373), .A(n2372), .ZN(n3849) );
  NOR2_X1 U2436 ( .A1(n4469), .A2(n4470), .ZN(n4468) );
  NAND2_X1 U2437 ( .A1(n4452), .A2(n2180), .ZN(n4469) );
  NAND2_X1 U2438 ( .A1(n4490), .A2(n2181), .ZN(n2180) );
  AOI21_X1 U2439 ( .B1(n4462), .B2(n4461), .A(n4460), .ZN(n4467) );
  NOR2_X1 U2440 ( .A1(n3058), .A2(n3067), .ZN(n3064) );
  INV_X1 U2441 ( .A(n3057), .ZN(n3058) );
  INV_X1 U2442 ( .A(n3559), .ZN(n2228) );
  AOI21_X1 U2443 ( .B1(n3798), .B2(n3800), .A(n2238), .ZN(n2544) );
  AND2_X1 U2444 ( .A1(n2723), .A2(REG1_REG_2__SCAN_IN), .ZN(n2238) );
  NAND2_X1 U2445 ( .A1(n2262), .A2(n2556), .ZN(n2557) );
  NAND2_X1 U2446 ( .A1(n2554), .A2(REG2_REG_3__SCAN_IN), .ZN(n2262) );
  AOI21_X1 U2447 ( .B1(n2559), .B2(REG2_REG_5__SCAN_IN), .A(n2623), .ZN(n2609)
         );
  NAND2_X1 U2448 ( .A1(n2699), .A2(n2304), .ZN(n2701) );
  OR2_X1 U2449 ( .A1(n4402), .A2(n3814), .ZN(n3815) );
  AOI21_X1 U2450 ( .B1(n4409), .B2(n3835), .A(n2257), .ZN(n3837) );
  AND2_X1 U2451 ( .A1(n4407), .A2(REG2_REG_13__SCAN_IN), .ZN(n2257) );
  INV_X1 U2452 ( .A(n3900), .ZN(n2291) );
  NAND2_X1 U2453 ( .A1(n2764), .A2(n2938), .ZN(n3706) );
  OR2_X1 U2454 ( .A1(n2467), .A2(n2343), .ZN(n2345) );
  AND2_X1 U2455 ( .A1(n3774), .A2(n3703), .ZN(n2442) );
  NAND2_X1 U2456 ( .A1(n3905), .A2(n3990), .ZN(n2202) );
  NAND2_X1 U2457 ( .A1(n3265), .A2(n3249), .ZN(n3253) );
  INV_X1 U2458 ( .A(IR_REG_28__SCAN_IN), .ZN(n4798) );
  AND2_X1 U2459 ( .A1(n2194), .A2(n2313), .ZN(n3328) );
  INV_X1 U2460 ( .A(IR_REG_17__SCAN_IN), .ZN(n2313) );
  INV_X1 U2461 ( .A(IR_REG_14__SCAN_IN), .ZN(n4797) );
  AND2_X1 U2462 ( .A1(n2653), .A2(n2652), .ZN(n3434) );
  NOR2_X1 U2463 ( .A1(n2231), .A2(n2167), .ZN(n2230) );
  INV_X1 U2464 ( .A(n3401), .ZN(n2231) );
  OAI21_X1 U2465 ( .B1(n3445), .B2(n2663), .A(n2582), .ZN(n2583) );
  AND2_X1 U2466 ( .A1(n3354), .A2(n3353), .ZN(n3561) );
  AND2_X1 U2467 ( .A1(n3348), .A2(n3347), .ZN(n2227) );
  OR2_X1 U2468 ( .A1(n2226), .A2(n2157), .ZN(n2224) );
  INV_X1 U2469 ( .A(n3488), .ZN(n2226) );
  NAND2_X1 U2470 ( .A1(n2228), .A2(n2227), .ZN(n2225) );
  NAND2_X1 U2471 ( .A1(n2222), .A2(n2218), .ZN(n3568) );
  NAND2_X1 U2472 ( .A1(n2220), .A2(n2219), .ZN(n2218) );
  NAND2_X1 U2473 ( .A1(n3488), .A2(n2217), .ZN(n2222) );
  INV_X1 U2474 ( .A(n2305), .ZN(n2219) );
  XNOR2_X1 U2475 ( .A(n2724), .B(n3446), .ZN(n2742) );
  OAI22_X1 U2476 ( .A1(n2764), .A2(n2649), .B1(n2761), .B2(n3448), .ZN(n2724)
         );
  NAND2_X1 U2477 ( .A1(n2210), .A2(n2209), .ZN(n3599) );
  AOI21_X1 U2478 ( .B1(n2140), .B2(n2214), .A(n2168), .ZN(n2209) );
  AND2_X1 U2479 ( .A1(n4348), .A2(n4349), .ZN(n2324) );
  OAI21_X1 U2480 ( .B1(n2191), .B2(n2612), .A(n2188), .ZN(n2687) );
  NAND2_X1 U2481 ( .A1(n2611), .A2(n2189), .ZN(n2188) );
  NOR2_X1 U2482 ( .A1(n2612), .A2(n2190), .ZN(n2189) );
  XNOR2_X1 U2483 ( .A(n2609), .B(n4353), .ZN(n2611) );
  AOI21_X1 U2484 ( .B1(n2559), .B2(REG1_REG_5__SCAN_IN), .A(n2629), .ZN(n2603)
         );
  INV_X1 U2485 ( .A(IR_REG_9__SCAN_IN), .ZN(n2684) );
  OR2_X1 U2486 ( .A1(n2687), .A2(n2264), .ZN(n2263) );
  AND2_X1 U2487 ( .A1(n4352), .A2(REG2_REG_7__SCAN_IN), .ZN(n2264) );
  NAND2_X1 U2488 ( .A1(n2701), .A2(n2254), .ZN(n2256) );
  AND2_X1 U2489 ( .A1(n2700), .A2(n2255), .ZN(n2254) );
  INV_X1 U2490 ( .A(n4499), .ZN(n2255) );
  XNOR2_X1 U2491 ( .A(n2240), .B(n3832), .ZN(n4394) );
  NOR2_X1 U2492 ( .A1(n4394), .A2(n4395), .ZN(n4393) );
  OR2_X1 U2493 ( .A1(n4430), .A2(n4431), .ZN(n2186) );
  XNOR2_X1 U2494 ( .A(n2131), .B(n3311), .ZN(n4443) );
  NAND2_X1 U2495 ( .A1(n4443), .A2(n4442), .ZN(n4441) );
  OR2_X1 U2496 ( .A1(n3437), .A2(n3436), .ZN(n3853) );
  NOR2_X2 U2497 ( .A1(n3936), .A2(n3923), .ZN(n4211) );
  OR2_X1 U2498 ( .A1(n3427), .A2(n4777), .ZN(n3437) );
  INV_X1 U2499 ( .A(n3913), .ZN(n3954) );
  NAND2_X1 U2500 ( .A1(n2133), .A2(n2161), .ZN(n2280) );
  NAND2_X1 U2501 ( .A1(n2296), .A2(n2298), .ZN(n2293) );
  OR2_X1 U2502 ( .A1(n2295), .A2(n2297), .ZN(n2294) );
  INV_X1 U2503 ( .A(n2298), .ZN(n2295) );
  NAND2_X1 U2504 ( .A1(n4123), .A2(n4125), .ZN(n4122) );
  NAND2_X1 U2505 ( .A1(n4188), .A2(n4172), .ZN(n3893) );
  INV_X1 U2506 ( .A(n4155), .ZN(n4148) );
  NOR2_X1 U2507 ( .A1(n3237), .A2(n3228), .ZN(n3230) );
  NOR2_X1 U2508 ( .A1(n3690), .A2(n2285), .ZN(n2284) );
  INV_X1 U2509 ( .A(n2286), .ZN(n2285) );
  OR2_X1 U2510 ( .A1(n3138), .A2(n3137), .ZN(n2286) );
  NOR2_X1 U2511 ( .A1(n3087), .A2(n3091), .ZN(n2306) );
  NOR2_X1 U2512 ( .A1(n2902), .A2(n2445), .ZN(n2904) );
  NAND2_X1 U2513 ( .A1(n2833), .A2(REG3_REG_6__SCAN_IN), .ZN(n2902) );
  AND2_X1 U2514 ( .A1(n2856), .A2(n2855), .ZN(n2857) );
  INV_X1 U2515 ( .A(n3703), .ZN(n3696) );
  AND2_X1 U2516 ( .A1(n3349), .A2(DATAI_30_), .ZN(n4217) );
  NOR2_X1 U2517 ( .A1(n4090), .A2(n4062), .ZN(n4067) );
  INV_X1 U2518 ( .A(n4349), .ZN(n2409) );
  INV_X1 U2519 ( .A(IR_REG_24__SCAN_IN), .ZN(n2318) );
  INV_X1 U2520 ( .A(IR_REG_23__SCAN_IN), .ZN(n2325) );
  AND2_X1 U2521 ( .A1(n2316), .A2(n2300), .ZN(n2299) );
  INV_X1 U2522 ( .A(IR_REG_16__SCAN_IN), .ZN(n3309) );
  AND2_X1 U2523 ( .A1(n3105), .A2(n3109), .ZN(n3830) );
  AND2_X1 U2524 ( .A1(n2308), .A2(n2269), .ZN(n2268) );
  INV_X1 U2525 ( .A(IR_REG_5__SCAN_IN), .ZN(n2269) );
  NAND2_X1 U2526 ( .A1(IR_REG_31__SCAN_IN), .A2(n2418), .ZN(n2548) );
  INV_X1 U2527 ( .A(n3136), .ZN(n3137) );
  AND4_X1 U2528 ( .A1(n2542), .A2(n2541), .A3(n2540), .A4(n2539), .ZN(n2865)
         );
  OR2_X1 U2529 ( .A1(n2537), .A2(n4826), .ZN(n2541) );
  INV_X1 U2530 ( .A(n4023), .ZN(n3987) );
  NAND2_X1 U2531 ( .A1(n2832), .A2(n2831), .ZN(n2946) );
  NAND2_X1 U2532 ( .A1(n2538), .A2(REG1_REG_1__SCAN_IN), .ZN(n2337) );
  OR2_X1 U2533 ( .A1(n2537), .A2(n2335), .ZN(n2338) );
  OR2_X1 U2534 ( .A1(n2662), .A2(n2661), .ZN(n3623) );
  OR2_X1 U2535 ( .A1(n2662), .A2(n2596), .ZN(n3626) );
  NAND4_X1 U2536 ( .A1(n2465), .A2(n2464), .A3(n2463), .A4(n2462), .ZN(n3585)
         );
  OR2_X1 U2537 ( .A1(n2536), .A2(n2718), .ZN(n2357) );
  AND3_X1 U2538 ( .A1(n2356), .A2(n2355), .A3(n2354), .ZN(n2358) );
  XNOR2_X1 U2539 ( .A(n2263), .B(n4499), .ZN(n4370) );
  NAND2_X1 U2540 ( .A1(n4370), .A2(REG2_REG_8__SCAN_IN), .ZN(n2179) );
  NAND2_X1 U2541 ( .A1(n4378), .A2(n3828), .ZN(n4388) );
  NAND2_X1 U2542 ( .A1(n4388), .A2(n4389), .ZN(n4387) );
  OAI21_X1 U2543 ( .B1(n4387), .B2(n3832), .A(n2182), .ZN(n4399) );
  AOI21_X1 U2544 ( .B1(n4387), .B2(n2184), .A(n2183), .ZN(n2182) );
  NOR2_X1 U2545 ( .A1(n4495), .A2(n2185), .ZN(n2184) );
  NOR2_X1 U2546 ( .A1(n3832), .A2(n3831), .ZN(n2183) );
  NAND2_X1 U2547 ( .A1(n4399), .A2(REG2_REG_12__SCAN_IN), .ZN(n4398) );
  NAND2_X1 U2548 ( .A1(n4453), .A2(n4454), .ZN(n4452) );
  AOI21_X1 U2549 ( .B1(n3844), .B2(REG2_REG_18__SCAN_IN), .A(n4468), .ZN(n3846) );
  AND2_X1 U2550 ( .A1(n2479), .A2(n3772), .ZN(n4472) );
  NAND2_X1 U2551 ( .A1(n4449), .A2(n2303), .ZN(n4462) );
  NAND2_X1 U2552 ( .A1(n3885), .A2(n3884), .ZN(n4222) );
  NAND2_X1 U2553 ( .A1(n3880), .A2(n4184), .ZN(n3885) );
  AND2_X1 U2554 ( .A1(n4104), .A2(n3641), .ZN(n3861) );
  OAI21_X1 U2555 ( .B1(n2731), .B2(n2207), .A(n2773), .ZN(n2205) );
  NOR2_X1 U2556 ( .A1(n2157), .A2(n2305), .ZN(n2217) );
  NAND2_X1 U2557 ( .A1(n2225), .A2(n2221), .ZN(n2220) );
  NOR2_X1 U2558 ( .A1(n3561), .A2(n2160), .ZN(n2221) );
  INV_X1 U2559 ( .A(n4426), .ZN(n2252) );
  OR2_X1 U2560 ( .A1(n4425), .A2(n3818), .ZN(n3820) );
  AND2_X1 U2561 ( .A1(n3946), .A2(n3937), .ZN(n3876) );
  AND2_X1 U2562 ( .A1(n3349), .A2(DATAI_27_), .ZN(n3913) );
  OR2_X1 U2563 ( .A1(n2280), .A2(n2279), .ZN(n2278) );
  NAND2_X1 U2564 ( .A1(n3780), .A2(n2990), .ZN(n3722) );
  AND2_X1 U2565 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2516) );
  AND3_X1 U2566 ( .A1(n4797), .A2(n3309), .A3(n3306), .ZN(n2194) );
  NOR2_X1 U2567 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2309)
         );
  INV_X1 U2568 ( .A(IR_REG_6__SCAN_IN), .ZN(n2606) );
  NAND2_X1 U2569 ( .A1(n3189), .A2(n2308), .ZN(n2266) );
  AND2_X1 U2570 ( .A1(n3481), .A2(n3482), .ZN(n3401) );
  OR2_X1 U2571 ( .A1(n3367), .A2(n3571), .ZN(n3378) );
  NAND2_X1 U2572 ( .A1(n3064), .A2(n3063), .ZN(n3100) );
  INV_X1 U2573 ( .A(n3062), .ZN(n3063) );
  NAND2_X1 U2574 ( .A1(n3061), .A2(n3060), .ZN(n3103) );
  NAND2_X1 U2575 ( .A1(n3632), .A2(REG2_REG_4__SCAN_IN), .ZN(n2539) );
  XNOR2_X1 U2576 ( .A(n2741), .B(n3446), .ZN(n2775) );
  NAND2_X1 U2577 ( .A1(n3355), .A2(REG3_REG_21__SCAN_IN), .ZN(n3367) );
  NOR2_X1 U2578 ( .A1(n2525), .A2(n4775), .ZN(n2526) );
  NAND2_X1 U2579 ( .A1(n2232), .A2(n3402), .ZN(n3535) );
  OR2_X1 U2580 ( .A1(n3479), .A2(n3403), .ZN(n2232) );
  INV_X1 U2581 ( .A(n2172), .ZN(n2237) );
  NAND2_X1 U2582 ( .A1(n3349), .A2(DATAI_22_), .ZN(n4052) );
  OAI22_X1 U2583 ( .A1(n2651), .A2(n3445), .B1(n2649), .B2(n2655), .ZN(n2726)
         );
  OAI21_X1 U2584 ( .B1(n2651), .B2(n2649), .A(n2650), .ZN(n2654) );
  NAND2_X1 U2585 ( .A1(n2760), .A2(n3417), .ZN(n2650) );
  INV_X1 U2586 ( .A(n2730), .ZN(n2208) );
  NAND2_X1 U2587 ( .A1(n2946), .A2(n2945), .ZN(n2982) );
  INV_X1 U2588 ( .A(n2950), .ZN(n2956) );
  AND3_X1 U2589 ( .A1(n3637), .A2(n3636), .A3(n3635), .ZN(n3679) );
  AND4_X1 U2590 ( .A1(n2501), .A2(n2500), .A3(n2499), .A4(n2498), .ZN(n4168)
         );
  OR2_X1 U2591 ( .A1(n2536), .A2(REG3_REG_3__SCAN_IN), .ZN(n2791) );
  OR2_X1 U2592 ( .A1(n3634), .A2(n2566), .ZN(n2795) );
  XNOR2_X1 U2593 ( .A(n2723), .B(n2476), .ZN(n3800) );
  NAND2_X1 U2594 ( .A1(n3802), .A2(n2485), .ZN(n2555) );
  XNOR2_X1 U2595 ( .A(n2557), .B(n2261), .ZN(n2558) );
  OR3_X1 U2596 ( .A1(n2681), .A2(IR_REG_7__SCAN_IN), .A3(IR_REG_8__SCAN_IN), 
        .ZN(n2683) );
  NAND2_X1 U2597 ( .A1(n3824), .A2(n2193), .ZN(n3827) );
  NAND2_X1 U2598 ( .A1(n4351), .A2(REG2_REG_9__SCAN_IN), .ZN(n2193) );
  NOR2_X1 U2599 ( .A1(n3809), .A2(n2301), .ZN(n3810) );
  INV_X1 U2600 ( .A(REG3_REG_11__SCAN_IN), .ZN(n4775) );
  NOR2_X1 U2601 ( .A1(n3813), .A2(n4393), .ZN(n4404) );
  INV_X1 U2602 ( .A(n2240), .ZN(n3812) );
  NAND2_X1 U2603 ( .A1(n2253), .A2(n3836), .ZN(n2250) );
  NAND2_X1 U2604 ( .A1(n3815), .A2(n4421), .ZN(n3816) );
  NAND2_X1 U2605 ( .A1(n3838), .A2(REG2_REG_14__SCAN_IN), .ZN(n2259) );
  NOR2_X1 U2606 ( .A1(n3837), .A2(n3836), .ZN(n3839) );
  XNOR2_X1 U2607 ( .A(n3820), .B(n4491), .ZN(n4440) );
  NAND2_X1 U2608 ( .A1(n4440), .A2(n4439), .ZN(n4438) );
  AND2_X1 U2609 ( .A1(n3349), .A2(n2443), .ZN(n2471) );
  AND2_X1 U2610 ( .A1(n2142), .A2(n2174), .ZN(n2247) );
  AOI21_X1 U2611 ( .B1(n4461), .B2(n2247), .A(n2246), .ZN(n2245) );
  NOR2_X1 U2612 ( .A1(n2142), .A2(n2174), .ZN(n2246) );
  AND2_X1 U2613 ( .A1(n3349), .A2(DATAI_29_), .ZN(n3923) );
  AND2_X1 U2614 ( .A1(n3433), .A2(n3432), .ZN(n3935) );
  INV_X1 U2615 ( .A(n3909), .ZN(n3910) );
  AOI21_X1 U2616 ( .B1(n2134), .B2(n2294), .A(n2158), .ZN(n2289) );
  AND2_X1 U2617 ( .A1(n3349), .A2(DATAI_21_), .ZN(n4062) );
  AND2_X1 U2618 ( .A1(n3668), .A2(n4017), .ZN(n4060) );
  AND2_X1 U2619 ( .A1(n3338), .A2(REG3_REG_20__SCAN_IN), .ZN(n3355) );
  OR2_X1 U2620 ( .A1(n3321), .A2(n4773), .ZN(n3337) );
  NOR2_X1 U2621 ( .A1(n3299), .A2(n3298), .ZN(n3300) );
  OR2_X1 U2622 ( .A1(n3165), .A2(n4770), .ZN(n3299) );
  AOI21_X1 U2623 ( .B1(n2273), .B2(n2272), .A(n2165), .ZN(n2271) );
  INV_X1 U2624 ( .A(n3253), .ZN(n2272) );
  INV_X1 U2625 ( .A(REG3_REG_14__SCAN_IN), .ZN(n3162) );
  INV_X1 U2626 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2459) );
  OR2_X1 U2627 ( .A1(n3716), .A2(n3009), .ZN(n3087) );
  AND2_X1 U2628 ( .A1(n2964), .A2(n3722), .ZN(n3716) );
  AND4_X1 U2629 ( .A1(n2909), .A2(n2908), .A3(n2907), .A4(n2906), .ZN(n3018)
         );
  INV_X1 U2630 ( .A(n4128), .ZN(n4187) );
  NAND2_X1 U2631 ( .A1(n2818), .A2(n2819), .ZN(n2868) );
  NAND2_X1 U2632 ( .A1(n2811), .A2(n3711), .ZN(n2861) );
  AND2_X1 U2633 ( .A1(n2803), .A2(n2806), .ZN(n2852) );
  OR2_X1 U2634 ( .A1(n2801), .A2(n2805), .ZN(n2856) );
  OR2_X1 U2635 ( .A1(n2923), .A2(n2849), .ZN(n2921) );
  INV_X1 U2636 ( .A(n2799), .ZN(n2793) );
  OR2_X1 U2637 ( .A1(n2635), .A2(n2587), .ZN(n4191) );
  NAND2_X1 U2638 ( .A1(n2345), .A2(n2344), .ZN(n2347) );
  NAND2_X1 U2639 ( .A1(n3973), .A2(n3954), .ZN(n2201) );
  NOR2_X1 U2640 ( .A1(n2144), .A2(n3937), .ZN(n3922) );
  NOR3_X1 U2641 ( .A1(n4028), .A2(n2202), .A3(n3677), .ZN(n3971) );
  NOR2_X1 U2642 ( .A1(n4028), .A2(n2202), .ZN(n3988) );
  OR2_X1 U2643 ( .A1(n4027), .A2(n3921), .ZN(n4028) );
  NAND2_X1 U2644 ( .A1(n3349), .A2(DATAI_23_), .ZN(n4029) );
  NAND2_X1 U2645 ( .A1(n4153), .A2(n2171), .ZN(n4090) );
  NAND2_X1 U2646 ( .A1(n4153), .A2(n2141), .ZN(n4115) );
  AND2_X1 U2647 ( .A1(n4153), .A2(n3896), .ZN(n4135) );
  NOR2_X1 U2648 ( .A1(n4270), .A2(n4148), .ZN(n4153) );
  NOR2_X1 U2649 ( .A1(n3269), .A2(n3887), .ZN(n4194) );
  AND2_X1 U2650 ( .A1(n2275), .A2(n3251), .ZN(n3254) );
  NAND2_X1 U2651 ( .A1(n2276), .A2(n3253), .ZN(n2275) );
  NAND2_X1 U2652 ( .A1(n2195), .A2(n3249), .ZN(n3269) );
  INV_X1 U2653 ( .A(n3203), .ZN(n2196) );
  INV_X1 U2654 ( .A(n3587), .ZN(n3207) );
  AND2_X1 U2655 ( .A1(n3080), .A2(n3137), .ZN(n3204) );
  NAND2_X1 U2656 ( .A1(n2894), .A2(n2135), .ZN(n2973) );
  NAND2_X1 U2657 ( .A1(n2177), .A2(n2894), .ZN(n3001) );
  INV_X1 U2658 ( .A(IR_REG_4__SCAN_IN), .ZN(n4799) );
  NOR2_X1 U2659 ( .A1(n2937), .A2(n2938), .ZN(n2936) );
  NAND2_X1 U2660 ( .A1(n2655), .A2(n2668), .ZN(n2937) );
  XNOR2_X1 U2661 ( .A(n2236), .B(n2317), .ZN(n2411) );
  NAND2_X1 U2662 ( .A1(n2148), .A2(IR_REG_31__SCAN_IN), .ZN(n2236) );
  INV_X1 U2663 ( .A(IR_REG_20__SCAN_IN), .ZN(n2370) );
  INV_X1 U2664 ( .A(IR_REG_15__SCAN_IN), .ZN(n3306) );
  AND2_X1 U2665 ( .A1(n3157), .A2(n3156), .ZN(n4407) );
  AND2_X1 U2666 ( .A1(n2239), .A2(n2418), .ZN(n2723) );
  INV_X1 U2667 ( .A(n2265), .ZN(n2239) );
  OAI21_X1 U2668 ( .B1(n2349), .B2(n2267), .A(n2266), .ZN(n2265) );
  NAND2_X1 U2669 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_2__SCAN_IN), .ZN(n2267)
         );
  MUX2_X1 U2670 ( .A(IR_REG_31__SCAN_IN), .B(n2348), .S(IR_REG_1__SCAN_IN), 
        .Z(n2351) );
  AOI21_X1 U2671 ( .B1(n3606), .B2(n3608), .A(n3607), .ZN(n3473) );
  AND4_X1 U2672 ( .A1(n3123), .A2(n3122), .A3(n3121), .A4(n3120), .ZN(n3265)
         );
  XNOR2_X1 U2673 ( .A(n2776), .B(n2775), .ZN(n2773) );
  AND2_X1 U2674 ( .A1(n3853), .A2(n3438), .ZN(n3938) );
  AND2_X1 U2675 ( .A1(n2224), .A2(n2169), .ZN(n3498) );
  AND4_X1 U2676 ( .A1(n2531), .A2(n2530), .A3(n2529), .A4(n2528), .ZN(n3141)
         );
  AOI21_X1 U2677 ( .B1(n3398), .B2(n3400), .A(n2234), .ZN(n2233) );
  AND2_X1 U2678 ( .A1(n3403), .A2(n3402), .ZN(n2234) );
  NAND2_X1 U2679 ( .A1(n2828), .A2(n2827), .ZN(n2832) );
  OR2_X1 U2680 ( .A1(n3296), .A2(n2214), .ZN(n2211) );
  AND4_X1 U2681 ( .A1(n2523), .A2(n2522), .A3(n2521), .A4(n2520), .ZN(n2955)
         );
  AOI21_X1 U2682 ( .B1(n3488), .B2(n3489), .A(n2227), .ZN(n3558) );
  AND4_X1 U2683 ( .A1(n3169), .A2(n3168), .A3(n3167), .A4(n3166), .ZN(n4192)
         );
  INV_X1 U2684 ( .A(n4052), .ZN(n4045) );
  INV_X1 U2685 ( .A(n3626), .ZN(n3583) );
  AND4_X1 U2686 ( .A1(n2882), .A2(n2881), .A3(n2880), .A4(n2879), .ZN(n3028)
         );
  AND2_X1 U2687 ( .A1(n2593), .A2(n4196), .ZN(n3624) );
  OR2_X1 U2688 ( .A1(n2662), .A2(n2590), .ZN(n3616) );
  INV_X1 U2689 ( .A(n3616), .ZN(n3621) );
  INV_X1 U2690 ( .A(n3614), .ZN(n3631) );
  NOR2_X1 U2691 ( .A1(n2649), .A2(n2595), .ZN(n3771) );
  INV_X1 U2692 ( .A(n3946), .ZN(n3916) );
  OAI211_X1 U2693 ( .C1(n3510), .C2(n3459), .A(n2621), .B(n2620), .ZN(n4005)
         );
  NAND2_X1 U2694 ( .A1(n2573), .A2(n2572), .ZN(n4023) );
  OAI211_X1 U2695 ( .C1(n4031), .C2(n3459), .A(n3382), .B(n3381), .ZN(n4044)
         );
  INV_X1 U2696 ( .A(n4130), .ZN(n4166) );
  INV_X1 U2697 ( .A(n4168), .ZN(n3890) );
  INV_X1 U2698 ( .A(n3265), .ZN(n3778) );
  INV_X1 U2699 ( .A(n3237), .ZN(n3584) );
  NAND4_X1 U2700 ( .A1(n2451), .A2(n2450), .A3(n2449), .A4(n2448), .ZN(n3088)
         );
  INV_X1 U2701 ( .A(n3018), .ZN(n3779) );
  INV_X1 U2702 ( .A(n3028), .ZN(n3780) );
  INV_X1 U2703 ( .A(n2651), .ZN(n2926) );
  AND2_X1 U2704 ( .A1(n2471), .A2(n2470), .ZN(n2479) );
  NAND2_X1 U2705 ( .A1(n2483), .A2(n2482), .ZN(n3785) );
  OR2_X1 U2706 ( .A1(n2481), .A2(REG2_REG_1__SCAN_IN), .ZN(n2483) );
  NAND2_X1 U2707 ( .A1(n2481), .A2(REG2_REG_1__SCAN_IN), .ZN(n2482) );
  NAND2_X1 U2708 ( .A1(n3803), .A2(n3804), .ZN(n3802) );
  OAI21_X1 U2709 ( .B1(n2723), .B2(n2480), .A(n2192), .ZN(n3804) );
  NAND2_X1 U2710 ( .A1(n2723), .A2(n2480), .ZN(n2192) );
  XNOR2_X1 U2711 ( .A(n2555), .B(n2490), .ZN(n2554) );
  INV_X1 U2712 ( .A(n2558), .ZN(n2641) );
  AND2_X1 U2713 ( .A1(n2187), .A2(n2191), .ZN(n2613) );
  NAND2_X1 U2714 ( .A1(n2611), .A2(REG2_REG_6__SCAN_IN), .ZN(n2187) );
  AOI22_X1 U2715 ( .A1(n2605), .A2(REG1_REG_6__SCAN_IN), .B1(n4353), .B2(n2604), .ZN(n2699) );
  NAND2_X1 U2716 ( .A1(n2179), .A2(n2694), .ZN(n2696) );
  INV_X1 U2717 ( .A(n2263), .ZN(n2693) );
  INV_X1 U2718 ( .A(n2256), .ZN(n2704) );
  XNOR2_X1 U2719 ( .A(n3827), .B(n4498), .ZN(n4379) );
  NAND2_X1 U2720 ( .A1(n4379), .A2(REG2_REG_10__SCAN_IN), .ZN(n4378) );
  XNOR2_X1 U2721 ( .A(n3810), .B(n4498), .ZN(n4374) );
  NOR2_X1 U2722 ( .A1(n4384), .A2(n4383), .ZN(n4382) );
  NAND2_X1 U2723 ( .A1(n4398), .A2(n3834), .ZN(n4409) );
  NOR2_X1 U2724 ( .A1(n4415), .A2(n4414), .ZN(n4413) );
  NAND2_X1 U2725 ( .A1(n2250), .A2(n3816), .ZN(n4415) );
  NOR2_X1 U2726 ( .A1(n3839), .A2(n2259), .ZN(n4417) );
  NAND2_X1 U2727 ( .A1(n2260), .A2(n3838), .ZN(n4418) );
  INV_X1 U2728 ( .A(n3839), .ZN(n2260) );
  NOR2_X1 U2729 ( .A1(n2258), .A2(n3839), .ZN(n4430) );
  INV_X1 U2730 ( .A(n2259), .ZN(n2258) );
  NAND2_X1 U2731 ( .A1(n4441), .A2(n3842), .ZN(n4453) );
  INV_X1 U2732 ( .A(n2247), .ZN(n2243) );
  NAND2_X1 U2733 ( .A1(n2245), .A2(n2248), .ZN(n2244) );
  OR2_X1 U2734 ( .A1(n4461), .A2(n2142), .ZN(n2248) );
  AOI21_X1 U2735 ( .B1(n4217), .B2(n4214), .A(n4213), .ZN(n4361) );
  NAND2_X1 U2736 ( .A1(n2281), .A2(n2280), .ZN(n3996) );
  NAND2_X1 U2737 ( .A1(n4037), .A2(n2130), .ZN(n2281) );
  NAND2_X1 U2738 ( .A1(n4037), .A2(n3903), .ZN(n4015) );
  OR2_X1 U2739 ( .A1(n4123), .A2(n2294), .ZN(n2292) );
  NAND2_X1 U2740 ( .A1(n4122), .A2(n3897), .ZN(n4100) );
  OR2_X1 U2741 ( .A1(n4171), .A2(n4172), .ZN(n4270) );
  NAND2_X1 U2742 ( .A1(n2287), .A2(n2286), .ZN(n3205) );
  OR2_X1 U2743 ( .A1(n3140), .A2(n3139), .ZN(n2287) );
  OR2_X1 U2744 ( .A1(n4477), .A2(n4350), .ZN(n4137) );
  INV_X1 U2745 ( .A(n4202), .ZN(n3953) );
  INV_X1 U2746 ( .A(n4479), .ZN(n4195) );
  OR2_X1 U2747 ( .A1(n2589), .A2(n2676), .ZN(n4196) );
  INV_X1 U2748 ( .A(n4216), .ZN(n4127) );
  NAND2_X1 U2749 ( .A1(n2361), .A2(n2360), .ZN(n2577) );
  OR2_X1 U2750 ( .A1(n3349), .A2(n2359), .ZN(n2361) );
  NAND2_X1 U2751 ( .A1(n3349), .A2(DATAI_0_), .ZN(n2360) );
  NOR2_X1 U2752 ( .A1(n2935), .A2(n2679), .ZN(n4547) );
  INV_X1 U2753 ( .A(n4242), .ZN(n4286) );
  INV_X1 U2754 ( .A(n4545), .ZN(n4544) );
  AND2_X1 U2755 ( .A1(n4544), .A2(n4536), .ZN(n4242) );
  INV_X1 U2756 ( .A(n4547), .ZN(n4545) );
  OAI211_X1 U2757 ( .C1(n2200), .C2(n4503), .A(n4223), .B(n2199), .ZN(n4291)
         );
  INV_X1 U2758 ( .A(n4221), .ZN(n2200) );
  INV_X1 U2759 ( .A(n4222), .ZN(n2199) );
  NAND2_X1 U2760 ( .A1(n2591), .A2(n2674), .ZN(n4485) );
  XNOR2_X1 U2761 ( .A(n2319), .B(IR_REG_26__SCAN_IN), .ZN(n4347) );
  OR2_X1 U2762 ( .A1(n2328), .A2(n3189), .ZN(n2319) );
  XNOR2_X1 U2763 ( .A(n2320), .B(IR_REG_25__SCAN_IN), .ZN(n4348) );
  XNOR2_X1 U2764 ( .A(n2323), .B(IR_REG_24__SCAN_IN), .ZN(n4349) );
  AND2_X1 U2765 ( .A1(n2748), .A2(STATE_REG_SCAN_IN), .ZN(n4487) );
  INV_X1 U2766 ( .A(n2411), .ZN(n3774) );
  AND2_X1 U2767 ( .A1(n2367), .A2(n2148), .ZN(n3703) );
  XNOR2_X1 U2768 ( .A(n2689), .B(IR_REG_7__SCAN_IN), .ZN(n4352) );
  INV_X1 U2769 ( .A(IR_REG_3__SCAN_IN), .ZN(n2547) );
  AOI21_X1 U2770 ( .B1(n2132), .B2(n4467), .A(n4466), .ZN(n4474) );
  NAND2_X1 U2771 ( .A1(n4457), .A2(n2244), .ZN(n2242) );
  AND3_X1 U2772 ( .A1(n2317), .A2(n2316), .A3(n2300), .ZN(n2129) );
  AND2_X1 U2773 ( .A1(n2133), .A2(n3903), .ZN(n2130) );
  NAND2_X1 U2774 ( .A1(n3778), .A2(n3250), .ZN(n3251) );
  AND2_X1 U2775 ( .A1(n2186), .A2(n2175), .ZN(n2131) );
  NAND2_X1 U2776 ( .A1(n3296), .A2(n3295), .ZN(n3516) );
  OR2_X1 U2777 ( .A1(n4462), .A2(n4461), .ZN(n2132) );
  INV_X1 U2778 ( .A(n3251), .ZN(n3252) );
  OR2_X1 U2779 ( .A1(n4009), .A2(n4029), .ZN(n2133) );
  AND2_X1 U2780 ( .A1(n2293), .A2(n2291), .ZN(n2134) );
  AND2_X1 U2781 ( .A1(n2956), .A2(n2990), .ZN(n2135) );
  INV_X1 U2782 ( .A(IR_REG_31__SCAN_IN), .ZN(n3189) );
  OAI21_X1 U2783 ( .B1(n3599), .B2(n3595), .A(n3596), .ZN(n3488) );
  AND2_X1 U2784 ( .A1(n2325), .A2(n2318), .ZN(n2136) );
  NOR2_X1 U2785 ( .A1(n3252), .A2(n2274), .ZN(n2273) );
  AND2_X1 U2786 ( .A1(n2147), .A2(n2331), .ZN(n2137) );
  AND2_X1 U2787 ( .A1(n2130), .A2(n3904), .ZN(n2138) );
  AND2_X1 U2788 ( .A1(n3518), .A2(n2215), .ZN(n2139) );
  AND2_X1 U2789 ( .A1(n2212), .A2(n2159), .ZN(n2140) );
  AND2_X1 U2790 ( .A1(n3896), .A2(n4116), .ZN(n2141) );
  NAND2_X1 U2791 ( .A1(n2208), .A2(n2731), .ZN(n2747) );
  XOR2_X1 U2792 ( .A(n4350), .B(REG1_REG_19__SCAN_IN), .Z(n2142) );
  INV_X1 U2793 ( .A(n4457), .ZN(n4460) );
  NAND2_X1 U2794 ( .A1(n2936), .A2(n2793), .ZN(n2817) );
  AND2_X1 U2795 ( .A1(n2252), .A2(REG1_REG_14__SCAN_IN), .ZN(n2143) );
  INV_X1 U2796 ( .A(n2865), .ZN(n2798) );
  OR3_X1 U2797 ( .A1(n4028), .A2(n2202), .A3(n2201), .ZN(n2144) );
  NAND2_X2 U2798 ( .A1(n2434), .A2(n4344), .ZN(n2536) );
  OR2_X1 U2799 ( .A1(n4080), .A2(n3862), .ZN(n2145) );
  NOR2_X1 U2800 ( .A1(n3296), .A2(n3295), .ZN(n2146) );
  NAND2_X1 U2801 ( .A1(n4347), .A2(n2324), .ZN(n2576) );
  AND4_X2 U2802 ( .A1(n2340), .A2(n2339), .A3(n2338), .A4(n2337), .ZN(n2651)
         );
  AND2_X1 U2803 ( .A1(n3259), .A2(n3733), .ZN(n3690) );
  NAND2_X1 U2804 ( .A1(n2351), .A2(n2350), .ZN(n2481) );
  NAND2_X1 U2805 ( .A1(n2229), .A2(n2233), .ZN(n3505) );
  AND2_X1 U2806 ( .A1(n2327), .A2(n4798), .ZN(n2147) );
  NAND2_X1 U2807 ( .A1(n2368), .A2(n2299), .ZN(n2148) );
  AND3_X2 U2808 ( .A1(n2315), .A2(n2197), .A3(n3327), .ZN(n2328) );
  NOR2_X1 U2809 ( .A1(n4413), .A2(n3817), .ZN(n2149) );
  NAND2_X1 U2810 ( .A1(n2368), .A2(n2316), .ZN(n2365) );
  NAND2_X1 U2811 ( .A1(n2419), .A2(n2302), .ZN(n2423) );
  NAND2_X1 U2812 ( .A1(n2358), .A2(n2357), .ZN(n2580) );
  AND2_X1 U2813 ( .A1(n2224), .A2(n2225), .ZN(n2150) );
  INV_X1 U2814 ( .A(IR_REG_2__SCAN_IN), .ZN(n2308) );
  INV_X1 U2815 ( .A(IR_REG_29__SCAN_IN), .ZN(n2331) );
  OAI21_X1 U2816 ( .B1(n4125), .B2(n2297), .A(n3899), .ZN(n2296) );
  AND4_X1 U2817 ( .A1(n2315), .A2(n3327), .A3(n2129), .A4(n2136), .ZN(n2151)
         );
  NAND2_X1 U2818 ( .A1(n3088), .A2(n3551), .ZN(n2152) );
  INV_X1 U2819 ( .A(n2746), .ZN(n2207) );
  NAND2_X1 U2820 ( .A1(n2349), .A2(n2308), .ZN(n2418) );
  INV_X1 U2821 ( .A(n2418), .ZN(n2419) );
  AND2_X1 U2822 ( .A1(n2136), .A2(n2198), .ZN(n2153) );
  AND2_X1 U2823 ( .A1(n2278), .A2(n3906), .ZN(n2154) );
  INV_X1 U2824 ( .A(IR_REG_22__SCAN_IN), .ZN(n2317) );
  INV_X1 U2825 ( .A(n3255), .ZN(n2274) );
  NOR2_X1 U2826 ( .A1(n4028), .A2(n4006), .ZN(n2155) );
  AND2_X1 U2827 ( .A1(n4166), .A2(n4148), .ZN(n2156) );
  NAND2_X1 U2828 ( .A1(n2290), .A2(n2289), .ZN(n4057) );
  NAND2_X1 U2829 ( .A1(n3489), .A2(n2228), .ZN(n2157) );
  NAND2_X1 U2830 ( .A1(n2211), .A2(n2212), .ZN(n3524) );
  NAND2_X1 U2831 ( .A1(n3108), .A2(n3107), .ZN(n3148) );
  NAND2_X1 U2832 ( .A1(n2292), .A2(n2293), .ZN(n4077) );
  INV_X1 U2833 ( .A(n3832), .ZN(n4495) );
  AND2_X1 U2834 ( .A1(n4066), .A2(n4091), .ZN(n2158) );
  OR2_X1 U2835 ( .A1(n3318), .A2(n3525), .ZN(n2159) );
  AND2_X1 U2836 ( .A1(n3496), .A2(n3495), .ZN(n2160) );
  NAND2_X1 U2837 ( .A1(n2275), .A2(n2273), .ZN(n3889) );
  INV_X1 U2838 ( .A(n3228), .ZN(n3229) );
  OR2_X1 U2839 ( .A1(n3188), .A2(n3187), .ZN(n3287) );
  INV_X1 U2840 ( .A(n3027), .ZN(n3005) );
  AND2_X1 U2841 ( .A1(n4009), .A2(n4029), .ZN(n2161) );
  AND2_X1 U2842 ( .A1(n2287), .A2(n2284), .ZN(n2162) );
  INV_X1 U2843 ( .A(n3904), .ZN(n2279) );
  AND2_X1 U2844 ( .A1(n3141), .A2(n3207), .ZN(n2163) );
  NOR2_X1 U2845 ( .A1(n3314), .A2(n3313), .ZN(n2164) );
  NOR2_X1 U2846 ( .A1(n3888), .A2(n3887), .ZN(n2165) );
  NAND2_X1 U2847 ( .A1(n3984), .A2(n3677), .ZN(n2166) );
  NOR2_X1 U2848 ( .A1(n3400), .A2(n3402), .ZN(n2167) );
  NOR2_X1 U2849 ( .A1(n3526), .A2(n3319), .ZN(n2168) );
  AND2_X1 U2850 ( .A1(n2225), .A2(n2223), .ZN(n2169) );
  AND2_X1 U2851 ( .A1(n2862), .A2(n2859), .ZN(n2801) );
  NAND2_X1 U2852 ( .A1(n2747), .A2(n2746), .ZN(n2774) );
  AOI21_X1 U2853 ( .B1(n3093), .B2(n2306), .A(n3092), .ZN(n3140) );
  OR2_X1 U2854 ( .A1(n2782), .A2(n2781), .ZN(n2828) );
  AND2_X1 U2855 ( .A1(n2894), .A2(n2956), .ZN(n2170) );
  NAND2_X1 U2856 ( .A1(n2196), .A2(n3228), .ZN(n3241) );
  INV_X1 U2857 ( .A(n3241), .ZN(n2195) );
  AND2_X1 U2858 ( .A1(n2141), .A2(n4091), .ZN(n2171) );
  NAND2_X1 U2859 ( .A1(n3112), .A2(n3113), .ZN(n2172) );
  NAND2_X1 U2860 ( .A1(n4194), .A2(n4193), .ZN(n4171) );
  AND2_X1 U2861 ( .A1(n2328), .A2(n2327), .ZN(n2382) );
  AND2_X1 U2862 ( .A1(n3830), .A2(REG1_REG_11__SCAN_IN), .ZN(n2173) );
  NAND2_X1 U2863 ( .A1(n3844), .A2(REG1_REG_18__SCAN_IN), .ZN(n2174) );
  INV_X1 U2864 ( .A(n2203), .ZN(n3080) );
  INV_X1 U2865 ( .A(n3990), .ZN(n3983) );
  NAND2_X1 U2866 ( .A1(n3349), .A2(DATAI_25_), .ZN(n3990) );
  NAND2_X1 U2867 ( .A1(n3841), .A2(REG2_REG_15__SCAN_IN), .ZN(n2175) );
  INV_X1 U2868 ( .A(n2817), .ZN(n2818) );
  NAND2_X1 U2869 ( .A1(n2245), .A2(n2243), .ZN(n2176) );
  AND2_X1 U2870 ( .A1(n2135), .A2(n3027), .ZN(n2177) );
  AND2_X1 U2871 ( .A1(n4457), .A2(n2176), .ZN(n2178) );
  INV_X1 U2872 ( .A(n3843), .ZN(n4490) );
  INV_X1 U2873 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2190) );
  INV_X1 U2874 ( .A(n2235), .ZN(n2667) );
  NAND2_X1 U2875 ( .A1(n3696), .A2(n2411), .ZN(n2235) );
  XNOR2_X1 U2876 ( .A(n2550), .B(IR_REG_4__SCAN_IN), .ZN(n4354) );
  INV_X1 U2877 ( .A(n4354), .ZN(n2261) );
  INV_X1 U2878 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2181) );
  OAI211_X1 U2879 ( .C1(n4370), .C2(REG2_REG_8__SCAN_IN), .A(n2179), .B(n4472), 
        .ZN(n4371) );
  NAND2_X1 U2880 ( .A1(n4387), .A2(n3831), .ZN(n3833) );
  INV_X1 U2881 ( .A(n3831), .ZN(n2185) );
  INV_X1 U2882 ( .A(n2186), .ZN(n4429) );
  NAND2_X1 U2883 ( .A1(n2610), .A2(n4353), .ZN(n2191) );
  NAND2_X1 U2884 ( .A1(n3327), .A2(n2194), .ZN(n3315) );
  NAND3_X1 U2885 ( .A1(n2315), .A2(n3327), .A3(n2129), .ZN(n2321) );
  NAND3_X1 U2886 ( .A1(n2177), .A2(n3085), .A3(n2894), .ZN(n2203) );
  NAND2_X1 U2887 ( .A1(n2206), .A2(n2204), .ZN(n2779) );
  INV_X1 U2888 ( .A(n2205), .ZN(n2204) );
  NAND2_X1 U2889 ( .A1(n2730), .A2(n2746), .ZN(n2206) );
  NAND2_X1 U2890 ( .A1(n3296), .A2(n2140), .ZN(n2210) );
  INV_X1 U2891 ( .A(n3619), .ZN(n2216) );
  AND2_X1 U2892 ( .A1(n3480), .A2(n3401), .ZN(n3479) );
  OR2_X1 U2893 ( .A1(n3479), .A2(n3398), .ZN(n3534) );
  NAND2_X1 U2894 ( .A1(n3480), .A2(n2230), .ZN(n2229) );
  OAI21_X1 U2895 ( .B1(n2982), .B2(n2981), .A(n2980), .ZN(n2984) );
  OR2_X2 U2896 ( .A1(n3448), .A2(n4536), .ZN(n3445) );
  NAND2_X1 U2897 ( .A1(n4462), .A2(n2178), .ZN(n2241) );
  OAI211_X1 U2898 ( .C1(n4462), .C2(n2242), .A(n2241), .B(n3852), .ZN(U3259)
         );
  NAND2_X1 U2899 ( .A1(n3817), .A2(n2252), .ZN(n2251) );
  NAND2_X1 U2900 ( .A1(n2251), .A2(n2249), .ZN(n4425) );
  NAND3_X1 U2901 ( .A1(n2250), .A2(n3816), .A3(n2143), .ZN(n2249) );
  INV_X1 U2902 ( .A(n3815), .ZN(n2253) );
  NAND2_X1 U2903 ( .A1(n2701), .A2(n2700), .ZN(n2702) );
  NAND2_X1 U2904 ( .A1(n2703), .A2(n2256), .ZN(n4366) );
  NAND2_X1 U2905 ( .A1(n3632), .A2(REG2_REG_2__SCAN_IN), .ZN(n2378) );
  NAND2_X1 U2906 ( .A1(n3632), .A2(REG2_REG_0__SCAN_IN), .ZN(n2355) );
  NAND2_X1 U2907 ( .A1(n3632), .A2(REG2_REG_8__SCAN_IN), .ZN(n2908) );
  NAND2_X1 U2908 ( .A1(n3632), .A2(REG2_REG_7__SCAN_IN), .ZN(n2882) );
  NAND2_X1 U2909 ( .A1(n3632), .A2(REG2_REG_6__SCAN_IN), .ZN(n2836) );
  NAND2_X1 U2910 ( .A1(n3632), .A2(REG2_REG_5__SCAN_IN), .ZN(n2522) );
  NAND2_X1 U2911 ( .A1(n3632), .A2(REG2_REG_9__SCAN_IN), .ZN(n2449) );
  NAND2_X1 U2912 ( .A1(n3632), .A2(REG2_REG_10__SCAN_IN), .ZN(n2462) );
  NAND2_X1 U2913 ( .A1(n3632), .A2(REG2_REG_25__SCAN_IN), .ZN(n2620) );
  AND3_X2 U2914 ( .A1(n2302), .A2(n2349), .A3(n2268), .ZN(n2422) );
  NAND2_X1 U2915 ( .A1(n3248), .A2(n2273), .ZN(n2270) );
  NAND2_X1 U2916 ( .A1(n2270), .A2(n2271), .ZN(n4179) );
  NAND2_X1 U2917 ( .A1(n4037), .A2(n2138), .ZN(n2277) );
  NAND2_X1 U2918 ( .A1(n2277), .A2(n2154), .ZN(n3979) );
  NAND2_X1 U2919 ( .A1(n3140), .A2(n2284), .ZN(n2283) );
  NAND2_X1 U2920 ( .A1(n2328), .A2(n2147), .ZN(n2330) );
  NAND2_X1 U2921 ( .A1(n2328), .A2(n2137), .ZN(n2288) );
  NAND2_X1 U2922 ( .A1(n4123), .A2(n2134), .ZN(n2290) );
  AND2_X1 U2923 ( .A1(n3327), .A2(n2315), .ZN(n2368) );
  NAND2_X1 U2924 ( .A1(n3701), .A2(n3705), .ZN(n2362) );
  OR2_X1 U2925 ( .A1(n2453), .A2(n2333), .ZN(n2340) );
  NAND2_X1 U2926 ( .A1(n2434), .A2(n2334), .ZN(n2453) );
  OR2_X1 U2927 ( .A1(n2935), .A2(n2934), .ZN(n4790) );
  AND2_X1 U2928 ( .A1(n4351), .A2(REG1_REG_9__SCAN_IN), .ZN(n2301) );
  OR2_X1 U2929 ( .A1(n3843), .A2(REG1_REG_17__SCAN_IN), .ZN(n2303) );
  OR2_X1 U2930 ( .A1(n2698), .A2(n4820), .ZN(n2304) );
  AND2_X1 U2931 ( .A1(n3366), .A2(n3365), .ZN(n2305) );
  OR2_X1 U2932 ( .A1(n2576), .A2(n2439), .ZN(n3783) );
  NAND2_X1 U2933 ( .A1(n2779), .A2(n2778), .ZN(n2782) );
  AOI21_X1 U2934 ( .B1(n2580), .B2(n3416), .A(n2578), .ZN(n2656) );
  NAND2_X1 U2935 ( .A1(n2584), .A2(n2583), .ZN(n2658) );
  INV_X1 U2936 ( .A(n2800), .ZN(n2928) );
  NAND2_X1 U2937 ( .A1(n3019), .A2(n3020), .ZN(n2307) );
  AND4_X1 U2938 ( .A1(n3305), .A2(n3304), .A3(n3303), .A4(n3302), .ZN(n4152)
         );
  INV_X1 U2939 ( .A(n4114), .ZN(n4149) );
  AND4_X1 U2940 ( .A1(n3326), .A2(n3325), .A3(n3324), .A4(n3323), .ZN(n4114)
         );
  NAND2_X1 U2941 ( .A1(n2362), .A2(n2363), .ZN(n2850) );
  INV_X1 U2942 ( .A(IR_REG_18__SCAN_IN), .ZN(n2314) );
  NAND2_X1 U2943 ( .A1(n3397), .A2(n3396), .ZN(n3398) );
  OR2_X1 U2944 ( .A1(n4352), .A2(REG1_REG_7__SCAN_IN), .ZN(n2700) );
  NAND2_X1 U2945 ( .A1(n2926), .A2(n2655), .ZN(n3701) );
  INV_X1 U2946 ( .A(IR_REG_27__SCAN_IN), .ZN(n2343) );
  NAND2_X1 U2947 ( .A1(n3935), .A2(n3954), .ZN(n3912) );
  INV_X1 U2948 ( .A(n3895), .ZN(n3896) );
  NAND2_X1 U2949 ( .A1(n2467), .A2(n4798), .ZN(n2344) );
  AND2_X1 U2950 ( .A1(n3379), .A2(n2618), .ZN(n3410) );
  AND2_X1 U2951 ( .A1(n3935), .A2(n3913), .ZN(n3874) );
  NAND2_X1 U2952 ( .A1(n4114), .A2(n3896), .ZN(n3897) );
  OR2_X1 U2953 ( .A1(n2460), .A2(n2459), .ZN(n2525) );
  INV_X1 U2954 ( .A(n4091), .ZN(n4083) );
  INV_X1 U2955 ( .A(n2884), .ZN(n2887) );
  AND2_X1 U2956 ( .A1(n2442), .A2(n2408), .ZN(n2750) );
  INV_X1 U2957 ( .A(n2971), .ZN(n2990) );
  NAND2_X1 U2958 ( .A1(n3349), .A2(DATAI_1_), .ZN(n2352) );
  INV_X1 U2959 ( .A(n4172), .ZN(n3892) );
  NAND2_X1 U2960 ( .A1(n3349), .A2(DATAI_24_), .ZN(n3905) );
  INV_X1 U2961 ( .A(REG3_REG_15__SCAN_IN), .ZN(n4770) );
  NOR2_X1 U2962 ( .A1(n3378), .A2(n3377), .ZN(n3379) );
  AND4_X1 U2963 ( .A1(n2507), .A2(n2506), .A3(n2505), .A4(n2504), .ZN(n4130)
         );
  AND4_X1 U2964 ( .A1(n2495), .A2(n2494), .A3(n2493), .A4(n2492), .ZN(n3237)
         );
  AOI22_X1 U2965 ( .A1(n2643), .A2(REG1_REG_4__SCAN_IN), .B1(n4354), .B2(n2552), .ZN(n2631) );
  INV_X1 U2966 ( .A(n2683), .ZN(n2685) );
  NOR2_X1 U2967 ( .A1(n3811), .A2(n4373), .ZN(n4384) );
  AOI21_X1 U2968 ( .B1(n4464), .B2(ADDR_REG_18__SCAN_IN), .A(n4463), .ZN(n4465) );
  AND2_X1 U2969 ( .A1(n3883), .A2(n3882), .ZN(n3884) );
  AND4_X1 U2970 ( .A1(n2513), .A2(n2512), .A3(n2511), .A4(n2510), .ZN(n4066)
         );
  AND2_X1 U2971 ( .A1(n3349), .A2(DATAI_28_), .ZN(n3937) );
  INV_X1 U2972 ( .A(n4029), .ZN(n3921) );
  INV_X1 U2973 ( .A(n3249), .ZN(n3250) );
  NAND2_X1 U2974 ( .A1(n4089), .A2(n4540), .ZN(n4525) );
  NOR2_X1 U2975 ( .A1(n2589), .A2(n2750), .ZN(n2678) );
  NAND2_X1 U2976 ( .A1(n2576), .A2(n4487), .ZN(n2589) );
  OR2_X1 U2977 ( .A1(n3163), .A2(n3162), .ZN(n3165) );
  NOR2_X1 U2978 ( .A1(n3337), .A2(n3336), .ZN(n3338) );
  AND2_X1 U2979 ( .A1(n2526), .A2(REG3_REG_12__SCAN_IN), .ZN(n3118) );
  INV_X1 U2980 ( .A(n3905), .ZN(n4006) );
  NAND2_X1 U2981 ( .A1(n3118), .A2(REG3_REG_13__SCAN_IN), .ZN(n3163) );
  INV_X1 U2982 ( .A(n3624), .ZN(n3588) );
  AND2_X1 U2983 ( .A1(n2516), .A2(REG3_REG_5__SCAN_IN), .ZN(n2833) );
  OR2_X1 U2984 ( .A1(n2755), .A2(n2754), .ZN(n3614) );
  AND4_X1 U2985 ( .A1(n3343), .A2(n3342), .A3(n3341), .A4(n3340), .ZN(n4129)
         );
  NAND2_X1 U2986 ( .A1(n2685), .A2(n2684), .ZN(n3154) );
  INV_X1 U2987 ( .A(n4465), .ZN(n4466) );
  AND2_X1 U2988 ( .A1(n2479), .A2(n2636), .ZN(n4457) );
  OAI22_X1 U2989 ( .A1(n3231), .A2(n3230), .B1(n3229), .B2(n3584), .ZN(n3248)
         );
  OAI21_X1 U2990 ( .B1(n2674), .B2(D_REG_0__SCAN_IN), .A(n2440), .ZN(n2679) );
  NAND2_X1 U2991 ( .A1(n3349), .A2(DATAI_26_), .ZN(n3973) );
  NAND2_X1 U2992 ( .A1(n3349), .A2(DATAI_20_), .ZN(n4091) );
  INV_X1 U2993 ( .A(n4110), .ZN(n4116) );
  INV_X1 U2994 ( .A(n4186), .ZN(n4193) );
  AND2_X1 U2995 ( .A1(n2809), .A2(n2808), .ZN(n4511) );
  AND2_X1 U2996 ( .A1(n2412), .A2(n2411), .ZN(n4510) );
  NAND2_X1 U2997 ( .A1(n2395), .A2(n4347), .ZN(n2674) );
  AND2_X1 U2998 ( .A1(n2444), .A2(n2470), .ZN(n4464) );
  INV_X1 U2999 ( .A(n3679), .ZN(n4207) );
  INV_X1 U3000 ( .A(n4192), .ZN(n3888) );
  OR2_X1 U3001 ( .A1(n4477), .A2(n2846), .ZN(n4202) );
  AND3_X1 U3002 ( .A1(n4530), .A2(n4529), .A3(n4528), .ZN(n4546) );
  INV_X1 U3003 ( .A(n4307), .ZN(n4342) );
  INV_X1 U3004 ( .A(n4485), .ZN(n4486) );
  INV_X1 U3005 ( .A(n2334), .ZN(n4344) );
  INV_X1 U3006 ( .A(n3849), .ZN(n4350) );
  INV_X1 U3007 ( .A(n4407), .ZN(n4494) );
  OR2_X1 U3008 ( .A1(n2151), .A2(n3189), .ZN(n2320) );
  NAND2_X1 U3009 ( .A1(n2321), .A2(IR_REG_31__SCAN_IN), .ZN(n2326) );
  NAND2_X1 U3010 ( .A1(n2326), .A2(n2325), .ZN(n2322) );
  NAND2_X1 U3011 ( .A1(n2322), .A2(IR_REG_31__SCAN_IN), .ZN(n2323) );
  XNOR2_X1 U3012 ( .A(n2326), .B(n2325), .ZN(n2748) );
  INV_X1 U3013 ( .A(n4487), .ZN(n2439) );
  INV_X2 U3014 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NOR2_X1 U3015 ( .A1(IR_REG_26__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2327)
         );
  INV_X1 U3016 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2333) );
  INV_X1 U3017 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2414) );
  OR2_X1 U3018 ( .A1(n2536), .A2(n2414), .ZN(n2339) );
  INV_X1 U3019 ( .A(n2434), .ZN(n2336) );
  INV_X1 U3020 ( .A(REG0_REG_1__SCAN_IN), .ZN(n2335) );
  INV_X1 U3021 ( .A(IR_REG_26__SCAN_IN), .ZN(n2341) );
  NAND2_X1 U3022 ( .A1(n2328), .A2(n2341), .ZN(n2342) );
  NAND2_X1 U3023 ( .A1(n4798), .A2(IR_REG_27__SCAN_IN), .ZN(n2346) );
  NAND2_X4 U3024 ( .A1(n2347), .A2(n2346), .ZN(n3349) );
  NAND2_X1 U3025 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2348)
         );
  INV_X1 U3026 ( .A(n2349), .ZN(n2350) );
  INV_X1 U3027 ( .A(n2481), .ZN(n4356) );
  OAI21_X2 U3028 ( .B1(n3349), .B2(n2481), .A(n2352), .ZN(n2760) );
  NAND2_X1 U3029 ( .A1(n2651), .A2(n2760), .ZN(n3705) );
  INV_X1 U3030 ( .A(REG0_REG_0__SCAN_IN), .ZN(n2353) );
  OR2_X1 U3031 ( .A1(n2537), .A2(n2353), .ZN(n2356) );
  NAND2_X1 U3032 ( .A1(n2538), .A2(REG1_REG_0__SCAN_IN), .ZN(n2354) );
  INV_X1 U3033 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2718) );
  INV_X1 U3034 ( .A(n4357), .ZN(n2359) );
  AND2_X1 U3035 ( .A1(n2580), .A2(n2577), .ZN(n2363) );
  OR2_X1 U3036 ( .A1(n2363), .A2(n2362), .ZN(n2364) );
  NAND2_X1 U3037 ( .A1(n2850), .A2(n2364), .ZN(n2712) );
  NAND2_X1 U3038 ( .A1(n2365), .A2(IR_REG_31__SCAN_IN), .ZN(n2366) );
  MUX2_X1 U3039 ( .A(IR_REG_31__SCAN_IN), .B(n2366), .S(IR_REG_21__SCAN_IN), 
        .Z(n2367) );
  INV_X1 U3040 ( .A(n2368), .ZN(n2369) );
  NAND2_X1 U3041 ( .A1(n2372), .A2(IR_REG_31__SCAN_IN), .ZN(n2371) );
  XNOR2_X1 U3042 ( .A(n2652), .B(n3774), .ZN(n2375) );
  NAND2_X1 U3043 ( .A1(n2375), .A2(n3849), .ZN(n4089) );
  INV_X1 U3044 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2376) );
  OR2_X1 U3045 ( .A1(n2536), .A2(n2376), .ZN(n2381) );
  NAND2_X1 U3046 ( .A1(n2538), .A2(REG1_REG_2__SCAN_IN), .ZN(n2380) );
  INV_X1 U3047 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2377) );
  OR2_X1 U3048 ( .A1(n2537), .A2(n2377), .ZN(n2379) );
  NOR2_X1 U3049 ( .A1(n2382), .A2(n3189), .ZN(n2383) );
  MUX2_X1 U3050 ( .A(n3189), .B(n2383), .S(IR_REG_28__SCAN_IN), .Z(n2384) );
  INV_X1 U3051 ( .A(n2384), .ZN(n2385) );
  NAND2_X1 U3052 ( .A1(n2385), .A2(n2330), .ZN(n2635) );
  NAND2_X1 U3053 ( .A1(n2635), .A2(n2442), .ZN(n4128) );
  INV_X1 U3054 ( .A(n3767), .ZN(n2432) );
  AND2_X2 U3055 ( .A1(n2667), .A2(n2432), .ZN(n4216) );
  NAND2_X1 U3056 ( .A1(n2760), .A2(n4216), .ZN(n2387) );
  INV_X1 U3057 ( .A(n2442), .ZN(n2587) );
  INV_X1 U3058 ( .A(n4191), .ZN(n3210) );
  NAND2_X1 U3059 ( .A1(n2580), .A2(n3210), .ZN(n2386) );
  OAI211_X1 U3060 ( .C1(n2764), .C2(n4128), .A(n2387), .B(n2386), .ZN(n2388)
         );
  INV_X1 U3061 ( .A(n2388), .ZN(n2393) );
  INV_X1 U3062 ( .A(n2580), .ZN(n2663) );
  NAND2_X1 U3063 ( .A1(n2663), .A2(n2577), .ZN(n3700) );
  XNOR2_X1 U3064 ( .A(n2362), .B(n3700), .ZN(n2391) );
  NAND2_X1 U3065 ( .A1(n3774), .A2(n4350), .ZN(n2390) );
  NAND2_X1 U3066 ( .A1(n3703), .A2(n2432), .ZN(n2389) );
  NAND2_X2 U3067 ( .A1(n2390), .A2(n2389), .ZN(n4184) );
  NAND2_X1 U3068 ( .A1(n2391), .A2(n4184), .ZN(n2392) );
  OAI211_X1 U3069 ( .C1(n2712), .C2(n4089), .A(n2393), .B(n2392), .ZN(n2714)
         );
  INV_X1 U3070 ( .A(n4348), .ZN(n2406) );
  NAND2_X1 U3071 ( .A1(n2406), .A2(n2409), .ZN(n2394) );
  MUX2_X1 U3072 ( .A(n2409), .B(n2394), .S(B_REG_SCAN_IN), .Z(n2395) );
  INV_X1 U3073 ( .A(n2674), .ZN(n2672) );
  NOR2_X1 U3074 ( .A1(D_REG_5__SCAN_IN), .A2(D_REG_24__SCAN_IN), .ZN(n4810) );
  NOR4_X1 U3075 ( .A1(D_REG_27__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_6__SCAN_IN), .A4(D_REG_7__SCAN_IN), .ZN(n2398) );
  NOR4_X1 U3076 ( .A1(D_REG_13__SCAN_IN), .A2(D_REG_16__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n2397) );
  NOR4_X1 U3077 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2396) );
  AND4_X1 U3078 ( .A1(n4810), .A2(n2398), .A3(n2397), .A4(n2396), .ZN(n2404)
         );
  NOR4_X1 U3079 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_3__SCAN_IN), .A4(D_REG_4__SCAN_IN), .ZN(n2402) );
  NOR4_X1 U3080 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_14__SCAN_IN), .A4(D_REG_2__SCAN_IN), .ZN(n2401) );
  NOR4_X1 U3081 ( .A1(D_REG_19__SCAN_IN), .A2(D_REG_21__SCAN_IN), .A3(
        D_REG_22__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2400) );
  NOR4_X1 U3082 ( .A1(D_REG_8__SCAN_IN), .A2(D_REG_17__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_15__SCAN_IN), .ZN(n2399) );
  AND4_X1 U3083 ( .A1(n2402), .A2(n2401), .A3(n2400), .A4(n2399), .ZN(n2403)
         );
  NAND2_X1 U3084 ( .A1(n2404), .A2(n2403), .ZN(n2671) );
  INV_X1 U3085 ( .A(n2671), .ZN(n2405) );
  NAND2_X1 U3086 ( .A1(n2405), .A2(D_REG_1__SCAN_IN), .ZN(n2407) );
  INV_X1 U3087 ( .A(n4347), .ZN(n2410) );
  NAND2_X1 U3088 ( .A1(n2410), .A2(n2406), .ZN(n2673) );
  INV_X1 U3089 ( .A(n2673), .ZN(n2438) );
  AOI21_X1 U3090 ( .B1(n2672), .B2(n2407), .A(n2438), .ZN(n2585) );
  NAND2_X1 U3091 ( .A1(n3767), .A2(n3849), .ZN(n2408) );
  NAND2_X1 U3092 ( .A1(n2410), .A2(n2409), .ZN(n2440) );
  NAND3_X1 U3093 ( .A1(n2585), .A2(n2678), .A3(n2679), .ZN(n2413) );
  AND2_X1 U3094 ( .A1(n3767), .A2(n4350), .ZN(n2412) );
  NAND2_X1 U3095 ( .A1(n4510), .A2(n3696), .ZN(n2676) );
  MUX2_X1 U3096 ( .A(n2714), .B(REG2_REG_1__SCAN_IN), .S(n4477), .Z(n2417) );
  INV_X1 U3097 ( .A(n4536), .ZN(n4503) );
  NOR2_X2 U3098 ( .A1(n4137), .A2(n4503), .ZN(n4479) );
  OAI21_X1 U3099 ( .B1(n2668), .B2(n2655), .A(n2937), .ZN(n2711) );
  NOR2_X1 U3100 ( .A1(n4195), .A2(n2711), .ZN(n2416) );
  OR2_X1 U3101 ( .A1(n2652), .A2(n3849), .ZN(n2845) );
  OR2_X1 U3102 ( .A1(n4477), .A2(n2845), .ZN(n4099) );
  OAI22_X1 U3103 ( .A1(n2712), .A2(n4099), .B1(n2414), .B2(n4196), .ZN(n2415)
         );
  OR3_X1 U3104 ( .A1(n2417), .A2(n2416), .A3(n2415), .ZN(U3289) );
  INV_X1 U3105 ( .A(DATAI_2_), .ZN(n2420) );
  INV_X1 U3106 ( .A(n2723), .ZN(n3796) );
  MUX2_X1 U3107 ( .A(n2420), .B(n3796), .S(STATE_REG_SCAN_IN), .Z(n2421) );
  INV_X1 U3108 ( .A(n2421), .ZN(U3350) );
  INV_X1 U3109 ( .A(n2422), .ZN(n2426) );
  NAND2_X1 U3110 ( .A1(n2423), .A2(IR_REG_31__SCAN_IN), .ZN(n2424) );
  MUX2_X1 U3111 ( .A(IR_REG_31__SCAN_IN), .B(n2424), .S(IR_REG_5__SCAN_IN), 
        .Z(n2425) );
  NAND2_X1 U3112 ( .A1(n2426), .A2(n2425), .ZN(n2829) );
  INV_X1 U3113 ( .A(DATAI_5_), .ZN(n2427) );
  MUX2_X1 U3114 ( .A(n2829), .B(n2427), .S(U3149), .Z(n2428) );
  INV_X1 U3115 ( .A(n2428), .ZN(U3347) );
  INV_X1 U3116 ( .A(DATAI_21_), .ZN(n4555) );
  NAND2_X1 U3117 ( .A1(n3703), .A2(STATE_REG_SCAN_IN), .ZN(n2429) );
  OAI21_X1 U3118 ( .B1(STATE_REG_SCAN_IN), .B2(n4555), .A(n2429), .ZN(U3331)
         );
  INV_X1 U3119 ( .A(DATAI_22_), .ZN(n2431) );
  NAND2_X1 U3120 ( .A1(n3774), .A2(STATE_REG_SCAN_IN), .ZN(n2430) );
  OAI21_X1 U3121 ( .B1(STATE_REG_SCAN_IN), .B2(n2431), .A(n2430), .ZN(U3330)
         );
  INV_X1 U3122 ( .A(DATAI_20_), .ZN(n4558) );
  NAND2_X1 U3123 ( .A1(n2432), .A2(STATE_REG_SCAN_IN), .ZN(n2433) );
  OAI21_X1 U3124 ( .B1(STATE_REG_SCAN_IN), .B2(n4558), .A(n2433), .ZN(U3332)
         );
  INV_X1 U3125 ( .A(DATAI_30_), .ZN(n2436) );
  NAND2_X1 U3126 ( .A1(n2434), .A2(STATE_REG_SCAN_IN), .ZN(n2435) );
  OAI21_X1 U3127 ( .B1(STATE_REG_SCAN_IN), .B2(n2436), .A(n2435), .ZN(U3322)
         );
  INV_X1 U3128 ( .A(DATAI_31_), .ZN(n4549) );
  OR4_X1 U3129 ( .A1(n2288), .A2(IR_REG_30__SCAN_IN), .A3(U3149), .A4(n3189), 
        .ZN(n2437) );
  OAI21_X1 U3130 ( .B1(STATE_REG_SCAN_IN), .B2(n4549), .A(n2437), .ZN(U3321)
         );
  INV_X1 U3131 ( .A(n2589), .ZN(n2591) );
  INV_X1 U3132 ( .A(D_REG_1__SCAN_IN), .ZN(n4605) );
  AOI22_X1 U3133 ( .A1(n4485), .A2(n4605), .B1(n2438), .B2(n4487), .ZN(U3459)
         );
  OAI22_X1 U3134 ( .A1(n4486), .A2(D_REG_0__SCAN_IN), .B1(n2440), .B2(n2439), 
        .ZN(n2441) );
  INV_X1 U3135 ( .A(n2441), .ZN(U3458) );
  NAND2_X1 U3136 ( .A1(n2442), .A2(n2748), .ZN(n2443) );
  INV_X1 U3137 ( .A(n2471), .ZN(n2444) );
  OR2_X1 U3138 ( .A1(n2748), .A2(U3149), .ZN(n3776) );
  NAND2_X1 U3139 ( .A1(n2589), .A2(n3776), .ZN(n2470) );
  NOR2_X1 U3140 ( .A1(n4464), .A2(U4043), .ZN(U3148) );
  INV_X1 U3141 ( .A(DATAO_REG_9__SCAN_IN), .ZN(n4746) );
  NAND2_X1 U3142 ( .A1(REG3_REG_7__SCAN_IN), .A2(REG3_REG_8__SCAN_IN), .ZN(
        n2445) );
  NAND2_X1 U3143 ( .A1(n2904), .A2(REG3_REG_9__SCAN_IN), .ZN(n2460) );
  OR2_X1 U3144 ( .A1(n2904), .A2(REG3_REG_9__SCAN_IN), .ZN(n2446) );
  NAND2_X1 U3145 ( .A1(n2460), .A2(n2446), .ZN(n3552) );
  OR2_X1 U3146 ( .A1(n2536), .A2(n3552), .ZN(n2451) );
  INV_X1 U3147 ( .A(REG0_REG_9__SCAN_IN), .ZN(n2447) );
  OR2_X1 U31480 ( .A1(n3634), .A2(n2447), .ZN(n2450) );
  NAND2_X1 U31490 ( .A1(n3297), .A2(REG1_REG_9__SCAN_IN), .ZN(n2448) );
  NAND2_X1 U3150 ( .A1(n3088), .A2(U4043), .ZN(n2452) );
  OAI21_X1 U3151 ( .B1(U4043), .B2(n4746), .A(n2452), .ZN(U3559) );
  INV_X1 U3152 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n4837) );
  INV_X1 U3153 ( .A(REG0_REG_30__SCAN_IN), .ZN(n2456) );
  INV_X4 U3154 ( .A(n2453), .ZN(n3632) );
  NAND2_X1 U3155 ( .A1(n3632), .A2(REG2_REG_30__SCAN_IN), .ZN(n2455) );
  NAND2_X1 U3156 ( .A1(n3297), .A2(REG1_REG_30__SCAN_IN), .ZN(n2454) );
  OAI211_X1 U3157 ( .C1(n3634), .C2(n2456), .A(n2455), .B(n2454), .ZN(n3881)
         );
  NAND2_X1 U3158 ( .A1(n3881), .A2(U4043), .ZN(n2457) );
  OAI21_X1 U3159 ( .B1(U4043), .B2(n4837), .A(n2457), .ZN(U3580) );
  INV_X1 U3160 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n4749) );
  INV_X1 U3161 ( .A(REG0_REG_10__SCAN_IN), .ZN(n2458) );
  OR2_X1 U3162 ( .A1(n3634), .A2(n2458), .ZN(n2465) );
  INV_X1 U3163 ( .A(n2536), .ZN(n3439) );
  NAND2_X1 U3164 ( .A1(n2460), .A2(n2459), .ZN(n2461) );
  NAND2_X1 U3165 ( .A1(n2525), .A2(n2461), .ZN(n3081) );
  OR2_X1 U3166 ( .A1(n3459), .A2(n3081), .ZN(n2464) );
  NAND2_X1 U3167 ( .A1(n3297), .A2(REG1_REG_10__SCAN_IN), .ZN(n2463) );
  NAND2_X1 U3168 ( .A1(n3585), .A2(U4043), .ZN(n2466) );
  OAI21_X1 U3169 ( .B1(U4043), .B2(n4749), .A(n2466), .ZN(U3560) );
  XNOR2_X1 U3170 ( .A(n2467), .B(IR_REG_27__SCAN_IN), .ZN(n4346) );
  INV_X1 U3171 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2719) );
  AND2_X1 U3172 ( .A1(n4346), .A2(n2719), .ZN(n2468) );
  NOR2_X1 U3173 ( .A1(n2635), .A2(n2468), .ZN(n2640) );
  OAI21_X1 U3174 ( .B1(REG1_REG_0__SCAN_IN), .B2(n4346), .A(n2640), .ZN(n2469)
         );
  MUX2_X1 U3175 ( .A(n2469), .B(n2640), .S(n4357), .Z(n2475) );
  INV_X1 U3176 ( .A(n2479), .ZN(n2474) );
  AOI22_X1 U3177 ( .A1(n4464), .A2(ADDR_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n2473) );
  INV_X1 U3178 ( .A(n4346), .ZN(n2636) );
  INV_X1 U3179 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4831) );
  NAND3_X1 U3180 ( .A1(n4457), .A2(n4357), .A3(n4831), .ZN(n2472) );
  OAI211_X1 U3181 ( .C1(n2475), .C2(n2474), .A(n2473), .B(n2472), .ZN(U3240)
         );
  XNOR2_X1 U3182 ( .A(n2548), .B(IR_REG_3__SCAN_IN), .ZN(n4355) );
  INV_X1 U3183 ( .A(n4355), .ZN(n2490) );
  NAND2_X1 U3184 ( .A1(n2479), .A2(n2635), .ZN(n4475) );
  INV_X1 U3185 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2476) );
  XNOR2_X1 U3186 ( .A(n2481), .B(REG1_REG_1__SCAN_IN), .ZN(n3788) );
  AND2_X1 U3187 ( .A1(n4357), .A2(REG1_REG_0__SCAN_IN), .ZN(n3787) );
  NAND2_X1 U3188 ( .A1(n3788), .A2(n3787), .ZN(n2478) );
  NAND2_X1 U3189 ( .A1(n4356), .A2(REG1_REG_1__SCAN_IN), .ZN(n2477) );
  NAND2_X1 U3190 ( .A1(n2478), .A2(n2477), .ZN(n3798) );
  XNOR2_X1 U3191 ( .A(n2544), .B(n4355), .ZN(n2546) );
  XOR2_X1 U3192 ( .A(n2546), .B(REG1_REG_3__SCAN_IN), .Z(n2487) );
  NOR2_X1 U3193 ( .A1(n2635), .A2(n2636), .ZN(n3772) );
  INV_X1 U3194 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2480) );
  AND2_X1 U3195 ( .A1(n4357), .A2(REG2_REG_0__SCAN_IN), .ZN(n3786) );
  NAND2_X1 U3196 ( .A1(n3785), .A2(n3786), .ZN(n3784) );
  NAND2_X1 U3197 ( .A1(n4356), .A2(REG2_REG_1__SCAN_IN), .ZN(n2484) );
  NAND2_X1 U3198 ( .A1(n3784), .A2(n2484), .ZN(n3803) );
  NAND2_X1 U3199 ( .A1(n2723), .A2(REG2_REG_2__SCAN_IN), .ZN(n2485) );
  INV_X1 U3200 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2768) );
  XNOR2_X1 U3201 ( .A(n2554), .B(n2768), .ZN(n2486) );
  AOI22_X1 U3202 ( .A1(n4457), .A2(n2487), .B1(n4472), .B2(n2486), .ZN(n2489)
         );
  AOI22_X1 U3203 ( .A1(n4464), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n2488) );
  OAI211_X1 U3204 ( .C1(n2490), .C2(n4475), .A(n2489), .B(n2488), .ZN(U3243)
         );
  INV_X1 U3205 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n4756) );
  NAND2_X1 U3206 ( .A1(n3632), .A2(REG2_REG_12__SCAN_IN), .ZN(n2495) );
  NAND2_X1 U3207 ( .A1(n3297), .A2(REG1_REG_12__SCAN_IN), .ZN(n2494) );
  NOR2_X1 U3208 ( .A1(n2526), .A2(REG3_REG_12__SCAN_IN), .ZN(n2491) );
  OR2_X1 U3209 ( .A1(n3118), .A2(n2491), .ZN(n3143) );
  OR2_X1 U32100 ( .A1(n3459), .A2(n3143), .ZN(n2493) );
  INV_X1 U32110 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4649) );
  OR2_X1 U32120 ( .A1(n3634), .A2(n4649), .ZN(n2492) );
  NAND2_X1 U32130 ( .A1(n3584), .A2(U4043), .ZN(n2496) );
  OAI21_X1 U32140 ( .B1(U4043), .B2(n4756), .A(n2496), .ZN(U3562) );
  INV_X1 U32150 ( .A(DATAO_REG_15__SCAN_IN), .ZN(n4755) );
  NAND2_X1 U32160 ( .A1(n3632), .A2(REG2_REG_15__SCAN_IN), .ZN(n2501) );
  NAND2_X1 U32170 ( .A1(n3297), .A2(REG1_REG_15__SCAN_IN), .ZN(n2500) );
  NAND2_X1 U32180 ( .A1(n3165), .A2(n4770), .ZN(n2497) );
  NAND2_X1 U32190 ( .A1(n3299), .A2(n2497), .ZN(n4197) );
  OR2_X1 U32200 ( .A1(n2536), .A2(n4197), .ZN(n2499) );
  INV_X1 U32210 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4332) );
  OR2_X1 U32220 ( .A1(n3634), .A2(n4332), .ZN(n2498) );
  NAND2_X1 U32230 ( .A1(n3890), .A2(U4043), .ZN(n2502) );
  OAI21_X1 U32240 ( .B1(U4043), .B2(n4755), .A(n2502), .ZN(U3565) );
  INV_X1 U32250 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n4759) );
  NAND2_X1 U32260 ( .A1(n3297), .A2(REG1_REG_17__SCAN_IN), .ZN(n2507) );
  NAND2_X1 U32270 ( .A1(n3632), .A2(REG2_REG_17__SCAN_IN), .ZN(n2506) );
  INV_X1 U32280 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4652) );
  OR2_X1 U32290 ( .A1(n3634), .A2(n4652), .ZN(n2505) );
  INV_X1 U32300 ( .A(REG3_REG_16__SCAN_IN), .ZN(n3298) );
  NAND2_X1 U32310 ( .A1(n3300), .A2(REG3_REG_17__SCAN_IN), .ZN(n3321) );
  OR2_X1 U32320 ( .A1(n3300), .A2(REG3_REG_17__SCAN_IN), .ZN(n2503) );
  NAND2_X1 U32330 ( .A1(n3321), .A2(n2503), .ZN(n4157) );
  OR2_X1 U32340 ( .A1(n2536), .A2(n4157), .ZN(n2504) );
  NAND2_X1 U32350 ( .A1(n4166), .A2(U4043), .ZN(n2508) );
  OAI21_X1 U32360 ( .B1(U4043), .B2(n4759), .A(n2508), .ZN(U3567) );
  INV_X1 U32370 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n4758) );
  NAND2_X1 U32380 ( .A1(n3297), .A2(REG1_REG_20__SCAN_IN), .ZN(n2513) );
  NAND2_X1 U32390 ( .A1(n3632), .A2(REG2_REG_20__SCAN_IN), .ZN(n2512) );
  INV_X1 U32400 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4773) );
  INV_X1 U32410 ( .A(REG3_REG_19__SCAN_IN), .ZN(n3336) );
  NOR2_X1 U32420 ( .A1(n3338), .A2(REG3_REG_20__SCAN_IN), .ZN(n2509) );
  OR2_X1 U32430 ( .A1(n3355), .A2(n2509), .ZN(n4093) );
  OR2_X1 U32440 ( .A1(n3459), .A2(n4093), .ZN(n2511) );
  INV_X1 U32450 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4319) );
  OR2_X1 U32460 ( .A1(n3634), .A2(n4319), .ZN(n2510) );
  INV_X1 U32470 ( .A(n4066), .ZN(n4111) );
  NAND2_X1 U32480 ( .A1(n4111), .A2(U4043), .ZN(n2514) );
  OAI21_X1 U32490 ( .B1(U4043), .B2(n4758), .A(n2514), .ZN(U3570) );
  INV_X1 U32500 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n4836) );
  NAND2_X1 U32510 ( .A1(n3297), .A2(REG1_REG_5__SCAN_IN), .ZN(n2523) );
  INV_X1 U32520 ( .A(REG0_REG_5__SCAN_IN), .ZN(n2515) );
  OR2_X1 U32530 ( .A1(n3634), .A2(n2515), .ZN(n2521) );
  INV_X1 U32540 ( .A(n2833), .ZN(n2519) );
  INV_X1 U32550 ( .A(n2516), .ZN(n2535) );
  INV_X1 U32560 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2517) );
  NAND2_X1 U32570 ( .A1(n2535), .A2(n2517), .ZN(n2518) );
  NAND2_X1 U32580 ( .A1(n2519), .A2(n2518), .ZN(n2870) );
  OR2_X1 U32590 ( .A1(n2536), .A2(n2870), .ZN(n2520) );
  INV_X1 U32600 ( .A(n2955), .ZN(n2888) );
  NAND2_X1 U32610 ( .A1(n2888), .A2(U4043), .ZN(n2524) );
  OAI21_X1 U32620 ( .B1(U4043), .B2(n4836), .A(n2524), .ZN(U3555) );
  INV_X1 U32630 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n4748) );
  NAND2_X1 U32640 ( .A1(n3297), .A2(REG1_REG_11__SCAN_IN), .ZN(n2531) );
  NAND2_X1 U32650 ( .A1(n3632), .A2(REG2_REG_11__SCAN_IN), .ZN(n2530) );
  INV_X1 U32660 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3216) );
  OR2_X1 U32670 ( .A1(n3634), .A2(n3216), .ZN(n2529) );
  AND2_X1 U32680 ( .A1(n2525), .A2(n4775), .ZN(n2527) );
  OR2_X1 U32690 ( .A1(n2527), .A2(n2526), .ZN(n3589) );
  OR2_X1 U32700 ( .A1(n3459), .A2(n3589), .ZN(n2528) );
  INV_X1 U32710 ( .A(n3141), .ZN(n3130) );
  NAND2_X1 U32720 ( .A1(n3130), .A2(U4043), .ZN(n2532) );
  OAI21_X1 U32730 ( .B1(U4043), .B2(n4748), .A(n2532), .ZN(U3561) );
  INV_X1 U32740 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n4740) );
  NAND2_X1 U32750 ( .A1(n2926), .A2(U4043), .ZN(n2533) );
  OAI21_X1 U32760 ( .B1(U4043), .B2(n4740), .A(n2533), .ZN(U3551) );
  INV_X1 U32770 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n4743) );
  NOR2_X1 U32780 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n4796) );
  INV_X1 U32790 ( .A(n4796), .ZN(n2534) );
  NAND2_X1 U32800 ( .A1(n2535), .A2(n2534), .ZN(n2820) );
  OR2_X1 U32810 ( .A1(n2536), .A2(n2820), .ZN(n2542) );
  NAND2_X1 U32820 ( .A1(n2538), .A2(REG1_REG_4__SCAN_IN), .ZN(n2540) );
  NAND2_X1 U32830 ( .A1(n2798), .A2(U4043), .ZN(n2543) );
  OAI21_X1 U32840 ( .B1(U4043), .B2(n4743), .A(n2543), .ZN(U3554) );
  INV_X1 U32850 ( .A(n2829), .ZN(n2559) );
  NOR2_X1 U32860 ( .A1(n2544), .A2(n2490), .ZN(n2545) );
  AOI21_X1 U32870 ( .B1(n2546), .B2(REG1_REG_3__SCAN_IN), .A(n2545), .ZN(n2551) );
  NAND2_X1 U32880 ( .A1(n2548), .A2(n2547), .ZN(n2549) );
  NAND2_X1 U32890 ( .A1(n2549), .A2(IR_REG_31__SCAN_IN), .ZN(n2550) );
  XNOR2_X1 U32900 ( .A(n2551), .B(n4354), .ZN(n2643) );
  INV_X1 U32910 ( .A(n2551), .ZN(n2552) );
  INV_X1 U32920 ( .A(REG1_REG_5__SCAN_IN), .ZN(n4534) );
  MUX2_X1 U32930 ( .A(REG1_REG_5__SCAN_IN), .B(n4534), .S(n2829), .Z(n2630) );
  NOR2_X1 U32940 ( .A1(n2631), .A2(n2630), .ZN(n2629) );
  OR2_X1 U32950 ( .A1(n2422), .A2(n3189), .ZN(n2553) );
  XNOR2_X1 U32960 ( .A(n2553), .B(IR_REG_6__SCAN_IN), .ZN(n4353) );
  XNOR2_X1 U32970 ( .A(n2603), .B(n4353), .ZN(n2605) );
  XNOR2_X1 U32980 ( .A(n2605), .B(REG1_REG_6__SCAN_IN), .ZN(n2565) );
  INV_X1 U32990 ( .A(REG3_REG_6__SCAN_IN), .ZN(n4828) );
  NOR2_X1 U33000 ( .A1(STATE_REG_SCAN_IN), .A2(n4828), .ZN(n2957) );
  INV_X1 U33010 ( .A(ADDR_REG_6__SCAN_IN), .ZN(n4731) );
  INV_X1 U33020 ( .A(n4464), .ZN(n4436) );
  NAND2_X1 U33030 ( .A1(n2555), .A2(n4355), .ZN(n2556) );
  AOI22_X1 U33040 ( .A1(n2558), .A2(REG2_REG_4__SCAN_IN), .B1(n4354), .B2(
        n2557), .ZN(n2625) );
  INV_X1 U33050 ( .A(REG2_REG_5__SCAN_IN), .ZN(n4693) );
  MUX2_X1 U33060 ( .A(REG2_REG_5__SCAN_IN), .B(n4693), .S(n2829), .Z(n2624) );
  NOR2_X1 U33070 ( .A1(n2625), .A2(n2624), .ZN(n2623) );
  XNOR2_X1 U33080 ( .A(n2611), .B(n2190), .ZN(n2560) );
  NAND2_X1 U33090 ( .A1(n2560), .A2(n4472), .ZN(n2561) );
  OAI21_X1 U33100 ( .B1(n4731), .B2(n4436), .A(n2561), .ZN(n2562) );
  NOR2_X1 U33110 ( .A1(n2957), .A2(n2562), .ZN(n2564) );
  INV_X1 U33120 ( .A(n4475), .ZN(n4422) );
  NAND2_X1 U33130 ( .A1(n4422), .A2(n4353), .ZN(n2563) );
  OAI211_X1 U33140 ( .C1(n2565), .C2(n4460), .A(n2564), .B(n2563), .ZN(U3246)
         );
  INV_X1 U33150 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n4744) );
  INV_X1 U33160 ( .A(REG0_REG_3__SCAN_IN), .ZN(n2566) );
  OR2_X1 U33170 ( .A1(n2453), .A2(n2768), .ZN(n2792) );
  NAND2_X1 U33180 ( .A1(n3297), .A2(REG1_REG_3__SCAN_IN), .ZN(n2790) );
  NAND2_X1 U33190 ( .A1(n2800), .A2(U4043), .ZN(n2567) );
  OAI21_X1 U33200 ( .B1(U4043), .B2(n4744), .A(n2567), .ZN(U3553) );
  INV_X1 U33210 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n4762) );
  INV_X1 U33220 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3571) );
  INV_X1 U33230 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3377) );
  INV_X1 U33240 ( .A(REG3_REG_24__SCAN_IN), .ZN(n2568) );
  XNOR2_X1 U33250 ( .A(n3379), .B(n2568), .ZN(n3998) );
  NAND2_X1 U33260 ( .A1(n3998), .A2(n3439), .ZN(n2573) );
  INV_X1 U33270 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4654) );
  NAND2_X1 U33280 ( .A1(n3632), .A2(REG2_REG_24__SCAN_IN), .ZN(n2570) );
  NAND2_X1 U33290 ( .A1(n3297), .A2(REG1_REG_24__SCAN_IN), .ZN(n2569) );
  OAI211_X1 U33300 ( .C1(n4654), .C2(n3634), .A(n2570), .B(n2569), .ZN(n2571)
         );
  INV_X1 U33310 ( .A(n2571), .ZN(n2572) );
  NAND2_X1 U33320 ( .A1(n4023), .A2(U4043), .ZN(n2574) );
  OAI21_X1 U33330 ( .B1(U4043), .B2(n4762), .A(n2574), .ZN(U3574) );
  INV_X1 U33340 ( .A(n2652), .ZN(n2575) );
  AND2_X1 U33350 ( .A1(n2577), .A2(n3417), .ZN(n2578) );
  INV_X1 U33360 ( .A(n2576), .ZN(n2581) );
  NAND2_X1 U33370 ( .A1(n2581), .A2(REG1_REG_0__SCAN_IN), .ZN(n2579) );
  NAND2_X1 U33380 ( .A1(n2656), .A2(n2579), .ZN(n2584) );
  AOI22_X1 U33390 ( .A1(n2577), .A2(n3416), .B1(n2581), .B2(n4357), .ZN(n2582)
         );
  OAI21_X1 U33400 ( .B1(n2584), .B2(n2583), .A(n2658), .ZN(n2637) );
  INV_X1 U33410 ( .A(n2679), .ZN(n2934) );
  NAND2_X1 U33420 ( .A1(n2934), .A2(n2585), .ZN(n2662) );
  NAND2_X1 U33430 ( .A1(n2667), .A2(n4350), .ZN(n2586) );
  NAND2_X1 U33440 ( .A1(n2587), .A2(n2586), .ZN(n2588) );
  OR2_X1 U33450 ( .A1(n2588), .A2(n4216), .ZN(n2597) );
  OR2_X1 U33460 ( .A1(n2589), .A2(n2597), .ZN(n2590) );
  INV_X1 U33470 ( .A(n2662), .ZN(n2592) );
  NAND3_X1 U33480 ( .A1(n2592), .A2(n4216), .A3(n2591), .ZN(n2593) );
  NAND2_X1 U33490 ( .A1(n3774), .A2(n3849), .ZN(n2653) );
  INV_X1 U33500 ( .A(n2653), .ZN(n2594) );
  NAND2_X1 U33510 ( .A1(n4487), .A2(n2594), .ZN(n2595) );
  NAND2_X1 U33520 ( .A1(n3771), .A2(n2635), .ZN(n2596) );
  AOI22_X1 U3353 ( .A1(n3588), .A2(n2577), .B1(n2926), .B2(n3583), .ZN(n2602)
         );
  NAND2_X1 U33540 ( .A1(n2597), .A2(n4127), .ZN(n2598) );
  NAND2_X1 U3355 ( .A1(n2662), .A2(n2598), .ZN(n2753) );
  INV_X1 U3356 ( .A(n2753), .ZN(n2600) );
  AND2_X1 U3357 ( .A1(n2662), .A2(n3771), .ZN(n2754) );
  INV_X1 U3358 ( .A(n2678), .ZN(n2599) );
  NOR3_X1 U3359 ( .A1(n2600), .A2(n2754), .A3(n2599), .ZN(n2734) );
  OR2_X1 U3360 ( .A1(n2734), .A2(n2718), .ZN(n2601) );
  OAI211_X1 U3361 ( .C1(n2637), .C2(n3616), .A(n2602), .B(n2601), .ZN(U3229)
         );
  INV_X1 U3362 ( .A(n2603), .ZN(n2604) );
  INV_X1 U3363 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4820) );
  NAND2_X1 U3364 ( .A1(n2422), .A2(n2606), .ZN(n2681) );
  NAND2_X1 U3365 ( .A1(n2681), .A2(IR_REG_31__SCAN_IN), .ZN(n2689) );
  MUX2_X1 U3366 ( .A(n4820), .B(REG1_REG_7__SCAN_IN), .S(n4352), .Z(n2607) );
  XNOR2_X1 U3367 ( .A(n2699), .B(n2607), .ZN(n2617) );
  AND2_X1 U3368 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n2987) );
  AOI21_X1 U3369 ( .B1(n4464), .B2(ADDR_REG_7__SCAN_IN), .A(n2987), .ZN(n2608)
         );
  INV_X1 U3370 ( .A(n2608), .ZN(n2615) );
  INV_X1 U3371 ( .A(n2609), .ZN(n2610) );
  INV_X1 U3372 ( .A(REG2_REG_7__SCAN_IN), .ZN(n4821) );
  MUX2_X1 U3373 ( .A(n4821), .B(REG2_REG_7__SCAN_IN), .S(n4352), .Z(n2612) );
  INV_X1 U3374 ( .A(n4472), .ZN(n4416) );
  AOI211_X1 U3375 ( .C1(n2613), .C2(n2612), .A(n4416), .B(n2687), .ZN(n2614)
         );
  AOI211_X1 U3376 ( .C1(n4422), .C2(n4352), .A(n2615), .B(n2614), .ZN(n2616)
         );
  OAI21_X1 U3377 ( .B1(n4460), .B2(n2617), .A(n2616), .ZN(U3247) );
  INV_X1 U3378 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n4761) );
  AND2_X1 U3379 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG3_REG_24__SCAN_IN), .ZN(
        n2618) );
  AOI21_X1 U3380 ( .B1(n3379), .B2(REG3_REG_24__SCAN_IN), .A(
        REG3_REG_25__SCAN_IN), .ZN(n2619) );
  OR2_X1 U3381 ( .A1(n3410), .A2(n2619), .ZN(n3510) );
  INV_X1 U3382 ( .A(n3634), .ZN(n3412) );
  AOI22_X1 U3383 ( .A1(n3412), .A2(REG0_REG_25__SCAN_IN), .B1(n3297), .B2(
        REG1_REG_25__SCAN_IN), .ZN(n2621) );
  NAND2_X1 U3384 ( .A1(n4005), .A2(U4043), .ZN(n2622) );
  OAI21_X1 U3385 ( .B1(U4043), .B2(n4761), .A(n2622), .ZN(U3575) );
  AND2_X1 U3386 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n2839) );
  INV_X1 U3387 ( .A(ADDR_REG_5__SCAN_IN), .ZN(n4730) );
  AOI211_X1 U3388 ( .C1(n2625), .C2(n2624), .A(n2623), .B(n4416), .ZN(n2626)
         );
  INV_X1 U3389 ( .A(n2626), .ZN(n2627) );
  OAI21_X1 U3390 ( .B1(n4730), .B2(n4436), .A(n2627), .ZN(n2628) );
  NOR2_X1 U3391 ( .A1(n2839), .A2(n2628), .ZN(n2634) );
  AOI211_X1 U3392 ( .C1(n2631), .C2(n2630), .A(n2629), .B(n4460), .ZN(n2632)
         );
  INV_X1 U3393 ( .A(n2632), .ZN(n2633) );
  OAI211_X1 U3394 ( .C1(n4475), .C2(n2829), .A(n2634), .B(n2633), .ZN(U3245)
         );
  INV_X1 U3395 ( .A(n2635), .ZN(n4345) );
  NAND3_X1 U3396 ( .A1(n2637), .A2(n4345), .A3(n2636), .ZN(n2639) );
  AOI21_X1 U3397 ( .B1(n3772), .B2(n3786), .A(n3783), .ZN(n2638) );
  OAI211_X1 U3398 ( .C1(n4357), .C2(n2640), .A(n2639), .B(n2638), .ZN(n3808)
         );
  XNOR2_X1 U3399 ( .A(n2641), .B(REG2_REG_4__SCAN_IN), .ZN(n2647) );
  NAND2_X1 U3400 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n2785) );
  NAND2_X1 U3401 ( .A1(n4464), .A2(ADDR_REG_4__SCAN_IN), .ZN(n2642) );
  OAI211_X1 U3402 ( .C1(n4475), .C2(n2261), .A(n2785), .B(n2642), .ZN(n2646)
         );
  XNOR2_X1 U3403 ( .A(n2643), .B(REG1_REG_4__SCAN_IN), .ZN(n2644) );
  NOR2_X1 U3404 ( .A1(n4460), .A2(n2644), .ZN(n2645) );
  AOI211_X1 U3405 ( .C1(n4472), .C2(n2647), .A(n2646), .B(n2645), .ZN(n2648)
         );
  NAND2_X1 U3406 ( .A1(n3808), .A2(n2648), .ZN(U3244) );
  XNOR2_X1 U3407 ( .A(n2654), .B(n3434), .ZN(n2725) );
  XNOR2_X1 U3408 ( .A(n2725), .B(n2726), .ZN(n2659) );
  NAND2_X1 U3409 ( .A1(n2656), .A2(n3434), .ZN(n2657) );
  NAND2_X1 U3410 ( .A1(n2658), .A2(n2657), .ZN(n2660) );
  NAND2_X1 U3411 ( .A1(n2660), .A2(n2659), .ZN(n2729) );
  OAI211_X1 U3412 ( .C1(n2659), .C2(n2660), .A(n2729), .B(n3621), .ZN(n2666)
         );
  NAND2_X1 U3413 ( .A1(n3771), .A2(n4345), .ZN(n2661) );
  OAI22_X1 U3414 ( .A1(n2663), .A2(n3623), .B1(n2764), .B2(n3626), .ZN(n2664)
         );
  AOI21_X1 U3415 ( .B1(n2760), .B2(n3588), .A(n2664), .ZN(n2665) );
  OAI211_X1 U3416 ( .C1(n2734), .C2(n2414), .A(n2666), .B(n2665), .ZN(U3219)
         );
  NAND2_X1 U3417 ( .A1(n2580), .A2(n2668), .ZN(n3702) );
  NAND2_X1 U3418 ( .A1(n3700), .A2(n3702), .ZN(n3684) );
  NOR2_X1 U3419 ( .A1(n2668), .A2(n2235), .ZN(n2670) );
  INV_X1 U3420 ( .A(n4089), .ZN(n2814) );
  OAI21_X1 U3421 ( .B1(n2814), .B2(n4184), .A(n3684), .ZN(n2669) );
  OAI21_X1 U3422 ( .B1(n2651), .B2(n4128), .A(n2669), .ZN(n2716) );
  AOI211_X1 U3423 ( .C1(n4510), .C2(n3684), .A(n2670), .B(n2716), .ZN(n4500)
         );
  NAND2_X1 U3424 ( .A1(n2672), .A2(n2671), .ZN(n2677) );
  OAI21_X1 U3425 ( .B1(n2674), .B2(D_REG_1__SCAN_IN), .A(n2673), .ZN(n2675) );
  NAND4_X1 U3426 ( .A1(n2678), .A2(n2677), .A3(n2676), .A4(n2675), .ZN(n2935)
         );
  NAND2_X1 U3427 ( .A1(n4545), .A2(REG1_REG_0__SCAN_IN), .ZN(n2680) );
  OAI21_X1 U3428 ( .B1(n4500), .B2(n4545), .A(n2680), .ZN(U3518) );
  NAND2_X1 U3429 ( .A1(n2683), .A2(IR_REG_31__SCAN_IN), .ZN(n2682) );
  MUX2_X1 U3430 ( .A(n2682), .B(IR_REG_31__SCAN_IN), .S(n2684), .Z(n2686) );
  NAND2_X1 U3431 ( .A1(n2686), .A2(n3154), .ZN(n3825) );
  INV_X1 U3432 ( .A(IR_REG_7__SCAN_IN), .ZN(n2688) );
  NAND2_X1 U3433 ( .A1(n2689), .A2(n2688), .ZN(n2690) );
  NAND2_X1 U3434 ( .A1(n2690), .A2(IR_REG_31__SCAN_IN), .ZN(n2692) );
  INV_X1 U3435 ( .A(IR_REG_8__SCAN_IN), .ZN(n2691) );
  XNOR2_X1 U3436 ( .A(n2692), .B(n2691), .ZN(n4499) );
  OR2_X1 U3437 ( .A1(n2693), .A2(n4499), .ZN(n2694) );
  INV_X1 U3438 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3003) );
  MUX2_X1 U3439 ( .A(n3003), .B(REG2_REG_9__SCAN_IN), .S(n3825), .Z(n2695) );
  NAND2_X1 U3440 ( .A1(n2696), .A2(n2695), .ZN(n3824) );
  OAI211_X1 U3441 ( .C1(n2696), .C2(n2695), .A(n3824), .B(n4472), .ZN(n2710)
         );
  INV_X1 U3442 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2697) );
  NOR2_X1 U3443 ( .A1(STATE_REG_SCAN_IN), .A2(n2697), .ZN(n3550) );
  INV_X1 U3444 ( .A(n4352), .ZN(n2698) );
  INV_X1 U3445 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4367) );
  NAND2_X1 U3446 ( .A1(n2702), .A2(n4499), .ZN(n2703) );
  NOR2_X1 U3447 ( .A1(n4367), .A2(n4366), .ZN(n4365) );
  NOR2_X1 U3448 ( .A1(n2704), .A2(n4365), .ZN(n2707) );
  INV_X1 U3449 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2705) );
  MUX2_X1 U3450 ( .A(REG1_REG_9__SCAN_IN), .B(n2705), .S(n3825), .Z(n2706) );
  NOR2_X1 U3451 ( .A1(n2707), .A2(n2706), .ZN(n3809) );
  AOI211_X1 U3452 ( .C1(n2707), .C2(n2706), .A(n3809), .B(n4460), .ZN(n2708)
         );
  AOI211_X1 U3453 ( .C1(n4464), .C2(ADDR_REG_9__SCAN_IN), .A(n3550), .B(n2708), 
        .ZN(n2709) );
  OAI211_X1 U3454 ( .C1(n4475), .C2(n3825), .A(n2710), .B(n2709), .ZN(U3249)
         );
  INV_X1 U3455 ( .A(n4510), .ZN(n4540) );
  OAI22_X1 U3456 ( .A1(n2712), .A2(n4540), .B1(n4503), .B2(n2711), .ZN(n2713)
         );
  NOR2_X1 U3457 ( .A1(n2714), .A2(n2713), .ZN(n4501) );
  NAND2_X1 U34580 ( .A1(n4545), .A2(REG1_REG_1__SCAN_IN), .ZN(n2715) );
  OAI21_X1 U34590 ( .B1(n4501), .B2(n4545), .A(n2715), .ZN(U3519) );
  OAI21_X1 U3460 ( .B1(n4350), .B2(n2235), .A(n4127), .ZN(n2717) );
  AOI21_X1 U3461 ( .B1(n2577), .B2(n2717), .A(n2716), .ZN(n2722) );
  INV_X1 U3462 ( .A(n4099), .ZN(n4480) );
  INV_X2 U3463 ( .A(n4477), .ZN(n4198) );
  OAI22_X1 U3464 ( .A1(n4198), .A2(n2719), .B1(n2718), .B2(n4196), .ZN(n2720)
         );
  AOI21_X1 U3465 ( .B1(n4480), .B2(n3684), .A(n2720), .ZN(n2721) );
  OAI21_X1 U3466 ( .B1(n2722), .B2(n4477), .A(n2721), .ZN(U3290) );
  MUX2_X1 U34670 ( .A(n2723), .B(DATAI_2_), .S(n3349), .Z(n2938) );
  INV_X1 U3468 ( .A(n2938), .ZN(n2761) );
  OAI22_X1 U34690 ( .A1(n2764), .A2(n3445), .B1(n2649), .B2(n2761), .ZN(n2743)
         );
  XNOR2_X1 U3470 ( .A(n2742), .B(n2743), .ZN(n2733) );
  INV_X1 U34710 ( .A(n2725), .ZN(n2727) );
  NAND2_X1 U3472 ( .A1(n2727), .A2(n2726), .ZN(n2728) );
  NAND2_X1 U34730 ( .A1(n2729), .A2(n2728), .ZN(n2730) );
  INV_X1 U3474 ( .A(n2733), .ZN(n2731) );
  INV_X1 U34750 ( .A(n2747), .ZN(n2732) );
  AOI21_X1 U3476 ( .B1(n2733), .B2(n2730), .A(n2732), .ZN(n2738) );
  OAI22_X1 U34770 ( .A1(n2928), .A2(n3626), .B1(n2651), .B2(n3623), .ZN(n2736)
         );
  NOR2_X1 U3478 ( .A1(n2734), .A2(n2376), .ZN(n2735) );
  AOI211_X1 U34790 ( .C1(n2938), .C2(n3588), .A(n2736), .B(n2735), .ZN(n2737)
         );
  OAI21_X1 U3480 ( .B1(n2738), .B2(n3616), .A(n2737), .ZN(U3234) );
  MUX2_X1 U34810 ( .A(n4355), .B(DATAI_3_), .S(n3349), .Z(n2799) );
  AOI22_X1 U3482 ( .A1(n2800), .A2(n3422), .B1(n2799), .B2(n3416), .ZN(n2776)
         );
  NAND2_X1 U34830 ( .A1(n2800), .A2(n3416), .ZN(n2740) );
  NAND2_X1 U3484 ( .A1(n2799), .A2(n3417), .ZN(n2739) );
  NAND2_X1 U34850 ( .A1(n2740), .A2(n2739), .ZN(n2741) );
  INV_X1 U3486 ( .A(n2742), .ZN(n2745) );
  INV_X1 U34870 ( .A(n2743), .ZN(n2744) );
  NAND2_X1 U3488 ( .A1(n2745), .A2(n2744), .ZN(n2746) );
  XOR2_X1 U34890 ( .A(n2773), .B(n2774), .Z(n2759) );
  OAI22_X1 U3490 ( .A1(n2764), .A2(n3623), .B1(n2865), .B2(n3626), .ZN(n2757)
         );
  INV_X1 U34910 ( .A(n2748), .ZN(n2749) );
  NOR2_X1 U3492 ( .A1(n2750), .A2(n2749), .ZN(n2751) );
  AND2_X1 U34930 ( .A1(n2576), .A2(n2751), .ZN(n2752) );
  AOI21_X1 U3494 ( .B1(n2753), .B2(n2752), .A(U3149), .ZN(n2755) );
  MUX2_X1 U34950 ( .A(n3614), .B(U3149), .S(REG3_REG_3__SCAN_IN), .Z(n2756) );
  AOI211_X1 U3496 ( .C1(n2799), .C2(n3588), .A(n2757), .B(n2756), .ZN(n2758)
         );
  OAI21_X1 U34970 ( .B1(n2759), .B2(n3616), .A(n2758), .ZN(U3215) );
  NAND2_X1 U3498 ( .A1(n2926), .A2(n2760), .ZN(n2847) );
  NAND2_X1 U34990 ( .A1(n2850), .A2(n2847), .ZN(n2923) );
  INV_X1 U3500 ( .A(n2764), .ZN(n3782) );
  NAND2_X1 U35010 ( .A1(n3782), .A2(n2761), .ZN(n3709) );
  AND2_X2 U3502 ( .A1(n3709), .A2(n3706), .ZN(n2849) );
  NAND2_X1 U35030 ( .A1(n2764), .A2(n2761), .ZN(n2797) );
  NAND2_X1 U3504 ( .A1(n2921), .A2(n2797), .ZN(n2762) );
  NAND2_X1 U35050 ( .A1(n2928), .A2(n2799), .ZN(n3711) );
  NAND2_X1 U35060 ( .A1(n2800), .A2(n2793), .ZN(n3708) );
  AND2_X2 U35070 ( .A1(n3711), .A2(n3708), .ZN(n3670) );
  XNOR2_X1 U35080 ( .A(n2762), .B(n3670), .ZN(n4504) );
  OAI21_X2 U35090 ( .B1(n2362), .B2(n3700), .A(n3705), .ZN(n2925) );
  NAND2_X1 U35100 ( .A1(n2925), .A2(n2849), .ZN(n2924) );
  NAND2_X1 U35110 ( .A1(n2924), .A2(n3706), .ZN(n2810) );
  XNOR2_X1 U35120 ( .A(n2810), .B(n3670), .ZN(n2766) );
  AOI22_X1 U35130 ( .A1(n2798), .A2(n4187), .B1(n4216), .B2(n2799), .ZN(n2763)
         );
  OAI21_X1 U35140 ( .B1(n2764), .B2(n4191), .A(n2763), .ZN(n2765) );
  AOI21_X1 U35150 ( .B1(n2766), .B2(n4184), .A(n2765), .ZN(n2767) );
  OAI21_X1 U35160 ( .B1(n4504), .B2(n4089), .A(n2767), .ZN(n4506) );
  NAND2_X1 U35170 ( .A1(n4506), .A2(n4198), .ZN(n2772) );
  OAI21_X1 U35180 ( .B1(n2936), .B2(n2793), .A(n2817), .ZN(n4502) );
  INV_X1 U35190 ( .A(n4502), .ZN(n2770) );
  OAI22_X1 U35200 ( .A1(n4198), .A2(n2768), .B1(REG3_REG_3__SCAN_IN), .B2(
        n4196), .ZN(n2769) );
  AOI21_X1 U35210 ( .B1(n2770), .B2(n4479), .A(n2769), .ZN(n2771) );
  OAI211_X1 U35220 ( .C1(n4504), .C2(n4099), .A(n2772), .B(n2771), .ZN(U3287)
         );
  INV_X1 U35230 ( .A(n2775), .ZN(n2777) );
  NAND2_X1 U35240 ( .A1(n2777), .A2(n2776), .ZN(n2778) );
  MUX2_X1 U35250 ( .A(n4354), .B(DATAI_4_), .S(n3349), .Z(n2854) );
  INV_X1 U35260 ( .A(n2854), .ZN(n2819) );
  OAI22_X1 U35270 ( .A1(n2865), .A2(n3373), .B1(n3448), .B2(n2819), .ZN(n2780)
         );
  XNOR2_X1 U35280 ( .A(n2780), .B(n3446), .ZN(n2826) );
  OAI22_X1 U35290 ( .A1(n2865), .A2(n3445), .B1(n3373), .B2(n2819), .ZN(n2825)
         );
  XNOR2_X1 U35300 ( .A(n2826), .B(n2825), .ZN(n2781) );
  AOI21_X1 U35310 ( .B1(n2782), .B2(n2781), .A(n3616), .ZN(n2783) );
  NAND2_X1 U35320 ( .A1(n2783), .A2(n2828), .ZN(n2789) );
  INV_X1 U35330 ( .A(n3623), .ZN(n3586) );
  NAND2_X1 U35340 ( .A1(n3586), .A2(n2800), .ZN(n2784) );
  OAI21_X1 U35350 ( .B1(n3624), .B2(n2819), .A(n2784), .ZN(n2787) );
  OAI21_X1 U35360 ( .B1(n2955), .B2(n3626), .A(n2785), .ZN(n2786) );
  NOR2_X1 U35370 ( .A1(n2787), .A2(n2786), .ZN(n2788) );
  OAI211_X1 U35380 ( .C1(n3631), .C2(n2820), .A(n2789), .B(n2788), .ZN(U3227)
         );
  NAND4_X1 U35390 ( .A1(n2795), .A2(n2794), .A3(n2793), .A4(n2792), .ZN(n2796)
         );
  AND2_X1 U35400 ( .A1(n2797), .A2(n2796), .ZN(n2803) );
  NAND2_X1 U35410 ( .A1(n2798), .A2(n2819), .ZN(n2862) );
  NAND2_X1 U35420 ( .A1(n2865), .A2(n2854), .ZN(n2859) );
  INV_X1 U35430 ( .A(n2801), .ZN(n2806) );
  NAND2_X1 U35440 ( .A1(n2921), .A2(n2852), .ZN(n2802) );
  NAND2_X1 U35450 ( .A1(n2800), .A2(n2799), .ZN(n2805) );
  AND2_X1 U35460 ( .A1(n2802), .A2(n2856), .ZN(n2809) );
  NAND2_X1 U35470 ( .A1(n2921), .A2(n2803), .ZN(n2804) );
  AND2_X1 U35480 ( .A1(n2805), .A2(n2804), .ZN(n2807) );
  NAND2_X1 U35490 ( .A1(n2807), .A2(n2801), .ZN(n2808) );
  INV_X1 U35500 ( .A(n4511), .ZN(n2824) );
  INV_X1 U35510 ( .A(n4184), .ZN(n4025) );
  NAND2_X1 U35520 ( .A1(n2810), .A2(n3670), .ZN(n2811) );
  XOR2_X1 U35530 ( .A(n2801), .B(n2861), .Z(n2816) );
  AOI22_X1 U35540 ( .A1(n2800), .A2(n3210), .B1(n4216), .B2(n2854), .ZN(n2812)
         );
  OAI21_X1 U35550 ( .B1(n2955), .B2(n4128), .A(n2812), .ZN(n2813) );
  AOI21_X1 U35560 ( .B1(n4511), .B2(n2814), .A(n2813), .ZN(n2815) );
  OAI21_X1 U35570 ( .B1(n4025), .B2(n2816), .A(n2815), .ZN(n4508) );
  OAI211_X1 U35580 ( .C1(n2818), .C2(n2819), .A(n4536), .B(n2868), .ZN(n4507)
         );
  OAI22_X1 U35590 ( .A1(n4507), .A2(n4350), .B1(n4196), .B2(n2820), .ZN(n2821)
         );
  OAI21_X1 U35600 ( .B1(n4508), .B2(n2821), .A(n4198), .ZN(n2823) );
  NAND2_X1 U35610 ( .A1(n4477), .A2(REG2_REG_4__SCAN_IN), .ZN(n2822) );
  OAI211_X1 U35620 ( .C1(n2824), .C2(n4099), .A(n2823), .B(n2822), .ZN(U3286)
         );
  NAND2_X1 U35630 ( .A1(n2826), .A2(n2825), .ZN(n2827) );
  MUX2_X1 U35640 ( .A(n2829), .B(n2427), .S(n3349), .Z(n2884) );
  OAI22_X1 U35650 ( .A1(n2955), .A2(n3373), .B1(n3448), .B2(n2884), .ZN(n2830)
         );
  XNOR2_X1 U35660 ( .A(n2830), .B(n3434), .ZN(n2942) );
  OAI22_X1 U35670 ( .A1(n2955), .A2(n3445), .B1(n3373), .B2(n2884), .ZN(n2943)
         );
  XNOR2_X1 U35680 ( .A(n2942), .B(n2943), .ZN(n2831) );
  OAI211_X1 U35690 ( .C1(n2832), .C2(n2831), .A(n2946), .B(n3621), .ZN(n2844)
         );
  NAND2_X1 U35700 ( .A1(n2798), .A2(n3586), .ZN(n2841) );
  OAI21_X1 U35710 ( .B1(n2833), .B2(REG3_REG_6__SCAN_IN), .A(n2902), .ZN(n2963) );
  OR2_X1 U35720 ( .A1(n3459), .A2(n2963), .ZN(n2838) );
  INV_X1 U35730 ( .A(REG0_REG_6__SCAN_IN), .ZN(n2834) );
  OR2_X1 U35740 ( .A1(n3634), .A2(n2834), .ZN(n2837) );
  NAND2_X1 U35750 ( .A1(n3297), .A2(REG1_REG_6__SCAN_IN), .ZN(n2835) );
  NAND4_X1 U35760 ( .A1(n2838), .A2(n2837), .A3(n2836), .A4(n2835), .ZN(n3781)
         );
  AOI21_X1 U35770 ( .B1(n3583), .B2(n3781), .A(n2839), .ZN(n2840) );
  OAI211_X1 U35780 ( .C1(n3624), .C2(n2884), .A(n2841), .B(n2840), .ZN(n2842)
         );
  INV_X1 U35790 ( .A(n2842), .ZN(n2843) );
  OAI211_X1 U35800 ( .C1(n3631), .C2(n2870), .A(n2844), .B(n2843), .ZN(U3224)
         );
  AND2_X1 U35810 ( .A1(n4089), .A2(n2845), .ZN(n2846) );
  INV_X1 U3582 ( .A(n2847), .ZN(n2848) );
  NOR2_X1 U3583 ( .A1(n2849), .A2(n2848), .ZN(n2851) );
  NAND2_X1 U3584 ( .A1(n2851), .A2(n2850), .ZN(n2853) );
  NAND2_X1 U3585 ( .A1(n2853), .A2(n2852), .ZN(n2858) );
  NAND2_X1 U3586 ( .A1(n2798), .A2(n2854), .ZN(n2855) );
  NAND2_X1 U3587 ( .A1(n2858), .A2(n2857), .ZN(n2886) );
  AND2_X1 U3588 ( .A1(n2888), .A2(n2884), .ZN(n2874) );
  INV_X1 U3589 ( .A(n2874), .ZN(n3713) );
  NAND2_X1 U3590 ( .A1(n2955), .A2(n2887), .ZN(n3723) );
  NAND2_X1 U3591 ( .A1(n3713), .A2(n3723), .ZN(n3689) );
  XNOR2_X1 U3592 ( .A(n2886), .B(n3689), .ZN(n4513) );
  INV_X1 U3593 ( .A(n2859), .ZN(n2860) );
  NAND2_X1 U3594 ( .A1(n2863), .A2(n2862), .ZN(n2875) );
  XNOR2_X1 U3595 ( .A(n2875), .B(n3689), .ZN(n2867) );
  AOI22_X1 U3596 ( .A1(n3781), .A2(n4187), .B1(n4216), .B2(n2887), .ZN(n2864)
         );
  OAI21_X1 U3597 ( .B1(n2865), .B2(n4191), .A(n2864), .ZN(n2866) );
  AOI21_X1 U3598 ( .B1(n2867), .B2(n4184), .A(n2866), .ZN(n4514) );
  MUX2_X1 U3599 ( .A(n4514), .B(n4693), .S(n4477), .Z(n2873) );
  AND2_X1 U3600 ( .A1(n2868), .A2(n2887), .ZN(n2869) );
  NOR2_X1 U3601 ( .A1(n2894), .A2(n2869), .ZN(n4517) );
  INV_X1 U3602 ( .A(n2870), .ZN(n2871) );
  INV_X1 U3603 ( .A(n4196), .ZN(n4476) );
  AOI22_X1 U3604 ( .A1(n4517), .A2(n4479), .B1(n2871), .B2(n4476), .ZN(n2872)
         );
  OAI211_X1 U3605 ( .C1(n4202), .C2(n4513), .A(n2873), .B(n2872), .ZN(U3285)
         );
  OAI21_X2 U3606 ( .B1(n2875), .B2(n2874), .A(n3723), .ZN(n2899) );
  INV_X1 U3607 ( .A(n3781), .ZN(n2876) );
  MUX2_X1 U3608 ( .A(n4353), .B(DATAI_6_), .S(n3349), .Z(n2950) );
  NAND2_X1 U3609 ( .A1(n2876), .A2(n2950), .ZN(n3715) );
  NAND2_X1 U3610 ( .A1(n3781), .A2(n2956), .ZN(n3725) );
  AND2_X1 U3611 ( .A1(n3715), .A2(n3725), .ZN(n3673) );
  XNOR2_X1 U3612 ( .A(n2899), .B(n3673), .ZN(n2893) );
  NAND2_X1 U3613 ( .A1(n3297), .A2(REG1_REG_7__SCAN_IN), .ZN(n2881) );
  INV_X1 U3614 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2877) );
  XNOR2_X1 U3615 ( .A(n2902), .B(n2877), .ZN(n2994) );
  OR2_X1 U3616 ( .A1(n2536), .A2(n2994), .ZN(n2880) );
  INV_X1 U3617 ( .A(REG0_REG_7__SCAN_IN), .ZN(n2878) );
  OR2_X1 U3618 ( .A1(n3634), .A2(n2878), .ZN(n2879) );
  AOI22_X1 U3619 ( .A1(n3780), .A2(n4187), .B1(n4216), .B2(n2950), .ZN(n2883)
         );
  OAI21_X1 U3620 ( .B1(n2955), .B2(n4191), .A(n2883), .ZN(n2892) );
  NAND2_X1 U3621 ( .A1(n2955), .A2(n2884), .ZN(n2885) );
  NAND2_X1 U3622 ( .A1(n2886), .A2(n2885), .ZN(n2890) );
  NAND2_X1 U3623 ( .A1(n2888), .A2(n2887), .ZN(n2889) );
  NAND2_X1 U3624 ( .A1(n2890), .A2(n2889), .ZN(n2918) );
  XOR2_X1 U3625 ( .A(n2918), .B(n3673), .Z(n4541) );
  NOR2_X1 U3626 ( .A1(n4541), .A2(n4089), .ZN(n2891) );
  AOI211_X1 U3627 ( .C1(n2893), .C2(n4184), .A(n2892), .B(n2891), .ZN(n4539)
         );
  INV_X1 U3628 ( .A(n2894), .ZN(n2895) );
  AOI21_X1 U3629 ( .B1(n2950), .B2(n2895), .A(n2170), .ZN(n4537) );
  OAI22_X1 U3630 ( .A1(n4198), .A2(n2190), .B1(n2963), .B2(n4196), .ZN(n2897)
         );
  NOR2_X1 U3631 ( .A1(n4541), .A2(n4099), .ZN(n2896) );
  AOI211_X1 U3632 ( .C1(n4479), .C2(n4537), .A(n2897), .B(n2896), .ZN(n2898)
         );
  OAI21_X1 U3633 ( .B1(n4539), .B2(n4477), .A(n2898), .ZN(U3284) );
  NAND2_X1 U3634 ( .A1(n2899), .A2(n3725), .ZN(n2900) );
  NAND2_X1 U3635 ( .A1(n2900), .A2(n3715), .ZN(n2966) );
  MUX2_X1 U3636 ( .A(n4352), .B(DATAI_7_), .S(n3349), .Z(n2971) );
  NAND2_X1 U3637 ( .A1(n3028), .A2(n2971), .ZN(n2964) );
  XNOR2_X1 U3638 ( .A(n2966), .B(n3716), .ZN(n2913) );
  NAND2_X1 U3639 ( .A1(n3297), .A2(REG1_REG_8__SCAN_IN), .ZN(n2909) );
  INV_X1 U3640 ( .A(REG0_REG_8__SCAN_IN), .ZN(n2901) );
  OR2_X1 U3641 ( .A1(n3634), .A2(n2901), .ZN(n2907) );
  INV_X1 U3642 ( .A(n2902), .ZN(n2903) );
  AOI21_X1 U3643 ( .B1(n2903), .B2(REG3_REG_7__SCAN_IN), .A(
        REG3_REG_8__SCAN_IN), .ZN(n2905) );
  OR2_X1 U3644 ( .A1(n2905), .A2(n2904), .ZN(n3033) );
  OR2_X1 U3645 ( .A1(n2536), .A2(n3033), .ZN(n2906) );
  NAND2_X1 U3646 ( .A1(n2971), .A2(n4216), .ZN(n2911) );
  NAND2_X1 U3647 ( .A1(n3781), .A2(n3210), .ZN(n2910) );
  OAI211_X1 U3648 ( .C1(n3018), .C2(n4128), .A(n2911), .B(n2910), .ZN(n2912)
         );
  AOI21_X1 U3649 ( .B1(n2913), .B2(n4184), .A(n2912), .ZN(n4524) );
  OAI211_X1 U3650 ( .C1(n2170), .C2(n2990), .A(n4536), .B(n2973), .ZN(n4521)
         );
  INV_X1 U3651 ( .A(n4521), .ZN(n2916) );
  INV_X1 U3652 ( .A(n4137), .ZN(n2915) );
  OAI22_X1 U3653 ( .A1(n4198), .A2(n4821), .B1(n2994), .B2(n4196), .ZN(n2914)
         );
  AOI21_X1 U3654 ( .B1(n2916), .B2(n2915), .A(n2914), .ZN(n2920) );
  AND2_X1 U3655 ( .A1(n3781), .A2(n2950), .ZN(n2917) );
  OAI22_X1 U3656 ( .A1(n2918), .A2(n2917), .B1(n2950), .B2(n3781), .ZN(n3084)
         );
  OR2_X1 U3657 ( .A1(n3084), .A2(n3716), .ZN(n4520) );
  NAND2_X1 U3658 ( .A1(n3084), .A2(n3716), .ZN(n4519) );
  NAND3_X1 U3659 ( .A1(n4520), .A2(n4519), .A3(n3953), .ZN(n2919) );
  OAI211_X1 U3660 ( .C1(n4524), .C2(n4477), .A(n2920), .B(n2919), .ZN(U3283)
         );
  INV_X1 U3661 ( .A(n2921), .ZN(n2922) );
  AOI21_X1 U3662 ( .B1(n2849), .B2(n2923), .A(n2922), .ZN(n2929) );
  INV_X1 U3663 ( .A(n2929), .ZN(n4481) );
  OAI21_X1 U3664 ( .B1(n2849), .B2(n2925), .A(n2924), .ZN(n2932) );
  AOI22_X1 U3665 ( .A1(n2926), .A2(n3210), .B1(n4216), .B2(n2938), .ZN(n2927)
         );
  OAI21_X1 U3666 ( .B1(n2928), .B2(n4128), .A(n2927), .ZN(n2931) );
  NOR2_X1 U3667 ( .A1(n2929), .A2(n4089), .ZN(n2930) );
  AOI211_X1 U3668 ( .C1(n4184), .C2(n2932), .A(n2931), .B(n2930), .ZN(n4484)
         );
  INV_X1 U3669 ( .A(n4484), .ZN(n2933) );
  AOI21_X1 U3670 ( .B1(n4510), .B2(n4481), .A(n2933), .ZN(n2941) );
  AOI21_X1 U3671 ( .B1(n2938), .B2(n2937), .A(n2936), .ZN(n4478) );
  INV_X2 U3672 ( .A(n4790), .ZN(n4518) );
  AND2_X1 U3673 ( .A1(n4518), .A2(n4536), .ZN(n4307) );
  AOI22_X1 U3674 ( .A1(n4478), .A2(n4307), .B1(n4790), .B2(REG0_REG_2__SCAN_IN), .ZN(n2939) );
  OAI21_X1 U3675 ( .B1(n2941), .B2(n4790), .A(n2939), .ZN(U3471) );
  AOI22_X1 U3676 ( .A1(n4478), .A2(n4242), .B1(REG1_REG_2__SCAN_IN), .B2(n4545), .ZN(n2940) );
  OAI21_X1 U3677 ( .B1(n2941), .B2(n4545), .A(n2940), .ZN(U3520) );
  INV_X1 U3678 ( .A(n2942), .ZN(n2944) );
  NAND2_X1 U3679 ( .A1(n2944), .A2(n2943), .ZN(n2945) );
  NAND2_X1 U3680 ( .A1(n3781), .A2(n3416), .ZN(n2948) );
  NAND2_X1 U3681 ( .A1(n2950), .A2(n3417), .ZN(n2947) );
  NAND2_X1 U3682 ( .A1(n2948), .A2(n2947), .ZN(n2949) );
  XNOR2_X1 U3683 ( .A(n2949), .B(n3446), .ZN(n2980) );
  NAND2_X1 U3684 ( .A1(n3781), .A2(n3422), .ZN(n2952) );
  NAND2_X1 U3685 ( .A1(n2950), .A2(n3416), .ZN(n2951) );
  NAND2_X1 U3686 ( .A1(n2952), .A2(n2951), .ZN(n2981) );
  XNOR2_X1 U3687 ( .A(n2980), .B(n2981), .ZN(n2953) );
  XNOR2_X1 U3688 ( .A(n2982), .B(n2953), .ZN(n2954) );
  NAND2_X1 U3689 ( .A1(n2954), .A2(n3621), .ZN(n2962) );
  OAI22_X1 U3690 ( .A1(n3624), .A2(n2956), .B1(n2955), .B2(n3623), .ZN(n2960)
         );
  INV_X1 U3691 ( .A(n2957), .ZN(n2958) );
  OAI21_X1 U3692 ( .B1(n3028), .B2(n3626), .A(n2958), .ZN(n2959) );
  NOR2_X1 U3693 ( .A1(n2960), .A2(n2959), .ZN(n2961) );
  OAI211_X1 U3694 ( .C1(n3631), .C2(n2963), .A(n2962), .B(n2961), .ZN(U3236)
         );
  INV_X1 U3695 ( .A(n2964), .ZN(n2965) );
  OAI21_X2 U3696 ( .B1(n2966), .B2(n2965), .A(n3722), .ZN(n2995) );
  INV_X1 U3697 ( .A(DATAI_8_), .ZN(n2967) );
  MUX2_X1 U3698 ( .A(n4499), .B(n2967), .S(n3349), .Z(n3027) );
  NAND2_X1 U3699 ( .A1(n3018), .A2(n3005), .ZN(n3720) );
  NAND2_X1 U3700 ( .A1(n3779), .A2(n3027), .ZN(n3726) );
  AND2_X1 U3701 ( .A1(n3720), .A2(n3726), .ZN(n3669) );
  XNOR2_X1 U3702 ( .A(n2995), .B(n3669), .ZN(n2970) );
  INV_X1 U3703 ( .A(n3088), .ZN(n3086) );
  OAI22_X1 U3704 ( .A1(n3086), .A2(n4128), .B1(n4127), .B2(n3027), .ZN(n2968)
         );
  AOI21_X1 U3705 ( .B1(n3210), .B2(n3780), .A(n2968), .ZN(n2969) );
  OAI21_X1 U3706 ( .B1(n2970), .B2(n4025), .A(n2969), .ZN(n3034) );
  INV_X1 U3707 ( .A(n3034), .ZN(n2979) );
  NAND2_X1 U3708 ( .A1(n3780), .A2(n2971), .ZN(n3007) );
  NAND2_X1 U3709 ( .A1(n4520), .A2(n3007), .ZN(n2972) );
  XNOR2_X1 U3710 ( .A(n2972), .B(n3669), .ZN(n3035) );
  INV_X1 U3711 ( .A(n2973), .ZN(n2974) );
  OAI21_X1 U3712 ( .B1(n2974), .B2(n3027), .A(n3001), .ZN(n3039) );
  NOR2_X1 U3713 ( .A1(n3039), .A2(n4195), .ZN(n2977) );
  INV_X1 U3714 ( .A(REG2_REG_8__SCAN_IN), .ZN(n2975) );
  OAI22_X1 U3715 ( .A1(n4198), .A2(n2975), .B1(n3033), .B2(n4196), .ZN(n2976)
         );
  AOI211_X1 U3716 ( .C1(n3035), .C2(n3953), .A(n2977), .B(n2976), .ZN(n2978)
         );
  OAI21_X1 U3717 ( .B1(n2979), .B2(n4477), .A(n2978), .ZN(U3282) );
  NAND2_X1 U3718 ( .A1(n2982), .A2(n2981), .ZN(n2983) );
  NAND2_X1 U3719 ( .A1(n2984), .A2(n2983), .ZN(n3061) );
  OAI22_X1 U3720 ( .A1(n3028), .A2(n3373), .B1(n3448), .B2(n2990), .ZN(n2985)
         );
  XNOR2_X1 U3721 ( .A(n2985), .B(n3434), .ZN(n3014) );
  OAI22_X1 U3722 ( .A1(n3028), .A2(n3445), .B1(n3373), .B2(n2990), .ZN(n3015)
         );
  XNOR2_X1 U3723 ( .A(n3014), .B(n3015), .ZN(n3059) );
  XOR2_X1 U3724 ( .A(n3061), .B(n3059), .Z(n2986) );
  NAND2_X1 U3725 ( .A1(n2986), .A2(n3621), .ZN(n2993) );
  NAND2_X1 U3726 ( .A1(n3779), .A2(n3583), .ZN(n2989) );
  AOI21_X1 U3727 ( .B1(n3586), .B2(n3781), .A(n2987), .ZN(n2988) );
  OAI211_X1 U3728 ( .C1(n3624), .C2(n2990), .A(n2989), .B(n2988), .ZN(n2991)
         );
  INV_X1 U3729 ( .A(n2991), .ZN(n2992) );
  OAI211_X1 U3730 ( .C1(n3631), .C2(n2994), .A(n2993), .B(n2992), .ZN(U3210)
         );
  NAND2_X1 U3731 ( .A1(n2995), .A2(n3720), .ZN(n2996) );
  NAND2_X1 U3732 ( .A1(n2996), .A2(n3726), .ZN(n3072) );
  INV_X1 U3733 ( .A(n3825), .ZN(n4351) );
  MUX2_X1 U3734 ( .A(n4351), .B(DATAI_9_), .S(n3349), .Z(n3551) );
  INV_X1 U3735 ( .A(n3551), .ZN(n3085) );
  AND2_X1 U3736 ( .A1(n3088), .A2(n3085), .ZN(n3731) );
  INV_X1 U3737 ( .A(n3731), .ZN(n3727) );
  NAND2_X1 U3738 ( .A1(n3086), .A2(n3551), .ZN(n3719) );
  AND2_X1 U3739 ( .A1(n3727), .A2(n3719), .ZN(n3671) );
  INV_X1 U3740 ( .A(n3671), .ZN(n2997) );
  XNOR2_X1 U3741 ( .A(n3072), .B(n2997), .ZN(n3000) );
  AOI22_X1 U3742 ( .A1(n3585), .A2(n4187), .B1(n4216), .B2(n3551), .ZN(n2998)
         );
  OAI21_X1 U3743 ( .B1(n3018), .B2(n4191), .A(n2998), .ZN(n2999) );
  AOI21_X1 U3744 ( .B1(n3000), .B2(n4184), .A(n2999), .ZN(n4530) );
  AND2_X1 U3745 ( .A1(n3001), .A2(n3551), .ZN(n3002) );
  NOR2_X1 U3746 ( .A1(n3080), .A2(n3002), .ZN(n4527) );
  OAI22_X1 U3747 ( .A1(n4198), .A2(n3003), .B1(n3552), .B2(n4196), .ZN(n3004)
         );
  AOI21_X1 U3748 ( .B1(n4527), .B2(n4479), .A(n3004), .ZN(n3013) );
  AND2_X1 U3749 ( .A1(n3018), .A2(n3027), .ZN(n3009) );
  OR2_X1 U3750 ( .A1(n3084), .A2(n3087), .ZN(n3010) );
  NAND2_X1 U3751 ( .A1(n3779), .A2(n3005), .ZN(n3006) );
  AND2_X1 U3752 ( .A1(n3007), .A2(n3006), .ZN(n3008) );
  OR2_X1 U3753 ( .A1(n3009), .A2(n3008), .ZN(n3089) );
  NAND2_X1 U3754 ( .A1(n3010), .A2(n3089), .ZN(n3011) );
  XNOR2_X1 U3755 ( .A(n3011), .B(n3671), .ZN(n4526) );
  NAND2_X1 U3756 ( .A1(n4526), .A2(n3953), .ZN(n3012) );
  OAI211_X1 U3757 ( .C1(n4530), .C2(n4477), .A(n3013), .B(n3012), .ZN(U3281)
         );
  NAND2_X1 U3758 ( .A1(n3061), .A2(n3059), .ZN(n3544) );
  INV_X1 U3759 ( .A(n3014), .ZN(n3016) );
  NAND2_X1 U3760 ( .A1(n3016), .A2(n3015), .ZN(n3046) );
  NAND2_X1 U3761 ( .A1(n3544), .A2(n3046), .ZN(n3024) );
  OAI22_X1 U3762 ( .A1(n3018), .A2(n3373), .B1(n3448), .B2(n3027), .ZN(n3017)
         );
  XNOR2_X1 U3763 ( .A(n3017), .B(n3446), .ZN(n3019) );
  OAI22_X1 U3764 ( .A1(n3018), .A2(n3445), .B1(n3373), .B2(n3027), .ZN(n3020)
         );
  INV_X1 U3765 ( .A(n3019), .ZN(n3022) );
  INV_X1 U3766 ( .A(n3020), .ZN(n3021) );
  NAND2_X1 U3767 ( .A1(n3022), .A2(n3021), .ZN(n3545) );
  NAND2_X1 U3768 ( .A1(n2307), .A2(n3545), .ZN(n3023) );
  XNOR2_X1 U3769 ( .A(n3024), .B(n3023), .ZN(n3025) );
  NAND2_X1 U3770 ( .A1(n3025), .A2(n3621), .ZN(n3032) );
  NAND2_X1 U3771 ( .A1(n3583), .A2(n3088), .ZN(n3026) );
  OAI21_X1 U3772 ( .B1(n3624), .B2(n3027), .A(n3026), .ZN(n3030) );
  NAND2_X1 U3773 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n4364) );
  OAI21_X1 U3774 ( .B1(n3028), .B2(n3623), .A(n4364), .ZN(n3029) );
  NOR2_X1 U3775 ( .A1(n3030), .A2(n3029), .ZN(n3031) );
  OAI211_X1 U3776 ( .C1(n3631), .C2(n3033), .A(n3032), .B(n3031), .ZN(U3218)
         );
  AOI21_X1 U3777 ( .B1(n3035), .B2(n4525), .A(n3034), .ZN(n3037) );
  MUX2_X1 U3778 ( .A(n2901), .B(n3037), .S(n4518), .Z(n3036) );
  OAI21_X1 U3779 ( .B1(n3039), .B2(n4342), .A(n3036), .ZN(U3483) );
  MUX2_X1 U3780 ( .A(n4367), .B(n3037), .S(n4547), .Z(n3038) );
  OAI21_X1 U3781 ( .B1(n3039), .B2(n4286), .A(n3038), .ZN(U3526) );
  INV_X1 U3782 ( .A(n3081), .ZN(n3070) );
  NAND2_X1 U3783 ( .A1(n3154), .A2(IR_REG_31__SCAN_IN), .ZN(n3040) );
  XNOR2_X1 U3784 ( .A(n3040), .B(IR_REG_10__SCAN_IN), .ZN(n3826) );
  MUX2_X1 U3785 ( .A(n3826), .B(DATAI_10_), .S(n3349), .Z(n3136) );
  NAND2_X1 U3786 ( .A1(n3130), .A2(n3583), .ZN(n3042) );
  AND2_X1 U3787 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4377) );
  AOI21_X1 U3788 ( .B1(n3586), .B2(n3088), .A(n4377), .ZN(n3041) );
  OAI211_X1 U3789 ( .C1(n3624), .C2(n3137), .A(n3042), .B(n3041), .ZN(n3069)
         );
  NAND2_X1 U3790 ( .A1(n3585), .A2(n3416), .ZN(n3044) );
  NAND2_X1 U3791 ( .A1(n3136), .A2(n3417), .ZN(n3043) );
  NAND2_X1 U3792 ( .A1(n3044), .A2(n3043), .ZN(n3045) );
  XNOR2_X1 U3793 ( .A(n3045), .B(n3434), .ZN(n3096) );
  AOI22_X1 U3794 ( .A1(n3585), .A2(n3422), .B1(n3416), .B2(n3136), .ZN(n3097)
         );
  XNOR2_X1 U3795 ( .A(n3096), .B(n3097), .ZN(n3067) );
  AND2_X1 U3796 ( .A1(n3046), .A2(n2307), .ZN(n3543) );
  NAND2_X1 U3797 ( .A1(n3088), .A2(n3416), .ZN(n3048) );
  NAND2_X1 U3798 ( .A1(n3551), .A2(n3417), .ZN(n3047) );
  NAND2_X1 U3799 ( .A1(n3048), .A2(n3047), .ZN(n3049) );
  XNOR2_X1 U3800 ( .A(n3049), .B(n3446), .ZN(n3051) );
  AOI22_X1 U3801 ( .A1(n3088), .A2(n3422), .B1(n3416), .B2(n3551), .ZN(n3052)
         );
  XNOR2_X1 U3802 ( .A(n3051), .B(n3052), .ZN(n3547) );
  AND2_X1 U3803 ( .A1(n3543), .A2(n3547), .ZN(n3062) );
  NAND2_X1 U3804 ( .A1(n3544), .A2(n3062), .ZN(n3056) );
  INV_X1 U3805 ( .A(n3545), .ZN(n3050) );
  NAND2_X1 U3806 ( .A1(n3547), .A2(n3050), .ZN(n3055) );
  INV_X1 U3807 ( .A(n3051), .ZN(n3053) );
  NAND2_X1 U3808 ( .A1(n3053), .A2(n3052), .ZN(n3054) );
  AND2_X1 U3809 ( .A1(n3055), .A2(n3054), .ZN(n3057) );
  NAND2_X1 U3810 ( .A1(n3056), .A2(n3057), .ZN(n3066) );
  AND2_X1 U3811 ( .A1(n3059), .A2(n3064), .ZN(n3060) );
  NAND2_X1 U3812 ( .A1(n3103), .A2(n3100), .ZN(n3065) );
  AOI211_X1 U3813 ( .C1(n3067), .C2(n3066), .A(n3616), .B(n3065), .ZN(n3068)
         );
  AOI211_X1 U3814 ( .C1(n3070), .C2(n3614), .A(n3069), .B(n3068), .ZN(n3071)
         );
  INV_X1 U3815 ( .A(n3071), .ZN(U3214) );
  INV_X1 U3816 ( .A(n3072), .ZN(n3073) );
  NAND2_X1 U3817 ( .A1(n3073), .A2(n3727), .ZN(n3074) );
  NAND2_X1 U3818 ( .A1(n3074), .A2(n3719), .ZN(n3128) );
  INV_X1 U3819 ( .A(n3585), .ZN(n3138) );
  NAND2_X1 U3820 ( .A1(n3138), .A2(n3136), .ZN(n3730) );
  NAND2_X1 U3821 ( .A1(n3585), .A2(n3137), .ZN(n3734) );
  NAND2_X1 U3822 ( .A1(n3730), .A2(n3734), .ZN(n3687) );
  INV_X1 U3823 ( .A(n3687), .ZN(n3075) );
  XNOR2_X1 U3824 ( .A(n3128), .B(n3075), .ZN(n3079) );
  NAND2_X1 U3825 ( .A1(n3136), .A2(n4216), .ZN(n3077) );
  NAND2_X1 U3826 ( .A1(n3088), .A2(n3210), .ZN(n3076) );
  OAI211_X1 U3827 ( .C1(n3141), .C2(n4128), .A(n3077), .B(n3076), .ZN(n3078)
         );
  AOI21_X1 U3828 ( .B1(n3079), .B2(n4184), .A(n3078), .ZN(n3178) );
  AOI21_X1 U3829 ( .B1(n3136), .B2(n2203), .A(n3204), .ZN(n3183) );
  INV_X1 U3830 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3082) );
  OAI22_X1 U3831 ( .A1(n4198), .A2(n3082), .B1(n3081), .B2(n4196), .ZN(n3083)
         );
  AOI21_X1 U3832 ( .B1(n3183), .B2(n4479), .A(n3083), .ZN(n3095) );
  INV_X1 U3833 ( .A(n3084), .ZN(n3093) );
  AND2_X1 U3834 ( .A1(n3086), .A2(n3085), .ZN(n3091) );
  AND2_X1 U3835 ( .A1(n2152), .A2(n3089), .ZN(n3090) );
  NOR2_X1 U3836 ( .A1(n3091), .A2(n3090), .ZN(n3092) );
  XNOR2_X1 U3837 ( .A(n3140), .B(n3687), .ZN(n3176) );
  NAND2_X1 U3838 ( .A1(n3176), .A2(n3953), .ZN(n3094) );
  OAI211_X1 U3839 ( .C1(n3178), .C2(n4477), .A(n3095), .B(n3094), .ZN(U3280)
         );
  INV_X1 U3840 ( .A(n3096), .ZN(n3099) );
  INV_X1 U3841 ( .A(n3097), .ZN(n3098) );
  NAND2_X1 U3842 ( .A1(n3099), .A2(n3098), .ZN(n3101) );
  AND2_X1 U3843 ( .A1(n3101), .A2(n3100), .ZN(n3102) );
  NAND2_X1 U3844 ( .A1(n3103), .A2(n3102), .ZN(n3581) );
  OAI21_X1 U3845 ( .B1(n3154), .B2(IR_REG_10__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n3104) );
  OR2_X1 U3846 ( .A1(n3104), .A2(n3152), .ZN(n3105) );
  NAND2_X1 U3847 ( .A1(n3104), .A2(n3152), .ZN(n3109) );
  MUX2_X1 U3848 ( .A(n3830), .B(DATAI_11_), .S(n3349), .Z(n3587) );
  OAI22_X1 U3849 ( .A1(n3141), .A2(n3445), .B1(n3373), .B2(n3207), .ZN(n3578)
         );
  OAI22_X1 U3850 ( .A1(n3141), .A2(n3373), .B1(n3448), .B2(n3207), .ZN(n3106)
         );
  XNOR2_X1 U3851 ( .A(n3106), .B(n3446), .ZN(n3579) );
  OAI21_X1 U3852 ( .B1(n3581), .B2(n3578), .A(n3579), .ZN(n3108) );
  NAND2_X1 U3853 ( .A1(n3581), .A2(n3578), .ZN(n3107) );
  NAND2_X1 U3854 ( .A1(n3109), .A2(IR_REG_31__SCAN_IN), .ZN(n3110) );
  XNOR2_X1 U3855 ( .A(n3110), .B(IR_REG_12__SCAN_IN), .ZN(n3832) );
  INV_X1 U3856 ( .A(DATAI_12_), .ZN(n4571) );
  MUX2_X1 U3857 ( .A(n4495), .B(n4571), .S(n3349), .Z(n3228) );
  OAI22_X1 U3858 ( .A1(n3237), .A2(n3373), .B1(n3448), .B2(n3228), .ZN(n3111)
         );
  XNOR2_X1 U3859 ( .A(n3111), .B(n3446), .ZN(n3112) );
  OAI22_X1 U3860 ( .A1(n3237), .A2(n3445), .B1(n3373), .B2(n3228), .ZN(n3113)
         );
  INV_X1 U3861 ( .A(n3112), .ZN(n3115) );
  INV_X1 U3862 ( .A(n3113), .ZN(n3114) );
  NAND2_X1 U3863 ( .A1(n3115), .A2(n3114), .ZN(n3149) );
  NAND2_X1 U3864 ( .A1(n2172), .A2(n3149), .ZN(n3116) );
  XNOR2_X1 U3865 ( .A(n3148), .B(n3116), .ZN(n3117) );
  NAND2_X1 U3866 ( .A1(n3117), .A2(n3621), .ZN(n3127) );
  NAND2_X1 U3867 ( .A1(n3297), .A2(REG1_REG_13__SCAN_IN), .ZN(n3123) );
  NAND2_X1 U3868 ( .A1(n3632), .A2(REG2_REG_13__SCAN_IN), .ZN(n3122) );
  INV_X1 U3869 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4340) );
  OR2_X1 U3870 ( .A1(n3634), .A2(n4340), .ZN(n3121) );
  OR2_X1 U3871 ( .A1(n3118), .A2(REG3_REG_13__SCAN_IN), .ZN(n3119) );
  NAND2_X1 U3872 ( .A1(n3163), .A2(n3119), .ZN(n3242) );
  OR2_X1 U3873 ( .A1(n3459), .A2(n3242), .ZN(n3120) );
  OAI22_X1 U3874 ( .A1(n3624), .A2(n3228), .B1(n3265), .B2(n3626), .ZN(n3125)
         );
  NAND2_X1 U3875 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4392) );
  OAI21_X1 U3876 ( .B1(n3141), .B2(n3623), .A(n4392), .ZN(n3124) );
  NOR2_X1 U3877 ( .A1(n3125), .A2(n3124), .ZN(n3126) );
  OAI211_X1 U3878 ( .C1(n3631), .C2(n3143), .A(n3127), .B(n3126), .ZN(U3221)
         );
  NAND2_X1 U3879 ( .A1(n3128), .A2(n3734), .ZN(n3129) );
  NAND2_X1 U3880 ( .A1(n3129), .A2(n3730), .ZN(n3206) );
  NAND2_X1 U3881 ( .A1(n3130), .A2(n3207), .ZN(n3733) );
  NAND2_X1 U3882 ( .A1(n3206), .A2(n3733), .ZN(n3263) );
  NAND2_X1 U3883 ( .A1(n3141), .A2(n3587), .ZN(n3259) );
  NAND2_X1 U3884 ( .A1(n3263), .A2(n3259), .ZN(n3234) );
  NAND2_X1 U3885 ( .A1(n3237), .A2(n3229), .ZN(n3258) );
  NAND2_X1 U3886 ( .A1(n3584), .A2(n3228), .ZN(n3257) );
  NAND2_X1 U3887 ( .A1(n3258), .A2(n3257), .ZN(n3688) );
  INV_X1 U3888 ( .A(n3688), .ZN(n3131) );
  XNOR2_X1 U3889 ( .A(n3234), .B(n3131), .ZN(n3135) );
  OAI22_X1 U3890 ( .A1(n3265), .A2(n4128), .B1(n4127), .B2(n3228), .ZN(n3133)
         );
  NOR2_X1 U3891 ( .A1(n3141), .A2(n4191), .ZN(n3132) );
  OR2_X1 U3892 ( .A1(n3133), .A2(n3132), .ZN(n3134) );
  AOI21_X1 U3893 ( .B1(n3135), .B2(n4184), .A(n3134), .ZN(n3219) );
  NOR2_X1 U3894 ( .A1(n3585), .A2(n3136), .ZN(n3139) );
  XNOR2_X1 U3895 ( .A(n3227), .B(n3688), .ZN(n3218) );
  NAND2_X1 U3896 ( .A1(n3204), .A2(n3207), .ZN(n3203) );
  NAND2_X1 U3897 ( .A1(n3203), .A2(n3229), .ZN(n3142) );
  NAND2_X1 U3898 ( .A1(n3241), .A2(n3142), .ZN(n3226) );
  NOR2_X1 U3899 ( .A1(n4196), .A2(n3143), .ZN(n3144) );
  AOI21_X1 U3900 ( .B1(n4477), .B2(REG2_REG_12__SCAN_IN), .A(n3144), .ZN(n3145) );
  OAI21_X1 U3901 ( .B1(n3226), .B2(n4195), .A(n3145), .ZN(n3146) );
  AOI21_X1 U3902 ( .B1(n3218), .B2(n3953), .A(n3146), .ZN(n3147) );
  OAI21_X1 U3903 ( .B1(n4477), .B2(n3219), .A(n3147), .ZN(U3278) );
  INV_X1 U3904 ( .A(IR_REG_10__SCAN_IN), .ZN(n3151) );
  INV_X1 U3905 ( .A(IR_REG_12__SCAN_IN), .ZN(n3150) );
  NAND3_X1 U3906 ( .A1(n3152), .A2(n3151), .A3(n3150), .ZN(n3153) );
  OAI21_X1 U3907 ( .B1(n3154), .B2(n3153), .A(IR_REG_31__SCAN_IN), .ZN(n3155)
         );
  MUX2_X1 U3908 ( .A(IR_REG_31__SCAN_IN), .B(n3155), .S(IR_REG_13__SCAN_IN), 
        .Z(n3157) );
  INV_X1 U3909 ( .A(n3327), .ZN(n3156) );
  INV_X1 U3910 ( .A(DATAI_13_), .ZN(n3158) );
  MUX2_X1 U3911 ( .A(n4494), .B(n3158), .S(n3349), .Z(n3249) );
  OAI22_X1 U3912 ( .A1(n3265), .A2(n3373), .B1(n3448), .B2(n3249), .ZN(n3159)
         );
  XNOR2_X1 U3913 ( .A(n3159), .B(n3434), .ZN(n3187) );
  OAI22_X1 U3914 ( .A1(n3265), .A2(n3445), .B1(n2649), .B2(n3249), .ZN(n3185)
         );
  XNOR2_X1 U3915 ( .A(n3187), .B(n3185), .ZN(n3160) );
  XNOR2_X1 U3916 ( .A(n3188), .B(n3160), .ZN(n3161) );
  NAND2_X1 U3917 ( .A1(n3161), .A2(n3621), .ZN(n3175) );
  OAI22_X1 U3918 ( .A1(n3624), .A2(n3249), .B1(n3237), .B2(n3623), .ZN(n3173)
         );
  NAND2_X1 U3919 ( .A1(n3632), .A2(REG2_REG_14__SCAN_IN), .ZN(n3169) );
  NAND2_X1 U3920 ( .A1(n3297), .A2(REG1_REG_14__SCAN_IN), .ZN(n3168) );
  NAND2_X1 U3921 ( .A1(n3163), .A2(n3162), .ZN(n3164) );
  NAND2_X1 U3922 ( .A1(n3165), .A2(n3164), .ZN(n3273) );
  OR2_X1 U3923 ( .A1(n3459), .A2(n3273), .ZN(n3167) );
  INV_X1 U3924 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4336) );
  OR2_X1 U3925 ( .A1(n3634), .A2(n4336), .ZN(n3166) );
  INV_X1 U3926 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3170) );
  NOR2_X1 U3927 ( .A1(STATE_REG_SCAN_IN), .A2(n3170), .ZN(n4406) );
  INV_X1 U3928 ( .A(n4406), .ZN(n3171) );
  OAI21_X1 U3929 ( .B1(n4192), .B2(n3626), .A(n3171), .ZN(n3172) );
  NOR2_X1 U3930 ( .A1(n3173), .A2(n3172), .ZN(n3174) );
  OAI211_X1 U3931 ( .C1(n3631), .C2(n3242), .A(n3175), .B(n3174), .ZN(U3231)
         );
  NAND2_X1 U3932 ( .A1(n3176), .A2(n4525), .ZN(n3177) );
  NAND2_X1 U3933 ( .A1(n3178), .A2(n3177), .ZN(n3181) );
  MUX2_X1 U3934 ( .A(REG0_REG_10__SCAN_IN), .B(n3181), .S(n4518), .Z(n3179) );
  AOI21_X1 U3935 ( .B1(n3183), .B2(n4307), .A(n3179), .ZN(n3180) );
  INV_X1 U3936 ( .A(n3180), .ZN(U3487) );
  MUX2_X1 U3937 ( .A(REG1_REG_10__SCAN_IN), .B(n3181), .S(n4544), .Z(n3182) );
  AOI21_X1 U3938 ( .B1(n4242), .B2(n3183), .A(n3182), .ZN(n3184) );
  INV_X1 U3939 ( .A(n3184), .ZN(U3528) );
  NAND2_X1 U3940 ( .A1(n3188), .A2(n3187), .ZN(n3186) );
  NAND2_X1 U3941 ( .A1(n3186), .A2(n3185), .ZN(n3290) );
  NAND2_X1 U3942 ( .A1(n3290), .A2(n3287), .ZN(n3197) );
  OR2_X1 U3943 ( .A1(n3327), .A2(n3189), .ZN(n3190) );
  XNOR2_X1 U3944 ( .A(n3190), .B(IR_REG_14__SCAN_IN), .ZN(n4421) );
  MUX2_X1 U3945 ( .A(n4421), .B(DATAI_14_), .S(n3349), .Z(n3887) );
  INV_X1 U3946 ( .A(n3887), .ZN(n3271) );
  OAI22_X1 U3947 ( .A1(n4192), .A2(n3373), .B1(n3448), .B2(n3271), .ZN(n3191)
         );
  XNOR2_X1 U3948 ( .A(n3191), .B(n3446), .ZN(n3192) );
  OAI22_X1 U3949 ( .A1(n4192), .A2(n3445), .B1(n2649), .B2(n3271), .ZN(n3193)
         );
  NAND2_X1 U3950 ( .A1(n3192), .A2(n3193), .ZN(n3286) );
  INV_X1 U3951 ( .A(n3192), .ZN(n3195) );
  INV_X1 U3952 ( .A(n3193), .ZN(n3194) );
  NAND2_X1 U3953 ( .A1(n3195), .A2(n3194), .ZN(n3288) );
  NAND2_X1 U3954 ( .A1(n3286), .A2(n3288), .ZN(n3196) );
  XNOR2_X1 U3955 ( .A(n3197), .B(n3196), .ZN(n3198) );
  NAND2_X1 U3956 ( .A1(n3198), .A2(n3621), .ZN(n3202) );
  OAI22_X1 U3957 ( .A1(n3624), .A2(n3271), .B1(n4168), .B2(n3626), .ZN(n3200)
         );
  NAND2_X1 U3958 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4423) );
  OAI21_X1 U3959 ( .B1(n3265), .B2(n3623), .A(n4423), .ZN(n3199) );
  NOR2_X1 U3960 ( .A1(n3200), .A2(n3199), .ZN(n3201) );
  OAI211_X1 U3961 ( .C1(n3631), .C2(n3273), .A(n3202), .B(n3201), .ZN(U3212)
         );
  OAI21_X1 U3962 ( .B1(n3204), .B2(n3207), .A(n3203), .ZN(n3280) );
  INV_X1 U3963 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4677) );
  AOI21_X1 U3964 ( .B1(n3690), .B2(n3205), .A(n2162), .ZN(n3285) );
  INV_X1 U3965 ( .A(n3285), .ZN(n3213) );
  XOR2_X1 U3966 ( .A(n3690), .B(n3206), .Z(n3212) );
  OAI22_X1 U3967 ( .A1(n3237), .A2(n4128), .B1(n4127), .B2(n3207), .ZN(n3209)
         );
  NOR2_X1 U3968 ( .A1(n3285), .A2(n4089), .ZN(n3208) );
  AOI211_X1 U3969 ( .C1(n3210), .C2(n3585), .A(n3209), .B(n3208), .ZN(n3211)
         );
  OAI21_X1 U3970 ( .B1(n4025), .B2(n3212), .A(n3211), .ZN(n3279) );
  AOI21_X1 U3971 ( .B1(n4510), .B2(n3213), .A(n3279), .ZN(n3215) );
  MUX2_X1 U3972 ( .A(n4677), .B(n3215), .S(n4547), .Z(n3214) );
  OAI21_X1 U3973 ( .B1(n4286), .B2(n3280), .A(n3214), .ZN(U3529) );
  MUX2_X1 U3974 ( .A(n3216), .B(n3215), .S(n4518), .Z(n3217) );
  OAI21_X1 U3975 ( .B1(n3280), .B2(n4342), .A(n3217), .ZN(U3489) );
  NAND2_X1 U3976 ( .A1(n3218), .A2(n4525), .ZN(n3220) );
  NAND2_X1 U3977 ( .A1(n3220), .A2(n3219), .ZN(n3223) );
  MUX2_X1 U3978 ( .A(n3223), .B(REG0_REG_12__SCAN_IN), .S(n4790), .Z(n3221) );
  INV_X1 U3979 ( .A(n3221), .ZN(n3222) );
  OAI21_X1 U3980 ( .B1(n3226), .B2(n4342), .A(n3222), .ZN(U3491) );
  MUX2_X1 U3981 ( .A(n3223), .B(REG1_REG_12__SCAN_IN), .S(n4545), .Z(n3224) );
  INV_X1 U3982 ( .A(n3224), .ZN(n3225) );
  OAI21_X1 U3983 ( .B1(n4286), .B2(n3226), .A(n3225), .ZN(U3530) );
  INV_X1 U3984 ( .A(n3227), .ZN(n3231) );
  NOR2_X1 U3985 ( .A1(n3778), .A2(n3249), .ZN(n3260) );
  NAND2_X1 U3986 ( .A1(n3778), .A2(n3249), .ZN(n3256) );
  INV_X1 U3987 ( .A(n3256), .ZN(n3232) );
  NOR2_X1 U3988 ( .A1(n3260), .A2(n3232), .ZN(n3683) );
  XNOR2_X1 U3989 ( .A(n3248), .B(n3683), .ZN(n4281) );
  INV_X1 U3990 ( .A(n3258), .ZN(n3233) );
  OAI21_X1 U3991 ( .B1(n3234), .B2(n3233), .A(n3257), .ZN(n3235) );
  XOR2_X1 U3992 ( .A(n3683), .B(n3235), .Z(n3239) );
  AOI22_X1 U3993 ( .A1(n3888), .A2(n4187), .B1(n4216), .B2(n3250), .ZN(n3236)
         );
  OAI21_X1 U3994 ( .B1(n3237), .B2(n4191), .A(n3236), .ZN(n3238) );
  AOI21_X1 U3995 ( .B1(n3239), .B2(n4184), .A(n3238), .ZN(n3240) );
  OAI21_X1 U3996 ( .B1(n4281), .B2(n4089), .A(n3240), .ZN(n4282) );
  NAND2_X1 U3997 ( .A1(n4282), .A2(n4198), .ZN(n3247) );
  OAI21_X1 U3998 ( .B1(n2195), .B2(n3249), .A(n3269), .ZN(n4343) );
  INV_X1 U3999 ( .A(n4343), .ZN(n3245) );
  INV_X1 U4000 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3243) );
  OAI22_X1 U4001 ( .A1(n4198), .A2(n3243), .B1(n3242), .B2(n4196), .ZN(n3244)
         );
  AOI21_X1 U4002 ( .B1(n3245), .B2(n4479), .A(n3244), .ZN(n3246) );
  OAI211_X1 U4003 ( .C1(n4281), .C2(n4099), .A(n3247), .B(n3246), .ZN(U3277)
         );
  NAND2_X1 U4004 ( .A1(n4192), .A2(n3887), .ZN(n4180) );
  NAND2_X1 U4005 ( .A1(n3888), .A2(n3271), .ZN(n3639) );
  NAND2_X1 U4006 ( .A1(n4180), .A2(n3639), .ZN(n3255) );
  OAI21_X1 U4007 ( .B1(n3254), .B2(n3255), .A(n3889), .ZN(n4279) );
  INV_X1 U4008 ( .A(n4279), .ZN(n3278) );
  NAND2_X1 U4009 ( .A1(n3257), .A2(n3256), .ZN(n3736) );
  NAND2_X1 U4010 ( .A1(n3259), .A2(n3258), .ZN(n3262) );
  INV_X1 U4011 ( .A(n3736), .ZN(n3261) );
  AOI21_X1 U4012 ( .B1(n3262), .B2(n3261), .A(n3260), .ZN(n3740) );
  OAI21_X2 U4013 ( .B1(n3263), .B2(n3736), .A(n3740), .ZN(n3638) );
  NAND2_X2 U4014 ( .A1(n3638), .A2(n2274), .ZN(n4181) );
  OAI21_X1 U4015 ( .B1(n2274), .B2(n3638), .A(n4181), .ZN(n3267) );
  AOI22_X1 U4016 ( .A1(n3890), .A2(n4187), .B1(n4216), .B2(n3887), .ZN(n3264)
         );
  OAI21_X1 U4017 ( .B1(n3265), .B2(n4191), .A(n3264), .ZN(n3266) );
  AOI21_X1 U4018 ( .B1(n3267), .B2(n4184), .A(n3266), .ZN(n3268) );
  OAI21_X1 U4019 ( .B1(n3278), .B2(n4089), .A(n3268), .ZN(n4278) );
  NAND2_X1 U4020 ( .A1(n4278), .A2(n4198), .ZN(n3277) );
  INV_X1 U4021 ( .A(n3269), .ZN(n3272) );
  INV_X1 U4022 ( .A(n4194), .ZN(n3270) );
  OAI21_X1 U4023 ( .B1(n3272), .B2(n3271), .A(n3270), .ZN(n4338) );
  INV_X1 U4024 ( .A(n4338), .ZN(n3275) );
  OAI22_X1 U4025 ( .A1(n4198), .A2(n4696), .B1(n3273), .B2(n4196), .ZN(n3274)
         );
  AOI21_X1 U4026 ( .B1(n3275), .B2(n4479), .A(n3274), .ZN(n3276) );
  OAI211_X1 U4027 ( .C1(n3278), .C2(n4099), .A(n3277), .B(n3276), .ZN(U3276)
         );
  NAND2_X1 U4028 ( .A1(n3279), .A2(n4198), .ZN(n3284) );
  INV_X1 U4029 ( .A(n3280), .ZN(n3282) );
  OAI22_X1 U4030 ( .A1(n4198), .A2(n3829), .B1(n3589), .B2(n4196), .ZN(n3281)
         );
  AOI21_X1 U4031 ( .B1(n3282), .B2(n4479), .A(n3281), .ZN(n3283) );
  OAI211_X1 U4032 ( .C1(n3285), .C2(n4099), .A(n3284), .B(n3283), .ZN(U3279)
         );
  NAND2_X1 U4033 ( .A1(n3327), .A2(n4797), .ZN(n3292) );
  NAND2_X1 U4034 ( .A1(n3292), .A2(IR_REG_31__SCAN_IN), .ZN(n3307) );
  XNOR2_X1 U4035 ( .A(n3307), .B(IR_REG_15__SCAN_IN), .ZN(n3841) );
  MUX2_X1 U4036 ( .A(n3841), .B(DATAI_15_), .S(n3349), .Z(n4186) );
  OAI22_X1 U4037 ( .A1(n4168), .A2(n3373), .B1(n3448), .B2(n4193), .ZN(n3293)
         );
  XNOR2_X1 U4038 ( .A(n3293), .B(n3446), .ZN(n3295) );
  AND2_X1 U4039 ( .A1(n4186), .A2(n3416), .ZN(n3294) );
  AOI21_X1 U4040 ( .B1(n3890), .B2(n3422), .A(n3294), .ZN(n3619) );
  NAND2_X1 U4041 ( .A1(n3632), .A2(REG2_REG_16__SCAN_IN), .ZN(n3305) );
  NAND2_X1 U4042 ( .A1(n3297), .A2(REG1_REG_16__SCAN_IN), .ZN(n3304) );
  AND2_X1 U40430 ( .A1(n3299), .A2(n3298), .ZN(n3301) );
  OR2_X1 U4044 ( .A1(n3301), .A2(n3300), .ZN(n4173) );
  OR2_X1 U4045 ( .A1(n3459), .A2(n4173), .ZN(n3303) );
  INV_X1 U4046 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4648) );
  OR2_X1 U4047 ( .A1(n3634), .A2(n4648), .ZN(n3302) );
  NAND2_X1 U4048 ( .A1(n3307), .A2(n3306), .ZN(n3308) );
  NAND2_X1 U4049 ( .A1(n3308), .A2(IR_REG_31__SCAN_IN), .ZN(n3310) );
  XNOR2_X1 U4050 ( .A(n3310), .B(n3309), .ZN(n4491) );
  INV_X1 U4051 ( .A(n4491), .ZN(n3311) );
  MUX2_X1 U4052 ( .A(n3311), .B(DATAI_16_), .S(n3349), .Z(n4172) );
  OAI22_X1 U4053 ( .A1(n4152), .A2(n3445), .B1(n3373), .B2(n3892), .ZN(n3313)
         );
  OAI22_X1 U4054 ( .A1(n4152), .A2(n3373), .B1(n3448), .B2(n3892), .ZN(n3312)
         );
  XNOR2_X1 U4055 ( .A(n3312), .B(n3446), .ZN(n3314) );
  XOR2_X1 U4056 ( .A(n3313), .B(n3314), .Z(n3518) );
  NAND2_X1 U4057 ( .A1(n3315), .A2(IR_REG_31__SCAN_IN), .ZN(n3316) );
  XNOR2_X1 U4058 ( .A(n3316), .B(IR_REG_17__SCAN_IN), .ZN(n3843) );
  INV_X1 U4059 ( .A(DATAI_17_), .ZN(n4565) );
  MUX2_X1 U4060 ( .A(n4490), .B(n4565), .S(n3349), .Z(n4155) );
  OAI22_X1 U4061 ( .A1(n4130), .A2(n3373), .B1(n3448), .B2(n4155), .ZN(n3317)
         );
  XOR2_X1 U4062 ( .A(n3446), .B(n3317), .Z(n3526) );
  INV_X1 U4063 ( .A(n3526), .ZN(n3318) );
  OAI22_X1 U4064 ( .A1(n4130), .A2(n3445), .B1(n2649), .B2(n4155), .ZN(n3525)
         );
  INV_X1 U4065 ( .A(n3525), .ZN(n3319) );
  NAND2_X1 U4066 ( .A1(n3297), .A2(REG1_REG_18__SCAN_IN), .ZN(n3326) );
  NAND2_X1 U4067 ( .A1(n3632), .A2(REG2_REG_18__SCAN_IN), .ZN(n3325) );
  INV_X1 U4068 ( .A(REG0_REG_18__SCAN_IN), .ZN(n3320) );
  OR2_X1 U4069 ( .A1(n3634), .A2(n3320), .ZN(n3324) );
  NAND2_X1 U4070 ( .A1(n3321), .A2(n4773), .ZN(n3322) );
  NAND2_X1 U4071 ( .A1(n3337), .A2(n3322), .ZN(n4138) );
  OR2_X1 U4072 ( .A1(n3459), .A2(n4138), .ZN(n3323) );
  NAND2_X1 U4073 ( .A1(n3327), .A2(n3328), .ZN(n3329) );
  NAND2_X1 U4074 ( .A1(n3329), .A2(IR_REG_31__SCAN_IN), .ZN(n3330) );
  XNOR2_X1 U4075 ( .A(n3330), .B(IR_REG_18__SCAN_IN), .ZN(n3844) );
  MUX2_X1 U4076 ( .A(n3844), .B(DATAI_18_), .S(n3349), .Z(n3895) );
  OAI22_X1 U4077 ( .A1(n4114), .A2(n3373), .B1(n3448), .B2(n3896), .ZN(n3331)
         );
  XNOR2_X1 U4078 ( .A(n3331), .B(n3446), .ZN(n3332) );
  OAI22_X1 U4079 ( .A1(n4114), .A2(n3445), .B1(n2649), .B2(n3896), .ZN(n3333)
         );
  AND2_X1 U4080 ( .A1(n3332), .A2(n3333), .ZN(n3595) );
  INV_X1 U4081 ( .A(n3332), .ZN(n3335) );
  INV_X1 U4082 ( .A(n3333), .ZN(n3334) );
  NAND2_X1 U4083 ( .A1(n3335), .A2(n3334), .ZN(n3596) );
  NAND2_X1 U4084 ( .A1(n3632), .A2(REG2_REG_19__SCAN_IN), .ZN(n3343) );
  NAND2_X1 U4085 ( .A1(n3297), .A2(REG1_REG_19__SCAN_IN), .ZN(n3342) );
  AND2_X1 U4086 ( .A1(n3337), .A2(n3336), .ZN(n3339) );
  OR2_X1 U4087 ( .A1(n3339), .A2(n3338), .ZN(n4117) );
  OR2_X1 U4088 ( .A1(n2536), .A2(n4117), .ZN(n3341) );
  INV_X1 U4089 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4323) );
  OR2_X1 U4090 ( .A1(n3634), .A2(n4323), .ZN(n3340) );
  MUX2_X1 U4091 ( .A(n4350), .B(DATAI_19_), .S(n3349), .Z(n4110) );
  OAI22_X1 U4092 ( .A1(n4129), .A2(n3445), .B1(n3373), .B2(n4116), .ZN(n3346)
         );
  OAI22_X1 U4093 ( .A1(n4129), .A2(n3373), .B1(n3448), .B2(n4116), .ZN(n3344)
         );
  XNOR2_X1 U4094 ( .A(n3344), .B(n3446), .ZN(n3345) );
  XOR2_X1 U4095 ( .A(n3346), .B(n3345), .Z(n3489) );
  INV_X1 U4096 ( .A(n3345), .ZN(n3348) );
  INV_X1 U4097 ( .A(n3346), .ZN(n3347) );
  OAI22_X1 U4098 ( .A1(n4066), .A2(n3373), .B1(n3448), .B2(n4091), .ZN(n3350)
         );
  XNOR2_X1 U4099 ( .A(n3350), .B(n3446), .ZN(n3351) );
  OAI22_X1 U4100 ( .A1(n4066), .A2(n3445), .B1(n3373), .B2(n4091), .ZN(n3352)
         );
  AND2_X1 U4101 ( .A1(n3351), .A2(n3352), .ZN(n3559) );
  INV_X1 U4102 ( .A(n3351), .ZN(n3354) );
  INV_X1 U4103 ( .A(n3352), .ZN(n3353) );
  OR2_X1 U4104 ( .A1(n3355), .A2(REG3_REG_21__SCAN_IN), .ZN(n3356) );
  NAND2_X1 U4105 ( .A1(n3367), .A2(n3356), .ZN(n4071) );
  OR2_X1 U4106 ( .A1(n2536), .A2(n4071), .ZN(n3360) );
  INV_X1 U4107 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4315) );
  OR2_X1 U4108 ( .A1(n3634), .A2(n4315), .ZN(n3359) );
  NAND2_X1 U4109 ( .A1(n3632), .A2(REG2_REG_21__SCAN_IN), .ZN(n3358) );
  NAND2_X1 U4110 ( .A1(n3297), .A2(REG1_REG_21__SCAN_IN), .ZN(n3357) );
  NAND4_X1 U4111 ( .A1(n3360), .A2(n3359), .A3(n3358), .A4(n3357), .ZN(n4084)
         );
  NAND2_X1 U4112 ( .A1(n4084), .A2(n3416), .ZN(n3362) );
  NAND2_X1 U4113 ( .A1(n4062), .A2(n3417), .ZN(n3361) );
  NAND2_X1 U4114 ( .A1(n3362), .A2(n3361), .ZN(n3363) );
  XNOR2_X1 U4115 ( .A(n3363), .B(n3434), .ZN(n3496) );
  AND2_X1 U4116 ( .A1(n4062), .A2(n3416), .ZN(n3364) );
  AOI21_X1 U4117 ( .B1(n4084), .B2(n3422), .A(n3364), .ZN(n3495) );
  INV_X1 U4118 ( .A(n3496), .ZN(n3366) );
  INV_X1 U4119 ( .A(n3495), .ZN(n3365) );
  NAND2_X1 U4120 ( .A1(n3367), .A2(n3571), .ZN(n3368) );
  NAND2_X1 U4121 ( .A1(n3378), .A2(n3368), .ZN(n3573) );
  OR2_X1 U4122 ( .A1(n3459), .A2(n3573), .ZN(n3372) );
  INV_X1 U4123 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4651) );
  OR2_X1 U4124 ( .A1(n3634), .A2(n4651), .ZN(n3371) );
  NAND2_X1 U4125 ( .A1(n3297), .A2(REG1_REG_22__SCAN_IN), .ZN(n3370) );
  NAND2_X1 U4126 ( .A1(n3632), .A2(REG2_REG_22__SCAN_IN), .ZN(n3369) );
  NAND4_X1 U4127 ( .A1(n3372), .A2(n3371), .A3(n3370), .A4(n3369), .ZN(n4063)
         );
  INV_X1 U4128 ( .A(n4063), .ZN(n4021) );
  OAI22_X1 U4129 ( .A1(n4021), .A2(n3445), .B1(n3373), .B2(n4052), .ZN(n3388)
         );
  NAND2_X1 U4130 ( .A1(n4063), .A2(n3416), .ZN(n3375) );
  NAND2_X1 U4131 ( .A1(n4045), .A2(n3417), .ZN(n3374) );
  NAND2_X1 U4132 ( .A1(n3375), .A2(n3374), .ZN(n3376) );
  XNOR2_X1 U4133 ( .A(n3376), .B(n3446), .ZN(n3387) );
  XOR2_X1 U4134 ( .A(n3388), .B(n3387), .Z(n3569) );
  NAND2_X1 U4135 ( .A1(n3568), .A2(n3569), .ZN(n3480) );
  AND2_X1 U4136 ( .A1(n3378), .A2(n3377), .ZN(n3380) );
  OR2_X1 U4137 ( .A1(n3380), .A2(n3379), .ZN(n4031) );
  AOI22_X1 U4138 ( .A1(n3412), .A2(REG0_REG_23__SCAN_IN), .B1(n3297), .B2(
        REG1_REG_23__SCAN_IN), .ZN(n3382) );
  NAND2_X1 U4139 ( .A1(n3632), .A2(REG2_REG_23__SCAN_IN), .ZN(n3381) );
  NAND2_X1 U4140 ( .A1(n4044), .A2(n3416), .ZN(n3384) );
  NAND2_X1 U4141 ( .A1(n3921), .A2(n3417), .ZN(n3383) );
  NAND2_X1 U4142 ( .A1(n3384), .A2(n3383), .ZN(n3385) );
  XNOR2_X1 U4143 ( .A(n3385), .B(n3446), .ZN(n3391) );
  NOR2_X1 U4144 ( .A1(n4029), .A2(n2649), .ZN(n3386) );
  AOI21_X1 U4145 ( .B1(n4044), .B2(n3422), .A(n3386), .ZN(n3392) );
  XNOR2_X1 U4146 ( .A(n3391), .B(n3392), .ZN(n3481) );
  INV_X1 U4147 ( .A(n3387), .ZN(n3390) );
  INV_X1 U4148 ( .A(n3388), .ZN(n3389) );
  NAND2_X1 U4149 ( .A1(n3390), .A2(n3389), .ZN(n3482) );
  INV_X1 U4150 ( .A(n3391), .ZN(n3393) );
  NOR2_X1 U4151 ( .A1(n3393), .A2(n3392), .ZN(n3403) );
  INV_X1 U4152 ( .A(n3403), .ZN(n3397) );
  NAND2_X1 U4153 ( .A1(n4023), .A2(n3422), .ZN(n3395) );
  NAND2_X1 U4154 ( .A1(n4006), .A2(n3416), .ZN(n3394) );
  NAND2_X1 U4155 ( .A1(n3395), .A2(n3394), .ZN(n3402) );
  INV_X1 U4156 ( .A(n3402), .ZN(n3396) );
  OAI22_X1 U4157 ( .A1(n3987), .A2(n3373), .B1(n3448), .B2(n3905), .ZN(n3399)
         );
  XOR2_X1 U4158 ( .A(n3446), .B(n3399), .Z(n3537) );
  INV_X1 U4159 ( .A(n3537), .ZN(n3400) );
  NAND2_X1 U4160 ( .A1(n4005), .A2(n3416), .ZN(n3405) );
  NAND2_X1 U4161 ( .A1(n3983), .A2(n3417), .ZN(n3404) );
  NAND2_X1 U4162 ( .A1(n3405), .A2(n3404), .ZN(n3406) );
  XNOR2_X1 U4163 ( .A(n3406), .B(n3434), .ZN(n3409) );
  NOR2_X1 U4164 ( .A1(n3990), .A2(n2649), .ZN(n3407) );
  AOI21_X1 U4165 ( .B1(n4005), .B2(n3422), .A(n3407), .ZN(n3408) );
  NAND2_X1 U4166 ( .A1(n3409), .A2(n3408), .ZN(n3506) );
  NOR2_X1 U4167 ( .A1(n3409), .A2(n3408), .ZN(n3508) );
  AOI21_X1 U4168 ( .B1(n3505), .B2(n3506), .A(n3508), .ZN(n3606) );
  INV_X1 U4169 ( .A(REG2_REG_26__SCAN_IN), .ZN(n3415) );
  NAND2_X1 U4170 ( .A1(n3410), .A2(REG3_REG_26__SCAN_IN), .ZN(n3427) );
  OR2_X1 U4171 ( .A1(n3410), .A2(REG3_REG_26__SCAN_IN), .ZN(n3411) );
  NAND2_X1 U4172 ( .A1(n3427), .A2(n3411), .ZN(n3611) );
  OR2_X1 U4173 ( .A1(n3611), .A2(n3459), .ZN(n3414) );
  AOI22_X1 U4174 ( .A1(n3412), .A2(REG0_REG_26__SCAN_IN), .B1(n3297), .B2(
        REG1_REG_26__SCAN_IN), .ZN(n3413) );
  OAI211_X1 U4175 ( .C1(n2453), .C2(n3415), .A(n3414), .B(n3413), .ZN(n3984)
         );
  NAND2_X1 U4176 ( .A1(n3984), .A2(n3416), .ZN(n3419) );
  INV_X1 U4177 ( .A(n3973), .ZN(n3677) );
  NAND2_X1 U4178 ( .A1(n3677), .A2(n3417), .ZN(n3418) );
  NAND2_X1 U4179 ( .A1(n3419), .A2(n3418), .ZN(n3420) );
  XNOR2_X1 U4180 ( .A(n3420), .B(n3434), .ZN(n3426) );
  INV_X1 U4181 ( .A(n3426), .ZN(n3424) );
  NOR2_X1 U4182 ( .A1(n3973), .A2(n2649), .ZN(n3421) );
  AOI21_X1 U4183 ( .B1(n3984), .B2(n3422), .A(n3421), .ZN(n3425) );
  INV_X1 U4184 ( .A(n3425), .ZN(n3423) );
  NAND2_X1 U4185 ( .A1(n3424), .A2(n3423), .ZN(n3608) );
  AND2_X1 U4186 ( .A1(n3426), .A2(n3425), .ZN(n3607) );
  INV_X1 U4187 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4777) );
  NAND2_X1 U4188 ( .A1(n3427), .A2(n4777), .ZN(n3428) );
  NAND2_X1 U4189 ( .A1(n3437), .A2(n3428), .ZN(n3955) );
  OR2_X1 U4190 ( .A1(n3955), .A2(n3459), .ZN(n3433) );
  INV_X1 U4191 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4669) );
  NAND2_X1 U4192 ( .A1(n3632), .A2(REG2_REG_27__SCAN_IN), .ZN(n3430) );
  NAND2_X1 U4193 ( .A1(n3297), .A2(REG1_REG_27__SCAN_IN), .ZN(n3429) );
  OAI211_X1 U4194 ( .C1(n3634), .C2(n4669), .A(n3430), .B(n3429), .ZN(n3431)
         );
  INV_X1 U4195 ( .A(n3431), .ZN(n3432) );
  OAI22_X1 U4196 ( .A1(n3935), .A2(n3373), .B1(n3954), .B2(n3448), .ZN(n3435)
         );
  XNOR2_X1 U4197 ( .A(n3435), .B(n3434), .ZN(n3453) );
  OAI22_X1 U4198 ( .A1(n3935), .A2(n3445), .B1(n3954), .B2(n2649), .ZN(n3451)
         );
  XNOR2_X1 U4199 ( .A(n3453), .B(n3451), .ZN(n3472) );
  NAND2_X1 U4200 ( .A1(n3473), .A2(n3472), .ZN(n3471) );
  INV_X1 U4201 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3436) );
  NAND2_X1 U4202 ( .A1(n3437), .A2(n3436), .ZN(n3438) );
  NAND2_X1 U4203 ( .A1(n3938), .A2(n3439), .ZN(n3444) );
  INV_X1 U4204 ( .A(REG0_REG_28__SCAN_IN), .ZN(n4668) );
  NAND2_X1 U4205 ( .A1(n3297), .A2(REG1_REG_28__SCAN_IN), .ZN(n3441) );
  NAND2_X1 U4206 ( .A1(n3632), .A2(REG2_REG_28__SCAN_IN), .ZN(n3440) );
  OAI211_X1 U4207 ( .C1(n3634), .C2(n4668), .A(n3441), .B(n3440), .ZN(n3442)
         );
  INV_X1 U4208 ( .A(n3442), .ZN(n3443) );
  INV_X1 U4209 ( .A(n3937), .ZN(n3655) );
  OAI22_X1 U4210 ( .A1(n3946), .A2(n3445), .B1(n3373), .B2(n3655), .ZN(n3447)
         );
  XNOR2_X1 U4211 ( .A(n3447), .B(n3446), .ZN(n3450) );
  OAI22_X1 U4212 ( .A1(n3946), .A2(n3373), .B1(n3448), .B2(n3655), .ZN(n3449)
         );
  XNOR2_X1 U4213 ( .A(n3450), .B(n3449), .ZN(n3462) );
  NAND2_X1 U4214 ( .A1(n3462), .A2(n3621), .ZN(n3470) );
  INV_X1 U4215 ( .A(n3451), .ZN(n3452) );
  NOR2_X1 U4216 ( .A1(n3453), .A2(n3452), .ZN(n3463) );
  NOR3_X1 U4217 ( .A1(n3462), .A2(n3463), .A3(n3616), .ZN(n3454) );
  NAND2_X1 U4218 ( .A1(n3471), .A2(n3454), .ZN(n3469) );
  INV_X1 U4219 ( .A(REG0_REG_29__SCAN_IN), .ZN(n4666) );
  NAND2_X1 U4220 ( .A1(n3632), .A2(REG2_REG_29__SCAN_IN), .ZN(n3456) );
  NAND2_X1 U4221 ( .A1(n3297), .A2(REG1_REG_29__SCAN_IN), .ZN(n3455) );
  OAI211_X1 U4222 ( .C1(n4666), .C2(n3634), .A(n3456), .B(n3455), .ZN(n3457)
         );
  INV_X1 U4223 ( .A(n3457), .ZN(n3458) );
  OAI21_X1 U4224 ( .B1(n3853), .B2(n3459), .A(n3458), .ZN(n3932) );
  AOI22_X1 U4225 ( .A1(n3932), .A2(n3583), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3461) );
  NAND2_X1 U4226 ( .A1(n3588), .A2(n3937), .ZN(n3460) );
  OAI211_X1 U4227 ( .C1(n3935), .C2(n3623), .A(n3461), .B(n3460), .ZN(n3467)
         );
  INV_X1 U4228 ( .A(n3462), .ZN(n3465) );
  INV_X1 U4229 ( .A(n3463), .ZN(n3464) );
  NOR3_X1 U4230 ( .A1(n3465), .A2(n3616), .A3(n3464), .ZN(n3466) );
  AOI211_X1 U4231 ( .C1(n3938), .C2(n3614), .A(n3467), .B(n3466), .ZN(n3468)
         );
  OAI211_X1 U4232 ( .C1(n3471), .C2(n3470), .A(n3469), .B(n3468), .ZN(U3217)
         );
  XNOR2_X1 U4233 ( .A(n3473), .B(n3472), .ZN(n3478) );
  INV_X1 U4234 ( .A(n3955), .ZN(n3476) );
  INV_X1 U4235 ( .A(n3984), .ZN(n3947) );
  OAI22_X1 U4236 ( .A1(n3947), .A2(n3623), .B1(n3624), .B2(n3954), .ZN(n3475)
         );
  OAI22_X1 U4237 ( .A1(n3946), .A2(n3626), .B1(STATE_REG_SCAN_IN), .B2(n4777), 
        .ZN(n3474) );
  AOI211_X1 U4238 ( .C1(n3476), .C2(n3614), .A(n3475), .B(n3474), .ZN(n3477)
         );
  OAI21_X1 U4239 ( .B1(n3478), .B2(n3616), .A(n3477), .ZN(U3211) );
  AOI21_X1 U4240 ( .B1(n3480), .B2(n3482), .A(n3481), .ZN(n3483) );
  NOR3_X1 U4241 ( .A1(n3479), .A2(n3483), .A3(n3616), .ZN(n3487) );
  AOI22_X1 U4242 ( .A1(n3588), .A2(n3921), .B1(n3586), .B2(n4063), .ZN(n3485)
         );
  AOI22_X1 U4243 ( .A1(n4023), .A2(n3583), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3484) );
  OAI211_X1 U4244 ( .C1(n3631), .C2(n4031), .A(n3485), .B(n3484), .ZN(n3486)
         );
  OR2_X1 U4245 ( .A1(n3487), .A2(n3486), .ZN(U3213) );
  XNOR2_X1 U4246 ( .A(n3488), .B(n3489), .ZN(n3490) );
  NAND2_X1 U4247 ( .A1(n3490), .A2(n3621), .ZN(n3494) );
  OAI22_X1 U4248 ( .A1(n3624), .A2(n4116), .B1(n4114), .B2(n3623), .ZN(n3492)
         );
  NAND2_X1 U4249 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3848) );
  OAI21_X1 U4250 ( .B1(n4066), .B2(n3626), .A(n3848), .ZN(n3491) );
  NOR2_X1 U4251 ( .A1(n3492), .A2(n3491), .ZN(n3493) );
  OAI211_X1 U4252 ( .C1(n3631), .C2(n4117), .A(n3494), .B(n3493), .ZN(U3216)
         );
  XNOR2_X1 U4253 ( .A(n3496), .B(n3495), .ZN(n3497) );
  XNOR2_X1 U4254 ( .A(n3498), .B(n3497), .ZN(n3499) );
  NAND2_X1 U4255 ( .A1(n3499), .A2(n3621), .ZN(n3504) );
  INV_X1 U4256 ( .A(n4062), .ZN(n4069) );
  OAI22_X1 U4257 ( .A1(n3624), .A2(n4069), .B1(n4066), .B2(n3623), .ZN(n3502)
         );
  INV_X1 U4258 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3500) );
  OAI22_X1 U4259 ( .A1(n4021), .A2(n3626), .B1(STATE_REG_SCAN_IN), .B2(n3500), 
        .ZN(n3501) );
  NOR2_X1 U4260 ( .A1(n3502), .A2(n3501), .ZN(n3503) );
  OAI211_X1 U4261 ( .C1(n3631), .C2(n4071), .A(n3504), .B(n3503), .ZN(U3220)
         );
  INV_X1 U4262 ( .A(n3506), .ZN(n3507) );
  NOR2_X1 U4263 ( .A1(n3508), .A2(n3507), .ZN(n3509) );
  XNOR2_X1 U4264 ( .A(n3505), .B(n3509), .ZN(n3515) );
  INV_X1 U4265 ( .A(n3510), .ZN(n3991) );
  OAI22_X1 U4266 ( .A1(n3987), .A2(n3623), .B1(n3624), .B2(n3990), .ZN(n3513)
         );
  INV_X1 U4267 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3511) );
  OAI22_X1 U4268 ( .A1(n3947), .A2(n3626), .B1(STATE_REG_SCAN_IN), .B2(n3511), 
        .ZN(n3512) );
  AOI211_X1 U4269 ( .C1(n3991), .C2(n3614), .A(n3513), .B(n3512), .ZN(n3514)
         );
  OAI21_X1 U4270 ( .B1(n3515), .B2(n3616), .A(n3514), .ZN(U3222) );
  AOI21_X1 U4271 ( .B1(n3619), .B2(n3516), .A(n2146), .ZN(n3517) );
  XOR2_X1 U4272 ( .A(n3518), .B(n3517), .Z(n3519) );
  NAND2_X1 U4273 ( .A1(n3519), .A2(n3621), .ZN(n3523) );
  OAI22_X1 U4274 ( .A1(n3624), .A2(n3892), .B1(n4168), .B2(n3623), .ZN(n3521)
         );
  NAND2_X1 U4275 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4435) );
  OAI21_X1 U4276 ( .B1(n4130), .B2(n3626), .A(n4435), .ZN(n3520) );
  NOR2_X1 U4277 ( .A1(n3521), .A2(n3520), .ZN(n3522) );
  OAI211_X1 U4278 ( .C1(n3631), .C2(n4173), .A(n3523), .B(n3522), .ZN(U3223)
         );
  XNOR2_X1 U4279 ( .A(n3526), .B(n3525), .ZN(n3527) );
  XNOR2_X1 U4280 ( .A(n3524), .B(n3527), .ZN(n3528) );
  NAND2_X1 U4281 ( .A1(n3528), .A2(n3621), .ZN(n3533) );
  OAI22_X1 U4282 ( .A1(n3624), .A2(n4155), .B1(n4152), .B2(n3623), .ZN(n3531)
         );
  AND2_X1 U4283 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4448) );
  INV_X1 U4284 ( .A(n4448), .ZN(n3529) );
  OAI21_X1 U4285 ( .B1(n4114), .B2(n3626), .A(n3529), .ZN(n3530) );
  NOR2_X1 U4286 ( .A1(n3531), .A2(n3530), .ZN(n3532) );
  OAI211_X1 U4287 ( .C1(n3631), .C2(n4157), .A(n3533), .B(n3532), .ZN(U3225)
         );
  NAND2_X1 U4288 ( .A1(n3535), .A2(n3534), .ZN(n3536) );
  XOR2_X1 U4289 ( .A(n3537), .B(n3536), .Z(n3538) );
  NAND2_X1 U4290 ( .A1(n3538), .A2(n3621), .ZN(n3542) );
  AOI22_X1 U4291 ( .A1(n4005), .A2(n3583), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3541) );
  AOI22_X1 U4292 ( .A1(n3588), .A2(n4006), .B1(n4044), .B2(n3586), .ZN(n3540)
         );
  NAND2_X1 U4293 ( .A1(n3614), .A2(n3998), .ZN(n3539) );
  NAND4_X1 U4294 ( .A1(n3542), .A2(n3541), .A3(n3540), .A4(n3539), .ZN(U3226)
         );
  NAND2_X1 U4295 ( .A1(n3544), .A2(n3543), .ZN(n3546) );
  NAND2_X1 U4296 ( .A1(n3546), .A2(n3545), .ZN(n3548) );
  XNOR2_X1 U4297 ( .A(n3548), .B(n3547), .ZN(n3549) );
  NAND2_X1 U4298 ( .A1(n3549), .A2(n3621), .ZN(n3557) );
  AOI21_X1 U4299 ( .B1(n3779), .B2(n3586), .A(n3550), .ZN(n3556) );
  AOI22_X1 U4300 ( .A1(n3588), .A2(n3551), .B1(n3583), .B2(n3585), .ZN(n3555)
         );
  INV_X1 U4301 ( .A(n3552), .ZN(n3553) );
  NAND2_X1 U4302 ( .A1(n3614), .A2(n3553), .ZN(n3554) );
  NAND4_X1 U4303 ( .A1(n3557), .A2(n3556), .A3(n3555), .A4(n3554), .ZN(U3228)
         );
  OAI21_X1 U4304 ( .B1(n3561), .B2(n3559), .A(n3558), .ZN(n3560) );
  OAI21_X1 U4305 ( .B1(n2150), .B2(n3561), .A(n3560), .ZN(n3562) );
  NAND2_X1 U4306 ( .A1(n3562), .A2(n3621), .ZN(n3567) );
  OAI22_X1 U4307 ( .A1(n3624), .A2(n4091), .B1(n4129), .B2(n3623), .ZN(n3565)
         );
  INV_X1 U4308 ( .A(n4084), .ZN(n4048) );
  INV_X1 U4309 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3563) );
  OAI22_X1 U4310 ( .A1(n4048), .A2(n3626), .B1(STATE_REG_SCAN_IN), .B2(n3563), 
        .ZN(n3564) );
  NOR2_X1 U4311 ( .A1(n3565), .A2(n3564), .ZN(n3566) );
  OAI211_X1 U4312 ( .C1(n3631), .C2(n4093), .A(n3567), .B(n3566), .ZN(U3230)
         );
  OAI21_X1 U4313 ( .B1(n3569), .B2(n3568), .A(n3480), .ZN(n3570) );
  NAND2_X1 U4314 ( .A1(n3570), .A2(n3621), .ZN(n3577) );
  NOR2_X1 U4315 ( .A1(n3571), .A2(STATE_REG_SCAN_IN), .ZN(n3572) );
  AOI21_X1 U4316 ( .B1(n4044), .B2(n3583), .A(n3572), .ZN(n3576) );
  AOI22_X1 U4317 ( .A1(n3588), .A2(n4045), .B1(n3586), .B2(n4084), .ZN(n3575)
         );
  INV_X1 U4318 ( .A(n3573), .ZN(n4051) );
  NAND2_X1 U4319 ( .A1(n3614), .A2(n4051), .ZN(n3574) );
  NAND4_X1 U4320 ( .A1(n3577), .A2(n3576), .A3(n3575), .A4(n3574), .ZN(U3232)
         );
  XNOR2_X1 U4321 ( .A(n3579), .B(n3578), .ZN(n3580) );
  XNOR2_X1 U4322 ( .A(n3581), .B(n3580), .ZN(n3582) );
  NAND2_X1 U4323 ( .A1(n3582), .A2(n3621), .ZN(n3594) );
  NOR2_X1 U4324 ( .A1(STATE_REG_SCAN_IN), .A2(n4775), .ZN(n4385) );
  AOI21_X1 U4325 ( .B1(n3584), .B2(n3583), .A(n4385), .ZN(n3593) );
  AOI22_X1 U4326 ( .A1(n3588), .A2(n3587), .B1(n3586), .B2(n3585), .ZN(n3592)
         );
  INV_X1 U4327 ( .A(n3589), .ZN(n3590) );
  NAND2_X1 U4328 ( .A1(n3614), .A2(n3590), .ZN(n3591) );
  NAND4_X1 U4329 ( .A1(n3594), .A2(n3593), .A3(n3592), .A4(n3591), .ZN(U3233)
         );
  INV_X1 U4330 ( .A(n3595), .ZN(n3597) );
  NAND2_X1 U4331 ( .A1(n3597), .A2(n3596), .ZN(n3598) );
  XNOR2_X1 U4332 ( .A(n3599), .B(n3598), .ZN(n3600) );
  NAND2_X1 U4333 ( .A1(n3600), .A2(n3621), .ZN(n3605) );
  OAI22_X1 U4334 ( .A1(n3624), .A2(n3896), .B1(n4130), .B2(n3623), .ZN(n3603)
         );
  AND2_X1 U4335 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4463) );
  INV_X1 U4336 ( .A(n4463), .ZN(n3601) );
  OAI21_X1 U4337 ( .B1(n4129), .B2(n3626), .A(n3601), .ZN(n3602) );
  NOR2_X1 U4338 ( .A1(n3603), .A2(n3602), .ZN(n3604) );
  OAI211_X1 U4339 ( .C1(n3631), .C2(n4138), .A(n3605), .B(n3604), .ZN(U3235)
         );
  INV_X1 U4340 ( .A(n3607), .ZN(n3609) );
  NAND2_X1 U4341 ( .A1(n3609), .A2(n3608), .ZN(n3610) );
  XNOR2_X1 U4342 ( .A(n3606), .B(n3610), .ZN(n3617) );
  INV_X1 U4343 ( .A(n3611), .ZN(n3974) );
  INV_X1 U4344 ( .A(n4005), .ZN(n3966) );
  OAI22_X1 U4345 ( .A1(n3966), .A2(n3623), .B1(n3624), .B2(n3973), .ZN(n3613)
         );
  INV_X1 U4346 ( .A(REG3_REG_26__SCAN_IN), .ZN(n4771) );
  OAI22_X1 U4347 ( .A1(n3935), .A2(n3626), .B1(STATE_REG_SCAN_IN), .B2(n4771), 
        .ZN(n3612) );
  AOI211_X1 U4348 ( .C1(n3974), .C2(n3614), .A(n3613), .B(n3612), .ZN(n3615)
         );
  OAI21_X1 U4349 ( .B1(n3617), .B2(n3616), .A(n3615), .ZN(U3237) );
  INV_X1 U4350 ( .A(n3516), .ZN(n3618) );
  NOR2_X1 U4351 ( .A1(n2146), .A2(n3618), .ZN(n3620) );
  XNOR2_X1 U4352 ( .A(n3620), .B(n3619), .ZN(n3622) );
  NAND2_X1 U4353 ( .A1(n3622), .A2(n3621), .ZN(n3630) );
  OAI22_X1 U4354 ( .A1(n3624), .A2(n4193), .B1(n4192), .B2(n3623), .ZN(n3628)
         );
  AND2_X1 U4355 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4428) );
  INV_X1 U4356 ( .A(n4428), .ZN(n3625) );
  OAI21_X1 U4357 ( .B1(n4152), .B2(n3626), .A(n3625), .ZN(n3627) );
  NOR2_X1 U4358 ( .A1(n3628), .A2(n3627), .ZN(n3629) );
  OAI211_X1 U4359 ( .C1(n3631), .C2(n4197), .A(n3630), .B(n3629), .ZN(U3238)
         );
  INV_X1 U4360 ( .A(n4217), .ZN(n4204) );
  NAND2_X1 U4361 ( .A1(n3297), .A2(REG1_REG_31__SCAN_IN), .ZN(n3637) );
  NAND2_X1 U4362 ( .A1(n3632), .A2(REG2_REG_31__SCAN_IN), .ZN(n3636) );
  INV_X1 U4363 ( .A(REG0_REG_31__SCAN_IN), .ZN(n3633) );
  OR2_X1 U4364 ( .A1(n3634), .A2(n3633), .ZN(n3635) );
  INV_X1 U4365 ( .A(n4180), .ZN(n3854) );
  NOR2_X1 U4366 ( .A1(n3638), .A2(n3854), .ZN(n3640) );
  NAND2_X1 U4367 ( .A1(n3890), .A2(n4193), .ZN(n3856) );
  NAND2_X1 U4368 ( .A1(n3856), .A2(n3639), .ZN(n3739) );
  NAND2_X1 U4369 ( .A1(n4152), .A2(n4172), .ZN(n3746) );
  NAND2_X1 U4370 ( .A1(n4168), .A2(n4186), .ZN(n3738) );
  OAI211_X1 U4371 ( .C1(n3640), .C2(n3739), .A(n3746), .B(n3738), .ZN(n3642)
         );
  NAND2_X1 U4372 ( .A1(n4149), .A2(n3896), .ZN(n4104) );
  INV_X1 U4373 ( .A(n4129), .ZN(n3898) );
  NAND2_X1 U4374 ( .A1(n3898), .A2(n4116), .ZN(n3641) );
  AND2_X1 U4375 ( .A1(n4111), .A2(n4091), .ZN(n3862) );
  INV_X1 U4376 ( .A(n3862), .ZN(n3646) );
  NAND2_X1 U4377 ( .A1(n4166), .A2(n4155), .ZN(n3860) );
  AND3_X1 U4378 ( .A1(n3861), .A2(n3646), .A3(n3860), .ZN(n3749) );
  INV_X1 U4379 ( .A(n4152), .ZN(n4188) );
  NAND2_X1 U4380 ( .A1(n4188), .A2(n3892), .ZN(n3745) );
  NAND3_X1 U4381 ( .A1(n3642), .A2(n3749), .A3(n3745), .ZN(n3648) );
  NAND2_X1 U4382 ( .A1(n4114), .A2(n3895), .ZN(n4106) );
  NAND2_X1 U4383 ( .A1(n4130), .A2(n4148), .ZN(n4101) );
  NAND2_X1 U4384 ( .A1(n4106), .A2(n4101), .ZN(n3643) );
  NAND2_X1 U4385 ( .A1(n3643), .A2(n3861), .ZN(n3645) );
  NAND2_X1 U4386 ( .A1(n4129), .A2(n4110), .ZN(n3644) );
  NAND2_X1 U4387 ( .A1(n3645), .A2(n3644), .ZN(n4078) );
  NOR2_X1 U4388 ( .A1(n4111), .A2(n4091), .ZN(n3647) );
  OAI21_X1 U4389 ( .B1(n4078), .B2(n3647), .A(n3646), .ZN(n4016) );
  NAND2_X1 U4390 ( .A1(n4021), .A2(n4045), .ZN(n4018) );
  NAND2_X1 U4391 ( .A1(n4048), .A2(n4062), .ZN(n4017) );
  AND2_X1 U4392 ( .A1(n4018), .A2(n4017), .ZN(n3752) );
  AND2_X1 U4393 ( .A1(n4016), .A2(n3752), .ZN(n3866) );
  NAND2_X1 U4394 ( .A1(n3648), .A2(n3866), .ZN(n3649) );
  AND2_X1 U4395 ( .A1(n4084), .A2(n4069), .ZN(n3753) );
  NAND2_X1 U4396 ( .A1(n4018), .A2(n3753), .ZN(n3863) );
  OR2_X1 U4397 ( .A1(n4023), .A2(n3905), .ZN(n3667) );
  OR2_X1 U4398 ( .A1(n4044), .A2(n4029), .ZN(n4000) );
  NAND2_X1 U4399 ( .A1(n3667), .A2(n4000), .ZN(n3868) );
  AOI21_X1 U4400 ( .B1(n3649), .B2(n3863), .A(n3868), .ZN(n3651) );
  NAND2_X1 U4401 ( .A1(n4044), .A2(n4029), .ZN(n3686) );
  NAND2_X1 U4402 ( .A1(n4063), .A2(n4052), .ZN(n3672) );
  AND2_X1 U4403 ( .A1(n3686), .A2(n3672), .ZN(n3864) );
  NAND2_X1 U4404 ( .A1(n4005), .A2(n3990), .ZN(n3869) );
  NAND2_X1 U4405 ( .A1(n4023), .A2(n3905), .ZN(n3867) );
  OAI211_X1 U4406 ( .C1(n3864), .C2(n3868), .A(n3869), .B(n3867), .ZN(n3699)
         );
  NAND2_X1 U4407 ( .A1(n3947), .A2(n3677), .ZN(n3650) );
  OR2_X1 U4408 ( .A1(n4005), .A2(n3990), .ZN(n3961) );
  AND2_X1 U4409 ( .A1(n3650), .A2(n3961), .ZN(n3755) );
  NOR2_X1 U4410 ( .A1(n3876), .A2(n3874), .ZN(n3658) );
  OAI211_X1 U4411 ( .C1(n3651), .C2(n3699), .A(n3755), .B(n3658), .ZN(n3661)
         );
  INV_X1 U4412 ( .A(n3923), .ZN(n3652) );
  OR2_X1 U4413 ( .A1(n3932), .A2(n3652), .ZN(n3654) );
  OR2_X1 U4414 ( .A1(n3881), .A2(n4204), .ZN(n3653) );
  AND2_X1 U4415 ( .A1(n3349), .A2(DATAI_31_), .ZN(n4208) );
  INV_X1 U4416 ( .A(n4208), .ZN(n4205) );
  NAND2_X1 U4417 ( .A1(n4207), .A2(n4205), .ZN(n3761) );
  AND2_X1 U4418 ( .A1(n3653), .A2(n3761), .ZN(n3680) );
  AND2_X1 U4419 ( .A1(n3654), .A2(n3680), .ZN(n3657) );
  INV_X1 U4420 ( .A(n3657), .ZN(n3660) );
  INV_X1 U4421 ( .A(n3932), .ZN(n3656) );
  NAND2_X1 U4422 ( .A1(n3916), .A2(n3655), .ZN(n3877) );
  OAI21_X1 U4423 ( .B1(n3656), .B2(n3923), .A(n3877), .ZN(n3758) );
  OAI21_X1 U4424 ( .B1(n3658), .B2(n3758), .A(n3657), .ZN(n3764) );
  AND2_X1 U4425 ( .A1(n3984), .A2(n3973), .ZN(n3871) );
  NOR2_X1 U4426 ( .A1(n3935), .A2(n3913), .ZN(n3760) );
  NOR2_X1 U4427 ( .A1(n3760), .A2(n3874), .ZN(n3952) );
  INV_X1 U4428 ( .A(n3952), .ZN(n3944) );
  NOR3_X1 U4429 ( .A1(n3871), .A2(n3944), .A3(n3758), .ZN(n3659) );
  OAI22_X1 U4430 ( .A1(n3661), .A2(n3660), .B1(n3764), .B2(n3659), .ZN(n3662)
         );
  OAI21_X1 U4431 ( .B1(n4204), .B2(n4207), .A(n3662), .ZN(n3665) );
  INV_X1 U4432 ( .A(n3881), .ZN(n3663) );
  NOR2_X1 U4433 ( .A1(n3663), .A2(n4217), .ZN(n3678) );
  OAI21_X1 U4434 ( .B1(n3678), .B2(n3679), .A(n4208), .ZN(n3664) );
  NAND2_X1 U4435 ( .A1(n3665), .A2(n3664), .ZN(n3698) );
  INV_X1 U4436 ( .A(n3876), .ZN(n3666) );
  NAND2_X1 U4437 ( .A1(n3666), .A2(n3877), .ZN(n3930) );
  INV_X1 U4438 ( .A(n3930), .ZN(n3927) );
  NAND2_X1 U4439 ( .A1(n3667), .A2(n3867), .ZN(n3997) );
  INV_X1 U4440 ( .A(n3997), .ZN(n4003) );
  INV_X1 U4441 ( .A(n3753), .ZN(n3668) );
  NAND4_X1 U4442 ( .A1(n3927), .A2(n3716), .A3(n4003), .A4(n4060), .ZN(n3676)
         );
  NAND2_X1 U4443 ( .A1(n3738), .A2(n3856), .ZN(n4178) );
  INV_X1 U4444 ( .A(n4178), .ZN(n4182) );
  NAND4_X1 U4445 ( .A1(n3671), .A2(n4182), .A3(n3670), .A4(n3669), .ZN(n3675)
         );
  NAND2_X1 U4446 ( .A1(n4018), .A2(n3672), .ZN(n4038) );
  INV_X1 U4447 ( .A(n4038), .ZN(n4040) );
  NAND2_X1 U4448 ( .A1(n3746), .A2(n3745), .ZN(n4164) );
  INV_X1 U4449 ( .A(n4164), .ZN(n3859) );
  NAND4_X1 U4450 ( .A1(n4040), .A2(n2274), .A3(n3859), .A4(n3673), .ZN(n3674)
         );
  NOR3_X1 U4451 ( .A1(n3676), .A2(n3675), .A3(n3674), .ZN(n3695) );
  NAND2_X1 U4452 ( .A1(n3947), .A2(n3973), .ZN(n3909) );
  NAND2_X1 U4453 ( .A1(n2166), .A2(n3909), .ZN(n3964) );
  NOR2_X1 U4454 ( .A1(n4066), .A2(n4091), .ZN(n3900) );
  NOR2_X1 U4455 ( .A1(n3900), .A2(n2158), .ZN(n4082) );
  NAND2_X1 U4456 ( .A1(n4106), .A2(n4104), .ZN(n4125) );
  XNOR2_X1 U4457 ( .A(n4129), .B(n4110), .ZN(n4108) );
  NAND2_X1 U4458 ( .A1(n4101), .A2(n3860), .ZN(n4146) );
  NOR4_X1 U4459 ( .A1(n4082), .A2(n4125), .A3(n4108), .A4(n4146), .ZN(n3682)
         );
  XNOR2_X1 U4460 ( .A(n3932), .B(n3923), .ZN(n3919) );
  AOI21_X1 U4461 ( .B1(n4208), .B2(n3679), .A(n3678), .ZN(n3765) );
  AND4_X1 U4462 ( .A1(n3919), .A2(n3952), .A3(n3765), .A4(n3680), .ZN(n3681)
         );
  NAND4_X1 U4463 ( .A1(n3964), .A2(n3683), .A3(n3682), .A4(n3681), .ZN(n3685)
         );
  NAND2_X1 U4464 ( .A1(n3869), .A2(n3961), .ZN(n3980) );
  NOR3_X1 U4465 ( .A1(n3685), .A2(n3980), .A3(n3684), .ZN(n3694) );
  NAND2_X1 U4466 ( .A1(n4000), .A2(n3686), .ZN(n4019) );
  NOR4_X1 U4467 ( .A1(n4019), .A2(n3689), .A3(n3688), .A4(n3687), .ZN(n3693)
         );
  INV_X1 U4468 ( .A(n2362), .ZN(n3691) );
  AND4_X1 U4469 ( .A1(n3691), .A2(n3690), .A3(n2801), .A4(n2849), .ZN(n3692)
         );
  NAND4_X1 U4470 ( .A1(n3695), .A2(n3694), .A3(n3693), .A4(n3692), .ZN(n3697)
         );
  MUX2_X1 U4471 ( .A(n3698), .B(n3697), .S(n3696), .Z(n3769) );
  INV_X1 U4472 ( .A(n3699), .ZN(n3757) );
  INV_X1 U4473 ( .A(n3700), .ZN(n3704) );
  OAI211_X1 U4474 ( .C1(n3704), .C2(n3703), .A(n3702), .B(n3701), .ZN(n3707)
         );
  NAND3_X1 U4475 ( .A1(n3707), .A2(n3706), .A3(n3705), .ZN(n3710) );
  NAND3_X1 U4476 ( .A1(n3710), .A2(n3709), .A3(n3708), .ZN(n3712) );
  NAND3_X1 U4477 ( .A1(n3712), .A2(n2859), .A3(n3711), .ZN(n3714) );
  NAND4_X1 U4478 ( .A1(n3714), .A2(n2862), .A3(n3725), .A4(n3713), .ZN(n3717)
         );
  NAND3_X1 U4479 ( .A1(n3717), .A2(n3716), .A3(n3715), .ZN(n3718) );
  NAND3_X1 U4480 ( .A1(n3718), .A2(n3722), .A3(n3726), .ZN(n3721) );
  AND3_X1 U4481 ( .A1(n3721), .A2(n3720), .A3(n3719), .ZN(n3732) );
  INV_X1 U4482 ( .A(n3722), .ZN(n3724) );
  NOR2_X1 U4483 ( .A1(n3724), .A2(n3723), .ZN(n3728) );
  NAND4_X1 U4484 ( .A1(n3728), .A2(n3727), .A3(n3726), .A4(n3725), .ZN(n3729)
         );
  OAI211_X1 U4485 ( .C1(n3732), .C2(n3731), .A(n3730), .B(n3729), .ZN(n3744)
         );
  INV_X1 U4486 ( .A(n3733), .ZN(n3737) );
  INV_X1 U4487 ( .A(n3734), .ZN(n3735) );
  NOR4_X1 U4488 ( .A1(n3737), .A2(n3736), .A3(n3739), .A4(n3735), .ZN(n3743)
         );
  INV_X1 U4489 ( .A(n3738), .ZN(n3742) );
  AOI21_X1 U4490 ( .B1(n3740), .B2(n4180), .A(n3739), .ZN(n3741) );
  AOI211_X1 U4491 ( .C1(n3744), .C2(n3743), .A(n3742), .B(n3741), .ZN(n3747)
         );
  INV_X1 U4492 ( .A(n3745), .ZN(n3858) );
  OAI21_X1 U4493 ( .B1(n3747), .B2(n3858), .A(n3746), .ZN(n3750) );
  INV_X1 U4494 ( .A(n4016), .ZN(n3748) );
  AOI21_X1 U4495 ( .B1(n3750), .B2(n3749), .A(n3748), .ZN(n3754) );
  INV_X1 U4496 ( .A(n3868), .ZN(n3751) );
  OAI211_X1 U4497 ( .C1(n3754), .C2(n3753), .A(n3752), .B(n3751), .ZN(n3756)
         );
  INV_X1 U4498 ( .A(n3755), .ZN(n3873) );
  AOI21_X1 U4499 ( .B1(n3757), .B2(n3756), .A(n3873), .ZN(n3759) );
  NOR4_X1 U4500 ( .A1(n3760), .A2(n3871), .A3(n3759), .A4(n3758), .ZN(n3766)
         );
  INV_X1 U4501 ( .A(n3765), .ZN(n3762) );
  NAND2_X1 U4502 ( .A1(n3762), .A2(n3761), .ZN(n3763) );
  AOI22_X1 U4503 ( .A1(n3766), .A2(n3765), .B1(n3764), .B2(n3763), .ZN(n3768)
         );
  MUX2_X1 U4504 ( .A(n3769), .B(n3768), .S(n3767), .Z(n3770) );
  XNOR2_X1 U4505 ( .A(n3770), .B(n3849), .ZN(n3777) );
  NAND2_X1 U4506 ( .A1(n3772), .A2(n3771), .ZN(n3773) );
  OAI211_X1 U4507 ( .C1(n3774), .C2(n3776), .A(n3773), .B(B_REG_SCAN_IN), .ZN(
        n3775) );
  OAI21_X1 U4508 ( .B1(n3777), .B2(n3776), .A(n3775), .ZN(U3239) );
  MUX2_X1 U4509 ( .A(n4207), .B(DATAO_REG_31__SCAN_IN), .S(n3783), .Z(U3581)
         );
  MUX2_X1 U4510 ( .A(DATAO_REG_29__SCAN_IN), .B(n3932), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4511 ( .A(n3916), .B(DATAO_REG_28__SCAN_IN), .S(n3783), .Z(U3578)
         );
  INV_X1 U4512 ( .A(n3935), .ZN(n3968) );
  MUX2_X1 U4513 ( .A(n3968), .B(DATAO_REG_27__SCAN_IN), .S(n3783), .Z(U3577)
         );
  MUX2_X1 U4514 ( .A(n3984), .B(DATAO_REG_26__SCAN_IN), .S(n3783), .Z(U3576)
         );
  MUX2_X1 U4515 ( .A(DATAO_REG_23__SCAN_IN), .B(n4044), .S(U4043), .Z(U3573)
         );
  MUX2_X1 U4516 ( .A(n4063), .B(DATAO_REG_22__SCAN_IN), .S(n3783), .Z(U3572)
         );
  MUX2_X1 U4517 ( .A(n4084), .B(DATAO_REG_21__SCAN_IN), .S(n3783), .Z(U3571)
         );
  MUX2_X1 U4518 ( .A(DATAO_REG_19__SCAN_IN), .B(n3898), .S(U4043), .Z(U3569)
         );
  MUX2_X1 U4519 ( .A(DATAO_REG_18__SCAN_IN), .B(n4149), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4520 ( .A(DATAO_REG_16__SCAN_IN), .B(n4188), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4521 ( .A(DATAO_REG_14__SCAN_IN), .B(n3888), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4522 ( .A(DATAO_REG_13__SCAN_IN), .B(n3778), .S(U4043), .Z(U3563)
         );
  MUX2_X1 U4523 ( .A(DATAO_REG_8__SCAN_IN), .B(n3779), .S(U4043), .Z(U3558) );
  MUX2_X1 U4524 ( .A(DATAO_REG_7__SCAN_IN), .B(n3780), .S(U4043), .Z(U3557) );
  MUX2_X1 U4525 ( .A(n3781), .B(DATAO_REG_6__SCAN_IN), .S(n3783), .Z(U3556) );
  MUX2_X1 U4526 ( .A(DATAO_REG_2__SCAN_IN), .B(n3782), .S(U4043), .Z(U3552) );
  MUX2_X1 U4527 ( .A(n2580), .B(DATAO_REG_0__SCAN_IN), .S(n3783), .Z(U3550) );
  NAND2_X1 U4528 ( .A1(n4422), .A2(n4356), .ZN(n3793) );
  AOI22_X1 U4529 ( .A1(n4464), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3792) );
  OAI211_X1 U4530 ( .C1(n3786), .C2(n3785), .A(n4472), .B(n3784), .ZN(n3791)
         );
  XOR2_X1 U4531 ( .A(n3788), .B(n3787), .Z(n3789) );
  NAND2_X1 U4532 ( .A1(n4457), .A2(n3789), .ZN(n3790) );
  NAND4_X1 U4533 ( .A1(n3793), .A2(n3792), .A3(n3791), .A4(n3790), .ZN(U3241)
         );
  NAND2_X1 U4534 ( .A1(U3149), .A2(REG3_REG_2__SCAN_IN), .ZN(n3795) );
  NAND2_X1 U4535 ( .A1(n4464), .A2(ADDR_REG_2__SCAN_IN), .ZN(n3794) );
  OAI211_X1 U4536 ( .C1(n4475), .C2(n3796), .A(n3795), .B(n3794), .ZN(n3797)
         );
  INV_X1 U4537 ( .A(n3797), .ZN(n3807) );
  INV_X1 U4538 ( .A(n3798), .ZN(n3799) );
  XNOR2_X1 U4539 ( .A(n3800), .B(n3799), .ZN(n3801) );
  NAND2_X1 U4540 ( .A1(n4457), .A2(n3801), .ZN(n3806) );
  OAI211_X1 U4541 ( .C1(n3804), .C2(n3803), .A(n4472), .B(n3802), .ZN(n3805)
         );
  NAND4_X1 U4542 ( .A1(n3808), .A2(n3807), .A3(n3806), .A4(n3805), .ZN(U3242)
         );
  INV_X1 U4543 ( .A(n3844), .ZN(n4489) );
  INV_X1 U4544 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4680) );
  AOI22_X1 U4545 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4489), .B1(n3844), .B2(
        n4680), .ZN(n4461) );
  INV_X1 U4546 ( .A(n3826), .ZN(n4498) );
  NOR2_X1 U4547 ( .A1(n3810), .A2(n4498), .ZN(n3811) );
  INV_X1 U4548 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4375) );
  NOR2_X1 U4549 ( .A1(n4375), .A2(n4374), .ZN(n4373) );
  INV_X1 U4550 ( .A(n3830), .ZN(n4496) );
  AOI22_X1 U4551 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4496), .B1(n3830), .B2(
        n4677), .ZN(n4383) );
  NOR2_X1 U4552 ( .A1(n3812), .A2(n4495), .ZN(n3813) );
  INV_X1 U4553 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4395) );
  INV_X1 U4554 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4284) );
  AOI22_X1 U4555 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4494), .B1(n4407), .B2(
        n4284), .ZN(n4403) );
  NOR2_X1 U4556 ( .A1(n4404), .A2(n4403), .ZN(n4402) );
  AND2_X1 U4557 ( .A1(n4407), .A2(REG1_REG_13__SCAN_IN), .ZN(n3814) );
  INV_X1 U4558 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4414) );
  INV_X1 U4559 ( .A(n3816), .ZN(n3817) );
  INV_X1 U4560 ( .A(n3841), .ZN(n4493) );
  INV_X1 U4561 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4276) );
  AOI22_X1 U4562 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4493), .B1(n3841), .B2(
        n4276), .ZN(n4426) );
  AND2_X1 U4563 ( .A1(n3841), .A2(REG1_REG_15__SCAN_IN), .ZN(n3818) );
  INV_X1 U4564 ( .A(n3820), .ZN(n3819) );
  NAND2_X1 U4565 ( .A1(n3819), .A2(n4491), .ZN(n3821) );
  INV_X1 U4566 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4439) );
  NAND2_X1 U4567 ( .A1(n3821), .A2(n4438), .ZN(n4450) );
  INV_X1 U4568 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4678) );
  AOI22_X1 U4569 ( .A1(n3843), .A2(REG1_REG_17__SCAN_IN), .B1(n4678), .B2(
        n4490), .ZN(n4451) );
  NAND2_X1 U4570 ( .A1(n4450), .A2(n4451), .ZN(n4449) );
  NAND2_X1 U4571 ( .A1(REG2_REG_18__SCAN_IN), .A2(n3844), .ZN(n3822) );
  OAI21_X1 U4572 ( .B1(REG2_REG_18__SCAN_IN), .B2(n3844), .A(n3822), .ZN(n4470) );
  NOR2_X1 U4573 ( .A1(n3843), .A2(REG2_REG_17__SCAN_IN), .ZN(n3823) );
  AOI21_X1 U4574 ( .B1(REG2_REG_17__SCAN_IN), .B2(n3843), .A(n3823), .ZN(n4454) );
  INV_X1 U4575 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4696) );
  NAND2_X1 U4576 ( .A1(n3826), .A2(n3827), .ZN(n3828) );
  INV_X1 U4577 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3829) );
  AOI22_X1 U4578 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3830), .B1(n4496), .B2(
        n3829), .ZN(n4389) );
  NAND2_X1 U4579 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3830), .ZN(n3831) );
  NAND2_X1 U4580 ( .A1(n3832), .A2(n3833), .ZN(n3834) );
  NAND2_X1 U4581 ( .A1(n3243), .A2(n4494), .ZN(n3835) );
  INV_X1 U4582 ( .A(n4421), .ZN(n3836) );
  NAND2_X1 U4583 ( .A1(n3837), .A2(n3836), .ZN(n3838) );
  INV_X1 U4584 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4585 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4493), .B1(n3841), .B2(
        n3840), .ZN(n4431) );
  NAND2_X1 U4586 ( .A1(n2131), .A2(n4491), .ZN(n3842) );
  INV_X1 U4587 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4442) );
  INV_X1 U4588 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4699) );
  MUX2_X1 U4589 ( .A(n4699), .B(REG2_REG_19__SCAN_IN), .S(n3849), .Z(n3845) );
  XNOR2_X1 U4590 ( .A(n3846), .B(n3845), .ZN(n3851) );
  NAND2_X1 U4591 ( .A1(n4464), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3847) );
  OAI211_X1 U4592 ( .C1(n4475), .C2(n3849), .A(n3848), .B(n3847), .ZN(n3850)
         );
  AOI21_X1 U4593 ( .B1(n3851), .B2(n4472), .A(n3850), .ZN(n3852) );
  INV_X1 U4594 ( .A(n3853), .ZN(n3886) );
  NOR2_X1 U4595 ( .A1(n4178), .A2(n3854), .ZN(n3855) );
  NAND2_X1 U4596 ( .A1(n4181), .A2(n3855), .ZN(n3857) );
  NAND2_X1 U4597 ( .A1(n3857), .A2(n3856), .ZN(n4165) );
  NAND2_X1 U4598 ( .A1(n4103), .A2(n3861), .ZN(n4080) );
  NAND2_X1 U4599 ( .A1(n3864), .A2(n3863), .ZN(n3865) );
  AOI21_X2 U4600 ( .B1(n2145), .B2(n3866), .A(n3865), .ZN(n4002) );
  OAI21_X1 U4601 ( .B1(n4002), .B2(n3868), .A(n3867), .ZN(n3981) );
  INV_X1 U4602 ( .A(n3869), .ZN(n3870) );
  NOR2_X2 U4603 ( .A1(n3981), .A2(n3870), .ZN(n3963) );
  INV_X1 U4604 ( .A(n3871), .ZN(n3872) );
  OAI21_X2 U4605 ( .B1(n3963), .B2(n3873), .A(n3872), .ZN(n3945) );
  INV_X1 U4606 ( .A(n3874), .ZN(n3875) );
  OAI21_X2 U4607 ( .B1(n3945), .B2(n3944), .A(n3875), .ZN(n3929) );
  AOI21_X1 U4608 ( .B1(n3929), .B2(n3877), .A(n3876), .ZN(n3878) );
  INV_X1 U4609 ( .A(n3878), .ZN(n3879) );
  XNOR2_X1 U4610 ( .A(n3879), .B(n3919), .ZN(n3880) );
  OR2_X1 U4611 ( .A1(n3946), .A2(n4191), .ZN(n3883) );
  AOI21_X1 U4612 ( .B1(B_REG_SCAN_IN), .B2(n4346), .A(n4128), .ZN(n4206) );
  AOI22_X1 U4613 ( .A1(n3881), .A2(n4206), .B1(n4216), .B2(n3923), .ZN(n3882)
         );
  AOI21_X1 U4614 ( .B1(n3886), .B2(n4476), .A(n4222), .ZN(n3926) );
  NAND2_X1 U4615 ( .A1(n3890), .A2(n4186), .ZN(n3891) );
  AOI22_X1 U4616 ( .A1(n4179), .A2(n3891), .B1(n4193), .B2(n4168), .ZN(n4163)
         );
  NAND2_X1 U4617 ( .A1(n4163), .A2(n4164), .ZN(n4162) );
  NAND2_X1 U4618 ( .A1(n4162), .A2(n3893), .ZN(n4144) );
  NAND2_X1 U4619 ( .A1(n4130), .A2(n4155), .ZN(n3894) );
  NAND2_X1 U4620 ( .A1(n3898), .A2(n4110), .ZN(n3899) );
  NAND2_X1 U4621 ( .A1(n4084), .A2(n4062), .ZN(n3902) );
  NOR2_X1 U4622 ( .A1(n4084), .A2(n4062), .ZN(n3901) );
  AOI21_X1 U4623 ( .B1(n4057), .B2(n3902), .A(n3901), .ZN(n4039) );
  NAND2_X1 U4624 ( .A1(n4039), .A2(n4038), .ZN(n4037) );
  NAND2_X1 U4625 ( .A1(n4063), .A2(n4045), .ZN(n3903) );
  INV_X1 U4626 ( .A(n4044), .ZN(n4009) );
  NAND2_X1 U4627 ( .A1(n4023), .A2(n4006), .ZN(n3904) );
  NAND2_X1 U4628 ( .A1(n3987), .A2(n3905), .ZN(n3906) );
  NOR2_X1 U4629 ( .A1(n4005), .A2(n3983), .ZN(n3908) );
  NAND2_X1 U4630 ( .A1(n4005), .A2(n3983), .ZN(n3907) );
  OAI21_X1 U4631 ( .B1(n3979), .B2(n3908), .A(n3907), .ZN(n3960) );
  INV_X1 U4632 ( .A(n3960), .ZN(n3911) );
  AOI21_X1 U4633 ( .B1(n3911), .B2(n2166), .A(n3910), .ZN(n3951) );
  NAND2_X1 U4634 ( .A1(n3951), .A2(n3912), .ZN(n3915) );
  NAND2_X1 U4635 ( .A1(n3968), .A2(n3913), .ZN(n3914) );
  NAND2_X1 U4636 ( .A1(n3915), .A2(n3914), .ZN(n3928) );
  NAND2_X1 U4637 ( .A1(n3928), .A2(n3930), .ZN(n3918) );
  NAND2_X1 U4638 ( .A1(n3916), .A2(n3937), .ZN(n3917) );
  NAND2_X1 U4639 ( .A1(n3918), .A2(n3917), .ZN(n3920) );
  XNOR2_X1 U4640 ( .A(n3920), .B(n3919), .ZN(n4220) );
  NAND2_X1 U4641 ( .A1(n4220), .A2(n3953), .ZN(n3925) );
  NAND2_X1 U4642 ( .A1(n4067), .A2(n4052), .ZN(n4027) );
  INV_X1 U4643 ( .A(n3922), .ZN(n3936) );
  AOI21_X1 U4644 ( .B1(n3923), .B2(n3936), .A(n4211), .ZN(n4221) );
  AOI22_X1 U4645 ( .A1(n4221), .A2(n4479), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4477), .ZN(n3924) );
  OAI211_X1 U4646 ( .C1(n4477), .C2(n3926), .A(n3925), .B(n3924), .ZN(U3354)
         );
  XNOR2_X1 U4647 ( .A(n3928), .B(n3927), .ZN(n4225) );
  INV_X1 U4648 ( .A(n4225), .ZN(n3943) );
  XOR2_X1 U4649 ( .A(n3930), .B(n3929), .Z(n3931) );
  NAND2_X1 U4650 ( .A1(n3931), .A2(n4184), .ZN(n3934) );
  AOI22_X1 U4651 ( .A1(n3932), .A2(n4187), .B1(n4216), .B2(n3937), .ZN(n3933)
         );
  OAI211_X1 U4652 ( .C1(n3935), .C2(n4191), .A(n3934), .B(n3933), .ZN(n4224)
         );
  AOI21_X1 U4653 ( .B1(n3937), .B2(n2144), .A(n3922), .ZN(n4293) );
  INV_X1 U4654 ( .A(n4293), .ZN(n3940) );
  AOI22_X1 U4655 ( .A1(n3938), .A2(n4476), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4477), .ZN(n3939) );
  OAI21_X1 U4656 ( .B1(n3940), .B2(n4195), .A(n3939), .ZN(n3941) );
  AOI21_X1 U4657 ( .B1(n4224), .B2(n4198), .A(n3941), .ZN(n3942) );
  OAI21_X1 U4658 ( .B1(n3943), .B2(n4202), .A(n3942), .ZN(U3262) );
  XNOR2_X1 U4659 ( .A(n3945), .B(n3944), .ZN(n3950) );
  NOR2_X1 U4660 ( .A1(n3946), .A2(n4128), .ZN(n3949) );
  OAI22_X1 U4661 ( .A1(n3947), .A2(n4191), .B1(n4127), .B2(n3954), .ZN(n3948)
         );
  AOI211_X1 U4662 ( .C1(n3950), .C2(n4184), .A(n3949), .B(n3948), .ZN(n4229)
         );
  XNOR2_X1 U4663 ( .A(n3951), .B(n3952), .ZN(n4228) );
  NAND2_X1 U4664 ( .A1(n4228), .A2(n3953), .ZN(n3959) );
  OAI21_X1 U4665 ( .B1(n3971), .B2(n3954), .A(n2144), .ZN(n4231) );
  INV_X1 U4666 ( .A(n4231), .ZN(n3957) );
  OAI22_X1 U4667 ( .A1(n3955), .A2(n4196), .B1(n4707), .B2(n4198), .ZN(n3956)
         );
  AOI21_X1 U4668 ( .B1(n3957), .B2(n4479), .A(n3956), .ZN(n3958) );
  OAI211_X1 U4669 ( .C1(n4229), .C2(n4477), .A(n3959), .B(n3958), .ZN(U3263)
         );
  XNOR2_X1 U4670 ( .A(n3960), .B(n3964), .ZN(n4233) );
  INV_X1 U4671 ( .A(n4233), .ZN(n3978) );
  INV_X1 U4672 ( .A(n3961), .ZN(n3962) );
  NOR2_X1 U4673 ( .A1(n3963), .A2(n3962), .ZN(n3965) );
  XNOR2_X1 U4674 ( .A(n3965), .B(n3964), .ZN(n3970) );
  OAI22_X1 U4675 ( .A1(n3966), .A2(n4191), .B1(n4127), .B2(n3973), .ZN(n3967)
         );
  AOI21_X1 U4676 ( .B1(n4187), .B2(n3968), .A(n3967), .ZN(n3969) );
  OAI21_X1 U4677 ( .B1(n3970), .B2(n4025), .A(n3969), .ZN(n4232) );
  INV_X1 U4678 ( .A(n3971), .ZN(n3972) );
  OAI21_X1 U4679 ( .B1(n3988), .B2(n3973), .A(n3972), .ZN(n4300) );
  AOI22_X1 U4680 ( .A1(n3974), .A2(n4476), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4477), .ZN(n3975) );
  OAI21_X1 U4681 ( .B1(n4300), .B2(n4195), .A(n3975), .ZN(n3976) );
  AOI21_X1 U4682 ( .B1(n4232), .B2(n4198), .A(n3976), .ZN(n3977) );
  OAI21_X1 U4683 ( .B1(n3978), .B2(n4202), .A(n3977), .ZN(U3264) );
  XNOR2_X1 U4684 ( .A(n3979), .B(n3980), .ZN(n4236) );
  INV_X1 U4685 ( .A(n4236), .ZN(n3995) );
  XNOR2_X1 U4686 ( .A(n3981), .B(n3980), .ZN(n3982) );
  NAND2_X1 U4687 ( .A1(n3982), .A2(n4184), .ZN(n3986) );
  AOI22_X1 U4688 ( .A1(n3984), .A2(n4187), .B1(n4216), .B2(n3983), .ZN(n3985)
         );
  OAI211_X1 U4689 ( .C1(n3987), .C2(n4191), .A(n3986), .B(n3985), .ZN(n4235)
         );
  INV_X1 U4690 ( .A(n3988), .ZN(n3989) );
  OAI21_X1 U4691 ( .B1(n2155), .B2(n3990), .A(n3989), .ZN(n4304) );
  AOI22_X1 U4692 ( .A1(n3991), .A2(n4476), .B1(REG2_REG_25__SCAN_IN), .B2(
        n4477), .ZN(n3992) );
  OAI21_X1 U4693 ( .B1(n4304), .B2(n4195), .A(n3992), .ZN(n3993) );
  AOI21_X1 U4694 ( .B1(n4235), .B2(n4198), .A(n3993), .ZN(n3994) );
  OAI21_X1 U4695 ( .B1(n3995), .B2(n4202), .A(n3994), .ZN(U3265) );
  XOR2_X1 U4696 ( .A(n3997), .B(n3996), .Z(n4240) );
  AOI21_X1 U4697 ( .B1(n4006), .B2(n4028), .A(n2155), .ZN(n4308) );
  INV_X1 U4698 ( .A(n3998), .ZN(n3999) );
  INV_X1 U4699 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4698) );
  OAI22_X1 U4700 ( .A1(n3999), .A2(n4196), .B1(n4198), .B2(n4698), .ZN(n4013)
         );
  INV_X1 U4701 ( .A(n4000), .ZN(n4001) );
  OR2_X1 U4702 ( .A1(n4002), .A2(n4001), .ZN(n4004) );
  XNOR2_X1 U4703 ( .A(n4004), .B(n4003), .ZN(n4011) );
  NAND2_X1 U4704 ( .A1(n4005), .A2(n4187), .ZN(n4008) );
  NAND2_X1 U4705 ( .A1(n4006), .A2(n4216), .ZN(n4007) );
  OAI211_X1 U4706 ( .C1(n4009), .C2(n4191), .A(n4008), .B(n4007), .ZN(n4010)
         );
  AOI21_X1 U4707 ( .B1(n4011), .B2(n4184), .A(n4010), .ZN(n4239) );
  NOR2_X1 U4708 ( .A1(n4239), .A2(n4477), .ZN(n4012) );
  AOI211_X1 U4709 ( .C1(n4308), .C2(n4479), .A(n4013), .B(n4012), .ZN(n4014)
         );
  OAI21_X1 U4710 ( .B1(n4240), .B2(n4202), .A(n4014), .ZN(U3266) );
  XOR2_X1 U4711 ( .A(n4019), .B(n4015), .Z(n4245) );
  INV_X1 U4712 ( .A(n4245), .ZN(n4036) );
  NAND2_X1 U4713 ( .A1(n2145), .A2(n4016), .ZN(n4059) );
  NAND2_X1 U4714 ( .A1(n4059), .A2(n4060), .ZN(n4058) );
  NAND2_X1 U4715 ( .A1(n4058), .A2(n4017), .ZN(n4041) );
  NAND2_X1 U4716 ( .A1(n4041), .A2(n4040), .ZN(n4043) );
  NAND2_X1 U4717 ( .A1(n4043), .A2(n4018), .ZN(n4020) );
  XNOR2_X1 U4718 ( .A(n4020), .B(n4019), .ZN(n4026) );
  OAI22_X1 U4719 ( .A1(n4021), .A2(n4191), .B1(n4127), .B2(n4029), .ZN(n4022)
         );
  AOI21_X1 U4720 ( .B1(n4187), .B2(n4023), .A(n4022), .ZN(n4024) );
  OAI21_X1 U4721 ( .B1(n4026), .B2(n4025), .A(n4024), .ZN(n4244) );
  INV_X1 U4722 ( .A(n4027), .ZN(n4030) );
  OAI21_X1 U4723 ( .B1(n4030), .B2(n4029), .A(n4028), .ZN(n4312) );
  INV_X1 U4724 ( .A(n4031), .ZN(n4032) );
  AOI22_X1 U4725 ( .A1(REG2_REG_23__SCAN_IN), .A2(n4477), .B1(n4032), .B2(
        n4476), .ZN(n4033) );
  OAI21_X1 U4726 ( .B1(n4312), .B2(n4195), .A(n4033), .ZN(n4034) );
  AOI21_X1 U4727 ( .B1(n4244), .B2(n4198), .A(n4034), .ZN(n4035) );
  OAI21_X1 U4728 ( .B1(n4036), .B2(n4202), .A(n4035), .ZN(U3267) );
  OAI21_X1 U4729 ( .B1(n4039), .B2(n4038), .A(n4037), .ZN(n4251) );
  OR2_X1 U4730 ( .A1(n4041), .A2(n4040), .ZN(n4042) );
  NAND2_X1 U4731 ( .A1(n4043), .A2(n4042), .ZN(n4050) );
  NAND2_X1 U4732 ( .A1(n4044), .A2(n4187), .ZN(n4047) );
  NAND2_X1 U4733 ( .A1(n4045), .A2(n4216), .ZN(n4046) );
  OAI211_X1 U4734 ( .C1(n4048), .C2(n4191), .A(n4047), .B(n4046), .ZN(n4049)
         );
  AOI21_X1 U4735 ( .B1(n4050), .B2(n4184), .A(n4049), .ZN(n4250) );
  AOI22_X1 U4736 ( .A1(n4477), .A2(REG2_REG_22__SCAN_IN), .B1(n4051), .B2(
        n4476), .ZN(n4054) );
  OR2_X1 U4737 ( .A1(n4067), .A2(n4052), .ZN(n4248) );
  NAND3_X1 U4738 ( .A1(n4027), .A2(n4248), .A3(n4479), .ZN(n4053) );
  OAI211_X1 U4739 ( .C1(n4250), .C2(n4477), .A(n4054), .B(n4053), .ZN(n4055)
         );
  INV_X1 U4740 ( .A(n4055), .ZN(n4056) );
  OAI21_X1 U4741 ( .B1(n4251), .B2(n4202), .A(n4056), .ZN(U3268) );
  XOR2_X1 U4742 ( .A(n4060), .B(n4057), .Z(n4253) );
  INV_X1 U4743 ( .A(n4253), .ZN(n4076) );
  OAI21_X1 U4744 ( .B1(n4060), .B2(n4059), .A(n4058), .ZN(n4061) );
  NAND2_X1 U4745 ( .A1(n4061), .A2(n4184), .ZN(n4065) );
  AOI22_X1 U4746 ( .A1(n4063), .A2(n4187), .B1(n4216), .B2(n4062), .ZN(n4064)
         );
  OAI211_X1 U4747 ( .C1(n4066), .C2(n4191), .A(n4065), .B(n4064), .ZN(n4252)
         );
  INV_X1 U4748 ( .A(n4090), .ZN(n4070) );
  INV_X1 U4749 ( .A(n4067), .ZN(n4068) );
  OAI21_X1 U4750 ( .B1(n4070), .B2(n4069), .A(n4068), .ZN(n4317) );
  INV_X1 U4751 ( .A(n4071), .ZN(n4072) );
  AOI22_X1 U4752 ( .A1(n4477), .A2(REG2_REG_21__SCAN_IN), .B1(n4072), .B2(
        n4476), .ZN(n4073) );
  OAI21_X1 U4753 ( .B1(n4317), .B2(n4195), .A(n4073), .ZN(n4074) );
  AOI21_X1 U4754 ( .B1(n4252), .B2(n4198), .A(n4074), .ZN(n4075) );
  OAI21_X1 U4755 ( .B1(n4076), .B2(n4202), .A(n4075), .ZN(U3269) );
  XNOR2_X1 U4756 ( .A(n4077), .B(n4082), .ZN(n4255) );
  INV_X1 U4757 ( .A(n4078), .ZN(n4079) );
  NAND2_X1 U4758 ( .A1(n4080), .A2(n4079), .ZN(n4081) );
  XOR2_X1 U4759 ( .A(n4082), .B(n4081), .Z(n4087) );
  AOI22_X1 U4760 ( .A1(n4084), .A2(n4187), .B1(n4216), .B2(n4083), .ZN(n4085)
         );
  OAI21_X1 U4761 ( .B1(n4129), .B2(n4191), .A(n4085), .ZN(n4086) );
  AOI21_X1 U4762 ( .B1(n4087), .B2(n4184), .A(n4086), .ZN(n4088) );
  OAI21_X1 U4763 ( .B1(n4255), .B2(n4089), .A(n4088), .ZN(n4256) );
  NAND2_X1 U4764 ( .A1(n4256), .A2(n4198), .ZN(n4098) );
  INV_X1 U4765 ( .A(n4115), .ZN(n4092) );
  OAI21_X1 U4766 ( .B1(n4092), .B2(n4091), .A(n4090), .ZN(n4321) );
  INV_X1 U4767 ( .A(n4321), .ZN(n4096) );
  INV_X1 U4768 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4094) );
  OAI22_X1 U4769 ( .A1(n4198), .A2(n4094), .B1(n4093), .B2(n4196), .ZN(n4095)
         );
  AOI21_X1 U4770 ( .B1(n4096), .B2(n4479), .A(n4095), .ZN(n4097) );
  OAI211_X1 U4771 ( .C1(n4255), .C2(n4099), .A(n4098), .B(n4097), .ZN(U3270)
         );
  XNOR2_X1 U4772 ( .A(n4100), .B(n4108), .ZN(n4261) );
  INV_X1 U4773 ( .A(n4261), .ZN(n4121) );
  INV_X1 U4774 ( .A(n4101), .ZN(n4102) );
  NOR2_X1 U4775 ( .A1(n4103), .A2(n4102), .ZN(n4126) );
  INV_X1 U4776 ( .A(n4104), .ZN(n4105) );
  AOI21_X1 U4777 ( .B1(n4126), .B2(n4106), .A(n4105), .ZN(n4107) );
  XOR2_X1 U4778 ( .A(n4108), .B(n4107), .Z(n4109) );
  NAND2_X1 U4779 ( .A1(n4109), .A2(n4184), .ZN(n4113) );
  AOI22_X1 U4780 ( .A1(n4111), .A2(n4187), .B1(n4216), .B2(n4110), .ZN(n4112)
         );
  OAI211_X1 U4781 ( .C1(n4114), .C2(n4191), .A(n4113), .B(n4112), .ZN(n4260)
         );
  OAI21_X1 U4782 ( .B1(n4135), .B2(n4116), .A(n4115), .ZN(n4325) );
  NOR2_X1 U4783 ( .A1(n4325), .A2(n4195), .ZN(n4119) );
  OAI22_X1 U4784 ( .A1(n4198), .A2(n4699), .B1(n4117), .B2(n4196), .ZN(n4118)
         );
  AOI211_X1 U4785 ( .C1(n4260), .C2(n4198), .A(n4119), .B(n4118), .ZN(n4120)
         );
  OAI21_X1 U4786 ( .B1(n4121), .B2(n4202), .A(n4120), .ZN(U3271) );
  OAI21_X1 U4787 ( .B1(n4123), .B2(n4125), .A(n4122), .ZN(n4124) );
  INV_X1 U4788 ( .A(n4124), .ZN(n4265) );
  XNOR2_X1 U4789 ( .A(n4126), .B(n4125), .ZN(n4134) );
  OAI22_X1 U4790 ( .A1(n4129), .A2(n4128), .B1(n4127), .B2(n3896), .ZN(n4132)
         );
  NOR2_X1 U4791 ( .A1(n4130), .A2(n4191), .ZN(n4131) );
  OR2_X1 U4792 ( .A1(n4132), .A2(n4131), .ZN(n4133) );
  AOI21_X1 U4793 ( .B1(n4134), .B2(n4184), .A(n4133), .ZN(n4264) );
  INV_X1 U4794 ( .A(n4264), .ZN(n4142) );
  INV_X1 U4795 ( .A(n4135), .ZN(n4136) );
  OAI211_X1 U4796 ( .C1(n4153), .C2(n3896), .A(n4136), .B(n4536), .ZN(n4263)
         );
  NOR2_X1 U4797 ( .A1(n4263), .A2(n4137), .ZN(n4141) );
  INV_X1 U4798 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4139) );
  OAI22_X1 U4799 ( .A1(n4198), .A2(n4139), .B1(n4138), .B2(n4196), .ZN(n4140)
         );
  AOI211_X1 U4800 ( .C1(n4142), .C2(n4198), .A(n4141), .B(n4140), .ZN(n4143)
         );
  OAI21_X1 U4801 ( .B1(n4265), .B2(n4202), .A(n4143), .ZN(U3272) );
  XOR2_X1 U4802 ( .A(n4146), .B(n4144), .Z(n4267) );
  INV_X1 U4803 ( .A(n4267), .ZN(n4161) );
  XOR2_X1 U4804 ( .A(n4146), .B(n4145), .Z(n4147) );
  NAND2_X1 U4805 ( .A1(n4147), .A2(n4184), .ZN(n4151) );
  AOI22_X1 U4806 ( .A1(n4149), .A2(n4187), .B1(n4216), .B2(n4148), .ZN(n4150)
         );
  OAI211_X1 U4807 ( .C1(n4152), .C2(n4191), .A(n4151), .B(n4150), .ZN(n4266)
         );
  INV_X1 U4808 ( .A(n4270), .ZN(n4156) );
  INV_X1 U4809 ( .A(n4153), .ZN(n4154) );
  OAI21_X1 U4810 ( .B1(n4156), .B2(n4155), .A(n4154), .ZN(n4329) );
  NOR2_X1 U4811 ( .A1(n4329), .A2(n4195), .ZN(n4159) );
  OAI22_X1 U4812 ( .A1(n4198), .A2(n2181), .B1(n4157), .B2(n4196), .ZN(n4158)
         );
  AOI211_X1 U4813 ( .C1(n4266), .C2(n4198), .A(n4159), .B(n4158), .ZN(n4160)
         );
  OAI21_X1 U4814 ( .B1(n4161), .B2(n4202), .A(n4160), .ZN(U3273) );
  OAI21_X1 U4815 ( .B1(n4163), .B2(n4164), .A(n4162), .ZN(n4273) );
  XNOR2_X1 U4816 ( .A(n4165), .B(n4164), .ZN(n4170) );
  AOI22_X1 U4817 ( .A1(n4166), .A2(n4187), .B1(n4216), .B2(n4172), .ZN(n4167)
         );
  OAI21_X1 U4818 ( .B1(n4168), .B2(n4191), .A(n4167), .ZN(n4169) );
  AOI21_X1 U4819 ( .B1(n4170), .B2(n4184), .A(n4169), .ZN(n4272) );
  INV_X1 U4820 ( .A(n4272), .ZN(n4176) );
  NAND2_X1 U4821 ( .A1(n4171), .A2(n4172), .ZN(n4269) );
  AND3_X1 U4822 ( .A1(n4270), .A2(n4479), .A3(n4269), .ZN(n4175) );
  OAI22_X1 U4823 ( .A1(n4198), .A2(n4442), .B1(n4173), .B2(n4196), .ZN(n4174)
         );
  AOI211_X1 U4824 ( .C1(n4176), .C2(n4198), .A(n4175), .B(n4174), .ZN(n4177)
         );
  OAI21_X1 U4825 ( .B1(n4273), .B2(n4202), .A(n4177), .ZN(U3274) );
  XNOR2_X1 U4826 ( .A(n4179), .B(n4178), .ZN(n4275) );
  INV_X1 U4827 ( .A(n4275), .ZN(n4203) );
  NAND2_X1 U4828 ( .A1(n4181), .A2(n4180), .ZN(n4183) );
  XNOR2_X1 U4829 ( .A(n4183), .B(n4182), .ZN(n4185) );
  NAND2_X1 U4830 ( .A1(n4185), .A2(n4184), .ZN(n4190) );
  AOI22_X1 U4831 ( .A1(n4188), .A2(n4187), .B1(n4216), .B2(n4186), .ZN(n4189)
         );
  OAI211_X1 U4832 ( .C1(n4192), .C2(n4191), .A(n4190), .B(n4189), .ZN(n4274)
         );
  OAI21_X1 U4833 ( .B1(n4194), .B2(n4193), .A(n4171), .ZN(n4334) );
  NOR2_X1 U4834 ( .A1(n4334), .A2(n4195), .ZN(n4200) );
  OAI22_X1 U4835 ( .A1(n4198), .A2(n3840), .B1(n4197), .B2(n4196), .ZN(n4199)
         );
  AOI211_X1 U4836 ( .C1(n4274), .C2(n4198), .A(n4200), .B(n4199), .ZN(n4201)
         );
  OAI21_X1 U4837 ( .B1(n4203), .B2(n4202), .A(n4201), .ZN(U3275) );
  NAND2_X1 U4838 ( .A1(n4211), .A2(n4204), .ZN(n4212) );
  XNOR2_X1 U4839 ( .A(n4212), .B(n4205), .ZN(n4358) );
  INV_X1 U4840 ( .A(n4358), .ZN(n4288) );
  INV_X1 U4841 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4209) );
  AND2_X1 U4842 ( .A1(n4207), .A2(n4206), .ZN(n4215) );
  AOI21_X1 U4843 ( .B1(n4208), .B2(n4216), .A(n4215), .ZN(n4360) );
  MUX2_X1 U4844 ( .A(n4209), .B(n4360), .S(n4544), .Z(n4210) );
  OAI21_X1 U4845 ( .B1(n4288), .B2(n4286), .A(n4210), .ZN(U3549) );
  INV_X1 U4846 ( .A(n4211), .ZN(n4214) );
  INV_X1 U4847 ( .A(n4212), .ZN(n4213) );
  INV_X1 U4848 ( .A(n4361), .ZN(n4290) );
  INV_X1 U4849 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4218) );
  AOI21_X1 U4850 ( .B1(n4217), .B2(n4216), .A(n4215), .ZN(n4363) );
  MUX2_X1 U4851 ( .A(n4218), .B(n4363), .S(n4544), .Z(n4219) );
  OAI21_X1 U4852 ( .B1(n4290), .B2(n4286), .A(n4219), .ZN(U3548) );
  NAND2_X1 U4853 ( .A1(n4220), .A2(n4525), .ZN(n4223) );
  MUX2_X1 U4854 ( .A(REG1_REG_29__SCAN_IN), .B(n4291), .S(n4544), .Z(U3547) );
  INV_X1 U4855 ( .A(REG1_REG_28__SCAN_IN), .ZN(n4686) );
  AOI21_X1 U4856 ( .B1(n4225), .B2(n4525), .A(n4224), .ZN(n4292) );
  MUX2_X1 U4857 ( .A(n4686), .B(n4292), .S(n4544), .Z(n4227) );
  NAND2_X1 U4858 ( .A1(n4293), .A2(n4242), .ZN(n4226) );
  NAND2_X1 U4859 ( .A1(n4227), .A2(n4226), .ZN(U3546) );
  NAND2_X1 U4860 ( .A1(n4228), .A2(n4525), .ZN(n4230) );
  OAI211_X1 U4861 ( .C1(n4503), .C2(n4231), .A(n4230), .B(n4229), .ZN(n4296)
         );
  MUX2_X1 U4862 ( .A(REG1_REG_27__SCAN_IN), .B(n4296), .S(n4544), .Z(U3545) );
  INV_X1 U4863 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4687) );
  AOI21_X1 U4864 ( .B1(n4233), .B2(n4525), .A(n4232), .ZN(n4297) );
  MUX2_X1 U4865 ( .A(n4687), .B(n4297), .S(n4547), .Z(n4234) );
  OAI21_X1 U4866 ( .B1(n4286), .B2(n4300), .A(n4234), .ZN(U3544) );
  INV_X1 U4867 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4237) );
  AOI21_X1 U4868 ( .B1(n4236), .B2(n4525), .A(n4235), .ZN(n4301) );
  MUX2_X1 U4869 ( .A(n4237), .B(n4301), .S(n4544), .Z(n4238) );
  OAI21_X1 U4870 ( .B1(n4286), .B2(n4304), .A(n4238), .ZN(U3543) );
  INV_X1 U4871 ( .A(n4525), .ZN(n4512) );
  OAI21_X1 U4872 ( .B1(n4240), .B2(n4512), .A(n4239), .ZN(n4305) );
  MUX2_X1 U4873 ( .A(REG1_REG_24__SCAN_IN), .B(n4305), .S(n4544), .Z(n4241) );
  AOI21_X1 U4874 ( .B1(n4242), .B2(n4308), .A(n4241), .ZN(n4243) );
  INV_X1 U4875 ( .A(n4243), .ZN(U3542) );
  INV_X1 U4876 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4246) );
  AOI21_X1 U4877 ( .B1(n4245), .B2(n4525), .A(n4244), .ZN(n4310) );
  MUX2_X1 U4878 ( .A(n4246), .B(n4310), .S(n4544), .Z(n4247) );
  OAI21_X1 U4879 ( .B1(n4286), .B2(n4312), .A(n4247), .ZN(U3541) );
  NAND3_X1 U4880 ( .A1(n4248), .A2(n4536), .A3(n4027), .ZN(n4249) );
  OAI211_X1 U4881 ( .C1(n4251), .C2(n4512), .A(n4250), .B(n4249), .ZN(n4313)
         );
  MUX2_X1 U4882 ( .A(REG1_REG_22__SCAN_IN), .B(n4313), .S(n4544), .Z(U3540) );
  INV_X1 U4883 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4684) );
  AOI21_X1 U4884 ( .B1(n4253), .B2(n4525), .A(n4252), .ZN(n4314) );
  MUX2_X1 U4885 ( .A(n4684), .B(n4314), .S(n4544), .Z(n4254) );
  OAI21_X1 U4886 ( .B1(n4286), .B2(n4317), .A(n4254), .ZN(U3539) );
  INV_X1 U4887 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4258) );
  INV_X1 U4888 ( .A(n4255), .ZN(n4257) );
  AOI21_X1 U4889 ( .B1(n4510), .B2(n4257), .A(n4256), .ZN(n4318) );
  MUX2_X1 U4890 ( .A(n4258), .B(n4318), .S(n4544), .Z(n4259) );
  OAI21_X1 U4891 ( .B1(n4286), .B2(n4321), .A(n4259), .ZN(U3538) );
  INV_X1 U4892 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4681) );
  AOI21_X1 U4893 ( .B1(n4261), .B2(n4525), .A(n4260), .ZN(n4322) );
  MUX2_X1 U4894 ( .A(n4681), .B(n4322), .S(n4547), .Z(n4262) );
  OAI21_X1 U4895 ( .B1(n4286), .B2(n4325), .A(n4262), .ZN(U3537) );
  OAI211_X1 U4896 ( .C1(n4265), .C2(n4512), .A(n4264), .B(n4263), .ZN(n4326)
         );
  MUX2_X1 U4897 ( .A(REG1_REG_18__SCAN_IN), .B(n4326), .S(n4544), .Z(U3536) );
  AOI21_X1 U4898 ( .B1(n4267), .B2(n4525), .A(n4266), .ZN(n4327) );
  MUX2_X1 U4899 ( .A(n4678), .B(n4327), .S(n4547), .Z(n4268) );
  OAI21_X1 U4900 ( .B1(n4286), .B2(n4329), .A(n4268), .ZN(U3535) );
  NAND3_X1 U4901 ( .A1(n4270), .A2(n4536), .A3(n4269), .ZN(n4271) );
  OAI211_X1 U4902 ( .C1(n4273), .C2(n4512), .A(n4272), .B(n4271), .ZN(n4330)
         );
  MUX2_X1 U4903 ( .A(REG1_REG_16__SCAN_IN), .B(n4330), .S(n4544), .Z(U3534) );
  AOI21_X1 U4904 ( .B1(n4275), .B2(n4525), .A(n4274), .ZN(n4331) );
  MUX2_X1 U4905 ( .A(n4276), .B(n4331), .S(n4547), .Z(n4277) );
  OAI21_X1 U4906 ( .B1(n4286), .B2(n4334), .A(n4277), .ZN(U3533) );
  AOI21_X1 U4907 ( .B1(n4510), .B2(n4279), .A(n4278), .ZN(n4335) );
  MUX2_X1 U4908 ( .A(n4414), .B(n4335), .S(n4547), .Z(n4280) );
  OAI21_X1 U4909 ( .B1(n4286), .B2(n4338), .A(n4280), .ZN(U3532) );
  INV_X1 U4910 ( .A(n4281), .ZN(n4283) );
  AOI21_X1 U4911 ( .B1(n4510), .B2(n4283), .A(n4282), .ZN(n4339) );
  MUX2_X1 U4912 ( .A(n4284), .B(n4339), .S(n4547), .Z(n4285) );
  OAI21_X1 U4913 ( .B1(n4286), .B2(n4343), .A(n4285), .ZN(U3531) );
  MUX2_X1 U4914 ( .A(n3633), .B(n4360), .S(n4518), .Z(n4287) );
  OAI21_X1 U4915 ( .B1(n4288), .B2(n4342), .A(n4287), .ZN(U3517) );
  MUX2_X1 U4916 ( .A(n2456), .B(n4363), .S(n4518), .Z(n4289) );
  OAI21_X1 U4917 ( .B1(n4290), .B2(n4342), .A(n4289), .ZN(U3516) );
  MUX2_X1 U4918 ( .A(REG0_REG_29__SCAN_IN), .B(n4291), .S(n4518), .Z(U3515) );
  MUX2_X1 U4919 ( .A(n4668), .B(n4292), .S(n4518), .Z(n4295) );
  NAND2_X1 U4920 ( .A1(n4293), .A2(n4307), .ZN(n4294) );
  NAND2_X1 U4921 ( .A1(n4295), .A2(n4294), .ZN(U3514) );
  MUX2_X1 U4922 ( .A(REG0_REG_27__SCAN_IN), .B(n4296), .S(n4518), .Z(U3513) );
  INV_X1 U4923 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4298) );
  MUX2_X1 U4924 ( .A(n4298), .B(n4297), .S(n4518), .Z(n4299) );
  OAI21_X1 U4925 ( .B1(n4300), .B2(n4342), .A(n4299), .ZN(U3512) );
  INV_X1 U4926 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4302) );
  MUX2_X1 U4927 ( .A(n4302), .B(n4301), .S(n4518), .Z(n4303) );
  OAI21_X1 U4928 ( .B1(n4304), .B2(n4342), .A(n4303), .ZN(U3511) );
  MUX2_X1 U4929 ( .A(REG0_REG_24__SCAN_IN), .B(n4305), .S(n4518), .Z(n4306) );
  AOI21_X1 U4930 ( .B1(n4308), .B2(n4307), .A(n4306), .ZN(n4309) );
  INV_X1 U4931 ( .A(n4309), .ZN(U3510) );
  INV_X1 U4932 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4655) );
  MUX2_X1 U4933 ( .A(n4655), .B(n4310), .S(n4518), .Z(n4311) );
  OAI21_X1 U4934 ( .B1(n4312), .B2(n4342), .A(n4311), .ZN(U3509) );
  MUX2_X1 U4935 ( .A(REG0_REG_22__SCAN_IN), .B(n4313), .S(n4518), .Z(U3508) );
  MUX2_X1 U4936 ( .A(n4315), .B(n4314), .S(n4518), .Z(n4316) );
  OAI21_X1 U4937 ( .B1(n4317), .B2(n4342), .A(n4316), .ZN(U3507) );
  MUX2_X1 U4938 ( .A(n4319), .B(n4318), .S(n4518), .Z(n4320) );
  OAI21_X1 U4939 ( .B1(n4321), .B2(n4342), .A(n4320), .ZN(U3506) );
  MUX2_X1 U4940 ( .A(n4323), .B(n4322), .S(n4518), .Z(n4324) );
  OAI21_X1 U4941 ( .B1(n4325), .B2(n4342), .A(n4324), .ZN(U3505) );
  MUX2_X1 U4942 ( .A(REG0_REG_18__SCAN_IN), .B(n4326), .S(n4518), .Z(U3503) );
  MUX2_X1 U4943 ( .A(n4652), .B(n4327), .S(n4518), .Z(n4328) );
  OAI21_X1 U4944 ( .B1(n4329), .B2(n4342), .A(n4328), .ZN(U3501) );
  MUX2_X1 U4945 ( .A(REG0_REG_16__SCAN_IN), .B(n4330), .S(n4518), .Z(U3499) );
  MUX2_X1 U4946 ( .A(n4332), .B(n4331), .S(n4518), .Z(n4333) );
  OAI21_X1 U4947 ( .B1(n4334), .B2(n4342), .A(n4333), .ZN(U3497) );
  MUX2_X1 U4948 ( .A(n4336), .B(n4335), .S(n4518), .Z(n4337) );
  OAI21_X1 U4949 ( .B1(n4338), .B2(n4342), .A(n4337), .ZN(U3495) );
  MUX2_X1 U4950 ( .A(n4340), .B(n4339), .S(n4518), .Z(n4341) );
  OAI21_X1 U4951 ( .B1(n4343), .B2(n4342), .A(n4341), .ZN(U3493) );
  MUX2_X1 U4952 ( .A(DATAI_29_), .B(n4344), .S(STATE_REG_SCAN_IN), .Z(U3323)
         );
  MUX2_X1 U4953 ( .A(DATAI_28_), .B(n4345), .S(STATE_REG_SCAN_IN), .Z(U3324)
         );
  MUX2_X1 U4954 ( .A(n4346), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U4955 ( .A(n4347), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U4956 ( .A(n4348), .B(DATAI_25_), .S(U3149), .Z(U3327) );
  MUX2_X1 U4957 ( .A(n4349), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U4958 ( .A(n4350), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U4959 ( .A(n4421), .B(DATAI_14_), .S(U3149), .Z(U3338) );
  MUX2_X1 U4960 ( .A(n4351), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  MUX2_X1 U4961 ( .A(DATAI_7_), .B(n4352), .S(STATE_REG_SCAN_IN), .Z(U3345) );
  MUX2_X1 U4962 ( .A(n4353), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U4963 ( .A(DATAI_4_), .B(n4354), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4964 ( .A(DATAI_3_), .B(n4355), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U4965 ( .A(n4356), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  MUX2_X1 U4966 ( .A(DATAI_0_), .B(n4357), .S(STATE_REG_SCAN_IN), .Z(U3352) );
  AOI22_X1 U4967 ( .A1(n4358), .A2(n4479), .B1(n4477), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n4359) );
  OAI21_X1 U4968 ( .B1(n4477), .B2(n4360), .A(n4359), .ZN(U3260) );
  AOI22_X1 U4969 ( .A1(n4361), .A2(n4479), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4477), .ZN(n4362) );
  OAI21_X1 U4970 ( .B1(n4477), .B2(n4363), .A(n4362), .ZN(U3261) );
  INV_X1 U4971 ( .A(n4364), .ZN(n4369) );
  AOI211_X1 U4972 ( .C1(n4367), .C2(n4366), .A(n4365), .B(n4460), .ZN(n4368)
         );
  AOI211_X1 U4973 ( .C1(n4464), .C2(ADDR_REG_8__SCAN_IN), .A(n4369), .B(n4368), 
        .ZN(n4372) );
  OAI211_X1 U4974 ( .C1(n4475), .C2(n4499), .A(n4372), .B(n4371), .ZN(U3248)
         );
  AOI211_X1 U4975 ( .C1(n4375), .C2(n4374), .A(n4373), .B(n4460), .ZN(n4376)
         );
  AOI211_X1 U4976 ( .C1(n4464), .C2(ADDR_REG_10__SCAN_IN), .A(n4377), .B(n4376), .ZN(n4381) );
  OAI211_X1 U4977 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4379), .A(n4472), .B(n4378), .ZN(n4380) );
  OAI211_X1 U4978 ( .C1(n4475), .C2(n4498), .A(n4381), .B(n4380), .ZN(U3250)
         );
  AOI211_X1 U4979 ( .C1(n4384), .C2(n4383), .A(n4382), .B(n4460), .ZN(n4386)
         );
  AOI211_X1 U4980 ( .C1(n4464), .C2(ADDR_REG_11__SCAN_IN), .A(n4386), .B(n4385), .ZN(n4391) );
  OAI211_X1 U4981 ( .C1(n4389), .C2(n4388), .A(n4472), .B(n4387), .ZN(n4390)
         );
  OAI211_X1 U4982 ( .C1(n4475), .C2(n4496), .A(n4391), .B(n4390), .ZN(U3251)
         );
  INV_X1 U4983 ( .A(n4392), .ZN(n4397) );
  AOI211_X1 U4984 ( .C1(n4395), .C2(n4394), .A(n4393), .B(n4460), .ZN(n4396)
         );
  AOI211_X1 U4985 ( .C1(n4464), .C2(ADDR_REG_12__SCAN_IN), .A(n4397), .B(n4396), .ZN(n4401) );
  OAI211_X1 U4986 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4399), .A(n4472), .B(n4398), .ZN(n4400) );
  OAI211_X1 U4987 ( .C1(n4475), .C2(n4495), .A(n4401), .B(n4400), .ZN(U3252)
         );
  AOI211_X1 U4988 ( .C1(n4404), .C2(n4403), .A(n4402), .B(n4460), .ZN(n4405)
         );
  AOI211_X1 U4989 ( .C1(n4464), .C2(ADDR_REG_13__SCAN_IN), .A(n4406), .B(n4405), .ZN(n4412) );
  AOI22_X1 U4990 ( .A1(REG2_REG_13__SCAN_IN), .A2(n4407), .B1(n4494), .B2(
        n3243), .ZN(n4410) );
  AOI21_X1 U4991 ( .B1(n4410), .B2(n4409), .A(n4416), .ZN(n4408) );
  OAI21_X1 U4992 ( .B1(n4410), .B2(n4409), .A(n4408), .ZN(n4411) );
  OAI211_X1 U4993 ( .C1(n4475), .C2(n4494), .A(n4412), .B(n4411), .ZN(U3253)
         );
  INV_X1 U4994 ( .A(ADDR_REG_14__SCAN_IN), .ZN(n4714) );
  AOI211_X1 U4995 ( .C1(n4415), .C2(n4414), .A(n4413), .B(n4460), .ZN(n4420)
         );
  AOI211_X1 U4996 ( .C1(n4418), .C2(n4696), .A(n4417), .B(n4416), .ZN(n4419)
         );
  AOI211_X1 U4997 ( .C1(n4422), .C2(n4421), .A(n4420), .B(n4419), .ZN(n4424)
         );
  OAI211_X1 U4998 ( .C1(n4436), .C2(n4714), .A(n4424), .B(n4423), .ZN(U3254)
         );
  AOI211_X1 U4999 ( .C1(n2149), .C2(n4426), .A(n4425), .B(n4460), .ZN(n4427)
         );
  AOI211_X1 U5000 ( .C1(n4464), .C2(ADDR_REG_15__SCAN_IN), .A(n4428), .B(n4427), .ZN(n4434) );
  AOI21_X1 U5001 ( .B1(n4431), .B2(n4430), .A(n4429), .ZN(n4432) );
  NAND2_X1 U5002 ( .A1(n4472), .A2(n4432), .ZN(n4433) );
  OAI211_X1 U5003 ( .C1(n4475), .C2(n4493), .A(n4434), .B(n4433), .ZN(U3255)
         );
  INV_X1 U5004 ( .A(ADDR_REG_16__SCAN_IN), .ZN(n4711) );
  OAI21_X1 U5005 ( .B1(n4436), .B2(n4711), .A(n4435), .ZN(n4437) );
  INV_X1 U5006 ( .A(n4437), .ZN(n4447) );
  OAI21_X1 U5007 ( .B1(n4440), .B2(n4439), .A(n4438), .ZN(n4445) );
  OAI21_X1 U5008 ( .B1(n4443), .B2(n4442), .A(n4441), .ZN(n4444) );
  AOI22_X1 U5009 ( .A1(n4457), .A2(n4445), .B1(n4472), .B2(n4444), .ZN(n4446)
         );
  OAI211_X1 U5010 ( .C1(n4491), .C2(n4475), .A(n4447), .B(n4446), .ZN(U3256)
         );
  AOI21_X1 U5011 ( .B1(n4464), .B2(ADDR_REG_17__SCAN_IN), .A(n4448), .ZN(n4459) );
  OAI21_X1 U5012 ( .B1(n4451), .B2(n4450), .A(n4449), .ZN(n4456) );
  OAI21_X1 U5013 ( .B1(n4454), .B2(n4453), .A(n4452), .ZN(n4455) );
  AOI22_X1 U5014 ( .A1(n4457), .A2(n4456), .B1(n4472), .B2(n4455), .ZN(n4458)
         );
  OAI211_X1 U5015 ( .C1(n4490), .C2(n4475), .A(n4459), .B(n4458), .ZN(U3257)
         );
  AOI21_X1 U5016 ( .B1(n4470), .B2(n4469), .A(n4468), .ZN(n4471) );
  NAND2_X1 U5017 ( .A1(n4472), .A2(n4471), .ZN(n4473) );
  OAI211_X1 U5018 ( .C1(n4475), .C2(n4489), .A(n4474), .B(n4473), .ZN(U3258)
         );
  AOI22_X1 U5019 ( .A1(REG2_REG_2__SCAN_IN), .A2(n4477), .B1(
        REG3_REG_2__SCAN_IN), .B2(n4476), .ZN(n4483) );
  AOI22_X1 U5020 ( .A1(n4481), .A2(n4480), .B1(n4479), .B2(n4478), .ZN(n4482)
         );
  OAI211_X1 U5021 ( .C1(n4477), .C2(n4484), .A(n4483), .B(n4482), .ZN(U3288)
         );
  INV_X1 U5022 ( .A(D_REG_31__SCAN_IN), .ZN(n4639) );
  NOR2_X1 U5023 ( .A1(n4486), .A2(n4639), .ZN(U3291) );
  AND2_X1 U5024 ( .A1(D_REG_30__SCAN_IN), .A2(n4485), .ZN(U3292) );
  INV_X1 U5025 ( .A(D_REG_29__SCAN_IN), .ZN(n4637) );
  NOR2_X1 U5026 ( .A1(n4486), .A2(n4637), .ZN(U3293) );
  INV_X1 U5027 ( .A(D_REG_28__SCAN_IN), .ZN(n4636) );
  NOR2_X1 U5028 ( .A1(n4486), .A2(n4636), .ZN(U3294) );
  AND2_X1 U5029 ( .A1(D_REG_27__SCAN_IN), .A2(n4485), .ZN(U3295) );
  INV_X1 U5030 ( .A(D_REG_26__SCAN_IN), .ZN(n4629) );
  NOR2_X1 U5031 ( .A1(n4486), .A2(n4629), .ZN(U3296) );
  AND2_X1 U5032 ( .A1(D_REG_25__SCAN_IN), .A2(n4485), .ZN(U3297) );
  INV_X1 U5033 ( .A(D_REG_24__SCAN_IN), .ZN(n4630) );
  NOR2_X1 U5034 ( .A1(n4486), .A2(n4630), .ZN(U3298) );
  INV_X1 U5035 ( .A(D_REG_23__SCAN_IN), .ZN(n4627) );
  NOR2_X1 U5036 ( .A1(n4486), .A2(n4627), .ZN(U3299) );
  AND2_X1 U5037 ( .A1(D_REG_22__SCAN_IN), .A2(n4485), .ZN(U3300) );
  AND2_X1 U5038 ( .A1(D_REG_21__SCAN_IN), .A2(n4485), .ZN(U3301) );
  INV_X1 U5039 ( .A(D_REG_20__SCAN_IN), .ZN(n4626) );
  NOR2_X1 U5040 ( .A1(n4486), .A2(n4626), .ZN(U3302) );
  AND2_X1 U5041 ( .A1(D_REG_19__SCAN_IN), .A2(n4485), .ZN(U3303) );
  INV_X1 U5042 ( .A(D_REG_18__SCAN_IN), .ZN(n4624) );
  NOR2_X1 U5043 ( .A1(n4486), .A2(n4624), .ZN(U3304) );
  AND2_X1 U5044 ( .A1(D_REG_17__SCAN_IN), .A2(n4485), .ZN(U3305) );
  INV_X1 U5045 ( .A(D_REG_16__SCAN_IN), .ZN(n4623) );
  NOR2_X1 U5046 ( .A1(n4486), .A2(n4623), .ZN(U3306) );
  AND2_X1 U5047 ( .A1(D_REG_15__SCAN_IN), .A2(n4485), .ZN(U3307) );
  INV_X1 U5048 ( .A(D_REG_14__SCAN_IN), .ZN(n4807) );
  NOR2_X1 U5049 ( .A1(n4486), .A2(n4807), .ZN(U3308) );
  INV_X1 U5050 ( .A(D_REG_13__SCAN_IN), .ZN(n4621) );
  NOR2_X1 U5051 ( .A1(n4486), .A2(n4621), .ZN(U3309) );
  AND2_X1 U5052 ( .A1(D_REG_12__SCAN_IN), .A2(n4485), .ZN(U3310) );
  INV_X1 U5053 ( .A(D_REG_11__SCAN_IN), .ZN(n4615) );
  NOR2_X1 U5054 ( .A1(n4486), .A2(n4615), .ZN(U3311) );
  INV_X1 U5055 ( .A(D_REG_10__SCAN_IN), .ZN(n4614) );
  NOR2_X1 U5056 ( .A1(n4486), .A2(n4614), .ZN(U3312) );
  INV_X1 U5057 ( .A(D_REG_9__SCAN_IN), .ZN(n4612) );
  NOR2_X1 U5058 ( .A1(n4486), .A2(n4612), .ZN(U3313) );
  AND2_X1 U5059 ( .A1(D_REG_8__SCAN_IN), .A2(n4485), .ZN(U3314) );
  INV_X1 U5060 ( .A(D_REG_7__SCAN_IN), .ZN(n4611) );
  NOR2_X1 U5061 ( .A1(n4486), .A2(n4611), .ZN(U3315) );
  INV_X1 U5062 ( .A(D_REG_6__SCAN_IN), .ZN(n4608) );
  NOR2_X1 U5063 ( .A1(n4486), .A2(n4608), .ZN(U3316) );
  INV_X1 U5064 ( .A(D_REG_5__SCAN_IN), .ZN(n4609) );
  NOR2_X1 U5065 ( .A1(n4486), .A2(n4609), .ZN(U3317) );
  AND2_X1 U5066 ( .A1(D_REG_4__SCAN_IN), .A2(n4485), .ZN(U3318) );
  AND2_X1 U5067 ( .A1(D_REG_3__SCAN_IN), .A2(n4485), .ZN(U3319) );
  INV_X1 U5068 ( .A(D_REG_2__SCAN_IN), .ZN(n4606) );
  NOR2_X1 U5069 ( .A1(n4486), .A2(n4606), .ZN(U3320) );
  INV_X1 U5070 ( .A(DATAI_23_), .ZN(n4488) );
  AOI21_X1 U5071 ( .B1(U3149), .B2(n4488), .A(n4487), .ZN(U3329) );
  INV_X1 U5072 ( .A(DATAI_18_), .ZN(n4566) );
  AOI22_X1 U5073 ( .A1(STATE_REG_SCAN_IN), .A2(n4489), .B1(n4566), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U5074 ( .A1(STATE_REG_SCAN_IN), .A2(n4490), .B1(n4565), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U5075 ( .A(DATAI_16_), .ZN(n4568) );
  AOI22_X1 U5076 ( .A1(STATE_REG_SCAN_IN), .A2(n4491), .B1(n4568), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5077 ( .A(DATAI_15_), .ZN(n4492) );
  AOI22_X1 U5078 ( .A1(STATE_REG_SCAN_IN), .A2(n4493), .B1(n4492), .B2(U3149), 
        .ZN(U3337) );
  AOI22_X1 U5079 ( .A1(STATE_REG_SCAN_IN), .A2(n4494), .B1(n3158), .B2(U3149), 
        .ZN(U3339) );
  AOI22_X1 U5080 ( .A1(STATE_REG_SCAN_IN), .A2(n4495), .B1(n4571), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5081 ( .A(DATAI_11_), .ZN(n4572) );
  AOI22_X1 U5082 ( .A1(STATE_REG_SCAN_IN), .A2(n4496), .B1(n4572), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5083 ( .A(DATAI_10_), .ZN(n4497) );
  AOI22_X1 U5084 ( .A1(STATE_REG_SCAN_IN), .A2(n4498), .B1(n4497), .B2(U3149), 
        .ZN(U3342) );
  AOI22_X1 U5085 ( .A1(STATE_REG_SCAN_IN), .A2(n4499), .B1(n2967), .B2(U3149), 
        .ZN(U3344) );
  AOI22_X1 U5086 ( .A1(n4518), .A2(n4500), .B1(n2353), .B2(n4790), .ZN(U3467)
         );
  AOI22_X1 U5087 ( .A1(n4518), .A2(n4501), .B1(n2335), .B2(n4790), .ZN(U3469)
         );
  OAI22_X1 U5088 ( .A1(n4504), .A2(n4540), .B1(n4503), .B2(n4502), .ZN(n4505)
         );
  NOR2_X1 U5089 ( .A1(n4506), .A2(n4505), .ZN(n4531) );
  AOI22_X1 U5090 ( .A1(n4518), .A2(n4531), .B1(n2566), .B2(n4790), .ZN(U3473)
         );
  INV_X1 U5091 ( .A(n4507), .ZN(n4509) );
  AOI211_X1 U5092 ( .C1(n4511), .C2(n4510), .A(n4509), .B(n4508), .ZN(n4533)
         );
  INV_X1 U5093 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4826) );
  AOI22_X1 U5094 ( .A1(n4518), .A2(n4533), .B1(n4826), .B2(n4790), .ZN(U3475)
         );
  NOR2_X1 U5095 ( .A1(n4513), .A2(n4512), .ZN(n4516) );
  INV_X1 U5096 ( .A(n4514), .ZN(n4515) );
  AOI211_X1 U5097 ( .C1(n4536), .C2(n4517), .A(n4516), .B(n4515), .ZN(n4535)
         );
  AOI22_X1 U5098 ( .A1(n4518), .A2(n4535), .B1(n2515), .B2(n4790), .ZN(U3477)
         );
  NAND3_X1 U5099 ( .A1(n4520), .A2(n4519), .A3(n4525), .ZN(n4522) );
  AND2_X1 U5100 ( .A1(n4522), .A2(n4521), .ZN(n4523) );
  AND2_X1 U5101 ( .A1(n4524), .A2(n4523), .ZN(n4543) );
  AOI22_X1 U5102 ( .A1(n4518), .A2(n4543), .B1(n2878), .B2(n4790), .ZN(U3481)
         );
  NAND2_X1 U5103 ( .A1(n4526), .A2(n4525), .ZN(n4529) );
  NAND2_X1 U5104 ( .A1(n4527), .A2(n4536), .ZN(n4528) );
  AOI22_X1 U5105 ( .A1(n4518), .A2(n4546), .B1(n2447), .B2(n4790), .ZN(U3485)
         );
  INV_X1 U5106 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4827) );
  AOI22_X1 U5107 ( .A1(n4544), .A2(n4531), .B1(n4827), .B2(n4545), .ZN(U3521)
         );
  INV_X1 U5108 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4532) );
  AOI22_X1 U5109 ( .A1(n4544), .A2(n4533), .B1(n4532), .B2(n4545), .ZN(U3522)
         );
  AOI22_X1 U5110 ( .A1(n4544), .A2(n4535), .B1(n4534), .B2(n4545), .ZN(U3523)
         );
  NAND2_X1 U5111 ( .A1(n4537), .A2(n4536), .ZN(n4538) );
  OAI211_X1 U5112 ( .C1(n4541), .C2(n4540), .A(n4539), .B(n4538), .ZN(n4791)
         );
  OAI22_X1 U5113 ( .A1(n4545), .A2(n4791), .B1(REG1_REG_6__SCAN_IN), .B2(n4544), .ZN(n4542) );
  INV_X1 U5114 ( .A(n4542), .ZN(U3524) );
  AOI22_X1 U5115 ( .A1(n4544), .A2(n4543), .B1(n4820), .B2(n4545), .ZN(U3525)
         );
  AOI22_X1 U5116 ( .A1(n4547), .A2(n4546), .B1(n2705), .B2(n4545), .ZN(U3527)
         );
  INV_X1 U5117 ( .A(DATAI_28_), .ZN(n4550) );
  AOI22_X1 U5118 ( .A1(n4550), .A2(keyinput85), .B1(keyinput96), .B2(n4549), 
        .ZN(n4548) );
  OAI221_X1 U5119 ( .B1(n4550), .B2(keyinput85), .C1(n4549), .C2(keyinput96), 
        .A(n4548), .ZN(n4563) );
  INV_X1 U5120 ( .A(DATAI_27_), .ZN(n4553) );
  INV_X1 U5121 ( .A(DATAI_26_), .ZN(n4552) );
  AOI22_X1 U5122 ( .A1(n4553), .A2(keyinput110), .B1(keyinput6), .B2(n4552), 
        .ZN(n4551) );
  OAI221_X1 U5123 ( .B1(n4553), .B2(keyinput110), .C1(n4552), .C2(keyinput6), 
        .A(n4551), .ZN(n4562) );
  INV_X1 U5124 ( .A(DATAI_24_), .ZN(n4556) );
  AOI22_X1 U5125 ( .A1(n4556), .A2(keyinput93), .B1(n4555), .B2(keyinput81), 
        .ZN(n4554) );
  OAI221_X1 U5126 ( .B1(n4556), .B2(keyinput93), .C1(n4555), .C2(keyinput81), 
        .A(n4554), .ZN(n4561) );
  INV_X1 U5127 ( .A(DATAI_19_), .ZN(n4559) );
  AOI22_X1 U5128 ( .A1(n4559), .A2(keyinput71), .B1(n4558), .B2(keyinput13), 
        .ZN(n4557) );
  OAI221_X1 U5129 ( .B1(n4559), .B2(keyinput71), .C1(n4558), .C2(keyinput13), 
        .A(n4557), .ZN(n4560) );
  NOR4_X1 U5130 ( .A1(n4563), .A2(n4562), .A3(n4561), .A4(n4560), .ZN(n4603)
         );
  AOI22_X1 U5131 ( .A1(n4566), .A2(keyinput66), .B1(n4565), .B2(keyinput80), 
        .ZN(n4564) );
  OAI221_X1 U5132 ( .B1(n4566), .B2(keyinput66), .C1(n4565), .C2(keyinput80), 
        .A(n4564), .ZN(n4579) );
  INV_X1 U5133 ( .A(DATAI_14_), .ZN(n4569) );
  AOI22_X1 U5134 ( .A1(n4569), .A2(keyinput62), .B1(n4568), .B2(keyinput60), 
        .ZN(n4567) );
  OAI221_X1 U5135 ( .B1(n4569), .B2(keyinput62), .C1(n4568), .C2(keyinput60), 
        .A(n4567), .ZN(n4578) );
  AOI22_X1 U5136 ( .A1(n4572), .A2(keyinput61), .B1(n4571), .B2(keyinput39), 
        .ZN(n4570) );
  OAI221_X1 U5137 ( .B1(n4572), .B2(keyinput61), .C1(n4571), .C2(keyinput39), 
        .A(n4570), .ZN(n4577) );
  INV_X1 U5138 ( .A(DATAI_6_), .ZN(n4575) );
  INV_X1 U5139 ( .A(DATAI_9_), .ZN(n4574) );
  AOI22_X1 U5140 ( .A1(n4575), .A2(keyinput38), .B1(n4574), .B2(keyinput123), 
        .ZN(n4573) );
  OAI221_X1 U5141 ( .B1(n4575), .B2(keyinput38), .C1(n4574), .C2(keyinput123), 
        .A(n4573), .ZN(n4576) );
  NOR4_X1 U5142 ( .A1(n4579), .A2(n4578), .A3(n4577), .A4(n4576), .ZN(n4602)
         );
  XOR2_X1 U5143 ( .A(n2718), .B(keyinput83), .Z(n4583) );
  XNOR2_X1 U5144 ( .A(REG3_REG_13__SCAN_IN), .B(keyinput90), .ZN(n4582) );
  XNOR2_X1 U5145 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput73), .ZN(n4581) );
  XNOR2_X1 U5146 ( .A(IR_REG_4__SCAN_IN), .B(keyinput28), .ZN(n4580) );
  NAND4_X1 U5147 ( .A1(n4583), .A2(n4582), .A3(n4581), .A4(n4580), .ZN(n4589)
         );
  XNOR2_X1 U5148 ( .A(STATE_REG_SCAN_IN), .B(keyinput117), .ZN(n4587) );
  XNOR2_X1 U5149 ( .A(DATAI_1_), .B(keyinput10), .ZN(n4586) );
  XNOR2_X1 U5150 ( .A(REG3_REG_21__SCAN_IN), .B(keyinput44), .ZN(n4585) );
  XNOR2_X1 U5151 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput48), .ZN(n4584) );
  NAND4_X1 U5152 ( .A1(n4587), .A2(n4586), .A3(n4585), .A4(n4584), .ZN(n4588)
         );
  NOR2_X1 U5153 ( .A1(n4589), .A2(n4588), .ZN(n4601) );
  XNOR2_X1 U5154 ( .A(IR_REG_8__SCAN_IN), .B(keyinput1), .ZN(n4593) );
  XNOR2_X1 U5155 ( .A(IR_REG_6__SCAN_IN), .B(keyinput12), .ZN(n4592) );
  XNOR2_X1 U5156 ( .A(IR_REG_10__SCAN_IN), .B(keyinput124), .ZN(n4591) );
  XNOR2_X1 U5157 ( .A(IR_REG_9__SCAN_IN), .B(keyinput36), .ZN(n4590) );
  NAND4_X1 U5158 ( .A1(n4593), .A2(n4592), .A3(n4591), .A4(n4590), .ZN(n4599)
         );
  XNOR2_X1 U5159 ( .A(IR_REG_16__SCAN_IN), .B(keyinput3), .ZN(n4597) );
  XNOR2_X1 U5160 ( .A(IR_REG_14__SCAN_IN), .B(keyinput114), .ZN(n4596) );
  XNOR2_X1 U5161 ( .A(IR_REG_28__SCAN_IN), .B(keyinput51), .ZN(n4595) );
  XNOR2_X1 U5162 ( .A(IR_REG_22__SCAN_IN), .B(keyinput104), .ZN(n4594) );
  NAND4_X1 U5163 ( .A1(n4597), .A2(n4596), .A3(n4595), .A4(n4594), .ZN(n4598)
         );
  NOR2_X1 U5164 ( .A1(n4599), .A2(n4598), .ZN(n4600) );
  NAND4_X1 U5165 ( .A1(n4603), .A2(n4602), .A3(n4601), .A4(n4600), .ZN(n4789)
         );
  AOI22_X1 U5166 ( .A1(n4606), .A2(keyinput50), .B1(n4605), .B2(keyinput25), 
        .ZN(n4604) );
  OAI221_X1 U5167 ( .B1(n4606), .B2(keyinput50), .C1(n4605), .C2(keyinput25), 
        .A(n4604), .ZN(n4619) );
  AOI22_X1 U5168 ( .A1(n4609), .A2(keyinput69), .B1(keyinput78), .B2(n4608), 
        .ZN(n4607) );
  OAI221_X1 U5169 ( .B1(n4609), .B2(keyinput69), .C1(n4608), .C2(keyinput78), 
        .A(n4607), .ZN(n4618) );
  AOI22_X1 U5170 ( .A1(n4612), .A2(keyinput94), .B1(n4611), .B2(keyinput103), 
        .ZN(n4610) );
  OAI221_X1 U5171 ( .B1(n4612), .B2(keyinput94), .C1(n4611), .C2(keyinput103), 
        .A(n4610), .ZN(n4617) );
  AOI22_X1 U5172 ( .A1(n4615), .A2(keyinput92), .B1(n4614), .B2(keyinput34), 
        .ZN(n4613) );
  OAI221_X1 U5173 ( .B1(n4615), .B2(keyinput92), .C1(n4614), .C2(keyinput34), 
        .A(n4613), .ZN(n4616) );
  NOR4_X1 U5174 ( .A1(n4619), .A2(n4618), .A3(n4617), .A4(n4616), .ZN(n4663)
         );
  AOI22_X1 U5175 ( .A1(n4807), .A2(keyinput32), .B1(n4621), .B2(keyinput29), 
        .ZN(n4620) );
  OAI221_X1 U5176 ( .B1(n4807), .B2(keyinput32), .C1(n4621), .C2(keyinput29), 
        .A(n4620), .ZN(n4634) );
  AOI22_X1 U5177 ( .A1(n4624), .A2(keyinput56), .B1(n4623), .B2(keyinput72), 
        .ZN(n4622) );
  OAI221_X1 U5178 ( .B1(n4624), .B2(keyinput56), .C1(n4623), .C2(keyinput72), 
        .A(n4622), .ZN(n4633) );
  AOI22_X1 U5179 ( .A1(n4627), .A2(keyinput8), .B1(n4626), .B2(keyinput0), 
        .ZN(n4625) );
  OAI221_X1 U5180 ( .B1(n4627), .B2(keyinput8), .C1(n4626), .C2(keyinput0), 
        .A(n4625), .ZN(n4632) );
  AOI22_X1 U5181 ( .A1(n4630), .A2(keyinput116), .B1(keyinput68), .B2(n4629), 
        .ZN(n4628) );
  OAI221_X1 U5182 ( .B1(n4630), .B2(keyinput116), .C1(n4629), .C2(keyinput68), 
        .A(n4628), .ZN(n4631) );
  NOR4_X1 U5183 ( .A1(n4634), .A2(n4633), .A3(n4632), .A4(n4631), .ZN(n4662)
         );
  AOI22_X1 U5184 ( .A1(n4637), .A2(keyinput20), .B1(n4636), .B2(keyinput54), 
        .ZN(n4635) );
  OAI221_X1 U5185 ( .B1(n4637), .B2(keyinput20), .C1(n4636), .C2(keyinput54), 
        .A(n4635), .ZN(n4645) );
  AOI22_X1 U5186 ( .A1(n2335), .A2(keyinput75), .B1(n4639), .B2(keyinput115), 
        .ZN(n4638) );
  OAI221_X1 U5187 ( .B1(n2335), .B2(keyinput75), .C1(n4639), .C2(keyinput115), 
        .A(n4638), .ZN(n4644) );
  AOI22_X1 U5188 ( .A1(n2377), .A2(keyinput14), .B1(keyinput86), .B2(n2566), 
        .ZN(n4640) );
  OAI221_X1 U5189 ( .B1(n2377), .B2(keyinput14), .C1(n2566), .C2(keyinput86), 
        .A(n4640), .ZN(n4643) );
  AOI22_X1 U5190 ( .A1(n2878), .A2(keyinput106), .B1(keyinput17), .B2(n4826), 
        .ZN(n4641) );
  OAI221_X1 U5191 ( .B1(n2878), .B2(keyinput106), .C1(n4826), .C2(keyinput17), 
        .A(n4641), .ZN(n4642) );
  NOR4_X1 U5192 ( .A1(n4645), .A2(n4644), .A3(n4643), .A4(n4642), .ZN(n4661)
         );
  AOI22_X1 U5193 ( .A1(n2901), .A2(keyinput87), .B1(n2447), .B2(keyinput126), 
        .ZN(n4646) );
  OAI221_X1 U5194 ( .B1(n2901), .B2(keyinput87), .C1(n2447), .C2(keyinput126), 
        .A(n4646), .ZN(n4659) );
  AOI22_X1 U5195 ( .A1(n4649), .A2(keyinput18), .B1(n4648), .B2(keyinput100), 
        .ZN(n4647) );
  OAI221_X1 U5196 ( .B1(n4649), .B2(keyinput18), .C1(n4648), .C2(keyinput100), 
        .A(n4647), .ZN(n4658) );
  AOI22_X1 U5197 ( .A1(n4652), .A2(keyinput99), .B1(n4651), .B2(keyinput46), 
        .ZN(n4650) );
  OAI221_X1 U5198 ( .B1(n4652), .B2(keyinput99), .C1(n4651), .C2(keyinput46), 
        .A(n4650), .ZN(n4657) );
  AOI22_X1 U5199 ( .A1(n4655), .A2(keyinput125), .B1(keyinput24), .B2(n4654), 
        .ZN(n4653) );
  OAI221_X1 U5200 ( .B1(n4655), .B2(keyinput125), .C1(n4654), .C2(keyinput24), 
        .A(n4653), .ZN(n4656) );
  NOR4_X1 U5201 ( .A1(n4659), .A2(n4658), .A3(n4657), .A4(n4656), .ZN(n4660)
         );
  NAND4_X1 U5202 ( .A1(n4663), .A2(n4662), .A3(n4661), .A4(n4660), .ZN(n4788)
         );
  AOI22_X1 U5203 ( .A1(n4827), .A2(keyinput101), .B1(n4820), .B2(keyinput120), 
        .ZN(n4664) );
  OAI221_X1 U5204 ( .B1(n4827), .B2(keyinput101), .C1(n4820), .C2(keyinput120), 
        .A(n4664), .ZN(n4675) );
  AOI22_X1 U5205 ( .A1(n4666), .A2(keyinput59), .B1(keyinput76), .B2(n2456), 
        .ZN(n4665) );
  OAI221_X1 U5206 ( .B1(n4666), .B2(keyinput59), .C1(n2456), .C2(keyinput76), 
        .A(n4665), .ZN(n4674) );
  AOI22_X1 U5207 ( .A1(n4669), .A2(keyinput47), .B1(n4668), .B2(keyinput15), 
        .ZN(n4667) );
  OAI221_X1 U5208 ( .B1(n4669), .B2(keyinput47), .C1(n4668), .C2(keyinput15), 
        .A(n4667), .ZN(n4673) );
  XNOR2_X1 U5209 ( .A(REG1_REG_2__SCAN_IN), .B(keyinput23), .ZN(n4671) );
  XNOR2_X1 U5210 ( .A(REG1_REG_0__SCAN_IN), .B(keyinput77), .ZN(n4670) );
  NAND2_X1 U5211 ( .A1(n4671), .A2(n4670), .ZN(n4672) );
  NOR4_X1 U5212 ( .A1(n4675), .A2(n4674), .A3(n4673), .A4(n4672), .ZN(n4722)
         );
  AOI22_X1 U5213 ( .A1(n4678), .A2(keyinput40), .B1(keyinput74), .B2(n4677), 
        .ZN(n4676) );
  OAI221_X1 U5214 ( .B1(n4678), .B2(keyinput40), .C1(n4677), .C2(keyinput74), 
        .A(n4676), .ZN(n4691) );
  AOI22_X1 U5215 ( .A1(n4681), .A2(keyinput122), .B1(keyinput95), .B2(n4680), 
        .ZN(n4679) );
  OAI221_X1 U5216 ( .B1(n4681), .B2(keyinput122), .C1(n4680), .C2(keyinput95), 
        .A(n4679), .ZN(n4690) );
  INV_X1 U5217 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4683) );
  AOI22_X1 U5218 ( .A1(n4684), .A2(keyinput65), .B1(n4683), .B2(keyinput30), 
        .ZN(n4682) );
  OAI221_X1 U5219 ( .B1(n4684), .B2(keyinput65), .C1(n4683), .C2(keyinput30), 
        .A(n4682), .ZN(n4689) );
  AOI22_X1 U5220 ( .A1(n4687), .A2(keyinput89), .B1(n4686), .B2(keyinput42), 
        .ZN(n4685) );
  OAI221_X1 U5221 ( .B1(n4687), .B2(keyinput89), .C1(n4686), .C2(keyinput42), 
        .A(n4685), .ZN(n4688) );
  NOR4_X1 U5222 ( .A1(n4691), .A2(n4690), .A3(n4689), .A4(n4688), .ZN(n4721)
         );
  AOI22_X1 U5223 ( .A1(n2480), .A2(keyinput112), .B1(n4693), .B2(keyinput11), 
        .ZN(n4692) );
  OAI221_X1 U5224 ( .B1(n2480), .B2(keyinput112), .C1(n4693), .C2(keyinput11), 
        .A(n4692), .ZN(n4703) );
  AOI22_X1 U5225 ( .A1(n2190), .A2(keyinput107), .B1(n4821), .B2(keyinput127), 
        .ZN(n4694) );
  OAI221_X1 U5226 ( .B1(n2190), .B2(keyinput107), .C1(n4821), .C2(keyinput127), 
        .A(n4694), .ZN(n4702) );
  AOI22_X1 U5227 ( .A1(n4139), .A2(keyinput119), .B1(n4696), .B2(keyinput45), 
        .ZN(n4695) );
  OAI221_X1 U5228 ( .B1(n4139), .B2(keyinput119), .C1(n4696), .C2(keyinput45), 
        .A(n4695), .ZN(n4701) );
  AOI22_X1 U5229 ( .A1(n4699), .A2(keyinput82), .B1(keyinput97), .B2(n4698), 
        .ZN(n4697) );
  OAI221_X1 U5230 ( .B1(n4699), .B2(keyinput82), .C1(n4698), .C2(keyinput97), 
        .A(n4697), .ZN(n4700) );
  NOR4_X1 U5231 ( .A1(n4703), .A2(n4702), .A3(n4701), .A4(n4700), .ZN(n4720)
         );
  INV_X1 U5232 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4705) );
  AOI22_X1 U5233 ( .A1(n4705), .A2(keyinput43), .B1(n3415), .B2(keyinput63), 
        .ZN(n4704) );
  OAI221_X1 U5234 ( .B1(n4705), .B2(keyinput43), .C1(n3415), .C2(keyinput63), 
        .A(n4704), .ZN(n4718) );
  INV_X1 U5235 ( .A(REG2_REG_28__SCAN_IN), .ZN(n4708) );
  INV_X1 U5236 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4707) );
  AOI22_X1 U5237 ( .A1(n4708), .A2(keyinput21), .B1(keyinput109), .B2(n4707), 
        .ZN(n4706) );
  OAI221_X1 U5238 ( .B1(n4708), .B2(keyinput21), .C1(n4707), .C2(keyinput109), 
        .A(n4706), .ZN(n4717) );
  INV_X1 U5239 ( .A(ADDR_REG_17__SCAN_IN), .ZN(n4710) );
  AOI22_X1 U5240 ( .A1(n4711), .A2(keyinput111), .B1(n4710), .B2(keyinput53), 
        .ZN(n4709) );
  OAI221_X1 U5241 ( .B1(n4711), .B2(keyinput111), .C1(n4710), .C2(keyinput53), 
        .A(n4709), .ZN(n4716) );
  INV_X1 U5242 ( .A(ADDR_REG_13__SCAN_IN), .ZN(n4713) );
  AOI22_X1 U5243 ( .A1(n4714), .A2(keyinput67), .B1(n4713), .B2(keyinput5), 
        .ZN(n4712) );
  OAI221_X1 U5244 ( .B1(n4714), .B2(keyinput67), .C1(n4713), .C2(keyinput5), 
        .A(n4712), .ZN(n4715) );
  NOR4_X1 U5245 ( .A1(n4718), .A2(n4717), .A3(n4716), .A4(n4715), .ZN(n4719)
         );
  NAND4_X1 U5246 ( .A1(n4722), .A2(n4721), .A3(n4720), .A4(n4719), .ZN(n4787)
         );
  INV_X1 U5247 ( .A(ADDR_REG_10__SCAN_IN), .ZN(n4725) );
  INV_X1 U5248 ( .A(ADDR_REG_12__SCAN_IN), .ZN(n4724) );
  AOI22_X1 U5249 ( .A1(n4725), .A2(keyinput108), .B1(keyinput102), .B2(n4724), 
        .ZN(n4723) );
  OAI221_X1 U5250 ( .B1(n4725), .B2(keyinput108), .C1(n4724), .C2(keyinput102), 
        .A(n4723), .ZN(n4738) );
  INV_X1 U5251 ( .A(ADDR_REG_8__SCAN_IN), .ZN(n4728) );
  INV_X1 U5252 ( .A(ADDR_REG_9__SCAN_IN), .ZN(n4727) );
  AOI22_X1 U5253 ( .A1(n4728), .A2(keyinput118), .B1(keyinput4), .B2(n4727), 
        .ZN(n4726) );
  OAI221_X1 U5254 ( .B1(n4728), .B2(keyinput118), .C1(n4727), .C2(keyinput4), 
        .A(n4726), .ZN(n4737) );
  AOI22_X1 U5255 ( .A1(n4731), .A2(keyinput105), .B1(n4730), .B2(keyinput98), 
        .ZN(n4729) );
  OAI221_X1 U5256 ( .B1(n4731), .B2(keyinput105), .C1(n4730), .C2(keyinput98), 
        .A(n4729), .ZN(n4736) );
  INV_X1 U5257 ( .A(ADDR_REG_4__SCAN_IN), .ZN(n4734) );
  INV_X1 U5258 ( .A(ADDR_REG_2__SCAN_IN), .ZN(n4733) );
  AOI22_X1 U5259 ( .A1(n4734), .A2(keyinput91), .B1(n4733), .B2(keyinput88), 
        .ZN(n4732) );
  OAI221_X1 U5260 ( .B1(n4734), .B2(keyinput91), .C1(n4733), .C2(keyinput88), 
        .A(n4732), .ZN(n4735) );
  NOR4_X1 U5261 ( .A1(n4738), .A2(n4737), .A3(n4736), .A4(n4735), .ZN(n4785)
         );
  INV_X1 U5262 ( .A(ADDR_REG_0__SCAN_IN), .ZN(n4741) );
  AOI22_X1 U5263 ( .A1(n4741), .A2(keyinput121), .B1(n4740), .B2(keyinput55), 
        .ZN(n4739) );
  OAI221_X1 U5264 ( .B1(n4741), .B2(keyinput121), .C1(n4740), .C2(keyinput55), 
        .A(n4739), .ZN(n4753) );
  AOI22_X1 U5265 ( .A1(n4744), .A2(keyinput57), .B1(keyinput35), .B2(n4743), 
        .ZN(n4742) );
  OAI221_X1 U5266 ( .B1(n4744), .B2(keyinput57), .C1(n4743), .C2(keyinput35), 
        .A(n4742), .ZN(n4752) );
  AOI22_X1 U5267 ( .A1(n4746), .A2(keyinput49), .B1(keyinput19), .B2(n4836), 
        .ZN(n4745) );
  OAI221_X1 U5268 ( .B1(n4746), .B2(keyinput49), .C1(n4836), .C2(keyinput19), 
        .A(n4745), .ZN(n4751) );
  AOI22_X1 U5269 ( .A1(n4749), .A2(keyinput7), .B1(n4748), .B2(keyinput70), 
        .ZN(n4747) );
  OAI221_X1 U5270 ( .B1(n4749), .B2(keyinput7), .C1(n4748), .C2(keyinput70), 
        .A(n4747), .ZN(n4750) );
  NOR4_X1 U5271 ( .A1(n4753), .A2(n4752), .A3(n4751), .A4(n4750), .ZN(n4784)
         );
  AOI22_X1 U5272 ( .A1(n4756), .A2(keyinput33), .B1(n4755), .B2(keyinput64), 
        .ZN(n4754) );
  OAI221_X1 U5273 ( .B1(n4756), .B2(keyinput33), .C1(n4755), .C2(keyinput64), 
        .A(n4754), .ZN(n4768) );
  AOI22_X1 U5274 ( .A1(n4759), .A2(keyinput52), .B1(n4758), .B2(keyinput26), 
        .ZN(n4757) );
  OAI221_X1 U5275 ( .B1(n4759), .B2(keyinput52), .C1(n4758), .C2(keyinput26), 
        .A(n4757), .ZN(n4767) );
  AOI22_X1 U5276 ( .A1(n4762), .A2(keyinput16), .B1(keyinput84), .B2(n4761), 
        .ZN(n4760) );
  OAI221_X1 U5277 ( .B1(n4762), .B2(keyinput16), .C1(n4761), .C2(keyinput84), 
        .A(n4760), .ZN(n4766) );
  INV_X1 U5278 ( .A(B_REG_SCAN_IN), .ZN(n4764) );
  AOI22_X1 U5279 ( .A1(n4764), .A2(keyinput37), .B1(keyinput41), .B2(n4837), 
        .ZN(n4763) );
  OAI221_X1 U5280 ( .B1(n4764), .B2(keyinput37), .C1(n4837), .C2(keyinput41), 
        .A(n4763), .ZN(n4765) );
  NOR4_X1 U5281 ( .A1(n4768), .A2(n4767), .A3(n4766), .A4(n4765), .ZN(n4783)
         );
  AOI22_X1 U5282 ( .A1(n4771), .A2(keyinput2), .B1(keyinput31), .B2(n4770), 
        .ZN(n4769) );
  OAI221_X1 U5283 ( .B1(n4771), .B2(keyinput2), .C1(n4770), .C2(keyinput31), 
        .A(n4769), .ZN(n4781) );
  AOI22_X1 U5284 ( .A1(n4773), .A2(keyinput9), .B1(keyinput113), .B2(n4828), 
        .ZN(n4772) );
  OAI221_X1 U5285 ( .B1(n4773), .B2(keyinput9), .C1(n4828), .C2(keyinput113), 
        .A(n4772), .ZN(n4780) );
  AOI22_X1 U5286 ( .A1(n4775), .A2(keyinput79), .B1(keyinput22), .B2(n2376), 
        .ZN(n4774) );
  OAI221_X1 U5287 ( .B1(n4775), .B2(keyinput79), .C1(n2376), .C2(keyinput22), 
        .A(n4774), .ZN(n4779) );
  AOI22_X1 U5288 ( .A1(n3511), .A2(keyinput27), .B1(n4777), .B2(keyinput58), 
        .ZN(n4776) );
  OAI221_X1 U5289 ( .B1(n3511), .B2(keyinput27), .C1(n4777), .C2(keyinput58), 
        .A(n4776), .ZN(n4778) );
  NOR4_X1 U5290 ( .A1(n4781), .A2(n4780), .A3(n4779), .A4(n4778), .ZN(n4782)
         );
  NAND4_X1 U5291 ( .A1(n4785), .A2(n4784), .A3(n4783), .A4(n4782), .ZN(n4786)
         );
  NOR4_X1 U5292 ( .A1(n4789), .A2(n4788), .A3(n4787), .A4(n4786), .ZN(n4793)
         );
  AOI22_X1 U5293 ( .A1(n4518), .A2(n4791), .B1(REG0_REG_6__SCAN_IN), .B2(n4790), .ZN(n4792) );
  XNOR2_X1 U5294 ( .A(n4793), .B(n4792), .ZN(n4855) );
  NAND4_X1 U5295 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n4795) );
  NAND4_X1 U5296 ( .A1(D_REG_13__SCAN_IN), .A2(D_REG_16__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n4794) );
  NOR2_X1 U5297 ( .A1(n4795), .A2(n4794), .ZN(n4803) );
  NAND4_X1 U5298 ( .A1(n4798), .A2(n4797), .A3(IR_REG_22__SCAN_IN), .A4(n4796), 
        .ZN(n4801) );
  NAND4_X1 U5299 ( .A1(n4799), .A2(IR_REG_6__SCAN_IN), .A3(IR_REG_8__SCAN_IN), 
        .A4(IR_REG_16__SCAN_IN), .ZN(n4800) );
  NOR2_X1 U5300 ( .A1(n4801), .A2(n4800), .ZN(n4802) );
  AND2_X1 U5301 ( .A1(n4803), .A2(n4802), .ZN(n4811) );
  NAND4_X1 U5302 ( .A1(n4804), .A2(STATE_REG_SCAN_IN), .A3(D_REG_29__SCAN_IN), 
        .A4(D_REG_28__SCAN_IN), .ZN(n4806) );
  NAND4_X1 U5303 ( .A1(B_REG_SCAN_IN), .A2(D_REG_1__SCAN_IN), .A3(
        D_REG_6__SCAN_IN), .A4(D_REG_7__SCAN_IN), .ZN(n4805) );
  NOR2_X1 U5304 ( .A1(n4806), .A2(n4805), .ZN(n4809) );
  AND4_X1 U5305 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(n4807), .ZN(n4808) );
  AND4_X1 U5306 ( .A1(n4811), .A2(n4810), .A3(n4809), .A4(n4808), .ZN(n4853)
         );
  NAND4_X1 U5307 ( .A1(DATAI_17_), .A2(ADDR_REG_12__SCAN_IN), .A3(
        ADDR_REG_9__SCAN_IN), .A4(ADDR_REG_4__SCAN_IN), .ZN(n4815) );
  NAND4_X1 U5308 ( .A1(REG0_REG_12__SCAN_IN), .A2(REG0_REG_8__SCAN_IN), .A3(
        ADDR_REG_17__SCAN_IN), .A4(ADDR_REG_10__SCAN_IN), .ZN(n4814) );
  NAND4_X1 U5309 ( .A1(REG2_REG_28__SCAN_IN), .A2(REG2_REG_27__SCAN_IN), .A3(
        REG2_REG_26__SCAN_IN), .A4(REG1_REG_18__SCAN_IN), .ZN(n4813) );
  NAND4_X1 U5310 ( .A1(DATAI_27_), .A2(DATAI_26_), .A3(DATAI_21_), .A4(
        DATAI_24_), .ZN(n4812) );
  NOR4_X1 U5311 ( .A1(n4815), .A2(n4814), .A3(n4813), .A4(n4812), .ZN(n4852)
         );
  NAND4_X1 U5312 ( .A1(REG0_REG_29__SCAN_IN), .A2(DATAO_REG_17__SCAN_IN), .A3(
        ADDR_REG_6__SCAN_IN), .A4(DATAO_REG_12__SCAN_IN), .ZN(n4819) );
  NAND4_X1 U5313 ( .A1(DATAI_31_), .A2(ADDR_REG_14__SCAN_IN), .A3(
        DATAO_REG_25__SCAN_IN), .A4(ADDR_REG_2__SCAN_IN), .ZN(n4818) );
  NAND4_X1 U5314 ( .A1(REG1_REG_21__SCAN_IN), .A2(REG0_REG_17__SCAN_IN), .A3(
        REG0_REG_9__SCAN_IN), .A4(REG2_REG_24__SCAN_IN), .ZN(n4817) );
  NAND4_X1 U5315 ( .A1(REG1_REG_26__SCAN_IN), .A2(REG0_REG_23__SCAN_IN), .A3(
        REG0_REG_24__SCAN_IN), .A4(DATAO_REG_10__SCAN_IN), .ZN(n4816) );
  NOR4_X1 U5316 ( .A1(n4819), .A2(n4818), .A3(n4817), .A4(n4816), .ZN(n4851)
         );
  NOR4_X1 U5317 ( .A1(REG3_REG_21__SCAN_IN), .A2(ADDR_REG_13__SCAN_IN), .A3(
        ADDR_REG_5__SCAN_IN), .A4(DATAO_REG_3__SCAN_IN), .ZN(n4825) );
  NOR4_X1 U5318 ( .A1(DATAI_20_), .A2(DATAI_9_), .A3(n4821), .A4(n4820), .ZN(
        n4824) );
  NOR4_X1 U5319 ( .A1(DATAI_16_), .A2(DATAO_REG_24__SCAN_IN), .A3(
        DATAO_REG_20__SCAN_IN), .A4(DATAO_REG_15__SCAN_IN), .ZN(n4823) );
  NOR4_X1 U5320 ( .A1(DATAO_REG_4__SCAN_IN), .A2(DATAO_REG_9__SCAN_IN), .A3(
        DATAO_REG_11__SCAN_IN), .A4(DATAO_REG_1__SCAN_IN), .ZN(n4822) );
  NAND4_X1 U5321 ( .A1(n4825), .A2(n4824), .A3(n4823), .A4(n4822), .ZN(n4849)
         );
  NOR4_X1 U5322 ( .A1(REG0_REG_3__SCAN_IN), .A2(REG2_REG_6__SCAN_IN), .A3(
        n2718), .A4(n2878), .ZN(n4835) );
  NOR4_X1 U5323 ( .A1(n4828), .A2(n4827), .A3(n4826), .A4(DATAI_6_), .ZN(n4834) );
  NOR4_X1 U5324 ( .A1(REG3_REG_2__SCAN_IN), .A2(n2480), .A3(n2377), .A4(n2335), 
        .ZN(n4830) );
  INV_X1 U5325 ( .A(DATAI_1_), .ZN(n4829) );
  NAND3_X1 U5326 ( .A1(n4830), .A2(REG1_REG_2__SCAN_IN), .A3(n4829), .ZN(n4832) );
  NOR3_X1 U5327 ( .A1(n4832), .A2(REG2_REG_5__SCAN_IN), .A3(n4831), .ZN(n4833)
         );
  NAND3_X1 U5328 ( .A1(n4835), .A2(n4834), .A3(n4833), .ZN(n4848) );
  NOR4_X1 U5329 ( .A1(DATAI_28_), .A2(DATAI_19_), .A3(DATAI_18_), .A4(n4836), 
        .ZN(n4841) );
  NOR4_X1 U5330 ( .A1(REG3_REG_13__SCAN_IN), .A2(REG3_REG_11__SCAN_IN), .A3(
        ADDR_REG_8__SCAN_IN), .A4(ADDR_REG_0__SCAN_IN), .ZN(n4840) );
  NOR4_X1 U5331 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG2_REG_25__SCAN_IN), .A3(
        REG1_REG_19__SCAN_IN), .A4(n4837), .ZN(n4839) );
  NOR4_X1 U5332 ( .A1(REG3_REG_27__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .A3(
        REG2_REG_19__SCAN_IN), .A4(REG2_REG_18__SCAN_IN), .ZN(n4838) );
  NAND4_X1 U5333 ( .A1(n4841), .A2(n4840), .A3(n4839), .A4(n4838), .ZN(n4847)
         );
  NOR4_X1 U5334 ( .A1(REG3_REG_18__SCAN_IN), .A2(REG0_REG_22__SCAN_IN), .A3(
        REG1_REG_22__SCAN_IN), .A4(REG0_REG_16__SCAN_IN), .ZN(n4845) );
  NOR4_X1 U5335 ( .A1(REG0_REG_28__SCAN_IN), .A2(REG1_REG_28__SCAN_IN), .A3(
        REG0_REG_27__SCAN_IN), .A4(REG0_REG_30__SCAN_IN), .ZN(n4844) );
  NOR4_X1 U5336 ( .A1(REG1_REG_17__SCAN_IN), .A2(REG2_REG_14__SCAN_IN), .A3(
        REG1_REG_11__SCAN_IN), .A4(ADDR_REG_16__SCAN_IN), .ZN(n4843) );
  NOR4_X1 U5337 ( .A1(REG3_REG_15__SCAN_IN), .A2(DATAI_14_), .A3(DATAI_12_), 
        .A4(DATAI_11_), .ZN(n4842) );
  NAND4_X1 U5338 ( .A1(n4845), .A2(n4844), .A3(n4843), .A4(n4842), .ZN(n4846)
         );
  NOR4_X1 U5339 ( .A1(n4849), .A2(n4848), .A3(n4847), .A4(n4846), .ZN(n4850)
         );
  NAND4_X1 U5340 ( .A1(n4853), .A2(n4852), .A3(n4851), .A4(n4850), .ZN(n4854)
         );
  XNOR2_X1 U5341 ( .A(n4855), .B(n4854), .ZN(U3479) );
endmodule

