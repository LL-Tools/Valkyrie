

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4261, n4262, n4263, n4264, n4265, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936;

  NOR2_X1 U4766 ( .A1(n8125), .A2(n8126), .ZN(n8124) );
  XNOR2_X1 U4767 ( .A(n8306), .B(n8132), .ZN(n8118) );
  NAND2_X1 U4768 ( .A1(n6956), .A2(n4614), .ZN(n4608) );
  CLKBUF_X1 U4769 ( .A(n6329), .Z(n7642) );
  INV_X2 U4770 ( .A(n7675), .ZN(n7762) );
  INV_X1 U4771 ( .A(n5678), .ZN(n7235) );
  INV_X1 U4772 ( .A(n7248), .ZN(n7080) );
  INV_X1 U4773 ( .A(n6026), .ZN(n6341) );
  INV_X4 U4774 ( .A(n5461), .ZN(n7244) );
  XNOR2_X1 U4775 ( .A(n4904), .B(SI_1_), .ZN(n4934) );
  INV_X1 U4776 ( .A(n7391), .ZN(n7384) );
  INV_X1 U4777 ( .A(n7040), .ZN(n4759) );
  INV_X1 U4778 ( .A(n6976), .ZN(n7079) );
  OAI21_X1 U4779 ( .B1(n6471), .B2(n7399), .A(n6470), .ZN(n6472) );
  INV_X1 U4780 ( .A(n6011), .ZN(n7538) );
  AND2_X1 U4781 ( .A1(n5415), .A2(n4294), .ZN(n6703) );
  INV_X1 U4782 ( .A(n5579), .ZN(n7222) );
  NAND2_X1 U4783 ( .A1(n5185), .A2(n5186), .ZN(n5669) );
  INV_X1 U4784 ( .A(n7678), .ZN(n7485) );
  NAND2_X1 U4785 ( .A1(n6878), .A2(n6877), .ZN(n6956) );
  AND2_X1 U4786 ( .A1(n5405), .A2(n5404), .ZN(n5786) );
  INV_X1 U4787 ( .A(n9501), .ZN(n6314) );
  OR2_X1 U4788 ( .A1(n6820), .A2(n8752), .ZN(n6939) );
  INV_X1 U4789 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n4835) );
  OR2_X1 U4790 ( .A1(n8424), .A2(n7697), .ZN(n8497) );
  NAND2_X1 U4791 ( .A1(n8610), .A2(n8609), .ZN(n9122) );
  AND2_X1 U4792 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n6692) );
  AND4_X1 U4793 ( .A1(n5558), .A2(n5557), .A3(n5556), .A4(n5559), .ZN(n8257)
         );
  XNOR2_X1 U4794 ( .A(n4874), .B(n4873), .ZN(n5370) );
  NAND2_X1 U4795 ( .A1(n5415), .A2(n6079), .ZN(n4261) );
  OAI21_X2 U4796 ( .B1(n7739), .B2(n8683), .A(n8642), .ZN(n9110) );
  OAI22_X2 U4797 ( .A1(n5745), .A2(n5744), .B1(n5691), .B2(n5690), .ZN(n9551)
         );
  INV_X4 U4798 ( .A(n6455), .ZN(n5576) );
  OAI21_X2 U4799 ( .B1(n8414), .B2(n8416), .A(n8415), .ZN(n7625) );
  INV_X1 U4800 ( .A(n4261), .ZN(n4262) );
  INV_X4 U4801 ( .A(n4261), .ZN(n4263) );
  INV_X2 U4802 ( .A(n9606), .ZN(n5718) );
  OR2_X1 U4803 ( .A1(n5452), .A2(n8727), .ZN(n4264) );
  OR2_X1 U4804 ( .A1(n5452), .A2(n8727), .ZN(n9519) );
  NOR3_X1 U4805 ( .A1(n4391), .A2(n8717), .A3(n4306), .ZN(n4390) );
  OAI22_X1 U4806 ( .A1(n7231), .A2(n4697), .B1(n4696), .B2(n7232), .ZN(n7241)
         );
  AND2_X1 U4807 ( .A1(n7863), .A2(n4295), .ZN(n4635) );
  NAND2_X1 U4808 ( .A1(n7070), .A2(n7069), .ZN(n8342) );
  NAND2_X1 U4809 ( .A1(n5882), .A2(n9480), .ZN(n8654) );
  NAND2_X1 U4810 ( .A1(n9488), .A2(n8820), .ZN(n6357) );
  NOR2_X1 U4811 ( .A1(n8823), .A2(n9427), .ZN(n6096) );
  NAND2_X1 U4812 ( .A1(n8817), .A2(n9511), .ZN(n8529) );
  INV_X1 U4813 ( .A(n8822), .ZN(n5882) );
  OAI211_X1 U4814 ( .C1(n6322), .C2(n5771), .A(n5770), .B(n5769), .ZN(n5784)
         );
  INV_X2 U4815 ( .A(n6011), .ZN(n4265) );
  INV_X1 U4816 ( .A(n9610), .ZN(n9669) );
  INV_X1 U4817 ( .A(n5887), .ZN(n9427) );
  INV_X1 U4818 ( .A(n8628), .ZN(n4267) );
  OAI211_X1 U4819 ( .C1(n6976), .C2(n5682), .A(n5681), .B(n5680), .ZN(n6309)
         );
  CLKBUF_X2 U4820 ( .A(n5577), .Z(n7228) );
  NAND2_X2 U4821 ( .A1(n5669), .A2(n7244), .ZN(n7248) );
  INV_X2 U4822 ( .A(n4913), .ZN(n5461) );
  AND2_X1 U4823 ( .A1(n4605), .A2(n4604), .ZN(n8454) );
  AND2_X1 U4824 ( .A1(n7456), .A2(n7455), .ZN(n4813) );
  NOR2_X1 U4825 ( .A1(n9126), .A2(n4416), .ZN(n4746) );
  NAND2_X1 U4826 ( .A1(n4390), .A2(n4724), .ZN(n8719) );
  AOI21_X1 U4827 ( .B1(n8930), .B2(n9117), .A(n8929), .ZN(n9134) );
  AND2_X1 U4828 ( .A1(n8623), .A2(n8619), .ZN(n8767) );
  NAND2_X1 U4829 ( .A1(n8168), .A2(n4579), .ZN(n8142) );
  AOI21_X1 U4830 ( .B1(n4796), .B2(n4276), .A(n4794), .ZN(n4793) );
  NAND2_X1 U4831 ( .A1(n7250), .A2(n7249), .ZN(n8272) );
  OAI21_X1 U4832 ( .B1(n4382), .B2(n8628), .A(n4381), .ZN(n8576) );
  NAND2_X1 U4833 ( .A1(n4606), .A2(n4609), .ZN(n8433) );
  NAND2_X1 U4834 ( .A1(n4594), .A2(n4592), .ZN(n6876) );
  NAND2_X1 U4835 ( .A1(n7144), .A2(n7143), .ZN(n8301) );
  AOI21_X1 U4836 ( .B1(n4629), .B2(n4634), .A(n4319), .ZN(n4627) );
  XNOR2_X1 U4837 ( .A(n6918), .B(n6917), .ZN(n7679) );
  NAND2_X1 U4838 ( .A1(n4720), .A2(n6832), .ZN(n6918) );
  AOI21_X1 U4839 ( .B1(n4635), .B2(n4633), .A(n7820), .ZN(n4632) );
  OR2_X1 U4840 ( .A1(n6500), .A2(n4730), .ZN(n4726) );
  NAND2_X1 U4841 ( .A1(n5824), .A2(n5823), .ZN(n5832) );
  NAND2_X1 U4842 ( .A1(n8779), .A2(n8644), .ZN(n6621) );
  NAND2_X1 U4843 ( .A1(n6979), .A2(n6978), .ZN(n7976) );
  NAND2_X1 U4844 ( .A1(n6804), .A2(n6803), .ZN(n9205) );
  NAND2_X1 U4845 ( .A1(n6891), .A2(n6890), .ZN(n9352) );
  NAND2_X2 U4846 ( .A1(n5965), .A2(n8238), .ZN(n8265) );
  NAND2_X1 U4847 ( .A1(n6764), .A2(n6763), .ZN(n6972) );
  AND2_X1 U4848 ( .A1(n7303), .A2(n7306), .ZN(n7407) );
  NAND2_X1 U4849 ( .A1(n6279), .A2(n6278), .ZN(n9703) );
  INV_X1 U4850 ( .A(n6067), .ZN(n9495) );
  NAND2_X1 U4851 ( .A1(n4312), .A2(n5413), .ZN(n8823) );
  AND2_X2 U4852 ( .A1(n5121), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  AND2_X1 U4853 ( .A1(n4424), .A2(n4422), .ZN(n6067) );
  OAI211_X1 U4854 ( .C1(n6322), .C2(n6148), .A(n6147), .B(n6146), .ZN(n9501)
         );
  AND3_X1 U4855 ( .A1(n5650), .A2(n5649), .A3(n4397), .ZN(n6090) );
  INV_X2 U4856 ( .A(n7497), .ZN(n6011) );
  NAND2_X1 U4857 ( .A1(n5658), .A2(n5657), .ZN(n8821) );
  NAND4_X1 U4858 ( .A1(n5993), .A2(n5992), .A3(n5991), .A4(n5990), .ZN(n8819)
         );
  CLKBUF_X1 U4859 ( .A(n6703), .Z(n7484) );
  AND2_X2 U4860 ( .A1(n5416), .A2(n5415), .ZN(n7497) );
  NAND4_X1 U4861 ( .A1(n5688), .A2(n5687), .A3(n5686), .A4(n5685), .ZN(n7994)
         );
  AOI21_X1 U4862 ( .B1(n4706), .B2(n4708), .A(n4704), .ZN(n4703) );
  INV_X2 U4863 ( .A(n7982), .ZN(P2_U3966) );
  INV_X1 U4864 ( .A(n6329), .ZN(n6322) );
  INV_X2 U4865 ( .A(n7635), .ZN(n7591) );
  CLKBUF_X3 U4866 ( .A(n5496), .Z(n8615) );
  OAI21_X1 U4867 ( .B1(n6932), .B2(n5420), .A(n5418), .ZN(n5887) );
  NAND2_X2 U4868 ( .A1(n5456), .A2(n6079), .ZN(n7675) );
  INV_X2 U4869 ( .A(n5712), .ZN(n7168) );
  CLKBUF_X1 U4870 ( .A(n5463), .Z(n6932) );
  AND2_X1 U4871 ( .A1(n9269), .A2(n5403), .ZN(n5496) );
  NAND2_X1 U4872 ( .A1(n4817), .A2(n4440), .ZN(n9644) );
  NAND2_X1 U4873 ( .A1(n8773), .A2(n5414), .ZN(n5452) );
  NAND2_X1 U4874 ( .A1(n4759), .A2(n5086), .ZN(n5696) );
  NAND2_X1 U4875 ( .A1(n8794), .A2(n8772), .ZN(n6079) );
  AND2_X2 U4876 ( .A1(n9639), .A2(n8286), .ZN(n9606) );
  XNOR2_X1 U4877 ( .A(n4865), .B(n4864), .ZN(n5414) );
  NAND2_X1 U4878 ( .A1(n5402), .A2(n5401), .ZN(n5405) );
  NAND2_X1 U4879 ( .A1(n4895), .A2(n4894), .ZN(n5603) );
  INV_X1 U4880 ( .A(n5404), .ZN(n9269) );
  MUX2_X1 U4881 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4890), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n4891) );
  AND2_X1 U4882 ( .A1(n4869), .A2(n4868), .ZN(n8794) );
  MUX2_X1 U4883 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5400), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5402) );
  NAND2_X1 U4884 ( .A1(n4868), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4865) );
  XNOR2_X1 U4885 ( .A(n5399), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5404) );
  MUX2_X1 U4886 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4893), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n4895) );
  XNOR2_X1 U4887 ( .A(n5393), .B(n5392), .ZN(n8772) );
  NAND2_X1 U4888 ( .A1(n5076), .A2(n5075), .ZN(n5077) );
  OAI21_X1 U4889 ( .B1(n5391), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n4867) );
  NAND2_X1 U4890 ( .A1(n5078), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5079) );
  INV_X2 U4891 ( .A(n6509), .ZN(n4268) );
  OR2_X2 U4892 ( .A1(n7244), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9275) );
  XNOR2_X1 U4893 ( .A(n4920), .B(SI_4_), .ZN(n4936) );
  NOR2_X1 U4894 ( .A1(n4860), .A2(n4861), .ZN(n4872) );
  XNOR2_X1 U4895 ( .A(n4935), .B(P2_IR_REG_1__SCAN_IN), .ZN(n9282) );
  NAND2_X1 U4896 ( .A1(n6692), .A2(n4899), .ZN(n4900) );
  NOR2_X1 U4897 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n6693) );
  INV_X1 U4898 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4734) );
  INV_X4 U4899 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U4900 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n4864) );
  NOR2_X1 U4901 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4857) );
  INV_X1 U4902 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5541) );
  INV_X1 U4903 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4836) );
  INV_X4 U4904 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NOR2_X1 U4905 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n4760) );
  AND2_X1 U4906 ( .A1(n5463), .A2(n7244), .ZN(n6329) );
  NAND3_X2 U4907 ( .A1(n6019), .A2(n6024), .A3(n6018), .ZN(n6414) );
  INV_X2 U4908 ( .A(n9606), .ZN(n4269) );
  OAI211_X2 U4909 ( .C1(n6322), .C2(n6321), .A(n6320), .B(n6319), .ZN(n8380)
         );
  AND2_X1 U4910 ( .A1(n7332), .A2(n7331), .ZN(n4469) );
  NAND2_X1 U4911 ( .A1(n9594), .A2(n4789), .ZN(n4792) );
  NOR2_X1 U4912 ( .A1(n7414), .A2(n4790), .ZN(n4789) );
  INV_X1 U4913 ( .A(n6780), .ZN(n4790) );
  NAND2_X1 U4914 ( .A1(n4830), .A2(n4478), .ZN(n4477) );
  INV_X1 U4915 ( .A(n5405), .ZN(n5403) );
  NAND2_X1 U4916 ( .A1(n4882), .A2(n4881), .ZN(n4399) );
  NAND2_X1 U4917 ( .A1(n4854), .A2(n4853), .ZN(n4992) );
  INV_X2 U4918 ( .A(n5463), .ZN(n7566) );
  AND2_X1 U4919 ( .A1(n4757), .A2(n4889), .ZN(n4755) );
  AND2_X2 U4920 ( .A1(n4984), .A2(n4852), .ZN(n4854) );
  INV_X1 U4921 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n4852) );
  NAND2_X1 U4922 ( .A1(n4469), .A2(n4313), .ZN(n4468) );
  NAND2_X1 U4923 ( .A1(n8576), .A2(n8569), .ZN(n4380) );
  NOR2_X1 U4924 ( .A1(n8074), .A2(n7253), .ZN(n4554) );
  NAND2_X1 U4925 ( .A1(n7230), .A2(n4307), .ZN(n4552) );
  NAND2_X1 U4926 ( .A1(n4324), .A2(n7386), .ZN(n4551) );
  NAND2_X1 U4927 ( .A1(n8822), .A2(n6090), .ZN(n8655) );
  NOR2_X1 U4928 ( .A1(n9215), .A2(n8813), .ZN(n4515) );
  AND2_X1 U4929 ( .A1(n4733), .A2(n6586), .ZN(n4732) );
  NAND2_X1 U4930 ( .A1(n6499), .A2(n6498), .ZN(n4733) );
  NAND2_X1 U4931 ( .A1(n4961), .A2(SI_7_), .ZN(n4965) );
  OR2_X1 U4932 ( .A1(n4646), .A2(n4643), .ZN(n4641) );
  NAND2_X1 U4933 ( .A1(n5549), .A2(n5963), .ZN(n5673) );
  OR2_X1 U4934 ( .A1(n8081), .A2(n7252), .ZN(n7389) );
  OR2_X1 U4935 ( .A1(n8287), .A2(n7884), .ZN(n7385) );
  NAND2_X1 U4936 ( .A1(n8104), .A2(n7901), .ZN(n4807) );
  OR2_X1 U4937 ( .A1(n8296), .A2(n7962), .ZN(n7378) );
  OR2_X1 U4938 ( .A1(n8306), .A2(n8132), .ZN(n4808) );
  OR2_X1 U4939 ( .A1(n8310), .A2(n7903), .ZN(n7368) );
  OR2_X1 U4940 ( .A1(n8327), .A2(n8199), .ZN(n7112) );
  NOR2_X1 U4941 ( .A1(n4780), .A2(n7418), .ZN(n4779) );
  INV_X1 U4942 ( .A(n4782), .ZN(n4780) );
  NOR2_X1 U4943 ( .A1(n4785), .A2(n7056), .ZN(n4784) );
  OR2_X1 U4944 ( .A1(n9693), .A2(n6519), .ZN(n7304) );
  OR2_X1 U4945 ( .A1(n9131), .A2(n8953), .ZN(n8728) );
  NAND2_X1 U4946 ( .A1(n9131), .A2(n8953), .ZN(n8909) );
  NAND2_X1 U4947 ( .A1(n8977), .A2(n4305), .ZN(n4412) );
  OR2_X1 U4948 ( .A1(n9141), .A2(n8952), .ZN(n8782) );
  NAND2_X1 U4949 ( .A1(n9148), .A2(n8501), .ZN(n8704) );
  OR2_X1 U4950 ( .A1(n9157), .A2(n8474), .ZN(n8730) );
  INV_X1 U4951 ( .A(n4492), .ZN(n4490) );
  AND2_X1 U4952 ( .A1(n6361), .A2(n6382), .ZN(n8737) );
  OR2_X1 U4953 ( .A1(n8944), .A2(n9131), .ZN(n8932) );
  XNOR2_X1 U4954 ( .A(n7241), .B(n7240), .ZN(n7238) );
  NOR2_X1 U4955 ( .A1(n4758), .A2(n4311), .ZN(n4757) );
  AND2_X1 U4956 ( .A1(n5871), .A2(n5837), .ZN(n5869) );
  AND2_X1 U4957 ( .A1(n5114), .A2(n5101), .ZN(n5112) );
  AND2_X1 U4958 ( .A1(n4347), .A2(n5016), .ZN(n5013) );
  AND2_X1 U4959 ( .A1(n4996), .A2(n4995), .ZN(n4997) );
  INV_X1 U4960 ( .A(n4999), .ZN(n5015) );
  NAND2_X1 U4961 ( .A1(n5566), .A2(n4903), .ZN(n4904) );
  NAND2_X1 U4962 ( .A1(n5548), .A2(n5547), .ZN(n7427) );
  AOI21_X1 U4963 ( .B1(n4470), .B2(n7395), .A(n7394), .ZN(n7396) );
  INV_X1 U4964 ( .A(n5696), .ZN(n5712) );
  NAND2_X1 U4965 ( .A1(n7040), .A2(n5086), .ZN(n6455) );
  NAND2_X1 U4966 ( .A1(n8130), .A2(n7368), .ZN(n8117) );
  NAND2_X1 U4967 ( .A1(n8142), .A2(n4577), .ZN(n8130) );
  NOR2_X1 U4968 ( .A1(n8127), .A2(n4578), .ZN(n4577) );
  INV_X1 U4969 ( .A(n7189), .ZN(n4578) );
  XNOR2_X1 U4970 ( .A(n8317), .B(n8166), .ZN(n8146) );
  OR2_X1 U4971 ( .A1(n8338), .A2(n8229), .ZN(n7089) );
  OR2_X1 U4972 ( .A1(n9352), .A2(n7972), .ZN(n7329) );
  OR2_X1 U4973 ( .A1(n9352), .A2(n7985), .ZN(n6973) );
  NAND2_X1 U4974 ( .A1(n6972), .A2(n7986), .ZN(n4791) );
  NAND2_X1 U4975 ( .A1(n5941), .A2(n4773), .ZN(n4772) );
  NOR2_X1 U4976 ( .A1(n7407), .A2(n4774), .ZN(n4773) );
  AND2_X1 U4977 ( .A1(n5961), .A2(n7253), .ZN(n9639) );
  NAND2_X1 U4978 ( .A1(n4473), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5059) );
  AND2_X1 U4979 ( .A1(n7578), .A2(n7577), .ZN(n7580) );
  NAND2_X1 U4980 ( .A1(n5459), .A2(n5458), .ZN(n5472) );
  XNOR2_X1 U4981 ( .A(n4582), .B(n7675), .ZN(n5778) );
  OAI21_X1 U4982 ( .B1(n6957), .B2(n5882), .A(n5651), .ZN(n4582) );
  OR2_X1 U4983 ( .A1(n9136), .A2(n8899), .ZN(n8908) );
  AND2_X1 U4984 ( .A1(n7653), .A2(n7652), .ZN(n8399) );
  NOR2_X1 U4985 ( .A1(n8932), .A2(n9128), .ZN(n8915) );
  NAND2_X1 U4986 ( .A1(n8901), .A2(n4524), .ZN(n8925) );
  NOR2_X1 U4987 ( .A1(n8922), .A2(n4525), .ZN(n4524) );
  INV_X1 U4988 ( .A(n8900), .ZN(n4525) );
  INV_X1 U4989 ( .A(n8896), .ZN(n8952) );
  OR2_X1 U4990 ( .A1(n9148), .A2(n8501), .ZN(n8781) );
  OR2_X1 U4991 ( .A1(n7665), .A2(n7664), .ZN(n7683) );
  AND2_X1 U4992 ( .A1(n9005), .A2(n8994), .ZN(n8990) );
  OR2_X1 U4993 ( .A1(n9161), .A2(n8808), .ZN(n7730) );
  INV_X1 U4994 ( .A(n9014), .ZN(n9041) );
  NAND2_X1 U4995 ( .A1(n7512), .A2(n7511), .ZN(n9195) );
  NAND2_X1 U4996 ( .A1(n5401), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5399) );
  XNOR2_X1 U4997 ( .A(n6834), .B(n6833), .ZN(n7661) );
  INV_X1 U4998 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4851) );
  OAI21_X1 U4999 ( .B1(n8067), .B2(n9576), .A(n4676), .ZN(n4675) );
  AOI21_X1 U5000 ( .B1(n8068), .B2(n9573), .A(n9295), .ZN(n4676) );
  INV_X1 U5001 ( .A(n7704), .ZN(n4584) );
  NOR2_X1 U5002 ( .A1(n7704), .A2(n7703), .ZN(n4585) );
  NAND2_X1 U5003 ( .A1(n4725), .A2(n8628), .ZN(n4724) );
  OAI22_X1 U5004 ( .A1(n8627), .A2(n8626), .B1(n8625), .B2(n8786), .ZN(n4725)
         );
  NAND2_X1 U5005 ( .A1(n4364), .A2(n4361), .ZN(n4360) );
  OR2_X1 U5006 ( .A1(n8877), .A2(n8855), .ZN(n4364) );
  INV_X1 U5007 ( .A(n4362), .ZN(n4361) );
  OAI21_X1 U5008 ( .B1(n8879), .B2(n8878), .A(n4363), .ZN(n4362) );
  NAND2_X1 U5009 ( .A1(n4450), .A2(n7391), .ZN(n4451) );
  AOI21_X1 U5010 ( .B1(n8533), .B2(n4292), .A(n4395), .ZN(n4394) );
  OR2_X1 U5011 ( .A1(n7326), .A2(n4467), .ZN(n4466) );
  NAND2_X1 U5012 ( .A1(n4468), .A2(n7391), .ZN(n4467) );
  OR2_X1 U5013 ( .A1(n7325), .A2(n4465), .ZN(n4464) );
  NAND2_X1 U5014 ( .A1(n4468), .A2(n7384), .ZN(n4465) );
  AOI21_X1 U5015 ( .B1(n4379), .B2(n4378), .A(n4318), .ZN(n8575) );
  NOR2_X1 U5016 ( .A1(n8570), .A2(n4406), .ZN(n4378) );
  NAND2_X1 U5017 ( .A1(n4380), .A2(n8579), .ZN(n4379) );
  AOI21_X1 U5018 ( .B1(n4460), .B2(n4459), .A(n4458), .ZN(n7375) );
  INV_X1 U5019 ( .A(n7372), .ZN(n4458) );
  AND2_X1 U5020 ( .A1(n7373), .A2(n7371), .ZN(n4459) );
  OR2_X1 U5021 ( .A1(n8272), .A2(n7251), .ZN(n7390) );
  NAND2_X1 U5022 ( .A1(n8748), .A2(n4287), .ZN(n4522) );
  NAND2_X1 U5023 ( .A1(n5021), .A2(n5020), .ZN(n5035) );
  NAND2_X1 U5024 ( .A1(n6598), .A2(n6599), .ZN(n4653) );
  AOI21_X1 U5025 ( .B1(n7889), .B2(n7890), .A(n7826), .ZN(n7827) );
  AND2_X1 U5026 ( .A1(n7825), .A2(n7824), .ZN(n7826) );
  NOR2_X1 U5027 ( .A1(n8257), .A2(n9606), .ZN(n5560) );
  NAND2_X1 U5028 ( .A1(n4550), .A2(n4280), .ZN(n4548) );
  OAI21_X1 U5029 ( .B1(n4472), .B2(n4471), .A(n4304), .ZN(n4470) );
  NAND2_X1 U5030 ( .A1(n7449), .A2(n4279), .ZN(n4471) );
  AOI21_X1 U5031 ( .B1(n7382), .B2(n7381), .A(n7380), .ZN(n4472) );
  INV_X1 U5032 ( .A(n7756), .ZN(n5086) );
  NOR2_X1 U5033 ( .A1(n4566), .A2(n4562), .ZN(n4561) );
  INV_X1 U5034 ( .A(n7190), .ZN(n4562) );
  OAI21_X1 U5035 ( .B1(n4803), .B2(n4566), .A(n8091), .ZN(n4565) );
  AND2_X1 U5036 ( .A1(n4798), .A2(n4797), .ZN(n4796) );
  INV_X1 U5037 ( .A(n8091), .ZN(n4797) );
  OR2_X1 U5038 ( .A1(n8301), .A2(n7901), .ZN(n7373) );
  INV_X1 U5039 ( .A(n8310), .ZN(n7175) );
  AND2_X1 U5040 ( .A1(n7260), .A2(n7259), .ZN(n7418) );
  OR2_X1 U5041 ( .A1(n7976), .A2(n7915), .ZN(n7334) );
  INV_X1 U5042 ( .A(n7293), .ZN(n4559) );
  OR2_X1 U5043 ( .A1(n7993), .A2(n9669), .ZN(n7272) );
  OR2_X1 U5044 ( .A1(n9623), .A2(n9663), .ZN(n7269) );
  INV_X1 U5045 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4776) );
  AND3_X1 U5046 ( .A1(n4826), .A2(n4827), .A3(n4828), .ZN(n4441) );
  NOR2_X1 U5047 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n4827) );
  NOR2_X1 U5048 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n4828) );
  AND4_X1 U5049 ( .A1(n4825), .A2(n5117), .A3(n5026), .A4(n4973), .ZN(n4829)
         );
  NOR2_X1 U5050 ( .A1(n8767), .A2(n8889), .ZN(n8622) );
  NAND2_X1 U5051 ( .A1(n4357), .A2(n4356), .ZN(n5129) );
  INV_X1 U5052 ( .A(n5614), .ZN(n4356) );
  INV_X1 U5053 ( .A(n5613), .ZN(n4357) );
  NOR2_X1 U5054 ( .A1(n6853), .A2(n4543), .ZN(n6854) );
  AND2_X1 U5055 ( .A1(n6861), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4543) );
  NOR2_X1 U5056 ( .A1(n9148), .A2(n9152), .ZN(n4754) );
  OR2_X1 U5057 ( .A1(n9152), .A2(n8399), .ZN(n8776) );
  NOR2_X1 U5058 ( .A1(n4491), .A2(n4488), .ZN(n4487) );
  INV_X1 U5059 ( .A(n4494), .ZN(n4488) );
  NAND2_X1 U5060 ( .A1(n4322), .A2(n4496), .ZN(n4492) );
  INV_X1 U5061 ( .A(n4287), .ZN(n4519) );
  NOR2_X1 U5062 ( .A1(n4521), .A2(n4515), .ZN(n4514) );
  NAND2_X1 U5063 ( .A1(n4514), .A2(n6735), .ZN(n4512) );
  OR2_X1 U5064 ( .A1(n9400), .A2(n6965), .ZN(n8537) );
  AND2_X1 U5065 ( .A1(n6149), .A2(n6143), .ZN(n4528) );
  NAND2_X1 U5066 ( .A1(n4516), .A2(n4513), .ZN(n6737) );
  INV_X1 U5067 ( .A(n4515), .ZN(n4513) );
  NAND2_X1 U5068 ( .A1(n6733), .A2(n4517), .ZN(n4516) );
  AOI21_X1 U5069 ( .B1(n4716), .B2(n4719), .A(n4715), .ZN(n4714) );
  AOI21_X1 U5070 ( .B1(n5833), .B2(n5834), .A(n4701), .ZN(n4700) );
  OAI21_X1 U5071 ( .B1(n5761), .B2(n5760), .A(n5759), .ZN(n5821) );
  NOR2_X1 U5072 ( .A1(n5298), .A2(n4711), .ZN(n4710) );
  INV_X1 U5073 ( .A(n5114), .ZN(n4711) );
  INV_X1 U5074 ( .A(n5294), .ZN(n5298) );
  OAI21_X1 U5075 ( .B1(n5046), .B2(n5045), .A(n5044), .ZN(n5097) );
  NAND2_X1 U5076 ( .A1(n5095), .A2(n5049), .ZN(n5096) );
  XNOR2_X1 U5077 ( .A(n5043), .B(n9873), .ZN(n5042) );
  NAND2_X1 U5078 ( .A1(n4691), .A2(n4689), .ZN(n5046) );
  OR2_X1 U5079 ( .A1(n4998), .A2(n4692), .ZN(n4691) );
  INV_X1 U5080 ( .A(n4690), .ZN(n4689) );
  NAND2_X1 U5081 ( .A1(n4688), .A2(n5033), .ZN(n4692) );
  AOI21_X1 U5082 ( .B1(n4688), .B2(n4687), .A(n4686), .ZN(n4695) );
  INV_X1 U5083 ( .A(n5016), .ZN(n4686) );
  INV_X1 U5084 ( .A(n4997), .ZN(n4687) );
  INV_X1 U5085 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n4853) );
  AND2_X1 U5086 ( .A1(n4293), .A2(n5008), .ZN(n4619) );
  INV_X1 U5087 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n4950) );
  OAI21_X1 U5088 ( .B1(n4936), .B2(n4684), .A(n4943), .ZN(n4683) );
  INV_X1 U5089 ( .A(n4683), .ZN(n4681) );
  INV_X1 U5090 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n4919) );
  INV_X1 U5091 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4898) );
  OAI21_X1 U5092 ( .B1(n6596), .B2(n4642), .A(n4640), .ZN(n4639) );
  OR2_X1 U5093 ( .A1(n4648), .A2(n4643), .ZN(n4642) );
  AND2_X1 U5094 ( .A1(n4641), .A2(n4328), .ZN(n4640) );
  INV_X1 U5095 ( .A(n7790), .ZN(n4661) );
  NAND2_X1 U5096 ( .A1(n7244), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4439) );
  INV_X1 U5097 ( .A(n4632), .ZN(n4630) );
  NAND2_X1 U5098 ( .A1(n4651), .A2(n4653), .ZN(n4650) );
  NAND2_X1 U5099 ( .A1(n4652), .A2(n6650), .ZN(n4651) );
  NAND2_X1 U5100 ( .A1(n6595), .A2(n4654), .ZN(n4652) );
  AOI21_X1 U5101 ( .B1(n7855), .B2(n7856), .A(n7834), .ZN(n7837) );
  NAND2_X1 U5102 ( .A1(n6515), .A2(n6514), .ZN(n9564) );
  OR2_X1 U5103 ( .A1(n5577), .A2(n8264), .ZN(n5557) );
  OR2_X1 U5104 ( .A1(n8352), .A2(n5959), .ZN(n5571) );
  CLKBUF_X1 U5105 ( .A(n6455), .Z(n7224) );
  INV_X1 U5106 ( .A(n8285), .ZN(n8081) );
  NAND2_X1 U5107 ( .A1(n7237), .A2(n7236), .ZN(n8287) );
  INV_X1 U5108 ( .A(n7373), .ZN(n4566) );
  NAND2_X1 U5109 ( .A1(n4799), .A2(n4807), .ZN(n4798) );
  INV_X1 U5110 ( .A(n4802), .ZN(n4799) );
  AOI21_X1 U5111 ( .B1(n4804), .B2(n8118), .A(n4803), .ZN(n4802) );
  INV_X1 U5112 ( .A(n4807), .ZN(n4800) );
  AND2_X1 U5113 ( .A1(n7378), .A2(n7379), .ZN(n8091) );
  XNOR2_X1 U5114 ( .A(n8310), .B(n8144), .ZN(n8126) );
  OR2_X1 U5115 ( .A1(n4428), .A2(n8166), .ZN(n4818) );
  NOR2_X1 U5116 ( .A1(n8146), .A2(n4580), .ZN(n4579) );
  INV_X1 U5117 ( .A(n7348), .ZN(n4580) );
  OR2_X1 U5118 ( .A1(n8189), .A2(n8327), .ZN(n8157) );
  INV_X1 U5119 ( .A(n4764), .ZN(n4763) );
  OAI21_X1 U5120 ( .B1(n4765), .B2(n4277), .A(n7112), .ZN(n4764) );
  NAND2_X1 U5121 ( .A1(n4766), .A2(n4289), .ZN(n4765) );
  INV_X1 U5122 ( .A(n8198), .ZN(n4766) );
  OR2_X1 U5123 ( .A1(n8205), .A2(n7953), .ZN(n4811) );
  AOI21_X1 U5124 ( .B1(n4572), .B2(n4574), .A(n4571), .ZN(n4570) );
  INV_X1 U5125 ( .A(n4574), .ZN(n4573) );
  INV_X1 U5126 ( .A(n7183), .ZN(n4572) );
  OAI21_X1 U5127 ( .B1(n8219), .B2(n7078), .A(n4815), .ZN(n8204) );
  OR2_X1 U5128 ( .A1(n8222), .A2(n8250), .ZN(n4815) );
  AND2_X1 U5129 ( .A1(n4282), .A2(n7260), .ZN(n4574) );
  OR2_X1 U5130 ( .A1(n8349), .A2(n7954), .ZN(n7260) );
  NAND2_X1 U5131 ( .A1(n9322), .A2(n7183), .ZN(n4575) );
  AOI21_X1 U5132 ( .B1(n4784), .B2(n7332), .A(n4321), .ZN(n4782) );
  INV_X1 U5133 ( .A(n4784), .ZN(n4783) );
  NAND2_X1 U5134 ( .A1(n4792), .A2(n4297), .ZN(n9353) );
  OR2_X1 U5135 ( .A1(n6459), .A2(n6458), .ZN(n6605) );
  AND2_X1 U5136 ( .A1(n6778), .A2(n6777), .ZN(n9595) );
  NAND2_X1 U5137 ( .A1(n9595), .A2(n6779), .ZN(n9594) );
  NOR2_X1 U5138 ( .A1(n5974), .A2(n4771), .ZN(n4770) );
  INV_X1 U5139 ( .A(n5955), .ZN(n4771) );
  OR2_X1 U5140 ( .A1(n9622), .A2(n9676), .ZN(n7293) );
  NAND2_X1 U5141 ( .A1(n6121), .A2(n7405), .ZN(n6120) );
  OR2_X1 U5143 ( .A1(n7994), .A2(n9657), .ZN(n6183) );
  OR2_X1 U5144 ( .A1(n8257), .A2(n9644), .ZN(n8256) );
  NAND2_X1 U5145 ( .A1(n4436), .A2(n4435), .ZN(n4434) );
  NAND2_X1 U5146 ( .A1(n8287), .A2(n9694), .ZN(n4435) );
  OR2_X1 U5147 ( .A1(n8289), .A2(n9652), .ZN(n4436) );
  INV_X1 U5148 ( .A(n9332), .ZN(n9362) );
  INV_X1 U5149 ( .A(n6127), .ZN(n9676) );
  NOR2_X1 U5150 ( .A1(n4314), .A2(n4477), .ZN(n4476) );
  OR2_X1 U5151 ( .A1(n5540), .A2(n5539), .ZN(n5545) );
  INV_X1 U5152 ( .A(n4477), .ZN(n4475) );
  XNOR2_X1 U5153 ( .A(n5774), .B(n7675), .ZN(n6002) );
  AOI21_X1 U5154 ( .B1(n8821), .B2(n6703), .A(n5775), .ZN(n6003) );
  NAND2_X1 U5155 ( .A1(n9473), .A2(n4263), .ZN(n5468) );
  NAND2_X1 U5156 ( .A1(n8408), .A2(n7585), .ZN(n4589) );
  INV_X1 U5157 ( .A(n7585), .ZN(n4590) );
  NOR2_X1 U5158 ( .A1(n7660), .A2(n4599), .ZN(n4598) );
  NOR2_X1 U5159 ( .A1(n4600), .A2(n7640), .ZN(n4599) );
  INV_X1 U5160 ( .A(n8397), .ZN(n4600) );
  NAND2_X1 U5161 ( .A1(n4598), .A2(n4601), .ZN(n4596) );
  NOR2_X1 U5162 ( .A1(n4602), .A2(n8397), .ZN(n4601) );
  NAND2_X1 U5163 ( .A1(n4388), .A2(n4387), .ZN(n8396) );
  AOI21_X1 U5164 ( .B1(n4270), .B2(n4273), .A(n4602), .ZN(n4387) );
  INV_X1 U5165 ( .A(n7641), .ZN(n4597) );
  AND2_X1 U5166 ( .A1(n7656), .A2(n7655), .ZN(n7657) );
  OR2_X1 U5167 ( .A1(n7747), .A2(n6011), .ZN(n7656) );
  OR2_X1 U5168 ( .A1(n6155), .A2(n6154), .ZN(n6339) );
  NAND2_X1 U5169 ( .A1(n7497), .A2(n8823), .ZN(n5424) );
  INV_X1 U5170 ( .A(n5421), .ZN(n4485) );
  AND2_X1 U5171 ( .A1(n7600), .A2(n7601), .ZN(n8461) );
  OR2_X1 U5172 ( .A1(n6623), .A2(n6622), .ZN(n6743) );
  NAND2_X1 U5173 ( .A1(n6697), .A2(n6696), .ZN(n4594) );
  NAND2_X1 U5174 ( .A1(n6368), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6574) );
  INV_X1 U5175 ( .A(n6370), .ZN(n6368) );
  AOI21_X1 U5176 ( .B1(n7506), .B2(n4613), .A(n4316), .ZN(n4371) );
  INV_X1 U5177 ( .A(n7506), .ZN(n4372) );
  AND2_X1 U5178 ( .A1(n7508), .A2(n4610), .ZN(n4609) );
  NAND2_X1 U5179 ( .A1(n5414), .A2(n8917), .ZN(n8628) );
  INV_X1 U5180 ( .A(n8772), .ZN(n8727) );
  AND2_X1 U5181 ( .A1(n8782), .A2(n8781), .ZN(n8906) );
  AND3_X1 U5182 ( .A1(n7483), .A2(n7482), .A3(n7481), .ZN(n8474) );
  NAND2_X1 U5183 ( .A1(n5496), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5654) );
  NAND2_X1 U5184 ( .A1(n5334), .A2(n5335), .ZN(n5333) );
  OR2_X1 U5185 ( .A1(n5164), .A2(n5165), .ZN(n4359) );
  NOR2_X1 U5186 ( .A1(n5516), .A2(n4538), .ZN(n5519) );
  NOR2_X1 U5187 ( .A1(n5348), .A2(n4539), .ZN(n4538) );
  INV_X1 U5188 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n4539) );
  NOR2_X1 U5189 ( .A1(n5519), .A2(n5518), .ZN(n5848) );
  OR2_X1 U5190 ( .A1(n7012), .A2(n7011), .ZN(n4537) );
  NAND2_X1 U5191 ( .A1(n9417), .A2(n4353), .ZN(n7013) );
  OR2_X1 U5192 ( .A1(n9412), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n4353) );
  OR2_X1 U5193 ( .A1(n8841), .A2(n8840), .ZN(n4350) );
  INV_X1 U5194 ( .A(n8912), .ZN(n4421) );
  AND2_X1 U5195 ( .A1(n4412), .A2(n4411), .ZN(n8950) );
  NOR2_X1 U5196 ( .A1(n4413), .A2(n8951), .ZN(n4411) );
  NAND2_X1 U5197 ( .A1(n4501), .A2(n4499), .ZN(n8941) );
  AOI21_X1 U5198 ( .B1(n4502), .B2(n4504), .A(n4500), .ZN(n4499) );
  NOR2_X1 U5199 ( .A1(n8897), .A2(n8952), .ZN(n4500) );
  NAND2_X1 U5200 ( .A1(n4272), .A2(n4308), .ZN(n4503) );
  NAND2_X1 U5201 ( .A1(n4507), .A2(n4506), .ZN(n4505) );
  NAND2_X1 U5202 ( .A1(n4272), .A2(n4507), .ZN(n4504) );
  AND2_X1 U5203 ( .A1(n4414), .A2(n8782), .ZN(n8763) );
  NAND2_X1 U5204 ( .A1(n7466), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n7665) );
  INV_X1 U5205 ( .A(n7646), .ZN(n7466) );
  AND2_X1 U5206 ( .A1(n8776), .A2(n8962), .ZN(n8978) );
  NAND2_X1 U5207 ( .A1(n8989), .A2(n7733), .ZN(n4508) );
  OR2_X1 U5208 ( .A1(n9021), .A2(n4406), .ZN(n4401) );
  INV_X1 U5209 ( .A(n4405), .ZN(n4404) );
  OAI21_X1 U5210 ( .B1(n8759), .B2(n4406), .A(n8731), .ZN(n4405) );
  NAND2_X1 U5211 ( .A1(n9029), .A2(n4816), .ZN(n9004) );
  OR2_X1 U5212 ( .A1(n9063), .A2(n9174), .ZN(n9042) );
  NOR2_X1 U5213 ( .A1(n9042), .A2(n9168), .ZN(n9019) );
  NAND2_X1 U5214 ( .A1(n8693), .A2(n8579), .ZN(n9027) );
  OR2_X1 U5215 ( .A1(n9184), .A2(n9059), .ZN(n9054) );
  NOR2_X1 U5216 ( .A1(n8810), .A2(n9205), .ZN(n6929) );
  OR2_X1 U5217 ( .A1(n6737), .A2(n8748), .ZN(n4523) );
  AND2_X1 U5218 ( .A1(n8537), .A2(n8539), .ZN(n8748) );
  OR2_X1 U5219 ( .A1(n6487), .A2(n6493), .ZN(n6489) );
  INV_X1 U5220 ( .A(n9060), .ZN(n9112) );
  AND2_X1 U5221 ( .A1(n5425), .A2(n5607), .ZN(n9114) );
  NAND2_X1 U5222 ( .A1(n8614), .A2(n8613), .ZN(n9396) );
  AND2_X1 U5223 ( .A1(n8932), .A2(n8931), .ZN(n9132) );
  NAND2_X1 U5224 ( .A1(n7681), .A2(n7680), .ZN(n9141) );
  NAND2_X1 U5225 ( .A1(n7679), .A2(n7642), .ZN(n7681) );
  NAND2_X1 U5226 ( .A1(n6935), .A2(n6934), .ZN(n9199) );
  INV_X1 U5227 ( .A(n6734), .ZN(n9215) );
  INV_X1 U5228 ( .A(n6629), .ZN(n6636) );
  NAND2_X1 U5229 ( .A1(n6843), .A2(n9505), .ZN(n9515) );
  XNOR2_X1 U5230 ( .A(n7238), .B(SI_30_), .ZN(n8611) );
  XNOR2_X1 U5231 ( .A(n7035), .B(n7034), .ZN(n7757) );
  NAND2_X1 U5232 ( .A1(n4756), .A2(n4757), .ZN(n4892) );
  NAND2_X1 U5233 ( .A1(n4374), .A2(n4373), .ZN(n4876) );
  AOI21_X1 U5234 ( .B1(n4376), .B2(n5306), .A(n5306), .ZN(n4373) );
  INV_X1 U5235 ( .A(n4377), .ZN(n4376) );
  NAND2_X1 U5236 ( .A1(n4726), .A2(n4727), .ZN(n6716) );
  AND2_X1 U5237 ( .A1(n6588), .A2(n6505), .ZN(n6586) );
  NAND2_X1 U5238 ( .A1(n4699), .A2(n5834), .ZN(n5870) );
  OR2_X1 U5239 ( .A1(n5832), .A2(n5833), .ZN(n4699) );
  OAI21_X1 U5240 ( .B1(n5115), .B2(n4708), .A(n4706), .ZN(n5486) );
  AND2_X1 U5241 ( .A1(n4998), .A2(n4997), .ZN(n5018) );
  INV_X1 U5242 ( .A(n4933), .ZN(n4685) );
  NOR2_X1 U5243 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n4941) );
  AOI21_X1 U5244 ( .B1(n4624), .B2(n4626), .A(n4338), .ZN(n4621) );
  XNOR2_X1 U5245 ( .A(n7874), .B(n7872), .ZN(n7876) );
  NAND2_X1 U5246 ( .A1(n7156), .A2(n7155), .ZN(n8296) );
  AND3_X1 U5247 ( .A1(n7050), .A2(n7049), .A3(n7048), .ZN(n7903) );
  NAND2_X1 U5248 ( .A1(n7133), .A2(n7132), .ZN(n8306) );
  NAND2_X1 U5249 ( .A1(n7661), .A2(n7235), .ZN(n7133) );
  XNOR2_X1 U5250 ( .A(n7837), .B(n7835), .ZN(n7927) );
  INV_X1 U5251 ( .A(n7985), .ZN(n7972) );
  INV_X1 U5252 ( .A(n7978), .ZN(n9566) );
  INV_X1 U5253 ( .A(n7983), .ZN(n8248) );
  OAI211_X1 U5254 ( .C1(n7431), .C2(n4457), .A(n4456), .B(n4455), .ZN(n4454)
         );
  NAND2_X1 U5255 ( .A1(n7434), .A2(n7433), .ZN(n4455) );
  INV_X1 U5256 ( .A(n7432), .ZN(n4457) );
  INV_X1 U5257 ( .A(n4669), .ZN(n8057) );
  OR2_X1 U5258 ( .A1(n8072), .A2(n8071), .ZN(n4673) );
  NAND2_X1 U5259 ( .A1(n4437), .A2(n4432), .ZN(n8357) );
  NAND2_X1 U5260 ( .A1(n8288), .A2(n9606), .ZN(n4437) );
  NOR2_X1 U5261 ( .A1(n4434), .A2(n4433), .ZN(n4432) );
  INV_X1 U5262 ( .A(n4813), .ZN(n4433) );
  NAND2_X1 U5263 ( .A1(n5065), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5067) );
  XNOR2_X1 U5264 ( .A(n5059), .B(n5058), .ZN(n5961) );
  NAND2_X1 U5265 ( .A1(n7462), .A2(n7461), .ZN(n9136) );
  INV_X1 U5266 ( .A(n8994), .ZN(n9157) );
  INV_X1 U5267 ( .A(n9068), .ZN(n9179) );
  NOR2_X1 U5268 ( .A1(n8454), .A2(n8453), .ZN(n8452) );
  NAND2_X1 U5269 ( .A1(n7628), .A2(n7627), .ZN(n9161) );
  INV_X1 U5270 ( .A(n8821), .ZN(n7215) );
  AND2_X1 U5271 ( .A1(n7672), .A2(n7671), .ZN(n8501) );
  OR2_X1 U5272 ( .A1(n8493), .A2(n8494), .ZN(n7697) );
  OR3_X1 U5273 ( .A1(n5427), .A2(n5425), .A3(n9216), .ZN(n8519) );
  OR2_X1 U5274 ( .A1(n8712), .A2(n8711), .ZN(n8713) );
  OR2_X1 U5275 ( .A1(n7614), .A2(n7613), .ZN(n9014) );
  AOI22_X1 U5276 ( .A1(n5161), .A2(n5162), .B1(n5138), .B2(n5139), .ZN(n5140)
         );
  XNOR2_X1 U5277 ( .A(n7013), .B(n7014), .ZN(n6862) );
  NOR2_X1 U5278 ( .A1(n6862), .A2(n6863), .ZN(n7015) );
  NAND2_X1 U5279 ( .A1(n8873), .A2(n4348), .ZN(n8876) );
  OR2_X1 U5280 ( .A1(n8874), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n4348) );
  OAI21_X1 U5281 ( .B1(n9426), .B2(n8883), .A(n8882), .ZN(n4546) );
  INV_X1 U5282 ( .A(n9396), .ZN(n8892) );
  OAI21_X1 U5283 ( .B1(n4420), .B2(n9229), .A(n4418), .ZN(n9126) );
  INV_X1 U5284 ( .A(n4419), .ZN(n4418) );
  XNOR2_X1 U5285 ( .A(n4421), .B(n8903), .ZN(n4420) );
  OAI22_X1 U5286 ( .A1(n8953), .A2(n9060), .B1(n8914), .B2(n8913), .ZN(n4419)
         );
  NAND2_X1 U5287 ( .A1(n8925), .A2(n8902), .ZN(n8904) );
  NAND2_X1 U5288 ( .A1(n8523), .A2(n8522), .ZN(n9128) );
  INV_X1 U5289 ( .A(n4423), .ZN(n4422) );
  NAND2_X1 U5290 ( .A1(n8612), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n4424) );
  OAI21_X1 U5291 ( .B1(n5996), .B2(n6322), .A(n5995), .ZN(n4423) );
  NAND2_X1 U5292 ( .A1(n6329), .A2(n4398), .ZN(n4397) );
  NAND2_X1 U5293 ( .A1(n5426), .A2(n8723), .ZN(n9436) );
  XNOR2_X1 U5294 ( .A(n5390), .B(n4863), .ZN(n9026) );
  INV_X1 U5295 ( .A(n5388), .ZN(n5389) );
  OAI21_X1 U5296 ( .B1(n7270), .B2(n7271), .A(n4281), .ZN(n4450) );
  NAND2_X1 U5297 ( .A1(n7275), .A2(n7270), .ZN(n7286) );
  NAND2_X1 U5298 ( .A1(n8535), .A2(n8747), .ZN(n4395) );
  NAND2_X1 U5299 ( .A1(n4468), .A2(n4463), .ZN(n4462) );
  NAND2_X1 U5300 ( .A1(n4469), .A2(n7414), .ZN(n4463) );
  NAND2_X1 U5301 ( .A1(n8567), .A2(n8628), .ZN(n4381) );
  INV_X1 U5302 ( .A(n8568), .ZN(n4382) );
  INV_X1 U5303 ( .A(n4554), .ZN(n4549) );
  INV_X1 U5304 ( .A(n8471), .ZN(n4389) );
  NAND2_X1 U5305 ( .A1(n9091), .A2(n8486), .ZN(n4496) );
  NOR2_X1 U5306 ( .A1(n7233), .A2(SI_29_), .ZN(n4697) );
  INV_X1 U5307 ( .A(n7233), .ZN(n4696) );
  INV_X1 U5308 ( .A(n7000), .ZN(n4715) );
  AND2_X1 U5309 ( .A1(n4722), .A2(n6917), .ZN(n4721) );
  NAND2_X1 U5310 ( .A1(n6833), .A2(n6832), .ZN(n4722) );
  INV_X1 U5311 ( .A(n5869), .ZN(n4701) );
  INV_X1 U5312 ( .A(n5485), .ZN(n4704) );
  NAND2_X1 U5313 ( .A1(n5047), .A2(n9832), .ZN(n5095) );
  NAND2_X1 U5314 ( .A1(n5001), .A2(n5000), .ZN(n5016) );
  INV_X1 U5315 ( .A(n6897), .ZN(n4643) );
  INV_X1 U5316 ( .A(n5673), .ZN(n7803) );
  AND2_X1 U5317 ( .A1(n5961), .A2(n5547), .ZN(n4479) );
  NOR2_X1 U5318 ( .A1(n4277), .A2(n4769), .ZN(n4762) );
  NOR2_X1 U5319 ( .A1(n4445), .A2(n8338), .ZN(n4444) );
  INV_X1 U5320 ( .A(n4446), .ZN(n4445) );
  NOR2_X1 U5321 ( .A1(n8342), .A2(n8349), .ZN(n4446) );
  AND2_X1 U5322 ( .A1(n9335), .A2(n9362), .ZN(n8234) );
  NAND2_X1 U5323 ( .A1(n5713), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5807) );
  NAND2_X1 U5324 ( .A1(n8260), .A2(n8256), .ZN(n6135) );
  NAND2_X1 U5325 ( .A1(n9596), .A2(n9380), .ZN(n9356) );
  AND2_X1 U5326 ( .A1(n9609), .A2(n9676), .ZN(n6123) );
  INV_X1 U5327 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5117) );
  INV_X1 U5328 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5026) );
  INV_X1 U5329 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n4973) );
  NAND2_X1 U5330 ( .A1(n6004), .A2(n6003), .ZN(n6016) );
  INV_X1 U5331 ( .A(n6955), .ZN(n4616) );
  NOR2_X1 U5332 ( .A1(n4612), .A2(n6881), .ZN(n4607) );
  OR2_X1 U5333 ( .A1(n7509), .A2(n4613), .ZN(n4612) );
  OR2_X1 U5334 ( .A1(n7509), .A2(n4611), .ZN(n4610) );
  NAND2_X1 U5335 ( .A1(n4615), .A2(n7488), .ZN(n4611) );
  AND2_X1 U5336 ( .A1(n4503), .A2(n4325), .ZN(n4502) );
  NOR2_X1 U5337 ( .A1(n4753), .A2(n9141), .ZN(n4752) );
  INV_X1 U5338 ( .A(n4754), .ZN(n4753) );
  INV_X1 U5339 ( .A(n7733), .ZN(n4506) );
  NAND2_X1 U5340 ( .A1(n4404), .A2(n4406), .ZN(n4402) );
  AND2_X1 U5341 ( .A1(n8730), .A2(n8995), .ZN(n8699) );
  AND2_X1 U5342 ( .A1(n4496), .A2(n9102), .ZN(n4494) );
  NAND2_X1 U5343 ( .A1(n4750), .A2(n9082), .ZN(n4749) );
  NOR2_X1 U5344 ( .A1(n9189), .A2(n9195), .ZN(n4750) );
  NOR2_X1 U5345 ( .A1(n9215), .A2(n9239), .ZN(n4739) );
  AND2_X1 U5346 ( .A1(n8671), .A2(n8674), .ZN(n8749) );
  INV_X1 U5347 ( .A(n8813), .ZN(n6739) );
  AND2_X1 U5348 ( .A1(n9222), .A2(n9231), .ZN(n9223) );
  NAND2_X1 U5349 ( .A1(n8990), .A2(n7747), .ZN(n8981) );
  AOI21_X1 U5350 ( .B1(n4721), .B2(n4718), .A(n4717), .ZN(n4716) );
  INV_X1 U5351 ( .A(n6919), .ZN(n4717) );
  INV_X1 U5352 ( .A(n6832), .ZN(n4718) );
  INV_X1 U5353 ( .A(n4721), .ZN(n4719) );
  OAI21_X1 U5354 ( .B1(n4886), .B2(n5306), .A(n4880), .ZN(n4377) );
  NAND2_X1 U5355 ( .A1(n4526), .A2(n4872), .ZN(n4758) );
  AND2_X1 U5356 ( .A1(n4870), .A2(n4527), .ZN(n4526) );
  AND2_X1 U5357 ( .A1(n4871), .A2(n4620), .ZN(n4527) );
  AOI21_X1 U5358 ( .B1(n4732), .B2(n4729), .A(n4728), .ZN(n4727) );
  INV_X1 U5359 ( .A(n6498), .ZN(n4729) );
  INV_X1 U5360 ( .A(n6588), .ZN(n4728) );
  INV_X1 U5361 ( .A(n4732), .ZN(n4730) );
  INV_X1 U5362 ( .A(n4707), .ZN(n4706) );
  OAI21_X1 U5363 ( .B1(n4710), .B2(n4708), .A(n5430), .ZN(n4707) );
  NAND2_X1 U5364 ( .A1(n4709), .A2(n5297), .ZN(n4708) );
  INV_X1 U5365 ( .A(n5431), .ZN(n4709) );
  OR2_X1 U5366 ( .A1(n5050), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n5105) );
  OR2_X1 U5367 ( .A1(n4967), .A2(n4966), .ZN(n4996) );
  NAND2_X1 U5368 ( .A1(n4970), .A2(SI_8_), .ZN(n4999) );
  AND2_X1 U5369 ( .A1(n7960), .A2(n4625), .ZN(n4624) );
  OR2_X1 U5370 ( .A1(n4626), .A2(n7899), .ZN(n4625) );
  INV_X1 U5371 ( .A(n7843), .ZN(n4626) );
  NAND2_X1 U5372 ( .A1(n7940), .A2(n7830), .ZN(n7833) );
  OR3_X1 U5373 ( .A1(n7166), .A2(n7848), .A3(n7882), .ZN(n7193) );
  NOR2_X1 U5374 ( .A1(n5664), .A2(n5562), .ZN(n5569) );
  AND2_X1 U5375 ( .A1(n5561), .A2(n5560), .ZN(n5562) );
  INV_X1 U5376 ( .A(n7822), .ZN(n4638) );
  INV_X1 U5377 ( .A(n7821), .ZN(n4637) );
  AND2_X1 U5378 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5713) );
  INV_X1 U5379 ( .A(n7951), .ZN(n4633) );
  INV_X1 U5380 ( .A(n4635), .ZN(n4634) );
  AOI21_X1 U5381 ( .B1(n4647), .B2(n4650), .A(n4310), .ZN(n4646) );
  NOR2_X1 U5382 ( .A1(n6760), .A2(n4288), .ZN(n4647) );
  NAND2_X1 U5383 ( .A1(n4650), .A2(n4649), .ZN(n4648) );
  INV_X1 U5384 ( .A(n6760), .ZN(n4649) );
  NAND2_X1 U5385 ( .A1(n6593), .A2(n4655), .ZN(n4654) );
  INV_X1 U5386 ( .A(n6594), .ZN(n4655) );
  NAND2_X1 U5387 ( .A1(n4659), .A2(n4658), .ZN(n4662) );
  NOR4_X1 U5388 ( .A1(n7425), .A2(n7424), .A3(n7448), .A4(n7423), .ZN(n7426)
         );
  AND2_X1 U5389 ( .A1(n4555), .A2(n4553), .ZN(n7254) );
  OR2_X1 U5390 ( .A1(n5226), .A2(n5225), .ZN(n4667) );
  NAND2_X1 U5391 ( .A1(n4667), .A2(n4666), .ZN(n4665) );
  NAND2_X1 U5392 ( .A1(n5942), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4666) );
  OR2_X1 U5393 ( .A1(n8044), .A2(n4345), .ZN(n4669) );
  NOR2_X1 U5394 ( .A1(n7444), .A2(n8287), .ZN(n8079) );
  NAND2_X1 U5395 ( .A1(n4560), .A2(n4564), .ZN(n7192) );
  INV_X1 U5396 ( .A(n4565), .ZN(n4564) );
  INV_X1 U5397 ( .A(n7441), .ZN(n7422) );
  NAND2_X1 U5398 ( .A1(n4795), .A2(n4793), .ZN(n7442) );
  NOR2_X1 U5399 ( .A1(n8296), .A2(n8107), .ZN(n4794) );
  NOR2_X1 U5400 ( .A1(n8098), .A2(n8296), .ZN(n8086) );
  NAND2_X1 U5401 ( .A1(n7175), .A2(n8160), .ZN(n4427) );
  NOR2_X1 U5402 ( .A1(n4425), .A2(n8157), .ZN(n8113) );
  OR2_X1 U5403 ( .A1(n4290), .A2(n8306), .ZN(n4425) );
  INV_X1 U5404 ( .A(n8126), .ZN(n8127) );
  NAND2_X1 U5405 ( .A1(n8142), .A2(n7189), .ZN(n8128) );
  NOR2_X1 U5406 ( .A1(n4426), .A2(n8157), .ZN(n8148) );
  OR2_X1 U5407 ( .A1(n8317), .A2(n8322), .ZN(n4426) );
  OR2_X1 U5408 ( .A1(n8322), .A2(n7892), .ZN(n7348) );
  NAND2_X1 U5409 ( .A1(n7348), .A2(n7360), .ZN(n8163) );
  CLKBUF_X1 U5410 ( .A(n8161), .Z(n8180) );
  NAND2_X1 U5411 ( .A1(n8234), .A2(n4442), .ZN(n8189) );
  NOR2_X1 U5412 ( .A1(n8332), .A2(n4443), .ZN(n4442) );
  INV_X1 U5413 ( .A(n4444), .ZN(n4443) );
  AND2_X1 U5414 ( .A1(n7350), .A2(n8196), .ZN(n8207) );
  OR2_X1 U5415 ( .A1(n7071), .A2(n9830), .ZN(n7095) );
  NAND2_X1 U5416 ( .A1(n8234), .A2(n4446), .ZN(n8220) );
  NAND2_X1 U5417 ( .A1(n4778), .A2(n4777), .ZN(n8219) );
  AOI21_X1 U5418 ( .B1(n4779), .B2(n4783), .A(n4274), .ZN(n4777) );
  NAND2_X1 U5419 ( .A1(n8234), .A2(n4787), .ZN(n8235) );
  NAND2_X1 U5420 ( .A1(n7181), .A2(n7333), .ZN(n9323) );
  AND2_X1 U5421 ( .A1(n7334), .A2(n7329), .ZN(n4576) );
  NAND2_X1 U5422 ( .A1(n4786), .A2(n4784), .ZN(n9324) );
  AND2_X1 U5423 ( .A1(n4786), .A2(n4788), .ZN(n9326) );
  NAND2_X1 U5424 ( .A1(n7057), .A2(n7416), .ZN(n4786) );
  OR2_X1 U5425 ( .A1(n9356), .A2(n9352), .ZN(n9357) );
  NOR2_X1 U5426 ( .A1(n9357), .A2(n7976), .ZN(n9335) );
  NAND2_X1 U5427 ( .A1(n6603), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6904) );
  AND2_X1 U5428 ( .A1(n7318), .A2(n7321), .ZN(n9593) );
  NOR2_X1 U5429 ( .A1(n4569), .A2(n4568), .ZN(n4567) );
  INV_X1 U5430 ( .A(n7265), .ZN(n4568) );
  INV_X1 U5431 ( .A(n7317), .ZN(n4569) );
  AND2_X1 U5432 ( .A1(n9598), .A2(n9720), .ZN(n9596) );
  NOR2_X1 U5433 ( .A1(n6294), .A2(n9703), .ZN(n6474) );
  AND2_X1 U5434 ( .A1(n6474), .A2(n9712), .ZN(n9598) );
  INV_X1 U5435 ( .A(n5976), .ZN(n5975) );
  AND2_X1 U5436 ( .A1(n7299), .A2(n7265), .ZN(n7399) );
  INV_X1 U5437 ( .A(n7990), .ZN(n6519) );
  NAND3_X1 U5438 ( .A1(n9609), .A2(n4448), .A3(n4271), .ZN(n6294) );
  NAND2_X1 U5439 ( .A1(n9609), .A2(n4278), .ZN(n6265) );
  NAND2_X1 U5440 ( .A1(n9609), .A2(n4271), .ZN(n6266) );
  OAI211_X1 U5441 ( .C1(n6121), .C2(n4557), .A(n4556), .B(n7305), .ZN(n6262)
         );
  INV_X1 U5442 ( .A(n4558), .ZN(n4557) );
  NOR2_X1 U5443 ( .A1(n5973), .A2(n4559), .ZN(n4558) );
  OR2_X1 U5444 ( .A1(n6306), .A2(n9552), .ZN(n9605) );
  NOR2_X1 U5445 ( .A1(n9605), .A2(n9610), .ZN(n9609) );
  NAND2_X1 U5446 ( .A1(n6183), .A2(n7284), .ZN(n7400) );
  XNOR2_X1 U5447 ( .A(n5963), .B(n5961), .ZN(n5962) );
  AND2_X1 U5448 ( .A1(n9639), .A2(n7435), .ZN(n9694) );
  INV_X1 U5449 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n9895) );
  AND2_X1 U5450 ( .A1(n4839), .A2(n4775), .ZN(n4581) );
  AND2_X1 U5451 ( .A1(n4330), .A2(n5066), .ZN(n4775) );
  OR2_X1 U5452 ( .A1(n5004), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5024) );
  OR2_X1 U5453 ( .A1(n6543), .A2(n6416), .ZN(n6413) );
  NAND2_X1 U5454 ( .A1(n6433), .A2(n6432), .ZN(n6530) );
  AND2_X1 U5455 ( .A1(n7620), .A2(n7621), .ZN(n8416) );
  AOI21_X1 U5456 ( .B1(n4371), .B2(n4372), .A(n4370), .ZN(n4369) );
  INV_X1 U5457 ( .A(n8508), .ZN(n4370) );
  AND2_X1 U5458 ( .A1(n7545), .A2(n7543), .ZN(n8442) );
  INV_X1 U5459 ( .A(n6941), .ZN(n6940) );
  NAND2_X1 U5460 ( .A1(n6532), .A2(n6533), .ZN(n6563) );
  OR2_X1 U5461 ( .A1(n6339), .A2(n6336), .ZN(n6370) );
  NAND2_X1 U5462 ( .A1(n6703), .A2(n8823), .ZN(n4484) );
  NAND2_X1 U5463 ( .A1(n4591), .A2(n7584), .ZN(n8406) );
  INV_X1 U5464 ( .A(n8405), .ZN(n4591) );
  NAND2_X1 U5465 ( .A1(n6741), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6806) );
  INV_X1 U5466 ( .A(n6743), .ZN(n6741) );
  NAND2_X1 U5467 ( .A1(n7464), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n7629) );
  INV_X1 U5468 ( .A(n7608), .ZN(n7464) );
  NAND2_X1 U5469 ( .A1(n6572), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6623) );
  INV_X1 U5470 ( .A(n6029), .ZN(n6027) );
  NAND2_X1 U5471 ( .A1(n5985), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6029) );
  INV_X1 U5472 ( .A(n5987), .ZN(n5985) );
  OR2_X1 U5473 ( .A1(n6806), .A2(n6805), .ZN(n6821) );
  OR2_X1 U5474 ( .A1(n6821), .A2(n8509), .ZN(n6941) );
  OAI21_X1 U5475 ( .B1(n8627), .B2(n8634), .A(n8790), .ZN(n4723) );
  NOR2_X1 U5476 ( .A1(n8607), .A2(n4392), .ZN(n4391) );
  NAND2_X1 U5477 ( .A1(n8804), .A2(n8628), .ZN(n4393) );
  AND2_X1 U5478 ( .A1(n8889), .A2(n8620), .ZN(n8717) );
  INV_X1 U5479 ( .A(n8717), .ZN(n8791) );
  INV_X1 U5480 ( .A(n5786), .ZN(n7635) );
  NAND2_X1 U5481 ( .A1(n5333), .A2(n5128), .ZN(n5613) );
  INV_X1 U5482 ( .A(n5129), .ZN(n5612) );
  NAND2_X1 U5483 ( .A1(n4359), .A2(n4358), .ZN(n5130) );
  NAND2_X1 U5484 ( .A1(n5994), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n4358) );
  NOR2_X1 U5485 ( .A1(n5130), .A2(n5131), .ZN(n5172) );
  NOR2_X1 U5486 ( .A1(n5848), .A2(n4336), .ZN(n8825) );
  NAND2_X1 U5487 ( .A1(n8825), .A2(n8826), .ZN(n8824) );
  NOR2_X1 U5488 ( .A1(n6241), .A2(n4544), .ZN(n6244) );
  AND2_X1 U5489 ( .A1(n6730), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4544) );
  NOR2_X1 U5490 ( .A1(n6244), .A2(n6243), .ZN(n6853) );
  NAND2_X1 U5491 ( .A1(n6237), .A2(n4351), .ZN(n6238) );
  OR2_X1 U5492 ( .A1(n6730), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n4351) );
  NAND2_X1 U5493 ( .A1(n6238), .A2(n6239), .ZN(n6860) );
  XNOR2_X1 U5494 ( .A(n6854), .B(n9412), .ZN(n9416) );
  AND2_X1 U5495 ( .A1(n4537), .A2(n4536), .ZN(n8847) );
  NAND2_X1 U5496 ( .A1(n8844), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4536) );
  NOR2_X1 U5497 ( .A1(n8847), .A2(n8846), .ZN(n8858) );
  INV_X1 U5498 ( .A(n4412), .ZN(n4410) );
  NAND2_X1 U5499 ( .A1(n4323), .A2(n4414), .ZN(n4413) );
  INV_X1 U5500 ( .A(n8572), .ZN(n4415) );
  NAND2_X1 U5501 ( .A1(n8976), .A2(n8572), .ZN(n8907) );
  AND2_X1 U5502 ( .A1(n7710), .A2(n7684), .ZN(n8498) );
  NAND2_X1 U5503 ( .A1(n8990), .A2(n4754), .ZN(n8967) );
  AND2_X1 U5504 ( .A1(n8990), .A2(n4752), .ZN(n8943) );
  NAND2_X1 U5505 ( .A1(n8977), .A2(n8978), .ZN(n8976) );
  OR2_X1 U5506 ( .A1(n7631), .A2(n7479), .ZN(n7646) );
  AND2_X1 U5507 ( .A1(n9019), .A2(n9010), .ZN(n9005) );
  NAND2_X1 U5508 ( .A1(n7463), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n7569) );
  INV_X1 U5509 ( .A(n7549), .ZN(n7463) );
  OR2_X1 U5510 ( .A1(n7569), .A2(n8409), .ZN(n7589) );
  AOI21_X1 U5511 ( .B1(n9075), .B2(n4490), .A(n4309), .ZN(n4489) );
  NAND2_X1 U5512 ( .A1(n4493), .A2(n4492), .ZN(n9076) );
  NAND2_X1 U5513 ( .A1(n9103), .A2(n4494), .ZN(n4493) );
  NOR2_X1 U5514 ( .A1(n9105), .A2(n4748), .ZN(n9087) );
  INV_X1 U5515 ( .A(n4750), .ZN(n4748) );
  NAND2_X1 U5516 ( .A1(n9110), .A2(n9111), .ZN(n9109) );
  NOR2_X1 U5517 ( .A1(n9105), .A2(n9195), .ZN(n9104) );
  NAND2_X1 U5518 ( .A1(n6939), .A2(n8547), .ZN(n7739) );
  OR2_X1 U5519 ( .A1(n6937), .A2(n9199), .ZN(n9105) );
  AND2_X1 U5520 ( .A1(n4512), .A2(n4518), .ZN(n4511) );
  AOI21_X1 U5521 ( .B1(n4520), .B2(n4519), .A(n4320), .ZN(n4518) );
  AND2_X1 U5522 ( .A1(n9235), .A2(n4735), .ZN(n6848) );
  NOR2_X1 U5523 ( .A1(n4737), .A2(n9210), .ZN(n4735) );
  AND2_X1 U5524 ( .A1(n8546), .A2(n8679), .ZN(n8541) );
  NAND2_X1 U5525 ( .A1(n9235), .A2(n4739), .ZN(n6752) );
  NAND2_X1 U5526 ( .A1(n9235), .A2(n9312), .ZN(n9236) );
  INV_X1 U5527 ( .A(n8749), .ZN(n9231) );
  NOR2_X1 U5528 ( .A1(n6489), .A2(n6636), .ZN(n9235) );
  OAI211_X1 U5529 ( .C1(n6347), .C2(n6334), .A(n6333), .B(n6332), .ZN(n6493)
         );
  NOR2_X1 U5530 ( .A1(n4743), .A2(n4742), .ZN(n4741) );
  NAND2_X1 U5531 ( .A1(n9511), .A2(n9488), .ZN(n4743) );
  NAND2_X1 U5532 ( .A1(n6144), .A2(n6143), .ZN(n6150) );
  NAND2_X1 U5533 ( .A1(n4744), .A2(n4285), .ZN(n6389) );
  NOR2_X1 U5534 ( .A1(n6062), .A2(n4745), .ZN(n6168) );
  NAND2_X1 U5535 ( .A1(n6067), .A2(n9488), .ZN(n4745) );
  NOR2_X1 U5536 ( .A1(n6062), .A2(n6209), .ZN(n6205) );
  NAND2_X1 U5537 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5987) );
  NAND2_X1 U5538 ( .A1(n4483), .A2(n5876), .ZN(n6078) );
  AND2_X1 U5539 ( .A1(n8650), .A2(n9427), .ZN(n6103) );
  INV_X1 U5540 ( .A(n5667), .ZN(n4398) );
  INV_X1 U5541 ( .A(n9114), .ZN(n9062) );
  OR2_X1 U5542 ( .A1(n8950), .A2(n8926), .ZN(n8928) );
  INV_X1 U5543 ( .A(n4523), .ZN(n6799) );
  AND3_X1 U5544 ( .A1(n9468), .A2(n5447), .A3(n5446), .ZN(n5891) );
  INV_X1 U5545 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4529) );
  XNOR2_X1 U5546 ( .A(n7231), .B(n7234), .ZN(n8521) );
  XNOR2_X1 U5547 ( .A(n7001), .B(n7000), .ZN(n7460) );
  NAND2_X1 U5548 ( .A1(n4713), .A2(n4716), .ZN(n7001) );
  OR2_X1 U5549 ( .A1(n6834), .A2(n4719), .ZN(n4713) );
  OR2_X1 U5550 ( .A1(n6834), .A2(n6833), .ZN(n4720) );
  INV_X1 U5551 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4886) );
  NOR2_X1 U5552 ( .A1(n4618), .A2(n4862), .ZN(n4617) );
  INV_X1 U5553 ( .A(n4619), .ZN(n4618) );
  NAND2_X1 U5554 ( .A1(n4705), .A2(n5297), .ZN(n5432) );
  NAND2_X1 U5555 ( .A1(n5115), .A2(n4710), .ZN(n4705) );
  NAND2_X1 U5556 ( .A1(n5115), .A2(n5114), .ZN(n5299) );
  NAND2_X1 U5557 ( .A1(n4694), .A2(n4695), .ZN(n5034) );
  OR2_X1 U5558 ( .A1(n4998), .A2(n5017), .ZN(n4694) );
  XNOR2_X1 U5559 ( .A(n4960), .B(SI_7_), .ZN(n4966) );
  INV_X1 U5560 ( .A(n4679), .ZN(n4678) );
  OAI21_X1 U5561 ( .B1(n4683), .B2(n4922), .A(n4317), .ZN(n4679) );
  XNOR2_X1 U5562 ( .A(n4948), .B(SI_6_), .ZN(n4954) );
  INV_X1 U5563 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n4367) );
  INV_X1 U5564 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4366) );
  INV_X1 U5565 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4365) );
  NAND2_X1 U5566 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n4542) );
  INV_X1 U5567 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4899) );
  NAND2_X1 U5568 ( .A1(n4662), .A2(n4660), .ZN(n7789) );
  INV_X1 U5569 ( .A(n8119), .ZN(n7901) );
  INV_X1 U5570 ( .A(n7988), .ZN(n6611) );
  NAND2_X1 U5571 ( .A1(n4636), .A2(n4635), .ZN(n7862) );
  AND2_X1 U5572 ( .A1(n4636), .A2(n4295), .ZN(n7864) );
  NAND2_X1 U5573 ( .A1(n7952), .A2(n7951), .ZN(n4636) );
  AND2_X1 U5574 ( .A1(n7874), .A2(n7873), .ZN(n7875) );
  NAND2_X1 U5575 ( .A1(n7165), .A2(n7164), .ZN(n8290) );
  AOI21_X1 U5576 ( .B1(n5803), .B2(n4660), .A(n6047), .ZN(n4657) );
  NAND2_X1 U5577 ( .A1(n5669), .A2(n4438), .ZN(n4440) );
  OAI21_X1 U5578 ( .B1(n5551), .B2(n7244), .A(n4439), .ZN(n4438) );
  NAND2_X1 U5579 ( .A1(n7104), .A2(n7103), .ZN(n8327) );
  INV_X1 U5580 ( .A(n4644), .ZN(n6761) );
  AOI21_X1 U5581 ( .B1(n6596), .B2(n4288), .A(n4645), .ZN(n4644) );
  INV_X1 U5582 ( .A(n4650), .ZN(n4645) );
  XNOR2_X1 U5583 ( .A(n7842), .B(n7840), .ZN(n7899) );
  AOI21_X1 U5584 ( .B1(n9551), .B2(n9548), .A(n9547), .ZN(n5801) );
  AND3_X1 U5585 ( .A1(n7130), .A2(n7129), .A3(n7128), .ZN(n8166) );
  NOR2_X1 U5586 ( .A1(n5571), .A2(n7435), .ZN(n9559) );
  NAND2_X1 U5587 ( .A1(n4632), .A2(n4631), .ZN(n7934) );
  OR2_X1 U5588 ( .A1(n7952), .A2(n4634), .ZN(n4631) );
  OAI21_X1 U5589 ( .B1(n6596), .B2(n4648), .A(n4646), .ZN(n6898) );
  OAI21_X1 U5590 ( .B1(n6596), .B2(n6595), .A(n4654), .ZN(n6651) );
  OR2_X1 U5591 ( .A1(n6455), .A2(n9794), .ZN(n5559) );
  OR2_X1 U5592 ( .A1(n5696), .A2(n5554), .ZN(n5558) );
  INV_X1 U5593 ( .A(n4662), .ZN(n6042) );
  NAND2_X1 U5594 ( .A1(n4623), .A2(n7843), .ZN(n7959) );
  NAND2_X1 U5595 ( .A1(n7898), .A2(n7899), .ZN(n4623) );
  OR2_X1 U5596 ( .A1(n5571), .A2(n5570), .ZN(n7978) );
  NAND4_X1 U5597 ( .A1(n5717), .A2(n5716), .A3(n5715), .A4(n5714), .ZN(n7993)
         );
  NAND4_X1 U5598 ( .A1(n5707), .A2(n5706), .A3(n5705), .A4(n5704), .ZN(n9623)
         );
  OR2_X1 U5599 ( .A1(n5577), .A2(n5683), .ZN(n5687) );
  OR2_X1 U5600 ( .A1(n5577), .A2(n5088), .ZN(n5090) );
  NAND2_X1 U5601 ( .A1(n5276), .A2(n5277), .ZN(n5275) );
  NOR2_X1 U5602 ( .A1(n5239), .A2(n5238), .ZN(n5237) );
  AND2_X1 U5603 ( .A1(n5275), .A2(n4677), .ZN(n5239) );
  NAND2_X1 U5604 ( .A1(n5796), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4677) );
  INV_X1 U5605 ( .A(n4667), .ZN(n5326) );
  AND2_X1 U5606 ( .A1(n4665), .A2(n4664), .ZN(n5596) );
  INV_X1 U5607 ( .A(n5328), .ZN(n4664) );
  INV_X1 U5608 ( .A(n4665), .ZN(n5329) );
  NOR2_X1 U5609 ( .A1(n5596), .A2(n4663), .ZN(n5599) );
  AND2_X1 U5610 ( .A1(n5908), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4663) );
  NOR2_X1 U5611 ( .A1(n5901), .A2(n4672), .ZN(n5904) );
  AND2_X1 U5612 ( .A1(n6600), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4672) );
  NAND2_X1 U5613 ( .A1(n5904), .A2(n5903), .ZN(n6227) );
  NAND2_X1 U5614 ( .A1(n6227), .A2(n4671), .ZN(n6231) );
  OR2_X1 U5615 ( .A1(n6762), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4671) );
  NAND2_X1 U5616 ( .A1(n6231), .A2(n6230), .ZN(n7996) );
  NOR2_X1 U5617 ( .A1(n8033), .A2(n4670), .ZN(n8037) );
  AND2_X1 U5618 ( .A1(n8034), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4670) );
  NOR2_X1 U5619 ( .A1(n8037), .A2(n8036), .ZN(n8044) );
  XNOR2_X1 U5620 ( .A(n4669), .B(n4668), .ZN(n8045) );
  INV_X1 U5621 ( .A(n8272), .ZN(n8075) );
  AND2_X1 U5622 ( .A1(n7221), .A2(n7220), .ZN(n8285) );
  NAND2_X1 U5623 ( .A1(n7451), .A2(n9619), .ZN(n7456) );
  INV_X1 U5624 ( .A(n4563), .ZN(n8090) );
  AOI21_X1 U5625 ( .B1(n8105), .B2(n4803), .A(n4566), .ZN(n4563) );
  OAI21_X1 U5626 ( .B1(n8124), .B2(n4276), .A(n4798), .ZN(n8085) );
  INV_X1 U5627 ( .A(n8301), .ZN(n8104) );
  NAND2_X1 U5628 ( .A1(n4801), .A2(n4804), .ZN(n8097) );
  NAND2_X1 U5629 ( .A1(n8124), .A2(n4806), .ZN(n4801) );
  NOR2_X1 U5630 ( .A1(n8124), .A2(n4809), .ZN(n8112) );
  NAND2_X1 U5631 ( .A1(n7053), .A2(n7052), .ZN(n8310) );
  NAND2_X1 U5632 ( .A1(n4767), .A2(n4765), .ZN(n8173) );
  NAND2_X1 U5633 ( .A1(n7090), .A2(n4768), .ZN(n4767) );
  NAND2_X1 U5634 ( .A1(n7090), .A2(n4811), .ZN(n8188) );
  NAND2_X1 U5635 ( .A1(n4575), .A2(n4574), .ZN(n8227) );
  NAND2_X1 U5636 ( .A1(n4781), .A2(n4782), .ZN(n8233) );
  OR2_X1 U5637 ( .A1(n7057), .A2(n4783), .ZN(n4781) );
  NAND2_X1 U5638 ( .A1(n7055), .A2(n7054), .ZN(n9332) );
  NAND2_X1 U5639 ( .A1(n9341), .A2(n7329), .ZN(n7180) );
  AND2_X1 U5640 ( .A1(n4792), .A2(n4791), .ZN(n9355) );
  NAND2_X1 U5641 ( .A1(n9594), .A2(n6780), .ZN(n6782) );
  NAND2_X1 U5642 ( .A1(n6602), .A2(n6601), .ZN(n9592) );
  NAND2_X1 U5643 ( .A1(n4772), .A2(n5955), .ZN(n5957) );
  NAND2_X1 U5644 ( .A1(n6120), .A2(n7293), .ZN(n6111) );
  OR2_X1 U5645 ( .A1(n9631), .A2(n8275), .ZN(n8238) );
  INV_X1 U5646 ( .A(n8237), .ZN(n9591) );
  INV_X1 U5647 ( .A(n8078), .ZN(n9337) );
  INV_X1 U5648 ( .A(n9632), .ZN(n9887) );
  XNOR2_X1 U5649 ( .A(n4833), .B(n4835), .ZN(n6589) );
  XNOR2_X1 U5650 ( .A(n5061), .B(n4474), .ZN(n7253) );
  INV_X1 U5651 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5679) );
  NAND2_X1 U5652 ( .A1(n4608), .A2(n7488), .ZN(n8389) );
  NAND2_X1 U5653 ( .A1(n7759), .A2(n7758), .ZN(n9131) );
  INV_X1 U5654 ( .A(n5472), .ZN(n5474) );
  INV_X1 U5655 ( .A(n4588), .ZN(n4587) );
  OAI21_X1 U5656 ( .B1(n8461), .B2(n4589), .A(n8462), .ZN(n4588) );
  INV_X1 U5657 ( .A(n6878), .ZN(n6880) );
  NAND2_X1 U5658 ( .A1(n8453), .A2(n7659), .ZN(n4603) );
  NAND2_X1 U5659 ( .A1(n7663), .A2(n7662), .ZN(n9148) );
  NAND2_X1 U5660 ( .A1(n7661), .A2(n7642), .ZN(n7663) );
  INV_X1 U5661 ( .A(n9113), .ZN(n8436) );
  INV_X1 U5662 ( .A(n9096), .ZN(n9059) );
  NAND2_X1 U5663 ( .A1(n8396), .A2(n8397), .ZN(n4604) );
  INV_X1 U5664 ( .A(n8814), .ZN(n6709) );
  NAND2_X1 U5665 ( .A1(n5463), .A2(n9276), .ZN(n5418) );
  NAND2_X1 U5666 ( .A1(n6956), .A2(n6955), .ZN(n7490) );
  NOR2_X1 U5667 ( .A1(n6707), .A2(n4593), .ZN(n4592) );
  INV_X1 U5668 ( .A(n6701), .ZN(n4593) );
  OR2_X1 U5669 ( .A1(n8511), .A2(n9062), .ZN(n8487) );
  NAND2_X1 U5670 ( .A1(n7548), .A2(n7547), .ZN(n9184) );
  OR2_X1 U5671 ( .A1(n8511), .A2(n9060), .ZN(n8500) );
  OAI21_X1 U5672 ( .B1(n4608), .B2(n4372), .A(n4371), .ZN(n8506) );
  INV_X1 U5673 ( .A(n8485), .ZN(n8517) );
  INV_X1 U5674 ( .A(n8719), .ZN(n8722) );
  NAND2_X1 U5675 ( .A1(n5496), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5790) );
  AND3_X1 U5676 ( .A1(n5656), .A2(n5655), .A3(n5654), .ZN(n5657) );
  NAND2_X1 U5677 ( .A1(n5496), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5480) );
  NAND2_X1 U5678 ( .A1(n5496), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5408) );
  INV_X1 U5679 ( .A(n4359), .ZN(n5163) );
  NAND2_X1 U5680 ( .A1(n5609), .A2(n4533), .ZN(n5161) );
  NAND2_X1 U5681 ( .A1(n4535), .A2(n4534), .ZN(n4533) );
  INV_X1 U5682 ( .A(n7202), .ZN(n4535) );
  NAND2_X1 U5683 ( .A1(n6145), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4531) );
  NOR2_X1 U5684 ( .A1(n5282), .A2(n5283), .ZN(n5345) );
  NAND2_X1 U5685 ( .A1(n4355), .A2(n4354), .ZN(n5346) );
  OR2_X1 U5686 ( .A1(n6331), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n4354) );
  INV_X1 U5687 ( .A(n5345), .ZN(n4355) );
  NAND2_X1 U5688 ( .A1(n5346), .A2(n5347), .ZN(n5511) );
  NAND2_X1 U5689 ( .A1(n5842), .A2(n5843), .ZN(n6237) );
  NAND2_X1 U5690 ( .A1(n8829), .A2(n4352), .ZN(n5842) );
  OR2_X1 U5691 ( .A1(n8828), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n4352) );
  AND2_X1 U5692 ( .A1(n5109), .A2(n5157), .ZN(n6861) );
  NOR2_X1 U5693 ( .A1(n7008), .A2(n7009), .ZN(n7012) );
  INV_X1 U5694 ( .A(n4537), .ZN(n8843) );
  NOR2_X1 U5695 ( .A1(n7015), .A2(n7016), .ZN(n7020) );
  INV_X1 U5696 ( .A(n4350), .ZN(n8853) );
  NAND2_X1 U5697 ( .A1(n8857), .A2(n8856), .ZN(n8873) );
  AND2_X1 U5698 ( .A1(n4350), .A2(n4349), .ZN(n8857) );
  NAND2_X1 U5699 ( .A1(n8859), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n4349) );
  INV_X1 U5700 ( .A(n9122), .ZN(n8889) );
  AND2_X1 U5701 ( .A1(n8925), .A2(n8924), .ZN(n9130) );
  NAND2_X1 U5702 ( .A1(n8901), .A2(n8900), .ZN(n8923) );
  INV_X1 U5703 ( .A(n9136), .ZN(n8949) );
  NAND2_X1 U5704 ( .A1(n4498), .A2(n4503), .ZN(n8898) );
  OR2_X1 U5705 ( .A1(n8989), .A2(n4504), .ZN(n4498) );
  AND2_X1 U5706 ( .A1(n7683), .A2(n7666), .ZN(n8969) );
  INV_X1 U5707 ( .A(n9148), .ZN(n8972) );
  NAND2_X1 U5708 ( .A1(n4508), .A2(n4507), .ZN(n8959) );
  AND2_X1 U5709 ( .A1(n4508), .A2(n4509), .ZN(n8975) );
  NAND2_X1 U5710 ( .A1(n4401), .A2(n4404), .ZN(n8996) );
  AND2_X1 U5711 ( .A1(n7478), .A2(n7477), .ZN(n8994) );
  NAND2_X1 U5712 ( .A1(n4403), .A2(n8693), .ZN(n9011) );
  NAND2_X1 U5713 ( .A1(n9021), .A2(n8759), .ZN(n4403) );
  INV_X1 U5714 ( .A(n9161), .ZN(n9010) );
  NAND2_X1 U5715 ( .A1(n7606), .A2(n7605), .ZN(n9168) );
  NAND2_X1 U5716 ( .A1(n7588), .A2(n7587), .ZN(n9174) );
  AND2_X1 U5717 ( .A1(n7568), .A2(n7567), .ZN(n9068) );
  NAND2_X1 U5718 ( .A1(n9076), .A2(n9075), .ZN(n9182) );
  AND2_X1 U5719 ( .A1(n4495), .A2(n4497), .ZN(n9086) );
  NAND2_X1 U5720 ( .A1(n9103), .A2(n9102), .ZN(n4495) );
  AND2_X1 U5721 ( .A1(n6619), .A2(n6618), .ZN(n6734) );
  AND2_X1 U5722 ( .A1(n6350), .A2(n6349), .ZN(n6629) );
  INV_X1 U5723 ( .A(n9429), .ZN(n9100) );
  INV_X1 U5724 ( .A(n9428), .ZN(n9031) );
  AOI211_X1 U5725 ( .C1(n9216), .C2(n9396), .A(n9395), .B(n9394), .ZN(n9407)
         );
  NAND2_X1 U5726 ( .A1(n4417), .A2(n4340), .ZN(n4416) );
  NOR2_X1 U5727 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n4530) );
  NAND2_X1 U5728 ( .A1(n4878), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4874) );
  OR2_X1 U5729 ( .A1(n4876), .A2(n4875), .ZN(n4877) );
  XNOR2_X1 U5730 ( .A(n6587), .B(n6586), .ZN(n7476) );
  NAND2_X1 U5731 ( .A1(n4731), .A2(n6498), .ZN(n6587) );
  OR2_X1 U5732 ( .A1(n6500), .A2(n6499), .ZN(n4731) );
  INV_X1 U5733 ( .A(n8794), .ZN(n8773) );
  AND2_X1 U5734 ( .A1(n4854), .A2(n4293), .ZN(n5007) );
  INV_X1 U5735 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9891) );
  INV_X1 U5736 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6334) );
  INV_X1 U5737 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n4991) );
  NAND2_X1 U5738 ( .A1(n4682), .A2(n4922), .ZN(n4944) );
  NAND2_X1 U5739 ( .A1(n4937), .A2(n4936), .ZN(n4682) );
  OR2_X1 U5740 ( .A1(n4941), .A2(n5306), .ZN(n4958) );
  NAND2_X1 U5741 ( .A1(n4942), .A2(n4540), .ZN(n5124) );
  INV_X1 U5742 ( .A(n4941), .ZN(n4942) );
  INV_X1 U5743 ( .A(n4541), .ZN(n4540) );
  OAI22_X1 U5744 ( .A1(n5420), .A2(n4542), .B1(P1_IR_REG_31__SCAN_IN), .B2(
        P1_IR_REG_1__SCAN_IN), .ZN(n4541) );
  INV_X1 U5745 ( .A(n4454), .ZN(n7439) );
  OAI211_X1 U5746 ( .C1(n8069), .C2(n5547), .A(n4674), .B(n4344), .ZN(P2_U3264) );
  NAND2_X1 U5747 ( .A1(n4675), .A2(n5547), .ZN(n4674) );
  NAND2_X1 U5748 ( .A1(n4431), .A2(n4342), .ZN(P2_U3517) );
  NAND2_X1 U5749 ( .A1(n8357), .A2(n9726), .ZN(n4431) );
  INV_X1 U5750 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n4430) );
  OAI222_X1 U5751 ( .A1(n8371), .A2(n7219), .B1(n4268), .B2(n9270), .C1(
        P2_U3152), .C2(n7040), .ZN(P2_U3328) );
  OAI222_X1 U5752 ( .A1(n8371), .A2(n7131), .B1(n4268), .B2(n6727), .C1(n6725), 
        .C2(P2_U3152), .ZN(P2_U3333) );
  OAI21_X1 U5753 ( .B1(n7033), .B2(n4268), .A(n4480), .ZN(P2_U3336) );
  INV_X1 U5754 ( .A(n4481), .ZN(n4480) );
  OAI222_X1 U5755 ( .A1(n8371), .A2(n5829), .B1(n4268), .B2(n5830), .C1(
        P2_U3152), .C2(n8213), .ZN(P2_U3339) );
  OAI222_X1 U5756 ( .A1(n8371), .A2(n5767), .B1(n4268), .B2(n5766), .C1(
        P2_U3152), .C2(n4668), .ZN(P2_U3340) );
  OAI222_X1 U5757 ( .A1(n8371), .A2(n6975), .B1(n4268), .B2(n5317), .C1(
        P2_U3152), .C2(n8019), .ZN(P2_U3343) );
  OAI222_X1 U5758 ( .A1(n8371), .A2(n5057), .B1(n4268), .B2(n5056), .C1(
        P2_U3152), .C2(n5860), .ZN(P2_U3346) );
  OAI222_X1 U5759 ( .A1(n8371), .A2(n5553), .B1(n4268), .B2(n5551), .C1(
        P2_U3152), .C2(n5552), .ZN(P2_U3357) );
  NOR2_X1 U5760 ( .A1(n7788), .A2(n4583), .ZN(n7721) );
  OAI211_X1 U5761 ( .C1(n8880), .C2(n8917), .A(n4547), .B(n4545), .ZN(P1_U3260) );
  INV_X1 U5762 ( .A(n4546), .ZN(n4545) );
  NAND2_X1 U5763 ( .A1(n4360), .A2(n8917), .ZN(n4547) );
  OR2_X1 U5764 ( .A1(n4389), .A2(n4284), .ZN(n4270) );
  AND2_X1 U5765 ( .A1(n4278), .A2(n4449), .ZN(n4271) );
  OR2_X1 U5766 ( .A1(n7735), .A2(n8963), .ZN(n4272) );
  AND2_X1 U5767 ( .A1(n4389), .A2(n4284), .ZN(n4273) );
  AND2_X1 U5768 ( .A1(n4787), .A2(n7954), .ZN(n4274) );
  INV_X1 U5769 ( .A(n5785), .ZN(n5989) );
  NAND2_X2 U5770 ( .A1(n5463), .A2(n5461), .ZN(n6347) );
  NAND3_X1 U5771 ( .A1(n4755), .A2(n4756), .A3(n4529), .ZN(n4275) );
  OR2_X1 U5772 ( .A1(n4805), .A2(n4800), .ZN(n4276) );
  NOR2_X1 U5773 ( .A1(n8177), .A2(n8165), .ZN(n4277) );
  NOR2_X1 U5774 ( .A1(n7976), .A2(n7984), .ZN(n7056) );
  AND2_X1 U5775 ( .A1(n9682), .A2(n9676), .ZN(n4278) );
  AOI211_X1 U5776 ( .C1(n8932), .C2(n9128), .A(n9519), .B(n8915), .ZN(n9127)
         );
  INV_X1 U5777 ( .A(n9127), .ZN(n4417) );
  AOI21_X1 U5778 ( .B1(n7586), .B2(n7235), .A(n7092), .ZN(n8194) );
  NAND2_X1 U5779 ( .A1(n4375), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4879) );
  OR2_X1 U5780 ( .A1(n7383), .A2(n7384), .ZN(n4279) );
  INV_X1 U5781 ( .A(n8118), .ZN(n4806) );
  INV_X1 U5782 ( .A(n7488), .ZN(n4613) );
  NOR2_X1 U5783 ( .A1(n7732), .A2(n4301), .ZN(n4507) );
  NAND2_X1 U5784 ( .A1(n6802), .A2(n6801), .ZN(n9210) );
  INV_X1 U5785 ( .A(n5803), .ZN(n4658) );
  AND2_X1 U5786 ( .A1(n9141), .A2(n8952), .ZN(n8905) );
  INV_X1 U5787 ( .A(n8905), .ZN(n4414) );
  OR2_X1 U5788 ( .A1(n8290), .A2(n7849), .ZN(n7383) );
  OR2_X1 U5789 ( .A1(n8285), .A2(n4549), .ZN(n4280) );
  AND2_X1 U5790 ( .A1(n7293), .A2(n7272), .ZN(n4281) );
  INV_X1 U5791 ( .A(n4922), .ZN(n4684) );
  INV_X1 U5792 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4939) );
  AND2_X1 U5793 ( .A1(n7343), .A2(n7263), .ZN(n4282) );
  AND3_X1 U5794 ( .A1(n4441), .A2(n4829), .A3(n4330), .ZN(n4283) );
  AND2_X1 U5795 ( .A1(n9195), .A2(n9095), .ZN(n7725) );
  INV_X1 U5796 ( .A(n8349), .ZN(n4787) );
  NAND2_X1 U5797 ( .A1(n4479), .A2(n7429), .ZN(n7391) );
  AND2_X1 U5798 ( .A1(n7637), .A2(n7636), .ZN(n4284) );
  AND3_X1 U5799 ( .A1(n6067), .A2(n6314), .A3(n9488), .ZN(n4285) );
  NAND2_X1 U5800 ( .A1(n6019), .A2(n6018), .ZN(n4286) );
  XNOR2_X1 U5801 ( .A(n5064), .B(n5063), .ZN(n5185) );
  INV_X1 U5802 ( .A(n6347), .ZN(n7524) );
  NAND2_X2 U5803 ( .A1(n7756), .A2(n7040), .ZN(n5579) );
  NAND2_X1 U5804 ( .A1(n4938), .A2(n4760), .ZN(n4925) );
  NAND2_X1 U5805 ( .A1(n5924), .A2(n5923), .ZN(n7273) );
  NAND2_X1 U5806 ( .A1(n9400), .A2(n8812), .ZN(n4287) );
  NAND2_X1 U5807 ( .A1(n4854), .A2(n4619), .ZN(n5010) );
  NAND2_X1 U5808 ( .A1(n5669), .A2(n5461), .ZN(n5678) );
  AND2_X1 U5809 ( .A1(n4653), .A2(n4654), .ZN(n4288) );
  INV_X1 U5810 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5306) );
  NAND2_X1 U5811 ( .A1(n5672), .A2(n5671), .ZN(n9649) );
  OR2_X1 U5812 ( .A1(n9168), .A2(n9041), .ZN(n8693) );
  INV_X1 U5813 ( .A(n8693), .ZN(n4406) );
  NAND2_X1 U5814 ( .A1(n8332), .A2(n8209), .ZN(n4289) );
  AND3_X1 U5815 ( .A1(n5465), .A2(n5467), .A3(n5466), .ZN(n8650) );
  INV_X1 U5816 ( .A(n8650), .ZN(n9473) );
  INV_X1 U5817 ( .A(n9075), .ZN(n4491) );
  INV_X1 U5818 ( .A(n7497), .ZN(n6957) );
  INV_X1 U5819 ( .A(n8317), .ZN(n4428) );
  NAND2_X1 U5820 ( .A1(n7123), .A2(n7122), .ZN(n8317) );
  OR2_X1 U5821 ( .A1(n8317), .A2(n4427), .ZN(n4290) );
  AND2_X1 U5822 ( .A1(n6044), .A2(n6043), .ZN(n4291) );
  NAND2_X1 U5823 ( .A1(n8406), .A2(n7585), .ZN(n8460) );
  AND2_X1 U5824 ( .A1(n4982), .A2(n4851), .ZN(n4984) );
  AND3_X1 U5825 ( .A1(n8671), .A2(n8669), .A3(n8628), .ZN(n4292) );
  NAND4_X1 U5826 ( .A1(n5481), .A2(n5480), .A3(n5479), .A4(n5478), .ZN(n8822)
         );
  NAND2_X1 U5827 ( .A1(n7115), .A2(n7114), .ZN(n8322) );
  INV_X1 U5828 ( .A(n9325), .ZN(n4785) );
  NOR2_X1 U5829 ( .A1(n4977), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n4982) );
  INV_X1 U5830 ( .A(n7263), .ZN(n4571) );
  AND2_X1 U5831 ( .A1(n4853), .A2(n4620), .ZN(n4293) );
  AND2_X1 U5832 ( .A1(n4264), .A2(n6079), .ZN(n4294) );
  NAND2_X1 U5833 ( .A1(n7816), .A2(n7817), .ZN(n4295) );
  OR2_X1 U5834 ( .A1(n9210), .A2(n8811), .ZN(n4296) );
  AND2_X1 U5835 ( .A1(n9354), .A2(n4791), .ZN(n4297) );
  NAND2_X1 U5836 ( .A1(n7526), .A2(n7525), .ZN(n9189) );
  NAND2_X1 U5837 ( .A1(n4938), .A2(n4939), .ZN(n4923) );
  NAND2_X1 U5838 ( .A1(n4941), .A2(n4734), .ZN(n4978) );
  AND2_X1 U5839 ( .A1(n4532), .A2(n4531), .ZN(n4298) );
  NAND2_X1 U5840 ( .A1(n7059), .A2(n7058), .ZN(n8349) );
  AND2_X1 U5841 ( .A1(n9189), .A2(n9115), .ZN(n4299) );
  OR2_X1 U5842 ( .A1(n4410), .A2(n4413), .ZN(n4300) );
  NOR2_X1 U5843 ( .A1(n7747), .A2(n8399), .ZN(n4301) );
  AND2_X1 U5844 ( .A1(n8168), .A2(n7348), .ZN(n4302) );
  OR2_X1 U5845 ( .A1(n8626), .A2(n8628), .ZN(n4303) );
  AND2_X1 U5846 ( .A1(n6567), .A2(n6566), .ZN(n9312) );
  AND3_X1 U5847 ( .A1(n7389), .A2(n7387), .A3(n7388), .ZN(n4304) );
  INV_X1 U5848 ( .A(n4805), .ZN(n4804) );
  OAI21_X1 U5849 ( .B1(n8118), .B2(n4810), .A(n4808), .ZN(n4805) );
  AND2_X1 U5850 ( .A1(n8906), .A2(n8978), .ZN(n4305) );
  AND2_X1 U5851 ( .A1(n4723), .A2(n4267), .ZN(n4306) );
  NOR2_X1 U5852 ( .A1(n5561), .A2(n5560), .ZN(n5664) );
  AND2_X1 U5853 ( .A1(n8728), .A2(n8909), .ZN(n8922) );
  AND2_X1 U5854 ( .A1(n7304), .A2(n7313), .ZN(n5974) );
  AND2_X1 U5855 ( .A1(n7386), .A2(n7422), .ZN(n4307) );
  AND2_X1 U5856 ( .A1(n8908), .A2(n8632), .ZN(n8942) );
  NAND2_X1 U5857 ( .A1(n7736), .A2(n4505), .ZN(n4308) );
  NAND2_X1 U5858 ( .A1(n7373), .A2(n7372), .ZN(n8106) );
  INV_X1 U5859 ( .A(n8106), .ZN(n4803) );
  AND2_X1 U5860 ( .A1(n7645), .A2(n7644), .ZN(n7747) );
  INV_X1 U5861 ( .A(n7747), .ZN(n9152) );
  NOR2_X1 U5862 ( .A1(n9082), .A2(n9059), .ZN(n4309) );
  NOR2_X1 U5863 ( .A1(n6759), .A2(n6758), .ZN(n4310) );
  INV_X1 U5864 ( .A(n5033), .ZN(n4693) );
  AND2_X1 U5865 ( .A1(n5035), .A2(n5023), .ZN(n5033) );
  NAND2_X1 U5866 ( .A1(n4887), .A2(n4886), .ZN(n4311) );
  NAND2_X1 U5867 ( .A1(n7385), .A2(n7386), .ZN(n7448) );
  INV_X1 U5868 ( .A(n4737), .ZN(n4736) );
  NAND2_X1 U5869 ( .A1(n4739), .A2(n4738), .ZN(n4737) );
  INV_X1 U5870 ( .A(n4521), .ZN(n4520) );
  NAND2_X1 U5871 ( .A1(n4522), .A2(n4296), .ZN(n4521) );
  AND3_X1 U5872 ( .A1(n5412), .A2(n5410), .A3(n5411), .ZN(n4312) );
  NAND2_X1 U5873 ( .A1(n9342), .A2(n7328), .ZN(n4313) );
  OR2_X1 U5874 ( .A1(n5015), .A2(n5014), .ZN(n5017) );
  INV_X1 U5875 ( .A(n5017), .ZN(n4688) );
  OR2_X1 U5876 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n4314) );
  AND2_X1 U5877 ( .A1(n4552), .A2(n4551), .ZN(n4315) );
  INV_X1 U5878 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4478) );
  INV_X1 U5879 ( .A(n4769), .ZN(n4768) );
  NAND2_X1 U5880 ( .A1(n4289), .A2(n4811), .ZN(n4769) );
  NAND2_X1 U5881 ( .A1(n7503), .A2(n7502), .ZN(n4316) );
  NAND2_X1 U5882 ( .A1(n4946), .A2(SI_5_), .ZN(n4317) );
  AND2_X1 U5883 ( .A1(n8730), .A2(n8571), .ZN(n4318) );
  INV_X1 U5884 ( .A(n4810), .ZN(n4809) );
  NAND2_X1 U5885 ( .A1(n7175), .A2(n7903), .ZN(n4810) );
  AND2_X1 U5886 ( .A1(n4638), .A2(n4637), .ZN(n4319) );
  NOR2_X1 U5887 ( .A1(n6971), .A2(n6818), .ZN(n4320) );
  NOR2_X1 U5888 ( .A1(n9362), .A2(n8248), .ZN(n4321) );
  INV_X1 U5889 ( .A(n8408), .ZN(n7584) );
  INV_X1 U5890 ( .A(n7424), .ZN(n4550) );
  OR2_X1 U5891 ( .A1(n7725), .A2(n4299), .ZN(n4322) );
  INV_X1 U5892 ( .A(n4615), .ZN(n4614) );
  OR2_X1 U5893 ( .A1(n7489), .A2(n4616), .ZN(n4615) );
  NAND2_X1 U5894 ( .A1(n8906), .A2(n4415), .ZN(n4323) );
  NAND2_X1 U5895 ( .A1(n7449), .A2(n7383), .ZN(n4324) );
  INV_X1 U5896 ( .A(n7625), .ZN(n8470) );
  OR2_X1 U5897 ( .A1(n9141), .A2(n8896), .ZN(n4325) );
  NOR2_X1 U5898 ( .A1(n4291), .A2(n4661), .ZN(n4660) );
  NOR2_X1 U5899 ( .A1(n8461), .A2(n4590), .ZN(n4326) );
  AND2_X1 U5900 ( .A1(n4476), .A2(n4474), .ZN(n4327) );
  NAND2_X1 U5901 ( .A1(n6896), .A2(n6895), .ZN(n4328) );
  AND2_X1 U5902 ( .A1(n4551), .A2(n4554), .ZN(n4329) );
  AND2_X1 U5903 ( .A1(n4842), .A2(n4776), .ZN(n4330) );
  OR2_X1 U5904 ( .A1(n8157), .A2(n4290), .ZN(n4331) );
  AND2_X1 U5905 ( .A1(n7280), .A2(n7273), .ZN(n4332) );
  AND2_X1 U5906 ( .A1(n8949), .A2(n4752), .ZN(n4333) );
  AND2_X1 U5907 ( .A1(n8699), .A2(n4402), .ZN(n4334) );
  AND2_X1 U5908 ( .A1(n4596), .A2(n4603), .ZN(n4335) );
  AND2_X1 U5909 ( .A1(n4854), .A2(n4617), .ZN(n5388) );
  INV_X1 U5910 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n4620) );
  NAND2_X1 U5911 ( .A1(n4597), .A2(n4602), .ZN(n4605) );
  INV_X1 U5912 ( .A(n9070), .ZN(n9433) );
  OAI211_X1 U5913 ( .C1(n6322), .C2(n7204), .A(n6007), .B(n6006), .ZN(n6209)
         );
  INV_X1 U5914 ( .A(n6209), .ZN(n9488) );
  INV_X1 U5915 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4474) );
  INV_X1 U5916 ( .A(n7640), .ZN(n4602) );
  NAND2_X1 U5917 ( .A1(n9028), .A2(n9027), .ZN(n9029) );
  XNOR2_X1 U5918 ( .A(n7247), .B(n7246), .ZN(n8608) );
  INV_X1 U5919 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5420) );
  NAND2_X1 U5920 ( .A1(n4831), .A2(n4830), .ZN(n5490) );
  AND2_X1 U5921 ( .A1(n6565), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4336) );
  AND2_X1 U5922 ( .A1(n4523), .A2(n4287), .ZN(n4337) );
  NAND2_X1 U5923 ( .A1(n4594), .A2(n6701), .ZN(n6706) );
  NOR3_X1 U5924 ( .A1(n9105), .A2(n4749), .A3(n9179), .ZN(n4751) );
  AND2_X1 U5925 ( .A1(n7846), .A2(n7845), .ZN(n4338) );
  INV_X1 U5926 ( .A(n5348), .ZN(n6348) );
  AND2_X1 U5927 ( .A1(n4575), .A2(n7260), .ZN(n4339) );
  NAND2_X1 U5928 ( .A1(n8234), .A2(n4444), .ZN(n4447) );
  NAND2_X1 U5929 ( .A1(n9128), .A2(n9216), .ZN(n4340) );
  INV_X1 U5930 ( .A(n6735), .ZN(n4517) );
  NOR2_X1 U5931 ( .A1(n6739), .A2(n6734), .ZN(n6735) );
  INV_X1 U5932 ( .A(n4747), .ZN(n9078) );
  NOR2_X1 U5933 ( .A1(n9105), .A2(n4749), .ZN(n4747) );
  AND2_X1 U5934 ( .A1(n4727), .A2(n6715), .ZN(n4341) );
  INV_X1 U5935 ( .A(n7056), .ZN(n4788) );
  INV_X1 U5936 ( .A(n7732), .ZN(n4509) );
  AND2_X1 U5937 ( .A1(n5584), .A2(n9694), .ZN(n9565) );
  AOI21_X1 U5938 ( .B1(n6380), .B2(n6385), .A(n6324), .ZN(n6641) );
  INV_X1 U5939 ( .A(n9413), .ZN(n4363) );
  NAND2_X1 U5940 ( .A1(n5944), .A2(n5943), .ZN(n6270) );
  INV_X1 U5941 ( .A(n6270), .ZN(n4449) );
  OR2_X1 U5942 ( .A1(n6075), .A2(n8736), .ZN(n6144) );
  OR2_X1 U5943 ( .A1(n9726), .A2(n4430), .ZN(n4342) );
  NAND2_X1 U5944 ( .A1(n6451), .A2(n7265), .ZN(n6784) );
  NAND2_X1 U5945 ( .A1(n4482), .A2(n5877), .ZN(n6070) );
  NAND2_X1 U5946 ( .A1(n4840), .A2(n4839), .ZN(n4844) );
  OR2_X1 U5947 ( .A1(n4844), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n4343) );
  NAND2_X1 U5948 ( .A1(n9235), .A2(n4736), .ZN(n4740) );
  INV_X1 U5949 ( .A(n7725), .ZN(n4497) );
  AND4_X1 U5950 ( .A1(n5583), .A2(n5582), .A3(n5581), .A4(n5580), .ZN(n5925)
         );
  INV_X1 U5951 ( .A(n8048), .ZN(n4668) );
  OR2_X1 U5952 ( .A1(n6086), .A2(n5784), .ZN(n6062) );
  INV_X1 U5953 ( .A(n6062), .ZN(n4744) );
  XNOR2_X1 U5954 ( .A(n5067), .B(n5066), .ZN(n5186) );
  AND2_X1 U5955 ( .A1(n5567), .A2(n9638), .ZN(n8266) );
  NAND2_X1 U5956 ( .A1(n7273), .A2(n7279), .ZN(n7403) );
  INV_X1 U5957 ( .A(n7403), .ZN(n5969) );
  NAND2_X1 U5958 ( .A1(n6732), .A2(n6731), .ZN(n9400) );
  INV_X1 U5959 ( .A(n9400), .ZN(n4738) );
  NAND2_X1 U5960 ( .A1(n5910), .A2(n5909), .ZN(n9693) );
  INV_X1 U5961 ( .A(n9693), .ZN(n4448) );
  AND2_X1 U5962 ( .A1(n5546), .A2(n5574), .ZN(n9624) );
  NAND2_X1 U5963 ( .A1(n5140), .A2(n5141), .ZN(n4532) );
  AND2_X1 U5964 ( .A1(n4673), .A2(n8070), .ZN(n4344) );
  AND2_X1 U5965 ( .A1(n8050), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4345) );
  AND2_X1 U5966 ( .A1(n4484), .A2(n4485), .ZN(n4346) );
  INV_X1 U5967 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n4534) );
  OAI222_X1 U5968 ( .A1(n8371), .A2(n9890), .B1(n4268), .B2(n5667), .C1(
        P2_U3152), .C2(n5668), .ZN(P2_U3356) );
  OAI222_X1 U5969 ( .A1(n8371), .A2(n5719), .B1(n4268), .B2(n5996), .C1(
        P2_U3152), .C2(n5722), .ZN(P2_U3353) );
  NAND2_X2 U5970 ( .A1(n7244), .A2(P2_U3152), .ZN(n8371) );
  OAI222_X1 U5971 ( .A1(n8371), .A2(n5692), .B1(n4268), .B2(n7204), .C1(
        P2_U3152), .C2(n5695), .ZN(P2_U3354) );
  OAI222_X1 U5972 ( .A1(n8371), .A2(n5679), .B1(n4268), .B2(n5771), .C1(
        P2_U3152), .C2(n5682), .ZN(P2_U3355) );
  OAI22_X1 U5973 ( .A1(n5961), .A2(P2_U3152), .B1(n8371), .B2(n7113), .ZN(
        n4481) );
  NAND2_X1 U5974 ( .A1(n5002), .A2(SI_9_), .ZN(n4347) );
  NOR2_X1 U5975 ( .A1(n4630), .A2(n7933), .ZN(n4629) );
  NAND2_X1 U5976 ( .A1(n4628), .A2(n4627), .ZN(n7889) );
  NAND2_X1 U5977 ( .A1(n4622), .A2(n4621), .ZN(n7877) );
  OAI21_X1 U5978 ( .B1(n4695), .B2(n4693), .A(n5035), .ZN(n4690) );
  OAI21_X1 U5979 ( .B1(n5097), .B2(n5096), .A(n5095), .ZN(n5113) );
  NAND2_X1 U5980 ( .A1(n6366), .A2(n8735), .ZN(n6195) );
  NAND2_X1 U5981 ( .A1(n6080), .A2(n8654), .ZN(n6366) );
  NAND2_X1 U5982 ( .A1(n8657), .A2(n8733), .ZN(n6080) );
  INV_X1 U5983 ( .A(n5881), .ZN(n8733) );
  NAND2_X1 U5984 ( .A1(n6097), .A2(n5880), .ZN(n8657) );
  NAND4_X1 U5985 ( .A1(n4734), .A2(n4367), .A3(n4366), .A4(n4365), .ZN(n4977)
         );
  NAND2_X1 U5986 ( .A1(n4608), .A2(n4371), .ZN(n4368) );
  NAND2_X1 U5987 ( .A1(n4368), .A2(n4369), .ZN(n8432) );
  NAND2_X1 U5988 ( .A1(n4888), .A2(n4376), .ZN(n4374) );
  NAND2_X1 U5989 ( .A1(n4888), .A2(n4886), .ZN(n4375) );
  INV_X1 U5990 ( .A(n6421), .ZN(n4386) );
  NAND2_X1 U5991 ( .A1(n4383), .A2(n6421), .ZN(n4384) );
  INV_X1 U5992 ( .A(n4822), .ZN(n4383) );
  OAI211_X1 U5993 ( .C1(n6414), .C2(n4386), .A(n4384), .B(n8378), .ZN(n8377)
         );
  NAND2_X1 U5994 ( .A1(n8377), .A2(n6429), .ZN(n6435) );
  NAND2_X1 U5995 ( .A1(n4385), .A2(n6421), .ZN(n8376) );
  NAND2_X1 U5996 ( .A1(n6414), .A2(n4822), .ZN(n4385) );
  OAI21_X1 U5997 ( .B1(n7625), .B2(n4273), .A(n4270), .ZN(n7641) );
  NAND2_X1 U5998 ( .A1(n7625), .A2(n4270), .ZN(n4388) );
  AND2_X2 U5999 ( .A1(n6876), .A2(n6875), .ZN(n6878) );
  NAND3_X1 U6000 ( .A1(n8629), .A2(n4303), .A3(n4393), .ZN(n4392) );
  AOI21_X1 U6001 ( .B1(n8540), .B2(n8678), .A(n8677), .ZN(n8542) );
  NAND2_X1 U6002 ( .A1(n4396), .A2(n4394), .ZN(n8540) );
  OR2_X1 U6003 ( .A1(n8534), .A2(n8628), .ZN(n4396) );
  INV_X1 U6004 ( .A(n6090), .ZN(n9480) );
  NAND3_X1 U6005 ( .A1(n4484), .A2(n4485), .A3(n5455), .ZN(n5459) );
  OR2_X2 U6006 ( .A1(n4399), .A2(n5370), .ZN(n5415) );
  INV_X1 U6007 ( .A(n4854), .ZN(n4989) );
  INV_X2 U6008 ( .A(n4992), .ZN(n4756) );
  NAND2_X1 U6009 ( .A1(n4400), .A2(n4334), .ZN(n7746) );
  NAND2_X1 U6010 ( .A1(n9021), .A2(n4404), .ZN(n4400) );
  NAND2_X2 U6011 ( .A1(n4407), .A2(n8667), .ZN(n9230) );
  NAND2_X1 U6012 ( .A1(n6621), .A2(n6620), .ZN(n4407) );
  AND2_X2 U6013 ( .A1(n4409), .A2(n4408), .ZN(n8779) );
  NAND2_X1 U6014 ( .A1(n6364), .A2(n6365), .ZN(n4408) );
  NAND2_X1 U6015 ( .A1(n8664), .A2(n6366), .ZN(n4409) );
  NAND2_X2 U6016 ( .A1(n5603), .A2(n5607), .ZN(n5463) );
  NAND2_X2 U6017 ( .A1(n4891), .A2(n4275), .ZN(n5607) );
  NAND2_X1 U6018 ( .A1(n8819), .A2(n6067), .ZN(n6353) );
  NOR2_X1 U6019 ( .A1(n8322), .A2(n8157), .ZN(n4429) );
  INV_X1 U6020 ( .A(n4429), .ZN(n8156) );
  AND4_X2 U6021 ( .A1(n4441), .A2(n4938), .A3(n4760), .A4(n4829), .ZN(n4840)
         );
  NAND4_X1 U6022 ( .A1(n4839), .A2(n4760), .A3(n4283), .A4(n4938), .ZN(n5065)
         );
  INV_X1 U6023 ( .A(n4447), .ZN(n8211) );
  NAND3_X1 U6024 ( .A1(n7272), .A2(n7384), .A3(n7269), .ZN(n7275) );
  NAND2_X1 U6025 ( .A1(n4452), .A2(n4451), .ZN(n7283) );
  NAND4_X1 U6026 ( .A1(n7282), .A2(n7281), .A3(n7286), .A4(n4453), .ZN(n4452)
         );
  NAND2_X1 U6027 ( .A1(n7384), .A2(n4332), .ZN(n4453) );
  NAND3_X1 U6028 ( .A1(n7431), .A2(n7397), .A3(n7427), .ZN(n4456) );
  NAND2_X1 U6029 ( .A1(n4840), .A2(n4836), .ZN(n5491) );
  NAND3_X1 U6030 ( .A1(n4461), .A2(n8118), .A3(n7370), .ZN(n4460) );
  NAND3_X1 U6031 ( .A1(n7367), .A2(n7366), .A3(n8126), .ZN(n4461) );
  NAND3_X1 U6032 ( .A1(n4466), .A2(n4464), .A3(n4462), .ZN(n7336) );
  AND2_X1 U6033 ( .A1(n4831), .A2(n4475), .ZN(n5540) );
  NAND2_X1 U6034 ( .A1(n4831), .A2(n4476), .ZN(n5060) );
  NAND2_X1 U6035 ( .A1(n4831), .A2(n4327), .ZN(n4473) );
  NAND3_X1 U6036 ( .A1(n5961), .A2(n5547), .A3(n8286), .ZN(n9696) );
  NAND2_X1 U6037 ( .A1(n6078), .A2(n5881), .ZN(n4482) );
  NAND2_X1 U6038 ( .A1(n6094), .A2(n6100), .ZN(n4483) );
  NAND2_X1 U6039 ( .A1(n9103), .A2(n4487), .ZN(n4486) );
  NAND2_X1 U6040 ( .A1(n4486), .A2(n4489), .ZN(n9050) );
  NAND2_X1 U6041 ( .A1(n8989), .A2(n4502), .ZN(n4501) );
  NAND2_X1 U6042 ( .A1(n6736), .A2(n4514), .ZN(n4510) );
  NAND2_X1 U6043 ( .A1(n4510), .A2(n4511), .ZN(n6927) );
  NAND2_X1 U6044 ( .A1(n6144), .A2(n4528), .ZN(n6317) );
  NAND2_X1 U6045 ( .A1(n4755), .A2(n4756), .ZN(n4894) );
  NAND3_X1 U6046 ( .A1(n4755), .A2(n4756), .A3(n4530), .ZN(n5401) );
  AOI21_X1 U6047 ( .B1(n7230), .B2(n7422), .A(n7229), .ZN(n7450) );
  NAND2_X1 U6048 ( .A1(n4315), .A2(n7389), .ZN(n4555) );
  AOI21_X1 U6049 ( .B1(n4552), .B2(n4329), .A(n4548), .ZN(n4553) );
  OAI21_X2 U6050 ( .B1(n6262), .B2(n6260), .A(n7306), .ZN(n6283) );
  NAND2_X1 U6051 ( .A1(n6119), .A2(n4558), .ZN(n4556) );
  NAND2_X1 U6052 ( .A1(n7191), .A2(n7190), .ZN(n8105) );
  NAND2_X1 U6053 ( .A1(n7191), .A2(n4561), .ZN(n4560) );
  NAND2_X1 U6054 ( .A1(n6451), .A2(n4567), .ZN(n9584) );
  NAND2_X1 U6055 ( .A1(n9584), .A2(n7323), .ZN(n6785) );
  OAI21_X1 U6056 ( .B1(n9322), .B2(n4573), .A(n4570), .ZN(n8206) );
  NAND2_X1 U6057 ( .A1(n9341), .A2(n4576), .ZN(n7181) );
  NAND2_X2 U6058 ( .A1(n9344), .A2(n6990), .ZN(n9341) );
  NAND2_X1 U6059 ( .A1(n4840), .A2(n4581), .ZN(n5071) );
  NAND2_X2 U6060 ( .A1(n8161), .A2(n7188), .ZN(n8168) );
  NAND2_X1 U6061 ( .A1(n7192), .A2(n7378), .ZN(n7230) );
  NAND2_X1 U6062 ( .A1(n5970), .A2(n5969), .ZN(n6134) );
  AOI21_X1 U6063 ( .B1(n8497), .B2(n7702), .A(n4584), .ZN(n4583) );
  AND2_X2 U6064 ( .A1(n8497), .A2(n4585), .ZN(n7788) );
  NAND2_X1 U6065 ( .A1(n8405), .A2(n4326), .ZN(n4586) );
  NAND2_X1 U6066 ( .A1(n4586), .A2(n4587), .ZN(n8414) );
  NAND2_X1 U6067 ( .A1(n7641), .A2(n4598), .ZN(n4595) );
  NAND2_X1 U6068 ( .A1(n4595), .A2(n4335), .ZN(n8426) );
  NAND2_X1 U6069 ( .A1(n6878), .A2(n4607), .ZN(n4606) );
  NAND2_X1 U6070 ( .A1(n7898), .A2(n4624), .ZN(n4622) );
  NAND2_X1 U6071 ( .A1(n7952), .A2(n4629), .ZN(n4628) );
  INV_X1 U6072 ( .A(n4639), .ZN(n6899) );
  INV_X1 U6073 ( .A(n5802), .ZN(n4659) );
  NAND2_X1 U6074 ( .A1(n4656), .A2(n4657), .ZN(n6049) );
  NAND2_X1 U6075 ( .A1(n5802), .A2(n4660), .ZN(n4656) );
  NOR2_X1 U6076 ( .A1(n6042), .A2(n4291), .ZN(n7791) );
  NAND2_X1 U6077 ( .A1(n4937), .A2(n4681), .ZN(n4680) );
  NAND2_X1 U6078 ( .A1(n4680), .A2(n4678), .ZN(n4955) );
  OAI21_X2 U6079 ( .B1(n4934), .B2(n4685), .A(n4905), .ZN(n4911) );
  NAND2_X1 U6080 ( .A1(n4698), .A2(n4700), .ZN(n5872) );
  NAND2_X1 U6081 ( .A1(n5832), .A2(n5834), .ZN(n4698) );
  NAND2_X1 U6082 ( .A1(n4702), .A2(n4703), .ZN(n5488) );
  NAND2_X1 U6083 ( .A1(n5115), .A2(n4706), .ZN(n4702) );
  NAND2_X1 U6084 ( .A1(n4712), .A2(n4714), .ZN(n7003) );
  NAND2_X1 U6085 ( .A1(n6834), .A2(n4716), .ZN(n4712) );
  NAND2_X1 U6086 ( .A1(n4726), .A2(n4341), .ZN(n6720) );
  INV_X1 U6087 ( .A(n4740), .ZN(n6847) );
  NAND2_X1 U6088 ( .A1(n6067), .A2(n6314), .ZN(n4742) );
  NAND2_X1 U6089 ( .A1(n4744), .A2(n4741), .ZN(n6487) );
  NAND2_X1 U6090 ( .A1(n9129), .A2(n4746), .ZN(n9243) );
  INV_X1 U6091 ( .A(n4751), .ZN(n9063) );
  NAND2_X1 U6092 ( .A1(n8990), .A2(n4333), .ZN(n8944) );
  NOR2_X1 U6093 ( .A1(n4992), .A2(n4758), .ZN(n4888) );
  NAND2_X1 U6094 ( .A1(n6103), .A2(n6090), .ZN(n6086) );
  NAND2_X2 U6095 ( .A1(n4759), .A2(n7756), .ZN(n5577) );
  NAND2_X1 U6096 ( .A1(n7090), .A2(n4762), .ZN(n4761) );
  NAND2_X1 U6097 ( .A1(n4761), .A2(n4763), .ZN(n8155) );
  NAND2_X1 U6098 ( .A1(n4772), .A2(n4770), .ZN(n6276) );
  NAND2_X1 U6099 ( .A1(n5941), .A2(n5940), .ZN(n6261) );
  INV_X1 U6100 ( .A(n5940), .ZN(n4774) );
  NAND2_X1 U6101 ( .A1(n7057), .A2(n4779), .ZN(n4778) );
  NAND2_X1 U6102 ( .A1(n8124), .A2(n4796), .ZN(n4795) );
  NAND2_X1 U6103 ( .A1(n6049), .A2(n6048), .ZN(n6515) );
  XNOR2_X1 U6104 ( .A(n7833), .B(n7831), .ZN(n7855) );
  NOR2_X1 U6105 ( .A1(n9393), .A2(n9519), .ZN(n9394) );
  XNOR2_X1 U6106 ( .A(n5673), .B(n9644), .ZN(n5561) );
  CLKBUF_X1 U6107 ( .A(n6134), .Z(n6301) );
  NAND2_X1 U6108 ( .A1(n5784), .A2(n4262), .ZN(n5772) );
  NAND2_X1 U6109 ( .A1(n6848), .A2(n6928), .ZN(n6937) );
  INV_X1 U6110 ( .A(n6435), .ZN(n6433) );
  NAND2_X1 U6111 ( .A1(n5647), .A2(n5646), .ZN(n5777) );
  NAND2_X1 U6112 ( .A1(n8821), .A2(n7497), .ZN(n5773) );
  OR2_X1 U6113 ( .A1(n6347), .A2(n5462), .ZN(n5466) );
  NAND2_X1 U6114 ( .A1(n5780), .A2(n5779), .ZN(n6005) );
  NAND2_X1 U6115 ( .A1(n5071), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5064) );
  OAI21_X2 U6116 ( .B1(n9564), .B2(n9560), .A(n9561), .ZN(n6596) );
  XNOR2_X1 U6117 ( .A(n7450), .B(n7449), .ZN(n7451) );
  NAND2_X1 U6118 ( .A1(n5404), .A2(n5403), .ZN(n6026) );
  AND2_X1 U6119 ( .A1(n7717), .A2(n7716), .ZN(n8953) );
  INV_X1 U6120 ( .A(n8810), .ZN(n6964) );
  OR2_X1 U6121 ( .A1(n9010), .A2(n8418), .ZN(n4812) );
  OR2_X1 U6122 ( .A1(n8513), .A2(n8436), .ZN(n4814) );
  OR2_X1 U6123 ( .A1(n7729), .A2(n9041), .ZN(n4816) );
  OR2_X1 U6124 ( .A1(n5669), .A2(n5552), .ZN(n4817) );
  NOR2_X1 U6125 ( .A1(n4917), .A2(n4929), .ZN(n4819) );
  NOR2_X1 U6126 ( .A1(n6639), .A2(n9223), .ZN(n4820) );
  OR2_X1 U6127 ( .A1(n5669), .A2(n5668), .ZN(n4821) );
  NAND2_X1 U6128 ( .A1(n7039), .A2(n7038), .ZN(n7231) );
  AND2_X1 U6129 ( .A1(n6549), .A2(n6413), .ZN(n4822) );
  INV_X1 U6130 ( .A(n9205), .ZN(n6928) );
  NAND2_X1 U6131 ( .A1(n7564), .A2(n8480), .ZN(n8405) );
  NAND2_X1 U6132 ( .A1(n7544), .A2(n8442), .ZN(n8445) );
  NAND2_X1 U6133 ( .A1(n6061), .A2(n9436), .ZN(n9070) );
  NOR2_X1 U6134 ( .A1(n6073), .A2(n6196), .ZN(n4823) );
  INV_X1 U6135 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n4825) );
  INV_X1 U6136 ( .A(n7448), .ZN(n7449) );
  NOR2_X1 U6137 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n4826) );
  INV_X1 U6138 ( .A(n8415), .ZN(n7624) );
  NOR2_X1 U6139 ( .A1(n7453), .A2(n7252), .ZN(n7454) );
  INV_X1 U6140 ( .A(n6135), .ZN(n5970) );
  OR2_X1 U6141 ( .A1(n7208), .A2(n7205), .ZN(n6018) );
  INV_X1 U6142 ( .A(n4263), .ZN(n6524) );
  INV_X1 U6143 ( .A(n6592), .ZN(n4881) );
  OR2_X1 U6144 ( .A1(n7829), .A2(n7828), .ZN(n7830) );
  INV_X1 U6145 ( .A(n6512), .ZN(n6513) );
  INV_X1 U6146 ( .A(n6605), .ZN(n6603) );
  INV_X1 U6147 ( .A(n9649), .ZN(n5923) );
  XNOR2_X1 U6148 ( .A(n5470), .B(n7675), .ZN(n5473) );
  INV_X1 U6149 ( .A(n7629), .ZN(n7465) );
  NAND2_X1 U6150 ( .A1(n7524), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5770) );
  INV_X1 U6151 ( .A(n5013), .ZN(n5014) );
  AND2_X1 U6152 ( .A1(n4962), .A2(n4965), .ZN(n4963) );
  OR2_X1 U6153 ( .A1(n7125), .A2(n7928), .ZN(n7134) );
  OR2_X1 U6154 ( .A1(n7134), .A2(n7900), .ZN(n7146) );
  OR3_X1 U6155 ( .A1(n6904), .A2(n6903), .A3(n6902), .ZN(n6981) );
  NAND2_X1 U6156 ( .A1(n5975), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6459) );
  INV_X1 U6157 ( .A(n9593), .ZN(n6779) );
  NOR2_X1 U6158 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4824) );
  INV_X1 U6159 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6154) );
  INV_X1 U6160 ( .A(n7206), .ZN(n7207) );
  OR2_X1 U6161 ( .A1(n7589), .A2(n9856), .ZN(n7608) );
  INV_X1 U6162 ( .A(n6574), .ZN(n6572) );
  OR2_X1 U6163 ( .A1(n7683), .A2(n7682), .ZN(n7710) );
  NAND2_X1 U6164 ( .A1(n7465), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n7631) );
  NAND2_X1 U6165 ( .A1(n9131), .A2(n8805), .ZN(n8902) );
  INV_X1 U6166 ( .A(n8737), .ZN(n6149) );
  INV_X1 U6167 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4863) );
  NAND2_X1 U6168 ( .A1(n5301), .A2(n5300), .ZN(n5430) );
  INV_X1 U6169 ( .A(n5042), .ZN(n5045) );
  NAND2_X1 U6170 ( .A1(n7460), .A2(n7235), .ZN(n7156) );
  NOR2_X1 U6171 ( .A1(n5807), .A2(n5806), .ZN(n5947) );
  AND2_X1 U6172 ( .A1(n7808), .A2(n7911), .ZN(n7809) );
  OR2_X1 U6173 ( .A1(n5579), .A2(n5555), .ZN(n5556) );
  OR2_X1 U6174 ( .A1(n7105), .A2(n7891), .ZN(n7124) );
  NAND2_X1 U6175 ( .A1(n7383), .A2(n7381), .ZN(n7441) );
  INV_X1 U6176 ( .A(n7984), .ZN(n7915) );
  AND2_X1 U6177 ( .A1(n7327), .A2(n9343), .ZN(n7414) );
  NAND2_X1 U6178 ( .A1(n7269), .A2(n9615), .ZN(n7402) );
  NAND2_X1 U6179 ( .A1(n5072), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5075) );
  OR2_X1 U6180 ( .A1(n7487), .A2(n7486), .ZN(n7488) );
  NAND2_X1 U6181 ( .A1(n6940), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7528) );
  OR2_X1 U6182 ( .A1(n7528), .A2(n7527), .ZN(n7549) );
  NAND2_X1 U6183 ( .A1(n6027), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6155) );
  INV_X1 U6184 ( .A(n5414), .ZN(n5449) );
  OR2_X1 U6185 ( .A1(n7778), .A2(n6026), .ZN(n7717) );
  INV_X1 U6186 ( .A(n8615), .ZN(n7772) );
  INV_X1 U6187 ( .A(n9073), .ZN(n9040) );
  INV_X1 U6188 ( .A(n9184), .ZN(n9082) );
  INV_X1 U6189 ( .A(n8812), .ZN(n6965) );
  AND2_X1 U6190 ( .A1(n6360), .A2(n6353), .ZN(n8736) );
  AND2_X1 U6191 ( .A1(n5879), .A2(n5878), .ZN(n9229) );
  OR2_X1 U6192 ( .A1(n9505), .A2(n8794), .ZN(n5446) );
  AND2_X1 U6193 ( .A1(n5487), .A2(n5436), .ZN(n5485) );
  XNOR2_X1 U6194 ( .A(n5295), .B(SI_14_), .ZN(n5294) );
  OR2_X1 U6195 ( .A1(n5949), .A2(n5912), .ZN(n5976) );
  OR3_X1 U6196 ( .A1(n6589), .A2(n6839), .A3(n6725), .ZN(n5736) );
  NAND2_X1 U6197 ( .A1(n5712), .A2(n5701), .ZN(n5706) );
  AND2_X1 U6198 ( .A1(n5188), .A2(n5187), .ZN(n9573) );
  INV_X1 U6199 ( .A(n8251), .ZN(n9621) );
  NAND2_X1 U6200 ( .A1(n7356), .A2(n7352), .ZN(n8198) );
  INV_X1 U6201 ( .A(n7418), .ZN(n8245) );
  INV_X1 U6202 ( .A(n9694), .ZN(n9719) );
  AND2_X1 U6203 ( .A1(n9691), .A2(n9696), .ZN(n9652) );
  AND2_X1 U6204 ( .A1(n5526), .A2(n5525), .ZN(n9630) );
  AND2_X1 U6205 ( .A1(n5028), .A2(n5036), .ZN(n6277) );
  AND2_X1 U6206 ( .A1(n7701), .A2(n7700), .ZN(n7703) );
  INV_X1 U6207 ( .A(n8519), .ZN(n8496) );
  AOI21_X1 U6208 ( .B1(n8947), .B2(n7571), .A(n7469), .ZN(n8899) );
  INV_X1 U6209 ( .A(n5124), .ZN(n5464) );
  INV_X1 U6210 ( .A(n9026), .ZN(n8917) );
  NAND2_X1 U6211 ( .A1(n8781), .A2(n8704), .ZN(n8963) );
  NAND2_X1 U6212 ( .A1(n8684), .A2(n9092), .ZN(n9102) );
  INV_X1 U6213 ( .A(n9229), .ZN(n9117) );
  AND2_X1 U6214 ( .A1(n5387), .A2(n9263), .ZN(n6391) );
  INV_X1 U6215 ( .A(n9515), .ZN(n9208) );
  OR2_X1 U6216 ( .A1(n8628), .A2(n8727), .ZN(n9505) );
  INV_X1 U6217 ( .A(n6391), .ZN(n6060) );
  AND2_X1 U6218 ( .A1(n5372), .A2(n5371), .ZN(n9262) );
  AND2_X1 U6219 ( .A1(n5507), .A2(n5762), .ZN(n8859) );
  XNOR2_X1 U6220 ( .A(n4945), .B(SI_5_), .ZN(n4943) );
  INV_X1 U6221 ( .A(n7903), .ZN(n8144) );
  NAND2_X1 U6222 ( .A1(n8265), .A2(n9628), .ZN(n8254) );
  OR2_X1 U6223 ( .A1(n8354), .A2(n8352), .ZN(n9742) );
  OR2_X1 U6224 ( .A1(n8354), .A2(n8353), .ZN(n9724) );
  AND2_X1 U6225 ( .A1(n5735), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9637) );
  INV_X1 U6226 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9835) );
  INV_X1 U6227 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5692) );
  INV_X1 U6228 ( .A(n9189), .ZN(n9091) );
  INV_X1 U6229 ( .A(n9210), .ZN(n6971) );
  INV_X1 U6230 ( .A(n9141), .ZN(n8897) );
  NAND2_X1 U6231 ( .A1(n7690), .A2(n7689), .ZN(n8896) );
  XNOR2_X1 U6232 ( .A(n8892), .B(n8915), .ZN(n9393) );
  OR3_X1 U6233 ( .A1(n9321), .A2(n8725), .A3(n7762), .ZN(n9121) );
  INV_X1 U6234 ( .A(n9544), .ZN(n9541) );
  INV_X1 U6235 ( .A(n9528), .ZN(n9526) );
  CLKBUF_X1 U6236 ( .A(n9453), .Z(n9467) );
  INV_X1 U6237 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5032) );
  NOR2_X1 U6238 ( .A1(n5350), .A2(n9930), .ZN(n9929) );
  NOR2_X1 U6239 ( .A1(n6687), .A2(n9929), .ZN(n9773) );
  NOR2_X2 U6240 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n4907) );
  AND2_X2 U6241 ( .A1(n4907), .A2(n4824), .ZN(n4938) );
  INV_X1 U6242 ( .A(n5491), .ZN(n4831) );
  INV_X2 U6243 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4830) );
  INV_X2 U6244 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5058) );
  NAND2_X1 U6245 ( .A1(n5059), .A2(n5058), .ZN(n4832) );
  NAND2_X1 U6246 ( .A1(n4832), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4847) );
  INV_X1 U6247 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9778) );
  NAND2_X1 U6248 ( .A1(n4847), .A2(n9778), .ZN(n4849) );
  NAND2_X1 U6249 ( .A1(n4849), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4833) );
  NOR2_X1 U6250 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n4834) );
  NAND4_X1 U6251 ( .A1(n4834), .A2(n4478), .A3(n4830), .A4(n5541), .ZN(n4838)
         );
  INV_X2 U6252 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5543) );
  NAND4_X1 U6253 ( .A1(n5058), .A2(n4836), .A3(n5543), .A4(n4835), .ZN(n4837)
         );
  NOR2_X1 U6254 ( .A1(n4838), .A2(n4837), .ZN(n4839) );
  NAND2_X1 U6255 ( .A1(n4343), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4841) );
  MUX2_X1 U6256 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4841), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n4843) );
  INV_X1 U6257 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4842) );
  NAND2_X1 U6258 ( .A1(n4843), .A2(n5065), .ZN(n6839) );
  NAND2_X1 U6259 ( .A1(n4844), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4845) );
  MUX2_X1 U6260 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4845), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n4846) );
  NAND2_X1 U6261 ( .A1(n4846), .A2(n4343), .ZN(n6725) );
  OR2_X1 U6262 ( .A1(n4847), .A2(n9778), .ZN(n4848) );
  NAND2_X1 U6263 ( .A1(n4849), .A2(n4848), .ZN(n5735) );
  INV_X1 U6264 ( .A(n9637), .ZN(n4850) );
  OR2_X1 U6265 ( .A1(n5736), .A2(n4850), .ZN(n7982) );
  INV_X1 U6266 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5008) );
  INV_X1 U6267 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5107) );
  INV_X1 U6268 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4856) );
  INV_X1 U6269 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4855) );
  NAND4_X1 U6270 ( .A1(n4857), .A2(n5107), .A3(n4856), .A4(n4855), .ZN(n4861)
         );
  INV_X1 U6271 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5309) );
  INV_X1 U6272 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5505) );
  INV_X1 U6273 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n4859) );
  INV_X1 U6274 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n4858) );
  NAND4_X1 U6275 ( .A1(n5309), .A2(n5505), .A3(n4859), .A4(n4858), .ZN(n4860)
         );
  INV_X1 U6276 ( .A(n4872), .ZN(n4862) );
  NAND2_X1 U6277 ( .A1(n5388), .A2(n4863), .ZN(n5391) );
  INV_X1 U6278 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n4866) );
  NAND2_X1 U6279 ( .A1(n4867), .A2(n4866), .ZN(n4868) );
  OR2_X1 U6280 ( .A1(n4867), .A2(n4866), .ZN(n4869) );
  NAND2_X1 U6281 ( .A1(n5449), .A2(n8794), .ZN(n8720) );
  NOR2_X1 U6282 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n4871) );
  NOR3_X1 U6283 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .A3(
        P1_IR_REG_9__SCAN_IN), .ZN(n4870) );
  INV_X1 U6284 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4880) );
  INV_X1 U6285 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4875) );
  NAND2_X1 U6286 ( .A1(n4876), .A2(n4875), .ZN(n4878) );
  INV_X1 U6287 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4873) );
  NAND2_X1 U6288 ( .A1(n4878), .A2(n4877), .ZN(n6726) );
  INV_X1 U6289 ( .A(n6726), .ZN(n4882) );
  XNOR2_X1 U6290 ( .A(n4879), .B(n4880), .ZN(n6592) );
  NAND2_X1 U6291 ( .A1(n8720), .A2(n5415), .ZN(n4885) );
  INV_X1 U6292 ( .A(n4888), .ZN(n4883) );
  NAND2_X1 U6293 ( .A1(n4883), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4884) );
  XNOR2_X1 U6294 ( .A(n4884), .B(n4886), .ZN(n6506) );
  NAND2_X1 U6295 ( .A1(n4885), .A2(n6506), .ZN(n5145) );
  NOR3_X1 U6296 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .A3(
        P1_IR_REG_25__SCAN_IN), .ZN(n4887) );
  INV_X1 U6297 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4889) );
  NAND2_X1 U6298 ( .A1(n4894), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4890) );
  NAND2_X1 U6299 ( .A1(n4892), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4893) );
  NAND2_X1 U6300 ( .A1(n5145), .A2(n6932), .ZN(n4896) );
  NAND2_X1 U6301 ( .A1(n4896), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U6302 ( .A(n6506), .ZN(n4897) );
  NOR2_X1 U6303 ( .A1(n5415), .A2(n4897), .ZN(n5121) );
  XNOR2_X1 U6304 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  NAND2_X1 U6305 ( .A1(n6693), .A2(n4898), .ZN(n4901) );
  NAND2_X4 U6306 ( .A1(n4901), .A2(n4900), .ZN(n4913) );
  INV_X1 U6307 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9890) );
  NOR2_X1 U6308 ( .A1(n7244), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6509) );
  AND2_X1 U6309 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4902) );
  NAND2_X1 U6310 ( .A1(n5461), .A2(n4902), .ZN(n5566) );
  NAND3_X1 U6311 ( .A1(n4913), .A2(SI_0_), .A3(P2_DATAO_REG_0__SCAN_IN), .ZN(
        n4903) );
  MUX2_X1 U6312 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n4913), .Z(n4933) );
  NAND2_X1 U6313 ( .A1(n4904), .A2(SI_1_), .ZN(n4905) );
  MUX2_X1 U6314 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n4913), .Z(n4912) );
  INV_X1 U6315 ( .A(SI_2_), .ZN(n4906) );
  XNOR2_X1 U6316 ( .A(n4912), .B(n4906), .ZN(n4910) );
  XNOR2_X1 U6317 ( .A(n4911), .B(n4910), .ZN(n5667) );
  INV_X1 U6318 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4909) );
  INV_X1 U6319 ( .A(n4907), .ZN(n4931) );
  NAND2_X1 U6320 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4931), .ZN(n4908) );
  XNOR2_X1 U6321 ( .A(n4909), .B(n4908), .ZN(n5668) );
  INV_X1 U6322 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n5719) );
  NAND2_X1 U6323 ( .A1(n4911), .A2(n4910), .ZN(n4928) );
  NAND2_X1 U6324 ( .A1(n4912), .A2(SI_2_), .ZN(n4927) );
  INV_X1 U6325 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n4981) );
  MUX2_X1 U6326 ( .A(n5679), .B(n4981), .S(n4913), .Z(n4916) );
  INV_X1 U6327 ( .A(n4916), .ZN(n4914) );
  NAND2_X1 U6328 ( .A1(n4914), .A2(SI_3_), .ZN(n4915) );
  AND2_X1 U6329 ( .A1(n4927), .A2(n4915), .ZN(n4918) );
  INV_X1 U6330 ( .A(n4915), .ZN(n4917) );
  XNOR2_X1 U6331 ( .A(n4916), .B(SI_3_), .ZN(n4929) );
  AOI21_X2 U6332 ( .B1(n4928), .B2(n4918), .A(n4819), .ZN(n4937) );
  MUX2_X1 U6333 ( .A(n5692), .B(n4919), .S(n4913), .Z(n4920) );
  INV_X1 U6334 ( .A(n4920), .ZN(n4921) );
  NAND2_X1 U6335 ( .A1(n4921), .A2(SI_4_), .ZN(n4922) );
  INV_X1 U6336 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n4986) );
  MUX2_X1 U6337 ( .A(n5719), .B(n4986), .S(n4913), .Z(n4945) );
  XNOR2_X1 U6338 ( .A(n4944), .B(n4943), .ZN(n5996) );
  NAND2_X1 U6339 ( .A1(n4923), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4924) );
  MUX2_X1 U6340 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4924), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n4926) );
  NAND2_X1 U6341 ( .A1(n4926), .A2(n4925), .ZN(n5722) );
  NAND2_X1 U6342 ( .A1(n4928), .A2(n4927), .ZN(n4930) );
  XNOR2_X1 U6343 ( .A(n4930), .B(n4929), .ZN(n5771) );
  OAI21_X1 U6344 ( .B1(P2_IR_REG_2__SCAN_IN), .B2(n4931), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n4932) );
  XNOR2_X1 U6345 ( .A(n4932), .B(P2_IR_REG_3__SCAN_IN), .ZN(n5220) );
  INV_X1 U6346 ( .A(n5220), .ZN(n5682) );
  INV_X1 U6347 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5553) );
  XNOR2_X1 U6348 ( .A(n4934), .B(n4933), .ZN(n5460) );
  INV_X1 U6349 ( .A(n5460), .ZN(n5551) );
  NAND2_X1 U6350 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4935) );
  INV_X1 U6351 ( .A(n9282), .ZN(n5552) );
  XNOR2_X1 U6352 ( .A(n4937), .B(n4936), .ZN(n7204) );
  OR2_X1 U6353 ( .A1(n4938), .A2(n5539), .ZN(n4940) );
  XNOR2_X1 U6354 ( .A(n4940), .B(n4939), .ZN(n5695) );
  NAND2_X1 U6355 ( .A1(n7244), .A2(P1_U3084), .ZN(n6728) );
  OAI222_X1 U6356 ( .A1(n9275), .A2(n5462), .B1(n6728), .B2(n5551), .C1(
        P1_U3084), .C2(n5124), .ZN(P1_U3352) );
  INV_X1 U6357 ( .A(n4945), .ZN(n4946) );
  INV_X1 U6358 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n4947) );
  INV_X1 U6359 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n4988) );
  MUX2_X1 U6360 ( .A(n4947), .B(n4988), .S(n7244), .Z(n4948) );
  NAND2_X1 U6361 ( .A1(n4955), .A2(n4954), .ZN(n4964) );
  INV_X1 U6362 ( .A(n4948), .ZN(n4949) );
  NAND2_X1 U6363 ( .A1(n4949), .A2(SI_6_), .ZN(n4962) );
  NAND2_X1 U6364 ( .A1(n4964), .A2(n4962), .ZN(n4951) );
  MUX2_X1 U6365 ( .A(n4950), .B(n4991), .S(n4913), .Z(n4960) );
  XNOR2_X1 U6366 ( .A(n4951), .B(n4966), .ZN(n6321) );
  NOR2_X1 U6367 ( .A1(n4925), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n4974) );
  INV_X1 U6368 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5539) );
  OR2_X1 U6369 ( .A1(n4974), .A2(n5539), .ZN(n4952) );
  XNOR2_X1 U6370 ( .A(n4952), .B(P2_IR_REG_7__SCAN_IN), .ZN(n5936) );
  INV_X1 U6371 ( .A(n8371), .ZN(n5494) );
  AOI22_X1 U6372 ( .A1(n5936), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n5494), .ZN(n4953) );
  OAI21_X1 U6373 ( .B1(n6321), .B2(n4268), .A(n4953), .ZN(P2_U3351) );
  XNOR2_X1 U6374 ( .A(n4955), .B(n4954), .ZN(n6148) );
  NAND2_X1 U6375 ( .A1(n4925), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4956) );
  XNOR2_X1 U6376 ( .A(n4956), .B(P2_IR_REG_6__SCAN_IN), .ZN(n5796) );
  AOI22_X1 U6377 ( .A1(n5796), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n5494), .ZN(n4957) );
  OAI21_X1 U6378 ( .B1(n6148), .B2(n4268), .A(n4957), .ZN(P2_U3352) );
  CLKBUF_X1 U6379 ( .A(n6728), .Z(n9273) );
  INV_X1 U6380 ( .A(n9275), .ZN(n9265) );
  XNOR2_X1 U6381 ( .A(n4958), .B(P1_IR_REG_2__SCAN_IN), .ZN(n5648) );
  AOI22_X1 U6382 ( .A1(n9265), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n5648), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n4959) );
  OAI21_X1 U6383 ( .B1(n5667), .B2(n9273), .A(n4959), .ZN(P1_U3351) );
  INV_X1 U6384 ( .A(n4960), .ZN(n4961) );
  NAND2_X1 U6385 ( .A1(n4964), .A2(n4963), .ZN(n4998) );
  INV_X1 U6386 ( .A(n4965), .ZN(n4967) );
  AND2_X1 U6387 ( .A1(n4998), .A2(n4996), .ZN(n4972) );
  INV_X1 U6388 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n4968) );
  MUX2_X1 U6389 ( .A(n4968), .B(n6334), .S(n4913), .Z(n4969) );
  INV_X1 U6390 ( .A(SI_8_), .ZN(n9846) );
  NAND2_X1 U6391 ( .A1(n4969), .A2(n9846), .ZN(n4995) );
  INV_X1 U6392 ( .A(n4969), .ZN(n4970) );
  NAND2_X1 U6393 ( .A1(n4995), .A2(n4999), .ZN(n4971) );
  XNOR2_X1 U6394 ( .A(n4972), .B(n4971), .ZN(n6330) );
  INV_X1 U6395 ( .A(n6330), .ZN(n4994) );
  NAND2_X1 U6396 ( .A1(n4974), .A2(n4973), .ZN(n5004) );
  NAND2_X1 U6397 ( .A1(n5004), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4975) );
  XNOR2_X1 U6398 ( .A(n4975), .B(P2_IR_REG_8__SCAN_IN), .ZN(n5942) );
  AOI22_X1 U6399 ( .A1(n5942), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n5494), .ZN(n4976) );
  OAI21_X1 U6400 ( .B1(n4994), .B2(n4268), .A(n4976), .ZN(P2_U3350) );
  NAND2_X1 U6401 ( .A1(n4978), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4979) );
  MUX2_X1 U6402 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4979), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n4980) );
  AND2_X1 U6403 ( .A1(n4977), .A2(n4980), .ZN(n5768) );
  INV_X1 U6404 ( .A(n5768), .ZN(n5337) );
  OAI222_X1 U6405 ( .A1(n9275), .A2(n4981), .B1(n9273), .B2(n5771), .C1(
        P1_U3084), .C2(n5337), .ZN(P1_U3350) );
  NOR2_X1 U6406 ( .A1(n4982), .A2(n5306), .ZN(n4983) );
  MUX2_X1 U6407 ( .A(n5306), .B(n4983), .S(P1_IR_REG_5__SCAN_IN), .Z(n4985) );
  OR2_X1 U6408 ( .A1(n4985), .A2(n4984), .ZN(n5139) );
  OAI222_X1 U6409 ( .A1(n9275), .A2(n4986), .B1(n9273), .B2(n5996), .C1(
        P1_U3084), .C2(n5139), .ZN(P1_U3348) );
  OR2_X1 U6410 ( .A1(n4984), .A2(n5306), .ZN(n4987) );
  XNOR2_X1 U6411 ( .A(n4987), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6145) );
  INV_X1 U6412 ( .A(n6145), .ZN(n5173) );
  OAI222_X1 U6413 ( .A1(n9275), .A2(n4988), .B1(n9273), .B2(n6148), .C1(
        P1_U3084), .C2(n5173), .ZN(P1_U3347) );
  NAND2_X1 U6414 ( .A1(n4989), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4990) );
  XNOR2_X1 U6415 ( .A(n4990), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6318) );
  INV_X1 U6416 ( .A(n6318), .ZN(n5281) );
  OAI222_X1 U6417 ( .A1(n9275), .A2(n4991), .B1(n9273), .B2(n6321), .C1(
        P1_U3084), .C2(n5281), .ZN(P1_U3346) );
  NAND2_X1 U6418 ( .A1(n4992), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4993) );
  XNOR2_X1 U6419 ( .A(n4993), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6331) );
  INV_X1 U6420 ( .A(n6331), .ZN(n5284) );
  OAI222_X1 U6421 ( .A1(n9275), .A2(n6334), .B1(n9273), .B2(n4994), .C1(
        P1_U3084), .C2(n5284), .ZN(P1_U3345) );
  NOR2_X1 U6422 ( .A1(n5018), .A2(n5015), .ZN(n5003) );
  MUX2_X1 U6423 ( .A(n9835), .B(n9891), .S(n4913), .Z(n5001) );
  INV_X1 U6424 ( .A(SI_9_), .ZN(n5000) );
  INV_X1 U6425 ( .A(n5001), .ZN(n5002) );
  XNOR2_X1 U6426 ( .A(n5003), .B(n5013), .ZN(n6346) );
  INV_X1 U6427 ( .A(n6346), .ZN(n5012) );
  NAND2_X1 U6428 ( .A1(n5024), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5005) );
  XNOR2_X1 U6429 ( .A(n5005), .B(P2_IR_REG_9__SCAN_IN), .ZN(n5908) );
  INV_X1 U6430 ( .A(n5908), .ZN(n5006) );
  OAI222_X1 U6431 ( .A1(n4268), .A2(n5012), .B1(n5006), .B2(P2_U3152), .C1(
        n9835), .C2(n8371), .ZN(P2_U3349) );
  OR2_X1 U6432 ( .A1(n5007), .A2(n5306), .ZN(n5009) );
  MUX2_X1 U6433 ( .A(n5009), .B(P1_IR_REG_31__SCAN_IN), .S(n5008), .Z(n5011)
         );
  NAND2_X1 U6434 ( .A1(n5011), .A2(n5010), .ZN(n5348) );
  OAI222_X1 U6435 ( .A1(n9275), .A2(n9891), .B1(n6728), .B2(n5012), .C1(n5348), 
        .C2(P1_U3084), .ZN(P1_U3344) );
  INV_X1 U6436 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5019) );
  MUX2_X1 U6437 ( .A(n5019), .B(n5032), .S(n7244), .Z(n5021) );
  INV_X1 U6438 ( .A(SI_10_), .ZN(n5020) );
  INV_X1 U6439 ( .A(n5021), .ZN(n5022) );
  NAND2_X1 U6440 ( .A1(n5022), .A2(SI_10_), .ZN(n5023) );
  XNOR2_X1 U6441 ( .A(n5034), .B(n5033), .ZN(n6564) );
  INV_X1 U6442 ( .A(n6564), .ZN(n5031) );
  NOR2_X1 U6443 ( .A1(n5024), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5054) );
  OR2_X1 U6444 ( .A1(n5054), .A2(n5539), .ZN(n5027) );
  INV_X1 U6445 ( .A(n5027), .ZN(n5025) );
  NAND2_X1 U6446 ( .A1(n5025), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n5028) );
  NAND2_X1 U6447 ( .A1(n5027), .A2(n5026), .ZN(n5036) );
  AOI22_X1 U6448 ( .A1(n6277), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n5494), .ZN(n5029) );
  OAI21_X1 U6449 ( .B1(n5031), .B2(n4268), .A(n5029), .ZN(P2_U3348) );
  NAND2_X1 U6450 ( .A1(n5010), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5030) );
  XNOR2_X1 U6451 ( .A(n5030), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6565) );
  INV_X1 U6452 ( .A(n6565), .ZN(n5515) );
  OAI222_X1 U6453 ( .A1(n9275), .A2(n5032), .B1(n6728), .B2(n5031), .C1(n5515), 
        .C2(P1_U3084), .ZN(P1_U3343) );
  MUX2_X1 U6454 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n7244), .Z(n5043) );
  INV_X1 U6455 ( .A(SI_11_), .ZN(n9873) );
  XNOR2_X1 U6456 ( .A(n5046), .B(n5042), .ZN(n6617) );
  INV_X1 U6457 ( .A(n6617), .ZN(n5040) );
  NAND2_X1 U6458 ( .A1(n5036), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5037) );
  XNOR2_X1 U6459 ( .A(n5037), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6452) );
  INV_X1 U6460 ( .A(n6452), .ZN(n5643) );
  INV_X1 U6461 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5038) );
  OAI222_X1 U6462 ( .A1(n4268), .A2(n5040), .B1(n5643), .B2(P2_U3152), .C1(
        n5038), .C2(n8371), .ZN(P2_U3347) );
  INV_X1 U6463 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5041) );
  OR2_X1 U6464 ( .A1(n5010), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5050) );
  NAND2_X1 U6465 ( .A1(n5050), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5039) );
  XNOR2_X1 U6466 ( .A(n5039), .B(P1_IR_REG_11__SCAN_IN), .ZN(n8828) );
  INV_X1 U6467 ( .A(n8828), .ZN(n5847) );
  OAI222_X1 U6468 ( .A1(n9275), .A2(n5041), .B1(n6728), .B2(n5040), .C1(n5847), 
        .C2(P1_U3084), .ZN(P1_U3342) );
  INV_X1 U6469 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5052) );
  NAND2_X1 U6470 ( .A1(n5043), .A2(SI_11_), .ZN(n5044) );
  INV_X1 U6471 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n5057) );
  MUX2_X1 U6472 ( .A(n5057), .B(n5052), .S(n7244), .Z(n5047) );
  INV_X1 U6473 ( .A(SI_12_), .ZN(n9832) );
  INV_X1 U6474 ( .A(n5047), .ZN(n5048) );
  NAND2_X1 U6475 ( .A1(n5048), .A2(SI_12_), .ZN(n5049) );
  XNOR2_X1 U6476 ( .A(n5097), .B(n5096), .ZN(n6729) );
  INV_X1 U6477 ( .A(n6729), .ZN(n5056) );
  NAND2_X1 U6478 ( .A1(n5105), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5051) );
  XNOR2_X1 U6479 ( .A(n5051), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6730) );
  INV_X1 U6480 ( .A(n6730), .ZN(n5845) );
  OAI222_X1 U6481 ( .A1(n9275), .A2(n5052), .B1(n6728), .B2(n5056), .C1(
        P1_U3084), .C2(n5845), .ZN(P1_U3341) );
  NOR2_X1 U6482 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5053) );
  NAND2_X1 U6483 ( .A1(n5054), .A2(n5053), .ZN(n5102) );
  NAND2_X1 U6484 ( .A1(n5102), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5055) );
  XNOR2_X1 U6485 ( .A(n5055), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6600) );
  INV_X1 U6486 ( .A(n6600), .ZN(n5860) );
  NAND2_X1 U6487 ( .A1(n5736), .A2(n9637), .ZN(n9631) );
  INV_X1 U6488 ( .A(n9631), .ZN(n8277) );
  INV_X1 U6489 ( .A(n5961), .ZN(n5548) );
  NAND2_X1 U6490 ( .A1(n5060), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5061) );
  INV_X1 U6491 ( .A(n7253), .ZN(n7429) );
  NAND2_X1 U6492 ( .A1(n5548), .A2(n7429), .ZN(n5575) );
  INV_X1 U6493 ( .A(n5575), .ZN(n5546) );
  NAND2_X1 U6494 ( .A1(n8277), .A2(n5546), .ZN(n5070) );
  INV_X1 U6495 ( .A(n5735), .ZN(n5062) );
  NAND2_X1 U6496 ( .A1(n5062), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7438) );
  NAND2_X1 U6497 ( .A1(n9631), .A2(n7438), .ZN(n5068) );
  INV_X1 U6498 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5063) );
  INV_X1 U6499 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5066) );
  NAND2_X1 U6500 ( .A1(n5068), .A2(n7079), .ZN(n5069) );
  AND2_X1 U6501 ( .A1(n5070), .A2(n5069), .ZN(n8072) );
  INV_X1 U6502 ( .A(n8072), .ZN(n9578) );
  NOR2_X1 U6503 ( .A1(n9578), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U6504 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n5085) );
  NOR2_X2 U6505 ( .A1(n5071), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n5073) );
  INV_X1 U6506 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5072) );
  NAND2_X1 U6507 ( .A1(n5073), .A2(n5072), .ZN(n5078) );
  OR2_X1 U6508 ( .A1(n5073), .A2(n5539), .ZN(n5074) );
  NAND2_X1 U6509 ( .A1(n5074), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n5076) );
  NAND2_X2 U6510 ( .A1(n5078), .A2(n5077), .ZN(n7756) );
  INV_X1 U6511 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8370) );
  XNOR2_X2 U6512 ( .A(n5079), .B(n8370), .ZN(n7040) );
  INV_X1 U6513 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n5083) );
  NAND2_X1 U6514 ( .A1(n7222), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5082) );
  INV_X1 U6515 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n5080) );
  OR2_X1 U6516 ( .A1(n7224), .A2(n5080), .ZN(n5081) );
  OAI211_X1 U6517 ( .C1(n7228), .C2(n5083), .A(n5082), .B(n5081), .ZN(n8074)
         );
  NAND2_X1 U6518 ( .A1(P2_U3966), .A2(n8074), .ZN(n5084) );
  OAI21_X1 U6519 ( .B1(P2_U3966), .B2(n5085), .A(n5084), .ZN(P2_U3583) );
  INV_X1 U6520 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5094) );
  INV_X1 U6521 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6175) );
  OR2_X1 U6522 ( .A1(n5696), .A2(n6175), .ZN(n5092) );
  INV_X1 U6523 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5087) );
  OR2_X1 U6524 ( .A1(n5579), .A2(n5087), .ZN(n5091) );
  INV_X1 U6525 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5088) );
  NAND2_X1 U6526 ( .A1(n5576), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5089) );
  NAND4_X2 U6527 ( .A1(n5092), .A2(n5091), .A3(n5090), .A4(n5089), .ZN(n5567)
         );
  NAND2_X1 U6528 ( .A1(P2_U3966), .A2(n5567), .ZN(n5093) );
  OAI21_X1 U6529 ( .B1(P2_U3966), .B2(n5094), .A(n5093), .ZN(P2_U3552) );
  INV_X1 U6530 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n5104) );
  INV_X1 U6531 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5111) );
  MUX2_X1 U6532 ( .A(n5104), .B(n5111), .S(n7244), .Z(n5099) );
  INV_X1 U6533 ( .A(SI_13_), .ZN(n5098) );
  NAND2_X1 U6534 ( .A1(n5099), .A2(n5098), .ZN(n5114) );
  INV_X1 U6535 ( .A(n5099), .ZN(n5100) );
  NAND2_X1 U6536 ( .A1(n5100), .A2(SI_13_), .ZN(n5101) );
  XNOR2_X1 U6537 ( .A(n5113), .B(n5112), .ZN(n6800) );
  INV_X1 U6538 ( .A(n6800), .ZN(n5110) );
  OR2_X1 U6539 ( .A1(n5102), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5103) );
  NAND2_X1 U6540 ( .A1(n5103), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5118) );
  XNOR2_X1 U6541 ( .A(n5118), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6762) );
  INV_X1 U6542 ( .A(n6762), .ZN(n5898) );
  OAI222_X1 U6543 ( .A1(n4268), .A2(n5110), .B1(n5898), .B2(P2_U3152), .C1(
        n5104), .C2(n8371), .ZN(P2_U3345) );
  NOR2_X1 U6544 ( .A1(n5105), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5305) );
  OR2_X1 U6545 ( .A1(n5305), .A2(n5306), .ZN(n5108) );
  INV_X1 U6546 ( .A(n5108), .ZN(n5106) );
  NAND2_X1 U6547 ( .A1(n5106), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n5109) );
  NAND2_X1 U6548 ( .A1(n5108), .A2(n5107), .ZN(n5157) );
  INV_X1 U6549 ( .A(n6861), .ZN(n6236) );
  OAI222_X1 U6550 ( .A1(n9275), .A2(n5111), .B1(n6728), .B2(n5110), .C1(n6236), 
        .C2(P1_U3084), .ZN(P1_U3340) );
  NAND2_X1 U6551 ( .A1(n5113), .A2(n5112), .ZN(n5115) );
  INV_X1 U6552 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n5116) );
  INV_X1 U6553 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n5160) );
  MUX2_X1 U6554 ( .A(n5116), .B(n5160), .S(n7244), .Z(n5295) );
  XNOR2_X1 U6555 ( .A(n5299), .B(n5294), .ZN(n6889) );
  INV_X1 U6556 ( .A(n6889), .ZN(n5159) );
  NAND2_X1 U6557 ( .A1(n5118), .A2(n5117), .ZN(n5119) );
  NAND2_X1 U6558 ( .A1(n5119), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5313) );
  XNOR2_X1 U6559 ( .A(n5313), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8000) );
  AOI22_X1 U6560 ( .A1(n8000), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n5494), .ZN(n5120) );
  OAI21_X1 U6561 ( .B1(n5159), .B2(n4268), .A(n5120), .ZN(P2_U3344) );
  INV_X1 U6562 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n5144) );
  OR2_X1 U6563 ( .A1(P1_U3083), .A2(n5121), .ZN(n9426) );
  NOR2_X1 U6564 ( .A1(n5603), .A2(P1_U3084), .ZN(n6925) );
  NAND2_X1 U6565 ( .A1(n5145), .A2(n6925), .ZN(n8878) );
  INV_X1 U6566 ( .A(n8878), .ZN(n5122) );
  AND2_X1 U6567 ( .A1(n5122), .A2(n5607), .ZN(n9413) );
  AND2_X1 U6568 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6554) );
  INV_X1 U6569 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9537) );
  MUX2_X1 U6570 ( .A(n9537), .B(P1_REG1_REG_6__SCAN_IN), .S(n6145), .Z(n5131)
         );
  INV_X1 U6571 ( .A(n5139), .ZN(n5994) );
  NAND2_X1 U6572 ( .A1(n4977), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5123) );
  XNOR2_X1 U6573 ( .A(n5123), .B(P1_IR_REG_4__SCAN_IN), .ZN(n7202) );
  XNOR2_X1 U6574 ( .A(n5124), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n5361) );
  AND2_X1 U6575 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n5360) );
  NAND2_X1 U6576 ( .A1(n5361), .A2(n5360), .ZN(n5359) );
  NAND2_X1 U6577 ( .A1(n5464), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5125) );
  NAND2_X1 U6578 ( .A1(n5359), .A2(n5125), .ZN(n5623) );
  INV_X1 U6579 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9531) );
  MUX2_X1 U6580 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9531), .S(n5648), .Z(n5624)
         );
  NAND2_X1 U6581 ( .A1(n5623), .A2(n5624), .ZN(n5622) );
  NAND2_X1 U6582 ( .A1(n5648), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5126) );
  NAND2_X1 U6583 ( .A1(n5622), .A2(n5126), .ZN(n5334) );
  INV_X1 U6584 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n5127) );
  XNOR2_X1 U6585 ( .A(n5768), .B(n5127), .ZN(n5335) );
  NAND2_X1 U6586 ( .A1(n5768), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5128) );
  INV_X1 U6587 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9533) );
  MUX2_X1 U6588 ( .A(n9533), .B(P1_REG1_REG_4__SCAN_IN), .S(n7202), .Z(n5614)
         );
  OAI21_X1 U6589 ( .B1(n7202), .B2(P1_REG1_REG_4__SCAN_IN), .A(n5129), .ZN(
        n5164) );
  XNOR2_X1 U6590 ( .A(n5994), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n5165) );
  AOI21_X1 U6591 ( .B1(n5131), .B2(n5130), .A(n5172), .ZN(n5133) );
  NOR2_X1 U6592 ( .A1(n5607), .A2(P1_U3084), .ZN(n7005) );
  AND2_X1 U6593 ( .A1(n7005), .A2(n5603), .ZN(n5132) );
  NAND2_X1 U6594 ( .A1(n5145), .A2(n5132), .ZN(n8855) );
  NOR2_X1 U6595 ( .A1(n5133), .A2(n8855), .ZN(n5134) );
  AOI211_X1 U6596 ( .C1(n9413), .C2(n6145), .A(n6554), .B(n5134), .ZN(n5143)
         );
  INV_X1 U6597 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n5135) );
  MUX2_X1 U6598 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n5135), .S(n6145), .Z(n5141)
         );
  XNOR2_X1 U6599 ( .A(n5464), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n5364) );
  NAND2_X1 U6600 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n5605) );
  NOR2_X1 U6601 ( .A1(n5364), .A2(n5605), .ZN(n5363) );
  AOI21_X1 U6602 ( .B1(n5464), .B2(P1_REG2_REG_1__SCAN_IN), .A(n5363), .ZN(
        n5628) );
  INV_X1 U6603 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5136) );
  MUX2_X1 U6604 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n5136), .S(n5648), .Z(n5137)
         );
  INV_X1 U6605 ( .A(n5137), .ZN(n5627) );
  NOR2_X1 U6606 ( .A1(n5628), .A2(n5627), .ZN(n5626) );
  AOI21_X1 U6607 ( .B1(n5648), .B2(P1_REG2_REG_2__SCAN_IN), .A(n5626), .ZN(
        n5340) );
  XNOR2_X1 U6608 ( .A(n5768), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n5339) );
  NOR2_X1 U6609 ( .A1(n5340), .A2(n5339), .ZN(n5338) );
  AOI21_X1 U6610 ( .B1(n5768), .B2(P1_REG2_REG_3__SCAN_IN), .A(n5338), .ZN(
        n5611) );
  MUX2_X1 U6611 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n4534), .S(n7202), .Z(n5610)
         );
  NAND2_X1 U6612 ( .A1(n5611), .A2(n5610), .ZN(n5609) );
  XNOR2_X1 U6613 ( .A(n5139), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n5162) );
  INV_X1 U6614 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5138) );
  NOR2_X1 U6615 ( .A1(n8878), .A2(n5607), .ZN(n9422) );
  OAI211_X1 U6616 ( .C1(n5141), .C2(n5140), .A(n4532), .B(n9422), .ZN(n5142)
         );
  OAI211_X1 U6617 ( .C1(n5144), .C2(n9426), .A(n5143), .B(n5142), .ZN(P1_U3247) );
  INV_X1 U6618 ( .A(n9426), .ZN(n8864) );
  INV_X1 U6619 ( .A(n5145), .ZN(n5153) );
  INV_X1 U6620 ( .A(n5607), .ZN(n8724) );
  INV_X1 U6621 ( .A(n5603), .ZN(n8885) );
  INV_X1 U6622 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5146) );
  NAND2_X1 U6623 ( .A1(n8885), .A2(n5146), .ZN(n5147) );
  NAND2_X1 U6624 ( .A1(n8724), .A2(n5147), .ZN(n5151) );
  NAND2_X1 U6625 ( .A1(n5151), .A2(n5420), .ZN(n5606) );
  NAND2_X1 U6626 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_STATE_REG_SCAN_IN), 
        .ZN(n5149) );
  INV_X1 U6627 ( .A(n6925), .ZN(n5148) );
  OAI21_X1 U6628 ( .B1(n5607), .B2(n5149), .A(n5148), .ZN(n5150) );
  OAI211_X1 U6629 ( .C1(n5151), .C2(n5420), .A(n5606), .B(n5150), .ZN(n5152)
         );
  INV_X1 U6630 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9435) );
  OAI22_X1 U6631 ( .A1(n5153), .A2(n5152), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9435), .ZN(n5155) );
  NOR3_X1 U6632 ( .A1(n8855), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n5420), .ZN(
        n5154) );
  AOI211_X1 U6633 ( .C1(P1_ADDR_REG_0__SCAN_IN), .C2(n8864), .A(n5155), .B(
        n5154), .ZN(n5156) );
  INV_X1 U6634 ( .A(n5156), .ZN(P1_U3241) );
  NAND2_X1 U6635 ( .A1(n5157), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5158) );
  XNOR2_X1 U6636 ( .A(n5158), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9412) );
  INV_X1 U6637 ( .A(n9412), .ZN(n6858) );
  OAI222_X1 U6638 ( .A1(n9275), .A2(n5160), .B1(n6728), .B2(n5159), .C1(n6858), 
        .C2(P1_U3084), .ZN(P1_U3339) );
  INV_X1 U6639 ( .A(n9422), .ZN(n8861) );
  XOR2_X1 U6640 ( .A(n5162), .B(n5161), .Z(n5169) );
  AND2_X1 U6641 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6037) );
  AOI211_X1 U6642 ( .C1(n5165), .C2(n5164), .A(n5163), .B(n8855), .ZN(n5166)
         );
  AOI211_X1 U6643 ( .C1(n9413), .C2(n5994), .A(n6037), .B(n5166), .ZN(n5168)
         );
  NAND2_X1 U6644 ( .A1(n8864), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n5167) );
  OAI211_X1 U6645 ( .C1(n8861), .C2(n5169), .A(n5168), .B(n5167), .ZN(P1_U3246) );
  INV_X1 U6646 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n5181) );
  INV_X1 U6647 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n5170) );
  MUX2_X1 U6648 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n5170), .S(n6318), .Z(n5171)
         );
  NAND2_X1 U6649 ( .A1(n4298), .A2(n5171), .ZN(n5287) );
  OAI21_X1 U6650 ( .B1(n4298), .B2(n5171), .A(n5287), .ZN(n5179) );
  INV_X1 U6651 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9539) );
  MUX2_X1 U6652 ( .A(n9539), .B(P1_REG1_REG_7__SCAN_IN), .S(n6318), .Z(n5175)
         );
  AOI21_X1 U6653 ( .B1(n5173), .B2(n9537), .A(n5172), .ZN(n5174) );
  NOR2_X1 U6654 ( .A1(n5174), .A2(n5175), .ZN(n5280) );
  AOI21_X1 U6655 ( .B1(n5175), .B2(n5174), .A(n5280), .ZN(n5177) );
  NAND2_X1 U6656 ( .A1(n9413), .A2(n6318), .ZN(n5176) );
  NAND2_X1 U6657 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n8383) );
  OAI211_X1 U6658 ( .C1(n5177), .C2(n8855), .A(n5176), .B(n8383), .ZN(n5178)
         );
  AOI21_X1 U6659 ( .B1(n9422), .B2(n5179), .A(n5178), .ZN(n5180) );
  OAI21_X1 U6660 ( .B1(n9426), .B2(n5181), .A(n5180), .ZN(P1_U3248) );
  OAI21_X1 U6661 ( .B1(n5736), .B2(P2_U3152), .A(n7438), .ZN(n5182) );
  INV_X1 U6662 ( .A(n5182), .ZN(n5183) );
  OAI21_X1 U6663 ( .B1(n9631), .B2(n5546), .A(n5183), .ZN(n5188) );
  NAND2_X1 U6664 ( .A1(n5188), .A2(n6976), .ZN(n5184) );
  NAND2_X1 U6665 ( .A1(n5184), .A2(n7982), .ZN(n5202) );
  AND2_X1 U6666 ( .A1(n5202), .A2(n5185), .ZN(n9295) );
  INV_X1 U6667 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6666) );
  AND2_X1 U6668 ( .A1(n6976), .A2(n5186), .ZN(n5187) );
  INV_X1 U6669 ( .A(n5668), .ZN(n9294) );
  INV_X1 U6670 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9581) );
  INV_X1 U6671 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9727) );
  XNOR2_X1 U6672 ( .A(n9282), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n9285) );
  NOR3_X1 U6673 ( .A1(n9581), .A2(n9727), .A3(n9285), .ZN(n9283) );
  AND2_X1 U6674 ( .A1(n9282), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5189) );
  NOR2_X1 U6675 ( .A1(n9283), .A2(n5189), .ZN(n9302) );
  INV_X1 U6676 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n5190) );
  MUX2_X1 U6677 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n5190), .S(n5668), .Z(n9301)
         );
  NOR2_X1 U6678 ( .A1(n9302), .A2(n9301), .ZN(n9300) );
  AOI21_X1 U6679 ( .B1(n9294), .B2(P2_REG1_REG_2__SCAN_IN), .A(n9300), .ZN(
        n5194) );
  OR2_X1 U6680 ( .A1(n5220), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5192) );
  NAND2_X1 U6681 ( .A1(n5220), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5191) );
  NAND2_X1 U6682 ( .A1(n5192), .A2(n5191), .ZN(n5193) );
  NOR2_X1 U6683 ( .A1(n5194), .A2(n5193), .ZN(n5208) );
  AOI21_X1 U6684 ( .B1(n5194), .B2(n5193), .A(n5208), .ZN(n5195) );
  NAND2_X1 U6685 ( .A1(n9573), .A2(n5195), .ZN(n5197) );
  NAND2_X1 U6686 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3152), .ZN(n5196) );
  OAI211_X1 U6687 ( .C1(n8072), .C2(n6666), .A(n5197), .B(n5196), .ZN(n5206)
         );
  OR2_X1 U6688 ( .A1(n9282), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5199) );
  NAND2_X1 U6689 ( .A1(n9282), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5198) );
  NAND2_X1 U6690 ( .A1(n5199), .A2(n5198), .ZN(n9278) );
  NOR3_X1 U6691 ( .A1(n9581), .A2(n5088), .A3(n9278), .ZN(n9279) );
  AOI21_X1 U6692 ( .B1(n9282), .B2(P2_REG2_REG_1__SCAN_IN), .A(n9279), .ZN(
        n9296) );
  INV_X1 U6693 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6140) );
  MUX2_X1 U6694 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n6140), .S(n5668), .Z(n9297)
         );
  NOR2_X1 U6695 ( .A1(n9296), .A2(n9297), .ZN(n9299) );
  AOI21_X1 U6696 ( .B1(n9294), .B2(P2_REG2_REG_2__SCAN_IN), .A(n9299), .ZN(
        n5204) );
  NAND2_X1 U6697 ( .A1(n5220), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5200) );
  OAI21_X1 U6698 ( .B1(n5220), .B2(P2_REG2_REG_3__SCAN_IN), .A(n5200), .ZN(
        n5203) );
  NOR2_X1 U6699 ( .A1(n5204), .A2(n5203), .ZN(n5219) );
  NOR2_X1 U6700 ( .A1(n5185), .A2(n5186), .ZN(n5201) );
  NAND2_X1 U6701 ( .A1(n5202), .A2(n5201), .ZN(n9576) );
  AOI211_X1 U6702 ( .C1(n5204), .C2(n5203), .A(n5219), .B(n9576), .ZN(n5205)
         );
  AOI211_X1 U6703 ( .C1(n9295), .C2(n5220), .A(n5206), .B(n5205), .ZN(n5207)
         );
  INV_X1 U6704 ( .A(n5207), .ZN(P2_U3248) );
  INV_X1 U6705 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n5218) );
  INV_X1 U6706 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5945) );
  MUX2_X1 U6707 ( .A(n5945), .B(P2_REG1_REG_8__SCAN_IN), .S(n5942), .Z(n5214)
         );
  XNOR2_X1 U6708 ( .A(n5722), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n5259) );
  INV_X1 U6709 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n5210) );
  AOI21_X1 U6710 ( .B1(n5220), .B2(P2_REG1_REG_3__SCAN_IN), .A(n5208), .ZN(
        n5244) );
  MUX2_X1 U6711 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n5210), .S(n5695), .Z(n5245)
         );
  NOR2_X1 U6712 ( .A1(n5244), .A2(n5245), .ZN(n5243) );
  INV_X1 U6713 ( .A(n5243), .ZN(n5209) );
  OAI21_X1 U6714 ( .B1(n5695), .B2(n5210), .A(n5209), .ZN(n5258) );
  NAND2_X1 U6715 ( .A1(n5259), .A2(n5258), .ZN(n5257) );
  INV_X1 U6716 ( .A(n5722), .ZN(n5267) );
  NAND2_X1 U6717 ( .A1(n5267), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5211) );
  NAND2_X1 U6718 ( .A1(n5257), .A2(n5211), .ZN(n5270) );
  INV_X1 U6719 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9735) );
  MUX2_X1 U6720 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n9735), .S(n5796), .Z(n5271)
         );
  NAND2_X1 U6721 ( .A1(n5270), .A2(n5271), .ZN(n5269) );
  NAND2_X1 U6722 ( .A1(n5796), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5212) );
  AND2_X1 U6723 ( .A1(n5269), .A2(n5212), .ZN(n5232) );
  INV_X1 U6724 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n5804) );
  MUX2_X1 U6725 ( .A(n5804), .B(P2_REG1_REG_7__SCAN_IN), .S(n5936), .Z(n5231)
         );
  NOR2_X1 U6726 ( .A1(n5232), .A2(n5231), .ZN(n5230) );
  AOI21_X1 U6727 ( .B1(n5936), .B2(P2_REG1_REG_7__SCAN_IN), .A(n5230), .ZN(
        n5213) );
  NOR2_X1 U6728 ( .A1(n5213), .A2(n5214), .ZN(n5320) );
  AOI21_X1 U6729 ( .B1(n5214), .B2(n5213), .A(n5320), .ZN(n5215) );
  NAND2_X1 U6730 ( .A1(n9573), .A2(n5215), .ZN(n5217) );
  NAND2_X1 U6731 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n5216) );
  OAI211_X1 U6732 ( .C1(n8072), .C2(n5218), .A(n5217), .B(n5216), .ZN(n5228)
         );
  INV_X1 U6733 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5711) );
  XOR2_X1 U6734 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n5722), .Z(n5263) );
  INV_X1 U6735 ( .A(n5695), .ZN(n5255) );
  AOI21_X1 U6736 ( .B1(n5220), .B2(P2_REG2_REG_3__SCAN_IN), .A(n5219), .ZN(
        n5252) );
  INV_X1 U6737 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5702) );
  MUX2_X1 U6738 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n5702), .S(n5695), .Z(n5251)
         );
  NOR2_X1 U6739 ( .A1(n5252), .A2(n5251), .ZN(n5250) );
  AOI21_X1 U6740 ( .B1(n5255), .B2(P2_REG2_REG_4__SCAN_IN), .A(n5250), .ZN(
        n5264) );
  NOR2_X1 U6741 ( .A1(n5263), .A2(n5264), .ZN(n5262) );
  INV_X1 U6742 ( .A(n5262), .ZN(n5221) );
  OAI21_X1 U6743 ( .B1(n5711), .B2(n5722), .A(n5221), .ZN(n5276) );
  INV_X1 U6744 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n5222) );
  MUX2_X1 U6745 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n5222), .S(n5796), .Z(n5277)
         );
  INV_X1 U6746 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n5223) );
  MUX2_X1 U6747 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n5223), .S(n5936), .Z(n5224)
         );
  INV_X1 U6748 ( .A(n5224), .ZN(n5238) );
  AOI21_X1 U6749 ( .B1(n5936), .B2(P2_REG2_REG_7__SCAN_IN), .A(n5237), .ZN(
        n5226) );
  INV_X1 U6750 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n5946) );
  MUX2_X1 U6751 ( .A(n5946), .B(P2_REG2_REG_8__SCAN_IN), .S(n5942), .Z(n5225)
         );
  AOI211_X1 U6752 ( .C1(n5226), .C2(n5225), .A(n5326), .B(n9576), .ZN(n5227)
         );
  AOI211_X1 U6753 ( .C1(n9295), .C2(n5942), .A(n5228), .B(n5227), .ZN(n5229)
         );
  INV_X1 U6754 ( .A(n5229), .ZN(P2_U3253) );
  INV_X1 U6755 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n5236) );
  AOI21_X1 U6756 ( .B1(n5232), .B2(n5231), .A(n5230), .ZN(n5233) );
  NAND2_X1 U6757 ( .A1(n9573), .A2(n5233), .ZN(n5235) );
  NAND2_X1 U6758 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3152), .ZN(n5234) );
  OAI211_X1 U6759 ( .C1(n8072), .C2(n5236), .A(n5235), .B(n5234), .ZN(n5241)
         );
  AOI211_X1 U6760 ( .C1(n5239), .C2(n5238), .A(n5237), .B(n9576), .ZN(n5240)
         );
  AOI211_X1 U6761 ( .C1(n9295), .C2(n5936), .A(n5241), .B(n5240), .ZN(n5242)
         );
  INV_X1 U6762 ( .A(n5242), .ZN(P2_U3252) );
  INV_X1 U6763 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n5249) );
  AOI21_X1 U6764 ( .B1(n5245), .B2(n5244), .A(n5243), .ZN(n5246) );
  NAND2_X1 U6765 ( .A1(n9573), .A2(n5246), .ZN(n5248) );
  NAND2_X1 U6766 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n5247) );
  OAI211_X1 U6767 ( .C1(n8072), .C2(n5249), .A(n5248), .B(n5247), .ZN(n5254)
         );
  AOI211_X1 U6768 ( .C1(n5252), .C2(n5251), .A(n5250), .B(n9576), .ZN(n5253)
         );
  AOI211_X1 U6769 ( .C1(n9295), .C2(n5255), .A(n5254), .B(n5253), .ZN(n5256)
         );
  INV_X1 U6770 ( .A(n5256), .ZN(P2_U3249) );
  INV_X1 U6771 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n5261) );
  OAI211_X1 U6772 ( .C1(n5259), .C2(n5258), .A(n9573), .B(n5257), .ZN(n5260)
         );
  NAND2_X1 U6773 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3152), .ZN(n5739) );
  OAI211_X1 U6774 ( .C1(n8072), .C2(n5261), .A(n5260), .B(n5739), .ZN(n5266)
         );
  AOI211_X1 U6775 ( .C1(n5264), .C2(n5263), .A(n5262), .B(n9576), .ZN(n5265)
         );
  AOI211_X1 U6776 ( .C1(n9295), .C2(n5267), .A(n5266), .B(n5265), .ZN(n5268)
         );
  INV_X1 U6777 ( .A(n5268), .ZN(P2_U3250) );
  INV_X1 U6778 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n5273) );
  OAI211_X1 U6779 ( .C1(n5271), .C2(n5270), .A(n9573), .B(n5269), .ZN(n5272)
         );
  NAND2_X1 U6780 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n5813) );
  OAI211_X1 U6781 ( .C1(n8072), .C2(n5273), .A(n5272), .B(n5813), .ZN(n5274)
         );
  AOI21_X1 U6782 ( .B1(n5796), .B2(n9295), .A(n5274), .ZN(n5279) );
  INV_X1 U6783 ( .A(n9576), .ZN(n9572) );
  OAI211_X1 U6784 ( .C1(n5277), .C2(n5276), .A(n9572), .B(n5275), .ZN(n5278)
         );
  NAND2_X1 U6785 ( .A1(n5279), .A2(n5278), .ZN(P2_U3251) );
  INV_X1 U6786 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9542) );
  MUX2_X1 U6787 ( .A(n9542), .B(P1_REG1_REG_8__SCAN_IN), .S(n6331), .Z(n5283)
         );
  AOI21_X1 U6788 ( .B1(n5281), .B2(n9539), .A(n5280), .ZN(n5282) );
  AOI21_X1 U6789 ( .B1(n5283), .B2(n5282), .A(n5345), .ZN(n5293) );
  NAND2_X1 U6790 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6446) );
  OAI21_X1 U6791 ( .B1(n4363), .B2(n5284), .A(n6446), .ZN(n5285) );
  AOI21_X1 U6792 ( .B1(n8864), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n5285), .ZN(
        n5292) );
  INV_X1 U6793 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5286) );
  MUX2_X1 U6794 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n5286), .S(n6331), .Z(n5289)
         );
  OAI21_X1 U6795 ( .B1(n6318), .B2(P1_REG2_REG_7__SCAN_IN), .A(n5287), .ZN(
        n5288) );
  NAND2_X1 U6796 ( .A1(n5288), .A2(n5289), .ZN(n5351) );
  OAI21_X1 U6797 ( .B1(n5289), .B2(n5288), .A(n5351), .ZN(n5290) );
  NAND2_X1 U6798 ( .A1(n5290), .A2(n9422), .ZN(n5291) );
  OAI211_X1 U6799 ( .C1(n5293), .C2(n8855), .A(n5292), .B(n5291), .ZN(P1_U3249) );
  INV_X1 U6800 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n9871) );
  INV_X1 U6801 ( .A(n5295), .ZN(n5296) );
  NAND2_X1 U6802 ( .A1(n5296), .A2(SI_14_), .ZN(n5297) );
  INV_X1 U6803 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6975) );
  MUX2_X1 U6804 ( .A(n6975), .B(n9871), .S(n7244), .Z(n5301) );
  INV_X1 U6805 ( .A(SI_15_), .ZN(n5300) );
  INV_X1 U6806 ( .A(n5301), .ZN(n5302) );
  NAND2_X1 U6807 ( .A1(n5302), .A2(SI_15_), .ZN(n5303) );
  NAND2_X1 U6808 ( .A1(n5430), .A2(n5303), .ZN(n5431) );
  XNOR2_X1 U6809 ( .A(n5432), .B(n5431), .ZN(n6974) );
  INV_X1 U6810 ( .A(n6974), .ZN(n5317) );
  NOR2_X1 U6811 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5304) );
  AND2_X1 U6812 ( .A1(n5305), .A2(n5304), .ZN(n5310) );
  NOR2_X1 U6813 ( .A1(n5310), .A2(n5306), .ZN(n5307) );
  MUX2_X1 U6814 ( .A(n5306), .B(n5307), .S(P1_IR_REG_15__SCAN_IN), .Z(n5308)
         );
  INV_X1 U6815 ( .A(n5308), .ZN(n5311) );
  NAND2_X1 U6816 ( .A1(n5310), .A2(n5309), .ZN(n5502) );
  NAND2_X1 U6817 ( .A1(n5311), .A2(n5502), .ZN(n7014) );
  OAI222_X1 U6818 ( .A1(n9275), .A2(n9871), .B1(n6728), .B2(n5317), .C1(
        P1_U3084), .C2(n7014), .ZN(P1_U3338) );
  INV_X1 U6819 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5312) );
  NAND2_X1 U6820 ( .A1(n5313), .A2(n5312), .ZN(n5314) );
  NAND2_X1 U6821 ( .A1(n5314), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5316) );
  INV_X1 U6822 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5315) );
  XNOR2_X1 U6823 ( .A(n5316), .B(n5315), .ZN(n8019) );
  INV_X1 U6824 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n6686) );
  OR2_X1 U6825 ( .A1(n5908), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5319) );
  NAND2_X1 U6826 ( .A1(n5908), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5318) );
  NAND2_X1 U6827 ( .A1(n5319), .A2(n5318), .ZN(n5322) );
  AOI21_X1 U6828 ( .B1(n5942), .B2(P2_REG1_REG_8__SCAN_IN), .A(n5320), .ZN(
        n5321) );
  NOR2_X1 U6829 ( .A1(n5321), .A2(n5322), .ZN(n5589) );
  AOI21_X1 U6830 ( .B1(n5322), .B2(n5321), .A(n5589), .ZN(n5323) );
  NAND2_X1 U6831 ( .A1(n9573), .A2(n5323), .ZN(n5325) );
  NAND2_X1 U6832 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n5324) );
  OAI211_X1 U6833 ( .C1(n8072), .C2(n6686), .A(n5325), .B(n5324), .ZN(n5331)
         );
  NAND2_X1 U6834 ( .A1(n5908), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5327) );
  OAI21_X1 U6835 ( .B1(n5908), .B2(P2_REG2_REG_9__SCAN_IN), .A(n5327), .ZN(
        n5328) );
  AOI211_X1 U6836 ( .C1(n5329), .C2(n5328), .A(n5596), .B(n9576), .ZN(n5330)
         );
  AOI211_X1 U6837 ( .C1(n9295), .C2(n5908), .A(n5331), .B(n5330), .ZN(n5332)
         );
  INV_X1 U6838 ( .A(n5332), .ZN(P2_U3254) );
  NAND2_X1 U6839 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3084), .ZN(n5783) );
  INV_X1 U6840 ( .A(n8855), .ZN(n9421) );
  OAI211_X1 U6841 ( .C1(n5335), .C2(n5334), .A(n9421), .B(n5333), .ZN(n5336)
         );
  OAI211_X1 U6842 ( .C1(n4363), .C2(n5337), .A(n5783), .B(n5336), .ZN(n5342)
         );
  AOI211_X1 U6843 ( .C1(n5340), .C2(n5339), .A(n5338), .B(n8861), .ZN(n5341)
         );
  AOI211_X1 U6844 ( .C1(P1_ADDR_REG_3__SCAN_IN), .C2(n8864), .A(n5342), .B(
        n5341), .ZN(n5343) );
  INV_X1 U6845 ( .A(n5343), .ZN(P1_U3244) );
  INV_X1 U6846 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5344) );
  MUX2_X1 U6847 ( .A(n5344), .B(P1_REG1_REG_9__SCAN_IN), .S(n5348), .Z(n5347)
         );
  OAI21_X1 U6848 ( .B1(n5347), .B2(n5346), .A(n5511), .ZN(n5357) );
  INV_X1 U6849 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n5350) );
  AND2_X1 U6850 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n6537) );
  AOI21_X1 U6851 ( .B1(n9413), .B2(n6348), .A(n6537), .ZN(n5349) );
  OAI21_X1 U6852 ( .B1(n9426), .B2(n5350), .A(n5349), .ZN(n5356) );
  OAI21_X1 U6853 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n6331), .A(n5351), .ZN(
        n5354) );
  NAND2_X1 U6854 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(n6348), .ZN(n5352) );
  OAI21_X1 U6855 ( .B1(n6348), .B2(P1_REG2_REG_9__SCAN_IN), .A(n5352), .ZN(
        n5353) );
  NOR2_X1 U6856 ( .A1(n5354), .A2(n5353), .ZN(n5516) );
  AOI211_X1 U6857 ( .C1(n5354), .C2(n5353), .A(n8861), .B(n5516), .ZN(n5355)
         );
  AOI211_X1 U6858 ( .C1(n9421), .C2(n5357), .A(n5356), .B(n5355), .ZN(n5358)
         );
  INV_X1 U6859 ( .A(n5358), .ZN(P1_U3250) );
  INV_X1 U6860 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n5368) );
  INV_X1 U6861 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6106) );
  OAI211_X1 U6862 ( .C1(n5361), .C2(n5360), .A(n9421), .B(n5359), .ZN(n5362)
         );
  OAI21_X1 U6863 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6106), .A(n5362), .ZN(n5366) );
  AOI211_X1 U6864 ( .C1(n5605), .C2(n5364), .A(n5363), .B(n8861), .ZN(n5365)
         );
  AOI211_X1 U6865 ( .C1(n9413), .C2(n5464), .A(n5366), .B(n5365), .ZN(n5367)
         );
  OAI21_X1 U6866 ( .B1(n9426), .B2(n5368), .A(n5367), .ZN(P1_U3242) );
  NAND2_X1 U6867 ( .A1(n6726), .A2(P1_B_REG_SCAN_IN), .ZN(n5369) );
  MUX2_X1 U6868 ( .A(n5369), .B(P1_B_REG_SCAN_IN), .S(n4881), .Z(n5372) );
  INV_X1 U6869 ( .A(n5370), .ZN(n5371) );
  INV_X1 U6870 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9469) );
  NAND2_X1 U6871 ( .A1(n9262), .A2(n9469), .ZN(n5374) );
  NAND2_X1 U6872 ( .A1(n5370), .A2(n6726), .ZN(n5373) );
  NAND2_X1 U6873 ( .A1(n5374), .A2(n5373), .ZN(n5444) );
  INV_X1 U6874 ( .A(n5444), .ZN(n5385) );
  NOR4_X1 U6875 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5378) );
  NOR4_X1 U6876 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n5377) );
  NOR4_X1 U6877 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5376) );
  NOR4_X1 U6878 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n5375) );
  NAND4_X1 U6879 ( .A1(n5378), .A2(n5377), .A3(n5376), .A4(n5375), .ZN(n5384)
         );
  NOR2_X1 U6880 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .ZN(
        n5382) );
  NOR4_X1 U6881 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n5381) );
  NOR4_X1 U6882 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n5380) );
  NOR4_X1 U6883 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n5379) );
  NAND4_X1 U6884 ( .A1(n5382), .A2(n5381), .A3(n5380), .A4(n5379), .ZN(n5383)
         );
  OAI21_X1 U6885 ( .B1(n5384), .B2(n5383), .A(n9262), .ZN(n5445) );
  NAND2_X1 U6886 ( .A1(n5385), .A2(n5445), .ZN(n5397) );
  INV_X1 U6887 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5386) );
  NAND2_X1 U6888 ( .A1(n9262), .A2(n5386), .ZN(n5387) );
  NAND2_X1 U6889 ( .A1(n5370), .A2(n6592), .ZN(n9263) );
  NAND2_X1 U6890 ( .A1(n5389), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5390) );
  NAND2_X1 U6891 ( .A1(n5391), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5393) );
  INV_X1 U6892 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5392) );
  OAI21_X1 U6893 ( .B1(n5397), .B2(n6060), .A(n5446), .ZN(n5395) );
  AND2_X1 U6894 ( .A1(n8772), .A2(n9026), .ZN(n5398) );
  OR2_X1 U6895 ( .A1(n8720), .A2(n5398), .ZN(n6059) );
  AND3_X1 U6896 ( .A1(n6059), .A2(n5415), .A3(n6506), .ZN(n5394) );
  NAND2_X1 U6897 ( .A1(n5395), .A2(n5394), .ZN(n5782) );
  NOR2_X1 U6898 ( .A1(n5782), .A2(P1_U3084), .ZN(n5659) );
  AND2_X1 U6899 ( .A1(n6506), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5396) );
  NAND2_X1 U6900 ( .A1(n5415), .A2(n5396), .ZN(n9470) );
  NOR2_X1 U6901 ( .A1(n5397), .A2(n9470), .ZN(n6393) );
  NAND2_X1 U6902 ( .A1(n6393), .A2(n6391), .ZN(n5427) );
  INV_X1 U6903 ( .A(n5398), .ZN(n8716) );
  OR2_X1 U6904 ( .A1(n5427), .A2(n8716), .ZN(n8511) );
  INV_X1 U6905 ( .A(n8720), .ZN(n5425) );
  INV_X1 U6906 ( .A(n8487), .ZN(n8503) );
  NAND2_X1 U6907 ( .A1(n4275), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5400) );
  NAND2_X1 U6908 ( .A1(n6341), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5409) );
  NAND2_X1 U6909 ( .A1(n5786), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5407) );
  AND2_X4 U6910 ( .A1(n9269), .A2(n5405), .ZN(n5785) );
  NAND2_X1 U6911 ( .A1(n5785), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5406) );
  NAND4_X2 U6912 ( .A1(n5409), .A2(n5408), .A3(n5407), .A4(n5406), .ZN(n5875)
         );
  NAND2_X1 U6913 ( .A1(n5496), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5413) );
  NAND2_X1 U6914 ( .A1(n6341), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5412) );
  NAND2_X1 U6915 ( .A1(n5786), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5411) );
  NAND2_X1 U6916 ( .A1(n5785), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5410) );
  INV_X1 U6917 ( .A(n6079), .ZN(n5416) );
  NAND2_X1 U6918 ( .A1(n7244), .A2(SI_0_), .ZN(n5417) );
  XNOR2_X1 U6919 ( .A(n5417), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9276) );
  NAND2_X1 U6920 ( .A1(n7497), .A2(n5887), .ZN(n5419) );
  OAI21_X1 U6921 ( .B1(n5415), .B2(n5420), .A(n5419), .ZN(n5421) );
  INV_X1 U6922 ( .A(n5415), .ZN(n5422) );
  AOI22_X1 U6923 ( .A1(n5887), .A2(n4262), .B1(P1_REG1_REG_0__SCAN_IN), .B2(
        n5422), .ZN(n5423) );
  NAND2_X1 U6924 ( .A1(n5424), .A2(n5423), .ZN(n5455) );
  OAI21_X1 U6925 ( .B1(n4346), .B2(n5455), .A(n5459), .ZN(n5604) );
  INV_X1 U6926 ( .A(n5452), .ZN(n5450) );
  NAND2_X1 U6927 ( .A1(n5450), .A2(n8716), .ZN(n9517) );
  INV_X2 U6928 ( .A(n9517), .ZN(n9216) );
  AOI22_X1 U6929 ( .A1(n8503), .A2(n5875), .B1(n5604), .B2(n8496), .ZN(n5429)
         );
  OR2_X1 U6930 ( .A1(n5452), .A2(n8772), .ZN(n6064) );
  INV_X1 U6931 ( .A(n5446), .ZN(n5426) );
  INV_X1 U6932 ( .A(n9470), .ZN(n8723) );
  OAI21_X2 U6933 ( .B1(n5427), .B2(n6064), .A(n9436), .ZN(n8490) );
  NAND2_X1 U6934 ( .A1(n8490), .A2(n5887), .ZN(n5428) );
  OAI211_X1 U6935 ( .C1(n5659), .C2(n9435), .A(n5429), .B(n5428), .ZN(P1_U3230) );
  INV_X1 U6936 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5440) );
  INV_X1 U6937 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5443) );
  MUX2_X1 U6938 ( .A(n5440), .B(n5443), .S(n7244), .Z(n5434) );
  INV_X1 U6939 ( .A(SI_16_), .ZN(n5433) );
  NAND2_X1 U6940 ( .A1(n5434), .A2(n5433), .ZN(n5487) );
  INV_X1 U6941 ( .A(n5434), .ZN(n5435) );
  NAND2_X1 U6942 ( .A1(n5435), .A2(SI_16_), .ZN(n5436) );
  XNOR2_X1 U6943 ( .A(n5486), .B(n5485), .ZN(n7510) );
  INV_X1 U6944 ( .A(n7510), .ZN(n5442) );
  NOR2_X1 U6945 ( .A1(n4840), .A2(n5539), .ZN(n5437) );
  MUX2_X1 U6946 ( .A(n5539), .B(n5437), .S(P2_IR_REG_16__SCAN_IN), .Z(n5438)
         );
  INV_X1 U6947 ( .A(n5438), .ZN(n5439) );
  AND2_X1 U6948 ( .A1(n5439), .A2(n5491), .ZN(n8034) );
  INV_X1 U6949 ( .A(n8034), .ZN(n8017) );
  OAI222_X1 U6950 ( .A1(n4268), .A2(n5442), .B1(n8017), .B2(P2_U3152), .C1(
        n5440), .C2(n8371), .ZN(P2_U3342) );
  NAND2_X1 U6951 ( .A1(n5502), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5441) );
  XNOR2_X1 U6952 ( .A(n5441), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8844) );
  INV_X1 U6953 ( .A(n8844), .ZN(n7017) );
  OAI222_X1 U6954 ( .A1(n9275), .A2(n5443), .B1(n9273), .B2(n5442), .C1(n7017), 
        .C2(P1_U3084), .ZN(P1_U3337) );
  AND2_X1 U6955 ( .A1(n5444), .A2(n8723), .ZN(n9468) );
  AND2_X1 U6956 ( .A1(n5445), .A2(n6059), .ZN(n5447) );
  AND2_X2 U6957 ( .A1(n5891), .A2(n6060), .ZN(n9528) );
  INV_X1 U6958 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5454) );
  NAND2_X1 U6959 ( .A1(n8823), .A2(n9427), .ZN(n8652) );
  INV_X1 U6960 ( .A(n8652), .ZN(n5448) );
  NOR2_X1 U6961 ( .A1(n6096), .A2(n5448), .ZN(n8734) );
  NAND2_X1 U6962 ( .A1(n5449), .A2(n9026), .ZN(n5456) );
  OR2_X1 U6963 ( .A1(n5456), .A2(n6079), .ZN(n5883) );
  INV_X1 U6964 ( .A(n5883), .ZN(n8725) );
  NOR3_X1 U6965 ( .A1(n8734), .A2(n8725), .A3(n5450), .ZN(n5451) );
  AOI21_X1 U6966 ( .B1(n9114), .B2(n5875), .A(n5451), .ZN(n9430) );
  OAI21_X1 U6967 ( .B1(n9427), .B2(n5452), .A(n9430), .ZN(n9241) );
  NAND2_X1 U6968 ( .A1(n9241), .A2(n9528), .ZN(n5453) );
  OAI21_X1 U6969 ( .B1(n9528), .B2(n5454), .A(n5453), .ZN(P1_U3454) );
  INV_X1 U6970 ( .A(n5455), .ZN(n5457) );
  NAND2_X1 U6971 ( .A1(n5457), .A2(n7675), .ZN(n5458) );
  NAND2_X1 U6972 ( .A1(n5875), .A2(n4265), .ZN(n5469) );
  NAND2_X1 U6973 ( .A1(n6329), .A2(n5460), .ZN(n5467) );
  INV_X1 U6974 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5462) );
  NAND2_X1 U6975 ( .A1(n7566), .A2(n5464), .ZN(n5465) );
  NAND2_X1 U6976 ( .A1(n5469), .A2(n5468), .ZN(n5470) );
  INV_X1 U6977 ( .A(n5473), .ZN(n5471) );
  NAND2_X1 U6978 ( .A1(n5472), .A2(n5471), .ZN(n5646) );
  NAND2_X1 U6979 ( .A1(n5474), .A2(n5473), .ZN(n5645) );
  NAND2_X1 U6980 ( .A1(n5646), .A2(n5645), .ZN(n5477) );
  NAND2_X1 U6981 ( .A1(n5875), .A2(n6703), .ZN(n5476) );
  OR2_X1 U6982 ( .A1(n8650), .A2(n7678), .ZN(n5475) );
  AND2_X1 U6983 ( .A1(n5476), .A2(n5475), .ZN(n5644) );
  XNOR2_X1 U6984 ( .A(n5477), .B(n5644), .ZN(n5484) );
  OR2_X1 U6985 ( .A1(n8720), .A2(n5607), .ZN(n9060) );
  NAND2_X1 U6986 ( .A1(n6341), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5481) );
  NAND2_X1 U6987 ( .A1(n5786), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5479) );
  NAND2_X1 U6988 ( .A1(n5785), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5478) );
  AOI22_X1 U6989 ( .A1(n9112), .A2(n8823), .B1(n8822), .B2(n9114), .ZN(n6101)
         );
  OAI22_X1 U6990 ( .A1(n5659), .A2(n6106), .B1(n8511), .B2(n6101), .ZN(n5482)
         );
  AOI21_X1 U6991 ( .B1(n9473), .B2(n8490), .A(n5482), .ZN(n5483) );
  OAI21_X1 U6992 ( .B1(n5484), .B2(n8519), .A(n5483), .ZN(P1_U3220) );
  NAND2_X1 U6993 ( .A1(n5488), .A2(n5487), .ZN(n5761) );
  INV_X1 U6994 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n5489) );
  INV_X1 U6995 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5509) );
  MUX2_X1 U6996 ( .A(n5489), .B(n5509), .S(n7244), .Z(n5757) );
  XNOR2_X1 U6997 ( .A(n5757), .B(SI_17_), .ZN(n5756) );
  XNOR2_X1 U6998 ( .A(n5761), .B(n5756), .ZN(n7523) );
  INV_X1 U6999 ( .A(n7523), .ZN(n5508) );
  NAND2_X1 U7000 ( .A1(n5491), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5492) );
  MUX2_X1 U7001 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5492), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n5493) );
  AND2_X1 U7002 ( .A1(n5490), .A2(n5493), .ZN(n8050) );
  AOI22_X1 U7003 ( .A1(n8050), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n5494), .ZN(n5495) );
  OAI21_X1 U7004 ( .B1(n5508), .B2(n4268), .A(n5495), .ZN(P2_U3341) );
  INV_X1 U7005 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n5501) );
  NAND2_X1 U7006 ( .A1(n8615), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n5499) );
  NAND2_X1 U7007 ( .A1(n5785), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U7008 ( .A1(n7591), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n5497) );
  AND3_X1 U7009 ( .A1(n5499), .A2(n5498), .A3(n5497), .ZN(n8887) );
  INV_X1 U7010 ( .A(n8887), .ZN(n8620) );
  NAND2_X1 U7011 ( .A1(n8620), .A2(P1_U4006), .ZN(n5500) );
  OAI21_X1 U7012 ( .B1(P1_U4006), .B2(n5501), .A(n5500), .ZN(P1_U3586) );
  OR2_X1 U7013 ( .A1(n5502), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n5503) );
  NAND2_X1 U7014 ( .A1(n5503), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5506) );
  INV_X1 U7015 ( .A(n5506), .ZN(n5504) );
  NAND2_X1 U7016 ( .A1(n5504), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n5507) );
  NAND2_X1 U7017 ( .A1(n5506), .A2(n5505), .ZN(n5762) );
  INV_X1 U7018 ( .A(n8859), .ZN(n8839) );
  OAI222_X1 U7019 ( .A1(n9275), .A2(n5509), .B1(n9273), .B2(n5508), .C1(n8839), 
        .C2(P1_U3084), .ZN(P1_U3336) );
  INV_X1 U7020 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n5510) );
  AOI22_X1 U7021 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n6565), .B1(n5515), .B2(
        n5510), .ZN(n5513) );
  OAI21_X1 U7022 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n6348), .A(n5511), .ZN(
        n5512) );
  NAND2_X1 U7023 ( .A1(n5513), .A2(n5512), .ZN(n5841) );
  OAI21_X1 U7024 ( .B1(n5513), .B2(n5512), .A(n5841), .ZN(n5522) );
  NAND2_X1 U7025 ( .A1(n8864), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n5514) );
  NAND2_X1 U7026 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6580) );
  OAI211_X1 U7027 ( .C1(n4363), .C2(n5515), .A(n5514), .B(n6580), .ZN(n5521)
         );
  NAND2_X1 U7028 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n6565), .ZN(n5517) );
  OAI21_X1 U7029 ( .B1(n6565), .B2(P1_REG2_REG_10__SCAN_IN), .A(n5517), .ZN(
        n5518) );
  AOI211_X1 U7030 ( .C1(n5519), .C2(n5518), .A(n5848), .B(n8861), .ZN(n5520)
         );
  AOI211_X1 U7031 ( .C1(n5522), .C2(n9421), .A(n5521), .B(n5520), .ZN(n5523)
         );
  INV_X1 U7032 ( .A(n5523), .ZN(P1_U3251) );
  INV_X1 U7033 ( .A(n5567), .ZN(n5587) );
  XNOR2_X1 U7034 ( .A(n6589), .B(P2_B_REG_SCAN_IN), .ZN(n5524) );
  NAND2_X1 U7035 ( .A1(n5524), .A2(n6725), .ZN(n5526) );
  INV_X1 U7036 ( .A(n6839), .ZN(n5525) );
  INV_X1 U7037 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9634) );
  NAND2_X1 U7038 ( .A1(n9630), .A2(n9634), .ZN(n5528) );
  AND2_X1 U7039 ( .A1(n6589), .A2(n6839), .ZN(n9633) );
  INV_X1 U7040 ( .A(n9633), .ZN(n5527) );
  NAND2_X1 U7041 ( .A1(n5528), .A2(n5527), .ZN(n8352) );
  INV_X1 U7042 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9635) );
  AND2_X1 U7043 ( .A1(n6839), .A2(n6725), .ZN(n9636) );
  AOI21_X1 U7044 ( .B1(n9630), .B2(n9635), .A(n9636), .ZN(n8280) );
  NOR2_X1 U7045 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .ZN(
        n5532) );
  NOR4_X1 U7046 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5531) );
  NOR4_X1 U7047 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n5530) );
  NOR4_X1 U7048 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n5529) );
  NAND4_X1 U7049 ( .A1(n5532), .A2(n5531), .A3(n5530), .A4(n5529), .ZN(n5538)
         );
  NOR4_X1 U7050 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n5536) );
  NOR4_X1 U7051 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n5535) );
  NOR4_X1 U7052 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5534) );
  NOR4_X1 U7053 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n5533) );
  NAND4_X1 U7054 ( .A1(n5536), .A2(n5535), .A3(n5534), .A4(n5533), .ZN(n5537)
         );
  OAI21_X1 U7055 ( .B1(n5538), .B2(n5537), .A(n9630), .ZN(n8278) );
  AND2_X1 U7056 ( .A1(n8280), .A2(n8278), .ZN(n5733) );
  NAND2_X1 U7057 ( .A1(n8277), .A2(n5733), .ZN(n5959) );
  NAND2_X1 U7058 ( .A1(n5545), .A2(n5541), .ZN(n5542) );
  NAND2_X1 U7059 ( .A1(n5542), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5544) );
  XNOR2_X2 U7060 ( .A(n5544), .B(n5543), .ZN(n8286) );
  XNOR2_X2 U7061 ( .A(n5545), .B(P2_IR_REG_19__SCAN_IN), .ZN(n5547) );
  INV_X1 U7062 ( .A(n5547), .ZN(n8213) );
  AND2_X1 U7063 ( .A1(n8286), .A2(n8213), .ZN(n5572) );
  INV_X1 U7064 ( .A(n5572), .ZN(n7435) );
  INV_X1 U7065 ( .A(n5185), .ZN(n5574) );
  NAND2_X1 U7066 ( .A1(n9559), .A2(n9624), .ZN(n7973) );
  INV_X1 U7067 ( .A(n9639), .ZN(n7397) );
  NAND3_X1 U7068 ( .A1(n7397), .A2(n7427), .A3(n7253), .ZN(n5549) );
  NAND2_X1 U7069 ( .A1(n8286), .A2(n7429), .ZN(n5963) );
  INV_X1 U7071 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9794) );
  INV_X1 U7072 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n5554) );
  INV_X1 U7073 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n8264) );
  INV_X1 U7074 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5555) );
  INV_X1 U7075 ( .A(SI_0_), .ZN(n5564) );
  INV_X1 U7076 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5563) );
  OAI21_X1 U7077 ( .B1(n7244), .B2(n5564), .A(n5563), .ZN(n5565) );
  AND2_X1 U7078 ( .A1(n5566), .A2(n5565), .ZN(n8375) );
  MUX2_X1 U7079 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8375), .S(n5669), .Z(n9638) );
  INV_X1 U7080 ( .A(n9638), .ZN(n5750) );
  AOI22_X1 U7081 ( .A1(n8266), .A2(n4269), .B1(n7803), .B2(n5750), .ZN(n5568)
         );
  NAND2_X1 U7082 ( .A1(n5569), .A2(n5568), .ZN(n5666) );
  OAI21_X1 U7083 ( .B1(n5569), .B2(n5568), .A(n5666), .ZN(n5573) );
  NAND2_X1 U7084 ( .A1(n9719), .A2(n5575), .ZN(n5570) );
  NAND2_X1 U7085 ( .A1(n9606), .A2(n5547), .ZN(n8275) );
  NAND2_X1 U7086 ( .A1(n5571), .A2(n8238), .ZN(n5584) );
  OR2_X1 U7087 ( .A1(n5572), .A2(n5575), .ZN(n8276) );
  NAND2_X1 U7088 ( .A1(n5584), .A2(n8276), .ZN(n7030) );
  AOI22_X1 U7089 ( .A1(n5573), .A2(n9566), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n7030), .ZN(n5586) );
  OR2_X1 U7090 ( .A1(n5575), .A2(n5574), .ZN(n8251) );
  NAND2_X1 U7091 ( .A1(n9559), .A2(n9621), .ZN(n7970) );
  INV_X1 U7092 ( .A(n7970), .ZN(n7869) );
  INV_X1 U7093 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n9904) );
  OR2_X1 U7094 ( .A1(n5696), .A2(n9904), .ZN(n5583) );
  NAND2_X1 U7095 ( .A1(n5576), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5582) );
  OR2_X1 U7096 ( .A1(n5577), .A2(n6140), .ZN(n5581) );
  INV_X1 U7097 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5578) );
  OR2_X1 U7098 ( .A1(n5579), .A2(n5578), .ZN(n5580) );
  AOI22_X1 U7099 ( .A1(n7869), .A2(n5924), .B1(n9565), .B2(n9644), .ZN(n5585)
         );
  OAI211_X1 U7100 ( .C1(n5587), .C2(n7973), .A(n5586), .B(n5585), .ZN(P2_U3224) );
  INV_X1 U7101 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n5595) );
  INV_X1 U7102 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n5588) );
  MUX2_X1 U7103 ( .A(n5588), .B(P2_REG1_REG_10__SCAN_IN), .S(n6277), .Z(n5591)
         );
  AOI21_X1 U7104 ( .B1(n5908), .B2(P2_REG1_REG_9__SCAN_IN), .A(n5589), .ZN(
        n5590) );
  NOR2_X1 U7105 ( .A1(n5590), .A2(n5591), .ZN(n5637) );
  AOI21_X1 U7106 ( .B1(n5591), .B2(n5590), .A(n5637), .ZN(n5592) );
  NAND2_X1 U7107 ( .A1(n9573), .A2(n5592), .ZN(n5594) );
  NAND2_X1 U7108 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n5593) );
  OAI211_X1 U7109 ( .C1(n8072), .C2(n5595), .A(n5594), .B(n5593), .ZN(n5601)
         );
  NAND2_X1 U7110 ( .A1(n6277), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5597) );
  OAI21_X1 U7111 ( .B1(n6277), .B2(P2_REG2_REG_10__SCAN_IN), .A(n5597), .ZN(
        n5598) );
  NOR2_X1 U7112 ( .A1(n5599), .A2(n5598), .ZN(n5633) );
  AOI211_X1 U7113 ( .C1(n5599), .C2(n5598), .A(n5633), .B(n9576), .ZN(n5600)
         );
  AOI211_X1 U7114 ( .C1(n9295), .C2(n6277), .A(n5601), .B(n5600), .ZN(n5602)
         );
  INV_X1 U7115 ( .A(n5602), .ZN(P2_U3255) );
  INV_X1 U7116 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n6665) );
  MUX2_X1 U7117 ( .A(n5605), .B(n5604), .S(n5603), .Z(n5608) );
  OAI211_X1 U7118 ( .C1(n5608), .C2(n5607), .A(P1_U4006), .B(n5606), .ZN(n5631) );
  OAI21_X1 U7119 ( .B1(n5611), .B2(n5610), .A(n5609), .ZN(n5620) );
  NAND2_X1 U7120 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3084), .ZN(n7214) );
  INV_X1 U7121 ( .A(n7214), .ZN(n5617) );
  AOI21_X1 U7122 ( .B1(n5614), .B2(n5613), .A(n5612), .ZN(n5615) );
  NOR2_X1 U7123 ( .A1(n8855), .A2(n5615), .ZN(n5616) );
  AOI211_X1 U7124 ( .C1(n9413), .C2(n7202), .A(n5617), .B(n5616), .ZN(n5618)
         );
  INV_X1 U7125 ( .A(n5618), .ZN(n5619) );
  AOI21_X1 U7126 ( .B1(n9422), .B2(n5620), .A(n5619), .ZN(n5621) );
  OAI211_X1 U7127 ( .C1(n6665), .C2(n9426), .A(n5631), .B(n5621), .ZN(P1_U3245) );
  INV_X1 U7128 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6667) );
  INV_X1 U7129 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6089) );
  OAI211_X1 U7130 ( .C1(n5624), .C2(n5623), .A(n9421), .B(n5622), .ZN(n5625)
         );
  OAI21_X1 U7131 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6089), .A(n5625), .ZN(n5630) );
  AOI211_X1 U7132 ( .C1(n5628), .C2(n5627), .A(n5626), .B(n8861), .ZN(n5629)
         );
  AOI211_X1 U7133 ( .C1(n9413), .C2(n5648), .A(n5630), .B(n5629), .ZN(n5632)
         );
  OAI211_X1 U7134 ( .C1(n6667), .C2(n9426), .A(n5632), .B(n5631), .ZN(P1_U3243) );
  INV_X1 U7135 ( .A(n9295), .ZN(n9575) );
  INV_X1 U7136 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n9781) );
  AOI22_X1 U7137 ( .A1(n6452), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n9781), .B2(
        n5643), .ZN(n5635) );
  AOI21_X1 U7138 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n6277), .A(n5633), .ZN(
        n5634) );
  NAND2_X1 U7139 ( .A1(n5634), .A2(n5635), .ZN(n5861) );
  OAI21_X1 U7140 ( .B1(n5635), .B2(n5634), .A(n5861), .ZN(n5636) );
  NAND2_X1 U7141 ( .A1(n5636), .A2(n9572), .ZN(n5642) );
  AND2_X1 U7142 ( .A1(P2_U3152), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6652) );
  AOI21_X1 U7143 ( .B1(n6277), .B2(P2_REG1_REG_10__SCAN_IN), .A(n5637), .ZN(
        n5639) );
  INV_X1 U7144 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6285) );
  MUX2_X1 U7145 ( .A(n6285), .B(P2_REG1_REG_11__SCAN_IN), .S(n6452), .Z(n5638)
         );
  NOR2_X1 U7146 ( .A1(n5639), .A2(n5638), .ZN(n5856) );
  INV_X1 U7147 ( .A(n9573), .ZN(n8030) );
  AOI211_X1 U7148 ( .C1(n5639), .C2(n5638), .A(n5856), .B(n8030), .ZN(n5640)
         );
  AOI211_X1 U7149 ( .C1(P2_ADDR_REG_11__SCAN_IN), .C2(n9578), .A(n6652), .B(
        n5640), .ZN(n5641) );
  OAI211_X1 U7150 ( .C1(n9575), .C2(n5643), .A(n5642), .B(n5641), .ZN(P2_U3256) );
  NAND2_X1 U7151 ( .A1(n5645), .A2(n5644), .ZN(n5647) );
  NAND2_X1 U7152 ( .A1(n7524), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5650) );
  NAND2_X1 U7153 ( .A1(n7566), .A2(n5648), .ZN(n5649) );
  NAND2_X1 U7154 ( .A1(n9480), .A2(n4263), .ZN(n5651) );
  AND2_X1 U7155 ( .A1(n9480), .A2(n7497), .ZN(n5652) );
  AOI21_X1 U7156 ( .B1(n8822), .B2(n6703), .A(n5652), .ZN(n5779) );
  XNOR2_X1 U7157 ( .A(n5778), .B(n5779), .ZN(n5776) );
  XNOR2_X1 U7158 ( .A(n5777), .B(n5776), .ZN(n5662) );
  INV_X1 U7159 ( .A(n5875), .ZN(n6081) );
  INV_X1 U7160 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5653) );
  NAND2_X1 U7161 ( .A1(n6341), .A2(n5653), .ZN(n5658) );
  NAND2_X1 U7162 ( .A1(n5785), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5656) );
  NAND2_X1 U7163 ( .A1(n5786), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5655) );
  OAI22_X1 U7164 ( .A1(n6081), .A2(n8500), .B1(n8487), .B2(n7215), .ZN(n5661)
         );
  INV_X1 U7165 ( .A(n8490), .ZN(n8512) );
  OAI22_X1 U7166 ( .A1(n8512), .A2(n6090), .B1(n5659), .B2(n6089), .ZN(n5660)
         );
  AOI211_X1 U7167 ( .C1(n5662), .C2(n8496), .A(n5661), .B(n5660), .ZN(n5663)
         );
  INV_X1 U7168 ( .A(n5663), .ZN(P1_U3235) );
  INV_X1 U7169 ( .A(n5664), .ZN(n5665) );
  NAND2_X1 U7170 ( .A1(n5666), .A2(n5665), .ZN(n7027) );
  NOR2_X1 U7171 ( .A1(n5925), .A2(n9606), .ZN(n5675) );
  OR2_X1 U7172 ( .A1(n5678), .A2(n5667), .ZN(n5670) );
  AND2_X1 U7173 ( .A1(n5670), .A2(n4821), .ZN(n5672) );
  OR2_X1 U7174 ( .A1(n7248), .A2(n9890), .ZN(n5671) );
  XNOR2_X1 U7175 ( .A(n5673), .B(n9649), .ZN(n5674) );
  NOR2_X1 U7176 ( .A1(n5675), .A2(n5674), .ZN(n5676) );
  AOI21_X1 U7177 ( .B1(n5675), .B2(n5674), .A(n5676), .ZN(n7028) );
  NAND2_X1 U7178 ( .A1(n7027), .A2(n7028), .ZN(n7026) );
  INV_X1 U7179 ( .A(n5676), .ZN(n5677) );
  NAND2_X1 U7180 ( .A1(n7026), .A2(n5677), .ZN(n5745) );
  OR2_X1 U7181 ( .A1(n5678), .A2(n5771), .ZN(n5681) );
  OR2_X1 U7182 ( .A1(n7248), .A2(n5679), .ZN(n5680) );
  XNOR2_X1 U7183 ( .A(n6309), .B(n5673), .ZN(n5689) );
  NAND2_X1 U7184 ( .A1(n5576), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5688) );
  INV_X1 U7185 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5683) );
  INV_X1 U7186 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5684) );
  OR2_X1 U7187 ( .A1(n5579), .A2(n5684), .ZN(n5686) );
  OR2_X1 U7188 ( .A1(n5696), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U7189 ( .A1(n7994), .A2(n5718), .ZN(n5690) );
  XOR2_X1 U7190 ( .A(n5689), .B(n5690), .Z(n5744) );
  INV_X1 U7191 ( .A(n5689), .ZN(n5691) );
  OR2_X1 U7192 ( .A1(n5678), .A2(n7204), .ZN(n5694) );
  OR2_X1 U7193 ( .A1(n7248), .A2(n5692), .ZN(n5693) );
  OAI211_X1 U7194 ( .C1(n6976), .C2(n5695), .A(n5694), .B(n5693), .ZN(n9552)
         );
  XOR2_X1 U7195 ( .A(n7847), .B(n9552), .Z(n5709) );
  NAND2_X1 U7196 ( .A1(n5576), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5707) );
  INV_X1 U7197 ( .A(n5713), .ZN(n5700) );
  INV_X1 U7198 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5698) );
  INV_X1 U7199 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5697) );
  NAND2_X1 U7200 ( .A1(n5698), .A2(n5697), .ZN(n5699) );
  NAND2_X1 U7201 ( .A1(n5700), .A2(n5699), .ZN(n9556) );
  INV_X1 U7202 ( .A(n9556), .ZN(n5701) );
  OR2_X1 U7203 ( .A1(n5577), .A2(n5702), .ZN(n5705) );
  INV_X1 U7204 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5703) );
  OR2_X1 U7205 ( .A1(n5579), .A2(n5703), .ZN(n5704) );
  NAND2_X1 U7206 ( .A1(n9623), .A2(n5718), .ZN(n5708) );
  NAND2_X1 U7207 ( .A1(n5709), .A2(n5708), .ZN(n9548) );
  NOR2_X1 U7208 ( .A1(n5709), .A2(n5708), .ZN(n9547) );
  NAND2_X1 U7209 ( .A1(n7222), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5717) );
  INV_X1 U7210 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5710) );
  OR2_X1 U7211 ( .A1(n7224), .A2(n5710), .ZN(n5716) );
  OR2_X1 U7212 ( .A1(n7228), .A2(n5711), .ZN(n5715) );
  OAI21_X1 U7213 ( .B1(n5713), .B2(P2_REG3_REG_5__SCAN_IN), .A(n5807), .ZN(
        n5732) );
  OR2_X1 U7214 ( .A1(n7168), .A2(n5732), .ZN(n5714) );
  AND2_X1 U7215 ( .A1(n7993), .A2(n5718), .ZN(n5724) );
  OR2_X1 U7216 ( .A1(n5996), .A2(n5678), .ZN(n5721) );
  OR2_X1 U7217 ( .A1(n7248), .A2(n5719), .ZN(n5720) );
  OAI211_X1 U7218 ( .C1(n6976), .C2(n5722), .A(n5721), .B(n5720), .ZN(n9610)
         );
  INV_X2 U7219 ( .A(n7803), .ZN(n7847) );
  XNOR2_X1 U7220 ( .A(n9610), .B(n7847), .ZN(n5723) );
  NOR2_X1 U7221 ( .A1(n5724), .A2(n5723), .ZN(n5800) );
  INV_X1 U7222 ( .A(n5800), .ZN(n5725) );
  NAND2_X1 U7223 ( .A1(n5724), .A2(n5723), .ZN(n5799) );
  NAND2_X1 U7224 ( .A1(n5725), .A2(n5799), .ZN(n5726) );
  XNOR2_X1 U7225 ( .A(n5801), .B(n5726), .ZN(n5743) );
  INV_X1 U7226 ( .A(n7973), .ZN(n7792) );
  NAND2_X1 U7227 ( .A1(n7222), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5731) );
  OR2_X1 U7228 ( .A1(n7224), .A2(n9735), .ZN(n5730) );
  OR2_X1 U7229 ( .A1(n7228), .A2(n5222), .ZN(n5729) );
  INV_X1 U7230 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5727) );
  XNOR2_X1 U7231 ( .A(n5807), .B(n5727), .ZN(n6125) );
  OR2_X1 U7232 ( .A1(n7168), .A2(n6125), .ZN(n5728) );
  NAND4_X1 U7233 ( .A1(n5731), .A2(n5730), .A3(n5729), .A4(n5728), .ZN(n9622)
         );
  AOI22_X1 U7234 ( .A1(n7792), .A2(n9623), .B1(n7869), .B2(n9622), .ZN(n5742)
         );
  INV_X1 U7235 ( .A(n5732), .ZN(n9612) );
  INV_X1 U7236 ( .A(n5733), .ZN(n5734) );
  OAI21_X1 U7237 ( .B1(n8352), .B2(n5734), .A(n8275), .ZN(n5737) );
  NAND4_X1 U7238 ( .A1(n5737), .A2(n5736), .A3(n5735), .A4(n8276), .ZN(n5738)
         );
  NAND2_X1 U7239 ( .A1(n5738), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9571) );
  INV_X1 U7240 ( .A(n9571), .ZN(n7947) );
  INV_X1 U7241 ( .A(n9565), .ZN(n7950) );
  OAI21_X1 U7242 ( .B1(n7950), .B2(n9669), .A(n5739), .ZN(n5740) );
  AOI21_X1 U7243 ( .B1(n9612), .B2(n7947), .A(n5740), .ZN(n5741) );
  OAI211_X1 U7244 ( .C1(n5743), .C2(n7978), .A(n5742), .B(n5741), .ZN(P2_U3229) );
  XNOR2_X1 U7245 ( .A(n5745), .B(n5744), .ZN(n5749) );
  AOI22_X1 U7246 ( .A1(n7792), .A2(n5924), .B1(n7869), .B2(n9623), .ZN(n5748)
         );
  INV_X1 U7247 ( .A(n6309), .ZN(n9657) );
  OAI22_X1 U7248 ( .A1(n7950), .A2(n9657), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5698), .ZN(n5746) );
  AOI21_X1 U7249 ( .B1(n7947), .B2(n5698), .A(n5746), .ZN(n5747) );
  OAI211_X1 U7250 ( .C1(n5749), .C2(n7978), .A(n5748), .B(n5747), .ZN(P2_U3220) );
  INV_X1 U7251 ( .A(n7030), .ZN(n5755) );
  INV_X1 U7252 ( .A(n8257), .ZN(n7995) );
  AOI22_X1 U7253 ( .A1(n7869), .A2(n7995), .B1(n9565), .B2(n9638), .ZN(n5754)
         );
  OR2_X1 U7254 ( .A1(n5567), .A2(n5750), .ZN(n6174) );
  INV_X1 U7255 ( .A(n6174), .ZN(n8258) );
  NAND2_X1 U7256 ( .A1(n5567), .A2(n5750), .ZN(n7277) );
  INV_X1 U7257 ( .A(n7277), .ZN(n5751) );
  MUX2_X1 U7258 ( .A(n9638), .B(n5751), .S(n5718), .Z(n5752) );
  OAI21_X1 U7259 ( .B1(n8258), .B2(n5752), .A(n9566), .ZN(n5753) );
  OAI211_X1 U7260 ( .C1(n5755), .C2(n6175), .A(n5754), .B(n5753), .ZN(P2_U3234) );
  INV_X1 U7261 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5764) );
  INV_X1 U7262 ( .A(n5756), .ZN(n5760) );
  INV_X1 U7263 ( .A(n5757), .ZN(n5758) );
  NAND2_X1 U7264 ( .A1(n5758), .A2(SI_17_), .ZN(n5759) );
  MUX2_X1 U7265 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7244), .Z(n5822) );
  XNOR2_X1 U7266 ( .A(n5822), .B(SI_18_), .ZN(n5819) );
  XNOR2_X1 U7267 ( .A(n5821), .B(n5819), .ZN(n7546) );
  INV_X1 U7268 ( .A(n7546), .ZN(n5766) );
  NAND2_X1 U7269 ( .A1(n5762), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5763) );
  XNOR2_X1 U7270 ( .A(n5763), .B(P1_IR_REG_18__SCAN_IN), .ZN(n8874) );
  INV_X1 U7271 ( .A(n8874), .ZN(n8867) );
  OAI222_X1 U7272 ( .A1(n9275), .A2(n5764), .B1(n6728), .B2(n5766), .C1(
        P1_U3084), .C2(n8867), .ZN(P1_U3335) );
  INV_X1 U7273 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n5767) );
  NAND2_X1 U7274 ( .A1(n5490), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5765) );
  XNOR2_X1 U7275 ( .A(n5765), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8048) );
  NAND2_X1 U7276 ( .A1(n7566), .A2(n5768), .ZN(n5769) );
  NAND2_X1 U7277 ( .A1(n5773), .A2(n5772), .ZN(n5774) );
  AND2_X1 U7278 ( .A1(n5784), .A2(n7497), .ZN(n5775) );
  XNOR2_X1 U7279 ( .A(n6002), .B(n6003), .ZN(n6015) );
  NAND2_X1 U7280 ( .A1(n5777), .A2(n5776), .ZN(n6014) );
  INV_X1 U7281 ( .A(n5778), .ZN(n5780) );
  NAND2_X1 U7282 ( .A1(n6014), .A2(n6005), .ZN(n5781) );
  XOR2_X1 U7283 ( .A(n6015), .B(n5781), .Z(n5795) );
  INV_X1 U7284 ( .A(n8500), .ZN(n5793) );
  NAND2_X1 U7285 ( .A1(n5782), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8485) );
  OAI21_X1 U7286 ( .B1(n8485), .B2(P1_REG3_REG_3__SCAN_IN), .A(n5783), .ZN(
        n5792) );
  INV_X1 U7287 ( .A(n5784), .ZN(n6213) );
  OAI21_X1 U7288 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n5987), .ZN(n6204) );
  INV_X1 U7289 ( .A(n6204), .ZN(n7212) );
  NAND2_X1 U7290 ( .A1(n6341), .A2(n7212), .ZN(n5789) );
  NAND2_X1 U7291 ( .A1(n5785), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5788) );
  NAND2_X1 U7292 ( .A1(n5786), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5787) );
  NAND4_X1 U7293 ( .A1(n5790), .A2(n5789), .A3(n5788), .A4(n5787), .ZN(n8820)
         );
  INV_X1 U7294 ( .A(n8820), .ZN(n6071) );
  OAI22_X1 U7295 ( .A1(n8512), .A2(n6213), .B1(n6071), .B2(n8487), .ZN(n5791)
         );
  AOI211_X1 U7296 ( .C1(n5793), .C2(n8822), .A(n5792), .B(n5791), .ZN(n5794)
         );
  OAI21_X1 U7297 ( .B1(n5795), .B2(n8519), .A(n5794), .ZN(P1_U3216) );
  NAND2_X1 U7298 ( .A1(n9622), .A2(n5718), .ZN(n6043) );
  OR2_X1 U7299 ( .A1(n6148), .A2(n5678), .ZN(n5798) );
  AOI22_X1 U7300 ( .A1(n7080), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n7079), .B2(
        n5796), .ZN(n5797) );
  NAND2_X1 U7301 ( .A1(n5798), .A2(n5797), .ZN(n6127) );
  XNOR2_X1 U7302 ( .A(n6127), .B(n7847), .ZN(n6041) );
  XOR2_X1 U7303 ( .A(n6043), .B(n6041), .Z(n5803) );
  OAI21_X1 U7304 ( .B1(n5801), .B2(n5800), .A(n5799), .ZN(n5802) );
  AOI21_X1 U7305 ( .B1(n5803), .B2(n5802), .A(n6042), .ZN(n5818) );
  NAND2_X1 U7306 ( .A1(n7222), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5812) );
  OR2_X1 U7307 ( .A1(n7224), .A2(n5804), .ZN(n5811) );
  OR2_X1 U7308 ( .A1(n7228), .A2(n5223), .ZN(n5810) );
  INV_X1 U7309 ( .A(n5807), .ZN(n5805) );
  AOI21_X1 U7310 ( .B1(n5805), .B2(P2_REG3_REG_6__SCAN_IN), .A(
        P2_REG3_REG_7__SCAN_IN), .ZN(n5808) );
  NAND2_X1 U7311 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_REG3_REG_6__SCAN_IN), 
        .ZN(n5806) );
  OR2_X1 U7312 ( .A1(n5808), .A2(n5947), .ZN(n7793) );
  OR2_X1 U7313 ( .A1(n7168), .A2(n7793), .ZN(n5809) );
  NAND4_X1 U7314 ( .A1(n5812), .A2(n5811), .A3(n5810), .A4(n5809), .ZN(n7992)
         );
  AOI22_X1 U7315 ( .A1(n7792), .A2(n7993), .B1(n7869), .B2(n7992), .ZN(n5817)
         );
  INV_X1 U7316 ( .A(n6125), .ZN(n5815) );
  OAI21_X1 U7317 ( .B1(n7950), .B2(n9676), .A(n5813), .ZN(n5814) );
  AOI21_X1 U7318 ( .B1(n5815), .B2(n7947), .A(n5814), .ZN(n5816) );
  OAI211_X1 U7319 ( .C1(n5818), .C2(n7978), .A(n5817), .B(n5816), .ZN(P2_U3241) );
  INV_X1 U7320 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n5829) );
  INV_X1 U7321 ( .A(n5819), .ZN(n5820) );
  NAND2_X1 U7322 ( .A1(n5821), .A2(n5820), .ZN(n5824) );
  NAND2_X1 U7323 ( .A1(n5822), .A2(SI_18_), .ZN(n5823) );
  INV_X1 U7324 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n5831) );
  MUX2_X1 U7325 ( .A(n5829), .B(n5831), .S(n7244), .Z(n5826) );
  INV_X1 U7326 ( .A(SI_19_), .ZN(n5825) );
  NAND2_X1 U7327 ( .A1(n5826), .A2(n5825), .ZN(n5834) );
  INV_X1 U7328 ( .A(n5826), .ZN(n5827) );
  NAND2_X1 U7329 ( .A1(n5827), .A2(SI_19_), .ZN(n5828) );
  NAND2_X1 U7330 ( .A1(n5834), .A2(n5828), .ZN(n5833) );
  XNOR2_X1 U7331 ( .A(n5832), .B(n5833), .ZN(n7565) );
  INV_X1 U7332 ( .A(n7565), .ZN(n5830) );
  OAI222_X1 U7333 ( .A1(n9275), .A2(n5831), .B1(n9273), .B2(n5830), .C1(
        P1_U3084), .C2(n9026), .ZN(P1_U3334) );
  INV_X1 U7334 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7091) );
  INV_X1 U7335 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n5839) );
  MUX2_X1 U7336 ( .A(n7091), .B(n5839), .S(n7244), .Z(n5835) );
  INV_X1 U7337 ( .A(SI_20_), .ZN(n9834) );
  NAND2_X1 U7338 ( .A1(n5835), .A2(n9834), .ZN(n5871) );
  INV_X1 U7339 ( .A(n5835), .ZN(n5836) );
  NAND2_X1 U7340 ( .A1(n5836), .A2(SI_20_), .ZN(n5837) );
  XNOR2_X1 U7341 ( .A(n5870), .B(n5869), .ZN(n7586) );
  INV_X1 U7342 ( .A(n7586), .ZN(n5838) );
  OAI222_X1 U7343 ( .A1(n4268), .A2(n5838), .B1(n8286), .B2(P2_U3152), .C1(
        n7091), .C2(n8371), .ZN(P2_U3338) );
  OAI222_X1 U7344 ( .A1(n9275), .A2(n5839), .B1(n9273), .B2(n5838), .C1(n8772), 
        .C2(P1_U3084), .ZN(P1_U3333) );
  INV_X1 U7345 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9405) );
  AOI22_X1 U7346 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n6730), .B1(n5845), .B2(
        n9405), .ZN(n5843) );
  INV_X1 U7347 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n5840) );
  AOI22_X1 U7348 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n8828), .B1(n5847), .B2(
        n5840), .ZN(n8831) );
  OAI21_X1 U7349 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n6565), .A(n5841), .ZN(
        n8830) );
  NAND2_X1 U7350 ( .A1(n8831), .A2(n8830), .ZN(n8829) );
  OAI21_X1 U7351 ( .B1(n5843), .B2(n5842), .A(n6237), .ZN(n5854) );
  NAND2_X1 U7352 ( .A1(n8864), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n5844) );
  NAND2_X1 U7353 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6883) );
  OAI211_X1 U7354 ( .C1(n4363), .C2(n5845), .A(n5844), .B(n6883), .ZN(n5853)
         );
  INV_X1 U7355 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n5846) );
  AOI22_X1 U7356 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n8828), .B1(n5847), .B2(
        n5846), .ZN(n8826) );
  OAI21_X1 U7357 ( .B1(n8828), .B2(P1_REG2_REG_11__SCAN_IN), .A(n8824), .ZN(
        n5851) );
  NAND2_X1 U7358 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n6730), .ZN(n5849) );
  OAI21_X1 U7359 ( .B1(n6730), .B2(P1_REG2_REG_12__SCAN_IN), .A(n5849), .ZN(
        n5850) );
  NOR2_X1 U7360 ( .A1(n5851), .A2(n5850), .ZN(n6241) );
  AOI211_X1 U7361 ( .C1(n5851), .C2(n5850), .A(n6241), .B(n8861), .ZN(n5852)
         );
  AOI211_X1 U7362 ( .C1(n5854), .C2(n9421), .A(n5853), .B(n5852), .ZN(n5855)
         );
  INV_X1 U7363 ( .A(n5855), .ZN(P1_U3253) );
  AOI21_X1 U7364 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n6452), .A(n5856), .ZN(
        n5858) );
  INV_X1 U7365 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9743) );
  AOI22_X1 U7366 ( .A1(n6600), .A2(P2_REG1_REG_12__SCAN_IN), .B1(n9743), .B2(
        n5860), .ZN(n5857) );
  NAND2_X1 U7367 ( .A1(n5858), .A2(n5857), .ZN(n5894) );
  OAI21_X1 U7368 ( .B1(n5858), .B2(n5857), .A(n5894), .ZN(n5867) );
  NAND2_X1 U7369 ( .A1(P2_U3152), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6613) );
  NAND2_X1 U7370 ( .A1(n9578), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n5859) );
  OAI211_X1 U7371 ( .C1(n9575), .C2(n5860), .A(n6613), .B(n5859), .ZN(n5866)
         );
  OAI21_X1 U7372 ( .B1(n6452), .B2(P2_REG2_REG_11__SCAN_IN), .A(n5861), .ZN(
        n5864) );
  NAND2_X1 U7373 ( .A1(n6600), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5862) );
  OAI21_X1 U7374 ( .B1(n6600), .B2(P2_REG2_REG_12__SCAN_IN), .A(n5862), .ZN(
        n5863) );
  NOR2_X1 U7375 ( .A1(n5863), .A2(n5864), .ZN(n5901) );
  AOI211_X1 U7376 ( .C1(n5864), .C2(n5863), .A(n5901), .B(n9576), .ZN(n5865)
         );
  AOI211_X1 U7377 ( .C1(n5867), .C2(n9573), .A(n5866), .B(n5865), .ZN(n5868)
         );
  INV_X1 U7378 ( .A(n5868), .ZN(P2_U3257) );
  NAND2_X1 U7379 ( .A1(n5872), .A2(n5871), .ZN(n6254) );
  INV_X1 U7380 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7102) );
  INV_X1 U7381 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n5874) );
  MUX2_X1 U7382 ( .A(n7102), .B(n5874), .S(n7244), .Z(n6250) );
  XNOR2_X1 U7383 ( .A(n6250), .B(SI_21_), .ZN(n6249) );
  XNOR2_X1 U7384 ( .A(n6254), .B(n6249), .ZN(n7604) );
  INV_X1 U7385 ( .A(n7604), .ZN(n5873) );
  OAI222_X1 U7386 ( .A1(n4268), .A2(n5873), .B1(n7253), .B2(P2_U3152), .C1(
        n7102), .C2(n8371), .ZN(P2_U3337) );
  OAI222_X1 U7387 ( .A1(n9275), .A2(n5874), .B1(n6728), .B2(n5873), .C1(n8773), 
        .C2(P1_U3084), .ZN(P1_U3332) );
  INV_X1 U7388 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5890) );
  XNOR2_X2 U7389 ( .A(n5875), .B(n8650), .ZN(n6100) );
  NAND2_X1 U7390 ( .A1(n8823), .A2(n5887), .ZN(n6094) );
  NAND2_X1 U7391 ( .A1(n6081), .A2(n8650), .ZN(n5876) );
  NAND2_X1 U7392 ( .A1(n8654), .A2(n8655), .ZN(n5881) );
  NAND2_X1 U7393 ( .A1(n5882), .A2(n6090), .ZN(n5877) );
  NAND2_X1 U7394 ( .A1(n7215), .A2(n5784), .ZN(n8658) );
  NAND2_X1 U7395 ( .A1(n8821), .A2(n6213), .ZN(n6356) );
  NAND2_X1 U7396 ( .A1(n8658), .A2(n6356), .ZN(n6069) );
  INV_X1 U7397 ( .A(n6069), .ZN(n8735) );
  XNOR2_X1 U7398 ( .A(n6070), .B(n8735), .ZN(n6214) );
  NAND2_X1 U7399 ( .A1(n5449), .A2(n8917), .ZN(n5879) );
  NAND2_X1 U7400 ( .A1(n8794), .A2(n8727), .ZN(n5878) );
  INV_X1 U7401 ( .A(n6100), .ZN(n8741) );
  NAND2_X1 U7402 ( .A1(n8741), .A2(n6096), .ZN(n6097) );
  NAND2_X1 U7403 ( .A1(n6081), .A2(n9473), .ZN(n5880) );
  OAI21_X1 U7404 ( .B1(n8735), .B2(n6366), .A(n6195), .ZN(n5886) );
  OAI22_X1 U7405 ( .A1(n5882), .A2(n9060), .B1(n6071), .B2(n9062), .ZN(n5885)
         );
  NAND3_X1 U7406 ( .A1(n5883), .A2(n7675), .A3(n9026), .ZN(n6843) );
  NOR2_X1 U7407 ( .A1(n6214), .A2(n6843), .ZN(n5884) );
  AOI211_X1 U7408 ( .C1(n9117), .C2(n5886), .A(n5885), .B(n5884), .ZN(n6219)
         );
  AOI21_X1 U7409 ( .B1(n5784), .B2(n6086), .A(n4744), .ZN(n6217) );
  INV_X1 U7410 ( .A(n9519), .ZN(n9502) );
  AOI22_X1 U7411 ( .A1(n6217), .A2(n9502), .B1(n9216), .B2(n5784), .ZN(n5888)
         );
  OAI211_X1 U7412 ( .C1(n6214), .C2(n9505), .A(n6219), .B(n5888), .ZN(n5892)
         );
  NAND2_X1 U7413 ( .A1(n5892), .A2(n9528), .ZN(n5889) );
  OAI21_X1 U7414 ( .B1(n9528), .B2(n5890), .A(n5889), .ZN(P1_U3463) );
  AND2_X2 U7415 ( .A1(n5891), .A2(n6391), .ZN(n9544) );
  NAND2_X1 U7416 ( .A1(n5892), .A2(n9544), .ZN(n5893) );
  OAI21_X1 U7417 ( .B1(n9544), .B2(n5127), .A(n5893), .ZN(P1_U3526) );
  INV_X1 U7418 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9385) );
  AOI22_X1 U7419 ( .A1(n6762), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n9385), .B2(
        n5898), .ZN(n5896) );
  OAI21_X1 U7420 ( .B1(n6600), .B2(P2_REG1_REG_12__SCAN_IN), .A(n5894), .ZN(
        n5895) );
  NAND2_X1 U7421 ( .A1(n5896), .A2(n5895), .ZN(n6220) );
  OAI21_X1 U7422 ( .B1(n5896), .B2(n5895), .A(n6220), .ZN(n5900) );
  NAND2_X1 U7423 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6771) );
  NAND2_X1 U7424 ( .A1(n9578), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n5897) );
  OAI211_X1 U7425 ( .C1(n9575), .C2(n5898), .A(n6771), .B(n5897), .ZN(n5899)
         );
  AOI21_X1 U7426 ( .B1(n5900), .B2(n9573), .A(n5899), .ZN(n5907) );
  NOR2_X1 U7427 ( .A1(n6762), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5902) );
  AOI21_X1 U7428 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n6762), .A(n5902), .ZN(
        n5903) );
  OAI21_X1 U7429 ( .B1(n5904), .B2(n5903), .A(n6227), .ZN(n5905) );
  NAND2_X1 U7430 ( .A1(n5905), .A2(n9572), .ZN(n5906) );
  NAND2_X1 U7431 ( .A1(n5907), .A2(n5906), .ZN(P2_U3258) );
  NAND2_X1 U7432 ( .A1(n6346), .A2(n7235), .ZN(n5910) );
  AOI22_X1 U7433 ( .A1(n7080), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7079), .B2(
        n5908), .ZN(n5909) );
  NAND2_X1 U7434 ( .A1(n5576), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5917) );
  INV_X1 U7435 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5966) );
  OR2_X1 U7436 ( .A1(n7228), .A2(n5966), .ZN(n5916) );
  INV_X1 U7437 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5911) );
  OR2_X1 U7438 ( .A1(n5579), .A2(n5911), .ZN(n5915) );
  NAND2_X1 U7439 ( .A1(n5947), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5949) );
  INV_X1 U7440 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5912) );
  NAND2_X1 U7441 ( .A1(n5949), .A2(n5912), .ZN(n5913) );
  NAND2_X1 U7442 ( .A1(n5976), .A2(n5913), .ZN(n9570) );
  OR2_X1 U7443 ( .A1(n7168), .A2(n9570), .ZN(n5914) );
  NAND4_X1 U7444 ( .A1(n5917), .A2(n5916), .A3(n5915), .A4(n5914), .ZN(n7990)
         );
  NAND2_X1 U7445 ( .A1(n9693), .A2(n6519), .ZN(n7313) );
  NAND2_X1 U7446 ( .A1(n8266), .A2(n9644), .ZN(n5918) );
  NAND2_X1 U7447 ( .A1(n5918), .A2(n8257), .ZN(n5922) );
  INV_X1 U7448 ( .A(n8266), .ZN(n5920) );
  INV_X1 U7449 ( .A(n9644), .ZN(n5919) );
  NAND2_X1 U7450 ( .A1(n5920), .A2(n5919), .ZN(n5921) );
  NAND2_X1 U7451 ( .A1(n5922), .A2(n5921), .ZN(n6131) );
  INV_X1 U7452 ( .A(n5925), .ZN(n5924) );
  NAND2_X1 U7453 ( .A1(n5925), .A2(n9649), .ZN(n7279) );
  NAND2_X1 U7454 ( .A1(n6131), .A2(n7403), .ZN(n5927) );
  NAND2_X1 U7455 ( .A1(n5925), .A2(n5923), .ZN(n5926) );
  NAND2_X1 U7456 ( .A1(n5927), .A2(n5926), .ZN(n6300) );
  NAND2_X1 U7457 ( .A1(n7994), .A2(n9657), .ZN(n7284) );
  NAND2_X1 U7458 ( .A1(n6300), .A2(n7400), .ZN(n5929) );
  OR2_X1 U7459 ( .A1(n7994), .A2(n6309), .ZN(n5928) );
  NAND2_X1 U7460 ( .A1(n5929), .A2(n5928), .ZN(n6181) );
  INV_X1 U7461 ( .A(n9552), .ZN(n9663) );
  NAND2_X1 U7462 ( .A1(n9623), .A2(n9663), .ZN(n9615) );
  NAND2_X1 U7463 ( .A1(n6181), .A2(n7402), .ZN(n5931) );
  OR2_X1 U7464 ( .A1(n9623), .A2(n9552), .ZN(n5930) );
  NAND2_X1 U7465 ( .A1(n5931), .A2(n5930), .ZN(n9604) );
  NAND2_X1 U7466 ( .A1(n7993), .A2(n9669), .ZN(n7287) );
  NAND2_X1 U7467 ( .A1(n7272), .A2(n7287), .ZN(n9617) );
  NAND2_X1 U7468 ( .A1(n9604), .A2(n9617), .ZN(n5933) );
  OR2_X1 U7469 ( .A1(n7993), .A2(n9610), .ZN(n5932) );
  NAND2_X1 U7470 ( .A1(n5933), .A2(n5932), .ZN(n6118) );
  NAND2_X1 U7471 ( .A1(n9622), .A2(n9676), .ZN(n7288) );
  NAND2_X1 U7472 ( .A1(n7293), .A2(n7288), .ZN(n6119) );
  NAND2_X1 U7473 ( .A1(n6118), .A2(n6119), .ZN(n5935) );
  OR2_X1 U7474 ( .A1(n9622), .A2(n6127), .ZN(n5934) );
  NAND2_X1 U7475 ( .A1(n5935), .A2(n5934), .ZN(n6110) );
  INV_X1 U7476 ( .A(n7992), .ZN(n5939) );
  OR2_X1 U7477 ( .A1(n6321), .A2(n5678), .ZN(n5938) );
  AOI22_X1 U7478 ( .A1(n7080), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7079), .B2(
        n5936), .ZN(n5937) );
  NAND2_X1 U7479 ( .A1(n5938), .A2(n5937), .ZN(n6114) );
  OR2_X1 U7480 ( .A1(n5939), .A2(n6114), .ZN(n7305) );
  NAND2_X1 U7481 ( .A1(n5939), .A2(n6114), .ZN(n7298) );
  NAND2_X1 U7482 ( .A1(n7305), .A2(n7298), .ZN(n7295) );
  NAND2_X1 U7483 ( .A1(n6110), .A2(n7295), .ZN(n5941) );
  OR2_X1 U7484 ( .A1(n7992), .A2(n6114), .ZN(n5940) );
  NAND2_X1 U7485 ( .A1(n6330), .A2(n7235), .ZN(n5944) );
  AOI22_X1 U7486 ( .A1(n7080), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7079), .B2(
        n5942), .ZN(n5943) );
  NAND2_X1 U7487 ( .A1(n7222), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5953) );
  OR2_X1 U7488 ( .A1(n7224), .A2(n5945), .ZN(n5952) );
  OR2_X1 U7489 ( .A1(n7228), .A2(n5946), .ZN(n5951) );
  OR2_X1 U7490 ( .A1(n5947), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5948) );
  NAND2_X1 U7491 ( .A1(n5949), .A2(n5948), .ZN(n6268) );
  OR2_X1 U7492 ( .A1(n7168), .A2(n6268), .ZN(n5950) );
  NAND4_X1 U7493 ( .A1(n5953), .A2(n5952), .A3(n5951), .A4(n5950), .ZN(n7991)
         );
  INV_X1 U7494 ( .A(n7991), .ZN(n5954) );
  OR2_X1 U7495 ( .A1(n6270), .A2(n5954), .ZN(n7303) );
  NAND2_X1 U7496 ( .A1(n6270), .A2(n5954), .ZN(n7306) );
  NAND2_X1 U7497 ( .A1(n6270), .A2(n7991), .ZN(n5955) );
  INV_X1 U7498 ( .A(n6276), .ZN(n5956) );
  AOI21_X1 U7499 ( .B1(n5974), .B2(n5957), .A(n5956), .ZN(n9697) );
  INV_X1 U7500 ( .A(n8276), .ZN(n5958) );
  NOR2_X1 U7501 ( .A1(n5959), .A2(n5958), .ZN(n5960) );
  NAND2_X1 U7502 ( .A1(n8352), .A2(n5960), .ZN(n5965) );
  OR2_X1 U7503 ( .A1(n5962), .A2(n5547), .ZN(n9691) );
  OR2_X1 U7504 ( .A1(n5963), .A2(n8213), .ZN(n6281) );
  NAND2_X1 U7505 ( .A1(n9691), .A2(n6281), .ZN(n9628) );
  NOR2_X1 U7506 ( .A1(n9644), .A2(n9638), .ZN(n8255) );
  AND2_X1 U7507 ( .A1(n8255), .A2(n5923), .ZN(n6307) );
  NAND2_X1 U7508 ( .A1(n6307), .A2(n9657), .ZN(n6306) );
  INV_X1 U7509 ( .A(n6114), .ZN(n9682) );
  INV_X1 U7510 ( .A(n6294), .ZN(n5964) );
  AOI211_X1 U7511 ( .C1(n9693), .C2(n6266), .A(n4269), .B(n5964), .ZN(n9692)
         );
  OR2_X1 U7512 ( .A1(n5965), .A2(n5547), .ZN(n6478) );
  INV_X1 U7513 ( .A(n6478), .ZN(n9600) );
  INV_X1 U7514 ( .A(n8286), .ZN(n7428) );
  AND2_X1 U7515 ( .A1(n9639), .A2(n7428), .ZN(n9611) );
  NAND2_X1 U7516 ( .A1(n8265), .A2(n9611), .ZN(n8237) );
  NOR2_X1 U7517 ( .A1(n8237), .A2(n4448), .ZN(n5968) );
  OAI22_X1 U7518 ( .A1(n8265), .A2(n5966), .B1(n9570), .B2(n8238), .ZN(n5967)
         );
  AOI211_X1 U7519 ( .C1(n9692), .C2(n9600), .A(n5968), .B(n5967), .ZN(n5984)
         );
  NAND2_X1 U7520 ( .A1(n8257), .A2(n9644), .ZN(n7278) );
  NAND2_X1 U7521 ( .A1(n7278), .A2(n6174), .ZN(n8260) );
  NAND2_X1 U7522 ( .A1(n6134), .A2(n7279), .ZN(n5971) );
  INV_X1 U7523 ( .A(n7400), .ZN(n7281) );
  NAND2_X1 U7524 ( .A1(n5971), .A2(n7281), .ZN(n6182) );
  AND2_X1 U7525 ( .A1(n7269), .A2(n6183), .ZN(n7271) );
  NAND2_X1 U7526 ( .A1(n6182), .A2(n7271), .ZN(n9616) );
  AND2_X1 U7527 ( .A1(n9615), .A2(n7287), .ZN(n7268) );
  NAND2_X1 U7528 ( .A1(n9616), .A2(n7268), .ZN(n5972) );
  NAND2_X1 U7529 ( .A1(n5972), .A2(n7272), .ZN(n6121) );
  INV_X1 U7530 ( .A(n6119), .ZN(n7405) );
  INV_X1 U7531 ( .A(n7298), .ZN(n5973) );
  INV_X1 U7532 ( .A(n7407), .ZN(n6260) );
  INV_X1 U7533 ( .A(n5974), .ZN(n7409) );
  XNOR2_X1 U7534 ( .A(n6283), .B(n7409), .ZN(n5982) );
  OR2_X1 U7535 ( .A1(n8286), .A2(n7253), .ZN(n7256) );
  NAND2_X1 U7536 ( .A1(n7427), .A2(n7256), .ZN(n9619) );
  INV_X1 U7537 ( .A(n9619), .ZN(n9345) );
  NAND2_X1 U7538 ( .A1(n7222), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U7539 ( .A1(n5576), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5980) );
  INV_X1 U7540 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9791) );
  NAND2_X1 U7541 ( .A1(n5976), .A2(n9791), .ZN(n5977) );
  NAND2_X1 U7542 ( .A1(n6459), .A2(n5977), .ZN(n6518) );
  OR2_X1 U7543 ( .A1(n7168), .A2(n6518), .ZN(n5979) );
  INV_X1 U7544 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6293) );
  OR2_X1 U7545 ( .A1(n7228), .A2(n6293), .ZN(n5978) );
  NAND4_X1 U7546 ( .A1(n5981), .A2(n5980), .A3(n5979), .A4(n5978), .ZN(n7989)
         );
  AOI22_X1 U7547 ( .A1(n9621), .A2(n7989), .B1(n7991), .B2(n9624), .ZN(n9557)
         );
  OAI21_X1 U7548 ( .B1(n5982), .B2(n9345), .A(n9557), .ZN(n9699) );
  NAND2_X1 U7549 ( .A1(n9699), .A2(n8265), .ZN(n5983) );
  OAI211_X1 U7550 ( .C1(n9697), .C2(n8254), .A(n5984), .B(n5983), .ZN(P2_U3287) );
  NAND2_X1 U7551 ( .A1(n8615), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5993) );
  INV_X2 U7552 ( .A(n6026), .ZN(n7571) );
  INV_X1 U7553 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U7554 ( .A1(n5987), .A2(n5986), .ZN(n5988) );
  AND2_X1 U7555 ( .A1(n6029), .A2(n5988), .ZN(n6065) );
  NAND2_X1 U7556 ( .A1(n7571), .A2(n6065), .ZN(n5992) );
  NAND2_X1 U7557 ( .A1(n5786), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5991) );
  NAND2_X1 U7558 ( .A1(n5785), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U7559 ( .A1(n8819), .A2(n6703), .ZN(n5998) );
  INV_X2 U7560 ( .A(n6347), .ZN(n8612) );
  NAND2_X1 U7561 ( .A1(n7566), .A2(n5994), .ZN(n5995) );
  NAND2_X1 U7562 ( .A1(n9495), .A2(n7538), .ZN(n5997) );
  NAND2_X1 U7563 ( .A1(n5998), .A2(n5997), .ZN(n6416) );
  NAND2_X1 U7564 ( .A1(n8819), .A2(n4265), .ZN(n6000) );
  NAND2_X1 U7565 ( .A1(n9495), .A2(n4263), .ZN(n5999) );
  NAND2_X1 U7566 ( .A1(n6000), .A2(n5999), .ZN(n6001) );
  XNOR2_X1 U7567 ( .A(n6001), .B(n7675), .ZN(n6543) );
  INV_X1 U7568 ( .A(n6002), .ZN(n6004) );
  NAND2_X1 U7569 ( .A1(n6005), .A2(n6016), .ZN(n7206) );
  NAND2_X1 U7570 ( .A1(n8820), .A2(n7497), .ZN(n6009) );
  NAND2_X1 U7571 ( .A1(n7524), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U7572 ( .A1(n7566), .A2(n7202), .ZN(n6006) );
  NAND2_X1 U7573 ( .A1(n6209), .A2(n4263), .ZN(n6008) );
  NAND2_X1 U7574 ( .A1(n6009), .A2(n6008), .ZN(n6010) );
  XNOR2_X1 U7575 ( .A(n6010), .B(n7762), .ZN(n6020) );
  AND2_X1 U7576 ( .A1(n6209), .A2(n7497), .ZN(n6012) );
  AOI21_X1 U7577 ( .B1(n8820), .B2(n6703), .A(n6012), .ZN(n6021) );
  XNOR2_X1 U7578 ( .A(n6020), .B(n6021), .ZN(n7205) );
  NOR2_X1 U7579 ( .A1(n7206), .A2(n7205), .ZN(n6013) );
  NAND2_X1 U7580 ( .A1(n6014), .A2(n6013), .ZN(n6019) );
  INV_X1 U7581 ( .A(n6015), .ZN(n6017) );
  NAND2_X1 U7582 ( .A1(n6017), .A2(n6016), .ZN(n7208) );
  INV_X1 U7583 ( .A(n6020), .ZN(n6023) );
  INV_X1 U7584 ( .A(n6021), .ZN(n6022) );
  NAND2_X1 U7585 ( .A1(n6023), .A2(n6022), .ZN(n6024) );
  XNOR2_X1 U7586 ( .A(n6543), .B(n6414), .ZN(n6025) );
  NOR2_X1 U7587 ( .A1(n6025), .A2(n6416), .ZN(n6544) );
  AOI21_X1 U7588 ( .B1(n6416), .B2(n6025), .A(n6544), .ZN(n6040) );
  INV_X1 U7589 ( .A(n8511), .ZN(n8419) );
  NAND2_X1 U7590 ( .A1(n8615), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6034) );
  INV_X1 U7591 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6028) );
  NAND2_X1 U7592 ( .A1(n6029), .A2(n6028), .ZN(n6030) );
  AND2_X1 U7593 ( .A1(n6155), .A2(n6030), .ZN(n6555) );
  NAND2_X1 U7594 ( .A1(n7571), .A2(n6555), .ZN(n6033) );
  NAND2_X1 U7595 ( .A1(n5785), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6032) );
  NAND2_X1 U7596 ( .A1(n5786), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6031) );
  NAND4_X1 U7597 ( .A1(n6034), .A2(n6033), .A3(n6032), .A4(n6031), .ZN(n8818)
         );
  NAND2_X1 U7598 ( .A1(n8818), .A2(n9114), .ZN(n6036) );
  NAND2_X1 U7599 ( .A1(n8820), .A2(n9112), .ZN(n6035) );
  NAND2_X1 U7600 ( .A1(n6036), .A2(n6035), .ZN(n6057) );
  AOI21_X1 U7601 ( .B1(n8419), .B2(n6057), .A(n6037), .ZN(n6039) );
  AOI22_X1 U7602 ( .A1(n8490), .A2(n9495), .B1(n8517), .B2(n6065), .ZN(n6038)
         );
  OAI211_X1 U7603 ( .C1(n6040), .C2(n8519), .A(n6039), .B(n6038), .ZN(P1_U3225) );
  INV_X1 U7604 ( .A(n6041), .ZN(n6044) );
  XNOR2_X1 U7605 ( .A(n6114), .B(n7803), .ZN(n6046) );
  NAND2_X1 U7606 ( .A1(n7992), .A2(n5718), .ZN(n6045) );
  NOR2_X1 U7607 ( .A1(n6046), .A2(n6045), .ZN(n6047) );
  AOI21_X1 U7608 ( .B1(n6046), .B2(n6045), .A(n6047), .ZN(n7790) );
  XNOR2_X1 U7609 ( .A(n6270), .B(n7847), .ZN(n6511) );
  NAND2_X1 U7610 ( .A1(n7991), .A2(n5718), .ZN(n6512) );
  XNOR2_X1 U7611 ( .A(n6511), .B(n6512), .ZN(n6048) );
  OAI211_X1 U7612 ( .C1(n6049), .C2(n6048), .A(n6515), .B(n9566), .ZN(n6055)
         );
  INV_X1 U7613 ( .A(n9559), .ZN(n6052) );
  NAND2_X1 U7614 ( .A1(n7990), .A2(n9621), .ZN(n6051) );
  NAND2_X1 U7615 ( .A1(n7992), .A2(n9624), .ZN(n6050) );
  AND2_X1 U7616 ( .A1(n6051), .A2(n6050), .ZN(n6263) );
  INV_X1 U7617 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9780) );
  OAI22_X1 U7618 ( .A1(n6052), .A2(n6263), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9780), .ZN(n6053) );
  AOI21_X1 U7619 ( .B1(n9565), .B2(n6270), .A(n6053), .ZN(n6054) );
  OAI211_X1 U7620 ( .C1(n9571), .C2(n6268), .A(n6055), .B(n6054), .ZN(P2_U3223) );
  INV_X1 U7621 ( .A(n8819), .ZN(n7211) );
  NAND2_X1 U7622 ( .A1(n7211), .A2(n9495), .ZN(n6360) );
  NAND2_X1 U7623 ( .A1(n6071), .A2(n6209), .ZN(n8661) );
  AND2_X1 U7624 ( .A1(n8658), .A2(n8661), .ZN(n6363) );
  NAND2_X1 U7625 ( .A1(n6195), .A2(n6363), .ZN(n6200) );
  NAND2_X1 U7626 ( .A1(n6200), .A2(n6357), .ZN(n6056) );
  XOR2_X1 U7627 ( .A(n8736), .B(n6056), .Z(n6058) );
  AOI21_X1 U7628 ( .B1(n6058), .B2(n9117), .A(n6057), .ZN(n9499) );
  NAND3_X1 U7629 ( .A1(n6393), .A2(n6060), .A3(n6059), .ZN(n6061) );
  OAI21_X1 U7630 ( .B1(n6205), .B2(n6067), .A(n9502), .ZN(n6063) );
  NOR2_X1 U7631 ( .A1(n6063), .A2(n6168), .ZN(n9494) );
  INV_X1 U7632 ( .A(n9070), .ZN(n9321) );
  OR2_X1 U7633 ( .A1(n9321), .A2(n8917), .ZN(n6085) );
  INV_X1 U7634 ( .A(n6085), .ZN(n9064) );
  OR2_X2 U7635 ( .A1(n9433), .A2(n6064), .ZN(n9428) );
  INV_X1 U7636 ( .A(n9436), .ZN(n9309) );
  AOI22_X1 U7637 ( .A1(n9321), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n6065), .B2(
        n9309), .ZN(n6066) );
  OAI21_X1 U7638 ( .B1(n9428), .B2(n6067), .A(n6066), .ZN(n6068) );
  AOI21_X1 U7639 ( .B1(n9494), .B2(n9064), .A(n6068), .ZN(n6077) );
  NAND2_X1 U7640 ( .A1(n6070), .A2(n6069), .ZN(n6193) );
  NAND2_X1 U7641 ( .A1(n7215), .A2(n6213), .ZN(n6192) );
  NAND2_X1 U7642 ( .A1(n6071), .A2(n9488), .ZN(n6072) );
  AND2_X1 U7643 ( .A1(n6192), .A2(n6072), .ZN(n6074) );
  INV_X1 U7644 ( .A(n6072), .ZN(n6073) );
  NAND2_X1 U7645 ( .A1(n8661), .A2(n6357), .ZN(n6196) );
  AOI21_X1 U7646 ( .B1(n6193), .B2(n6074), .A(n4823), .ZN(n6075) );
  NAND2_X1 U7647 ( .A1(n6075), .A2(n8736), .ZN(n9496) );
  INV_X1 U7648 ( .A(n9121), .ZN(n9077) );
  NAND3_X1 U7649 ( .A1(n6144), .A2(n9496), .A3(n9077), .ZN(n6076) );
  OAI211_X1 U7650 ( .C1(n9499), .C2(n9433), .A(n6077), .B(n6076), .ZN(P1_U3286) );
  XNOR2_X1 U7651 ( .A(n6078), .B(n8733), .ZN(n9484) );
  OR3_X1 U7652 ( .A1(n9030), .A2(n6079), .A3(n9026), .ZN(n9313) );
  OAI21_X1 U7653 ( .B1(n8733), .B2(n8657), .A(n6080), .ZN(n6084) );
  OAI22_X1 U7654 ( .A1(n6081), .A2(n9060), .B1(n7215), .B2(n9062), .ZN(n6083)
         );
  NOR2_X1 U7655 ( .A1(n9484), .A2(n6843), .ZN(n6082) );
  AOI211_X1 U7656 ( .C1(n9117), .C2(n6084), .A(n6083), .B(n6082), .ZN(n9483)
         );
  MUX2_X1 U7657 ( .A(n5136), .B(n9483), .S(n9070), .Z(n6093) );
  OR2_X1 U7658 ( .A1(n6085), .A2(n9519), .ZN(n9429) );
  INV_X1 U7659 ( .A(n6103), .ZN(n6088) );
  INV_X1 U7660 ( .A(n6086), .ZN(n6087) );
  AOI21_X1 U7661 ( .B1(n9480), .B2(n6088), .A(n6087), .ZN(n9481) );
  OAI22_X1 U7662 ( .A1(n9428), .A2(n6090), .B1(n6089), .B2(n9436), .ZN(n6091)
         );
  AOI21_X1 U7663 ( .B1(n9100), .B2(n9481), .A(n6091), .ZN(n6092) );
  OAI211_X1 U7664 ( .C1(n9484), .C2(n9313), .A(n6093), .B(n6092), .ZN(P1_U3289) );
  INV_X1 U7665 ( .A(n6094), .ZN(n6095) );
  XNOR2_X1 U7666 ( .A(n6100), .B(n6095), .ZN(n9475) );
  INV_X1 U7667 ( .A(n6096), .ZN(n6099) );
  INV_X1 U7668 ( .A(n6097), .ZN(n6098) );
  AOI21_X1 U7669 ( .B1(n6100), .B2(n6099), .A(n6098), .ZN(n6102) );
  OAI21_X1 U7670 ( .B1(n6102), .B2(n9229), .A(n6101), .ZN(n9471) );
  OAI21_X1 U7671 ( .B1(n8650), .B2(n9427), .A(n9502), .ZN(n6104) );
  NOR2_X1 U7672 ( .A1(n6104), .A2(n6103), .ZN(n9472) );
  NAND2_X1 U7673 ( .A1(n9472), .A2(n9026), .ZN(n6105) );
  OAI21_X1 U7674 ( .B1(n9436), .B2(n6106), .A(n6105), .ZN(n6107) );
  OAI21_X1 U7675 ( .B1(n9471), .B2(n6107), .A(n9070), .ZN(n6109) );
  INV_X1 U7676 ( .A(n9070), .ZN(n9030) );
  AOI22_X1 U7677 ( .A1(n9031), .A2(n9473), .B1(P1_REG2_REG_1__SCAN_IN), .B2(
        n9030), .ZN(n6108) );
  OAI211_X1 U7678 ( .C1(n9121), .C2(n9475), .A(n6109), .B(n6108), .ZN(P1_U3290) );
  XNOR2_X1 U7679 ( .A(n6110), .B(n7295), .ZN(n9684) );
  INV_X1 U7680 ( .A(n9684), .ZN(n6117) );
  INV_X1 U7681 ( .A(n7295), .ZN(n7406) );
  XNOR2_X1 U7682 ( .A(n6111), .B(n7406), .ZN(n6112) );
  AOI222_X1 U7683 ( .A1(n9619), .A2(n6112), .B1(n9622), .B2(n9624), .C1(n7991), 
        .C2(n9621), .ZN(n9681) );
  MUX2_X1 U7684 ( .A(n5223), .B(n9681), .S(n8265), .Z(n6116) );
  OAI211_X1 U7685 ( .C1(n6123), .C2(n9682), .A(n9606), .B(n6265), .ZN(n9680)
         );
  OAI22_X1 U7686 ( .A1(n9680), .A2(n6478), .B1(n7793), .B2(n8238), .ZN(n6113)
         );
  AOI21_X1 U7687 ( .B1(n9591), .B2(n6114), .A(n6113), .ZN(n6115) );
  OAI211_X1 U7688 ( .C1(n6117), .C2(n8254), .A(n6116), .B(n6115), .ZN(P2_U3289) );
  XNOR2_X1 U7689 ( .A(n6118), .B(n6119), .ZN(n9678) );
  INV_X1 U7690 ( .A(n9678), .ZN(n6130) );
  OAI21_X1 U7691 ( .B1(n7405), .B2(n6121), .A(n6120), .ZN(n6122) );
  AOI222_X1 U7692 ( .A1(n9619), .A2(n6122), .B1(n7992), .B2(n9621), .C1(n7993), 
        .C2(n9624), .ZN(n9675) );
  MUX2_X1 U7693 ( .A(n5222), .B(n9675), .S(n8265), .Z(n6129) );
  OAI21_X1 U7694 ( .B1(n9609), .B2(n9676), .A(n9606), .ZN(n6124) );
  OR2_X1 U7695 ( .A1(n6124), .A2(n6123), .ZN(n9674) );
  OAI22_X1 U7696 ( .A1(n9674), .A2(n6478), .B1(n6125), .B2(n8238), .ZN(n6126)
         );
  AOI21_X1 U7697 ( .B1(n9591), .B2(n6127), .A(n6126), .ZN(n6128) );
  OAI211_X1 U7698 ( .C1(n6130), .C2(n8254), .A(n6129), .B(n6128), .ZN(P2_U3290) );
  XNOR2_X1 U7699 ( .A(n6131), .B(n5969), .ZN(n9653) );
  OAI21_X1 U7700 ( .B1(n8255), .B2(n5923), .A(n9606), .ZN(n6132) );
  OR2_X1 U7701 ( .A1(n6132), .A2(n6307), .ZN(n9651) );
  OAI22_X1 U7702 ( .A1(n6478), .A2(n9651), .B1(n9904), .B2(n8238), .ZN(n6133)
         );
  AOI21_X1 U7703 ( .B1(n9591), .B2(n9649), .A(n6133), .ZN(n6142) );
  NAND2_X1 U7704 ( .A1(n6135), .A2(n7403), .ZN(n6136) );
  NAND2_X1 U7705 ( .A1(n6301), .A2(n6136), .ZN(n6139) );
  INV_X1 U7706 ( .A(n9624), .ZN(n8249) );
  NAND2_X1 U7707 ( .A1(n7994), .A2(n9621), .ZN(n6137) );
  OAI21_X1 U7708 ( .B1(n8257), .B2(n8249), .A(n6137), .ZN(n6138) );
  AOI21_X1 U7709 ( .B1(n6139), .B2(n9619), .A(n6138), .ZN(n9656) );
  MUX2_X1 U7710 ( .A(n9656), .B(n6140), .S(n8217), .Z(n6141) );
  OAI211_X1 U7711 ( .C1(n9653), .C2(n8254), .A(n6142), .B(n6141), .ZN(P2_U3294) );
  NAND2_X1 U7712 ( .A1(n8819), .A2(n9495), .ZN(n6143) );
  INV_X1 U7713 ( .A(n8818), .ZN(n6315) );
  NAND2_X1 U7714 ( .A1(n8612), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U7715 ( .A1(n7566), .A2(n6145), .ZN(n6146) );
  NAND2_X1 U7716 ( .A1(n6315), .A2(n9501), .ZN(n6361) );
  NAND2_X1 U7717 ( .A1(n8818), .A2(n6314), .ZN(n6382) );
  NAND2_X1 U7718 ( .A1(n6150), .A2(n8737), .ZN(n6151) );
  NAND2_X1 U7719 ( .A1(n6317), .A2(n6151), .ZN(n6152) );
  INV_X1 U7720 ( .A(n6152), .ZN(n9506) );
  INV_X1 U7721 ( .A(n6843), .ZN(n9478) );
  NAND2_X1 U7722 ( .A1(n6152), .A2(n9478), .ZN(n6166) );
  AND2_X1 U7723 ( .A1(n6357), .A2(n6353), .ZN(n6359) );
  NAND2_X1 U7724 ( .A1(n6200), .A2(n6359), .ZN(n6381) );
  NAND2_X1 U7725 ( .A1(n6381), .A2(n6360), .ZN(n6153) );
  XNOR2_X1 U7726 ( .A(n6153), .B(n8737), .ZN(n6164) );
  NAND2_X1 U7727 ( .A1(n8615), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6160) );
  NAND2_X1 U7728 ( .A1(n6155), .A2(n6154), .ZN(n6156) );
  AND2_X1 U7729 ( .A1(n6339), .A2(n6156), .ZN(n8379) );
  NAND2_X1 U7730 ( .A1(n7571), .A2(n8379), .ZN(n6159) );
  NAND2_X1 U7731 ( .A1(n5785), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6158) );
  NAND2_X1 U7732 ( .A1(n5786), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6157) );
  NAND4_X1 U7733 ( .A1(n6160), .A2(n6159), .A3(n6158), .A4(n6157), .ZN(n8817)
         );
  NAND2_X1 U7734 ( .A1(n8817), .A2(n9114), .ZN(n6162) );
  NAND2_X1 U7735 ( .A1(n8819), .A2(n9112), .ZN(n6161) );
  NAND2_X1 U7736 ( .A1(n6162), .A2(n6161), .ZN(n6163) );
  AOI21_X1 U7737 ( .B1(n6164), .B2(n9117), .A(n6163), .ZN(n6165) );
  NAND2_X1 U7738 ( .A1(n6166), .A2(n6165), .ZN(n9507) );
  MUX2_X1 U7739 ( .A(n9507), .B(P1_REG2_REG_6__SCAN_IN), .S(n9433), .Z(n6167)
         );
  INV_X1 U7740 ( .A(n6167), .ZN(n6173) );
  OR2_X1 U7741 ( .A1(n6168), .A2(n6314), .ZN(n6169) );
  AND2_X1 U7742 ( .A1(n6389), .A2(n6169), .ZN(n9503) );
  INV_X1 U7743 ( .A(n6555), .ZN(n6170) );
  OAI22_X1 U7744 ( .A1(n9428), .A2(n6314), .B1(n9436), .B2(n6170), .ZN(n6171)
         );
  AOI21_X1 U7745 ( .B1(n9503), .B2(n9100), .A(n6171), .ZN(n6172) );
  OAI211_X1 U7746 ( .C1(n9506), .C2(n9313), .A(n6173), .B(n6172), .ZN(P1_U3285) );
  NAND2_X1 U7747 ( .A1(n6174), .A2(n7277), .ZN(n9640) );
  INV_X1 U7748 ( .A(n9640), .ZN(n6180) );
  OR2_X1 U7749 ( .A1(n6478), .A2(n5718), .ZN(n8078) );
  OAI21_X1 U7750 ( .B1(n9337), .B2(n9591), .A(n9638), .ZN(n6179) );
  AOI22_X1 U7751 ( .A1(n9640), .A2(n9619), .B1(n7995), .B2(n9621), .ZN(n9642)
         );
  OAI21_X1 U7752 ( .B1(n6175), .B2(n8238), .A(n9642), .ZN(n6177) );
  NOR2_X1 U7753 ( .A1(n8265), .A2(n5088), .ZN(n6176) );
  AOI21_X1 U7754 ( .B1(n8265), .B2(n6177), .A(n6176), .ZN(n6178) );
  OAI211_X1 U7755 ( .C1(n6180), .C2(n8254), .A(n6179), .B(n6178), .ZN(P2_U3296) );
  XNOR2_X1 U7756 ( .A(n6181), .B(n7402), .ZN(n9666) );
  INV_X1 U7757 ( .A(n9666), .ZN(n6191) );
  NAND2_X1 U7758 ( .A1(n6182), .A2(n6183), .ZN(n6184) );
  XNOR2_X1 U7759 ( .A(n7402), .B(n6184), .ZN(n6185) );
  AOI22_X1 U7760 ( .A1(n9621), .A2(n7993), .B1(n7994), .B2(n9624), .ZN(n9545)
         );
  OAI21_X1 U7761 ( .B1(n6185), .B2(n9345), .A(n9545), .ZN(n9664) );
  NAND2_X1 U7762 ( .A1(n9664), .A2(n8265), .ZN(n6190) );
  NOR2_X1 U7763 ( .A1(n8265), .A2(n5702), .ZN(n6188) );
  AOI21_X1 U7764 ( .B1(n6306), .B2(n9552), .A(n4269), .ZN(n6186) );
  NAND2_X1 U7765 ( .A1(n6186), .A2(n9605), .ZN(n9662) );
  OAI22_X1 U7766 ( .A1(n6478), .A2(n9662), .B1(n9556), .B2(n8238), .ZN(n6187)
         );
  AOI211_X1 U7767 ( .C1(n9591), .C2(n9552), .A(n6188), .B(n6187), .ZN(n6189)
         );
  OAI211_X1 U7768 ( .C1(n6191), .C2(n8254), .A(n6190), .B(n6189), .ZN(P2_U3292) );
  NAND2_X1 U7769 ( .A1(n6193), .A2(n6192), .ZN(n6194) );
  INV_X1 U7770 ( .A(n6196), .ZN(n8738) );
  XNOR2_X1 U7771 ( .A(n6194), .B(n8738), .ZN(n9487) );
  INV_X1 U7772 ( .A(n6357), .ZN(n6201) );
  INV_X1 U7773 ( .A(n6195), .ZN(n6198) );
  INV_X1 U7774 ( .A(n8658), .ZN(n6197) );
  OAI21_X1 U7775 ( .B1(n6198), .B2(n6197), .A(n6196), .ZN(n6199) );
  OAI211_X1 U7776 ( .C1(n6201), .C2(n6200), .A(n6199), .B(n9117), .ZN(n6203)
         );
  AOI22_X1 U7777 ( .A1(n9112), .A2(n8821), .B1(n8819), .B2(n9114), .ZN(n6202)
         );
  OAI211_X1 U7778 ( .C1(n9487), .C2(n6843), .A(n6203), .B(n6202), .ZN(n9490)
         );
  NAND2_X1 U7779 ( .A1(n9490), .A2(n9070), .ZN(n6211) );
  OAI22_X1 U7780 ( .A1(n9070), .A2(n4534), .B1(n6204), .B2(n9436), .ZN(n6208)
         );
  INV_X1 U7781 ( .A(n6205), .ZN(n6206) );
  OAI21_X1 U7782 ( .B1(n9488), .B2(n4744), .A(n6206), .ZN(n9489) );
  NOR2_X1 U7783 ( .A1(n9489), .A2(n9429), .ZN(n6207) );
  AOI211_X1 U7784 ( .C1(n9031), .C2(n6209), .A(n6208), .B(n6207), .ZN(n6210)
         );
  OAI211_X1 U7785 ( .C1(n9487), .C2(n9313), .A(n6211), .B(n6210), .ZN(P1_U3287) );
  AOI22_X1 U7786 ( .A1(n9030), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9309), .B2(
        n5653), .ZN(n6212) );
  OAI21_X1 U7787 ( .B1(n9428), .B2(n6213), .A(n6212), .ZN(n6216) );
  NOR2_X1 U7788 ( .A1(n6214), .A2(n9313), .ZN(n6215) );
  AOI211_X1 U7789 ( .C1(n6217), .C2(n9100), .A(n6216), .B(n6215), .ZN(n6218)
         );
  OAI21_X1 U7790 ( .B1(n6219), .B2(n9030), .A(n6218), .ZN(P1_U3288) );
  OAI21_X1 U7791 ( .B1(n6762), .B2(P2_REG1_REG_13__SCAN_IN), .A(n6220), .ZN(
        n6222) );
  INV_X1 U7792 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n6765) );
  MUX2_X1 U7793 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n6765), .S(n8000), .Z(n6221)
         );
  NAND2_X1 U7794 ( .A1(n6221), .A2(n6222), .ZN(n7999) );
  OAI21_X1 U7795 ( .B1(n6222), .B2(n6221), .A(n7999), .ZN(n6226) );
  INV_X1 U7796 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n6224) );
  NAND2_X1 U7797 ( .A1(n9295), .A2(n8000), .ZN(n6223) );
  NAND2_X1 U7798 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n6912) );
  OAI211_X1 U7799 ( .C1(n8072), .C2(n6224), .A(n6223), .B(n6912), .ZN(n6225)
         );
  AOI21_X1 U7800 ( .B1(n6226), .B2(n9573), .A(n6225), .ZN(n6234) );
  INV_X1 U7801 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6228) );
  MUX2_X1 U7802 ( .A(n6228), .B(P2_REG2_REG_14__SCAN_IN), .S(n8000), .Z(n6229)
         );
  INV_X1 U7803 ( .A(n6229), .ZN(n6230) );
  OAI21_X1 U7804 ( .B1(n6231), .B2(n6230), .A(n7996), .ZN(n6232) );
  NAND2_X1 U7805 ( .A1(n6232), .A2(n9572), .ZN(n6233) );
  NAND2_X1 U7806 ( .A1(n6234), .A2(n6233), .ZN(P2_U3259) );
  INV_X1 U7807 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n6248) );
  INV_X1 U7808 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6235) );
  AOI22_X1 U7809 ( .A1(P1_REG1_REG_13__SCAN_IN), .A2(n6861), .B1(n6236), .B2(
        n6235), .ZN(n6239) );
  OAI21_X1 U7810 ( .B1(n6239), .B2(n6238), .A(n6860), .ZN(n6240) );
  NAND2_X1 U7811 ( .A1(n6240), .A2(n9421), .ZN(n6247) );
  AND2_X1 U7812 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6967) );
  NAND2_X1 U7813 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n6861), .ZN(n6242) );
  OAI21_X1 U7814 ( .B1(n6861), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6242), .ZN(
        n6243) );
  AOI211_X1 U7815 ( .C1(n6244), .C2(n6243), .A(n6853), .B(n8861), .ZN(n6245)
         );
  AOI211_X1 U7816 ( .C1(n9413), .C2(n6861), .A(n6967), .B(n6245), .ZN(n6246)
         );
  OAI211_X1 U7817 ( .C1(n9426), .C2(n6248), .A(n6247), .B(n6246), .ZN(P1_U3254) );
  INV_X1 U7818 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n6259) );
  INV_X1 U7819 ( .A(n6249), .ZN(n6253) );
  INV_X1 U7820 ( .A(n6250), .ZN(n6251) );
  NAND2_X1 U7821 ( .A1(n6251), .A2(SI_21_), .ZN(n6252) );
  OAI21_X2 U7822 ( .B1(n6254), .B2(n6253), .A(n6252), .ZN(n6500) );
  INV_X1 U7823 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7113) );
  MUX2_X1 U7824 ( .A(n7113), .B(n6259), .S(n7244), .Z(n6256) );
  INV_X1 U7825 ( .A(SI_22_), .ZN(n6255) );
  NAND2_X1 U7826 ( .A1(n6256), .A2(n6255), .ZN(n6498) );
  INV_X1 U7827 ( .A(n6256), .ZN(n6257) );
  NAND2_X1 U7828 ( .A1(n6257), .A2(SI_22_), .ZN(n6258) );
  NAND2_X1 U7829 ( .A1(n6498), .A2(n6258), .ZN(n6499) );
  XNOR2_X1 U7830 ( .A(n6500), .B(n6499), .ZN(n7626) );
  INV_X1 U7831 ( .A(n7626), .ZN(n7033) );
  OAI222_X1 U7832 ( .A1(n9275), .A2(n6259), .B1(n6728), .B2(n7033), .C1(
        P1_U3084), .C2(n5414), .ZN(P1_U3331) );
  XNOR2_X1 U7833 ( .A(n6261), .B(n6260), .ZN(n9689) );
  INV_X1 U7834 ( .A(n9689), .ZN(n6274) );
  XNOR2_X1 U7835 ( .A(n6262), .B(n7407), .ZN(n6264) );
  OAI21_X1 U7836 ( .B1(n6264), .B2(n9345), .A(n6263), .ZN(n9687) );
  INV_X1 U7837 ( .A(n6265), .ZN(n6267) );
  OAI21_X1 U7838 ( .B1(n6267), .B2(n4449), .A(n6266), .ZN(n9686) );
  OAI22_X1 U7839 ( .A1(n8265), .A2(n5946), .B1(n6268), .B2(n8238), .ZN(n6269)
         );
  AOI21_X1 U7840 ( .B1(n9591), .B2(n6270), .A(n6269), .ZN(n6271) );
  OAI21_X1 U7841 ( .B1(n9686), .B2(n8078), .A(n6271), .ZN(n6272) );
  AOI21_X1 U7842 ( .B1(n9687), .B2(n8265), .A(n6272), .ZN(n6273) );
  OAI21_X1 U7843 ( .B1(n8254), .B2(n6274), .A(n6273), .ZN(P2_U3288) );
  OR2_X1 U7844 ( .A1(n9693), .A2(n7990), .ZN(n6275) );
  NAND2_X1 U7845 ( .A1(n6276), .A2(n6275), .ZN(n6471) );
  NAND2_X1 U7846 ( .A1(n6564), .A2(n7235), .ZN(n6279) );
  AOI22_X1 U7847 ( .A1(n7080), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7079), .B2(
        n6277), .ZN(n6278) );
  INV_X1 U7848 ( .A(n7989), .ZN(n6280) );
  OR2_X1 U7849 ( .A1(n9703), .A2(n6280), .ZN(n7299) );
  NAND2_X1 U7850 ( .A1(n9703), .A2(n6280), .ZN(n7265) );
  XNOR2_X1 U7851 ( .A(n6471), .B(n7399), .ZN(n9702) );
  INV_X1 U7852 ( .A(n6281), .ZN(n6282) );
  AND2_X1 U7853 ( .A1(n8265), .A2(n6282), .ZN(n9338) );
  INV_X1 U7854 ( .A(n9338), .ZN(n6798) );
  NAND2_X1 U7855 ( .A1(n6283), .A2(n7304), .ZN(n6284) );
  NAND2_X1 U7856 ( .A1(n6284), .A2(n7313), .ZN(n6450) );
  XNOR2_X1 U7857 ( .A(n6450), .B(n7399), .ZN(n6291) );
  NAND2_X1 U7858 ( .A1(n7222), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6289) );
  OR2_X1 U7859 ( .A1(n6455), .A2(n6285), .ZN(n6288) );
  OR2_X1 U7860 ( .A1(n7228), .A2(n9781), .ZN(n6287) );
  INV_X1 U7861 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n6457) );
  XNOR2_X1 U7862 ( .A(n6459), .B(n6457), .ZN(n6656) );
  OR2_X1 U7863 ( .A1(n7168), .A2(n6656), .ZN(n6286) );
  NAND4_X1 U7864 ( .A1(n6289), .A2(n6288), .A3(n6287), .A4(n6286), .ZN(n7988)
         );
  OAI22_X1 U7865 ( .A1(n6519), .A2(n8249), .B1(n6611), .B2(n8251), .ZN(n6290)
         );
  AOI21_X1 U7866 ( .B1(n6291), .B2(n9619), .A(n6290), .ZN(n6292) );
  OAI21_X1 U7867 ( .B1(n9702), .B2(n9691), .A(n6292), .ZN(n9706) );
  NAND2_X1 U7868 ( .A1(n9706), .A2(n8265), .ZN(n6299) );
  OAI22_X1 U7869 ( .A1(n8265), .A2(n6293), .B1(n6518), .B2(n8238), .ZN(n6297)
         );
  AND2_X1 U7870 ( .A1(n6294), .A2(n9703), .ZN(n6295) );
  OR2_X1 U7871 ( .A1(n6295), .A2(n6474), .ZN(n9705) );
  NOR2_X1 U7872 ( .A1(n9705), .A2(n8078), .ZN(n6296) );
  AOI211_X1 U7873 ( .C1(n9591), .C2(n9703), .A(n6297), .B(n6296), .ZN(n6298)
         );
  OAI211_X1 U7874 ( .C1(n9702), .C2(n6798), .A(n6299), .B(n6298), .ZN(P2_U3286) );
  XNOR2_X1 U7875 ( .A(n6300), .B(n7281), .ZN(n6308) );
  INV_X1 U7876 ( .A(n6182), .ZN(n6303) );
  AND3_X1 U7877 ( .A1(n6301), .A2(n7279), .A3(n7400), .ZN(n6302) );
  OAI21_X1 U7878 ( .B1(n6303), .B2(n6302), .A(n9619), .ZN(n6305) );
  AOI22_X1 U7879 ( .A1(n5924), .A2(n9624), .B1(n9621), .B2(n9623), .ZN(n6304)
         );
  OAI211_X1 U7880 ( .C1(n6308), .C2(n9691), .A(n6305), .B(n6304), .ZN(n9659)
         );
  OAI21_X1 U7881 ( .B1(n6307), .B2(n9657), .A(n6306), .ZN(n9658) );
  INV_X1 U7882 ( .A(n6308), .ZN(n9661) );
  AOI22_X1 U7883 ( .A1(n9661), .A2(n9338), .B1(n9591), .B2(n6309), .ZN(n6311)
         );
  INV_X1 U7884 ( .A(n8265), .ZN(n8217) );
  INV_X1 U7885 ( .A(n8238), .ZN(n9613) );
  AOI22_X1 U7886 ( .A1(n8217), .A2(P2_REG2_REG_3__SCAN_IN), .B1(n9613), .B2(
        n5698), .ZN(n6310) );
  OAI211_X1 U7887 ( .C1(n8078), .C2(n9658), .A(n6311), .B(n6310), .ZN(n6312)
         );
  AOI21_X1 U7888 ( .B1(n8265), .B2(n9659), .A(n6312), .ZN(n6313) );
  INV_X1 U7889 ( .A(n6313), .ZN(P2_U3293) );
  NAND2_X1 U7890 ( .A1(n6315), .A2(n6314), .ZN(n6316) );
  NAND2_X1 U7891 ( .A1(n6317), .A2(n6316), .ZN(n6380) );
  INV_X1 U7892 ( .A(n8817), .ZN(n6323) );
  NAND2_X1 U7893 ( .A1(n8612), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n6320) );
  NAND2_X1 U7894 ( .A1(n7566), .A2(n6318), .ZN(n6319) );
  NAND2_X1 U7895 ( .A1(n6323), .A2(n8380), .ZN(n6482) );
  INV_X1 U7896 ( .A(n8380), .ZN(n9511) );
  NAND2_X1 U7897 ( .A1(n6482), .A2(n8529), .ZN(n6385) );
  NOR2_X1 U7898 ( .A1(n8817), .A2(n8380), .ZN(n6324) );
  NAND2_X1 U7899 ( .A1(n8615), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6328) );
  XNOR2_X1 U7900 ( .A(n6339), .B(P1_REG3_REG_8__SCAN_IN), .ZN(n6490) );
  NAND2_X1 U7901 ( .A1(n7571), .A2(n6490), .ZN(n6327) );
  NAND2_X1 U7902 ( .A1(n5785), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6326) );
  NAND2_X1 U7903 ( .A1(n7591), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6325) );
  NAND4_X1 U7904 ( .A1(n6328), .A2(n6327), .A3(n6326), .A4(n6325), .ZN(n8816)
         );
  INV_X1 U7905 ( .A(n8816), .ZN(n6535) );
  NAND2_X1 U7906 ( .A1(n7642), .A2(n6330), .ZN(n6333) );
  NAND2_X1 U7907 ( .A1(n7566), .A2(n6331), .ZN(n6332) );
  NAND2_X1 U7908 ( .A1(n6535), .A2(n6493), .ZN(n8531) );
  INV_X1 U7909 ( .A(n6493), .ZN(n9518) );
  NAND2_X1 U7910 ( .A1(n8816), .A2(n9518), .ZN(n8666) );
  NAND2_X1 U7911 ( .A1(n8531), .A2(n8666), .ZN(n6631) );
  NAND2_X1 U7912 ( .A1(n6641), .A2(n6631), .ZN(n6335) );
  NAND2_X1 U7913 ( .A1(n8816), .A2(n6493), .ZN(n6634) );
  NAND2_X1 U7914 ( .A1(n6335), .A2(n6634), .ZN(n6351) );
  NAND2_X1 U7915 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .ZN(n6336) );
  INV_X1 U7916 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6338) );
  INV_X1 U7917 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6337) );
  OAI21_X1 U7918 ( .B1(n6339), .B2(n6338), .A(n6337), .ZN(n6340) );
  AND2_X1 U7919 ( .A1(n6370), .A2(n6340), .ZN(n6538) );
  NAND2_X1 U7920 ( .A1(n6341), .A2(n6538), .ZN(n6345) );
  NAND2_X1 U7921 ( .A1(n8615), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6344) );
  NAND2_X1 U7922 ( .A1(n7591), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6343) );
  NAND2_X1 U7923 ( .A1(n5785), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6342) );
  NAND4_X1 U7924 ( .A1(n6345), .A2(n6344), .A3(n6343), .A4(n6342), .ZN(n8815)
         );
  INV_X1 U7925 ( .A(n8815), .ZN(n6630) );
  NAND2_X1 U7926 ( .A1(n6346), .A2(n7642), .ZN(n6350) );
  AOI22_X1 U7927 ( .A1(n8612), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7566), .B2(
        n6348), .ZN(n6349) );
  NAND2_X1 U7928 ( .A1(n6630), .A2(n6636), .ZN(n8667) );
  NAND2_X1 U7929 ( .A1(n8815), .A2(n6629), .ZN(n8669) );
  NAND2_X1 U7930 ( .A1(n8667), .A2(n8669), .ZN(n8745) );
  XNOR2_X1 U7931 ( .A(n6351), .B(n8745), .ZN(n6404) );
  AOI21_X1 U7932 ( .B1(n6636), .B2(n6489), .A(n9235), .ZN(n6401) );
  AOI22_X1 U7933 ( .A1(n9030), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n6538), .B2(
        n9309), .ZN(n6352) );
  OAI21_X1 U7934 ( .B1(n9428), .B2(n6629), .A(n6352), .ZN(n6378) );
  INV_X1 U7935 ( .A(n6353), .ZN(n6354) );
  NAND2_X1 U7936 ( .A1(n6361), .A2(n6354), .ZN(n6355) );
  AND2_X1 U7937 ( .A1(n8529), .A2(n6382), .ZN(n6365) );
  NAND2_X1 U7938 ( .A1(n6355), .A2(n6365), .ZN(n8660) );
  NAND2_X1 U7939 ( .A1(n6357), .A2(n6356), .ZN(n6358) );
  NOR2_X1 U7940 ( .A1(n8660), .A2(n6358), .ZN(n8664) );
  INV_X1 U7941 ( .A(n6359), .ZN(n6362) );
  AND2_X1 U7942 ( .A1(n6361), .A2(n6360), .ZN(n8662) );
  OAI21_X1 U7943 ( .B1(n6363), .B2(n6362), .A(n8662), .ZN(n6364) );
  AND2_X1 U7944 ( .A1(n6482), .A2(n8531), .ZN(n8644) );
  NAND2_X1 U7945 ( .A1(n6621), .A2(n8666), .ZN(n6367) );
  XNOR2_X1 U7946 ( .A(n6367), .B(n8745), .ZN(n6376) );
  NAND2_X1 U7947 ( .A1(n8615), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6375) );
  INV_X1 U7948 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6369) );
  NAND2_X1 U7949 ( .A1(n6370), .A2(n6369), .ZN(n6371) );
  AND2_X1 U7950 ( .A1(n6574), .A2(n6371), .ZN(n9310) );
  NAND2_X1 U7951 ( .A1(n7571), .A2(n9310), .ZN(n6374) );
  NAND2_X1 U7952 ( .A1(n5785), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6373) );
  NAND2_X1 U7953 ( .A1(n7591), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6372) );
  NAND4_X1 U7954 ( .A1(n6375), .A2(n6374), .A3(n6373), .A4(n6372), .ZN(n8814)
         );
  AOI222_X1 U7955 ( .A1(n9117), .A2(n6376), .B1(n8814), .B2(n9114), .C1(n8816), 
        .C2(n9112), .ZN(n6403) );
  NOR2_X1 U7956 ( .A1(n6403), .A2(n9321), .ZN(n6377) );
  AOI211_X1 U7957 ( .C1(n6401), .C2(n9100), .A(n6378), .B(n6377), .ZN(n6379)
         );
  OAI21_X1 U7958 ( .B1(n9121), .B2(n6404), .A(n6379), .ZN(P1_U3282) );
  XNOR2_X1 U7959 ( .A(n6380), .B(n6385), .ZN(n9514) );
  INV_X1 U7960 ( .A(n9514), .ZN(n6400) );
  NAND2_X1 U7961 ( .A1(n6381), .A2(n8662), .ZN(n6383) );
  NAND2_X1 U7962 ( .A1(n6383), .A2(n6382), .ZN(n6386) );
  NAND2_X1 U7963 ( .A1(n6386), .A2(n6482), .ZN(n8530) );
  INV_X1 U7964 ( .A(n8529), .ZN(n6384) );
  NOR2_X1 U7965 ( .A1(n8530), .A2(n6384), .ZN(n6388) );
  INV_X1 U7966 ( .A(n6385), .ZN(n8743) );
  OAI21_X1 U7967 ( .B1(n6386), .B2(n8743), .A(n9117), .ZN(n6387) );
  AOI22_X1 U7968 ( .A1(n9112), .A2(n8818), .B1(n8816), .B2(n9114), .ZN(n8381)
         );
  OAI21_X1 U7969 ( .B1(n6388), .B2(n6387), .A(n8381), .ZN(n9512) );
  AOI21_X1 U7970 ( .B1(n6389), .B2(n8380), .A(n9519), .ZN(n6390) );
  NAND2_X1 U7971 ( .A1(n6390), .A2(n6487), .ZN(n9510) );
  NOR2_X1 U7972 ( .A1(n6391), .A2(n8917), .ZN(n6392) );
  AND2_X1 U7973 ( .A1(n6393), .A2(n6392), .ZN(n9317) );
  INV_X1 U7974 ( .A(n9317), .ZN(n6397) );
  INV_X1 U7975 ( .A(n8379), .ZN(n6394) );
  OAI22_X1 U7976 ( .A1(n9070), .A2(n5170), .B1(n6394), .B2(n9436), .ZN(n6395)
         );
  AOI21_X1 U7977 ( .B1(n9031), .B2(n8380), .A(n6395), .ZN(n6396) );
  OAI21_X1 U7978 ( .B1(n9510), .B2(n6397), .A(n6396), .ZN(n6398) );
  AOI21_X1 U7979 ( .B1(n9512), .B2(n9070), .A(n6398), .ZN(n6399) );
  OAI21_X1 U7980 ( .B1(n6400), .B2(n9121), .A(n6399), .ZN(P1_U3284) );
  AOI22_X1 U7981 ( .A1(n6401), .A2(n9502), .B1(n9216), .B2(n6636), .ZN(n6402)
         );
  OAI211_X1 U7982 ( .C1(n6404), .C2(n9208), .A(n6403), .B(n6402), .ZN(n6406)
         );
  NAND2_X1 U7983 ( .A1(n6406), .A2(n9544), .ZN(n6405) );
  OAI21_X1 U7984 ( .B1(n9544), .B2(n5344), .A(n6405), .ZN(P1_U3532) );
  INV_X1 U7985 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9803) );
  NAND2_X1 U7986 ( .A1(n6406), .A2(n9528), .ZN(n6407) );
  OAI21_X1 U7987 ( .B1(n9528), .B2(n9803), .A(n6407), .ZN(P1_U3481) );
  NAND2_X1 U7988 ( .A1(n8818), .A2(n7538), .ZN(n6409) );
  NAND2_X1 U7989 ( .A1(n9501), .A2(n4263), .ZN(n6408) );
  NAND2_X1 U7990 ( .A1(n6409), .A2(n6408), .ZN(n6410) );
  XNOR2_X1 U7991 ( .A(n6410), .B(n7762), .ZN(n6415) );
  NAND2_X1 U7992 ( .A1(n8818), .A2(n6703), .ZN(n6412) );
  NAND2_X1 U7993 ( .A1(n9501), .A2(n7538), .ZN(n6411) );
  AND2_X1 U7994 ( .A1(n6412), .A2(n6411), .ZN(n6418) );
  NAND2_X1 U7995 ( .A1(n6415), .A2(n6418), .ZN(n6549) );
  INV_X1 U7996 ( .A(n6415), .ZN(n6542) );
  NAND2_X1 U7997 ( .A1(n6543), .A2(n6416), .ZN(n6417) );
  NAND2_X1 U7998 ( .A1(n6417), .A2(n6418), .ZN(n6420) );
  INV_X1 U7999 ( .A(n6417), .ZN(n6419) );
  INV_X1 U8000 ( .A(n6418), .ZN(n6541) );
  AOI22_X1 U8001 ( .A1(n6542), .A2(n6420), .B1(n6419), .B2(n6541), .ZN(n6421)
         );
  NAND2_X1 U8002 ( .A1(n8817), .A2(n4265), .ZN(n6423) );
  NAND2_X1 U8003 ( .A1(n8380), .A2(n4263), .ZN(n6422) );
  NAND2_X1 U8004 ( .A1(n6423), .A2(n6422), .ZN(n6424) );
  XNOR2_X1 U8005 ( .A(n6424), .B(n7675), .ZN(n6428) );
  AND2_X1 U8006 ( .A1(n8380), .A2(n7538), .ZN(n6425) );
  AOI21_X1 U8007 ( .B1(n8817), .B2(n6703), .A(n6425), .ZN(n6426) );
  XNOR2_X1 U8008 ( .A(n6428), .B(n6426), .ZN(n8378) );
  INV_X1 U8009 ( .A(n6426), .ZN(n6427) );
  NAND2_X1 U8010 ( .A1(n6428), .A2(n6427), .ZN(n6429) );
  NAND2_X1 U8011 ( .A1(n8816), .A2(n6703), .ZN(n6431) );
  NAND2_X1 U8012 ( .A1(n6493), .A2(n7538), .ZN(n6430) );
  NAND2_X1 U8013 ( .A1(n6431), .A2(n6430), .ZN(n6434) );
  INV_X1 U8014 ( .A(n6434), .ZN(n6432) );
  INV_X1 U8015 ( .A(n6530), .ZN(n6439) );
  NAND2_X1 U8016 ( .A1(n6435), .A2(n6434), .ZN(n6441) );
  NAND2_X1 U8017 ( .A1(n8816), .A2(n4265), .ZN(n6437) );
  NAND2_X1 U8018 ( .A1(n6493), .A2(n4263), .ZN(n6436) );
  NAND2_X1 U8019 ( .A1(n6437), .A2(n6436), .ZN(n6438) );
  XNOR2_X1 U8020 ( .A(n6438), .B(n7762), .ZN(n6440) );
  NAND2_X1 U8021 ( .A1(n6441), .A2(n6440), .ZN(n6531) );
  NOR2_X1 U8022 ( .A1(n6439), .A2(n6531), .ZN(n6443) );
  AOI21_X1 U8023 ( .B1(n6530), .B2(n6441), .A(n6440), .ZN(n6442) );
  OAI21_X1 U8024 ( .B1(n6443), .B2(n6442), .A(n8496), .ZN(n6449) );
  NAND2_X1 U8025 ( .A1(n8815), .A2(n9114), .ZN(n6445) );
  NAND2_X1 U8026 ( .A1(n8817), .A2(n9112), .ZN(n6444) );
  AND2_X1 U8027 ( .A1(n6445), .A2(n6444), .ZN(n6484) );
  OAI21_X1 U8028 ( .B1(n8511), .B2(n6484), .A(n6446), .ZN(n6447) );
  AOI21_X1 U8029 ( .B1(n6490), .B2(n8517), .A(n6447), .ZN(n6448) );
  OAI211_X1 U8030 ( .C1(n9518), .C2(n8512), .A(n6449), .B(n6448), .ZN(P1_U3219) );
  NAND2_X1 U8031 ( .A1(n6450), .A2(n7299), .ZN(n6451) );
  NAND2_X1 U8032 ( .A1(n6617), .A2(n7235), .ZN(n6454) );
  AOI22_X1 U8033 ( .A1(n7080), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n7079), .B2(
        n6452), .ZN(n6453) );
  NAND2_X1 U8034 ( .A1(n6454), .A2(n6453), .ZN(n6776) );
  OR2_X1 U8035 ( .A1(n6776), .A2(n6611), .ZN(n9583) );
  NAND2_X1 U8036 ( .A1(n6776), .A2(n6611), .ZN(n7317) );
  NAND2_X1 U8037 ( .A1(n9583), .A2(n7317), .ZN(n7412) );
  XNOR2_X1 U8038 ( .A(n6784), .B(n7412), .ZN(n6469) );
  NAND2_X1 U8039 ( .A1(n7989), .A2(n9624), .ZN(n6467) );
  NAND2_X1 U8040 ( .A1(n7222), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6465) );
  OR2_X1 U8041 ( .A1(n6455), .A2(n9743), .ZN(n6464) );
  INV_X1 U8042 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6456) );
  OAI21_X1 U8043 ( .B1(n6459), .B2(n6457), .A(n6456), .ZN(n6460) );
  NAND2_X1 U8044 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_REG3_REG_11__SCAN_IN), 
        .ZN(n6458) );
  NAND2_X1 U8045 ( .A1(n6460), .A2(n6605), .ZN(n9588) );
  OR2_X1 U8046 ( .A1(n7168), .A2(n9588), .ZN(n6463) );
  INV_X1 U8047 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6461) );
  OR2_X1 U8048 ( .A1(n7228), .A2(n6461), .ZN(n6462) );
  NAND4_X1 U8049 ( .A1(n6465), .A2(n6464), .A3(n6463), .A4(n6462), .ZN(n7987)
         );
  NAND2_X1 U8050 ( .A1(n7987), .A2(n9621), .ZN(n6466) );
  NAND2_X1 U8051 ( .A1(n6467), .A2(n6466), .ZN(n6653) );
  INV_X1 U8052 ( .A(n6653), .ZN(n6468) );
  OAI21_X1 U8053 ( .B1(n6469), .B2(n9345), .A(n6468), .ZN(n9713) );
  INV_X1 U8054 ( .A(n9713), .ZN(n6481) );
  NAND2_X1 U8055 ( .A1(n9703), .A2(n7989), .ZN(n6470) );
  NAND2_X1 U8056 ( .A1(n6472), .A2(n7412), .ZN(n6778) );
  OAI21_X1 U8057 ( .B1(n6472), .B2(n7412), .A(n6778), .ZN(n6473) );
  INV_X1 U8058 ( .A(n6473), .ZN(n9715) );
  INV_X1 U8059 ( .A(n8254), .ZN(n9601) );
  INV_X1 U8060 ( .A(n6776), .ZN(n9712) );
  OAI21_X1 U8061 ( .B1(n6474), .B2(n9712), .A(n9606), .ZN(n6475) );
  OR2_X1 U8062 ( .A1(n9598), .A2(n6475), .ZN(n9711) );
  OAI22_X1 U8063 ( .A1(n8265), .A2(n9781), .B1(n6656), .B2(n8238), .ZN(n6476)
         );
  AOI21_X1 U8064 ( .B1(n9591), .B2(n6776), .A(n6476), .ZN(n6477) );
  OAI21_X1 U8065 ( .B1(n9711), .B2(n6478), .A(n6477), .ZN(n6479) );
  AOI21_X1 U8066 ( .B1(n9715), .B2(n9601), .A(n6479), .ZN(n6480) );
  OAI21_X1 U8067 ( .B1(n6481), .B2(n8217), .A(n6480), .ZN(P2_U3285) );
  INV_X1 U8068 ( .A(n6631), .ZN(n8742) );
  XNOR2_X1 U8069 ( .A(n6641), .B(n8742), .ZN(n9523) );
  NAND2_X1 U8070 ( .A1(n8779), .A2(n6482), .ZN(n6483) );
  XNOR2_X1 U8071 ( .A(n6483), .B(n6631), .ZN(n6485) );
  OAI21_X1 U8072 ( .B1(n6485), .B2(n9229), .A(n6484), .ZN(n6486) );
  AOI21_X1 U8073 ( .B1(n9523), .B2(n9478), .A(n6486), .ZN(n9525) );
  INV_X1 U8074 ( .A(n9313), .ZN(n6496) );
  NAND2_X1 U8075 ( .A1(n6487), .A2(n6493), .ZN(n6488) );
  NAND2_X1 U8076 ( .A1(n6489), .A2(n6488), .ZN(n9520) );
  INV_X1 U8077 ( .A(n6490), .ZN(n6491) );
  OAI22_X1 U8078 ( .A1(n9070), .A2(n5286), .B1(n6491), .B2(n9436), .ZN(n6492)
         );
  AOI21_X1 U8079 ( .B1(n9031), .B2(n6493), .A(n6492), .ZN(n6494) );
  OAI21_X1 U8080 ( .B1(n9520), .B2(n9429), .A(n6494), .ZN(n6495) );
  AOI21_X1 U8081 ( .B1(n9523), .B2(n6496), .A(n6495), .ZN(n6497) );
  OAI21_X1 U8082 ( .B1(n9525), .B2(n9030), .A(n6497), .ZN(P1_U3283) );
  INV_X1 U8083 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7121) );
  INV_X1 U8084 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n6501) );
  MUX2_X1 U8085 ( .A(n7121), .B(n6501), .S(n7244), .Z(n6503) );
  INV_X1 U8086 ( .A(SI_23_), .ZN(n6502) );
  NAND2_X1 U8087 ( .A1(n6503), .A2(n6502), .ZN(n6588) );
  INV_X1 U8088 ( .A(n6503), .ZN(n6504) );
  NAND2_X1 U8089 ( .A1(n6504), .A2(SI_23_), .ZN(n6505) );
  INV_X1 U8090 ( .A(n7476), .ZN(n6508) );
  OR2_X1 U8091 ( .A1(n6506), .A2(P1_U3084), .ZN(n8770) );
  NAND2_X1 U8092 ( .A1(n9265), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6507) );
  OAI211_X1 U8093 ( .C1(n6508), .C2(n9273), .A(n8770), .B(n6507), .ZN(P1_U3330) );
  NAND2_X1 U8094 ( .A1(n7476), .A2(n6509), .ZN(n6510) );
  OAI211_X1 U8095 ( .C1(n7121), .C2(n8371), .A(n6510), .B(n7438), .ZN(P2_U3335) );
  NAND2_X1 U8096 ( .A1(n6511), .A2(n6513), .ZN(n6514) );
  XNOR2_X1 U8097 ( .A(n9693), .B(n7803), .ZN(n6517) );
  NAND2_X1 U8098 ( .A1(n7990), .A2(n5718), .ZN(n6516) );
  NOR2_X1 U8099 ( .A1(n6517), .A2(n6516), .ZN(n9560) );
  NAND2_X1 U8100 ( .A1(n6517), .A2(n6516), .ZN(n9561) );
  NAND2_X1 U8101 ( .A1(n7989), .A2(n5718), .ZN(n6594) );
  XNOR2_X1 U8102 ( .A(n9703), .B(n7847), .ZN(n6593) );
  XOR2_X1 U8103 ( .A(n6594), .B(n6593), .Z(n6595) );
  XNOR2_X1 U8104 ( .A(n6596), .B(n6595), .ZN(n6523) );
  OAI22_X1 U8105 ( .A1(n7970), .A2(n6611), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9791), .ZN(n6521) );
  OAI22_X1 U8106 ( .A1(n7973), .A2(n6519), .B1(n9571), .B2(n6518), .ZN(n6520)
         );
  AOI211_X1 U8107 ( .C1(n9565), .C2(n9703), .A(n6521), .B(n6520), .ZN(n6522)
         );
  OAI21_X1 U8108 ( .B1(n6523), .B2(n7978), .A(n6522), .ZN(P2_U3219) );
  NAND2_X1 U8109 ( .A1(n8815), .A2(n7538), .ZN(n6526) );
  OR2_X1 U8110 ( .A1(n6629), .A2(n6524), .ZN(n6525) );
  NAND2_X1 U8111 ( .A1(n6526), .A2(n6525), .ZN(n6527) );
  XNOR2_X1 U8112 ( .A(n6527), .B(n7762), .ZN(n6561) );
  NAND2_X1 U8113 ( .A1(n8815), .A2(n6703), .ZN(n6529) );
  INV_X1 U8114 ( .A(n7497), .ZN(n7678) );
  OR2_X1 U8115 ( .A1(n6629), .A2(n6011), .ZN(n6528) );
  NAND2_X1 U8116 ( .A1(n6529), .A2(n6528), .ZN(n6559) );
  XNOR2_X1 U8117 ( .A(n6561), .B(n6559), .ZN(n6533) );
  NAND2_X1 U8118 ( .A1(n6531), .A2(n6530), .ZN(n6532) );
  OAI21_X1 U8119 ( .B1(n6533), .B2(n6532), .A(n6563), .ZN(n6534) );
  NAND2_X1 U8120 ( .A1(n6534), .A2(n8496), .ZN(n6540) );
  OAI22_X1 U8121 ( .A1(n6535), .A2(n8500), .B1(n8487), .B2(n6709), .ZN(n6536)
         );
  AOI211_X1 U8122 ( .C1(n8517), .C2(n6538), .A(n6537), .B(n6536), .ZN(n6539)
         );
  OAI211_X1 U8123 ( .C1(n6629), .C2(n8512), .A(n6540), .B(n6539), .ZN(P1_U3229) );
  NAND2_X1 U8124 ( .A1(n6542), .A2(n6541), .ZN(n6547) );
  INV_X1 U8125 ( .A(n6547), .ZN(n6552) );
  INV_X1 U8126 ( .A(n6543), .ZN(n6546) );
  INV_X1 U8127 ( .A(n6414), .ZN(n6545) );
  AOI21_X1 U8128 ( .B1(n6546), .B2(n6545), .A(n6544), .ZN(n6551) );
  AOI21_X1 U8129 ( .B1(n6549), .B2(n6547), .A(n6551), .ZN(n6548) );
  AOI21_X1 U8130 ( .B1(n6551), .B2(n6549), .A(n6548), .ZN(n6550) );
  AOI21_X1 U8131 ( .B1(n6552), .B2(n6551), .A(n6550), .ZN(n6558) );
  AOI22_X1 U8132 ( .A1(n8503), .A2(n8817), .B1(n8490), .B2(n9501), .ZN(n6557)
         );
  NOR2_X1 U8133 ( .A1(n8500), .A2(n7211), .ZN(n6553) );
  AOI211_X1 U8134 ( .C1(n8517), .C2(n6555), .A(n6554), .B(n6553), .ZN(n6556)
         );
  OAI211_X1 U8135 ( .C1(n6558), .C2(n8519), .A(n6557), .B(n6556), .ZN(P1_U3237) );
  INV_X1 U8136 ( .A(n6559), .ZN(n6560) );
  NAND2_X1 U8137 ( .A1(n6561), .A2(n6560), .ZN(n6562) );
  NAND2_X1 U8138 ( .A1(n6563), .A2(n6562), .ZN(n6697) );
  NAND2_X1 U8139 ( .A1(n6564), .A2(n7642), .ZN(n6567) );
  AOI22_X1 U8140 ( .A1(n8612), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n7566), .B2(
        n6565), .ZN(n6566) );
  NAND2_X1 U8141 ( .A1(n8814), .A2(n4265), .ZN(n6568) );
  OAI21_X1 U8142 ( .B1(n9312), .B2(n6524), .A(n6568), .ZN(n6569) );
  XNOR2_X1 U8143 ( .A(n6569), .B(n7762), .ZN(n6700) );
  OR2_X1 U8144 ( .A1(n9312), .A2(n6011), .ZN(n6571) );
  NAND2_X1 U8145 ( .A1(n8814), .A2(n6703), .ZN(n6570) );
  NAND2_X1 U8146 ( .A1(n6571), .A2(n6570), .ZN(n6698) );
  XNOR2_X1 U8147 ( .A(n6700), .B(n6698), .ZN(n6696) );
  XOR2_X1 U8148 ( .A(n6697), .B(n6696), .Z(n6585) );
  INV_X1 U8149 ( .A(n9312), .ZN(n9239) );
  INV_X1 U8150 ( .A(n9310), .ZN(n6582) );
  NAND2_X1 U8151 ( .A1(n8615), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6579) );
  INV_X1 U8152 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6573) );
  NAND2_X1 U8153 ( .A1(n6574), .A2(n6573), .ZN(n6575) );
  AND2_X1 U8154 ( .A1(n6623), .A2(n6575), .ZN(n6712) );
  NAND2_X1 U8155 ( .A1(n7571), .A2(n6712), .ZN(n6578) );
  NAND2_X1 U8156 ( .A1(n5785), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6577) );
  NAND2_X1 U8157 ( .A1(n7591), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6576) );
  NAND4_X1 U8158 ( .A1(n6579), .A2(n6578), .A3(n6577), .A4(n6576), .ZN(n8813)
         );
  OAI22_X1 U8159 ( .A1(n6739), .A2(n9062), .B1(n6630), .B2(n9060), .ZN(n9233)
         );
  NAND2_X1 U8160 ( .A1(n8419), .A2(n9233), .ZN(n6581) );
  OAI211_X1 U8161 ( .C1(n8485), .C2(n6582), .A(n6581), .B(n6580), .ZN(n6583)
         );
  AOI21_X1 U8162 ( .B1(n9239), .B2(n8490), .A(n6583), .ZN(n6584) );
  OAI21_X1 U8163 ( .B1(n6585), .B2(n8519), .A(n6584), .ZN(P1_U3215) );
  INV_X1 U8164 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7051) );
  INV_X1 U8165 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n6590) );
  MUX2_X1 U8166 ( .A(n7051), .B(n6590), .S(n7244), .Z(n6717) );
  XNOR2_X1 U8167 ( .A(n6717), .B(SI_24_), .ZN(n6715) );
  XNOR2_X1 U8168 ( .A(n6716), .B(n6715), .ZN(n7643) );
  INV_X1 U8169 ( .A(n7643), .ZN(n6591) );
  OAI222_X1 U8170 ( .A1(n4268), .A2(n6591), .B1(P2_U3152), .B2(n6589), .C1(
        n7051), .C2(n8371), .ZN(P2_U3334) );
  OAI222_X1 U8171 ( .A1(P1_U3084), .A2(n6592), .B1(n6728), .B2(n6591), .C1(
        n6590), .C2(n9275), .ZN(P1_U3329) );
  XNOR2_X1 U8172 ( .A(n6776), .B(n7847), .ZN(n6598) );
  NAND2_X1 U8173 ( .A1(n7988), .A2(n5718), .ZN(n6597) );
  XNOR2_X1 U8174 ( .A(n6598), .B(n6597), .ZN(n6650) );
  INV_X1 U8175 ( .A(n6597), .ZN(n6599) );
  NAND2_X1 U8176 ( .A1(n7987), .A2(n5718), .ZN(n6758) );
  NAND2_X1 U8177 ( .A1(n6729), .A2(n7235), .ZN(n6602) );
  AOI22_X1 U8178 ( .A1(n7080), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7079), .B2(
        n6600), .ZN(n6601) );
  XNOR2_X1 U8179 ( .A(n9592), .B(n7847), .ZN(n6757) );
  XOR2_X1 U8180 ( .A(n6758), .B(n6757), .Z(n6760) );
  XNOR2_X1 U8181 ( .A(n6761), .B(n6760), .ZN(n6616) );
  NAND2_X1 U8182 ( .A1(n7222), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6610) );
  OR2_X1 U8183 ( .A1(n7224), .A2(n9385), .ZN(n6609) );
  INV_X1 U8184 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6604) );
  NAND2_X1 U8185 ( .A1(n6605), .A2(n6604), .ZN(n6606) );
  NAND2_X1 U8186 ( .A1(n6904), .A2(n6606), .ZN(n6791) );
  OR2_X1 U8187 ( .A1(n7168), .A2(n6791), .ZN(n6608) );
  INV_X1 U8188 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6792) );
  OR2_X1 U8189 ( .A1(n7228), .A2(n6792), .ZN(n6607) );
  NAND4_X1 U8190 ( .A1(n6610), .A2(n6609), .A3(n6608), .A4(n6607), .ZN(n7986)
         );
  INV_X1 U8191 ( .A(n7986), .ZN(n6781) );
  OAI22_X1 U8192 ( .A1(n6611), .A2(n8249), .B1(n6781), .B2(n8251), .ZN(n9586)
         );
  NAND2_X1 U8193 ( .A1(n9559), .A2(n9586), .ZN(n6612) );
  OAI211_X1 U8194 ( .C1(n9571), .C2(n9588), .A(n6613), .B(n6612), .ZN(n6614)
         );
  AOI21_X1 U8195 ( .B1(n9565), .B2(n9592), .A(n6614), .ZN(n6615) );
  OAI21_X1 U8196 ( .B1(n6616), .B2(n7978), .A(n6615), .ZN(P2_U3226) );
  NAND2_X1 U8197 ( .A1(n6617), .A2(n7642), .ZN(n6619) );
  AOI22_X1 U8198 ( .A1(n8612), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7566), .B2(
        n8828), .ZN(n6618) );
  XNOR2_X1 U8199 ( .A(n6734), .B(n6739), .ZN(n8747) );
  AND2_X1 U8200 ( .A1(n8666), .A2(n8669), .ZN(n6620) );
  NAND2_X1 U8201 ( .A1(n9312), .A2(n8814), .ZN(n8671) );
  NAND2_X1 U8202 ( .A1(n6709), .A2(n9239), .ZN(n8674) );
  OR2_X2 U8203 ( .A1(n9230), .A2(n9231), .ZN(n9227) );
  NAND2_X1 U8204 ( .A1(n9227), .A2(n8671), .ZN(n6738) );
  XOR2_X1 U8205 ( .A(n8747), .B(n6738), .Z(n6644) );
  NAND2_X1 U8206 ( .A1(n8615), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6628) );
  INV_X1 U8207 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6622) );
  NAND2_X1 U8208 ( .A1(n6623), .A2(n6622), .ZN(n6624) );
  AND2_X1 U8209 ( .A1(n6743), .A2(n6624), .ZN(n6882) );
  NAND2_X1 U8210 ( .A1(n7571), .A2(n6882), .ZN(n6627) );
  NAND2_X1 U8211 ( .A1(n5785), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6626) );
  NAND2_X1 U8212 ( .A1(n7591), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6625) );
  NAND4_X1 U8213 ( .A1(n6628), .A2(n6627), .A3(n6626), .A4(n6625), .ZN(n8812)
         );
  OAI22_X1 U8214 ( .A1(n6709), .A2(n9060), .B1(n6965), .B2(n9062), .ZN(n6643)
         );
  NAND2_X1 U8215 ( .A1(n6630), .A2(n6629), .ZN(n6633) );
  AND2_X1 U8216 ( .A1(n6631), .A2(n6633), .ZN(n9221) );
  NAND2_X1 U8217 ( .A1(n9312), .A2(n6709), .ZN(n6632) );
  AND2_X1 U8218 ( .A1(n9221), .A2(n6632), .ZN(n6640) );
  INV_X1 U8219 ( .A(n6632), .ZN(n6639) );
  INV_X1 U8220 ( .A(n6633), .ZN(n6635) );
  OR2_X1 U8221 ( .A1(n6635), .A2(n6634), .ZN(n6638) );
  NAND2_X1 U8222 ( .A1(n8815), .A2(n6636), .ZN(n6637) );
  AND2_X1 U8223 ( .A1(n6638), .A2(n6637), .ZN(n9222) );
  AOI21_X1 U8224 ( .B1(n6641), .B2(n6640), .A(n4820), .ZN(n6733) );
  XNOR2_X1 U8225 ( .A(n6733), .B(n8747), .ZN(n9220) );
  NOR2_X1 U8226 ( .A1(n9220), .A2(n6843), .ZN(n6642) );
  AOI211_X1 U8227 ( .C1(n6644), .C2(n9117), .A(n6643), .B(n6642), .ZN(n9219)
         );
  INV_X1 U8228 ( .A(n6752), .ZN(n6645) );
  AOI21_X1 U8229 ( .B1(n9215), .B2(n9236), .A(n6645), .ZN(n9217) );
  AOI22_X1 U8230 ( .A1(n9030), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n6712), .B2(
        n9309), .ZN(n6646) );
  OAI21_X1 U8231 ( .B1(n9428), .B2(n6734), .A(n6646), .ZN(n6648) );
  NOR2_X1 U8232 ( .A1(n9220), .A2(n9313), .ZN(n6647) );
  AOI211_X1 U8233 ( .C1(n9217), .C2(n9100), .A(n6648), .B(n6647), .ZN(n6649)
         );
  OAI21_X1 U8234 ( .B1(n9219), .B2(n9030), .A(n6649), .ZN(P1_U3280) );
  XOR2_X1 U8235 ( .A(n6651), .B(n6650), .Z(n6658) );
  AOI21_X1 U8236 ( .B1(n9559), .B2(n6653), .A(n6652), .ZN(n6655) );
  NAND2_X1 U8237 ( .A1(n9565), .A2(n6776), .ZN(n6654) );
  OAI211_X1 U8238 ( .C1(n9571), .C2(n6656), .A(n6655), .B(n6654), .ZN(n6657)
         );
  AOI21_X1 U8239 ( .B1(n6658), .B2(n9566), .A(n6657), .ZN(n6659) );
  INV_X1 U8240 ( .A(n6659), .ZN(P2_U3238) );
  INV_X1 U8241 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n9927) );
  NOR2_X1 U8242 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n6660) );
  AOI21_X1 U8243 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n6660), .ZN(n9752) );
  NOR2_X1 U8244 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n6661) );
  AOI21_X1 U8245 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n6661), .ZN(n9755) );
  NOR2_X1 U8246 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n6662) );
  AOI21_X1 U8247 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n6662), .ZN(n9758) );
  NOR2_X1 U8248 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n6663) );
  AOI21_X1 U8249 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n6663), .ZN(n9761) );
  NOR2_X1 U8250 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n6664) );
  AOI21_X1 U8251 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n6664), .ZN(n9764) );
  NOR2_X1 U8252 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n6673) );
  XOR2_X1 U8253 ( .A(n6665), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n9936) );
  NAND2_X1 U8254 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n6671) );
  XNOR2_X1 U8255 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n6666), .ZN(n9934) );
  NAND2_X1 U8256 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n6669) );
  XNOR2_X1 U8257 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n6667), .ZN(n9932) );
  AOI21_X1 U8258 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9746) );
  INV_X1 U8259 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9897) );
  NAND3_X1 U8260 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9748) );
  OAI21_X1 U8261 ( .B1(n9746), .B2(n9897), .A(n9748), .ZN(n9931) );
  NAND2_X1 U8262 ( .A1(n9932), .A2(n9931), .ZN(n6668) );
  NAND2_X1 U8263 ( .A1(n6669), .A2(n6668), .ZN(n9933) );
  NAND2_X1 U8264 ( .A1(n9934), .A2(n9933), .ZN(n6670) );
  NAND2_X1 U8265 ( .A1(n6671), .A2(n6670), .ZN(n9935) );
  NOR2_X1 U8266 ( .A1(n9936), .A2(n9935), .ZN(n6672) );
  NOR2_X1 U8267 ( .A1(n6673), .A2(n6672), .ZN(n6674) );
  NOR2_X1 U8268 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n6674), .ZN(n9923) );
  AND2_X1 U8269 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n6674), .ZN(n9922) );
  NOR2_X1 U8270 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n9922), .ZN(n6675) );
  NOR2_X1 U8271 ( .A1(n9923), .A2(n6675), .ZN(n6676) );
  NAND2_X1 U8272 ( .A1(n6676), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n6678) );
  XOR2_X1 U8273 ( .A(n6676), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n9920) );
  NAND2_X1 U8274 ( .A1(n9920), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n6677) );
  NAND2_X1 U8275 ( .A1(n6678), .A2(n6677), .ZN(n6679) );
  NAND2_X1 U8276 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n6679), .ZN(n6681) );
  XNOR2_X1 U8277 ( .A(n5181), .B(n6679), .ZN(n9919) );
  NAND2_X1 U8278 ( .A1(n9919), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n6680) );
  NAND2_X1 U8279 ( .A1(n6681), .A2(n6680), .ZN(n6682) );
  NAND2_X1 U8280 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n6682), .ZN(n6684) );
  XOR2_X1 U8281 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n6682), .Z(n9921) );
  NAND2_X1 U8282 ( .A1(n9921), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n6683) );
  NAND2_X1 U8283 ( .A1(n6684), .A2(n6683), .ZN(n6685) );
  AND2_X1 U8284 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n6685), .ZN(n6687) );
  XOR2_X1 U8285 ( .A(n6686), .B(n6685), .Z(n9930) );
  NAND2_X1 U8286 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n6688) );
  OAI21_X1 U8287 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n6688), .ZN(n9772) );
  NOR2_X1 U8288 ( .A1(n9773), .A2(n9772), .ZN(n9771) );
  AOI21_X1 U8289 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9771), .ZN(n9770) );
  NAND2_X1 U8290 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n6689) );
  OAI21_X1 U8291 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n6689), .ZN(n9769) );
  NOR2_X1 U8292 ( .A1(n9770), .A2(n9769), .ZN(n9768) );
  AOI21_X1 U8293 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9768), .ZN(n9767) );
  NOR2_X1 U8294 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n6690) );
  AOI21_X1 U8295 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n6690), .ZN(n9766) );
  NAND2_X1 U8296 ( .A1(n9767), .A2(n9766), .ZN(n9765) );
  OAI21_X1 U8297 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9765), .ZN(n9763) );
  NAND2_X1 U8298 ( .A1(n9764), .A2(n9763), .ZN(n9762) );
  OAI21_X1 U8299 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9762), .ZN(n9760) );
  NAND2_X1 U8300 ( .A1(n9761), .A2(n9760), .ZN(n9759) );
  OAI21_X1 U8301 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9759), .ZN(n9757) );
  NAND2_X1 U8302 ( .A1(n9758), .A2(n9757), .ZN(n9756) );
  OAI21_X1 U8303 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9756), .ZN(n9754) );
  NAND2_X1 U8304 ( .A1(n9755), .A2(n9754), .ZN(n9753) );
  OAI21_X1 U8305 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9753), .ZN(n9751) );
  NAND2_X1 U8306 ( .A1(n9752), .A2(n9751), .ZN(n9750) );
  OAI21_X1 U8307 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9750), .ZN(n9926) );
  NOR2_X1 U8308 ( .A1(n9927), .A2(n9926), .ZN(n6691) );
  NAND2_X1 U8309 ( .A1(n9927), .A2(n9926), .ZN(n9925) );
  OAI21_X1 U8310 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n6691), .A(n9925), .ZN(
        n6695) );
  NOR2_X1 U8311 ( .A1(n6693), .A2(n6692), .ZN(n6694) );
  XNOR2_X1 U8312 ( .A(n6695), .B(n6694), .ZN(ADD_1071_U4) );
  INV_X1 U8313 ( .A(n6698), .ZN(n6699) );
  NAND2_X1 U8314 ( .A1(n6700), .A2(n6699), .ZN(n6701) );
  OAI22_X1 U8315 ( .A1(n6734), .A2(n6524), .B1(n6739), .B2(n6011), .ZN(n6702)
         );
  XNOR2_X1 U8316 ( .A(n6702), .B(n7675), .ZN(n6874) );
  OR2_X1 U8317 ( .A1(n6734), .A2(n6011), .ZN(n6705) );
  NAND2_X1 U8318 ( .A1(n8813), .A2(n7484), .ZN(n6704) );
  NAND2_X1 U8319 ( .A1(n6705), .A2(n6704), .ZN(n6873) );
  XNOR2_X1 U8320 ( .A(n6874), .B(n6873), .ZN(n6707) );
  AOI21_X1 U8321 ( .B1(n6706), .B2(n6707), .A(n8519), .ZN(n6708) );
  NAND2_X1 U8322 ( .A1(n6708), .A2(n6876), .ZN(n6714) );
  NOR2_X1 U8323 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6573), .ZN(n6711) );
  OAI22_X1 U8324 ( .A1(n6709), .A2(n8500), .B1(n8487), .B2(n6965), .ZN(n6710)
         );
  AOI211_X1 U8325 ( .C1(n8517), .C2(n6712), .A(n6711), .B(n6710), .ZN(n6713)
         );
  OAI211_X1 U8326 ( .C1(n6734), .C2(n8512), .A(n6714), .B(n6713), .ZN(P1_U3234) );
  INV_X1 U8327 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7131) );
  INV_X1 U8328 ( .A(n6717), .ZN(n6718) );
  NAND2_X1 U8329 ( .A1(n6718), .A2(SI_24_), .ZN(n6719) );
  NAND2_X1 U8330 ( .A1(n6720), .A2(n6719), .ZN(n6834) );
  INV_X1 U8331 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n9808) );
  MUX2_X1 U8332 ( .A(n7131), .B(n9808), .S(n7244), .Z(n6722) );
  INV_X1 U8333 ( .A(SI_25_), .ZN(n6721) );
  NAND2_X1 U8334 ( .A1(n6722), .A2(n6721), .ZN(n6832) );
  INV_X1 U8335 ( .A(n6722), .ZN(n6723) );
  NAND2_X1 U8336 ( .A1(n6723), .A2(SI_25_), .ZN(n6724) );
  NAND2_X1 U8337 ( .A1(n6832), .A2(n6724), .ZN(n6833) );
  INV_X1 U8338 ( .A(n7661), .ZN(n6727) );
  OAI222_X1 U8339 ( .A1(n9275), .A2(n9808), .B1(n6728), .B2(n6727), .C1(
        P1_U3084), .C2(n6726), .ZN(P1_U3328) );
  NAND2_X1 U8340 ( .A1(n6729), .A2(n7642), .ZN(n6732) );
  AOI22_X1 U8341 ( .A1(n8612), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n7566), .B2(
        n6730), .ZN(n6731) );
  NAND2_X1 U8342 ( .A1(n9400), .A2(n6965), .ZN(n8539) );
  INV_X1 U8343 ( .A(n6733), .ZN(n6736) );
  AOI21_X1 U8344 ( .B1(n8748), .B2(n6737), .A(n6799), .ZN(n9404) );
  INV_X1 U8345 ( .A(n9404), .ZN(n9402) );
  NAND2_X1 U8346 ( .A1(n9215), .A2(n6739), .ZN(n8536) );
  NAND2_X1 U8347 ( .A1(n6738), .A2(n8536), .ZN(n6816) );
  OR2_X1 U8348 ( .A1(n9215), .A2(n6739), .ZN(n6815) );
  NAND2_X1 U8349 ( .A1(n6816), .A2(n6815), .ZN(n6740) );
  XNOR2_X1 U8350 ( .A(n6740), .B(n8748), .ZN(n6751) );
  NAND2_X1 U8351 ( .A1(n8615), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6748) );
  INV_X1 U8352 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6742) );
  NAND2_X1 U8353 ( .A1(n6743), .A2(n6742), .ZN(n6744) );
  AND2_X1 U8354 ( .A1(n6806), .A2(n6744), .ZN(n6968) );
  NAND2_X1 U8355 ( .A1(n7571), .A2(n6968), .ZN(n6747) );
  NAND2_X1 U8356 ( .A1(n5785), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6746) );
  NAND2_X1 U8357 ( .A1(n7591), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6745) );
  NAND4_X1 U8358 ( .A1(n6748), .A2(n6747), .A3(n6746), .A4(n6745), .ZN(n8811)
         );
  NAND2_X1 U8359 ( .A1(n8811), .A2(n9114), .ZN(n6750) );
  NAND2_X1 U8360 ( .A1(n8813), .A2(n9112), .ZN(n6749) );
  AND2_X1 U8361 ( .A1(n6750), .A2(n6749), .ZN(n6885) );
  OAI21_X1 U8362 ( .B1(n6751), .B2(n9229), .A(n6885), .ZN(n9398) );
  AOI211_X1 U8363 ( .C1(n9400), .C2(n6752), .A(n9519), .B(n6847), .ZN(n9399)
         );
  NAND2_X1 U8364 ( .A1(n9399), .A2(n9317), .ZN(n6754) );
  AOI22_X1 U8365 ( .A1(n9030), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n6882), .B2(
        n9309), .ZN(n6753) );
  OAI211_X1 U8366 ( .C1(n4738), .C2(n9428), .A(n6754), .B(n6753), .ZN(n6755)
         );
  AOI21_X1 U8367 ( .B1(n9070), .B2(n9398), .A(n6755), .ZN(n6756) );
  OAI21_X1 U8368 ( .B1(n9402), .B2(n9121), .A(n6756), .ZN(P1_U3279) );
  INV_X1 U8369 ( .A(n6757), .ZN(n6759) );
  NAND2_X1 U8370 ( .A1(n6800), .A2(n7235), .ZN(n6764) );
  AOI22_X1 U8371 ( .A1(n7080), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7079), .B2(
        n6762), .ZN(n6763) );
  XNOR2_X1 U8372 ( .A(n6972), .B(n7847), .ZN(n6896) );
  NAND2_X1 U8373 ( .A1(n7986), .A2(n5718), .ZN(n6894) );
  XNOR2_X1 U8374 ( .A(n6896), .B(n6894), .ZN(n6897) );
  XNOR2_X1 U8375 ( .A(n6898), .B(n6897), .ZN(n6775) );
  INV_X1 U8376 ( .A(n5577), .ZN(n7127) );
  NAND2_X1 U8377 ( .A1(n7127), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6770) );
  OR2_X1 U8378 ( .A1(n7224), .A2(n6765), .ZN(n6769) );
  INV_X1 U8379 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n6766) );
  OR2_X1 U8380 ( .A1(n5579), .A2(n6766), .ZN(n6768) );
  INV_X1 U8381 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n6903) );
  XNOR2_X1 U8382 ( .A(n6904), .B(n6903), .ZN(n9350) );
  OR2_X1 U8383 ( .A1(n7168), .A2(n9350), .ZN(n6767) );
  NAND4_X1 U8384 ( .A1(n6770), .A2(n6769), .A3(n6768), .A4(n6767), .ZN(n7985)
         );
  OAI21_X1 U8385 ( .B1(n7970), .B2(n7972), .A(n6771), .ZN(n6773) );
  INV_X1 U8386 ( .A(n7987), .ZN(n6787) );
  OAI22_X1 U8387 ( .A1(n7973), .A2(n6787), .B1(n9571), .B2(n6791), .ZN(n6772)
         );
  AOI211_X1 U8388 ( .C1(n9565), .C2(n6972), .A(n6773), .B(n6772), .ZN(n6774)
         );
  OAI21_X1 U8389 ( .B1(n6775), .B2(n7978), .A(n6774), .ZN(P2_U3236) );
  NAND2_X1 U8390 ( .A1(n6776), .A2(n7988), .ZN(n6777) );
  OR2_X1 U8391 ( .A1(n9592), .A2(n6787), .ZN(n7318) );
  NAND2_X1 U8392 ( .A1(n9592), .A2(n6787), .ZN(n7321) );
  OR2_X1 U8393 ( .A1(n9592), .A2(n7987), .ZN(n6780) );
  OR2_X1 U8394 ( .A1(n6972), .A2(n6781), .ZN(n7327) );
  NAND2_X1 U8395 ( .A1(n6972), .A2(n6781), .ZN(n9343) );
  NAND2_X1 U8396 ( .A1(n6782), .A2(n7414), .ZN(n6783) );
  NAND2_X1 U8397 ( .A1(n4792), .A2(n6783), .ZN(n9379) );
  AND2_X1 U8398 ( .A1(n7318), .A2(n9583), .ZN(n7323) );
  NAND2_X1 U8399 ( .A1(n6785), .A2(n7321), .ZN(n6786) );
  NAND2_X1 U8400 ( .A1(n6786), .A2(n7414), .ZN(n9344) );
  OAI21_X1 U8401 ( .B1(n7414), .B2(n6786), .A(n9344), .ZN(n6789) );
  OAI22_X1 U8402 ( .A1(n6787), .A2(n8249), .B1(n7972), .B2(n8251), .ZN(n6788)
         );
  AOI21_X1 U8403 ( .B1(n6789), .B2(n9619), .A(n6788), .ZN(n6790) );
  OAI21_X1 U8404 ( .B1(n9379), .B2(n9691), .A(n6790), .ZN(n9382) );
  NAND2_X1 U8405 ( .A1(n9382), .A2(n8265), .ZN(n6797) );
  OAI22_X1 U8406 ( .A1(n8265), .A2(n6792), .B1(n6791), .B2(n8238), .ZN(n6795)
         );
  INV_X1 U8407 ( .A(n9592), .ZN(n9720) );
  INV_X1 U8408 ( .A(n6972), .ZN(n9380) );
  OR2_X1 U8409 ( .A1(n9596), .A2(n9380), .ZN(n6793) );
  NAND2_X1 U8410 ( .A1(n9356), .A2(n6793), .ZN(n9381) );
  NOR2_X1 U8411 ( .A1(n9381), .A2(n8078), .ZN(n6794) );
  AOI211_X1 U8412 ( .C1(n9591), .C2(n6972), .A(n6795), .B(n6794), .ZN(n6796)
         );
  OAI211_X1 U8413 ( .C1(n9379), .C2(n6798), .A(n6797), .B(n6796), .ZN(P2_U3283) );
  NAND2_X1 U8414 ( .A1(n6800), .A2(n7642), .ZN(n6802) );
  AOI22_X1 U8415 ( .A1(n8612), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n7566), .B2(
        n6861), .ZN(n6801) );
  INV_X1 U8416 ( .A(n8811), .ZN(n6818) );
  NAND2_X1 U8417 ( .A1(n6889), .A2(n7642), .ZN(n6804) );
  AOI22_X1 U8418 ( .A1(n8612), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n9412), .B2(
        n7566), .ZN(n6803) );
  NAND2_X1 U8419 ( .A1(n8615), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6811) );
  INV_X1 U8420 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6805) );
  NAND2_X1 U8421 ( .A1(n6806), .A2(n6805), .ZN(n6807) );
  AND2_X1 U8422 ( .A1(n6821), .A2(n6807), .ZN(n8390) );
  NAND2_X1 U8423 ( .A1(n7571), .A2(n8390), .ZN(n6810) );
  NAND2_X1 U8424 ( .A1(n5785), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6809) );
  NAND2_X1 U8425 ( .A1(n7591), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6808) );
  NAND4_X1 U8426 ( .A1(n6811), .A2(n6810), .A3(n6809), .A4(n6808), .ZN(n8810)
         );
  OR2_X1 U8427 ( .A1(n9205), .A2(n6964), .ZN(n8547) );
  NAND2_X1 U8428 ( .A1(n9205), .A2(n6964), .ZN(n8641) );
  NAND2_X1 U8429 ( .A1(n8547), .A2(n8641), .ZN(n8752) );
  XNOR2_X1 U8430 ( .A(n6927), .B(n8752), .ZN(n9209) );
  INV_X1 U8431 ( .A(n6848), .ZN(n6813) );
  INV_X1 U8432 ( .A(n6937), .ZN(n6812) );
  AOI211_X1 U8433 ( .C1(n9205), .C2(n6813), .A(n9519), .B(n6812), .ZN(n9204)
         );
  AOI22_X1 U8434 ( .A1(n9030), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8390), .B2(
        n9309), .ZN(n6814) );
  OAI21_X1 U8435 ( .B1(n6928), .B2(n9428), .A(n6814), .ZN(n6830) );
  AND2_X1 U8436 ( .A1(n8537), .A2(n6815), .ZN(n8678) );
  NAND2_X1 U8437 ( .A1(n6816), .A2(n8678), .ZN(n6817) );
  NAND2_X1 U8438 ( .A1(n6817), .A2(n8539), .ZN(n6842) );
  OR2_X1 U8439 ( .A1(n9210), .A2(n6818), .ZN(n8546) );
  NAND2_X1 U8440 ( .A1(n9210), .A2(n6818), .ZN(n8679) );
  NAND2_X1 U8441 ( .A1(n6842), .A2(n8541), .ZN(n6819) );
  NAND2_X1 U8442 ( .A1(n6819), .A2(n8679), .ZN(n6820) );
  AOI21_X1 U8443 ( .B1(n6820), .B2(n8752), .A(n9229), .ZN(n6828) );
  NAND2_X1 U8444 ( .A1(n8615), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6826) );
  INV_X1 U8445 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8509) );
  NAND2_X1 U8446 ( .A1(n6821), .A2(n8509), .ZN(n6822) );
  AND2_X1 U8447 ( .A1(n6941), .A2(n6822), .ZN(n8516) );
  NAND2_X1 U8448 ( .A1(n7571), .A2(n8516), .ZN(n6825) );
  NAND2_X1 U8449 ( .A1(n7591), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6824) );
  NAND2_X1 U8450 ( .A1(n5785), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6823) );
  NAND4_X1 U8451 ( .A1(n6826), .A2(n6825), .A3(n6824), .A4(n6823), .ZN(n9113)
         );
  AOI22_X1 U8452 ( .A1(n9112), .A2(n8811), .B1(n9113), .B2(n9114), .ZN(n8392)
         );
  INV_X1 U8453 ( .A(n8392), .ZN(n6827) );
  AOI21_X1 U8454 ( .B1(n6828), .B2(n6939), .A(n6827), .ZN(n9207) );
  NOR2_X1 U8455 ( .A1(n9207), .A2(n9030), .ZN(n6829) );
  AOI211_X1 U8456 ( .C1(n9317), .C2(n9204), .A(n6830), .B(n6829), .ZN(n6831)
         );
  OAI21_X1 U8457 ( .B1(n9209), .B2(n9121), .A(n6831), .ZN(P1_U3277) );
  INV_X1 U8458 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7142) );
  INV_X1 U8459 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n6840) );
  MUX2_X1 U8460 ( .A(n7142), .B(n6840), .S(n7244), .Z(n6836) );
  INV_X1 U8461 ( .A(SI_26_), .ZN(n6835) );
  NAND2_X1 U8462 ( .A1(n6836), .A2(n6835), .ZN(n6919) );
  INV_X1 U8463 ( .A(n6836), .ZN(n6837) );
  NAND2_X1 U8464 ( .A1(n6837), .A2(SI_26_), .ZN(n6838) );
  AND2_X1 U8465 ( .A1(n6919), .A2(n6838), .ZN(n6917) );
  INV_X1 U8466 ( .A(n7679), .ZN(n6841) );
  OAI222_X1 U8467 ( .A1(n4268), .A2(n6841), .B1(P2_U3152), .B2(n6839), .C1(
        n7142), .C2(n8371), .ZN(P2_U3332) );
  OAI222_X1 U8468 ( .A1(P1_U3084), .A2(n5370), .B1(n9273), .B2(n6841), .C1(
        n6840), .C2(n9275), .ZN(P1_U3327) );
  XNOR2_X1 U8469 ( .A(n6842), .B(n8541), .ZN(n6846) );
  OAI22_X1 U8470 ( .A1(n6965), .A2(n9060), .B1(n6964), .B2(n9062), .ZN(n6845)
         );
  XNOR2_X1 U8471 ( .A(n4337), .B(n8541), .ZN(n9214) );
  NOR2_X1 U8472 ( .A1(n9214), .A2(n6843), .ZN(n6844) );
  AOI211_X1 U8473 ( .C1(n6846), .C2(n9117), .A(n6845), .B(n6844), .ZN(n9213)
         );
  AOI21_X1 U8474 ( .B1(n9210), .B2(n4740), .A(n6848), .ZN(n9211) );
  AOI22_X1 U8475 ( .A1(n9321), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n6968), .B2(
        n9309), .ZN(n6849) );
  OAI21_X1 U8476 ( .B1(n6971), .B2(n9428), .A(n6849), .ZN(n6851) );
  NOR2_X1 U8477 ( .A1(n9214), .A2(n9313), .ZN(n6850) );
  AOI211_X1 U8478 ( .C1(n9211), .C2(n9100), .A(n6851), .B(n6850), .ZN(n6852)
         );
  OAI21_X1 U8479 ( .B1(n9213), .B2(n9321), .A(n6852), .ZN(P1_U3278) );
  NAND2_X1 U8480 ( .A1(n6854), .A2(n6858), .ZN(n6855) );
  INV_X1 U8481 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9415) );
  NAND2_X1 U8482 ( .A1(n9416), .A2(n9415), .ZN(n9414) );
  NAND2_X1 U8483 ( .A1(n6855), .A2(n9414), .ZN(n7007) );
  XNOR2_X1 U8484 ( .A(n7007), .B(n7014), .ZN(n6857) );
  INV_X1 U8485 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n6856) );
  NOR2_X1 U8486 ( .A1(n6856), .A2(n6857), .ZN(n7008) );
  AOI211_X1 U8487 ( .C1(n6857), .C2(n6856), .A(n7008), .B(n8861), .ZN(n6868)
         );
  INV_X1 U8488 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n6863) );
  INV_X1 U8489 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6859) );
  AOI22_X1 U8490 ( .A1(n9412), .A2(P1_REG1_REG_14__SCAN_IN), .B1(n6859), .B2(
        n6858), .ZN(n9419) );
  OAI21_X1 U8491 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n6861), .A(n6860), .ZN(
        n9418) );
  NAND2_X1 U8492 ( .A1(n9419), .A2(n9418), .ZN(n9417) );
  AOI211_X1 U8493 ( .C1(n6863), .C2(n6862), .A(n7015), .B(n8855), .ZN(n6867)
         );
  NAND2_X1 U8494 ( .A1(n8864), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n6865) );
  NAND2_X1 U8495 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3084), .ZN(n6864) );
  OAI211_X1 U8496 ( .C1(n4363), .C2(n7014), .A(n6865), .B(n6864), .ZN(n6866)
         );
  OR3_X1 U8497 ( .A1(n6868), .A2(n6867), .A3(n6866), .ZN(P1_U3256) );
  NAND2_X1 U8498 ( .A1(n9400), .A2(n4263), .ZN(n6870) );
  NAND2_X1 U8499 ( .A1(n8812), .A2(n7485), .ZN(n6869) );
  NAND2_X1 U8500 ( .A1(n6870), .A2(n6869), .ZN(n6871) );
  XNOR2_X1 U8501 ( .A(n6871), .B(n7762), .ZN(n6954) );
  AND2_X1 U8502 ( .A1(n8812), .A2(n6703), .ZN(n6872) );
  AOI21_X1 U8503 ( .B1(n9400), .B2(n7485), .A(n6872), .ZN(n6953) );
  XNOR2_X1 U8504 ( .A(n6954), .B(n6953), .ZN(n6881) );
  NAND2_X1 U8505 ( .A1(n6874), .A2(n6873), .ZN(n6875) );
  INV_X1 U8506 ( .A(n6881), .ZN(n6877) );
  INV_X1 U8507 ( .A(n6956), .ZN(n6879) );
  AOI21_X1 U8508 ( .B1(n6881), .B2(n6880), .A(n6879), .ZN(n6888) );
  NAND2_X1 U8509 ( .A1(n8517), .A2(n6882), .ZN(n6884) );
  OAI211_X1 U8510 ( .C1(n8511), .C2(n6885), .A(n6884), .B(n6883), .ZN(n6886)
         );
  AOI21_X1 U8511 ( .B1(n9400), .B2(n8490), .A(n6886), .ZN(n6887) );
  OAI21_X1 U8512 ( .B1(n6888), .B2(n8519), .A(n6887), .ZN(P1_U3222) );
  NAND2_X1 U8513 ( .A1(n6889), .A2(n7235), .ZN(n6891) );
  AOI22_X1 U8514 ( .A1(n8000), .A2(n7079), .B1(n7080), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n6890) );
  INV_X1 U8515 ( .A(n9352), .ZN(n9376) );
  AND2_X1 U8516 ( .A1(n7985), .A2(n5718), .ZN(n6893) );
  XNOR2_X1 U8517 ( .A(n9352), .B(n7847), .ZN(n6892) );
  NOR2_X1 U8518 ( .A1(n6892), .A2(n6893), .ZN(n7800) );
  AOI21_X1 U8519 ( .B1(n6893), .B2(n6892), .A(n7800), .ZN(n6900) );
  INV_X1 U8520 ( .A(n6894), .ZN(n6895) );
  NAND2_X1 U8521 ( .A1(n6899), .A2(n6900), .ZN(n7802) );
  OAI21_X1 U8522 ( .B1(n6900), .B2(n6899), .A(n7802), .ZN(n6901) );
  NAND2_X1 U8523 ( .A1(n6901), .A2(n9566), .ZN(n6916) );
  NAND2_X1 U8524 ( .A1(n5576), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6909) );
  NAND2_X1 U8525 ( .A1(n7222), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6908) );
  INV_X1 U8526 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6902) );
  OAI21_X1 U8527 ( .B1(n6904), .B2(n6903), .A(n6902), .ZN(n6905) );
  NAND2_X1 U8528 ( .A1(n6905), .A2(n6981), .ZN(n7971) );
  OR2_X1 U8529 ( .A1(n7168), .A2(n7971), .ZN(n6907) );
  INV_X1 U8530 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n6994) );
  OR2_X1 U8531 ( .A1(n7228), .A2(n6994), .ZN(n6906) );
  NAND4_X1 U8532 ( .A1(n6909), .A2(n6908), .A3(n6907), .A4(n6906), .ZN(n7984)
         );
  NAND2_X1 U8533 ( .A1(n7984), .A2(n9621), .ZN(n6911) );
  NAND2_X1 U8534 ( .A1(n7986), .A2(n9624), .ZN(n6910) );
  NAND2_X1 U8535 ( .A1(n6911), .A2(n6910), .ZN(n9348) );
  INV_X1 U8536 ( .A(n6912), .ZN(n6914) );
  NOR2_X1 U8537 ( .A1(n9571), .A2(n9350), .ZN(n6913) );
  AOI211_X1 U8538 ( .C1(n9559), .C2(n9348), .A(n6914), .B(n6913), .ZN(n6915)
         );
  OAI211_X1 U8539 ( .C1(n9376), .C2(n7950), .A(n6916), .B(n6915), .ZN(P2_U3217) );
  INV_X1 U8540 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7154) );
  INV_X1 U8541 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n6920) );
  MUX2_X1 U8542 ( .A(n7154), .B(n6920), .S(n7244), .Z(n6922) );
  INV_X1 U8543 ( .A(SI_27_), .ZN(n6921) );
  NAND2_X1 U8544 ( .A1(n6922), .A2(n6921), .ZN(n7002) );
  INV_X1 U8545 ( .A(n6922), .ZN(n6923) );
  NAND2_X1 U8546 ( .A1(n6923), .A2(SI_27_), .ZN(n6924) );
  AND2_X1 U8547 ( .A1(n7002), .A2(n6924), .ZN(n7000) );
  INV_X1 U8548 ( .A(n7460), .ZN(n6952) );
  AOI21_X1 U8549 ( .B1(n9265), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n6925), .ZN(
        n6926) );
  OAI21_X1 U8550 ( .B1(n6952), .B2(n9273), .A(n6926), .ZN(P1_U3326) );
  INV_X1 U8551 ( .A(n6927), .ZN(n6931) );
  NAND2_X1 U8552 ( .A1(n9205), .A2(n8810), .ZN(n6930) );
  AOI21_X1 U8553 ( .B1(n6931), .B2(n6930), .A(n6929), .ZN(n7723) );
  NAND2_X1 U8554 ( .A1(n6974), .A2(n7642), .ZN(n6935) );
  OAI22_X1 U8555 ( .A1(n7014), .A2(n6932), .B1(n6347), .B2(n9871), .ZN(n6933)
         );
  INV_X1 U8556 ( .A(n6933), .ZN(n6934) );
  XNOR2_X1 U8557 ( .A(n9199), .B(n8436), .ZN(n8755) );
  XNOR2_X1 U8558 ( .A(n7723), .B(n8755), .ZN(n9203) );
  INV_X1 U8559 ( .A(n9105), .ZN(n6936) );
  AOI21_X1 U8560 ( .B1(n9199), .B2(n6937), .A(n6936), .ZN(n9200) );
  INV_X1 U8561 ( .A(n9199), .ZN(n8513) );
  AOI22_X1 U8562 ( .A1(n9030), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8516), .B2(
        n9309), .ZN(n6938) );
  OAI21_X1 U8563 ( .B1(n8513), .B2(n9428), .A(n6938), .ZN(n6950) );
  XNOR2_X1 U8564 ( .A(n7739), .B(n8755), .ZN(n6948) );
  NAND2_X1 U8565 ( .A1(n8615), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6946) );
  INV_X1 U8566 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9869) );
  NAND2_X1 U8567 ( .A1(n6941), .A2(n9869), .ZN(n6942) );
  AND2_X1 U8568 ( .A1(n7528), .A2(n6942), .ZN(n9106) );
  NAND2_X1 U8569 ( .A1(n7571), .A2(n9106), .ZN(n6945) );
  NAND2_X1 U8570 ( .A1(n5785), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6944) );
  NAND2_X1 U8571 ( .A1(n7591), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6943) );
  NAND4_X1 U8572 ( .A1(n6946), .A2(n6945), .A3(n6944), .A4(n6943), .ZN(n9095)
         );
  AOI22_X1 U8573 ( .A1(n9112), .A2(n8810), .B1(n9095), .B2(n9114), .ZN(n8510)
         );
  INV_X1 U8574 ( .A(n8510), .ZN(n6947) );
  AOI21_X1 U8575 ( .B1(n6948), .B2(n9117), .A(n6947), .ZN(n9202) );
  NOR2_X1 U8576 ( .A1(n9202), .A2(n9433), .ZN(n6949) );
  AOI211_X1 U8577 ( .C1(n9200), .C2(n9100), .A(n6950), .B(n6949), .ZN(n6951)
         );
  OAI21_X1 U8578 ( .B1(n9203), .B2(n9121), .A(n6951), .ZN(P1_U3276) );
  OAI222_X1 U8579 ( .A1(n4268), .A2(n6952), .B1(n5186), .B2(P2_U3152), .C1(
        n7154), .C2(n8371), .ZN(P2_U3331) );
  NAND2_X1 U8580 ( .A1(n6954), .A2(n6953), .ZN(n6955) );
  AND2_X1 U8581 ( .A1(n8811), .A2(n6703), .ZN(n6958) );
  AOI21_X1 U8582 ( .B1(n9210), .B2(n7485), .A(n6958), .ZN(n7486) );
  NAND2_X1 U8583 ( .A1(n9210), .A2(n4263), .ZN(n6960) );
  NAND2_X1 U8584 ( .A1(n8811), .A2(n7497), .ZN(n6959) );
  NAND2_X1 U8585 ( .A1(n6960), .A2(n6959), .ZN(n6961) );
  XNOR2_X1 U8586 ( .A(n6961), .B(n7762), .ZN(n7487) );
  XOR2_X1 U8587 ( .A(n7486), .B(n7487), .Z(n6962) );
  XNOR2_X1 U8588 ( .A(n7490), .B(n6962), .ZN(n6963) );
  NAND2_X1 U8589 ( .A1(n6963), .A2(n8496), .ZN(n6970) );
  OAI22_X1 U8590 ( .A1(n6965), .A2(n8500), .B1(n8487), .B2(n6964), .ZN(n6966)
         );
  AOI211_X1 U8591 ( .C1(n8517), .C2(n6968), .A(n6967), .B(n6966), .ZN(n6969)
         );
  OAI211_X1 U8592 ( .C1(n6971), .C2(n8512), .A(n6970), .B(n6969), .ZN(P1_U3232) );
  NAND2_X1 U8593 ( .A1(n9352), .A2(n7972), .ZN(n7330) );
  NAND2_X1 U8594 ( .A1(n7329), .A2(n7330), .ZN(n9354) );
  NAND2_X1 U8595 ( .A1(n9353), .A2(n6973), .ZN(n7057) );
  NAND2_X1 U8596 ( .A1(n6974), .A2(n7235), .ZN(n6979) );
  OAI22_X1 U8597 ( .A1(n8019), .A2(n6976), .B1(n7248), .B2(n6975), .ZN(n6977)
         );
  INV_X1 U8598 ( .A(n6977), .ZN(n6978) );
  NAND2_X1 U8599 ( .A1(n7976), .A2(n7915), .ZN(n7333) );
  NAND2_X1 U8600 ( .A1(n7334), .A2(n7333), .ZN(n7416) );
  XNOR2_X1 U8601 ( .A(n7057), .B(n7416), .ZN(n9372) );
  INV_X1 U8602 ( .A(n9372), .ZN(n6999) );
  NAND2_X1 U8603 ( .A1(n7222), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6988) );
  INV_X1 U8604 ( .A(n6981), .ZN(n6980) );
  NAND2_X1 U8605 ( .A1(n6980), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n7062) );
  INV_X1 U8606 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9805) );
  NAND2_X1 U8607 ( .A1(n6981), .A2(n9805), .ZN(n6982) );
  NAND2_X1 U8608 ( .A1(n7062), .A2(n6982), .ZN(n9330) );
  OR2_X1 U8609 ( .A1(n7168), .A2(n9330), .ZN(n6987) );
  INV_X1 U8610 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n6983) );
  OR2_X1 U8611 ( .A1(n7224), .A2(n6983), .ZN(n6986) );
  INV_X1 U8612 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n6984) );
  OR2_X1 U8613 ( .A1(n7228), .A2(n6984), .ZN(n6985) );
  NAND4_X1 U8614 ( .A1(n6988), .A2(n6987), .A3(n6986), .A4(n6985), .ZN(n7983)
         );
  INV_X1 U8615 ( .A(n9343), .ZN(n6989) );
  NOR2_X1 U8616 ( .A1(n9354), .A2(n6989), .ZN(n6990) );
  INV_X1 U8617 ( .A(n7416), .ZN(n7332) );
  XNOR2_X1 U8618 ( .A(n7180), .B(n7332), .ZN(n6991) );
  OAI222_X1 U8619 ( .A1(n8249), .A2(n7972), .B1(n8251), .B2(n8248), .C1(n9345), 
        .C2(n6991), .ZN(n9371) );
  INV_X1 U8620 ( .A(n7976), .ZN(n9368) );
  INV_X1 U8621 ( .A(n9357), .ZN(n6993) );
  INV_X1 U8622 ( .A(n9335), .ZN(n6992) );
  OAI21_X1 U8623 ( .B1(n9368), .B2(n6993), .A(n6992), .ZN(n9369) );
  OAI22_X1 U8624 ( .A1(n8265), .A2(n6994), .B1(n7971), .B2(n8238), .ZN(n6995)
         );
  AOI21_X1 U8625 ( .B1(n7976), .B2(n9591), .A(n6995), .ZN(n6996) );
  OAI21_X1 U8626 ( .B1(n9369), .B2(n8078), .A(n6996), .ZN(n6997) );
  AOI21_X1 U8627 ( .B1(n9371), .B2(n8265), .A(n6997), .ZN(n6998) );
  OAI21_X1 U8628 ( .B1(n6999), .B2(n8254), .A(n6998), .ZN(P2_U3281) );
  NAND2_X1 U8629 ( .A1(n7003), .A2(n7002), .ZN(n7035) );
  INV_X1 U8630 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7163) );
  INV_X1 U8631 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7004) );
  MUX2_X1 U8632 ( .A(n7163), .B(n7004), .S(n7244), .Z(n7037) );
  XNOR2_X1 U8633 ( .A(n7037), .B(SI_28_), .ZN(n7034) );
  INV_X1 U8634 ( .A(n7757), .ZN(n7041) );
  AOI21_X1 U8635 ( .B1(n9265), .B2(P2_DATAO_REG_28__SCAN_IN), .A(n7005), .ZN(
        n7006) );
  OAI21_X1 U8636 ( .B1(n7041), .B2(n9273), .A(n7006), .ZN(P1_U3325) );
  NOR2_X1 U8637 ( .A1(n7014), .A2(n7007), .ZN(n7009) );
  NAND2_X1 U8638 ( .A1(n8844), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7010) );
  OAI21_X1 U8639 ( .B1(n8844), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7010), .ZN(
        n7011) );
  AOI211_X1 U8640 ( .C1(n7012), .C2(n7011), .A(n8843), .B(n8861), .ZN(n7025)
         );
  NOR2_X1 U8641 ( .A1(n7014), .A2(n7013), .ZN(n7016) );
  INV_X1 U8642 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7018) );
  AOI22_X1 U8643 ( .A1(n8844), .A2(n7018), .B1(P1_REG1_REG_16__SCAN_IN), .B2(
        n7017), .ZN(n7019) );
  NOR2_X1 U8644 ( .A1(n7020), .A2(n7019), .ZN(n8837) );
  AOI211_X1 U8645 ( .C1(n7020), .C2(n7019), .A(n8837), .B(n8855), .ZN(n7024)
         );
  INV_X1 U8646 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7022) );
  NOR2_X1 U8647 ( .A1(n9869), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8438) );
  AOI21_X1 U8648 ( .B1(n9413), .B2(n8844), .A(n8438), .ZN(n7021) );
  OAI21_X1 U8649 ( .B1(n9426), .B2(n7022), .A(n7021), .ZN(n7023) );
  OR3_X1 U8650 ( .A1(n7025), .A2(n7024), .A3(n7023), .ZN(P1_U3257) );
  OAI21_X1 U8651 ( .B1(n7028), .B2(n7027), .A(n7026), .ZN(n7029) );
  AOI22_X1 U8652 ( .A1(n7029), .A2(n9566), .B1(n7869), .B2(n7994), .ZN(n7032)
         );
  AOI22_X1 U8653 ( .A1(n9565), .A2(n9649), .B1(n7030), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n7031) );
  OAI211_X1 U8654 ( .C1(n8257), .C2(n7973), .A(n7032), .B(n7031), .ZN(P2_U3239) );
  INV_X1 U8655 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7219) );
  NAND2_X1 U8656 ( .A1(n7035), .A2(n7034), .ZN(n7039) );
  INV_X1 U8657 ( .A(SI_28_), .ZN(n7036) );
  NAND2_X1 U8658 ( .A1(n7037), .A2(n7036), .ZN(n7038) );
  INV_X1 U8659 ( .A(SI_29_), .ZN(n7232) );
  MUX2_X1 U8660 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n7244), .Z(n7233) );
  MUX2_X1 U8661 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n7244), .Z(n7240) );
  INV_X1 U8662 ( .A(n8611), .ZN(n9270) );
  OAI222_X1 U8663 ( .A1(n4268), .A2(n7041), .B1(n5185), .B2(P2_U3152), .C1(
        n7163), .C2(n8371), .ZN(P2_U3330) );
  INV_X1 U8664 ( .A(n7062), .ZN(n7042) );
  NAND2_X1 U8665 ( .A1(n7042), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n7071) );
  INV_X1 U8666 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9830) );
  INV_X1 U8667 ( .A(n7095), .ZN(n7044) );
  AND2_X1 U8668 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_REG3_REG_20__SCAN_IN), 
        .ZN(n7043) );
  NAND2_X1 U8669 ( .A1(n7044), .A2(n7043), .ZN(n7105) );
  INV_X1 U8670 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n7891) );
  INV_X1 U8671 ( .A(n7124), .ZN(n7046) );
  AND2_X1 U8672 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(P2_REG3_REG_22__SCAN_IN), 
        .ZN(n7045) );
  NAND2_X1 U8673 ( .A1(n7046), .A2(n7045), .ZN(n7125) );
  INV_X1 U8674 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n7928) );
  NAND2_X1 U8675 ( .A1(n7125), .A2(n7928), .ZN(n7047) );
  NAND2_X1 U8676 ( .A1(n7134), .A2(n7047), .ZN(n8135) );
  OR2_X1 U8677 ( .A1(n8135), .A2(n7168), .ZN(n7050) );
  AOI22_X1 U8678 ( .A1(n7127), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n5576), .B2(
        P2_REG1_REG_24__SCAN_IN), .ZN(n7049) );
  NAND2_X1 U8679 ( .A1(n7222), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n7048) );
  NAND2_X1 U8680 ( .A1(n7643), .A2(n7235), .ZN(n7053) );
  OR2_X1 U8681 ( .A1(n7248), .A2(n7051), .ZN(n7052) );
  NAND2_X1 U8682 ( .A1(n7510), .A2(n7235), .ZN(n7055) );
  AOI22_X1 U8683 ( .A1(n7080), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n7079), .B2(
        n8034), .ZN(n7054) );
  OR2_X1 U8684 ( .A1(n9332), .A2(n8248), .ZN(n7338) );
  NAND2_X1 U8685 ( .A1(n9332), .A2(n8248), .ZN(n8244) );
  NAND2_X1 U8686 ( .A1(n7338), .A2(n8244), .ZN(n9325) );
  NAND2_X1 U8687 ( .A1(n7523), .A2(n7235), .ZN(n7059) );
  AOI22_X1 U8688 ( .A1(n7080), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n7079), .B2(
        n8050), .ZN(n7058) );
  NAND2_X1 U8689 ( .A1(n7127), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7068) );
  INV_X1 U8690 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n7060) );
  OR2_X1 U8691 ( .A1(n7224), .A2(n7060), .ZN(n7067) );
  INV_X1 U8692 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n7061) );
  NAND2_X1 U8693 ( .A1(n7062), .A2(n7061), .ZN(n7063) );
  NAND2_X1 U8694 ( .A1(n7071), .A2(n7063), .ZN(n8239) );
  OR2_X1 U8695 ( .A1(n7168), .A2(n8239), .ZN(n7066) );
  INV_X1 U8696 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n7064) );
  OR2_X1 U8697 ( .A1(n5579), .A2(n7064), .ZN(n7065) );
  NAND4_X1 U8698 ( .A1(n7068), .A2(n7067), .A3(n7066), .A4(n7065), .ZN(n8228)
         );
  INV_X1 U8699 ( .A(n8228), .ZN(n7954) );
  NAND2_X1 U8700 ( .A1(n8349), .A2(n7954), .ZN(n7259) );
  NAND2_X1 U8701 ( .A1(n7546), .A2(n7235), .ZN(n7070) );
  AOI22_X1 U8702 ( .A1(n7080), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n7079), .B2(
        n8048), .ZN(n7069) );
  NAND2_X1 U8703 ( .A1(n7127), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n7077) );
  INV_X1 U8704 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8062) );
  OR2_X1 U8705 ( .A1(n7224), .A2(n8062), .ZN(n7076) );
  NAND2_X1 U8706 ( .A1(n7071), .A2(n9830), .ZN(n7072) );
  NAND2_X1 U8707 ( .A1(n7095), .A2(n7072), .ZN(n8223) );
  OR2_X1 U8708 ( .A1(n7168), .A2(n8223), .ZN(n7075) );
  INV_X1 U8709 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n7073) );
  OR2_X1 U8710 ( .A1(n5579), .A2(n7073), .ZN(n7074) );
  NAND4_X1 U8711 ( .A1(n7077), .A2(n7076), .A3(n7075), .A4(n7074), .ZN(n8208)
         );
  NOR2_X1 U8712 ( .A1(n8342), .A2(n8208), .ZN(n7078) );
  INV_X1 U8713 ( .A(n8342), .ZN(n8222) );
  INV_X1 U8714 ( .A(n8208), .ZN(n8250) );
  NAND2_X1 U8715 ( .A1(n7565), .A2(n7235), .ZN(n7082) );
  AOI22_X1 U8716 ( .A1(n7080), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5547), .B2(
        n7079), .ZN(n7081) );
  NAND2_X2 U8717 ( .A1(n7082), .A2(n7081), .ZN(n8338) );
  XNOR2_X1 U8718 ( .A(n7095), .B(P2_REG3_REG_19__SCAN_IN), .ZN(n8212) );
  NAND2_X1 U8719 ( .A1(n5712), .A2(n8212), .ZN(n7088) );
  INV_X1 U8720 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n7083) );
  OR2_X1 U8721 ( .A1(n7224), .A2(n7083), .ZN(n7087) );
  INV_X1 U8722 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n7084) );
  OR2_X1 U8723 ( .A1(n5579), .A2(n7084), .ZN(n7086) );
  INV_X1 U8724 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8061) );
  OR2_X1 U8725 ( .A1(n7228), .A2(n8061), .ZN(n7085) );
  NAND4_X1 U8726 ( .A1(n7088), .A2(n7087), .A3(n7086), .A4(n7085), .ZN(n8229)
         );
  NAND2_X1 U8727 ( .A1(n8204), .A2(n7089), .ZN(n7090) );
  INV_X1 U8728 ( .A(n8338), .ZN(n8205) );
  INV_X1 U8729 ( .A(n8229), .ZN(n7953) );
  NOR2_X1 U8730 ( .A1(n7248), .A2(n7091), .ZN(n7092) );
  NAND2_X1 U8731 ( .A1(n5576), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n7101) );
  INV_X1 U8732 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n7093) );
  OR2_X1 U8733 ( .A1(n7228), .A2(n7093), .ZN(n7100) );
  INV_X1 U8734 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n7094) );
  INV_X1 U8735 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n7935) );
  OAI21_X1 U8736 ( .B1(n7095), .B2(n7094), .A(n7935), .ZN(n7096) );
  NAND2_X1 U8737 ( .A1(n7105), .A2(n7096), .ZN(n8191) );
  OR2_X1 U8738 ( .A1(n8191), .A2(n7168), .ZN(n7099) );
  INV_X1 U8739 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n7097) );
  OR2_X1 U8740 ( .A1(n5579), .A2(n7097), .ZN(n7098) );
  NAND4_X1 U8741 ( .A1(n7101), .A2(n7100), .A3(n7099), .A4(n7098), .ZN(n8209)
         );
  NAND2_X1 U8742 ( .A1(n8194), .A2(n8209), .ZN(n7356) );
  OR2_X1 U8743 ( .A1(n8194), .A2(n8209), .ZN(n7352) );
  INV_X1 U8744 ( .A(n8194), .ZN(n8332) );
  NAND2_X1 U8745 ( .A1(n7604), .A2(n7235), .ZN(n7104) );
  OR2_X1 U8746 ( .A1(n7248), .A2(n7102), .ZN(n7103) );
  INV_X1 U8747 ( .A(n8327), .ZN(n8177) );
  NAND2_X1 U8748 ( .A1(n7105), .A2(n7891), .ZN(n7106) );
  NAND2_X1 U8749 ( .A1(n7124), .A2(n7106), .ZN(n8174) );
  NAND2_X1 U8750 ( .A1(n5576), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n7108) );
  NAND2_X1 U8751 ( .A1(n7222), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n7107) );
  AND2_X1 U8752 ( .A1(n7108), .A2(n7107), .ZN(n7111) );
  INV_X1 U8753 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n7109) );
  OR2_X1 U8754 ( .A1(n7228), .A2(n7109), .ZN(n7110) );
  OAI211_X1 U8755 ( .C1(n8174), .C2(n7168), .A(n7111), .B(n7110), .ZN(n8199)
         );
  INV_X1 U8756 ( .A(n8199), .ZN(n8165) );
  NAND2_X1 U8757 ( .A1(n7626), .A2(n7235), .ZN(n7115) );
  OR2_X1 U8758 ( .A1(n7248), .A2(n7113), .ZN(n7114) );
  XNOR2_X1 U8759 ( .A(n7124), .B(P2_REG3_REG_22__SCAN_IN), .ZN(n8158) );
  NAND2_X1 U8760 ( .A1(n8158), .A2(n5712), .ZN(n7120) );
  INV_X1 U8761 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9858) );
  NAND2_X1 U8762 ( .A1(n5576), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n7117) );
  NAND2_X1 U8763 ( .A1(n7127), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n7116) );
  OAI211_X1 U8764 ( .C1(n5579), .C2(n9858), .A(n7117), .B(n7116), .ZN(n7118)
         );
  INV_X1 U8765 ( .A(n7118), .ZN(n7119) );
  NAND2_X1 U8766 ( .A1(n7120), .A2(n7119), .ZN(n8183) );
  INV_X1 U8767 ( .A(n8183), .ZN(n7892) );
  NAND2_X1 U8768 ( .A1(n8322), .A2(n7892), .ZN(n7360) );
  INV_X1 U8769 ( .A(n8322), .ZN(n8160) );
  AOI22_X1 U8770 ( .A1(n8155), .A2(n8163), .B1(n8160), .B2(n7892), .ZN(n8147)
         );
  NAND2_X1 U8771 ( .A1(n7476), .A2(n7235), .ZN(n7123) );
  OR2_X1 U8772 ( .A1(n7248), .A2(n7121), .ZN(n7122) );
  INV_X1 U8773 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n7944) );
  INV_X1 U8774 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n7857) );
  OAI21_X1 U8775 ( .B1(n7124), .B2(n7944), .A(n7857), .ZN(n7126) );
  NAND2_X1 U8776 ( .A1(n7126), .A2(n7125), .ZN(n8149) );
  OR2_X1 U8777 ( .A1(n8149), .A2(n7168), .ZN(n7130) );
  AOI22_X1 U8778 ( .A1(n7127), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n5576), .B2(
        P2_REG1_REG_23__SCAN_IN), .ZN(n7129) );
  NAND2_X1 U8779 ( .A1(n7222), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n7128) );
  NAND2_X1 U8780 ( .A1(n8147), .A2(n8146), .ZN(n8315) );
  NAND2_X1 U8781 ( .A1(n8315), .A2(n4818), .ZN(n8125) );
  OR2_X1 U8782 ( .A1(n7248), .A2(n7131), .ZN(n7132) );
  INV_X1 U8783 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n7900) );
  NAND2_X1 U8784 ( .A1(n7134), .A2(n7900), .ZN(n7135) );
  AND2_X1 U8785 ( .A1(n7146), .A2(n7135), .ZN(n8114) );
  NAND2_X1 U8786 ( .A1(n8114), .A2(n5712), .ZN(n7141) );
  INV_X1 U8787 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n7138) );
  NAND2_X1 U8788 ( .A1(n5576), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n7137) );
  NAND2_X1 U8789 ( .A1(n7222), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n7136) );
  OAI211_X1 U8790 ( .C1(n7228), .C2(n7138), .A(n7137), .B(n7136), .ZN(n7139)
         );
  INV_X1 U8791 ( .A(n7139), .ZN(n7140) );
  NAND2_X1 U8792 ( .A1(n7141), .A2(n7140), .ZN(n8132) );
  NAND2_X1 U8793 ( .A1(n7679), .A2(n7235), .ZN(n7144) );
  OR2_X1 U8794 ( .A1(n7248), .A2(n7142), .ZN(n7143) );
  INV_X1 U8795 ( .A(n7146), .ZN(n7145) );
  NAND2_X1 U8796 ( .A1(n7145), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n7166) );
  INV_X1 U8797 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n7961) );
  NAND2_X1 U8798 ( .A1(n7146), .A2(n7961), .ZN(n7147) );
  NAND2_X1 U8799 ( .A1(n7166), .A2(n7147), .ZN(n8101) );
  OR2_X1 U8800 ( .A1(n8101), .A2(n7168), .ZN(n7153) );
  INV_X1 U8801 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n7150) );
  NAND2_X1 U8802 ( .A1(n5576), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n7149) );
  NAND2_X1 U8803 ( .A1(n7222), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n7148) );
  OAI211_X1 U8804 ( .C1(n7150), .C2(n7228), .A(n7149), .B(n7148), .ZN(n7151)
         );
  INV_X1 U8805 ( .A(n7151), .ZN(n7152) );
  NAND2_X1 U8806 ( .A1(n7153), .A2(n7152), .ZN(n8119) );
  NAND2_X1 U8807 ( .A1(n8301), .A2(n7901), .ZN(n7372) );
  OR2_X1 U8808 ( .A1(n7248), .A2(n7154), .ZN(n7155) );
  XNOR2_X1 U8809 ( .A(n7166), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8087) );
  NAND2_X1 U8810 ( .A1(n8087), .A2(n5712), .ZN(n7162) );
  INV_X1 U8811 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n7159) );
  NAND2_X1 U8812 ( .A1(n7222), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n7158) );
  NAND2_X1 U8813 ( .A1(n5576), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n7157) );
  OAI211_X1 U8814 ( .C1(n7159), .C2(n7228), .A(n7158), .B(n7157), .ZN(n7160)
         );
  INV_X1 U8815 ( .A(n7160), .ZN(n7161) );
  NAND2_X1 U8816 ( .A1(n7162), .A2(n7161), .ZN(n8107) );
  INV_X1 U8817 ( .A(n8107), .ZN(n7962) );
  NAND2_X1 U8818 ( .A1(n8296), .A2(n7962), .ZN(n7379) );
  NAND2_X1 U8819 ( .A1(n7757), .A2(n7235), .ZN(n7165) );
  OR2_X1 U8820 ( .A1(n7248), .A2(n7163), .ZN(n7164) );
  INV_X1 U8821 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n7848) );
  INV_X1 U8822 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n7882) );
  OAI21_X1 U8823 ( .B1(n7166), .B2(n7848), .A(n7882), .ZN(n7167) );
  NAND2_X1 U8824 ( .A1(n7167), .A2(n7193), .ZN(n7883) );
  OR2_X1 U8825 ( .A1(n7883), .A2(n7168), .ZN(n7174) );
  INV_X1 U8826 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n7171) );
  NAND2_X1 U8827 ( .A1(n7222), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n7170) );
  NAND2_X1 U8828 ( .A1(n5576), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n7169) );
  OAI211_X1 U8829 ( .C1(n7171), .C2(n7228), .A(n7170), .B(n7169), .ZN(n7172)
         );
  INV_X1 U8830 ( .A(n7172), .ZN(n7173) );
  NAND2_X1 U8831 ( .A1(n7174), .A2(n7173), .ZN(n8092) );
  INV_X1 U8832 ( .A(n8092), .ZN(n7849) );
  NAND2_X1 U8833 ( .A1(n8290), .A2(n7849), .ZN(n7381) );
  XNOR2_X1 U8834 ( .A(n7442), .B(n7422), .ZN(n8294) );
  NAND2_X1 U8835 ( .A1(n8104), .A2(n8113), .ZN(n8098) );
  INV_X1 U8836 ( .A(n8086), .ZN(n7177) );
  INV_X1 U8837 ( .A(n8290), .ZN(n7440) );
  NAND2_X1 U8838 ( .A1(n7440), .A2(n8086), .ZN(n7444) );
  INV_X1 U8839 ( .A(n7444), .ZN(n7176) );
  AOI21_X1 U8840 ( .B1(n8290), .B2(n7177), .A(n7176), .ZN(n8291) );
  INV_X1 U8841 ( .A(n8265), .ZN(n9590) );
  INV_X1 U8842 ( .A(n7883), .ZN(n7178) );
  AOI22_X1 U8843 ( .A1(P2_REG2_REG_28__SCAN_IN), .A2(n9590), .B1(n7178), .B2(
        n9613), .ZN(n7179) );
  OAI21_X1 U8844 ( .B1(n7440), .B2(n8237), .A(n7179), .ZN(n7200) );
  NAND2_X1 U8845 ( .A1(n9323), .A2(n4785), .ZN(n9322) );
  INV_X1 U8846 ( .A(n8244), .ZN(n7182) );
  NOR2_X1 U8847 ( .A1(n8245), .A2(n7182), .ZN(n7183) );
  OR2_X1 U8848 ( .A1(n8342), .A2(n8250), .ZN(n7343) );
  NAND2_X1 U8849 ( .A1(n8342), .A2(n8250), .ZN(n7263) );
  OR2_X1 U8850 ( .A1(n8338), .A2(n7953), .ZN(n7350) );
  NAND2_X1 U8851 ( .A1(n8338), .A2(n7953), .ZN(n8196) );
  NAND2_X1 U8852 ( .A1(n8206), .A2(n8207), .ZN(n8195) );
  INV_X1 U8853 ( .A(n8196), .ZN(n7184) );
  NOR2_X1 U8854 ( .A1(n8198), .A2(n7184), .ZN(n7185) );
  NAND2_X1 U8855 ( .A1(n8195), .A2(n7185), .ZN(n7186) );
  NAND2_X1 U8856 ( .A1(n7186), .A2(n7356), .ZN(n8178) );
  OR2_X1 U8857 ( .A1(n8327), .A2(n8165), .ZN(n7357) );
  NAND2_X1 U8858 ( .A1(n8327), .A2(n8165), .ZN(n8162) );
  NAND2_X1 U8859 ( .A1(n7357), .A2(n8162), .ZN(n8179) );
  OR2_X2 U8860 ( .A1(n8178), .A2(n8179), .ZN(n8161) );
  INV_X1 U8861 ( .A(n8162), .ZN(n7187) );
  NOR2_X1 U8862 ( .A1(n8163), .A2(n7187), .ZN(n7188) );
  NAND2_X1 U8863 ( .A1(n8317), .A2(n8166), .ZN(n7189) );
  NAND2_X1 U8864 ( .A1(n8117), .A2(n8118), .ZN(n7191) );
  INV_X1 U8865 ( .A(n8132), .ZN(n7963) );
  OR2_X1 U8866 ( .A1(n8306), .A2(n7963), .ZN(n7190) );
  XNOR2_X1 U8867 ( .A(n7230), .B(n7441), .ZN(n7198) );
  INV_X1 U8868 ( .A(n7193), .ZN(n7445) );
  INV_X1 U8869 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n7196) );
  NAND2_X1 U8870 ( .A1(n7222), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n7195) );
  NAND2_X1 U8871 ( .A1(n5576), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n7194) );
  OAI211_X1 U8872 ( .C1(n7196), .C2(n7228), .A(n7195), .B(n7194), .ZN(n7197)
         );
  AOI21_X1 U8873 ( .B1(n7445), .B2(n5712), .A(n7197), .ZN(n7884) );
  INV_X1 U8874 ( .A(n7884), .ZN(n7981) );
  AOI222_X1 U8875 ( .A1(n9619), .A2(n7198), .B1(n8107), .B2(n9624), .C1(n7981), 
        .C2(n9621), .ZN(n8293) );
  NOR2_X1 U8876 ( .A1(n8293), .A2(n8217), .ZN(n7199) );
  AOI211_X1 U8877 ( .C1(n9337), .C2(n8291), .A(n7200), .B(n7199), .ZN(n7201)
         );
  OAI21_X1 U8878 ( .B1(n8294), .B2(n8254), .A(n7201), .ZN(P2_U3268) );
  AOI22_X1 U8879 ( .A1(n7202), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n9265), .ZN(n7203) );
  OAI21_X1 U8880 ( .B1(n7204), .B2(n9273), .A(n7203), .ZN(P1_U3349) );
  NAND2_X1 U8881 ( .A1(n6014), .A2(n7207), .ZN(n7209) );
  AND2_X1 U8882 ( .A1(n7209), .A2(n7208), .ZN(n7210) );
  AOI211_X1 U8883 ( .C1(n7205), .C2(n7210), .A(n8519), .B(n4286), .ZN(n7218)
         );
  OAI22_X1 U8884 ( .A1(n8512), .A2(n9488), .B1(n7211), .B2(n8487), .ZN(n7217)
         );
  NAND2_X1 U8885 ( .A1(n8517), .A2(n7212), .ZN(n7213) );
  OAI211_X1 U8886 ( .C1(n8500), .C2(n7215), .A(n7214), .B(n7213), .ZN(n7216)
         );
  OR3_X1 U8887 ( .A1(n7218), .A2(n7217), .A3(n7216), .ZN(P1_U3228) );
  NAND2_X1 U8888 ( .A1(n8611), .A2(n7235), .ZN(n7221) );
  OR2_X1 U8889 ( .A1(n7248), .A2(n7219), .ZN(n7220) );
  INV_X1 U8890 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n7227) );
  NAND2_X1 U8891 ( .A1(n7222), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n7226) );
  INV_X1 U8892 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n7223) );
  OR2_X1 U8893 ( .A1(n7224), .A2(n7223), .ZN(n7225) );
  OAI211_X1 U8894 ( .C1(n7228), .C2(n7227), .A(n7226), .B(n7225), .ZN(n7980)
         );
  INV_X1 U8895 ( .A(n7980), .ZN(n7252) );
  INV_X1 U8896 ( .A(n7383), .ZN(n7229) );
  XNOR2_X1 U8897 ( .A(n7233), .B(n7232), .ZN(n7234) );
  NAND2_X1 U8898 ( .A1(n8521), .A2(n7235), .ZN(n7237) );
  INV_X1 U8899 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7755) );
  OR2_X1 U8900 ( .A1(n7248), .A2(n7755), .ZN(n7236) );
  NAND2_X1 U8901 ( .A1(n8287), .A2(n7884), .ZN(n7386) );
  INV_X1 U8902 ( .A(n7238), .ZN(n7239) );
  NAND2_X1 U8903 ( .A1(n7239), .A2(SI_30_), .ZN(n7243) );
  NAND2_X1 U8904 ( .A1(n7241), .A2(n7240), .ZN(n7242) );
  NAND2_X1 U8905 ( .A1(n7243), .A2(n7242), .ZN(n7247) );
  MUX2_X1 U8906 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7244), .Z(n7245) );
  XNOR2_X1 U8907 ( .A(n7245), .B(SI_31_), .ZN(n7246) );
  NAND2_X1 U8908 ( .A1(n8608), .A2(n7235), .ZN(n7250) );
  OR2_X1 U8909 ( .A1(n7248), .A2(n5501), .ZN(n7249) );
  INV_X1 U8910 ( .A(n8074), .ZN(n7251) );
  NAND2_X1 U8911 ( .A1(n8081), .A2(n7252), .ZN(n7388) );
  NAND2_X1 U8912 ( .A1(n7390), .A2(n7388), .ZN(n7424) );
  NOR2_X1 U8913 ( .A1(n8075), .A2(n8074), .ZN(n7393) );
  NOR2_X1 U8914 ( .A1(n7254), .A2(n7393), .ZN(n7255) );
  XNOR2_X1 U8915 ( .A(n7255), .B(n8213), .ZN(n7434) );
  NAND2_X1 U8916 ( .A1(n4269), .A2(n7256), .ZN(n7433) );
  INV_X1 U8917 ( .A(n7389), .ZN(n7257) );
  NOR2_X1 U8918 ( .A1(n7393), .A2(n7257), .ZN(n7398) );
  MUX2_X1 U8919 ( .A(n4550), .B(n7398), .S(n7391), .Z(n7395) );
  NAND2_X1 U8920 ( .A1(n8306), .A2(n7963), .ZN(n7258) );
  AOI21_X1 U8921 ( .B1(n7372), .B2(n7258), .A(n7384), .ZN(n7376) );
  INV_X1 U8922 ( .A(n7259), .ZN(n7262) );
  NAND2_X1 U8923 ( .A1(n7343), .A2(n7260), .ZN(n7261) );
  MUX2_X1 U8924 ( .A(n7262), .B(n7261), .S(n7391), .Z(n7264) );
  NOR2_X1 U8925 ( .A1(n7264), .A2(n4571), .ZN(n7342) );
  NAND2_X1 U8926 ( .A1(n7317), .A2(n7265), .ZN(n7302) );
  NAND2_X1 U8927 ( .A1(n7299), .A2(n7304), .ZN(n7267) );
  NAND2_X1 U8928 ( .A1(n7399), .A2(n7313), .ZN(n7266) );
  MUX2_X1 U8929 ( .A(n7267), .B(n7266), .S(n7391), .Z(n7312) );
  NAND2_X1 U8930 ( .A1(n7268), .A2(n7391), .ZN(n7270) );
  AND2_X1 U8931 ( .A1(n7277), .A2(n7429), .ZN(n7274) );
  OAI211_X1 U8932 ( .C1(n8260), .C2(n7274), .A(n7273), .B(n8256), .ZN(n7276)
         );
  NAND3_X1 U8933 ( .A1(n7276), .A2(n7279), .A3(n7275), .ZN(n7282) );
  NAND2_X1 U8934 ( .A1(n8256), .A2(n7277), .ZN(n7401) );
  NAND3_X1 U8935 ( .A1(n7401), .A2(n7279), .A3(n7278), .ZN(n7280) );
  NAND2_X1 U8936 ( .A1(n7283), .A2(n7288), .ZN(n7292) );
  NAND2_X1 U8937 ( .A1(n9615), .A2(n7284), .ZN(n7285) );
  NAND2_X1 U8938 ( .A1(n7286), .A2(n7285), .ZN(n7289) );
  NAND3_X1 U8939 ( .A1(n7289), .A2(n7288), .A3(n7287), .ZN(n7290) );
  NAND2_X1 U8940 ( .A1(n7290), .A2(n7384), .ZN(n7291) );
  NAND2_X1 U8941 ( .A1(n7292), .A2(n7291), .ZN(n7297) );
  NOR2_X1 U8942 ( .A1(n7293), .A2(n7391), .ZN(n7294) );
  NOR2_X1 U8943 ( .A1(n7295), .A2(n7294), .ZN(n7296) );
  NAND2_X1 U8944 ( .A1(n7297), .A2(n7296), .ZN(n7309) );
  NAND3_X1 U8945 ( .A1(n7309), .A2(n7407), .A3(n7298), .ZN(n7300) );
  OAI211_X1 U8946 ( .C1(n7312), .C2(n7300), .A(n9583), .B(n7299), .ZN(n7301)
         );
  MUX2_X1 U8947 ( .A(n7302), .B(n7301), .S(n7391), .Z(n7316) );
  AND2_X1 U8948 ( .A1(n7304), .A2(n7303), .ZN(n7311) );
  AND2_X1 U8949 ( .A1(n7407), .A2(n7305), .ZN(n7308) );
  INV_X1 U8950 ( .A(n7306), .ZN(n7307) );
  AOI21_X1 U8951 ( .B1(n7309), .B2(n7308), .A(n7307), .ZN(n7310) );
  MUX2_X1 U8952 ( .A(n7311), .B(n7310), .S(n7384), .Z(n7314) );
  AOI21_X1 U8953 ( .B1(n7314), .B2(n7313), .A(n7312), .ZN(n7315) );
  OR2_X1 U8954 ( .A1(n7316), .A2(n7315), .ZN(n7324) );
  AND2_X1 U8955 ( .A1(n7321), .A2(n7317), .ZN(n7320) );
  INV_X1 U8956 ( .A(n7318), .ZN(n7319) );
  AOI21_X1 U8957 ( .B1(n7324), .B2(n7320), .A(n7319), .ZN(n7326) );
  INV_X1 U8958 ( .A(n7321), .ZN(n7322) );
  AOI21_X1 U8959 ( .B1(n7324), .B2(n7323), .A(n7322), .ZN(n7325) );
  INV_X1 U8960 ( .A(n9354), .ZN(n9342) );
  MUX2_X1 U8961 ( .A(n9343), .B(n7327), .S(n7384), .Z(n7328) );
  MUX2_X1 U8962 ( .A(n7330), .B(n7329), .S(n7391), .Z(n7331) );
  MUX2_X1 U8963 ( .A(n7334), .B(n7333), .S(n7391), .Z(n7335) );
  NAND2_X1 U8964 ( .A1(n7336), .A2(n7335), .ZN(n7337) );
  NAND2_X1 U8965 ( .A1(n7337), .A2(n4785), .ZN(n7340) );
  MUX2_X1 U8966 ( .A(n7338), .B(n8244), .S(n7391), .Z(n7339) );
  NAND3_X1 U8967 ( .A1(n7340), .A2(n7418), .A3(n7339), .ZN(n7341) );
  NAND2_X1 U8968 ( .A1(n7342), .A2(n7341), .ZN(n7355) );
  NAND3_X1 U8969 ( .A1(n7355), .A2(n7350), .A3(n7343), .ZN(n7344) );
  NAND2_X1 U8970 ( .A1(n7344), .A2(n8196), .ZN(n7345) );
  NAND2_X1 U8971 ( .A1(n7345), .A2(n7356), .ZN(n7346) );
  NAND3_X1 U8972 ( .A1(n7346), .A2(n8162), .A3(n7352), .ZN(n7347) );
  NAND3_X1 U8973 ( .A1(n7347), .A2(n7384), .A3(n7357), .ZN(n7349) );
  MUX2_X1 U8974 ( .A(n7384), .B(n7349), .S(n7348), .Z(n7363) );
  INV_X1 U8975 ( .A(n8146), .ZN(n8143) );
  INV_X1 U8976 ( .A(n7350), .ZN(n7354) );
  NAND2_X1 U8977 ( .A1(n7350), .A2(n4571), .ZN(n7351) );
  AND2_X1 U8978 ( .A1(n7351), .A2(n8196), .ZN(n7353) );
  OAI211_X1 U8979 ( .C1(n7355), .C2(n7354), .A(n7353), .B(n7352), .ZN(n7358)
         );
  NAND3_X1 U8980 ( .A1(n7358), .A2(n7357), .A3(n7356), .ZN(n7359) );
  NAND3_X1 U8981 ( .A1(n7359), .A2(n7360), .A3(n8162), .ZN(n7361) );
  MUX2_X1 U8982 ( .A(n7361), .B(n7360), .S(n7384), .Z(n7362) );
  NAND3_X1 U8983 ( .A1(n7363), .A2(n8143), .A3(n7362), .ZN(n7367) );
  OR2_X1 U8984 ( .A1(n8166), .A2(n7391), .ZN(n7365) );
  NAND2_X1 U8985 ( .A1(n8166), .A2(n7391), .ZN(n7364) );
  MUX2_X1 U8986 ( .A(n7365), .B(n7364), .S(n8317), .Z(n7366) );
  NAND2_X1 U8987 ( .A1(n8310), .A2(n7903), .ZN(n7369) );
  MUX2_X1 U8988 ( .A(n7369), .B(n7368), .S(n7391), .Z(n7370) );
  OR3_X1 U8989 ( .A1(n8306), .A2(n7963), .A3(n7391), .ZN(n7371) );
  OR2_X1 U8990 ( .A1(n7373), .A2(n7384), .ZN(n7374) );
  OAI211_X1 U8991 ( .C1(n7376), .C2(n7375), .A(n8091), .B(n7374), .ZN(n7377)
         );
  OAI211_X1 U8992 ( .C1(n7378), .C2(n7391), .A(n7377), .B(n7383), .ZN(n7382)
         );
  AOI21_X1 U8993 ( .B1(n7381), .B2(n7379), .A(n7384), .ZN(n7380) );
  MUX2_X1 U8994 ( .A(n7386), .B(n7385), .S(n7384), .Z(n7387) );
  INV_X1 U8995 ( .A(n7390), .ZN(n7392) );
  MUX2_X1 U8996 ( .A(n7393), .B(n7392), .S(n7391), .Z(n7394) );
  NOR2_X1 U8997 ( .A1(n7396), .A2(n7428), .ZN(n7431) );
  INV_X1 U8998 ( .A(n7398), .ZN(n7425) );
  INV_X1 U8999 ( .A(n7399), .ZN(n7411) );
  OR4_X1 U9000 ( .A1(n7401), .A2(n7400), .A3(n8260), .A4(n8286), .ZN(n7404) );
  NOR4_X1 U9001 ( .A1(n7404), .A2(n9617), .A3(n7403), .A4(n7402), .ZN(n7408)
         );
  NAND4_X1 U9002 ( .A1(n7408), .A2(n7407), .A3(n7406), .A4(n7405), .ZN(n7410)
         );
  NOR4_X1 U9003 ( .A1(n7412), .A2(n7411), .A3(n7410), .A4(n7409), .ZN(n7413)
         );
  NAND3_X1 U9004 ( .A1(n7414), .A2(n7413), .A3(n9593), .ZN(n7415) );
  NOR4_X1 U9005 ( .A1(n9325), .A2(n7416), .A3(n9354), .A4(n7415), .ZN(n7417)
         );
  NAND4_X1 U9006 ( .A1(n8207), .A2(n4282), .A3(n7418), .A4(n7417), .ZN(n7419)
         );
  OR4_X1 U9007 ( .A1(n8163), .A2(n8179), .A3(n8198), .A4(n7419), .ZN(n7420) );
  NOR4_X1 U9008 ( .A1(n8106), .A2(n8146), .A3(n8127), .A4(n7420), .ZN(n7421)
         );
  NAND4_X1 U9009 ( .A1(n7422), .A2(n8091), .A3(n7421), .A4(n8118), .ZN(n7423)
         );
  XNOR2_X1 U9010 ( .A(n7426), .B(n5547), .ZN(n7430) );
  OAI22_X1 U9011 ( .A1(n7430), .A2(n7429), .B1(n7428), .B2(n7427), .ZN(n7432)
         );
  NOR4_X1 U9012 ( .A1(n9631), .A2(n8249), .A3(n7435), .A4(n5186), .ZN(n7437)
         );
  OAI21_X1 U9013 ( .B1(n7438), .B2(n5548), .A(P2_B_REG_SCAN_IN), .ZN(n7436) );
  OAI22_X1 U9014 ( .A1(n7439), .A2(n7438), .B1(n7437), .B2(n7436), .ZN(
        P2_U3244) );
  AOI22_X1 U9015 ( .A1(n7442), .A2(n7441), .B1(n7440), .B2(n7849), .ZN(n7443)
         );
  XNOR2_X1 U9016 ( .A(n7443), .B(n7448), .ZN(n8289) );
  AOI21_X1 U9017 ( .B1(n8287), .B2(n7444), .A(n8079), .ZN(n8288) );
  INV_X1 U9018 ( .A(n8287), .ZN(n7447) );
  AOI22_X1 U9019 ( .A1(n8217), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n7445), .B2(
        n9613), .ZN(n7446) );
  OAI21_X1 U9020 ( .B1(n7447), .B2(n8237), .A(n7446), .ZN(n7458) );
  INV_X1 U9021 ( .A(P2_B_REG_SCAN_IN), .ZN(n9892) );
  NOR2_X1 U9022 ( .A1(n5186), .A2(n9892), .ZN(n7452) );
  NOR2_X1 U9023 ( .A1(n8251), .A2(n7452), .ZN(n8073) );
  INV_X1 U9024 ( .A(n8073), .ZN(n7453) );
  AOI21_X1 U9025 ( .B1(n8092), .B2(n9624), .A(n7454), .ZN(n7455) );
  NOR2_X1 U9026 ( .A1(n4813), .A2(n8217), .ZN(n7457) );
  AOI211_X1 U9027 ( .C1(n8288), .C2(n9337), .A(n7458), .B(n7457), .ZN(n7459)
         );
  OAI21_X1 U9028 ( .B1(n8289), .B2(n8254), .A(n7459), .ZN(P2_U3267) );
  NAND2_X1 U9029 ( .A1(n7460), .A2(n7642), .ZN(n7462) );
  NAND2_X1 U9030 ( .A1(n8612), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n7461) );
  NAND2_X1 U9031 ( .A1(n9136), .A2(n4263), .ZN(n7471) );
  INV_X1 U9032 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n7527) );
  INV_X1 U9033 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8409) );
  INV_X1 U9034 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9856) );
  INV_X1 U9035 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n7479) );
  INV_X1 U9036 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n7664) );
  INV_X1 U9037 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n7682) );
  XNOR2_X1 U9038 ( .A(n7710), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n8947) );
  INV_X1 U9039 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9843) );
  NAND2_X1 U9040 ( .A1(n7591), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n7468) );
  NAND2_X1 U9041 ( .A1(n5785), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n7467) );
  OAI211_X1 U9042 ( .C1(n7772), .C2(n9843), .A(n7468), .B(n7467), .ZN(n7469)
         );
  OR2_X1 U9043 ( .A1(n8899), .A2(n6011), .ZN(n7470) );
  NAND2_X1 U9044 ( .A1(n7471), .A2(n7470), .ZN(n7472) );
  XNOR2_X1 U9045 ( .A(n7472), .B(n7762), .ZN(n7475) );
  INV_X1 U9046 ( .A(n6703), .ZN(n7677) );
  NOR2_X1 U9047 ( .A1(n8899), .A2(n7677), .ZN(n7473) );
  AOI21_X1 U9048 ( .B1(n9136), .B2(n7485), .A(n7473), .ZN(n7474) );
  NAND2_X1 U9049 ( .A1(n7475), .A2(n7474), .ZN(n7781) );
  OAI21_X1 U9050 ( .B1(n7475), .B2(n7474), .A(n7781), .ZN(n7704) );
  NAND2_X1 U9051 ( .A1(n7476), .A2(n7642), .ZN(n7478) );
  NAND2_X1 U9052 ( .A1(n8612), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7477) );
  NAND2_X1 U9053 ( .A1(n7631), .A2(n7479), .ZN(n7480) );
  AND2_X1 U9054 ( .A1(n7646), .A2(n7480), .ZN(n8992) );
  NAND2_X1 U9055 ( .A1(n8992), .A2(n7571), .ZN(n7483) );
  AOI22_X1 U9056 ( .A1(n8615), .A2(P1_REG1_REG_23__SCAN_IN), .B1(n5785), .B2(
        P1_REG0_REG_23__SCAN_IN), .ZN(n7482) );
  NAND2_X1 U9057 ( .A1(n7591), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n7481) );
  INV_X1 U9058 ( .A(n8474), .ZN(n9013) );
  AOI22_X1 U9059 ( .A1(n9157), .A2(n7485), .B1(n7484), .B2(n9013), .ZN(n8397)
         );
  AND2_X1 U9060 ( .A1(n7487), .A2(n7486), .ZN(n7489) );
  NAND2_X1 U9061 ( .A1(n9205), .A2(n4263), .ZN(n7492) );
  NAND2_X1 U9062 ( .A1(n8810), .A2(n7485), .ZN(n7491) );
  NAND2_X1 U9063 ( .A1(n7492), .A2(n7491), .ZN(n7493) );
  XNOR2_X1 U9064 ( .A(n7493), .B(n7675), .ZN(n8387) );
  INV_X1 U9065 ( .A(n8387), .ZN(n7496) );
  NAND2_X1 U9066 ( .A1(n9205), .A2(n7485), .ZN(n7495) );
  NAND2_X1 U9067 ( .A1(n8810), .A2(n7484), .ZN(n7494) );
  NAND2_X1 U9068 ( .A1(n7495), .A2(n7494), .ZN(n7501) );
  INV_X1 U9069 ( .A(n7501), .ZN(n8386) );
  NAND2_X1 U9070 ( .A1(n7496), .A2(n8386), .ZN(n7506) );
  NAND2_X1 U9071 ( .A1(n9199), .A2(n4263), .ZN(n7499) );
  NAND2_X1 U9072 ( .A1(n9113), .A2(n7485), .ZN(n7498) );
  NAND2_X1 U9073 ( .A1(n7499), .A2(n7498), .ZN(n7500) );
  XNOR2_X1 U9074 ( .A(n7500), .B(n7675), .ZN(n7507) );
  INV_X1 U9075 ( .A(n7507), .ZN(n7503) );
  AND2_X1 U9076 ( .A1(n8387), .A2(n7501), .ZN(n7509) );
  INV_X1 U9077 ( .A(n7509), .ZN(n7502) );
  NAND2_X1 U9078 ( .A1(n9199), .A2(n7485), .ZN(n7505) );
  NAND2_X1 U9079 ( .A1(n9113), .A2(n7484), .ZN(n7504) );
  NAND2_X1 U9080 ( .A1(n7505), .A2(n7504), .ZN(n8508) );
  AND2_X1 U9081 ( .A1(n7507), .A2(n7506), .ZN(n7508) );
  NAND2_X1 U9082 ( .A1(n7510), .A2(n7642), .ZN(n7512) );
  AOI22_X1 U9083 ( .A1(n7566), .A2(n8844), .B1(n7524), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n7511) );
  NAND2_X1 U9084 ( .A1(n9195), .A2(n4263), .ZN(n7514) );
  NAND2_X1 U9085 ( .A1(n9095), .A2(n7485), .ZN(n7513) );
  NAND2_X1 U9086 ( .A1(n7514), .A2(n7513), .ZN(n7515) );
  XNOR2_X1 U9087 ( .A(n7515), .B(n7762), .ZN(n7517) );
  AND2_X1 U9088 ( .A1(n9095), .A2(n7484), .ZN(n7516) );
  AOI21_X1 U9089 ( .B1(n9195), .B2(n7485), .A(n7516), .ZN(n7518) );
  NAND2_X1 U9090 ( .A1(n7517), .A2(n7518), .ZN(n8441) );
  INV_X1 U9091 ( .A(n7517), .ZN(n7520) );
  INV_X1 U9092 ( .A(n7518), .ZN(n7519) );
  NAND2_X1 U9093 ( .A1(n7520), .A2(n7519), .ZN(n7521) );
  AND2_X1 U9094 ( .A1(n8441), .A2(n7521), .ZN(n8434) );
  AND2_X1 U9095 ( .A1(n8433), .A2(n8434), .ZN(n7522) );
  NAND2_X1 U9096 ( .A1(n8432), .A2(n7522), .ZN(n8431) );
  NAND2_X1 U9097 ( .A1(n8431), .A2(n8441), .ZN(n7544) );
  NAND2_X1 U9098 ( .A1(n7523), .A2(n7642), .ZN(n7526) );
  AOI22_X1 U9099 ( .A1(n8859), .A2(n7566), .B1(n7524), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n7525) );
  NAND2_X1 U9100 ( .A1(n9189), .A2(n4263), .ZN(n7535) );
  NAND2_X1 U9101 ( .A1(n8615), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n7533) );
  NAND2_X1 U9102 ( .A1(n7528), .A2(n7527), .ZN(n7529) );
  AND2_X1 U9103 ( .A1(n7549), .A2(n7529), .ZN(n9089) );
  NAND2_X1 U9104 ( .A1(n7571), .A2(n9089), .ZN(n7532) );
  NAND2_X1 U9105 ( .A1(n5785), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n7531) );
  NAND2_X1 U9106 ( .A1(n7591), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7530) );
  NAND4_X1 U9107 ( .A1(n7533), .A2(n7532), .A3(n7531), .A4(n7530), .ZN(n9115)
         );
  NAND2_X1 U9108 ( .A1(n9115), .A2(n7485), .ZN(n7534) );
  NAND2_X1 U9109 ( .A1(n7535), .A2(n7534), .ZN(n7536) );
  XNOR2_X1 U9110 ( .A(n7536), .B(n7762), .ZN(n7539) );
  AND2_X1 U9111 ( .A1(n9115), .A2(n7484), .ZN(n7537) );
  AOI21_X1 U9112 ( .B1(n9189), .B2(n7485), .A(n7537), .ZN(n7540) );
  NAND2_X1 U9113 ( .A1(n7539), .A2(n7540), .ZN(n7545) );
  INV_X1 U9114 ( .A(n7539), .ZN(n7542) );
  INV_X1 U9115 ( .A(n7540), .ZN(n7541) );
  NAND2_X1 U9116 ( .A1(n7542), .A2(n7541), .ZN(n7543) );
  NAND2_X1 U9117 ( .A1(n8445), .A2(n7545), .ZN(n7560) );
  NAND2_X1 U9118 ( .A1(n7546), .A2(n7642), .ZN(n7548) );
  AOI22_X1 U9119 ( .A1(n8874), .A2(n7566), .B1(n8612), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n7547) );
  NAND2_X1 U9120 ( .A1(n9184), .A2(n4263), .ZN(n7556) );
  NAND2_X1 U9121 ( .A1(n8615), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n7554) );
  INV_X1 U9122 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8483) );
  NAND2_X1 U9123 ( .A1(n7549), .A2(n8483), .ZN(n7550) );
  AND2_X1 U9124 ( .A1(n7569), .A2(n7550), .ZN(n9080) );
  NAND2_X1 U9125 ( .A1(n7571), .A2(n9080), .ZN(n7553) );
  NAND2_X1 U9126 ( .A1(n5785), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n7552) );
  NAND2_X1 U9127 ( .A1(n7591), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7551) );
  NAND4_X1 U9128 ( .A1(n7554), .A2(n7553), .A3(n7552), .A4(n7551), .ZN(n9096)
         );
  NAND2_X1 U9129 ( .A1(n9096), .A2(n7485), .ZN(n7555) );
  NAND2_X1 U9130 ( .A1(n7556), .A2(n7555), .ZN(n7557) );
  XNOR2_X1 U9131 ( .A(n7557), .B(n7762), .ZN(n7561) );
  NAND2_X1 U9132 ( .A1(n7560), .A2(n7561), .ZN(n8479) );
  NAND2_X1 U9133 ( .A1(n9184), .A2(n7485), .ZN(n7559) );
  NAND2_X1 U9134 ( .A1(n9096), .A2(n7484), .ZN(n7558) );
  NAND2_X1 U9135 ( .A1(n7559), .A2(n7558), .ZN(n8482) );
  NAND2_X1 U9136 ( .A1(n8479), .A2(n8482), .ZN(n7564) );
  INV_X1 U9137 ( .A(n7560), .ZN(n7563) );
  INV_X1 U9138 ( .A(n7561), .ZN(n7562) );
  NAND2_X1 U9139 ( .A1(n7563), .A2(n7562), .ZN(n8480) );
  NAND2_X1 U9140 ( .A1(n7565), .A2(n7642), .ZN(n7568) );
  AOI22_X1 U9141 ( .A1(n8612), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n8917), .B2(
        n7566), .ZN(n7567) );
  NAND2_X1 U9142 ( .A1(n8615), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n7575) );
  NAND2_X1 U9143 ( .A1(n7569), .A2(n8409), .ZN(n7570) );
  AND2_X1 U9144 ( .A1(n7589), .A2(n7570), .ZN(n9065) );
  NAND2_X1 U9145 ( .A1(n7571), .A2(n9065), .ZN(n7574) );
  NAND2_X1 U9146 ( .A1(n5785), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n7573) );
  NAND2_X1 U9147 ( .A1(n7591), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n7572) );
  NAND4_X1 U9148 ( .A1(n7575), .A2(n7574), .A3(n7573), .A4(n7572), .ZN(n9073)
         );
  OAI22_X1 U9149 ( .A1(n9068), .A2(n6524), .B1(n9040), .B2(n6011), .ZN(n7576)
         );
  XNOR2_X1 U9150 ( .A(n7576), .B(n7762), .ZN(n7579) );
  OR2_X1 U9151 ( .A1(n9068), .A2(n6011), .ZN(n7578) );
  NAND2_X1 U9152 ( .A1(n9073), .A2(n7484), .ZN(n7577) );
  NAND2_X1 U9153 ( .A1(n7579), .A2(n7580), .ZN(n7585) );
  INV_X1 U9154 ( .A(n7579), .ZN(n7582) );
  INV_X1 U9155 ( .A(n7580), .ZN(n7581) );
  NAND2_X1 U9156 ( .A1(n7582), .A2(n7581), .ZN(n7583) );
  NAND2_X1 U9157 ( .A1(n7585), .A2(n7583), .ZN(n8408) );
  NAND2_X1 U9158 ( .A1(n7586), .A2(n7642), .ZN(n7588) );
  NAND2_X1 U9159 ( .A1(n8612), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7587) );
  NAND2_X1 U9160 ( .A1(n9174), .A2(n4263), .ZN(n7597) );
  NAND2_X1 U9161 ( .A1(n8615), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n7595) );
  NAND2_X1 U9162 ( .A1(n7589), .A2(n9856), .ZN(n7590) );
  NAND2_X1 U9163 ( .A1(n7608), .A2(n7590), .ZN(n8465) );
  INV_X1 U9164 ( .A(n8465), .ZN(n9044) );
  NAND2_X1 U9165 ( .A1(n7571), .A2(n9044), .ZN(n7594) );
  NAND2_X1 U9166 ( .A1(n5785), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n7593) );
  NAND2_X1 U9167 ( .A1(n7591), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n7592) );
  NAND4_X1 U9168 ( .A1(n7595), .A2(n7594), .A3(n7593), .A4(n7592), .ZN(n8809)
         );
  NAND2_X1 U9169 ( .A1(n8809), .A2(n7485), .ZN(n7596) );
  NAND2_X1 U9170 ( .A1(n7597), .A2(n7596), .ZN(n7598) );
  XNOR2_X1 U9171 ( .A(n7598), .B(n7762), .ZN(n7600) );
  AND2_X1 U9172 ( .A1(n8809), .A2(n7484), .ZN(n7599) );
  AOI21_X1 U9173 ( .B1(n9174), .B2(n7485), .A(n7599), .ZN(n7601) );
  INV_X1 U9174 ( .A(n7600), .ZN(n7603) );
  INV_X1 U9175 ( .A(n7601), .ZN(n7602) );
  NAND2_X1 U9176 ( .A1(n7603), .A2(n7602), .ZN(n8462) );
  NAND2_X1 U9177 ( .A1(n7604), .A2(n7642), .ZN(n7606) );
  NAND2_X1 U9178 ( .A1(n8612), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n7605) );
  NAND2_X1 U9179 ( .A1(n9168), .A2(n4263), .ZN(n7616) );
  INV_X1 U9180 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n7607) );
  NAND2_X1 U9181 ( .A1(n7608), .A2(n7607), .ZN(n7609) );
  NAND2_X1 U9182 ( .A1(n7629), .A2(n7609), .ZN(n9020) );
  INV_X1 U9183 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n7610) );
  OAI22_X1 U9184 ( .A1(n9020), .A2(n6026), .B1(n7635), .B2(n7610), .ZN(n7614)
         );
  INV_X1 U9185 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n7612) );
  INV_X1 U9186 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n7611) );
  OAI22_X1 U9187 ( .A1(n7772), .A2(n7612), .B1(n5989), .B2(n7611), .ZN(n7613)
         );
  NAND2_X1 U9188 ( .A1(n9014), .A2(n7485), .ZN(n7615) );
  NAND2_X1 U9189 ( .A1(n7616), .A2(n7615), .ZN(n7617) );
  XNOR2_X1 U9190 ( .A(n7617), .B(n7675), .ZN(n7620) );
  NAND2_X1 U9191 ( .A1(n9168), .A2(n7485), .ZN(n7619) );
  NAND2_X1 U9192 ( .A1(n9014), .A2(n7484), .ZN(n7618) );
  NAND2_X1 U9193 ( .A1(n7619), .A2(n7618), .ZN(n7621) );
  INV_X1 U9194 ( .A(n7620), .ZN(n7623) );
  INV_X1 U9195 ( .A(n7621), .ZN(n7622) );
  NAND2_X1 U9196 ( .A1(n7623), .A2(n7622), .ZN(n8415) );
  NAND2_X1 U9197 ( .A1(n7626), .A2(n7642), .ZN(n7628) );
  NAND2_X1 U9198 ( .A1(n8612), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n7627) );
  NAND2_X1 U9199 ( .A1(n9161), .A2(n7485), .ZN(n7637) );
  INV_X1 U9200 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n7634) );
  AOI22_X1 U9201 ( .A1(n8615), .A2(P1_REG1_REG_22__SCAN_IN), .B1(n5785), .B2(
        P1_REG0_REG_22__SCAN_IN), .ZN(n7633) );
  INV_X1 U9202 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8473) );
  NAND2_X1 U9203 ( .A1(n7629), .A2(n8473), .ZN(n7630) );
  NAND2_X1 U9204 ( .A1(n7631), .A2(n7630), .ZN(n9007) );
  OR2_X1 U9205 ( .A1(n9007), .A2(n6026), .ZN(n7632) );
  OAI211_X1 U9206 ( .C1(n7635), .C2(n7634), .A(n7633), .B(n7632), .ZN(n8808)
         );
  NAND2_X1 U9207 ( .A1(n8808), .A2(n7484), .ZN(n7636) );
  INV_X1 U9208 ( .A(n8808), .ZN(n8418) );
  OAI22_X1 U9209 ( .A1(n9010), .A2(n6524), .B1(n8418), .B2(n6011), .ZN(n7638)
         );
  XNOR2_X1 U9210 ( .A(n7638), .B(n7675), .ZN(n8471) );
  OAI22_X1 U9211 ( .A1(n8994), .A2(n6524), .B1(n8474), .B2(n6011), .ZN(n7639)
         );
  XNOR2_X1 U9212 ( .A(n7639), .B(n7675), .ZN(n7640) );
  NAND2_X1 U9213 ( .A1(n7643), .A2(n7642), .ZN(n7645) );
  NAND2_X1 U9214 ( .A1(n8612), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n7644) );
  INV_X1 U9215 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8455) );
  NAND2_X1 U9216 ( .A1(n7646), .A2(n8455), .ZN(n7647) );
  NAND2_X1 U9217 ( .A1(n7665), .A2(n7647), .ZN(n8985) );
  OR2_X1 U9218 ( .A1(n8985), .A2(n6026), .ZN(n7653) );
  INV_X1 U9219 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n7650) );
  NAND2_X1 U9220 ( .A1(n5785), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n7649) );
  NAND2_X1 U9221 ( .A1(n7591), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n7648) );
  OAI211_X1 U9222 ( .C1(n7772), .C2(n7650), .A(n7649), .B(n7648), .ZN(n7651)
         );
  INV_X1 U9223 ( .A(n7651), .ZN(n7652) );
  OAI22_X1 U9224 ( .A1(n7747), .A2(n6524), .B1(n8399), .B2(n6011), .ZN(n7654)
         );
  XNOR2_X1 U9225 ( .A(n7654), .B(n7762), .ZN(n7658) );
  INV_X1 U9226 ( .A(n8399), .ZN(n8807) );
  NAND2_X1 U9227 ( .A1(n8807), .A2(n7484), .ZN(n7655) );
  NAND2_X1 U9228 ( .A1(n7658), .A2(n7657), .ZN(n7659) );
  OAI21_X1 U9229 ( .B1(n7658), .B2(n7657), .A(n7659), .ZN(n8453) );
  INV_X1 U9230 ( .A(n7659), .ZN(n7660) );
  NAND2_X1 U9231 ( .A1(n8612), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n7662) );
  NAND2_X1 U9232 ( .A1(n9148), .A2(n4263), .ZN(n7674) );
  NAND2_X1 U9233 ( .A1(n7665), .A2(n7664), .ZN(n7666) );
  NAND2_X1 U9234 ( .A1(n8969), .A2(n7571), .ZN(n7672) );
  INV_X1 U9235 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n7669) );
  NAND2_X1 U9236 ( .A1(n5785), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n7668) );
  NAND2_X1 U9237 ( .A1(n7591), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n7667) );
  OAI211_X1 U9238 ( .C1(n7772), .C2(n7669), .A(n7668), .B(n7667), .ZN(n7670)
         );
  INV_X1 U9239 ( .A(n7670), .ZN(n7671) );
  INV_X1 U9240 ( .A(n8501), .ZN(n8979) );
  NAND2_X1 U9241 ( .A1(n8979), .A2(n7485), .ZN(n7673) );
  NAND2_X1 U9242 ( .A1(n7674), .A2(n7673), .ZN(n7676) );
  XNOR2_X1 U9243 ( .A(n7676), .B(n7675), .ZN(n7696) );
  OAI22_X1 U9244 ( .A1(n8972), .A2(n6011), .B1(n8501), .B2(n7677), .ZN(n7695)
         );
  XNOR2_X1 U9245 ( .A(n7696), .B(n7695), .ZN(n8425) );
  NOR2_X1 U9246 ( .A1(n8426), .A2(n8425), .ZN(n8424) );
  NAND2_X1 U9247 ( .A1(n7524), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n7680) );
  NAND2_X1 U9248 ( .A1(n9141), .A2(n4263), .ZN(n7692) );
  NAND2_X1 U9249 ( .A1(n7683), .A2(n7682), .ZN(n7684) );
  NAND2_X1 U9250 ( .A1(n8498), .A2(n7571), .ZN(n7690) );
  INV_X1 U9251 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n7687) );
  NAND2_X1 U9252 ( .A1(n5785), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n7686) );
  NAND2_X1 U9253 ( .A1(n7591), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n7685) );
  OAI211_X1 U9254 ( .C1(n7772), .C2(n7687), .A(n7686), .B(n7685), .ZN(n7688)
         );
  INV_X1 U9255 ( .A(n7688), .ZN(n7689) );
  NAND2_X1 U9256 ( .A1(n8896), .A2(n7485), .ZN(n7691) );
  NAND2_X1 U9257 ( .A1(n7692), .A2(n7691), .ZN(n7693) );
  XNOR2_X1 U9258 ( .A(n7693), .B(n7762), .ZN(n7698) );
  AND2_X1 U9259 ( .A1(n8896), .A2(n7484), .ZN(n7694) );
  AOI21_X1 U9260 ( .B1(n9141), .B2(n7485), .A(n7694), .ZN(n7699) );
  XNOR2_X1 U9261 ( .A(n7698), .B(n7699), .ZN(n8493) );
  NOR2_X1 U9262 ( .A1(n7696), .A2(n7695), .ZN(n8494) );
  INV_X1 U9263 ( .A(n7698), .ZN(n7701) );
  INV_X1 U9264 ( .A(n7699), .ZN(n7700) );
  INV_X1 U9265 ( .A(n7703), .ZN(n7702) );
  INV_X1 U9266 ( .A(n8947), .ZN(n7705) );
  INV_X1 U9267 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n7709) );
  OAI22_X1 U9268 ( .A1(n7705), .A2(n8485), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7709), .ZN(n7719) );
  INV_X1 U9269 ( .A(n7710), .ZN(n7707) );
  AND2_X1 U9270 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P1_REG3_REG_27__SCAN_IN), 
        .ZN(n7706) );
  NAND2_X1 U9271 ( .A1(n7707), .A2(n7706), .ZN(n8916) );
  INV_X1 U9272 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7708) );
  OAI21_X1 U9273 ( .B1(n7710), .B2(n7709), .A(n7708), .ZN(n7711) );
  NAND2_X1 U9274 ( .A1(n8916), .A2(n7711), .ZN(n7778) );
  INV_X1 U9275 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n7714) );
  NAND2_X1 U9276 ( .A1(n5785), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n7713) );
  NAND2_X1 U9277 ( .A1(n7591), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n7712) );
  OAI211_X1 U9278 ( .C1(n7772), .C2(n7714), .A(n7713), .B(n7712), .ZN(n7715)
         );
  INV_X1 U9279 ( .A(n7715), .ZN(n7716) );
  OAI22_X1 U9280 ( .A1(n8953), .A2(n8487), .B1(n8952), .B2(n8500), .ZN(n7718)
         );
  AOI211_X1 U9281 ( .C1(n9136), .C2(n8490), .A(n7719), .B(n7718), .ZN(n7720)
         );
  OAI21_X1 U9282 ( .B1(n7721), .B2(n8519), .A(n7720), .ZN(P1_U3212) );
  OR2_X1 U9283 ( .A1(n9199), .A2(n9113), .ZN(n7722) );
  NAND2_X1 U9284 ( .A1(n7723), .A2(n7722), .ZN(n7724) );
  NAND2_X1 U9285 ( .A1(n7724), .A2(n4814), .ZN(n9103) );
  INV_X1 U9286 ( .A(n9095), .ZN(n8448) );
  OR2_X1 U9287 ( .A1(n9195), .A2(n8448), .ZN(n8684) );
  NAND2_X1 U9288 ( .A1(n9195), .A2(n8448), .ZN(n9092) );
  INV_X1 U9289 ( .A(n9115), .ZN(n8486) );
  NAND2_X1 U9290 ( .A1(n9184), .A2(n9059), .ZN(n8640) );
  NAND2_X1 U9291 ( .A1(n9054), .A2(n8640), .ZN(n9075) );
  NAND2_X1 U9292 ( .A1(n9068), .A2(n9040), .ZN(n7726) );
  AOI22_X1 U9293 ( .A1(n9050), .A2(n7726), .B1(n9073), .B2(n9179), .ZN(n9035)
         );
  NAND2_X1 U9294 ( .A1(n9174), .A2(n8809), .ZN(n7728) );
  NOR2_X1 U9295 ( .A1(n9174), .A2(n8809), .ZN(n7727) );
  AOI21_X1 U9296 ( .B1(n9035), .B2(n7728), .A(n7727), .ZN(n9028) );
  NAND2_X1 U9297 ( .A1(n9168), .A2(n9041), .ZN(n8579) );
  INV_X1 U9298 ( .A(n9168), .ZN(n7729) );
  NAND2_X1 U9299 ( .A1(n9004), .A2(n7730), .ZN(n7731) );
  NAND2_X1 U9300 ( .A1(n7731), .A2(n4812), .ZN(n8989) );
  NAND2_X1 U9301 ( .A1(n8994), .A2(n8474), .ZN(n7733) );
  NOR2_X1 U9302 ( .A1(n8994), .A2(n8474), .ZN(n7732) );
  NAND2_X1 U9303 ( .A1(n7747), .A2(n8399), .ZN(n8960) );
  NAND2_X1 U9304 ( .A1(n8972), .A2(n8501), .ZN(n7734) );
  AND2_X1 U9305 ( .A1(n8960), .A2(n7734), .ZN(n7736) );
  INV_X1 U9306 ( .A(n7734), .ZN(n7735) );
  XNOR2_X1 U9307 ( .A(n8898), .B(n8763), .ZN(n9145) );
  AND2_X1 U9308 ( .A1(n8967), .A2(n9141), .ZN(n7737) );
  NOR2_X1 U9309 ( .A1(n8943), .A2(n7737), .ZN(n9142) );
  INV_X1 U9310 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n7738) );
  OAI22_X1 U9311 ( .A1(n8897), .A2(n9428), .B1(n7738), .B2(n9070), .ZN(n7753)
         );
  NOR2_X1 U9312 ( .A1(n9199), .A2(n8436), .ZN(n8683) );
  NAND2_X1 U9313 ( .A1(n9199), .A2(n8436), .ZN(n8642) );
  INV_X1 U9314 ( .A(n9102), .ZN(n9111) );
  OR2_X1 U9315 ( .A1(n9189), .A2(n8486), .ZN(n8560) );
  NAND2_X1 U9316 ( .A1(n9189), .A2(n8486), .ZN(n8638) );
  NAND2_X1 U9317 ( .A1(n8560), .A2(n8638), .ZN(n8732) );
  INV_X1 U9318 ( .A(n9092), .ZN(n8556) );
  NOR2_X1 U9319 ( .A1(n8732), .A2(n8556), .ZN(n7740) );
  NAND2_X1 U9320 ( .A1(n9109), .A2(n7740), .ZN(n7741) );
  NAND2_X1 U9321 ( .A1(n7741), .A2(n8560), .ZN(n9072) );
  NAND2_X1 U9322 ( .A1(n9072), .A2(n4491), .ZN(n9055) );
  OR2_X1 U9323 ( .A1(n9179), .A2(n9040), .ZN(n8565) );
  NAND2_X1 U9324 ( .A1(n9179), .A2(n9040), .ZN(n9036) );
  NAND2_X1 U9325 ( .A1(n8565), .A2(n9036), .ZN(n9051) );
  INV_X1 U9326 ( .A(n9054), .ZN(n7742) );
  NOR2_X1 U9327 ( .A1(n9051), .A2(n7742), .ZN(n7743) );
  NAND2_X1 U9328 ( .A1(n9055), .A2(n7743), .ZN(n9052) );
  INV_X1 U9329 ( .A(n8809), .ZN(n9061) );
  OR2_X1 U9330 ( .A1(n9174), .A2(n9061), .ZN(n8569) );
  NAND2_X1 U9331 ( .A1(n9174), .A2(n9061), .ZN(n8577) );
  NAND2_X1 U9332 ( .A1(n8569), .A2(n8577), .ZN(n9037) );
  INV_X1 U9333 ( .A(n9036), .ZN(n8637) );
  NOR2_X1 U9334 ( .A1(n9037), .A2(n8637), .ZN(n7744) );
  NAND2_X1 U9335 ( .A1(n9052), .A2(n7744), .ZN(n7745) );
  NAND2_X1 U9336 ( .A1(n7745), .A2(n8569), .ZN(n9021) );
  INV_X1 U9337 ( .A(n9027), .ZN(n8759) );
  NAND2_X1 U9338 ( .A1(n9161), .A2(n8418), .ZN(n8731) );
  OR2_X1 U9339 ( .A1(n9161), .A2(n8418), .ZN(n8995) );
  NAND2_X1 U9340 ( .A1(n9157), .A2(n8474), .ZN(n8729) );
  NAND2_X1 U9341 ( .A1(n7746), .A2(n8729), .ZN(n8977) );
  NAND2_X1 U9342 ( .A1(n9152), .A2(n8399), .ZN(n8962) );
  AND2_X1 U9343 ( .A1(n8704), .A2(n8962), .ZN(n8572) );
  NAND2_X1 U9344 ( .A1(n8907), .A2(n8781), .ZN(n7749) );
  INV_X1 U9345 ( .A(n8763), .ZN(n7748) );
  XNOR2_X1 U9346 ( .A(n7749), .B(n7748), .ZN(n7750) );
  INV_X1 U9347 ( .A(n8899), .ZN(n8806) );
  AOI222_X1 U9348 ( .A1(n9117), .A2(n7750), .B1(n8806), .B2(n9114), .C1(n8979), 
        .C2(n9112), .ZN(n9144) );
  NAND2_X1 U9349 ( .A1(n8498), .A2(n9309), .ZN(n7751) );
  AOI21_X1 U9350 ( .B1(n9144), .B2(n7751), .A(n9321), .ZN(n7752) );
  AOI211_X1 U9351 ( .C1(n9100), .C2(n9142), .A(n7753), .B(n7752), .ZN(n7754)
         );
  OAI21_X1 U9352 ( .B1(n9145), .B2(n9121), .A(n7754), .ZN(P1_U3265) );
  INV_X1 U9353 ( .A(n8521), .ZN(n9272) );
  OAI222_X1 U9354 ( .A1(n4268), .A2(n9272), .B1(n7756), .B2(P2_U3152), .C1(
        n7755), .C2(n8371), .ZN(P2_U3329) );
  NAND2_X1 U9355 ( .A1(n7757), .A2(n7642), .ZN(n7759) );
  NAND2_X1 U9356 ( .A1(n8612), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n7758) );
  NAND2_X1 U9357 ( .A1(n9131), .A2(n7485), .ZN(n7761) );
  INV_X1 U9358 ( .A(n8953), .ZN(n8805) );
  NAND2_X1 U9359 ( .A1(n8805), .A2(n7484), .ZN(n7760) );
  NAND2_X1 U9360 ( .A1(n7761), .A2(n7760), .ZN(n7763) );
  XNOR2_X1 U9361 ( .A(n7763), .B(n7762), .ZN(n7766) );
  NAND2_X1 U9362 ( .A1(n9131), .A2(n4263), .ZN(n7764) );
  OAI21_X1 U9363 ( .B1(n8953), .B2(n6011), .A(n7764), .ZN(n7765) );
  XNOR2_X1 U9364 ( .A(n7766), .B(n7765), .ZN(n7767) );
  INV_X1 U9365 ( .A(n7767), .ZN(n7782) );
  NAND3_X1 U9366 ( .A1(n7782), .A2(n8496), .A3(n7781), .ZN(n7787) );
  AND2_X1 U9367 ( .A1(n7767), .A2(n8496), .ZN(n7768) );
  NAND2_X1 U9368 ( .A1(n7788), .A2(n7768), .ZN(n7786) );
  OR2_X1 U9369 ( .A1(n8899), .A2(n9060), .ZN(n7777) );
  OR2_X1 U9370 ( .A1(n8916), .A2(n6026), .ZN(n7775) );
  INV_X1 U9371 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n7771) );
  NAND2_X1 U9372 ( .A1(n7591), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n7770) );
  NAND2_X1 U9373 ( .A1(n5785), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7769) );
  OAI211_X1 U9374 ( .C1(n7772), .C2(n7771), .A(n7770), .B(n7769), .ZN(n7773)
         );
  INV_X1 U9375 ( .A(n7773), .ZN(n7774) );
  NAND2_X1 U9376 ( .A1(n7775), .A2(n7774), .ZN(n8804) );
  NAND2_X1 U9377 ( .A1(n8804), .A2(n9114), .ZN(n7776) );
  NAND2_X1 U9378 ( .A1(n7777), .A2(n7776), .ZN(n8929) );
  INV_X1 U9379 ( .A(n8929), .ZN(n7780) );
  INV_X1 U9380 ( .A(n7778), .ZN(n8933) );
  AOI22_X1 U9381 ( .A1(n8933), .A2(n8517), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n7779) );
  OAI21_X1 U9382 ( .B1(n7780), .B2(n8511), .A(n7779), .ZN(n7784) );
  NOR3_X1 U9383 ( .A1(n7782), .A2(n8519), .A3(n7781), .ZN(n7783) );
  AOI211_X1 U9384 ( .C1(n9131), .C2(n8490), .A(n7784), .B(n7783), .ZN(n7785)
         );
  OAI211_X1 U9385 ( .C1(n7788), .C2(n7787), .A(n7786), .B(n7785), .ZN(P1_U3218) );
  OAI211_X1 U9386 ( .C1(n7791), .C2(n7790), .A(n7789), .B(n9566), .ZN(n7799)
         );
  AOI22_X1 U9387 ( .A1(n7869), .A2(n7991), .B1(n7792), .B2(n9622), .ZN(n7798)
         );
  INV_X1 U9388 ( .A(n7793), .ZN(n7796) );
  INV_X1 U9389 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7794) );
  OAI22_X1 U9390 ( .A1(n7950), .A2(n9682), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7794), .ZN(n7795) );
  AOI21_X1 U9391 ( .B1(n7796), .B2(n7947), .A(n7795), .ZN(n7797) );
  NAND3_X1 U9392 ( .A1(n7799), .A2(n7798), .A3(n7797), .ZN(P2_U3215) );
  XNOR2_X1 U9393 ( .A(n8349), .B(n7847), .ZN(n7811) );
  INV_X1 U9394 ( .A(n7811), .ZN(n7814) );
  NAND2_X1 U9395 ( .A1(n8228), .A2(n5718), .ZN(n7813) );
  INV_X1 U9396 ( .A(n7800), .ZN(n7801) );
  NAND2_X1 U9397 ( .A1(n7802), .A2(n7801), .ZN(n7908) );
  AND2_X1 U9398 ( .A1(n7984), .A2(n5718), .ZN(n7968) );
  XNOR2_X1 U9399 ( .A(n7976), .B(n7847), .ZN(n7909) );
  XNOR2_X1 U9400 ( .A(n9332), .B(n7803), .ZN(n7804) );
  NAND2_X1 U9401 ( .A1(n7983), .A2(n5718), .ZN(n7805) );
  NAND2_X1 U9402 ( .A1(n7804), .A2(n7805), .ZN(n7912) );
  OAI21_X1 U9403 ( .B1(n7968), .B2(n7909), .A(n7912), .ZN(n7810) );
  NAND3_X1 U9404 ( .A1(n7912), .A2(n7968), .A3(n7909), .ZN(n7808) );
  INV_X1 U9405 ( .A(n7804), .ZN(n7807) );
  INV_X1 U9406 ( .A(n7805), .ZN(n7806) );
  NAND2_X1 U9407 ( .A1(n7807), .A2(n7806), .ZN(n7911) );
  OAI21_X1 U9408 ( .B1(n7908), .B2(n7810), .A(n7809), .ZN(n7921) );
  XNOR2_X1 U9409 ( .A(n7811), .B(n7813), .ZN(n7920) );
  NAND2_X1 U9410 ( .A1(n7921), .A2(n7920), .ZN(n7812) );
  OAI21_X1 U9411 ( .B1(n7814), .B2(n7813), .A(n7812), .ZN(n7952) );
  XNOR2_X1 U9412 ( .A(n8342), .B(n7847), .ZN(n7816) );
  NAND2_X1 U9413 ( .A1(n8208), .A2(n5718), .ZN(n7815) );
  XNOR2_X1 U9414 ( .A(n7816), .B(n7815), .ZN(n7951) );
  INV_X1 U9415 ( .A(n7815), .ZN(n7817) );
  AND2_X1 U9416 ( .A1(n8229), .A2(n5718), .ZN(n7819) );
  XNOR2_X1 U9417 ( .A(n8338), .B(n7847), .ZN(n7818) );
  NOR2_X1 U9418 ( .A1(n7818), .A2(n7819), .ZN(n7820) );
  AOI21_X1 U9419 ( .B1(n7819), .B2(n7818), .A(n7820), .ZN(n7863) );
  XNOR2_X1 U9420 ( .A(n8194), .B(n7847), .ZN(n7822) );
  NAND2_X1 U9421 ( .A1(n8209), .A2(n5718), .ZN(n7821) );
  XNOR2_X1 U9422 ( .A(n7822), .B(n7821), .ZN(n7933) );
  XNOR2_X1 U9423 ( .A(n8327), .B(n7847), .ZN(n7825) );
  NAND2_X1 U9424 ( .A1(n8199), .A2(n5718), .ZN(n7823) );
  XNOR2_X1 U9425 ( .A(n7825), .B(n7823), .ZN(n7890) );
  INV_X1 U9426 ( .A(n7823), .ZN(n7824) );
  XNOR2_X1 U9427 ( .A(n8322), .B(n7847), .ZN(n7828) );
  XNOR2_X1 U9428 ( .A(n7827), .B(n7828), .ZN(n7942) );
  NAND2_X1 U9429 ( .A1(n8183), .A2(n4269), .ZN(n7941) );
  NAND2_X1 U9430 ( .A1(n7942), .A2(n7941), .ZN(n7940) );
  INV_X1 U9431 ( .A(n7827), .ZN(n7829) );
  XNOR2_X1 U9432 ( .A(n8317), .B(n5673), .ZN(n7831) );
  NOR2_X1 U9433 ( .A1(n8166), .A2(n9606), .ZN(n7856) );
  INV_X1 U9434 ( .A(n7831), .ZN(n7832) );
  NOR2_X1 U9435 ( .A1(n7833), .A2(n7832), .ZN(n7834) );
  XNOR2_X1 U9436 ( .A(n8310), .B(n7847), .ZN(n7835) );
  NOR2_X1 U9437 ( .A1(n7903), .A2(n9606), .ZN(n7926) );
  NAND2_X1 U9438 ( .A1(n7927), .A2(n7926), .ZN(n7839) );
  INV_X1 U9439 ( .A(n7835), .ZN(n7836) );
  OR2_X1 U9440 ( .A1(n7837), .A2(n7836), .ZN(n7838) );
  NAND2_X1 U9441 ( .A1(n7839), .A2(n7838), .ZN(n7898) );
  XNOR2_X1 U9442 ( .A(n8306), .B(n7847), .ZN(n7842) );
  NAND2_X1 U9443 ( .A1(n8132), .A2(n5718), .ZN(n7840) );
  INV_X1 U9444 ( .A(n7840), .ZN(n7841) );
  NAND2_X1 U9445 ( .A1(n7842), .A2(n7841), .ZN(n7843) );
  XNOR2_X1 U9446 ( .A(n8301), .B(n7847), .ZN(n7846) );
  NAND2_X1 U9447 ( .A1(n8119), .A2(n4269), .ZN(n7844) );
  XNOR2_X1 U9448 ( .A(n7846), .B(n7844), .ZN(n7960) );
  INV_X1 U9449 ( .A(n7844), .ZN(n7845) );
  XNOR2_X1 U9450 ( .A(n8296), .B(n7847), .ZN(n7874) );
  NAND2_X1 U9451 ( .A1(n8107), .A2(n4269), .ZN(n7872) );
  XNOR2_X1 U9452 ( .A(n7877), .B(n7876), .ZN(n7854) );
  OAI22_X1 U9453 ( .A1(n7849), .A2(n7970), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7848), .ZN(n7852) );
  INV_X1 U9454 ( .A(n8087), .ZN(n7850) );
  OAI22_X1 U9455 ( .A1(n7973), .A2(n7901), .B1(n9571), .B2(n7850), .ZN(n7851)
         );
  AOI211_X1 U9456 ( .C1(n8296), .C2(n9565), .A(n7852), .B(n7851), .ZN(n7853)
         );
  OAI21_X1 U9457 ( .B1(n7854), .B2(n7978), .A(n7853), .ZN(P2_U3216) );
  XNOR2_X1 U9458 ( .A(n7855), .B(n7856), .ZN(n7861) );
  OAI22_X1 U9459 ( .A1(n7970), .A2(n7903), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7857), .ZN(n7859) );
  OAI22_X1 U9460 ( .A1(n7973), .A2(n7892), .B1(n9571), .B2(n8149), .ZN(n7858)
         );
  AOI211_X1 U9461 ( .C1(n8317), .C2(n9565), .A(n7859), .B(n7858), .ZN(n7860)
         );
  OAI21_X1 U9462 ( .B1(n7861), .B2(n7978), .A(n7860), .ZN(P2_U3218) );
  OAI21_X1 U9463 ( .B1(n7864), .B2(n7863), .A(n7862), .ZN(n7865) );
  NAND2_X1 U9464 ( .A1(n7865), .A2(n9566), .ZN(n7871) );
  NAND2_X1 U9465 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8070) );
  INV_X1 U9466 ( .A(n8070), .ZN(n7868) );
  INV_X1 U9467 ( .A(n8212), .ZN(n7866) );
  OAI22_X1 U9468 ( .A1(n7973), .A2(n8250), .B1(n9571), .B2(n7866), .ZN(n7867)
         );
  AOI211_X1 U9469 ( .C1(n7869), .C2(n8209), .A(n7868), .B(n7867), .ZN(n7870)
         );
  OAI211_X1 U9470 ( .C1(n8205), .C2(n7950), .A(n7871), .B(n7870), .ZN(P2_U3221) );
  INV_X1 U9471 ( .A(n7872), .ZN(n7873) );
  AOI21_X1 U9472 ( .B1(n7877), .B2(n7876), .A(n7875), .ZN(n7881) );
  NAND2_X1 U9473 ( .A1(n8092), .A2(n5718), .ZN(n7878) );
  XOR2_X1 U9474 ( .A(n7847), .B(n7878), .Z(n7879) );
  XNOR2_X1 U9475 ( .A(n8290), .B(n7879), .ZN(n7880) );
  XNOR2_X1 U9476 ( .A(n7881), .B(n7880), .ZN(n7888) );
  OAI22_X1 U9477 ( .A1(n7962), .A2(n7973), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7882), .ZN(n7886) );
  OAI22_X1 U9478 ( .A1(n7970), .A2(n7884), .B1(n9571), .B2(n7883), .ZN(n7885)
         );
  AOI211_X1 U9479 ( .C1(n8290), .C2(n9565), .A(n7886), .B(n7885), .ZN(n7887)
         );
  OAI21_X1 U9480 ( .B1(n7888), .B2(n7978), .A(n7887), .ZN(P2_U3222) );
  XNOR2_X1 U9481 ( .A(n7889), .B(n7890), .ZN(n7897) );
  OAI22_X1 U9482 ( .A1(n7970), .A2(n7892), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7891), .ZN(n7895) );
  INV_X1 U9483 ( .A(n8209), .ZN(n7893) );
  OAI22_X1 U9484 ( .A1(n7973), .A2(n7893), .B1(n9571), .B2(n8174), .ZN(n7894)
         );
  AOI211_X1 U9485 ( .C1(n8327), .C2(n9565), .A(n7895), .B(n7894), .ZN(n7896)
         );
  OAI21_X1 U9486 ( .B1(n7897), .B2(n7978), .A(n7896), .ZN(P2_U3225) );
  XNOR2_X1 U9487 ( .A(n7898), .B(n7899), .ZN(n7907) );
  OAI22_X1 U9488 ( .A1(n7970), .A2(n7901), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7900), .ZN(n7905) );
  INV_X1 U9489 ( .A(n8114), .ZN(n7902) );
  OAI22_X1 U9490 ( .A1(n7973), .A2(n7903), .B1(n9571), .B2(n7902), .ZN(n7904)
         );
  AOI211_X1 U9491 ( .C1(n8306), .C2(n9565), .A(n7905), .B(n7904), .ZN(n7906)
         );
  OAI21_X1 U9492 ( .B1(n7907), .B2(n7978), .A(n7906), .ZN(P2_U3227) );
  XNOR2_X1 U9493 ( .A(n7908), .B(n7909), .ZN(n7969) );
  INV_X1 U9494 ( .A(n7908), .ZN(n7910) );
  AOI22_X1 U9495 ( .A1(n7969), .A2(n7968), .B1(n7910), .B2(n7909), .ZN(n7914)
         );
  NAND2_X1 U9496 ( .A1(n7912), .A2(n7911), .ZN(n7913) );
  XNOR2_X1 U9497 ( .A(n7914), .B(n7913), .ZN(n7919) );
  OAI22_X1 U9498 ( .A1(n7915), .A2(n8249), .B1(n7954), .B2(n8251), .ZN(n9328)
         );
  NOR2_X1 U9499 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9805), .ZN(n8015) );
  AOI21_X1 U9500 ( .B1(n9559), .B2(n9328), .A(n8015), .ZN(n7916) );
  OAI21_X1 U9501 ( .B1(n9330), .B2(n9571), .A(n7916), .ZN(n7917) );
  AOI21_X1 U9502 ( .B1(n9332), .B2(n9565), .A(n7917), .ZN(n7918) );
  OAI21_X1 U9503 ( .B1(n7919), .B2(n7978), .A(n7918), .ZN(P2_U3228) );
  XNOR2_X1 U9504 ( .A(n7921), .B(n7920), .ZN(n7925) );
  OAI22_X1 U9505 ( .A1(n7970), .A2(n8250), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7061), .ZN(n7923) );
  OAI22_X1 U9506 ( .A1(n7973), .A2(n8248), .B1(n9571), .B2(n8239), .ZN(n7922)
         );
  AOI211_X1 U9507 ( .C1(n8349), .C2(n9565), .A(n7923), .B(n7922), .ZN(n7924)
         );
  OAI21_X1 U9508 ( .B1(n7925), .B2(n7978), .A(n7924), .ZN(P2_U3230) );
  XNOR2_X1 U9509 ( .A(n7927), .B(n7926), .ZN(n7932) );
  OAI22_X1 U9510 ( .A1(n7970), .A2(n7963), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7928), .ZN(n7930) );
  OAI22_X1 U9511 ( .A1(n7973), .A2(n8166), .B1(n9571), .B2(n8135), .ZN(n7929)
         );
  AOI211_X1 U9512 ( .C1(n8310), .C2(n9565), .A(n7930), .B(n7929), .ZN(n7931)
         );
  OAI21_X1 U9513 ( .B1(n7932), .B2(n7978), .A(n7931), .ZN(P2_U3231) );
  XNOR2_X1 U9514 ( .A(n7934), .B(n7933), .ZN(n7939) );
  OAI22_X1 U9515 ( .A1(n7970), .A2(n8165), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7935), .ZN(n7937) );
  OAI22_X1 U9516 ( .A1(n7973), .A2(n7953), .B1(n9571), .B2(n8191), .ZN(n7936)
         );
  AOI211_X1 U9517 ( .C1(n8332), .C2(n9565), .A(n7937), .B(n7936), .ZN(n7938)
         );
  OAI21_X1 U9518 ( .B1(n7939), .B2(n7978), .A(n7938), .ZN(P2_U3235) );
  OAI21_X1 U9519 ( .B1(n7942), .B2(n7941), .A(n7940), .ZN(n7943) );
  NAND2_X1 U9520 ( .A1(n7943), .A2(n9566), .ZN(n7949) );
  NOR2_X1 U9521 ( .A1(n7973), .A2(n8165), .ZN(n7946) );
  OAI22_X1 U9522 ( .A1(n7970), .A2(n8166), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7944), .ZN(n7945) );
  AOI211_X1 U9523 ( .C1(n7947), .C2(n8158), .A(n7946), .B(n7945), .ZN(n7948)
         );
  OAI211_X1 U9524 ( .C1(n8160), .C2(n7950), .A(n7949), .B(n7948), .ZN(P2_U3237) );
  XNOR2_X1 U9525 ( .A(n7952), .B(n7951), .ZN(n7958) );
  NAND2_X1 U9526 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8046) );
  OAI21_X1 U9527 ( .B1(n7970), .B2(n7953), .A(n8046), .ZN(n7956) );
  OAI22_X1 U9528 ( .A1(n7973), .A2(n7954), .B1(n9571), .B2(n8223), .ZN(n7955)
         );
  AOI211_X1 U9529 ( .C1(n8342), .C2(n9565), .A(n7956), .B(n7955), .ZN(n7957)
         );
  OAI21_X1 U9530 ( .B1(n7958), .B2(n7978), .A(n7957), .ZN(P2_U3240) );
  XNOR2_X1 U9531 ( .A(n7959), .B(n7960), .ZN(n7967) );
  OAI22_X1 U9532 ( .A1(n7962), .A2(n7970), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7961), .ZN(n7965) );
  OAI22_X1 U9533 ( .A1(n7973), .A2(n7963), .B1(n9571), .B2(n8101), .ZN(n7964)
         );
  AOI211_X1 U9534 ( .C1(n8301), .C2(n9565), .A(n7965), .B(n7964), .ZN(n7966)
         );
  OAI21_X1 U9535 ( .B1(n7967), .B2(n7978), .A(n7966), .ZN(P2_U3242) );
  XNOR2_X1 U9536 ( .A(n7969), .B(n7968), .ZN(n7979) );
  OAI22_X1 U9537 ( .A1(n7970), .A2(n8248), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6902), .ZN(n7975) );
  OAI22_X1 U9538 ( .A1(n7973), .A2(n7972), .B1(n9571), .B2(n7971), .ZN(n7974)
         );
  AOI211_X1 U9539 ( .C1(n7976), .C2(n9565), .A(n7975), .B(n7974), .ZN(n7977)
         );
  OAI21_X1 U9540 ( .B1(n7979), .B2(n7978), .A(n7977), .ZN(P2_U3243) );
  MUX2_X1 U9541 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n7980), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U9542 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n7981), .S(P2_U3966), .Z(
        P2_U3581) );
  MUX2_X1 U9543 ( .A(n8092), .B(P2_DATAO_REG_28__SCAN_IN), .S(n7982), .Z(
        P2_U3580) );
  MUX2_X1 U9544 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8107), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U9545 ( .A(n8119), .B(P2_DATAO_REG_26__SCAN_IN), .S(n7982), .Z(
        P2_U3578) );
  MUX2_X1 U9546 ( .A(n8132), .B(P2_DATAO_REG_25__SCAN_IN), .S(n7982), .Z(
        P2_U3577) );
  MUX2_X1 U9547 ( .A(n8144), .B(P2_DATAO_REG_24__SCAN_IN), .S(n7982), .Z(
        P2_U3576) );
  INV_X1 U9548 ( .A(n8166), .ZN(n8131) );
  MUX2_X1 U9549 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8131), .S(P2_U3966), .Z(
        P2_U3575) );
  MUX2_X1 U9550 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8183), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U9551 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8199), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U9552 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8209), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U9553 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8229), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U9554 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8208), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U9555 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8228), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9556 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n7983), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9557 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n7984), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9558 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n7985), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9559 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n7986), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9560 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n7987), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U9561 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n7988), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U9562 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n7989), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U9563 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n7990), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U9564 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n7991), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U9565 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n7992), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U9566 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n9622), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U9567 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n7993), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U9568 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n9623), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U9569 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n7994), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U9570 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n5924), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U9571 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n7995), .S(P2_U3966), .Z(
        P2_U3553) );
  OAI21_X1 U9572 ( .B1(n8000), .B2(P2_REG2_REG_14__SCAN_IN), .A(n7996), .ZN(
        n8018) );
  XOR2_X1 U9573 ( .A(n8019), .B(n8018), .Z(n7997) );
  NAND2_X1 U9574 ( .A1(n7997), .A2(n6994), .ZN(n8020) );
  OAI21_X1 U9575 ( .B1(n7997), .B2(n6994), .A(n8020), .ZN(n7998) );
  NAND2_X1 U9576 ( .A1(n7998), .A2(n9572), .ZN(n8009) );
  INV_X1 U9577 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8006) );
  OAI21_X1 U9578 ( .B1(n8000), .B2(P2_REG1_REG_14__SCAN_IN), .A(n7999), .ZN(
        n8010) );
  XNOR2_X1 U9579 ( .A(n8019), .B(n8010), .ZN(n8001) );
  INV_X1 U9580 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9373) );
  NAND2_X1 U9581 ( .A1(n8001), .A2(n9373), .ZN(n8003) );
  NOR2_X1 U9582 ( .A1(n9373), .A2(n8001), .ZN(n8011) );
  INV_X1 U9583 ( .A(n8011), .ZN(n8002) );
  NAND3_X1 U9584 ( .A1(n9573), .A2(n8003), .A3(n8002), .ZN(n8005) );
  NAND2_X1 U9585 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8004) );
  OAI211_X1 U9586 ( .C1(n8072), .C2(n8006), .A(n8005), .B(n8004), .ZN(n8007)
         );
  INV_X1 U9587 ( .A(n8007), .ZN(n8008) );
  OAI211_X1 U9588 ( .C1(n9575), .C2(n8019), .A(n8009), .B(n8008), .ZN(P2_U3260) );
  NOR2_X1 U9589 ( .A1(n8019), .A2(n8010), .ZN(n8012) );
  NOR2_X1 U9590 ( .A1(n8012), .A2(n8011), .ZN(n8014) );
  AOI22_X1 U9591 ( .A1(n8034), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n6983), .B2(
        n8017), .ZN(n8013) );
  NAND2_X1 U9592 ( .A1(n8013), .A2(n8014), .ZN(n8029) );
  OAI21_X1 U9593 ( .B1(n8014), .B2(n8013), .A(n8029), .ZN(n8027) );
  AOI21_X1 U9594 ( .B1(n9578), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8015), .ZN(
        n8016) );
  OAI21_X1 U9595 ( .B1(n9575), .B2(n8017), .A(n8016), .ZN(n8026) );
  NAND2_X1 U9596 ( .A1(n8019), .A2(n8018), .ZN(n8021) );
  NAND2_X1 U9597 ( .A1(n8021), .A2(n8020), .ZN(n8024) );
  NAND2_X1 U9598 ( .A1(n8034), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8022) );
  OAI21_X1 U9599 ( .B1(n8034), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8022), .ZN(
        n8023) );
  NOR2_X1 U9600 ( .A1(n8023), .A2(n8024), .ZN(n8033) );
  AOI211_X1 U9601 ( .C1(n8024), .C2(n8023), .A(n8033), .B(n9576), .ZN(n8025)
         );
  AOI211_X1 U9602 ( .C1(n8027), .C2(n9573), .A(n8026), .B(n8025), .ZN(n8028)
         );
  INV_X1 U9603 ( .A(n8028), .ZN(P2_U3261) );
  OAI21_X1 U9604 ( .B1(n8034), .B2(P2_REG1_REG_16__SCAN_IN), .A(n8029), .ZN(
        n8032) );
  XNOR2_X1 U9605 ( .A(n8050), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8031) );
  NOR2_X1 U9606 ( .A1(n8031), .A2(n8032), .ZN(n8049) );
  AOI211_X1 U9607 ( .C1(n8032), .C2(n8031), .A(n8049), .B(n8030), .ZN(n8043)
         );
  NAND2_X1 U9608 ( .A1(n8050), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8035) );
  OAI21_X1 U9609 ( .B1(n8050), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8035), .ZN(
        n8036) );
  AOI211_X1 U9610 ( .C1(n8037), .C2(n8036), .A(n8044), .B(n9576), .ZN(n8042)
         );
  INV_X1 U9611 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8040) );
  NAND2_X1 U9612 ( .A1(n9295), .A2(n8050), .ZN(n8039) );
  NAND2_X1 U9613 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3152), .ZN(n8038) );
  OAI211_X1 U9614 ( .C1(n8072), .C2(n8040), .A(n8039), .B(n8038), .ZN(n8041)
         );
  OR3_X1 U9615 ( .A1(n8043), .A2(n8042), .A3(n8041), .ZN(P2_U3262) );
  INV_X1 U9616 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8224) );
  NAND2_X1 U9617 ( .A1(n8045), .A2(n8224), .ZN(n8058) );
  OAI21_X1 U9618 ( .B1(n8045), .B2(n8224), .A(n8058), .ZN(n8055) );
  INV_X1 U9619 ( .A(n8046), .ZN(n8047) );
  AOI21_X1 U9620 ( .B1(n9578), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8047), .ZN(
        n8053) );
  XNOR2_X1 U9621 ( .A(n8048), .B(n8062), .ZN(n8064) );
  AOI21_X1 U9622 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8050), .A(n8049), .ZN(
        n8063) );
  XNOR2_X1 U9623 ( .A(n8064), .B(n8063), .ZN(n8051) );
  NAND2_X1 U9624 ( .A1(n9573), .A2(n8051), .ZN(n8052) );
  OAI211_X1 U9625 ( .C1(n9575), .C2(n4668), .A(n8053), .B(n8052), .ZN(n8054)
         );
  AOI21_X1 U9626 ( .B1(n9572), .B2(n8055), .A(n8054), .ZN(n8056) );
  INV_X1 U9627 ( .A(n8056), .ZN(P2_U3263) );
  INV_X1 U9628 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8071) );
  NAND2_X1 U9629 ( .A1(n8057), .A2(n4668), .ZN(n8059) );
  NAND2_X1 U9630 ( .A1(n8059), .A2(n8058), .ZN(n8060) );
  XOR2_X1 U9631 ( .A(n8061), .B(n8060), .Z(n8067) );
  AOI22_X1 U9632 ( .A1(n8064), .A2(n8063), .B1(n4668), .B2(n8062), .ZN(n8065)
         );
  XNOR2_X1 U9633 ( .A(n8065), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8068) );
  INV_X1 U9634 ( .A(n8068), .ZN(n8066) );
  AOI22_X1 U9635 ( .A1(n8067), .A2(n9572), .B1(n8066), .B2(n9573), .ZN(n8069)
         );
  NAND2_X1 U9636 ( .A1(n8285), .A2(n8079), .ZN(n8281) );
  XNOR2_X1 U9637 ( .A(n8281), .B(n8272), .ZN(n8274) );
  NAND2_X1 U9638 ( .A1(n8074), .A2(n8073), .ZN(n8283) );
  NOR2_X1 U9639 ( .A1(n9590), .A2(n8283), .ZN(n8082) );
  NOR2_X1 U9640 ( .A1(n8075), .A2(n8237), .ZN(n8076) );
  AOI211_X1 U9641 ( .C1(n8217), .C2(P2_REG2_REG_31__SCAN_IN), .A(n8082), .B(
        n8076), .ZN(n8077) );
  OAI21_X1 U9642 ( .B1(n8274), .B2(n8078), .A(n8077), .ZN(P2_U3265) );
  INV_X1 U9643 ( .A(n8079), .ZN(n8080) );
  NAND2_X1 U9644 ( .A1(n8081), .A2(n8080), .ZN(n8282) );
  NAND3_X1 U9645 ( .A1(n8282), .A2(n9337), .A3(n8281), .ZN(n8084) );
  AOI21_X1 U9646 ( .B1(n8217), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8082), .ZN(
        n8083) );
  OAI211_X1 U9647 ( .C1(n8285), .C2(n8237), .A(n8084), .B(n8083), .ZN(P2_U3266) );
  XOR2_X1 U9648 ( .A(n8091), .B(n8085), .Z(n8299) );
  AOI211_X1 U9649 ( .C1(n8296), .C2(n8098), .A(n4269), .B(n8086), .ZN(n8295)
         );
  INV_X1 U9650 ( .A(n8296), .ZN(n8089) );
  AOI22_X1 U9651 ( .A1(n8217), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8087), .B2(
        n9613), .ZN(n8088) );
  OAI21_X1 U9652 ( .B1(n8089), .B2(n8237), .A(n8088), .ZN(n8095) );
  XOR2_X1 U9653 ( .A(n8090), .B(n8091), .Z(n8093) );
  AOI222_X1 U9654 ( .A1(n9619), .A2(n8093), .B1(n8119), .B2(n9624), .C1(n8092), 
        .C2(n9621), .ZN(n8298) );
  NOR2_X1 U9655 ( .A1(n8298), .A2(n8217), .ZN(n8094) );
  AOI211_X1 U9656 ( .C1(n9600), .C2(n8295), .A(n8095), .B(n8094), .ZN(n8096)
         );
  OAI21_X1 U9657 ( .B1(n8299), .B2(n8254), .A(n8096), .ZN(P2_U3269) );
  XNOR2_X1 U9658 ( .A(n8097), .B(n4803), .ZN(n8304) );
  INV_X1 U9659 ( .A(n8113), .ZN(n8100) );
  INV_X1 U9660 ( .A(n8098), .ZN(n8099) );
  AOI211_X1 U9661 ( .C1(n8301), .C2(n8100), .A(n4269), .B(n8099), .ZN(n8300)
         );
  NOR2_X1 U9662 ( .A1(n9590), .A2(n5547), .ZN(n8243) );
  INV_X1 U9663 ( .A(n8101), .ZN(n8102) );
  AOI22_X1 U9664 ( .A1(n9590), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n8102), .B2(
        n9613), .ZN(n8103) );
  OAI21_X1 U9665 ( .B1(n8104), .B2(n8237), .A(n8103), .ZN(n8110) );
  XNOR2_X1 U9666 ( .A(n8105), .B(n8106), .ZN(n8108) );
  AOI222_X1 U9667 ( .A1(n9619), .A2(n8108), .B1(n8107), .B2(n9621), .C1(n8132), 
        .C2(n9624), .ZN(n8303) );
  NOR2_X1 U9668 ( .A1(n8303), .A2(n8217), .ZN(n8109) );
  AOI211_X1 U9669 ( .C1(n8300), .C2(n8243), .A(n8110), .B(n8109), .ZN(n8111)
         );
  OAI21_X1 U9670 ( .B1(n8304), .B2(n8254), .A(n8111), .ZN(P2_U3270) );
  XOR2_X1 U9671 ( .A(n8118), .B(n8112), .Z(n8309) );
  AOI211_X1 U9672 ( .C1(n8306), .C2(n4331), .A(n5718), .B(n8113), .ZN(n8305)
         );
  INV_X1 U9673 ( .A(n8306), .ZN(n8116) );
  AOI22_X1 U9674 ( .A1(n8217), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8114), .B2(
        n9613), .ZN(n8115) );
  OAI21_X1 U9675 ( .B1(n8116), .B2(n8237), .A(n8115), .ZN(n8122) );
  XOR2_X1 U9676 ( .A(n8118), .B(n8117), .Z(n8120) );
  AOI222_X1 U9677 ( .A1(n9619), .A2(n8120), .B1(n8119), .B2(n9621), .C1(n8144), 
        .C2(n9624), .ZN(n8308) );
  NOR2_X1 U9678 ( .A1(n8308), .A2(n8217), .ZN(n8121) );
  AOI211_X1 U9679 ( .C1(n8243), .C2(n8305), .A(n8122), .B(n8121), .ZN(n8123)
         );
  OAI21_X1 U9680 ( .B1(n8309), .B2(n8254), .A(n8123), .ZN(P2_U3271) );
  AOI21_X1 U9681 ( .B1(n8126), .B2(n8125), .A(n8124), .ZN(n8314) );
  NAND2_X1 U9682 ( .A1(n8128), .A2(n8127), .ZN(n8129) );
  NAND3_X1 U9683 ( .A1(n8130), .A2(n9619), .A3(n8129), .ZN(n8134) );
  AOI22_X1 U9684 ( .A1(n8132), .A2(n9621), .B1(n8131), .B2(n9624), .ZN(n8133)
         );
  AND2_X1 U9685 ( .A1(n8134), .A2(n8133), .ZN(n8313) );
  INV_X1 U9686 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8136) );
  OAI22_X1 U9687 ( .A1(n8265), .A2(n8136), .B1(n8135), .B2(n8238), .ZN(n8137)
         );
  AOI21_X1 U9688 ( .B1(n8310), .B2(n9591), .A(n8137), .ZN(n8139) );
  XNOR2_X1 U9689 ( .A(n8148), .B(n8310), .ZN(n8311) );
  NAND2_X1 U9690 ( .A1(n8311), .A2(n9337), .ZN(n8138) );
  OAI211_X1 U9691 ( .C1(n8313), .C2(n9590), .A(n8139), .B(n8138), .ZN(n8140)
         );
  INV_X1 U9692 ( .A(n8140), .ZN(n8141) );
  OAI21_X1 U9693 ( .B1(n8314), .B2(n8254), .A(n8141), .ZN(P2_U3272) );
  OAI21_X1 U9694 ( .B1(n4302), .B2(n8143), .A(n8142), .ZN(n8145) );
  AOI222_X1 U9695 ( .A1(n9619), .A2(n8145), .B1(n8183), .B2(n9624), .C1(n8144), 
        .C2(n9621), .ZN(n8320) );
  OR2_X1 U9696 ( .A1(n8147), .A2(n8146), .ZN(n8316) );
  NAND3_X1 U9697 ( .A1(n8316), .A2(n8315), .A3(n9601), .ZN(n8154) );
  AOI21_X1 U9698 ( .B1(n8317), .B2(n8156), .A(n8148), .ZN(n8318) );
  INV_X1 U9699 ( .A(n8149), .ZN(n8150) );
  AOI22_X1 U9700 ( .A1(n8217), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8150), .B2(
        n9613), .ZN(n8151) );
  OAI21_X1 U9701 ( .B1(n4428), .B2(n8237), .A(n8151), .ZN(n8152) );
  AOI21_X1 U9702 ( .B1(n8318), .B2(n9337), .A(n8152), .ZN(n8153) );
  OAI211_X1 U9703 ( .C1(n8217), .C2(n8320), .A(n8154), .B(n8153), .ZN(P2_U3273) );
  XOR2_X1 U9704 ( .A(n8155), .B(n8163), .Z(n8326) );
  AOI21_X1 U9705 ( .B1(n8322), .B2(n8157), .A(n4429), .ZN(n8323) );
  AOI22_X1 U9706 ( .A1(n8217), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8158), .B2(
        n9613), .ZN(n8159) );
  OAI21_X1 U9707 ( .B1(n8160), .B2(n8237), .A(n8159), .ZN(n8171) );
  NAND2_X1 U9708 ( .A1(n8180), .A2(n8162), .ZN(n8164) );
  AOI21_X1 U9709 ( .B1(n8164), .B2(n8163), .A(n9345), .ZN(n8169) );
  OAI22_X1 U9710 ( .A1(n8166), .A2(n8251), .B1(n8165), .B2(n8249), .ZN(n8167)
         );
  AOI21_X1 U9711 ( .B1(n8169), .B2(n8168), .A(n8167), .ZN(n8325) );
  NOR2_X1 U9712 ( .A1(n8325), .A2(n8217), .ZN(n8170) );
  AOI211_X1 U9713 ( .C1(n8323), .C2(n9337), .A(n8171), .B(n8170), .ZN(n8172)
         );
  OAI21_X1 U9714 ( .B1(n8326), .B2(n8254), .A(n8172), .ZN(P2_U3274) );
  XOR2_X1 U9715 ( .A(n8173), .B(n8179), .Z(n8331) );
  XNOR2_X1 U9716 ( .A(n8177), .B(n8189), .ZN(n8328) );
  INV_X1 U9717 ( .A(n8174), .ZN(n8175) );
  AOI22_X1 U9718 ( .A1(n8217), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8175), .B2(
        n9613), .ZN(n8176) );
  OAI21_X1 U9719 ( .B1(n8177), .B2(n8237), .A(n8176), .ZN(n8186) );
  INV_X1 U9720 ( .A(n8178), .ZN(n8182) );
  INV_X1 U9721 ( .A(n8179), .ZN(n8181) );
  OAI21_X1 U9722 ( .B1(n8182), .B2(n8181), .A(n8180), .ZN(n8184) );
  AOI222_X1 U9723 ( .A1(n9619), .A2(n8184), .B1(n8183), .B2(n9621), .C1(n8209), 
        .C2(n9624), .ZN(n8330) );
  NOR2_X1 U9724 ( .A1(n8330), .A2(n8217), .ZN(n8185) );
  AOI211_X1 U9725 ( .C1(n8328), .C2(n9337), .A(n8186), .B(n8185), .ZN(n8187)
         );
  OAI21_X1 U9726 ( .B1(n8331), .B2(n8254), .A(n8187), .ZN(P2_U3275) );
  XNOR2_X1 U9727 ( .A(n8188), .B(n8198), .ZN(n8336) );
  INV_X1 U9728 ( .A(n8189), .ZN(n8190) );
  AOI21_X1 U9729 ( .B1(n8332), .B2(n4447), .A(n8190), .ZN(n8333) );
  INV_X1 U9730 ( .A(n8191), .ZN(n8192) );
  AOI22_X1 U9731 ( .A1(n8217), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8192), .B2(
        n9613), .ZN(n8193) );
  OAI21_X1 U9732 ( .B1(n8194), .B2(n8237), .A(n8193), .ZN(n8202) );
  NAND2_X1 U9733 ( .A1(n8195), .A2(n8196), .ZN(n8197) );
  XOR2_X1 U9734 ( .A(n8198), .B(n8197), .Z(n8200) );
  AOI222_X1 U9735 ( .A1(n9619), .A2(n8200), .B1(n8199), .B2(n9621), .C1(n8229), 
        .C2(n9624), .ZN(n8335) );
  NOR2_X1 U9736 ( .A1(n8335), .A2(n8217), .ZN(n8201) );
  AOI211_X1 U9737 ( .C1(n8333), .C2(n9337), .A(n8202), .B(n8201), .ZN(n8203)
         );
  OAI21_X1 U9738 ( .B1(n8254), .B2(n8336), .A(n8203), .ZN(P2_U3276) );
  XOR2_X1 U9739 ( .A(n8204), .B(n8207), .Z(n8341) );
  NOR2_X1 U9740 ( .A1(n8205), .A2(n8237), .ZN(n8216) );
  OAI21_X1 U9741 ( .B1(n8207), .B2(n8206), .A(n8195), .ZN(n8210) );
  AOI222_X1 U9742 ( .A1(n9619), .A2(n8210), .B1(n8209), .B2(n9621), .C1(n8208), 
        .C2(n9624), .ZN(n8340) );
  AOI211_X1 U9743 ( .C1(n8338), .C2(n8220), .A(n5718), .B(n8211), .ZN(n8337)
         );
  AOI22_X1 U9744 ( .A1(n8337), .A2(n8213), .B1(n9613), .B2(n8212), .ZN(n8214)
         );
  AOI21_X1 U9745 ( .B1(n8340), .B2(n8214), .A(n9590), .ZN(n8215) );
  AOI211_X1 U9746 ( .C1(n8217), .C2(P2_REG2_REG_19__SCAN_IN), .A(n8216), .B(
        n8215), .ZN(n8218) );
  OAI21_X1 U9747 ( .B1(n8341), .B2(n8254), .A(n8218), .ZN(P2_U3277) );
  XNOR2_X1 U9748 ( .A(n8219), .B(n4282), .ZN(n8346) );
  INV_X1 U9749 ( .A(n8220), .ZN(n8221) );
  AOI21_X1 U9750 ( .B1(n8342), .B2(n8235), .A(n8221), .ZN(n8343) );
  NOR2_X1 U9751 ( .A1(n8222), .A2(n8237), .ZN(n8226) );
  OAI22_X1 U9752 ( .A1(n8265), .A2(n8224), .B1(n8223), .B2(n8238), .ZN(n8225)
         );
  AOI211_X1 U9753 ( .C1(n8343), .C2(n9337), .A(n8226), .B(n8225), .ZN(n8232)
         );
  OAI21_X1 U9754 ( .B1(n4339), .B2(n4282), .A(n8227), .ZN(n8230) );
  AOI222_X1 U9755 ( .A1(n9619), .A2(n8230), .B1(n8229), .B2(n9621), .C1(n8228), 
        .C2(n9624), .ZN(n8345) );
  OR2_X1 U9756 ( .A1(n8345), .A2(n8217), .ZN(n8231) );
  OAI211_X1 U9757 ( .C1(n8346), .C2(n8254), .A(n8232), .B(n8231), .ZN(P2_U3278) );
  XNOR2_X1 U9758 ( .A(n8233), .B(n8245), .ZN(n8351) );
  INV_X1 U9759 ( .A(n8234), .ZN(n9334) );
  INV_X1 U9760 ( .A(n8235), .ZN(n8236) );
  AOI211_X1 U9761 ( .C1(n8349), .C2(n9334), .A(n4269), .B(n8236), .ZN(n8348)
         );
  NOR2_X1 U9762 ( .A1(n4787), .A2(n8237), .ZN(n8242) );
  INV_X1 U9763 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8240) );
  OAI22_X1 U9764 ( .A1(n8265), .A2(n8240), .B1(n8239), .B2(n8238), .ZN(n8241)
         );
  AOI211_X1 U9765 ( .C1(n8348), .C2(n8243), .A(n8242), .B(n8241), .ZN(n8253)
         );
  NAND2_X1 U9766 ( .A1(n9322), .A2(n8244), .ZN(n8246) );
  XNOR2_X1 U9767 ( .A(n8246), .B(n8245), .ZN(n8247) );
  OAI222_X1 U9768 ( .A1(n8251), .A2(n8250), .B1(n8249), .B2(n8248), .C1(n8247), 
        .C2(n9345), .ZN(n8347) );
  NAND2_X1 U9769 ( .A1(n8347), .A2(n8265), .ZN(n8252) );
  OAI211_X1 U9770 ( .C1(n8351), .C2(n8254), .A(n8253), .B(n8252), .ZN(P2_U3279) );
  AOI21_X1 U9771 ( .B1(n9638), .B2(n9644), .A(n8255), .ZN(n9643) );
  AOI22_X1 U9772 ( .A1(n9643), .A2(n9337), .B1(n9591), .B2(n9644), .ZN(n8271)
         );
  INV_X1 U9773 ( .A(n8256), .ZN(n8261) );
  XNOR2_X1 U9774 ( .A(n8257), .B(n9644), .ZN(n8267) );
  NAND2_X1 U9775 ( .A1(n8267), .A2(n8258), .ZN(n8259) );
  OAI211_X1 U9776 ( .C1(n8261), .C2(n8260), .A(n8259), .B(n9619), .ZN(n8263)
         );
  AOI22_X1 U9777 ( .A1(n5924), .A2(n9621), .B1(n9624), .B2(n5567), .ZN(n8262)
         );
  NAND2_X1 U9778 ( .A1(n8263), .A2(n8262), .ZN(n9646) );
  AOI22_X1 U9779 ( .A1(n9646), .A2(n8265), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n9613), .ZN(n8270) );
  OR2_X1 U9780 ( .A1(n8265), .A2(n8264), .ZN(n8269) );
  XOR2_X1 U9781 ( .A(n8266), .B(n8267), .Z(n9648) );
  NAND2_X1 U9782 ( .A1(n9601), .A2(n9648), .ZN(n8268) );
  NAND4_X1 U9783 ( .A1(n8271), .A2(n8270), .A3(n8269), .A4(n8268), .ZN(
        P2_U3295) );
  NAND2_X1 U9784 ( .A1(n8272), .A2(n9694), .ZN(n8273) );
  OAI211_X1 U9785 ( .C1(n8274), .C2(n4269), .A(n8273), .B(n8283), .ZN(n8355)
         );
  NAND4_X1 U9786 ( .A1(n8278), .A2(n8277), .A3(n8276), .A4(n8275), .ZN(n8279)
         );
  OR2_X1 U9787 ( .A1(n8280), .A2(n8279), .ZN(n8354) );
  INV_X2 U9788 ( .A(n9742), .ZN(n9745) );
  MUX2_X1 U9789 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8355), .S(n9745), .Z(
        P2_U3551) );
  NAND3_X1 U9790 ( .A1(n8282), .A2(n9606), .A3(n8281), .ZN(n8284) );
  OAI211_X1 U9791 ( .C1(n8285), .C2(n9719), .A(n8284), .B(n8283), .ZN(n8356)
         );
  MUX2_X1 U9792 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8356), .S(n9745), .Z(
        P2_U3550) );
  MUX2_X1 U9793 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8357), .S(n9745), .Z(
        P2_U3549) );
  AOI22_X1 U9794 ( .A1(n8291), .A2(n9606), .B1(n9694), .B2(n8290), .ZN(n8292)
         );
  OAI211_X1 U9795 ( .C1(n8294), .C2(n9652), .A(n8293), .B(n8292), .ZN(n8358)
         );
  MUX2_X1 U9796 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8358), .S(n9745), .Z(
        P2_U3548) );
  AOI21_X1 U9797 ( .B1(n9694), .B2(n8296), .A(n8295), .ZN(n8297) );
  OAI211_X1 U9798 ( .C1(n8299), .C2(n9652), .A(n8298), .B(n8297), .ZN(n8359)
         );
  MUX2_X1 U9799 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8359), .S(n9745), .Z(
        P2_U3547) );
  AOI21_X1 U9800 ( .B1(n9694), .B2(n8301), .A(n8300), .ZN(n8302) );
  OAI211_X1 U9801 ( .C1(n8304), .C2(n9652), .A(n8303), .B(n8302), .ZN(n8360)
         );
  MUX2_X1 U9802 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8360), .S(n9745), .Z(
        P2_U3546) );
  AOI21_X1 U9803 ( .B1(n9694), .B2(n8306), .A(n8305), .ZN(n8307) );
  OAI211_X1 U9804 ( .C1(n8309), .C2(n9652), .A(n8308), .B(n8307), .ZN(n8361)
         );
  MUX2_X1 U9805 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8361), .S(n9745), .Z(
        P2_U3545) );
  AOI22_X1 U9806 ( .A1(n8311), .A2(n9606), .B1(n9694), .B2(n8310), .ZN(n8312)
         );
  OAI211_X1 U9807 ( .C1(n8314), .C2(n9652), .A(n8313), .B(n8312), .ZN(n8362)
         );
  MUX2_X1 U9808 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8362), .S(n9745), .Z(
        P2_U3544) );
  INV_X1 U9809 ( .A(n9652), .ZN(n9723) );
  NAND3_X1 U9810 ( .A1(n8316), .A2(n8315), .A3(n9723), .ZN(n8321) );
  AOI22_X1 U9811 ( .A1(n8318), .A2(n9606), .B1(n9694), .B2(n8317), .ZN(n8319)
         );
  NAND3_X1 U9812 ( .A1(n8321), .A2(n8320), .A3(n8319), .ZN(n8363) );
  MUX2_X1 U9813 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8363), .S(n9745), .Z(
        P2_U3543) );
  AOI22_X1 U9814 ( .A1(n8323), .A2(n9606), .B1(n9694), .B2(n8322), .ZN(n8324)
         );
  OAI211_X1 U9815 ( .C1(n8326), .C2(n9652), .A(n8325), .B(n8324), .ZN(n8364)
         );
  MUX2_X1 U9816 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8364), .S(n9745), .Z(
        P2_U3542) );
  AOI22_X1 U9817 ( .A1(n8328), .A2(n9606), .B1(n9694), .B2(n8327), .ZN(n8329)
         );
  OAI211_X1 U9818 ( .C1(n8331), .C2(n9652), .A(n8330), .B(n8329), .ZN(n8365)
         );
  MUX2_X1 U9819 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8365), .S(n9745), .Z(
        P2_U3541) );
  AOI22_X1 U9820 ( .A1(n8333), .A2(n9606), .B1(n9694), .B2(n8332), .ZN(n8334)
         );
  OAI211_X1 U9821 ( .C1(n8336), .C2(n9652), .A(n8335), .B(n8334), .ZN(n8366)
         );
  MUX2_X1 U9822 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8366), .S(n9745), .Z(
        P2_U3540) );
  AOI21_X1 U9823 ( .B1(n9694), .B2(n8338), .A(n8337), .ZN(n8339) );
  OAI211_X1 U9824 ( .C1(n8341), .C2(n9652), .A(n8340), .B(n8339), .ZN(n8367)
         );
  MUX2_X1 U9825 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8367), .S(n9745), .Z(
        P2_U3539) );
  AOI22_X1 U9826 ( .A1(n8343), .A2(n9606), .B1(n9694), .B2(n8342), .ZN(n8344)
         );
  OAI211_X1 U9827 ( .C1(n8346), .C2(n9652), .A(n8345), .B(n8344), .ZN(n8368)
         );
  MUX2_X1 U9828 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8368), .S(n9745), .Z(
        P2_U3538) );
  AOI211_X1 U9829 ( .C1(n9694), .C2(n8349), .A(n8348), .B(n8347), .ZN(n8350)
         );
  OAI21_X1 U9830 ( .B1(n8351), .B2(n9652), .A(n8350), .ZN(n8369) );
  MUX2_X1 U9831 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8369), .S(n9745), .Z(
        P2_U3537) );
  INV_X1 U9832 ( .A(n8352), .ZN(n8353) );
  INV_X2 U9833 ( .A(n9724), .ZN(n9726) );
  MUX2_X1 U9834 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8355), .S(n9726), .Z(
        P2_U3519) );
  MUX2_X1 U9835 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8356), .S(n9726), .Z(
        P2_U3518) );
  MUX2_X1 U9836 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8358), .S(n9726), .Z(
        P2_U3516) );
  MUX2_X1 U9837 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8359), .S(n9726), .Z(
        P2_U3515) );
  MUX2_X1 U9838 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8360), .S(n9726), .Z(
        P2_U3514) );
  MUX2_X1 U9839 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8361), .S(n9726), .Z(
        P2_U3513) );
  MUX2_X1 U9840 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8362), .S(n9726), .Z(
        P2_U3512) );
  MUX2_X1 U9841 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8363), .S(n9726), .Z(
        P2_U3511) );
  MUX2_X1 U9842 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8364), .S(n9726), .Z(
        P2_U3510) );
  MUX2_X1 U9843 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8365), .S(n9726), .Z(
        P2_U3509) );
  MUX2_X1 U9844 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8366), .S(n9726), .Z(
        P2_U3508) );
  MUX2_X1 U9845 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8367), .S(n9726), .Z(
        P2_U3507) );
  MUX2_X1 U9846 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8368), .S(n9726), .Z(
        P2_U3505) );
  MUX2_X1 U9847 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8369), .S(n9726), .Z(
        P2_U3502) );
  INV_X1 U9848 ( .A(n8608), .ZN(n9267) );
  NAND3_X1 U9849 ( .A1(n8370), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n8372) );
  OAI22_X1 U9850 ( .A1(n5078), .A2(n8372), .B1(n5501), .B2(n8371), .ZN(n8373)
         );
  INV_X1 U9851 ( .A(n8373), .ZN(n8374) );
  OAI21_X1 U9852 ( .B1(n9267), .B2(n4268), .A(n8374), .ZN(P2_U3327) );
  MUX2_X1 U9853 ( .A(n8375), .B(P2_IR_REG_0__SCAN_IN), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  OAI211_X1 U9854 ( .C1(n8376), .C2(n8378), .A(n8377), .B(n8496), .ZN(n8385)
         );
  AOI22_X1 U9855 ( .A1(n8490), .A2(n8380), .B1(n8517), .B2(n8379), .ZN(n8384)
         );
  OR2_X1 U9856 ( .A1(n8511), .A2(n8381), .ZN(n8382) );
  NAND4_X1 U9857 ( .A1(n8385), .A2(n8384), .A3(n8383), .A4(n8382), .ZN(
        P1_U3211) );
  XNOR2_X1 U9858 ( .A(n8387), .B(n8386), .ZN(n8388) );
  XNOR2_X1 U9859 ( .A(n8389), .B(n8388), .ZN(n8395) );
  NAND2_X1 U9860 ( .A1(n8517), .A2(n8390), .ZN(n8391) );
  NAND2_X1 U9861 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9410) );
  OAI211_X1 U9862 ( .C1(n8511), .C2(n8392), .A(n8391), .B(n9410), .ZN(n8393)
         );
  AOI21_X1 U9863 ( .B1(n9205), .B2(n8490), .A(n8393), .ZN(n8394) );
  OAI21_X1 U9864 ( .B1(n8395), .B2(n8519), .A(n8394), .ZN(P1_U3213) );
  NAND2_X1 U9865 ( .A1(n4605), .A2(n8396), .ZN(n8398) );
  XNOR2_X1 U9866 ( .A(n8398), .B(n8397), .ZN(n8404) );
  INV_X1 U9867 ( .A(n8992), .ZN(n8401) );
  OAI22_X1 U9868 ( .A1(n8399), .A2(n9062), .B1(n8418), .B2(n9060), .ZN(n8999)
         );
  AOI22_X1 U9869 ( .A1(n8999), .A2(n8419), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8400) );
  OAI21_X1 U9870 ( .B1(n8401), .B2(n8485), .A(n8400), .ZN(n8402) );
  AOI21_X1 U9871 ( .B1(n9157), .B2(n8490), .A(n8402), .ZN(n8403) );
  OAI21_X1 U9872 ( .B1(n8404), .B2(n8519), .A(n8403), .ZN(P1_U3214) );
  INV_X1 U9873 ( .A(n8406), .ZN(n8407) );
  AOI21_X1 U9874 ( .B1(n8408), .B2(n8405), .A(n8407), .ZN(n8413) );
  NOR2_X1 U9875 ( .A1(n8409), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8881) );
  OAI22_X1 U9876 ( .A1(n9059), .A2(n8500), .B1(n8487), .B2(n9061), .ZN(n8410)
         );
  AOI211_X1 U9877 ( .C1(n8517), .C2(n9065), .A(n8881), .B(n8410), .ZN(n8412)
         );
  NAND2_X1 U9878 ( .A1(n9179), .A2(n8490), .ZN(n8411) );
  OAI211_X1 U9879 ( .C1(n8413), .C2(n8519), .A(n8412), .B(n8411), .ZN(P1_U3217) );
  NOR2_X1 U9880 ( .A1(n7624), .A2(n8416), .ZN(n8417) );
  XNOR2_X1 U9881 ( .A(n8414), .B(n8417), .ZN(n8423) );
  OAI22_X1 U9882 ( .A1(n8418), .A2(n9062), .B1(n9061), .B2(n9060), .ZN(n9022)
         );
  AOI22_X1 U9883 ( .A1(n9022), .A2(n8419), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8420) );
  OAI21_X1 U9884 ( .B1(n9020), .B2(n8485), .A(n8420), .ZN(n8421) );
  AOI21_X1 U9885 ( .B1(n9168), .B2(n8490), .A(n8421), .ZN(n8422) );
  OAI21_X1 U9886 ( .B1(n8423), .B2(n8519), .A(n8422), .ZN(P1_U3221) );
  AOI21_X1 U9887 ( .B1(n8426), .B2(n8425), .A(n8424), .ZN(n8430) );
  AOI22_X1 U9888 ( .A1(n8896), .A2(n9114), .B1(n9112), .B2(n8807), .ZN(n8965)
         );
  AOI22_X1 U9889 ( .A1(n8517), .A2(n8969), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8427) );
  OAI21_X1 U9890 ( .B1(n8965), .B2(n8511), .A(n8427), .ZN(n8428) );
  AOI21_X1 U9891 ( .B1(n9148), .B2(n8490), .A(n8428), .ZN(n8429) );
  OAI21_X1 U9892 ( .B1(n8430), .B2(n8519), .A(n8429), .ZN(P1_U3223) );
  INV_X1 U9893 ( .A(n9195), .ZN(n9108) );
  INV_X1 U9894 ( .A(n8431), .ZN(n8444) );
  AOI21_X1 U9895 ( .B1(n8432), .B2(n8433), .A(n8434), .ZN(n8435) );
  OAI21_X1 U9896 ( .B1(n8444), .B2(n8435), .A(n8496), .ZN(n8440) );
  OAI22_X1 U9897 ( .A1(n8436), .A2(n8500), .B1(n8487), .B2(n8486), .ZN(n8437)
         );
  AOI211_X1 U9898 ( .C1(n8517), .C2(n9106), .A(n8438), .B(n8437), .ZN(n8439)
         );
  OAI211_X1 U9899 ( .C1(n9108), .C2(n8512), .A(n8440), .B(n8439), .ZN(P1_U3224) );
  INV_X1 U9900 ( .A(n8441), .ZN(n8443) );
  NOR3_X1 U9901 ( .A1(n8444), .A2(n8443), .A3(n8442), .ZN(n8447) );
  INV_X1 U9902 ( .A(n8445), .ZN(n8446) );
  OAI21_X1 U9903 ( .B1(n8447), .B2(n8446), .A(n8496), .ZN(n8451) );
  AND2_X1 U9904 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8849) );
  OAI22_X1 U9905 ( .A1(n8448), .A2(n8500), .B1(n8487), .B2(n9059), .ZN(n8449)
         );
  AOI211_X1 U9906 ( .C1(n8517), .C2(n9089), .A(n8849), .B(n8449), .ZN(n8450)
         );
  OAI211_X1 U9907 ( .C1(n9091), .C2(n8512), .A(n8451), .B(n8450), .ZN(P1_U3226) );
  AOI21_X1 U9908 ( .B1(n8454), .B2(n8453), .A(n8452), .ZN(n8459) );
  OAI22_X1 U9909 ( .A1(n8485), .A2(n8985), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8455), .ZN(n8457) );
  OAI22_X1 U9910 ( .A1(n8501), .A2(n8487), .B1(n8474), .B2(n8500), .ZN(n8456)
         );
  AOI211_X1 U9911 ( .C1(n9152), .C2(n8490), .A(n8457), .B(n8456), .ZN(n8458)
         );
  OAI21_X1 U9912 ( .B1(n8459), .B2(n8519), .A(n8458), .ZN(P1_U3227) );
  INV_X1 U9913 ( .A(n8461), .ZN(n8463) );
  NAND2_X1 U9914 ( .A1(n8463), .A2(n8462), .ZN(n8464) );
  XNOR2_X1 U9915 ( .A(n8460), .B(n8464), .ZN(n8469) );
  OAI22_X1 U9916 ( .A1(n8485), .A2(n8465), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9856), .ZN(n8467) );
  OAI22_X1 U9917 ( .A1(n9040), .A2(n8500), .B1(n8487), .B2(n9041), .ZN(n8466)
         );
  AOI211_X1 U9918 ( .C1(n9174), .C2(n8490), .A(n8467), .B(n8466), .ZN(n8468)
         );
  OAI21_X1 U9919 ( .B1(n8469), .B2(n8519), .A(n8468), .ZN(P1_U3231) );
  XNOR2_X1 U9920 ( .A(n8471), .B(n4284), .ZN(n8472) );
  XNOR2_X1 U9921 ( .A(n8470), .B(n8472), .ZN(n8478) );
  OAI22_X1 U9922 ( .A1(n8485), .A2(n9007), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8473), .ZN(n8476) );
  OAI22_X1 U9923 ( .A1(n8474), .A2(n8487), .B1(n8500), .B2(n9041), .ZN(n8475)
         );
  AOI211_X1 U9924 ( .C1(n9161), .C2(n8490), .A(n8476), .B(n8475), .ZN(n8477)
         );
  OAI21_X1 U9925 ( .B1(n8478), .B2(n8519), .A(n8477), .ZN(P1_U3233) );
  NAND2_X1 U9926 ( .A1(n8480), .A2(n8479), .ZN(n8481) );
  XOR2_X1 U9927 ( .A(n8482), .B(n8481), .Z(n8492) );
  INV_X1 U9928 ( .A(n9080), .ZN(n8484) );
  OAI22_X1 U9929 ( .A1(n8485), .A2(n8484), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8483), .ZN(n8489) );
  OAI22_X1 U9930 ( .A1(n9040), .A2(n8487), .B1(n8500), .B2(n8486), .ZN(n8488)
         );
  AOI211_X1 U9931 ( .C1(n9184), .C2(n8490), .A(n8489), .B(n8488), .ZN(n8491)
         );
  OAI21_X1 U9932 ( .B1(n8492), .B2(n8519), .A(n8491), .ZN(P1_U3236) );
  OAI21_X1 U9933 ( .B1(n8424), .B2(n8494), .A(n8493), .ZN(n8495) );
  NAND3_X1 U9934 ( .A1(n8497), .A2(n8496), .A3(n8495), .ZN(n8505) );
  AOI22_X1 U9935 ( .A1(n8498), .A2(n8517), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n8499) );
  OAI21_X1 U9936 ( .B1(n8501), .B2(n8500), .A(n8499), .ZN(n8502) );
  AOI21_X1 U9937 ( .B1(n8806), .B2(n8503), .A(n8502), .ZN(n8504) );
  OAI211_X1 U9938 ( .C1(n8897), .C2(n8512), .A(n8505), .B(n8504), .ZN(P1_U3238) );
  NAND2_X1 U9939 ( .A1(n8433), .A2(n8506), .ZN(n8507) );
  XOR2_X1 U9940 ( .A(n8508), .B(n8507), .Z(n8520) );
  OAI22_X1 U9941 ( .A1(n8511), .A2(n8510), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8509), .ZN(n8515) );
  NOR2_X1 U9942 ( .A1(n8513), .A2(n8512), .ZN(n8514) );
  AOI211_X1 U9943 ( .C1(n8517), .C2(n8516), .A(n8515), .B(n8514), .ZN(n8518)
         );
  OAI21_X1 U9944 ( .B1(n8520), .B2(n8519), .A(n8518), .ZN(P1_U3239) );
  NAND2_X1 U9945 ( .A1(n8521), .A2(n7642), .ZN(n8523) );
  NAND2_X1 U9946 ( .A1(n8612), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8522) );
  INV_X1 U9947 ( .A(n9128), .ZN(n8626) );
  INV_X1 U9948 ( .A(n8908), .ZN(n8926) );
  OAI21_X1 U9949 ( .B1(n8926), .B2(n8628), .A(n8728), .ZN(n8524) );
  OAI21_X1 U9950 ( .B1(n8728), .B2(n8628), .A(n8524), .ZN(n8527) );
  NOR2_X1 U9951 ( .A1(n8909), .A2(n8628), .ZN(n8593) );
  INV_X1 U9952 ( .A(n8593), .ZN(n8526) );
  NAND2_X1 U9953 ( .A1(n9136), .A2(n8899), .ZN(n8632) );
  NAND3_X1 U9954 ( .A1(n8909), .A2(n8628), .A3(n8632), .ZN(n8525) );
  NAND3_X1 U9955 ( .A1(n8527), .A2(n8526), .A3(n8525), .ZN(n8606) );
  INV_X1 U9956 ( .A(n8731), .ZN(n8571) );
  AND2_X1 U9957 ( .A1(n8547), .A2(n8628), .ZN(n8548) );
  INV_X1 U9958 ( .A(n9230), .ZN(n8528) );
  NAND2_X1 U9959 ( .A1(n8528), .A2(n8674), .ZN(n8534) );
  NAND3_X1 U9960 ( .A1(n8530), .A2(n8666), .A3(n8529), .ZN(n8532) );
  NAND3_X1 U9961 ( .A1(n8532), .A2(n8531), .A3(n8667), .ZN(n8533) );
  MUX2_X1 U9962 ( .A(n8671), .B(n8674), .S(n8628), .Z(n8535) );
  AND2_X1 U9963 ( .A1(n8539), .A2(n8536), .ZN(n8643) );
  NAND2_X1 U9964 ( .A1(n8540), .A2(n8643), .ZN(n8538) );
  NAND2_X1 U9965 ( .A1(n8641), .A2(n4267), .ZN(n8545) );
  AOI21_X1 U9966 ( .B1(n8538), .B2(n8537), .A(n8545), .ZN(n8544) );
  INV_X1 U9967 ( .A(n8539), .ZN(n8677) );
  INV_X1 U9968 ( .A(n8541), .ZN(n8753) );
  INV_X1 U9969 ( .A(n8679), .ZN(n8646) );
  OAI22_X1 U9970 ( .A1(n8542), .A2(n8753), .B1(n8646), .B2(n8628), .ZN(n8543)
         );
  OAI21_X1 U9971 ( .B1(n8548), .B2(n8544), .A(n8543), .ZN(n8555) );
  INV_X1 U9972 ( .A(n8545), .ZN(n8551) );
  NAND2_X1 U9973 ( .A1(n8547), .A2(n8546), .ZN(n8682) );
  INV_X1 U9974 ( .A(n8548), .ZN(n8549) );
  AOI21_X1 U9975 ( .B1(n8679), .B2(n8641), .A(n8549), .ZN(n8550) );
  AOI211_X1 U9976 ( .C1(n8551), .C2(n8682), .A(n8755), .B(n8550), .ZN(n8554)
         );
  INV_X1 U9977 ( .A(n8642), .ZN(n8552) );
  MUX2_X1 U9978 ( .A(n8552), .B(n8683), .S(n8628), .Z(n8553) );
  AOI211_X1 U9979 ( .C1(n8555), .C2(n8554), .A(n8553), .B(n9102), .ZN(n8559)
         );
  INV_X1 U9980 ( .A(n8684), .ZN(n8557) );
  MUX2_X1 U9981 ( .A(n8557), .B(n8556), .S(n8628), .Z(n8558) );
  NOR3_X1 U9982 ( .A1(n8559), .A2(n8558), .A3(n8732), .ZN(n8563) );
  NAND2_X1 U9983 ( .A1(n8640), .A2(n8638), .ZN(n8561) );
  NAND2_X1 U9984 ( .A1(n9054), .A2(n8560), .ZN(n8691) );
  MUX2_X1 U9985 ( .A(n8561), .B(n8691), .S(n8628), .Z(n8562) );
  NOR2_X1 U9986 ( .A1(n8563), .A2(n8562), .ZN(n8566) );
  NAND2_X1 U9987 ( .A1(n8565), .A2(n9054), .ZN(n8564) );
  OAI211_X1 U9988 ( .C1(n8566), .C2(n8564), .A(n9036), .B(n8577), .ZN(n8568)
         );
  NAND2_X1 U9989 ( .A1(n9036), .A2(n8640), .ZN(n8694) );
  AND2_X1 U9990 ( .A1(n8569), .A2(n8565), .ZN(n8692) );
  OAI21_X1 U9991 ( .B1(n8566), .B2(n8694), .A(n8692), .ZN(n8567) );
  INV_X1 U9992 ( .A(n8699), .ZN(n8570) );
  INV_X1 U9993 ( .A(n8978), .ZN(n8574) );
  INV_X1 U9994 ( .A(n8704), .ZN(n8573) );
  NAND2_X1 U9995 ( .A1(n8572), .A2(n8729), .ZN(n8708) );
  OAI21_X1 U9996 ( .B1(n8573), .B2(n8776), .A(n8708), .ZN(n8775) );
  OAI21_X1 U9997 ( .B1(n8575), .B2(n8574), .A(n8775), .ZN(n8588) );
  INV_X1 U9998 ( .A(n8962), .ZN(n8586) );
  INV_X1 U9999 ( .A(n8576), .ZN(n8582) );
  INV_X1 U10000 ( .A(n8577), .ZN(n8578) );
  NAND2_X1 U10001 ( .A1(n8693), .A2(n8578), .ZN(n8580) );
  AND2_X1 U10002 ( .A1(n8580), .A2(n8579), .ZN(n8581) );
  NAND2_X1 U10003 ( .A1(n8581), .A2(n8731), .ZN(n8690) );
  AOI21_X1 U10004 ( .B1(n8582), .B2(n8693), .A(n8690), .ZN(n8584) );
  INV_X1 U10005 ( .A(n8995), .ZN(n8583) );
  OAI211_X1 U10006 ( .C1(n8584), .C2(n8583), .A(n8978), .B(n8729), .ZN(n8585)
         );
  AND2_X1 U10007 ( .A1(n8781), .A2(n8776), .ZN(n8703) );
  OAI211_X1 U10008 ( .C1(n8586), .C2(n8730), .A(n8585), .B(n8703), .ZN(n8587)
         );
  MUX2_X1 U10009 ( .A(n8588), .B(n8587), .S(n8628), .Z(n8597) );
  INV_X1 U10010 ( .A(n8597), .ZN(n8596) );
  NAND2_X1 U10011 ( .A1(n9141), .A2(n8781), .ZN(n8590) );
  NAND2_X1 U10012 ( .A1(n8704), .A2(n8896), .ZN(n8589) );
  MUX2_X1 U10013 ( .A(n8590), .B(n8589), .S(n8628), .Z(n8595) );
  NOR2_X1 U10014 ( .A1(n9141), .A2(n4267), .ZN(n8600) );
  INV_X1 U10015 ( .A(n8600), .ZN(n8591) );
  OAI211_X1 U10016 ( .C1(n8952), .C2(n8591), .A(n8728), .B(n8942), .ZN(n8592)
         );
  NOR2_X1 U10017 ( .A1(n8593), .A2(n8592), .ZN(n8594) );
  OAI21_X1 U10018 ( .B1(n8596), .B2(n8595), .A(n8594), .ZN(n8605) );
  OAI21_X1 U10019 ( .B1(n4267), .B2(n8704), .A(n8597), .ZN(n8603) );
  INV_X1 U10020 ( .A(n8728), .ZN(n8599) );
  OAI211_X1 U10021 ( .C1(n9141), .C2(n8781), .A(n8952), .B(n4267), .ZN(n8598)
         );
  OR3_X1 U10022 ( .A1(n8599), .A2(n8926), .A3(n8598), .ZN(n8602) );
  NAND3_X1 U10023 ( .A1(n8909), .A2(n8600), .A3(n8632), .ZN(n8601) );
  AOI22_X1 U10024 ( .A1(n8603), .A2(n8897), .B1(n8602), .B2(n8601), .ZN(n8604)
         );
  AOI21_X1 U10025 ( .B1(n8606), .B2(n8605), .A(n8604), .ZN(n8621) );
  NOR3_X1 U10026 ( .A1(n8621), .A2(n9128), .A3(n8804), .ZN(n8607) );
  NAND2_X1 U10027 ( .A1(n8608), .A2(n7642), .ZN(n8610) );
  NAND2_X1 U10028 ( .A1(n8612), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8609) );
  NAND2_X1 U10029 ( .A1(n9122), .A2(n8887), .ZN(n8623) );
  NAND2_X1 U10030 ( .A1(n8611), .A2(n7642), .ZN(n8614) );
  NAND2_X1 U10031 ( .A1(n8612), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8613) );
  NAND2_X1 U10032 ( .A1(n8615), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8618) );
  NAND2_X1 U10033 ( .A1(n7591), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8617) );
  NAND2_X1 U10034 ( .A1(n5785), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8616) );
  AND3_X1 U10035 ( .A1(n8618), .A2(n8617), .A3(n8616), .ZN(n8913) );
  OR2_X1 U10036 ( .A1(n9396), .A2(n8913), .ZN(n8619) );
  INV_X1 U10037 ( .A(n8913), .ZN(n8803) );
  AOI21_X1 U10038 ( .B1(n8803), .B2(n8620), .A(n8892), .ZN(n8624) );
  NOR2_X1 U10039 ( .A1(n8622), .A2(n8624), .ZN(n8629) );
  NAND2_X1 U10040 ( .A1(n8621), .A2(n8629), .ZN(n8627) );
  INV_X1 U10041 ( .A(n8804), .ZN(n8634) );
  INV_X1 U10042 ( .A(n8622), .ZN(n8790) );
  INV_X1 U10043 ( .A(n8623), .ZN(n8625) );
  INV_X1 U10044 ( .A(n8624), .ZN(n8786) );
  NAND2_X1 U10045 ( .A1(n8772), .A2(n8917), .ZN(n8715) );
  INV_X1 U10046 ( .A(n8767), .ZN(n8712) );
  NAND2_X1 U10047 ( .A1(n9396), .A2(n8913), .ZN(n8765) );
  OR2_X1 U10048 ( .A1(n9128), .A2(n8634), .ZN(n8630) );
  NAND2_X1 U10049 ( .A1(n8630), .A2(n8728), .ZN(n8788) );
  NAND2_X1 U10050 ( .A1(n8908), .A2(n8905), .ZN(n8631) );
  AND3_X1 U10051 ( .A1(n8909), .A2(n8632), .A3(n8631), .ZN(n8633) );
  OR2_X1 U10052 ( .A1(n8788), .A2(n8633), .ZN(n8636) );
  NAND2_X1 U10053 ( .A1(n9128), .A2(n8634), .ZN(n8635) );
  AND2_X1 U10054 ( .A1(n8636), .A2(n8635), .ZN(n8785) );
  INV_X1 U10055 ( .A(n8942), .ZN(n8951) );
  OR2_X1 U10056 ( .A1(n8690), .A2(n8637), .ZN(n8701) );
  AND2_X1 U10057 ( .A1(n8638), .A2(n9092), .ZN(n8639) );
  AND2_X1 U10058 ( .A1(n8640), .A2(n8639), .ZN(n8689) );
  INV_X1 U10059 ( .A(n8689), .ZN(n8648) );
  NAND2_X1 U10060 ( .A1(n8642), .A2(n8641), .ZN(n8686) );
  INV_X1 U10061 ( .A(n8643), .ZN(n8676) );
  NAND3_X1 U10062 ( .A1(n8644), .A2(n8674), .A3(n8667), .ZN(n8645) );
  OR4_X1 U10063 ( .A1(n8686), .A2(n8646), .A3(n8676), .A4(n8645), .ZN(n8647)
         );
  OR2_X1 U10064 ( .A1(n8648), .A2(n8647), .ZN(n8649) );
  NOR2_X1 U10065 ( .A1(n8701), .A2(n8649), .ZN(n8780) );
  NAND2_X1 U10066 ( .A1(n5875), .A2(n8650), .ZN(n8651) );
  NAND3_X1 U10067 ( .A1(n8652), .A2(n8794), .A3(n8651), .ZN(n8653) );
  NAND2_X1 U10068 ( .A1(n8654), .A2(n8653), .ZN(n8656) );
  OAI21_X1 U10069 ( .B1(n8657), .B2(n8656), .A(n8655), .ZN(n8659) );
  NAND2_X1 U10070 ( .A1(n8659), .A2(n8658), .ZN(n8665) );
  AOI21_X1 U10071 ( .B1(n8662), .B2(n8661), .A(n8660), .ZN(n8663) );
  AOI21_X1 U10072 ( .B1(n8665), .B2(n8664), .A(n8663), .ZN(n8702) );
  INV_X1 U10073 ( .A(n8666), .ZN(n8668) );
  NAND2_X1 U10074 ( .A1(n8668), .A2(n8667), .ZN(n8670) );
  NAND2_X1 U10075 ( .A1(n8670), .A2(n8669), .ZN(n8673) );
  INV_X1 U10076 ( .A(n8671), .ZN(n8672) );
  AOI21_X1 U10077 ( .B1(n8674), .B2(n8673), .A(n8672), .ZN(n8675) );
  OAI22_X1 U10078 ( .A1(n8678), .A2(n8677), .B1(n8676), .B2(n8675), .ZN(n8680)
         );
  AND2_X1 U10079 ( .A1(n8680), .A2(n8679), .ZN(n8681) );
  NOR2_X1 U10080 ( .A1(n8682), .A2(n8681), .ZN(n8687) );
  INV_X1 U10081 ( .A(n8683), .ZN(n8685) );
  OAI211_X1 U10082 ( .C1(n8687), .C2(n8686), .A(n8685), .B(n8684), .ZN(n8688)
         );
  NAND2_X1 U10083 ( .A1(n8689), .A2(n8688), .ZN(n8700) );
  INV_X1 U10084 ( .A(n8690), .ZN(n8697) );
  INV_X1 U10085 ( .A(n8691), .ZN(n8695) );
  OAI211_X1 U10086 ( .C1(n8695), .C2(n8694), .A(n8693), .B(n8692), .ZN(n8696)
         );
  NAND2_X1 U10087 ( .A1(n8697), .A2(n8696), .ZN(n8698) );
  OAI211_X1 U10088 ( .C1(n8701), .C2(n8700), .A(n8699), .B(n8698), .ZN(n8777)
         );
  AOI21_X1 U10089 ( .B1(n8780), .B2(n8702), .A(n8777), .ZN(n8707) );
  INV_X1 U10090 ( .A(n8703), .ZN(n8705) );
  NAND2_X1 U10091 ( .A1(n8705), .A2(n8704), .ZN(n8706) );
  OAI211_X1 U10092 ( .C1(n8708), .C2(n8707), .A(n8782), .B(n8706), .ZN(n8709)
         );
  OR3_X1 U10093 ( .A1(n8788), .A2(n8951), .A3(n8709), .ZN(n8710) );
  AND3_X1 U10094 ( .A1(n8765), .A2(n8785), .A3(n8710), .ZN(n8711) );
  NAND2_X1 U10095 ( .A1(n8713), .A2(n8791), .ZN(n8714) );
  MUX2_X1 U10096 ( .A(n8716), .B(n8715), .S(n8714), .Z(n8797) );
  NOR4_X1 U10097 ( .A1(n8717), .A2(n5449), .A3(n8773), .A4(n8770), .ZN(n8718)
         );
  NAND3_X1 U10098 ( .A1(n8719), .A2(n8797), .A3(n8718), .ZN(n8802) );
  NOR3_X1 U10099 ( .A1(n8720), .A2(n9026), .A3(n8770), .ZN(n8721) );
  NAND3_X1 U10100 ( .A1(n8722), .A2(n8797), .A3(n8721), .ZN(n8801) );
  NAND4_X1 U10101 ( .A1(n8725), .A2(n8724), .A3(n8885), .A4(n8723), .ZN(n8726)
         );
  OAI211_X1 U10102 ( .C1(n5449), .C2(n8770), .A(n8726), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8800) );
  NAND2_X1 U10103 ( .A1(n8727), .A2(n8917), .ZN(n8768) );
  INV_X1 U10104 ( .A(n8768), .ZN(n8771) );
  XNOR2_X1 U10105 ( .A(n9128), .B(n8804), .ZN(n8903) );
  INV_X1 U10106 ( .A(n8903), .ZN(n8911) );
  INV_X1 U10107 ( .A(n8922), .ZN(n8927) );
  INV_X1 U10108 ( .A(n8963), .ZN(n8762) );
  NAND2_X1 U10109 ( .A1(n8730), .A2(n8729), .ZN(n8997) );
  AND2_X1 U10110 ( .A1(n8995), .A2(n8731), .ZN(n9012) );
  INV_X1 U10111 ( .A(n9051), .ZN(n9053) );
  INV_X1 U10112 ( .A(n8732), .ZN(n9093) );
  NAND3_X1 U10113 ( .A1(n8735), .A2(n8734), .A3(n8733), .ZN(n8740) );
  NAND3_X1 U10114 ( .A1(n8738), .A2(n8737), .A3(n8736), .ZN(n8739) );
  NOR2_X1 U10115 ( .A1(n8740), .A2(n8739), .ZN(n8744) );
  NAND4_X1 U10116 ( .A1(n8744), .A2(n8743), .A3(n8742), .A4(n8741), .ZN(n8746)
         );
  NOR2_X1 U10117 ( .A1(n8746), .A2(n8745), .ZN(n8750) );
  NAND4_X1 U10118 ( .A1(n8750), .A2(n8749), .A3(n8748), .A4(n8747), .ZN(n8751)
         );
  OR3_X1 U10119 ( .A1(n8753), .A2(n8752), .A3(n8751), .ZN(n8754) );
  NOR3_X1 U10120 ( .A1(n9102), .A2(n8755), .A3(n8754), .ZN(n8756) );
  NAND4_X1 U10121 ( .A1(n9053), .A2(n4491), .A3(n9093), .A4(n8756), .ZN(n8757)
         );
  NOR2_X1 U10122 ( .A1(n9037), .A2(n8757), .ZN(n8758) );
  NAND3_X1 U10123 ( .A1(n9012), .A2(n8759), .A3(n8758), .ZN(n8760) );
  NOR2_X1 U10124 ( .A1(n8997), .A2(n8760), .ZN(n8761) );
  NAND4_X1 U10125 ( .A1(n8763), .A2(n8762), .A3(n8978), .A4(n8761), .ZN(n8764)
         );
  NOR4_X1 U10126 ( .A1(n8911), .A2(n8927), .A3(n8951), .A4(n8764), .ZN(n8766)
         );
  NAND4_X1 U10127 ( .A1(n8767), .A2(n8766), .A3(n8765), .A4(n8791), .ZN(n8774)
         );
  NOR2_X1 U10128 ( .A1(n8774), .A2(n8768), .ZN(n8769) );
  AOI211_X1 U10129 ( .C1(n8794), .C2(n8771), .A(n8770), .B(n8769), .ZN(n8798)
         );
  NOR2_X1 U10130 ( .A1(n8772), .A2(n8917), .ZN(n8792) );
  NAND3_X1 U10131 ( .A1(n8774), .A2(n8792), .A3(n8773), .ZN(n8796) );
  INV_X1 U10132 ( .A(n8775), .ZN(n8784) );
  INV_X1 U10133 ( .A(n8776), .ZN(n8778) );
  AOI211_X1 U10134 ( .C1(n8780), .C2(n8779), .A(n8778), .B(n8777), .ZN(n8783)
         );
  OAI211_X1 U10135 ( .C1(n8784), .C2(n8783), .A(n8906), .B(n8908), .ZN(n8787)
         );
  OAI211_X1 U10136 ( .C1(n8788), .C2(n8787), .A(n8786), .B(n8785), .ZN(n8789)
         );
  NAND2_X1 U10137 ( .A1(n8790), .A2(n8789), .ZN(n8793) );
  NAND4_X1 U10138 ( .A1(n8794), .A2(n8793), .A3(n8792), .A4(n8791), .ZN(n8795)
         );
  NAND4_X1 U10139 ( .A1(n8798), .A2(n8797), .A3(n8796), .A4(n8795), .ZN(n8799)
         );
  NAND4_X1 U10140 ( .A1(n8802), .A2(n8801), .A3(n8800), .A4(n8799), .ZN(
        P1_U3240) );
  MUX2_X1 U10141 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n8803), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10142 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n8804), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10143 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n8805), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10144 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n8806), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10145 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n8896), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10146 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n8979), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10147 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n8807), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10148 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9013), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10149 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n8808), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10150 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9014), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10151 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n8809), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10152 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9073), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10153 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9096), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10154 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9115), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10155 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9095), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10156 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9113), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10157 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n8810), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10158 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n8811), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10159 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n8812), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10160 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n8813), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10161 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n8814), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10162 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n8815), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10163 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n8816), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10164 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n8817), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10165 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n8818), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10166 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n8819), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10167 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n8820), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10168 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n8821), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10169 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n8822), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10170 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n5875), .S(P1_U4006), .Z(
        P1_U3556) );
  MUX2_X1 U10171 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n8823), .S(P1_U4006), .Z(
        P1_U3555) );
  OAI21_X1 U10172 ( .B1(n8826), .B2(n8825), .A(n8824), .ZN(n8827) );
  NAND2_X1 U10173 ( .A1(n8827), .A2(n9422), .ZN(n8836) );
  AOI22_X1 U10174 ( .A1(n9413), .A2(n8828), .B1(P1_REG3_REG_11__SCAN_IN), .B2(
        P1_U3084), .ZN(n8835) );
  OAI21_X1 U10175 ( .B1(n8831), .B2(n8830), .A(n8829), .ZN(n8832) );
  NAND2_X1 U10176 ( .A1(n8832), .A2(n9421), .ZN(n8834) );
  NAND2_X1 U10177 ( .A1(n8864), .A2(P1_ADDR_REG_11__SCAN_IN), .ZN(n8833) );
  NAND4_X1 U10178 ( .A1(n8836), .A2(n8835), .A3(n8834), .A4(n8833), .ZN(
        P1_U3252) );
  INV_X1 U10179 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n8852) );
  AOI21_X1 U10180 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(n8844), .A(n8837), .ZN(
        n8841) );
  INV_X1 U10181 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n8838) );
  AOI22_X1 U10182 ( .A1(P1_REG1_REG_17__SCAN_IN), .A2(n8839), .B1(n8859), .B2(
        n8838), .ZN(n8840) );
  AOI211_X1 U10183 ( .C1(n8841), .C2(n8840), .A(n8853), .B(n8855), .ZN(n8842)
         );
  INV_X1 U10184 ( .A(n8842), .ZN(n8851) );
  NAND2_X1 U10185 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n8859), .ZN(n8845) );
  OAI21_X1 U10186 ( .B1(n8859), .B2(P1_REG2_REG_17__SCAN_IN), .A(n8845), .ZN(
        n8846) );
  AOI211_X1 U10187 ( .C1(n8847), .C2(n8846), .A(n8858), .B(n8861), .ZN(n8848)
         );
  AOI211_X1 U10188 ( .C1(n8859), .C2(n9413), .A(n8849), .B(n8848), .ZN(n8850)
         );
  OAI211_X1 U10189 ( .C1(n9426), .C2(n8852), .A(n8851), .B(n8850), .ZN(
        P1_U3258) );
  INV_X1 U10190 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n8854) );
  AOI22_X1 U10191 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n8874), .B1(n8867), .B2(
        n8854), .ZN(n8856) );
  AOI221_X1 U10192 ( .B1(n8857), .B2(n8873), .C1(n8856), .C2(n8873), .A(n8855), 
        .ZN(n8870) );
  AOI21_X1 U10193 ( .B1(n8859), .B2(P1_REG2_REG_17__SCAN_IN), .A(n8858), .ZN(
        n8863) );
  NAND2_X1 U10194 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n8874), .ZN(n8860) );
  OAI21_X1 U10195 ( .B1(n8874), .B2(P1_REG2_REG_18__SCAN_IN), .A(n8860), .ZN(
        n8862) );
  NOR2_X1 U10196 ( .A1(n8863), .A2(n8862), .ZN(n8871) );
  AOI211_X1 U10197 ( .C1(n8863), .C2(n8862), .A(n8871), .B(n8861), .ZN(n8869)
         );
  NAND2_X1 U10198 ( .A1(n8864), .A2(P1_ADDR_REG_18__SCAN_IN), .ZN(n8866) );
  NAND2_X1 U10199 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3084), .ZN(n8865) );
  OAI211_X1 U10200 ( .C1(n4363), .C2(n8867), .A(n8866), .B(n8865), .ZN(n8868)
         );
  OR3_X1 U10201 ( .A1(n8870), .A2(n8869), .A3(n8868), .ZN(P1_U3259) );
  INV_X1 U10202 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n8883) );
  AOI21_X1 U10203 ( .B1(n8874), .B2(P1_REG2_REG_18__SCAN_IN), .A(n8871), .ZN(
        n8872) );
  XNOR2_X1 U10204 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n8872), .ZN(n8879) );
  INV_X1 U10205 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n8875) );
  XOR2_X1 U10206 ( .A(n8876), .B(n8875), .Z(n8877) );
  AOI22_X1 U10207 ( .A1(n8879), .A2(n9422), .B1(n9421), .B2(n8877), .ZN(n8880)
         );
  INV_X1 U10208 ( .A(n8881), .ZN(n8882) );
  NAND2_X1 U10209 ( .A1(n8915), .A2(n8892), .ZN(n8884) );
  XNOR2_X1 U10210 ( .A(n8884), .B(n9122), .ZN(n9124) );
  NAND2_X1 U10211 ( .A1(n8885), .A2(P1_B_REG_SCAN_IN), .ZN(n8886) );
  NAND2_X1 U10212 ( .A1(n9114), .A2(n8886), .ZN(n8914) );
  NOR2_X1 U10213 ( .A1(n8887), .A2(n8914), .ZN(n9395) );
  INV_X1 U10214 ( .A(n9395), .ZN(n8888) );
  NOR2_X1 U10215 ( .A1(n9030), .A2(n8888), .ZN(n8894) );
  NOR2_X1 U10216 ( .A1(n8889), .A2(n9428), .ZN(n8890) );
  AOI211_X1 U10217 ( .C1(n9433), .C2(P1_REG2_REG_31__SCAN_IN), .A(n8894), .B(
        n8890), .ZN(n8891) );
  OAI21_X1 U10218 ( .B1(n9124), .B2(n9429), .A(n8891), .ZN(P1_U3261) );
  NOR2_X1 U10219 ( .A1(n8892), .A2(n9428), .ZN(n8893) );
  AOI211_X1 U10220 ( .C1(n9433), .C2(P1_REG2_REG_30__SCAN_IN), .A(n8894), .B(
        n8893), .ZN(n8895) );
  OAI21_X1 U10221 ( .B1(n9429), .B2(n9393), .A(n8895), .ZN(P1_U3262) );
  OR2_X1 U10222 ( .A1(n8941), .A2(n8942), .ZN(n8901) );
  NAND2_X1 U10223 ( .A1(n8949), .A2(n8899), .ZN(n8900) );
  INV_X1 U10224 ( .A(n9131), .ZN(n8936) );
  XNOR2_X1 U10225 ( .A(n8904), .B(n8903), .ZN(n9125) );
  INV_X1 U10226 ( .A(n9125), .ZN(n8921) );
  AOI22_X1 U10227 ( .A1(n9128), .A2(n9031), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9030), .ZN(n8920) );
  NAND2_X1 U10228 ( .A1(n8922), .A2(n8908), .ZN(n8910) );
  OAI21_X1 U10229 ( .B1(n8950), .B2(n8910), .A(n8909), .ZN(n8912) );
  OAI22_X1 U10230 ( .A1(n4417), .A2(n8917), .B1(n9436), .B2(n8916), .ZN(n8918)
         );
  OAI21_X1 U10231 ( .B1(n9126), .B2(n8918), .A(n9070), .ZN(n8919) );
  OAI211_X1 U10232 ( .C1(n8921), .C2(n9121), .A(n8920), .B(n8919), .ZN(
        P1_U3355) );
  NAND2_X1 U10233 ( .A1(n8923), .A2(n8922), .ZN(n8924) );
  INV_X1 U10234 ( .A(n9130), .ZN(n8940) );
  XNOR2_X1 U10235 ( .A(n8928), .B(n8927), .ZN(n8930) );
  INV_X1 U10236 ( .A(n9134), .ZN(n8938) );
  NAND2_X1 U10237 ( .A1(n8944), .A2(n9131), .ZN(n8931) );
  NAND2_X1 U10238 ( .A1(n9132), .A2(n9100), .ZN(n8935) );
  AOI22_X1 U10239 ( .A1(n8933), .A2(n9309), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9030), .ZN(n8934) );
  OAI211_X1 U10240 ( .C1(n8936), .C2(n9428), .A(n8935), .B(n8934), .ZN(n8937)
         );
  AOI21_X1 U10241 ( .B1(n8938), .B2(n9070), .A(n8937), .ZN(n8939) );
  OAI21_X1 U10242 ( .B1(n8940), .B2(n9121), .A(n8939), .ZN(P1_U3263) );
  XOR2_X1 U10243 ( .A(n8942), .B(n8941), .Z(n9140) );
  INV_X1 U10244 ( .A(n8943), .ZN(n8946) );
  INV_X1 U10245 ( .A(n8944), .ZN(n8945) );
  AOI21_X1 U10246 ( .B1(n9136), .B2(n8946), .A(n8945), .ZN(n9137) );
  AOI22_X1 U10247 ( .A1(n8947), .A2(n9309), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9030), .ZN(n8948) );
  OAI21_X1 U10248 ( .B1(n8949), .B2(n9428), .A(n8948), .ZN(n8957) );
  AOI211_X1 U10249 ( .C1(n8951), .C2(n4300), .A(n9229), .B(n8950), .ZN(n8955)
         );
  OAI22_X1 U10250 ( .A1(n8953), .A2(n9062), .B1(n8952), .B2(n9060), .ZN(n8954)
         );
  NOR2_X1 U10251 ( .A1(n8955), .A2(n8954), .ZN(n9139) );
  NOR2_X1 U10252 ( .A1(n9139), .A2(n9321), .ZN(n8956) );
  AOI211_X1 U10253 ( .C1(n9137), .C2(n9100), .A(n8957), .B(n8956), .ZN(n8958)
         );
  OAI21_X1 U10254 ( .B1(n9140), .B2(n9121), .A(n8958), .ZN(P1_U3264) );
  NAND2_X1 U10255 ( .A1(n8959), .A2(n8960), .ZN(n8961) );
  XOR2_X1 U10256 ( .A(n8963), .B(n8961), .Z(n9150) );
  NAND2_X1 U10257 ( .A1(n8976), .A2(n8962), .ZN(n8964) );
  XNOR2_X1 U10258 ( .A(n8964), .B(n8963), .ZN(n8966) );
  OAI21_X1 U10259 ( .B1(n8966), .B2(n9229), .A(n8965), .ZN(n9146) );
  INV_X1 U10260 ( .A(n8967), .ZN(n8968) );
  AOI211_X1 U10261 ( .C1(n9148), .C2(n8981), .A(n9519), .B(n8968), .ZN(n9147)
         );
  NAND2_X1 U10262 ( .A1(n9147), .A2(n9064), .ZN(n8971) );
  AOI22_X1 U10263 ( .A1(n8969), .A2(n9309), .B1(n9433), .B2(
        P1_REG2_REG_25__SCAN_IN), .ZN(n8970) );
  OAI211_X1 U10264 ( .C1(n8972), .C2(n9428), .A(n8971), .B(n8970), .ZN(n8973)
         );
  AOI21_X1 U10265 ( .B1(n9070), .B2(n9146), .A(n8973), .ZN(n8974) );
  OAI21_X1 U10266 ( .B1(n9150), .B2(n9121), .A(n8974), .ZN(P1_U3266) );
  XNOR2_X1 U10267 ( .A(n8975), .B(n8978), .ZN(n9155) );
  AOI22_X1 U10268 ( .A1(n9152), .A2(n9031), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9030), .ZN(n8988) );
  OAI21_X1 U10269 ( .B1(n8978), .B2(n8977), .A(n8976), .ZN(n8980) );
  AOI222_X1 U10270 ( .A1(n9117), .A2(n8980), .B1(n8979), .B2(n9114), .C1(n9013), .C2(n9112), .ZN(n9154) );
  INV_X1 U10271 ( .A(n8990), .ZN(n8983) );
  INV_X1 U10272 ( .A(n8981), .ZN(n8982) );
  AOI211_X1 U10273 ( .C1(n9152), .C2(n8983), .A(n9519), .B(n8982), .ZN(n9151)
         );
  NAND2_X1 U10274 ( .A1(n9151), .A2(n9026), .ZN(n8984) );
  OAI211_X1 U10275 ( .C1(n9436), .C2(n8985), .A(n9154), .B(n8984), .ZN(n8986)
         );
  NAND2_X1 U10276 ( .A1(n8986), .A2(n9070), .ZN(n8987) );
  OAI211_X1 U10277 ( .C1(n9155), .C2(n9121), .A(n8988), .B(n8987), .ZN(
        P1_U3267) );
  XNOR2_X1 U10278 ( .A(n8989), .B(n8997), .ZN(n9160) );
  INV_X1 U10279 ( .A(n9005), .ZN(n8991) );
  AOI211_X1 U10280 ( .C1(n9157), .C2(n8991), .A(n9519), .B(n8990), .ZN(n9156)
         );
  AOI22_X1 U10281 ( .A1(n9433), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n8992), .B2(
        n9309), .ZN(n8993) );
  OAI21_X1 U10282 ( .B1(n8994), .B2(n9428), .A(n8993), .ZN(n9002) );
  NAND2_X1 U10283 ( .A1(n8996), .A2(n8995), .ZN(n8998) );
  XNOR2_X1 U10284 ( .A(n8998), .B(n8997), .ZN(n9000) );
  AOI21_X1 U10285 ( .B1(n9000), .B2(n9117), .A(n8999), .ZN(n9159) );
  NOR2_X1 U10286 ( .A1(n9159), .A2(n9321), .ZN(n9001) );
  AOI211_X1 U10287 ( .C1(n9156), .C2(n9064), .A(n9002), .B(n9001), .ZN(n9003)
         );
  OAI21_X1 U10288 ( .B1(n9160), .B2(n9121), .A(n9003), .ZN(P1_U3268) );
  XOR2_X1 U10289 ( .A(n9012), .B(n9004), .Z(n9165) );
  INV_X1 U10290 ( .A(n9019), .ZN(n9006) );
  AOI21_X1 U10291 ( .B1(n9161), .B2(n9006), .A(n9005), .ZN(n9162) );
  INV_X1 U10292 ( .A(n9007), .ZN(n9008) );
  AOI22_X1 U10293 ( .A1(n9030), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9008), .B2(
        n9309), .ZN(n9009) );
  OAI21_X1 U10294 ( .B1(n9010), .B2(n9428), .A(n9009), .ZN(n9017) );
  XOR2_X1 U10295 ( .A(n9012), .B(n9011), .Z(n9015) );
  AOI222_X1 U10296 ( .A1(n9117), .A2(n9015), .B1(n9014), .B2(n9112), .C1(n9013), .C2(n9114), .ZN(n9164) );
  NOR2_X1 U10297 ( .A1(n9164), .A2(n9433), .ZN(n9016) );
  AOI211_X1 U10298 ( .C1(n9162), .C2(n9100), .A(n9017), .B(n9016), .ZN(n9018)
         );
  OAI21_X1 U10299 ( .B1(n9165), .B2(n9121), .A(n9018), .ZN(P1_U3269) );
  AOI211_X1 U10300 ( .C1(n9168), .C2(n9042), .A(n9519), .B(n9019), .ZN(n9167)
         );
  NOR2_X1 U10301 ( .A1(n9436), .A2(n9020), .ZN(n9025) );
  XNOR2_X1 U10302 ( .A(n9021), .B(n9027), .ZN(n9023) );
  AOI21_X1 U10303 ( .B1(n9023), .B2(n9117), .A(n9022), .ZN(n9170) );
  INV_X1 U10304 ( .A(n9170), .ZN(n9024) );
  AOI211_X1 U10305 ( .C1(n9167), .C2(n9026), .A(n9025), .B(n9024), .ZN(n9034)
         );
  OR2_X1 U10306 ( .A1(n9028), .A2(n9027), .ZN(n9166) );
  NAND3_X1 U10307 ( .A1(n9166), .A2(n9029), .A3(n9077), .ZN(n9033) );
  AOI22_X1 U10308 ( .A1(n9168), .A2(n9031), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9030), .ZN(n9032) );
  OAI211_X1 U10309 ( .C1(n9433), .C2(n9034), .A(n9033), .B(n9032), .ZN(
        P1_U3270) );
  XOR2_X1 U10310 ( .A(n9037), .B(n9035), .Z(n9176) );
  NAND2_X1 U10311 ( .A1(n9052), .A2(n9036), .ZN(n9038) );
  XNOR2_X1 U10312 ( .A(n9038), .B(n9037), .ZN(n9039) );
  OAI222_X1 U10313 ( .A1(n9062), .A2(n9041), .B1(n9060), .B2(n9040), .C1(n9039), .C2(n9229), .ZN(n9172) );
  INV_X1 U10314 ( .A(n9174), .ZN(n9047) );
  INV_X1 U10315 ( .A(n9042), .ZN(n9043) );
  AOI211_X1 U10316 ( .C1(n9174), .C2(n9063), .A(n9519), .B(n9043), .ZN(n9173)
         );
  NAND2_X1 U10317 ( .A1(n9173), .A2(n9064), .ZN(n9046) );
  AOI22_X1 U10318 ( .A1(n9030), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9044), .B2(
        n9309), .ZN(n9045) );
  OAI211_X1 U10319 ( .C1(n9047), .C2(n9428), .A(n9046), .B(n9045), .ZN(n9048)
         );
  AOI21_X1 U10320 ( .B1(n9172), .B2(n9070), .A(n9048), .ZN(n9049) );
  OAI21_X1 U10321 ( .B1(n9176), .B2(n9121), .A(n9049), .ZN(P1_U3271) );
  XNOR2_X1 U10322 ( .A(n9050), .B(n9051), .ZN(n9181) );
  INV_X1 U10323 ( .A(n9052), .ZN(n9057) );
  AOI21_X1 U10324 ( .B1(n9055), .B2(n9054), .A(n9053), .ZN(n9056) );
  NOR2_X1 U10325 ( .A1(n9057), .A2(n9056), .ZN(n9058) );
  OAI222_X1 U10326 ( .A1(n9062), .A2(n9061), .B1(n9060), .B2(n9059), .C1(n9229), .C2(n9058), .ZN(n9177) );
  AOI211_X1 U10327 ( .C1(n9179), .C2(n9078), .A(n9519), .B(n4751), .ZN(n9178)
         );
  NAND2_X1 U10328 ( .A1(n9178), .A2(n9064), .ZN(n9067) );
  AOI22_X1 U10329 ( .A1(n9321), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9065), .B2(
        n9309), .ZN(n9066) );
  OAI211_X1 U10330 ( .C1(n9068), .C2(n9428), .A(n9067), .B(n9066), .ZN(n9069)
         );
  AOI21_X1 U10331 ( .B1(n9177), .B2(n9070), .A(n9069), .ZN(n9071) );
  OAI21_X1 U10332 ( .B1(n9181), .B2(n9121), .A(n9071), .ZN(P1_U3272) );
  XNOR2_X1 U10333 ( .A(n9072), .B(n9075), .ZN(n9074) );
  AOI222_X1 U10334 ( .A1(n9117), .A2(n9074), .B1(n9115), .B2(n9112), .C1(n9073), .C2(n9114), .ZN(n9187) );
  OR2_X1 U10335 ( .A1(n9076), .A2(n9075), .ZN(n9183) );
  NAND3_X1 U10336 ( .A1(n9183), .A2(n9182), .A3(n9077), .ZN(n9085) );
  INV_X1 U10337 ( .A(n9087), .ZN(n9079) );
  AOI21_X1 U10338 ( .B1(n9184), .B2(n9079), .A(n4747), .ZN(n9185) );
  AOI22_X1 U10339 ( .A1(n9321), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9080), .B2(
        n9309), .ZN(n9081) );
  OAI21_X1 U10340 ( .B1(n9082), .B2(n9428), .A(n9081), .ZN(n9083) );
  AOI21_X1 U10341 ( .B1(n9185), .B2(n9100), .A(n9083), .ZN(n9084) );
  OAI211_X1 U10342 ( .C1(n9433), .C2(n9187), .A(n9085), .B(n9084), .ZN(
        P1_U3273) );
  XNOR2_X1 U10343 ( .A(n9086), .B(n9093), .ZN(n9193) );
  INV_X1 U10344 ( .A(n9104), .ZN(n9088) );
  AOI21_X1 U10345 ( .B1(n9189), .B2(n9088), .A(n9087), .ZN(n9190) );
  AOI22_X1 U10346 ( .A1(n9321), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9089), .B2(
        n9309), .ZN(n9090) );
  OAI21_X1 U10347 ( .B1(n9091), .B2(n9428), .A(n9090), .ZN(n9099) );
  NAND2_X1 U10348 ( .A1(n9109), .A2(n9092), .ZN(n9094) );
  XNOR2_X1 U10349 ( .A(n9094), .B(n9093), .ZN(n9097) );
  AOI222_X1 U10350 ( .A1(n9117), .A2(n9097), .B1(n9096), .B2(n9114), .C1(n9095), .C2(n9112), .ZN(n9192) );
  NOR2_X1 U10351 ( .A1(n9192), .A2(n9030), .ZN(n9098) );
  AOI211_X1 U10352 ( .C1(n9190), .C2(n9100), .A(n9099), .B(n9098), .ZN(n9101)
         );
  OAI21_X1 U10353 ( .B1(n9193), .B2(n9121), .A(n9101), .ZN(P1_U3274) );
  XNOR2_X1 U10354 ( .A(n9103), .B(n9102), .ZN(n9198) );
  AOI211_X1 U10355 ( .C1(n9195), .C2(n9105), .A(n9519), .B(n9104), .ZN(n9194)
         );
  AOI22_X1 U10356 ( .A1(n9321), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9106), .B2(
        n9309), .ZN(n9107) );
  OAI21_X1 U10357 ( .B1(n9108), .B2(n9428), .A(n9107), .ZN(n9119) );
  OAI21_X1 U10358 ( .B1(n9111), .B2(n9110), .A(n9109), .ZN(n9116) );
  AOI222_X1 U10359 ( .A1(n9117), .A2(n9116), .B1(n9115), .B2(n9114), .C1(n9113), .C2(n9112), .ZN(n9197) );
  NOR2_X1 U10360 ( .A1(n9197), .A2(n9030), .ZN(n9118) );
  AOI211_X1 U10361 ( .C1(n9194), .C2(n9317), .A(n9119), .B(n9118), .ZN(n9120)
         );
  OAI21_X1 U10362 ( .B1(n9198), .B2(n9121), .A(n9120), .ZN(P1_U3275) );
  AOI21_X1 U10363 ( .B1(n9122), .B2(n9216), .A(n9395), .ZN(n9123) );
  OAI21_X1 U10364 ( .B1(n9124), .B2(n9519), .A(n9123), .ZN(n9242) );
  MUX2_X1 U10365 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9242), .S(n9544), .Z(
        P1_U3554) );
  NAND2_X1 U10366 ( .A1(n9125), .A2(n9515), .ZN(n9129) );
  MUX2_X1 U10367 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9243), .S(n9544), .Z(
        P1_U3552) );
  NAND2_X1 U10368 ( .A1(n9130), .A2(n9515), .ZN(n9135) );
  AOI22_X1 U10369 ( .A1(n9132), .A2(n9502), .B1(n9216), .B2(n9131), .ZN(n9133)
         );
  NAND3_X1 U10370 ( .A1(n9135), .A2(n9134), .A3(n9133), .ZN(n9244) );
  MUX2_X1 U10371 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9244), .S(n9544), .Z(
        P1_U3551) );
  AOI22_X1 U10372 ( .A1(n9137), .A2(n9502), .B1(n9216), .B2(n9136), .ZN(n9138)
         );
  OAI211_X1 U10373 ( .C1(n9140), .C2(n9208), .A(n9139), .B(n9138), .ZN(n9245)
         );
  MUX2_X1 U10374 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9245), .S(n9544), .Z(
        P1_U3550) );
  AOI22_X1 U10375 ( .A1(n9142), .A2(n9502), .B1(n9216), .B2(n9141), .ZN(n9143)
         );
  OAI211_X1 U10376 ( .C1(n9145), .C2(n9208), .A(n9144), .B(n9143), .ZN(n9246)
         );
  MUX2_X1 U10377 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9246), .S(n9544), .Z(
        P1_U3549) );
  AOI211_X1 U10378 ( .C1(n9216), .C2(n9148), .A(n9147), .B(n9146), .ZN(n9149)
         );
  OAI21_X1 U10379 ( .B1(n9150), .B2(n9208), .A(n9149), .ZN(n9247) );
  MUX2_X1 U10380 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9247), .S(n9544), .Z(
        P1_U3548) );
  AOI21_X1 U10381 ( .B1(n9216), .B2(n9152), .A(n9151), .ZN(n9153) );
  OAI211_X1 U10382 ( .C1(n9155), .C2(n9208), .A(n9154), .B(n9153), .ZN(n9248)
         );
  MUX2_X1 U10383 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9248), .S(n9544), .Z(
        P1_U3547) );
  AOI21_X1 U10384 ( .B1(n9216), .B2(n9157), .A(n9156), .ZN(n9158) );
  OAI211_X1 U10385 ( .C1(n9160), .C2(n9208), .A(n9159), .B(n9158), .ZN(n9249)
         );
  MUX2_X1 U10386 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9249), .S(n9544), .Z(
        P1_U3546) );
  AOI22_X1 U10387 ( .A1(n9162), .A2(n9502), .B1(n9216), .B2(n9161), .ZN(n9163)
         );
  OAI211_X1 U10388 ( .C1(n9165), .C2(n9208), .A(n9164), .B(n9163), .ZN(n9250)
         );
  MUX2_X1 U10389 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9250), .S(n9544), .Z(
        P1_U3545) );
  NAND3_X1 U10390 ( .A1(n9166), .A2(n9029), .A3(n9515), .ZN(n9171) );
  AOI21_X1 U10391 ( .B1(n9216), .B2(n9168), .A(n9167), .ZN(n9169) );
  NAND3_X1 U10392 ( .A1(n9171), .A2(n9170), .A3(n9169), .ZN(n9251) );
  MUX2_X1 U10393 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9251), .S(n9544), .Z(
        P1_U3544) );
  AOI211_X1 U10394 ( .C1(n9216), .C2(n9174), .A(n9173), .B(n9172), .ZN(n9175)
         );
  OAI21_X1 U10395 ( .B1(n9176), .B2(n9208), .A(n9175), .ZN(n9252) );
  MUX2_X1 U10396 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9252), .S(n9544), .Z(
        P1_U3543) );
  AOI211_X1 U10397 ( .C1(n9216), .C2(n9179), .A(n9178), .B(n9177), .ZN(n9180)
         );
  OAI21_X1 U10398 ( .B1(n9181), .B2(n9208), .A(n9180), .ZN(n9253) );
  MUX2_X1 U10399 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9253), .S(n9544), .Z(
        P1_U3542) );
  NAND3_X1 U10400 ( .A1(n9183), .A2(n9182), .A3(n9515), .ZN(n9188) );
  AOI22_X1 U10401 ( .A1(n9185), .A2(n9502), .B1(n9216), .B2(n9184), .ZN(n9186)
         );
  NAND3_X1 U10402 ( .A1(n9188), .A2(n9187), .A3(n9186), .ZN(n9254) );
  MUX2_X1 U10403 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9254), .S(n9544), .Z(
        P1_U3541) );
  AOI22_X1 U10404 ( .A1(n9190), .A2(n9502), .B1(n9216), .B2(n9189), .ZN(n9191)
         );
  OAI211_X1 U10405 ( .C1(n9193), .C2(n9208), .A(n9192), .B(n9191), .ZN(n9255)
         );
  MUX2_X1 U10406 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9255), .S(n9544), .Z(
        P1_U3540) );
  AOI21_X1 U10407 ( .B1(n9216), .B2(n9195), .A(n9194), .ZN(n9196) );
  OAI211_X1 U10408 ( .C1(n9198), .C2(n9208), .A(n9197), .B(n9196), .ZN(n9256)
         );
  MUX2_X1 U10409 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9256), .S(n9544), .Z(
        P1_U3539) );
  AOI22_X1 U10410 ( .A1(n9200), .A2(n9502), .B1(n9216), .B2(n9199), .ZN(n9201)
         );
  OAI211_X1 U10411 ( .C1(n9203), .C2(n9208), .A(n9202), .B(n9201), .ZN(n9257)
         );
  MUX2_X1 U10412 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9257), .S(n9544), .Z(
        P1_U3538) );
  AOI21_X1 U10413 ( .B1(n9216), .B2(n9205), .A(n9204), .ZN(n9206) );
  OAI211_X1 U10414 ( .C1(n9209), .C2(n9208), .A(n9207), .B(n9206), .ZN(n9258)
         );
  MUX2_X1 U10415 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9258), .S(n9544), .Z(
        P1_U3537) );
  AOI22_X1 U10416 ( .A1(n9211), .A2(n9502), .B1(n9216), .B2(n9210), .ZN(n9212)
         );
  OAI211_X1 U10417 ( .C1(n9505), .C2(n9214), .A(n9213), .B(n9212), .ZN(n9259)
         );
  MUX2_X1 U10418 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9259), .S(n9544), .Z(
        P1_U3536) );
  AOI22_X1 U10419 ( .A1(n9217), .A2(n9502), .B1(n9216), .B2(n9215), .ZN(n9218)
         );
  OAI211_X1 U10420 ( .C1(n9505), .C2(n9220), .A(n9219), .B(n9218), .ZN(n9260)
         );
  MUX2_X1 U10421 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9260), .S(n9544), .Z(
        P1_U3534) );
  NAND2_X1 U10422 ( .A1(n6641), .A2(n9221), .ZN(n9224) );
  AND2_X1 U10423 ( .A1(n9224), .A2(n9222), .ZN(n9226) );
  NAND2_X1 U10424 ( .A1(n9224), .A2(n9223), .ZN(n9225) );
  OAI21_X1 U10425 ( .B1(n9226), .B2(n9231), .A(n9225), .ZN(n9234) );
  INV_X1 U10426 ( .A(n9234), .ZN(n9314) );
  INV_X1 U10427 ( .A(n9227), .ZN(n9228) );
  AOI211_X1 U10428 ( .C1(n9231), .C2(n9230), .A(n9229), .B(n9228), .ZN(n9232)
         );
  AOI211_X1 U10429 ( .C1(n9234), .C2(n9478), .A(n9233), .B(n9232), .ZN(n9320)
         );
  INV_X1 U10430 ( .A(n9235), .ZN(n9238) );
  INV_X1 U10431 ( .A(n9236), .ZN(n9237) );
  AOI211_X1 U10432 ( .C1(n9239), .C2(n9238), .A(n9519), .B(n9237), .ZN(n9318)
         );
  AOI21_X1 U10433 ( .B1(n9216), .B2(n9239), .A(n9318), .ZN(n9240) );
  OAI211_X1 U10434 ( .C1(n9314), .C2(n9505), .A(n9320), .B(n9240), .ZN(n9261)
         );
  MUX2_X1 U10435 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n9261), .S(n9544), .Z(
        P1_U3533) );
  MUX2_X1 U10436 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9241), .S(n9544), .Z(
        P1_U3523) );
  MUX2_X1 U10437 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9242), .S(n9528), .Z(
        P1_U3522) );
  MUX2_X1 U10438 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9243), .S(n9528), .Z(
        P1_U3520) );
  MUX2_X1 U10439 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9244), .S(n9528), .Z(
        P1_U3519) );
  MUX2_X1 U10440 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9245), .S(n9528), .Z(
        P1_U3518) );
  MUX2_X1 U10441 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9246), .S(n9528), .Z(
        P1_U3517) );
  MUX2_X1 U10442 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9247), .S(n9528), .Z(
        P1_U3516) );
  MUX2_X1 U10443 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9248), .S(n9528), .Z(
        P1_U3515) );
  MUX2_X1 U10444 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9249), .S(n9528), .Z(
        P1_U3514) );
  MUX2_X1 U10445 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9250), .S(n9528), .Z(
        P1_U3513) );
  MUX2_X1 U10446 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9251), .S(n9528), .Z(
        P1_U3512) );
  MUX2_X1 U10447 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9252), .S(n9528), .Z(
        P1_U3511) );
  MUX2_X1 U10448 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9253), .S(n9528), .Z(
        P1_U3510) );
  MUX2_X1 U10449 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9254), .S(n9528), .Z(
        P1_U3508) );
  MUX2_X1 U10450 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9255), .S(n9528), .Z(
        P1_U3505) );
  MUX2_X1 U10451 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9256), .S(n9528), .Z(
        P1_U3502) );
  MUX2_X1 U10452 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9257), .S(n9528), .Z(
        P1_U3499) );
  MUX2_X1 U10453 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9258), .S(n9528), .Z(
        P1_U3496) );
  MUX2_X1 U10454 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9259), .S(n9528), .Z(
        P1_U3493) );
  MUX2_X1 U10455 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n9260), .S(n9528), .Z(
        P1_U3487) );
  MUX2_X1 U10456 ( .A(P1_REG0_REG_10__SCAN_IN), .B(n9261), .S(n9528), .Z(
        P1_U3484) );
  NOR2_X1 U10457 ( .A1(n9470), .A2(n9262), .ZN(n9453) );
  MUX2_X1 U10458 ( .A(P1_D_REG_0__SCAN_IN), .B(n9263), .S(n9467), .Z(P1_U3440)
         );
  NOR4_X1 U10459 ( .A1(n5401), .A2(P1_IR_REG_30__SCAN_IN), .A3(n5306), .A4(
        P1_U3084), .ZN(n9264) );
  AOI21_X1 U10460 ( .B1(n9265), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9264), .ZN(
        n9266) );
  OAI21_X1 U10461 ( .B1(n9267), .B2(n9273), .A(n9266), .ZN(P1_U3322) );
  INV_X1 U10462 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9271) );
  OAI222_X1 U10463 ( .A1(n9275), .A2(n9271), .B1(n9273), .B2(n9270), .C1(n9269), .C2(P1_U3084), .ZN(P1_U3323) );
  INV_X1 U10464 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9274) );
  OAI222_X1 U10465 ( .A1(n9275), .A2(n9274), .B1(P1_U3084), .B2(n5405), .C1(
        n9273), .C2(n9272), .ZN(P1_U3324) );
  MUX2_X1 U10466 ( .A(n9276), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AOI22_X1 U10467 ( .A1(n9578), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n9293) );
  NAND2_X1 U10468 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9277) );
  NAND2_X1 U10469 ( .A1(n9278), .A2(n9277), .ZN(n9281) );
  INV_X1 U10470 ( .A(n9279), .ZN(n9280) );
  NAND2_X1 U10471 ( .A1(n9281), .A2(n9280), .ZN(n9290) );
  NAND2_X1 U10472 ( .A1(n9295), .A2(n9282), .ZN(n9289) );
  INV_X1 U10473 ( .A(n9283), .ZN(n9287) );
  NAND2_X1 U10474 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9284) );
  NAND2_X1 U10475 ( .A1(n9285), .A2(n9284), .ZN(n9286) );
  NAND3_X1 U10476 ( .A1(n9573), .A2(n9287), .A3(n9286), .ZN(n9288) );
  OAI211_X1 U10477 ( .C1(n9290), .C2(n9576), .A(n9289), .B(n9288), .ZN(n9291)
         );
  INV_X1 U10478 ( .A(n9291), .ZN(n9292) );
  NAND2_X1 U10479 ( .A1(n9293), .A2(n9292), .ZN(P2_U3246) );
  AOI22_X1 U10480 ( .A1(n9578), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9308) );
  NAND2_X1 U10481 ( .A1(n9295), .A2(n9294), .ZN(n9306) );
  AND2_X1 U10482 ( .A1(n9297), .A2(n9296), .ZN(n9298) );
  OR3_X1 U10483 ( .A1(n9576), .A2(n9299), .A3(n9298), .ZN(n9305) );
  AOI21_X1 U10484 ( .B1(n9302), .B2(n9301), .A(n9300), .ZN(n9303) );
  NAND2_X1 U10485 ( .A1(n9573), .A2(n9303), .ZN(n9304) );
  AND3_X1 U10486 ( .A1(n9306), .A2(n9305), .A3(n9304), .ZN(n9307) );
  NAND2_X1 U10487 ( .A1(n9308), .A2(n9307), .ZN(P2_U3247) );
  AOI22_X1 U10488 ( .A1(n9433), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n9310), .B2(
        n9309), .ZN(n9311) );
  OAI21_X1 U10489 ( .B1(n9428), .B2(n9312), .A(n9311), .ZN(n9316) );
  NOR2_X1 U10490 ( .A1(n9314), .A2(n9313), .ZN(n9315) );
  AOI211_X1 U10491 ( .C1(n9318), .C2(n9317), .A(n9316), .B(n9315), .ZN(n9319)
         );
  OAI21_X1 U10492 ( .B1(n9321), .B2(n9320), .A(n9319), .ZN(P1_U3281) );
  OAI21_X1 U10493 ( .B1(n4785), .B2(n9323), .A(n9322), .ZN(n9329) );
  OAI21_X1 U10494 ( .B1(n9326), .B2(n9325), .A(n9324), .ZN(n9333) );
  NOR2_X1 U10495 ( .A1(n9333), .A2(n9691), .ZN(n9327) );
  AOI211_X1 U10496 ( .C1(n9619), .C2(n9329), .A(n9328), .B(n9327), .ZN(n9364)
         );
  INV_X1 U10497 ( .A(n9330), .ZN(n9331) );
  AOI222_X1 U10498 ( .A1(n9332), .A2(n9591), .B1(P2_REG2_REG_16__SCAN_IN), 
        .B2(n9590), .C1(n9613), .C2(n9331), .ZN(n9340) );
  INV_X1 U10499 ( .A(n9333), .ZN(n9367) );
  OAI21_X1 U10500 ( .B1(n9362), .B2(n9335), .A(n9334), .ZN(n9363) );
  INV_X1 U10501 ( .A(n9363), .ZN(n9336) );
  AOI22_X1 U10502 ( .A1(n9367), .A2(n9338), .B1(n9337), .B2(n9336), .ZN(n9339)
         );
  OAI211_X1 U10503 ( .C1(n9590), .C2(n9364), .A(n9340), .B(n9339), .ZN(
        P2_U3280) );
  INV_X1 U10504 ( .A(n9341), .ZN(n9347) );
  AOI21_X1 U10505 ( .B1(n9344), .B2(n9343), .A(n9342), .ZN(n9346) );
  NOR3_X1 U10506 ( .A1(n9347), .A2(n9346), .A3(n9345), .ZN(n9349) );
  NOR2_X1 U10507 ( .A1(n9349), .A2(n9348), .ZN(n9375) );
  INV_X1 U10508 ( .A(n9350), .ZN(n9351) );
  AOI222_X1 U10509 ( .A1(n9352), .A2(n9591), .B1(P2_REG2_REG_14__SCAN_IN), 
        .B2(n9590), .C1(n9613), .C2(n9351), .ZN(n9361) );
  OAI21_X1 U10510 ( .B1(n9355), .B2(n9354), .A(n9353), .ZN(n9378) );
  INV_X1 U10511 ( .A(n9356), .ZN(n9358) );
  OAI211_X1 U10512 ( .C1(n9358), .C2(n9376), .A(n9606), .B(n9357), .ZN(n9374)
         );
  INV_X1 U10513 ( .A(n9374), .ZN(n9359) );
  AOI22_X1 U10514 ( .A1(n9378), .A2(n9601), .B1(n9600), .B2(n9359), .ZN(n9360)
         );
  OAI211_X1 U10515 ( .C1(n9590), .C2(n9375), .A(n9361), .B(n9360), .ZN(
        P2_U3282) );
  INV_X1 U10516 ( .A(n9696), .ZN(n9709) );
  OAI22_X1 U10517 ( .A1(n9363), .A2(n4269), .B1(n9362), .B2(n9719), .ZN(n9366)
         );
  INV_X1 U10518 ( .A(n9364), .ZN(n9365) );
  AOI211_X1 U10519 ( .C1(n9709), .C2(n9367), .A(n9366), .B(n9365), .ZN(n9387)
         );
  AOI22_X1 U10520 ( .A1(n9745), .A2(n9387), .B1(n6983), .B2(n9742), .ZN(
        P2_U3536) );
  OAI22_X1 U10521 ( .A1(n9369), .A2(n4269), .B1(n9368), .B2(n9719), .ZN(n9370)
         );
  AOI211_X1 U10522 ( .C1(n9372), .C2(n9723), .A(n9371), .B(n9370), .ZN(n9389)
         );
  AOI22_X1 U10523 ( .A1(n9745), .A2(n9389), .B1(n9373), .B2(n9742), .ZN(
        P2_U3535) );
  OAI211_X1 U10524 ( .C1(n9376), .C2(n9719), .A(n9375), .B(n9374), .ZN(n9377)
         );
  AOI21_X1 U10525 ( .B1(n9723), .B2(n9378), .A(n9377), .ZN(n9390) );
  AOI22_X1 U10526 ( .A1(n9745), .A2(n9390), .B1(n6765), .B2(n9742), .ZN(
        P2_U3534) );
  INV_X1 U10527 ( .A(n9379), .ZN(n9384) );
  OAI22_X1 U10528 ( .A1(n9381), .A2(n5718), .B1(n9380), .B2(n9719), .ZN(n9383)
         );
  AOI211_X1 U10529 ( .C1(n9709), .C2(n9384), .A(n9383), .B(n9382), .ZN(n9392)
         );
  AOI22_X1 U10530 ( .A1(n9745), .A2(n9392), .B1(n9385), .B2(n9742), .ZN(
        P2_U3533) );
  INV_X1 U10531 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9386) );
  AOI22_X1 U10532 ( .A1(n9726), .A2(n9387), .B1(n9386), .B2(n9724), .ZN(
        P2_U3499) );
  INV_X1 U10533 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9388) );
  AOI22_X1 U10534 ( .A1(n9726), .A2(n9389), .B1(n9388), .B2(n9724), .ZN(
        P2_U3496) );
  AOI22_X1 U10535 ( .A1(n9726), .A2(n9390), .B1(n6766), .B2(n9724), .ZN(
        P2_U3493) );
  INV_X1 U10536 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9391) );
  AOI22_X1 U10537 ( .A1(n9726), .A2(n9392), .B1(n9391), .B2(n9724), .ZN(
        P2_U3490) );
  INV_X1 U10538 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9397) );
  AOI22_X1 U10539 ( .A1(n9544), .A2(n9407), .B1(n9397), .B2(n9541), .ZN(
        P1_U3553) );
  AOI211_X1 U10540 ( .C1(n9216), .C2(n9400), .A(n9399), .B(n9398), .ZN(n9401)
         );
  OAI21_X1 U10541 ( .B1(n9402), .B2(n9505), .A(n9401), .ZN(n9403) );
  AOI21_X1 U10542 ( .B1(n9478), .B2(n9404), .A(n9403), .ZN(n9409) );
  AOI22_X1 U10543 ( .A1(n9544), .A2(n9409), .B1(n9405), .B2(n9541), .ZN(
        P1_U3535) );
  INV_X1 U10544 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9406) );
  AOI22_X1 U10545 ( .A1(n9528), .A2(n9407), .B1(n9406), .B2(n9526), .ZN(
        P1_U3521) );
  INV_X1 U10546 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9408) );
  AOI22_X1 U10547 ( .A1(n9528), .A2(n9409), .B1(n9408), .B2(n9526), .ZN(
        P1_U3490) );
  XNOR2_X1 U10548 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  INV_X1 U10549 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9859) );
  INV_X1 U10550 ( .A(n9410), .ZN(n9411) );
  AOI21_X1 U10551 ( .B1(n9413), .B2(n9412), .A(n9411), .ZN(n9425) );
  OAI21_X1 U10552 ( .B1(n9416), .B2(n9415), .A(n9414), .ZN(n9423) );
  OAI21_X1 U10553 ( .B1(n9419), .B2(n9418), .A(n9417), .ZN(n9420) );
  AOI22_X1 U10554 ( .A1(n9423), .A2(n9422), .B1(n9421), .B2(n9420), .ZN(n9424)
         );
  OAI211_X1 U10555 ( .C1(n9426), .C2(n9859), .A(n9425), .B(n9424), .ZN(
        P1_U3255) );
  AOI21_X1 U10556 ( .B1(n9429), .B2(n9428), .A(n9427), .ZN(n9432) );
  NOR2_X1 U10557 ( .A1(n9430), .A2(n9433), .ZN(n9431) );
  AOI211_X1 U10558 ( .C1(n9433), .C2(P1_REG2_REG_0__SCAN_IN), .A(n9432), .B(
        n9431), .ZN(n9434) );
  OAI21_X1 U10559 ( .B1(n9436), .B2(n9435), .A(n9434), .ZN(P1_U3291) );
  INV_X1 U10560 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n9437) );
  NOR2_X1 U10561 ( .A1(n9453), .A2(n9437), .ZN(P1_U3292) );
  INV_X1 U10562 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n9438) );
  NOR2_X1 U10563 ( .A1(n9453), .A2(n9438), .ZN(P1_U3293) );
  INV_X1 U10564 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n9439) );
  NOR2_X1 U10565 ( .A1(n9467), .A2(n9439), .ZN(P1_U3294) );
  INV_X1 U10566 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n9440) );
  NOR2_X1 U10567 ( .A1(n9467), .A2(n9440), .ZN(P1_U3295) );
  INV_X1 U10568 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n9441) );
  NOR2_X1 U10569 ( .A1(n9467), .A2(n9441), .ZN(P1_U3296) );
  INV_X1 U10570 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n9806) );
  NOR2_X1 U10571 ( .A1(n9467), .A2(n9806), .ZN(P1_U3297) );
  INV_X1 U10572 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n9442) );
  NOR2_X1 U10573 ( .A1(n9467), .A2(n9442), .ZN(P1_U3298) );
  INV_X1 U10574 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n9443) );
  NOR2_X1 U10575 ( .A1(n9467), .A2(n9443), .ZN(P1_U3299) );
  INV_X1 U10576 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n9444) );
  NOR2_X1 U10577 ( .A1(n9467), .A2(n9444), .ZN(P1_U3300) );
  INV_X1 U10578 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n9445) );
  NOR2_X1 U10579 ( .A1(n9453), .A2(n9445), .ZN(P1_U3301) );
  INV_X1 U10580 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n9446) );
  NOR2_X1 U10581 ( .A1(n9453), .A2(n9446), .ZN(P1_U3302) );
  INV_X1 U10582 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n9447) );
  NOR2_X1 U10583 ( .A1(n9453), .A2(n9447), .ZN(P1_U3303) );
  INV_X1 U10584 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n9448) );
  NOR2_X1 U10585 ( .A1(n9453), .A2(n9448), .ZN(P1_U3304) );
  INV_X1 U10586 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n9449) );
  NOR2_X1 U10587 ( .A1(n9453), .A2(n9449), .ZN(P1_U3305) );
  INV_X1 U10588 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n9450) );
  NOR2_X1 U10589 ( .A1(n9453), .A2(n9450), .ZN(P1_U3306) );
  INV_X1 U10590 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n9451) );
  NOR2_X1 U10591 ( .A1(n9453), .A2(n9451), .ZN(P1_U3307) );
  INV_X1 U10592 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n9452) );
  NOR2_X1 U10593 ( .A1(n9453), .A2(n9452), .ZN(P1_U3308) );
  INV_X1 U10594 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n9454) );
  NOR2_X1 U10595 ( .A1(n9467), .A2(n9454), .ZN(P1_U3309) );
  INV_X1 U10596 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n9455) );
  NOR2_X1 U10597 ( .A1(n9467), .A2(n9455), .ZN(P1_U3310) );
  INV_X1 U10598 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n9456) );
  NOR2_X1 U10599 ( .A1(n9467), .A2(n9456), .ZN(P1_U3311) );
  INV_X1 U10600 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n9457) );
  NOR2_X1 U10601 ( .A1(n9467), .A2(n9457), .ZN(P1_U3312) );
  INV_X1 U10602 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n9458) );
  NOR2_X1 U10603 ( .A1(n9467), .A2(n9458), .ZN(P1_U3313) );
  INV_X1 U10604 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n9459) );
  NOR2_X1 U10605 ( .A1(n9467), .A2(n9459), .ZN(P1_U3314) );
  INV_X1 U10606 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n9460) );
  NOR2_X1 U10607 ( .A1(n9467), .A2(n9460), .ZN(P1_U3315) );
  INV_X1 U10608 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n9461) );
  NOR2_X1 U10609 ( .A1(n9467), .A2(n9461), .ZN(P1_U3316) );
  INV_X1 U10610 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n9462) );
  NOR2_X1 U10611 ( .A1(n9467), .A2(n9462), .ZN(P1_U3317) );
  INV_X1 U10612 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n9463) );
  NOR2_X1 U10613 ( .A1(n9467), .A2(n9463), .ZN(P1_U3318) );
  INV_X1 U10614 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n9464) );
  NOR2_X1 U10615 ( .A1(n9467), .A2(n9464), .ZN(P1_U3319) );
  INV_X1 U10616 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n9465) );
  NOR2_X1 U10617 ( .A1(n9467), .A2(n9465), .ZN(P1_U3320) );
  INV_X1 U10618 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n9466) );
  NOR2_X1 U10619 ( .A1(n9467), .A2(n9466), .ZN(P1_U3321) );
  AOI21_X1 U10620 ( .B1(n9470), .B2(n9469), .A(n9468), .ZN(P1_U3441) );
  INV_X1 U10621 ( .A(n9475), .ZN(n9477) );
  AOI211_X1 U10622 ( .C1(n9216), .C2(n9473), .A(n9472), .B(n9471), .ZN(n9474)
         );
  OAI21_X1 U10623 ( .B1(n9505), .B2(n9475), .A(n9474), .ZN(n9476) );
  AOI21_X1 U10624 ( .B1(n9478), .B2(n9477), .A(n9476), .ZN(n9530) );
  INV_X1 U10625 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9479) );
  AOI22_X1 U10626 ( .A1(n9528), .A2(n9530), .B1(n9479), .B2(n9526), .ZN(
        P1_U3457) );
  AOI22_X1 U10627 ( .A1(n9481), .A2(n9502), .B1(n9216), .B2(n9480), .ZN(n9482)
         );
  OAI211_X1 U10628 ( .C1(n9484), .C2(n9505), .A(n9483), .B(n9482), .ZN(n9485)
         );
  INV_X1 U10629 ( .A(n9485), .ZN(n9532) );
  INV_X1 U10630 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9486) );
  AOI22_X1 U10631 ( .A1(n9528), .A2(n9532), .B1(n9486), .B2(n9526), .ZN(
        P1_U3460) );
  INV_X1 U10632 ( .A(n9505), .ZN(n9522) );
  INV_X1 U10633 ( .A(n9487), .ZN(n9492) );
  OAI22_X1 U10634 ( .A1(n9489), .A2(n9519), .B1(n9488), .B2(n9517), .ZN(n9491)
         );
  AOI211_X1 U10635 ( .C1(n9522), .C2(n9492), .A(n9491), .B(n9490), .ZN(n9534)
         );
  INV_X1 U10636 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9493) );
  AOI22_X1 U10637 ( .A1(n9528), .A2(n9534), .B1(n9493), .B2(n9526), .ZN(
        P1_U3466) );
  AOI21_X1 U10638 ( .B1(n9216), .B2(n9495), .A(n9494), .ZN(n9498) );
  NAND3_X1 U10639 ( .A1(n6144), .A2(n9496), .A3(n9515), .ZN(n9497) );
  AND3_X1 U10640 ( .A1(n9499), .A2(n9498), .A3(n9497), .ZN(n9536) );
  INV_X1 U10641 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9500) );
  AOI22_X1 U10642 ( .A1(n9528), .A2(n9536), .B1(n9500), .B2(n9526), .ZN(
        P1_U3469) );
  AOI22_X1 U10643 ( .A1(n9503), .A2(n9502), .B1(n9216), .B2(n9501), .ZN(n9504)
         );
  OAI21_X1 U10644 ( .B1(n9506), .B2(n9505), .A(n9504), .ZN(n9508) );
  NOR2_X1 U10645 ( .A1(n9508), .A2(n9507), .ZN(n9538) );
  INV_X1 U10646 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9509) );
  AOI22_X1 U10647 ( .A1(n9528), .A2(n9538), .B1(n9509), .B2(n9526), .ZN(
        P1_U3472) );
  OAI21_X1 U10648 ( .B1(n9511), .B2(n9517), .A(n9510), .ZN(n9513) );
  AOI211_X1 U10649 ( .C1(n9515), .C2(n9514), .A(n9513), .B(n9512), .ZN(n9540)
         );
  INV_X1 U10650 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9516) );
  AOI22_X1 U10651 ( .A1(n9528), .A2(n9540), .B1(n9516), .B2(n9526), .ZN(
        P1_U3475) );
  OAI22_X1 U10652 ( .A1(n9520), .A2(n9519), .B1(n9518), .B2(n9517), .ZN(n9521)
         );
  AOI21_X1 U10653 ( .B1(n9523), .B2(n9522), .A(n9521), .ZN(n9524) );
  AND2_X1 U10654 ( .A1(n9525), .A2(n9524), .ZN(n9543) );
  INV_X1 U10655 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9527) );
  AOI22_X1 U10656 ( .A1(n9528), .A2(n9543), .B1(n9527), .B2(n9526), .ZN(
        P1_U3478) );
  INV_X1 U10657 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9529) );
  AOI22_X1 U10658 ( .A1(n9544), .A2(n9530), .B1(n9529), .B2(n9541), .ZN(
        P1_U3524) );
  AOI22_X1 U10659 ( .A1(n9544), .A2(n9532), .B1(n9531), .B2(n9541), .ZN(
        P1_U3525) );
  AOI22_X1 U10660 ( .A1(n9544), .A2(n9534), .B1(n9533), .B2(n9541), .ZN(
        P1_U3527) );
  INV_X1 U10661 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9535) );
  AOI22_X1 U10662 ( .A1(n9544), .A2(n9536), .B1(n9535), .B2(n9541), .ZN(
        P1_U3528) );
  AOI22_X1 U10663 ( .A1(n9544), .A2(n9538), .B1(n9537), .B2(n9541), .ZN(
        P1_U3529) );
  AOI22_X1 U10664 ( .A1(n9544), .A2(n9540), .B1(n9539), .B2(n9541), .ZN(
        P1_U3530) );
  AOI22_X1 U10665 ( .A1(n9544), .A2(n9543), .B1(n9542), .B2(n9541), .ZN(
        P1_U3531) );
  INV_X1 U10666 ( .A(n9545), .ZN(n9546) );
  AOI22_X1 U10667 ( .A1(n9559), .A2(n9546), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3152), .ZN(n9555) );
  INV_X1 U10668 ( .A(n9547), .ZN(n9549) );
  NAND2_X1 U10669 ( .A1(n9549), .A2(n9548), .ZN(n9550) );
  XNOR2_X1 U10670 ( .A(n9551), .B(n9550), .ZN(n9553) );
  AOI22_X1 U10671 ( .A1(n9553), .A2(n9566), .B1(n9565), .B2(n9552), .ZN(n9554)
         );
  OAI211_X1 U10672 ( .C1(n9571), .C2(n9556), .A(n9555), .B(n9554), .ZN(
        P2_U3232) );
  INV_X1 U10673 ( .A(n9557), .ZN(n9558) );
  AOI22_X1 U10674 ( .A1(n9559), .A2(n9558), .B1(P2_REG3_REG_9__SCAN_IN), .B2(
        P2_U3152), .ZN(n9569) );
  INV_X1 U10675 ( .A(n9560), .ZN(n9562) );
  NAND2_X1 U10676 ( .A1(n9562), .A2(n9561), .ZN(n9563) );
  XNOR2_X1 U10677 ( .A(n9564), .B(n9563), .ZN(n9567) );
  AOI22_X1 U10678 ( .A1(n9567), .A2(n9566), .B1(n9565), .B2(n9693), .ZN(n9568)
         );
  OAI211_X1 U10679 ( .C1(n9571), .C2(n9570), .A(n9569), .B(n9568), .ZN(
        P2_U3233) );
  AOI22_X1 U10680 ( .A1(n9572), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9573), .ZN(n9582) );
  NAND2_X1 U10681 ( .A1(n9573), .A2(n9727), .ZN(n9574) );
  OAI211_X1 U10682 ( .C1(P2_REG2_REG_0__SCAN_IN), .C2(n9576), .A(n9575), .B(
        n9574), .ZN(n9577) );
  INV_X1 U10683 ( .A(n9577), .ZN(n9580) );
  AOI22_X1 U10684 ( .A1(n9578), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9579) );
  OAI221_X1 U10685 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9582), .C1(n9581), .C2(
        n9580), .A(n9579), .ZN(P2_U3245) );
  NAND2_X1 U10686 ( .A1(n9584), .A2(n9583), .ZN(n9585) );
  XOR2_X1 U10687 ( .A(n9593), .B(n9585), .Z(n9587) );
  AOI21_X1 U10688 ( .B1(n9587), .B2(n9619), .A(n9586), .ZN(n9718) );
  INV_X1 U10689 ( .A(n9588), .ZN(n9589) );
  AOI222_X1 U10690 ( .A1(n9592), .A2(n9591), .B1(P2_REG2_REG_12__SCAN_IN), 
        .B2(n9590), .C1(n9613), .C2(n9589), .ZN(n9603) );
  OAI21_X1 U10691 ( .B1(n9595), .B2(n6779), .A(n9594), .ZN(n9722) );
  INV_X1 U10692 ( .A(n9596), .ZN(n9597) );
  OAI211_X1 U10693 ( .C1(n9720), .C2(n9598), .A(n9597), .B(n9606), .ZN(n9717)
         );
  INV_X1 U10694 ( .A(n9717), .ZN(n9599) );
  AOI22_X1 U10695 ( .A1(n9722), .A2(n9601), .B1(n9600), .B2(n9599), .ZN(n9602)
         );
  OAI211_X1 U10696 ( .C1(n9590), .C2(n9718), .A(n9603), .B(n9602), .ZN(
        P2_U3284) );
  XNOR2_X1 U10697 ( .A(n9604), .B(n9617), .ZN(n9667) );
  NAND2_X1 U10698 ( .A1(n9605), .A2(n9610), .ZN(n9607) );
  NAND2_X1 U10699 ( .A1(n9607), .A2(n9606), .ZN(n9608) );
  OR2_X1 U10700 ( .A1(n9609), .A2(n9608), .ZN(n9668) );
  AOI22_X1 U10701 ( .A1(n9613), .A2(n9612), .B1(n9611), .B2(n9610), .ZN(n9614)
         );
  OAI21_X1 U10702 ( .B1(n9668), .B2(n5547), .A(n9614), .ZN(n9627) );
  NAND2_X1 U10703 ( .A1(n9616), .A2(n9615), .ZN(n9618) );
  XNOR2_X1 U10704 ( .A(n9618), .B(n9617), .ZN(n9620) );
  NAND2_X1 U10705 ( .A1(n9620), .A2(n9619), .ZN(n9626) );
  AOI22_X1 U10706 ( .A1(n9624), .A2(n9623), .B1(n9622), .B2(n9621), .ZN(n9625)
         );
  NAND2_X1 U10707 ( .A1(n9626), .A2(n9625), .ZN(n9672) );
  AOI211_X1 U10708 ( .C1(n9628), .C2(n9667), .A(n9627), .B(n9672), .ZN(n9629)
         );
  AOI22_X1 U10709 ( .A1(n8217), .A2(n5711), .B1(n9629), .B2(n8265), .ZN(
        P2_U3291) );
  NOR2_X1 U10710 ( .A1(n9631), .A2(n9630), .ZN(n9632) );
  AND2_X1 U10711 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9887), .ZN(P2_U3297) );
  AND2_X1 U10712 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9887), .ZN(P2_U3298) );
  AND2_X1 U10713 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9887), .ZN(P2_U3299) );
  AND2_X1 U10714 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9887), .ZN(P2_U3300) );
  INV_X1 U10715 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n9868) );
  NOR2_X1 U10716 ( .A1(n9632), .A2(n9868), .ZN(P2_U3301) );
  AND2_X1 U10717 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9887), .ZN(P2_U3302) );
  AND2_X1 U10718 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9887), .ZN(P2_U3303) );
  AND2_X1 U10719 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9887), .ZN(P2_U3304) );
  AND2_X1 U10720 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9887), .ZN(P2_U3305) );
  AND2_X1 U10721 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9887), .ZN(P2_U3306) );
  AND2_X1 U10722 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9887), .ZN(P2_U3307) );
  AND2_X1 U10723 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9887), .ZN(P2_U3308) );
  AND2_X1 U10724 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9887), .ZN(P2_U3309) );
  AND2_X1 U10725 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9887), .ZN(P2_U3310) );
  AND2_X1 U10726 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9887), .ZN(P2_U3311) );
  AND2_X1 U10727 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9887), .ZN(P2_U3312) );
  AND2_X1 U10728 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9887), .ZN(P2_U3313) );
  AND2_X1 U10729 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9887), .ZN(P2_U3314) );
  INV_X1 U10730 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n9802) );
  NOR2_X1 U10731 ( .A1(n9632), .A2(n9802), .ZN(P2_U3315) );
  AND2_X1 U10732 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9887), .ZN(P2_U3316) );
  AND2_X1 U10733 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9887), .ZN(P2_U3317) );
  AND2_X1 U10734 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9887), .ZN(P2_U3318) );
  AND2_X1 U10735 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9887), .ZN(P2_U3320) );
  AND2_X1 U10736 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9887), .ZN(P2_U3321) );
  AND2_X1 U10737 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9887), .ZN(P2_U3322) );
  AND2_X1 U10738 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9887), .ZN(P2_U3323) );
  AND2_X1 U10739 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9887), .ZN(P2_U3324) );
  AND2_X1 U10740 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9887), .ZN(P2_U3325) );
  AND2_X1 U10741 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9887), .ZN(P2_U3326) );
  AOI22_X1 U10742 ( .A1(n9634), .A2(n9887), .B1(n9637), .B2(n9633), .ZN(
        P2_U3437) );
  AOI22_X1 U10743 ( .A1(n9637), .A2(n9636), .B1(n9635), .B2(n9887), .ZN(
        P2_U3438) );
  AOI22_X1 U10744 ( .A1(n9640), .A2(n9723), .B1(n9639), .B2(n9638), .ZN(n9641)
         );
  AND2_X1 U10745 ( .A1(n9642), .A2(n9641), .ZN(n9728) );
  AOI22_X1 U10746 ( .A1(n9726), .A2(n9728), .B1(n5087), .B2(n9724), .ZN(
        P2_U3451) );
  INV_X1 U10747 ( .A(n9643), .ZN(n9645) );
  OAI22_X1 U10748 ( .A1(n9645), .A2(n4269), .B1(n5919), .B2(n9719), .ZN(n9647)
         );
  AOI211_X1 U10749 ( .C1(n9648), .C2(n9723), .A(n9647), .B(n9646), .ZN(n9729)
         );
  AOI22_X1 U10750 ( .A1(n9726), .A2(n9729), .B1(n5555), .B2(n9724), .ZN(
        P2_U3454) );
  NAND2_X1 U10751 ( .A1(n9649), .A2(n9694), .ZN(n9650) );
  AND2_X1 U10752 ( .A1(n9651), .A2(n9650), .ZN(n9655) );
  OR2_X1 U10753 ( .A1(n9653), .A2(n9652), .ZN(n9654) );
  AND3_X1 U10754 ( .A1(n9656), .A2(n9655), .A3(n9654), .ZN(n9730) );
  AOI22_X1 U10755 ( .A1(n9726), .A2(n9730), .B1(n5578), .B2(n9724), .ZN(
        P2_U3457) );
  OAI22_X1 U10756 ( .A1(n9658), .A2(n4269), .B1(n9657), .B2(n9719), .ZN(n9660)
         );
  AOI211_X1 U10757 ( .C1(n9709), .C2(n9661), .A(n9660), .B(n9659), .ZN(n9732)
         );
  AOI22_X1 U10758 ( .A1(n9726), .A2(n9732), .B1(n5684), .B2(n9724), .ZN(
        P2_U3460) );
  OAI21_X1 U10759 ( .B1(n9663), .B2(n9719), .A(n9662), .ZN(n9665) );
  AOI211_X1 U10760 ( .C1(n9723), .C2(n9666), .A(n9665), .B(n9664), .ZN(n9733)
         );
  AOI22_X1 U10761 ( .A1(n9726), .A2(n9733), .B1(n5703), .B2(n9724), .ZN(
        P2_U3463) );
  AND2_X1 U10762 ( .A1(n9667), .A2(n9723), .ZN(n9671) );
  OAI21_X1 U10763 ( .B1(n9669), .B2(n9719), .A(n9668), .ZN(n9670) );
  NOR3_X1 U10764 ( .A1(n9672), .A2(n9671), .A3(n9670), .ZN(n9734) );
  INV_X1 U10765 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9673) );
  AOI22_X1 U10766 ( .A1(n9726), .A2(n9734), .B1(n9673), .B2(n9724), .ZN(
        P2_U3466) );
  OAI211_X1 U10767 ( .C1(n9676), .C2(n9719), .A(n9675), .B(n9674), .ZN(n9677)
         );
  AOI21_X1 U10768 ( .B1(n9723), .B2(n9678), .A(n9677), .ZN(n9736) );
  INV_X1 U10769 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9679) );
  AOI22_X1 U10770 ( .A1(n9726), .A2(n9736), .B1(n9679), .B2(n9724), .ZN(
        P2_U3469) );
  OAI211_X1 U10771 ( .C1(n9682), .C2(n9719), .A(n9681), .B(n9680), .ZN(n9683)
         );
  AOI21_X1 U10772 ( .B1(n9723), .B2(n9684), .A(n9683), .ZN(n9737) );
  INV_X1 U10773 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9685) );
  AOI22_X1 U10774 ( .A1(n9726), .A2(n9737), .B1(n9685), .B2(n9724), .ZN(
        P2_U3472) );
  OAI22_X1 U10775 ( .A1(n9686), .A2(n5718), .B1(n4449), .B2(n9719), .ZN(n9688)
         );
  AOI211_X1 U10776 ( .C1(n9723), .C2(n9689), .A(n9688), .B(n9687), .ZN(n9738)
         );
  INV_X1 U10777 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9690) );
  AOI22_X1 U10778 ( .A1(n9726), .A2(n9738), .B1(n9690), .B2(n9724), .ZN(
        P2_U3475) );
  INV_X1 U10779 ( .A(n9691), .ZN(n9701) );
  INV_X1 U10780 ( .A(n9697), .ZN(n9700) );
  AOI21_X1 U10781 ( .B1(n9694), .B2(n9693), .A(n9692), .ZN(n9695) );
  OAI21_X1 U10782 ( .B1(n9697), .B2(n9696), .A(n9695), .ZN(n9698) );
  AOI211_X1 U10783 ( .C1(n9701), .C2(n9700), .A(n9699), .B(n9698), .ZN(n9739)
         );
  AOI22_X1 U10784 ( .A1(n9726), .A2(n9739), .B1(n5911), .B2(n9724), .ZN(
        P2_U3478) );
  INV_X1 U10785 ( .A(n9702), .ZN(n9708) );
  INV_X1 U10786 ( .A(n9703), .ZN(n9704) );
  OAI22_X1 U10787 ( .A1(n9705), .A2(n4269), .B1(n9704), .B2(n9719), .ZN(n9707)
         );
  AOI211_X1 U10788 ( .C1(n9709), .C2(n9708), .A(n9707), .B(n9706), .ZN(n9740)
         );
  INV_X1 U10789 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9710) );
  AOI22_X1 U10790 ( .A1(n9726), .A2(n9740), .B1(n9710), .B2(n9724), .ZN(
        P2_U3481) );
  OAI21_X1 U10791 ( .B1(n9712), .B2(n9719), .A(n9711), .ZN(n9714) );
  AOI211_X1 U10792 ( .C1(n9715), .C2(n9723), .A(n9714), .B(n9713), .ZN(n9741)
         );
  INV_X1 U10793 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9716) );
  AOI22_X1 U10794 ( .A1(n9726), .A2(n9741), .B1(n9716), .B2(n9724), .ZN(
        P2_U3484) );
  OAI211_X1 U10795 ( .C1(n9720), .C2(n9719), .A(n9718), .B(n9717), .ZN(n9721)
         );
  AOI21_X1 U10796 ( .B1(n9723), .B2(n9722), .A(n9721), .ZN(n9744) );
  INV_X1 U10797 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9725) );
  AOI22_X1 U10798 ( .A1(n9726), .A2(n9744), .B1(n9725), .B2(n9724), .ZN(
        P2_U3487) );
  AOI22_X1 U10799 ( .A1(n9745), .A2(n9728), .B1(n9727), .B2(n9742), .ZN(
        P2_U3520) );
  AOI22_X1 U10800 ( .A1(n9745), .A2(n9729), .B1(n9794), .B2(n9742), .ZN(
        P2_U3521) );
  AOI22_X1 U10801 ( .A1(n9745), .A2(n9730), .B1(n5190), .B2(n9742), .ZN(
        P2_U3522) );
  INV_X1 U10802 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9731) );
  AOI22_X1 U10803 ( .A1(n9745), .A2(n9732), .B1(n9731), .B2(n9742), .ZN(
        P2_U3523) );
  AOI22_X1 U10804 ( .A1(n9745), .A2(n9733), .B1(n5210), .B2(n9742), .ZN(
        P2_U3524) );
  AOI22_X1 U10805 ( .A1(n9745), .A2(n9734), .B1(n5710), .B2(n9742), .ZN(
        P2_U3525) );
  AOI22_X1 U10806 ( .A1(n9745), .A2(n9736), .B1(n9735), .B2(n9742), .ZN(
        P2_U3526) );
  AOI22_X1 U10807 ( .A1(n9745), .A2(n9737), .B1(n5804), .B2(n9742), .ZN(
        P2_U3527) );
  AOI22_X1 U10808 ( .A1(n9745), .A2(n9738), .B1(n5945), .B2(n9742), .ZN(
        P2_U3528) );
  INV_X1 U10809 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9855) );
  AOI22_X1 U10810 ( .A1(n9745), .A2(n9739), .B1(n9855), .B2(n9742), .ZN(
        P2_U3529) );
  AOI22_X1 U10811 ( .A1(n9745), .A2(n9740), .B1(n5588), .B2(n9742), .ZN(
        P2_U3530) );
  AOI22_X1 U10812 ( .A1(n9745), .A2(n9741), .B1(n6285), .B2(n9742), .ZN(
        P2_U3531) );
  AOI22_X1 U10813 ( .A1(n9745), .A2(n9744), .B1(n9743), .B2(n9742), .ZN(
        P2_U3532) );
  INV_X1 U10814 ( .A(n9746), .ZN(n9747) );
  NAND2_X1 U10815 ( .A1(n9748), .A2(n9747), .ZN(n9749) );
  XOR2_X1 U10816 ( .A(n9897), .B(n9749), .Z(ADD_1071_U5) );
  XOR2_X1 U10817 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U10818 ( .B1(n9752), .B2(n9751), .A(n9750), .ZN(ADD_1071_U56) );
  OAI21_X1 U10819 ( .B1(n9755), .B2(n9754), .A(n9753), .ZN(ADD_1071_U57) );
  OAI21_X1 U10820 ( .B1(n9758), .B2(n9757), .A(n9756), .ZN(ADD_1071_U58) );
  OAI21_X1 U10821 ( .B1(n9761), .B2(n9760), .A(n9759), .ZN(ADD_1071_U59) );
  OAI21_X1 U10822 ( .B1(n9764), .B2(n9763), .A(n9762), .ZN(ADD_1071_U60) );
  OAI21_X1 U10823 ( .B1(n9767), .B2(n9766), .A(n9765), .ZN(ADD_1071_U61) );
  AOI21_X1 U10824 ( .B1(n9770), .B2(n9769), .A(n9768), .ZN(ADD_1071_U62) );
  AOI21_X1 U10825 ( .B1(n9773), .B2(n9772), .A(n9771), .ZN(ADD_1071_U63) );
  INV_X1 U10826 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9775) );
  AOI22_X1 U10827 ( .A1(P2_U3152), .A2(keyinput57), .B1(keyinput61), .B2(n9775), .ZN(n9774) );
  OAI221_X1 U10828 ( .B1(P2_U3152), .B2(keyinput57), .C1(n9775), .C2(
        keyinput61), .A(n9774), .ZN(n9787) );
  AOI22_X1 U10829 ( .A1(n9778), .A2(keyinput5), .B1(n8883), .B2(keyinput6), 
        .ZN(n9777) );
  OAI221_X1 U10830 ( .B1(n9778), .B2(keyinput5), .C1(n8883), .C2(keyinput6), 
        .A(n9777), .ZN(n9786) );
  AOI22_X1 U10831 ( .A1(n9781), .A2(keyinput18), .B1(n9780), .B2(keyinput48), 
        .ZN(n9779) );
  OAI221_X1 U10832 ( .B1(n9781), .B2(keyinput18), .C1(n9780), .C2(keyinput48), 
        .A(n9779), .ZN(n9785) );
  XNOR2_X1 U10833 ( .A(P2_IR_REG_26__SCAN_IN), .B(keyinput8), .ZN(n9783) );
  XNOR2_X1 U10834 ( .A(P1_REG3_REG_14__SCAN_IN), .B(keyinput21), .ZN(n9782) );
  NAND2_X1 U10835 ( .A1(n9783), .A2(n9782), .ZN(n9784) );
  NOR4_X1 U10836 ( .A1(n9787), .A2(n9786), .A3(n9785), .A4(n9784), .ZN(n9828)
         );
  AOI22_X1 U10837 ( .A1(n9892), .A2(keyinput53), .B1(keyinput32), .B2(n5210), 
        .ZN(n9788) );
  OAI221_X1 U10838 ( .B1(n9892), .B2(keyinput53), .C1(n5210), .C2(keyinput32), 
        .A(n9788), .ZN(n9800) );
  INV_X1 U10839 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n9790) );
  AOI22_X1 U10840 ( .A1(n9791), .A2(keyinput24), .B1(keyinput46), .B2(n9790), 
        .ZN(n9789) );
  OAI221_X1 U10841 ( .B1(n9791), .B2(keyinput24), .C1(n9790), .C2(keyinput46), 
        .A(n9789), .ZN(n9799) );
  INV_X1 U10842 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9793) );
  AOI22_X1 U10843 ( .A1(n9794), .A2(keyinput55), .B1(n9793), .B2(keyinput39), 
        .ZN(n9792) );
  OAI221_X1 U10844 ( .B1(n9794), .B2(keyinput55), .C1(n9793), .C2(keyinput39), 
        .A(n9792), .ZN(n9798) );
  XOR2_X1 U10845 ( .A(n6766), .B(keyinput20), .Z(n9796) );
  XNOR2_X1 U10846 ( .A(P1_RD_REG_SCAN_IN), .B(keyinput29), .ZN(n9795) );
  NAND2_X1 U10847 ( .A1(n9796), .A2(n9795), .ZN(n9797) );
  NOR4_X1 U10848 ( .A1(n9800), .A2(n9799), .A3(n9798), .A4(n9797), .ZN(n9827)
         );
  AOI22_X1 U10849 ( .A1(n9803), .A2(keyinput2), .B1(keyinput17), .B2(n9802), 
        .ZN(n9801) );
  OAI221_X1 U10850 ( .B1(n9803), .B2(keyinput2), .C1(n9802), .C2(keyinput17), 
        .A(n9801), .ZN(n9813) );
  AOI22_X1 U10851 ( .A1(n9806), .A2(keyinput22), .B1(keyinput37), .B2(n9805), 
        .ZN(n9804) );
  OAI221_X1 U10852 ( .B1(n9806), .B2(keyinput22), .C1(n9805), .C2(keyinput37), 
        .A(n9804), .ZN(n9812) );
  AOI22_X1 U10853 ( .A1(n5350), .A2(keyinput0), .B1(n9808), .B2(keyinput56), 
        .ZN(n9807) );
  OAI221_X1 U10854 ( .B1(n5350), .B2(keyinput0), .C1(n9808), .C2(keyinput56), 
        .A(n9807), .ZN(n9811) );
  AOI22_X1 U10855 ( .A1(n9895), .A2(keyinput28), .B1(n7738), .B2(keyinput44), 
        .ZN(n9809) );
  OAI221_X1 U10856 ( .B1(n9895), .B2(keyinput28), .C1(n7738), .C2(keyinput44), 
        .A(n9809), .ZN(n9810) );
  NOR4_X1 U10857 ( .A1(n9813), .A2(n9812), .A3(n9811), .A4(n9810), .ZN(n9826)
         );
  INV_X1 U10858 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9815) );
  AOI22_X1 U10859 ( .A1(n9815), .A2(keyinput59), .B1(n9890), .B2(keyinput14), 
        .ZN(n9814) );
  OAI221_X1 U10860 ( .B1(n9815), .B2(keyinput59), .C1(n9890), .C2(keyinput14), 
        .A(n9814), .ZN(n9824) );
  AOI22_X1 U10861 ( .A1(n5344), .A2(keyinput15), .B1(n6573), .B2(keyinput43), 
        .ZN(n9816) );
  OAI221_X1 U10862 ( .B1(n5344), .B2(keyinput15), .C1(n6573), .C2(keyinput43), 
        .A(n9816), .ZN(n9823) );
  INV_X1 U10863 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9818) );
  AOI22_X1 U10864 ( .A1(n7232), .A2(keyinput25), .B1(keyinput41), .B2(n9818), 
        .ZN(n9817) );
  OAI221_X1 U10865 ( .B1(n7232), .B2(keyinput25), .C1(n9818), .C2(keyinput41), 
        .A(n9817), .ZN(n9822) );
  XNOR2_X1 U10866 ( .A(P1_REG1_REG_19__SCAN_IN), .B(keyinput45), .ZN(n9820) );
  XNOR2_X1 U10867 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput38), .ZN(n9819) );
  NAND2_X1 U10868 ( .A1(n9820), .A2(n9819), .ZN(n9821) );
  NOR4_X1 U10869 ( .A1(n9824), .A2(n9823), .A3(n9822), .A4(n9821), .ZN(n9825)
         );
  NAND4_X1 U10870 ( .A1(n9828), .A2(n9827), .A3(n9826), .A4(n9825), .ZN(n9886)
         );
  AOI22_X1 U10871 ( .A1(n9830), .A2(keyinput30), .B1(keyinput19), .B2(n5698), 
        .ZN(n9829) );
  OAI221_X1 U10872 ( .B1(n9830), .B2(keyinput30), .C1(n5698), .C2(keyinput19), 
        .A(n9829), .ZN(n9841) );
  AOI22_X1 U10873 ( .A1(n4830), .A2(keyinput47), .B1(n9832), .B2(keyinput31), 
        .ZN(n9831) );
  OAI221_X1 U10874 ( .B1(n4830), .B2(keyinput47), .C1(n9832), .C2(keyinput31), 
        .A(n9831), .ZN(n9840) );
  AOI22_X1 U10875 ( .A1(n9835), .A2(keyinput42), .B1(n9834), .B2(keyinput35), 
        .ZN(n9833) );
  OAI221_X1 U10876 ( .B1(n9835), .B2(keyinput42), .C1(n9834), .C2(keyinput35), 
        .A(n9833), .ZN(n9839) );
  XNOR2_X1 U10877 ( .A(P1_REG0_REG_14__SCAN_IN), .B(keyinput33), .ZN(n9837) );
  XNOR2_X1 U10878 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput60), .ZN(n9836) );
  NAND2_X1 U10879 ( .A1(n9837), .A2(n9836), .ZN(n9838) );
  NOR4_X1 U10880 ( .A1(n9841), .A2(n9840), .A3(n9839), .A4(n9838), .ZN(n9884)
         );
  AOI22_X1 U10881 ( .A1(n9843), .A2(keyinput16), .B1(keyinput50), .B2(n7109), 
        .ZN(n9842) );
  OAI221_X1 U10882 ( .B1(n9843), .B2(keyinput16), .C1(n7109), .C2(keyinput50), 
        .A(n9842), .ZN(n9853) );
  AOI22_X1 U10883 ( .A1(n9897), .A2(keyinput49), .B1(n9891), .B2(keyinput36), 
        .ZN(n9844) );
  OAI221_X1 U10884 ( .B1(n9897), .B2(keyinput49), .C1(n9891), .C2(keyinput36), 
        .A(n9844), .ZN(n9852) );
  INV_X1 U10885 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9847) );
  AOI22_X1 U10886 ( .A1(n9847), .A2(keyinput13), .B1(n9846), .B2(keyinput51), 
        .ZN(n9845) );
  OAI221_X1 U10887 ( .B1(n9847), .B2(keyinput13), .C1(n9846), .C2(keyinput51), 
        .A(n9845), .ZN(n9851) );
  XOR2_X1 U10888 ( .A(n5181), .B(keyinput7), .Z(n9849) );
  XNOR2_X1 U10889 ( .A(SI_2_), .B(keyinput27), .ZN(n9848) );
  NAND2_X1 U10890 ( .A1(n9849), .A2(n9848), .ZN(n9850) );
  NOR4_X1 U10891 ( .A1(n9853), .A2(n9852), .A3(n9851), .A4(n9850), .ZN(n9883)
         );
  AOI22_X1 U10892 ( .A1(n9856), .A2(keyinput4), .B1(keyinput10), .B2(n9855), 
        .ZN(n9854) );
  OAI221_X1 U10893 ( .B1(n9856), .B2(keyinput4), .C1(n9855), .C2(keyinput10), 
        .A(n9854), .ZN(n9866) );
  AOI22_X1 U10894 ( .A1(n9859), .A2(keyinput11), .B1(n9858), .B2(keyinput1), 
        .ZN(n9857) );
  OAI221_X1 U10895 ( .B1(n9859), .B2(keyinput11), .C1(n9858), .C2(keyinput1), 
        .A(n9857), .ZN(n9865) );
  XNOR2_X1 U10896 ( .A(P1_REG3_REG_10__SCAN_IN), .B(keyinput54), .ZN(n9863) );
  XNOR2_X1 U10897 ( .A(P2_IR_REG_29__SCAN_IN), .B(keyinput34), .ZN(n9862) );
  XNOR2_X1 U10898 ( .A(P2_IR_REG_5__SCAN_IN), .B(keyinput26), .ZN(n9861) );
  XNOR2_X1 U10899 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput62), .ZN(n9860) );
  NAND4_X1 U10900 ( .A1(n9863), .A2(n9862), .A3(n9861), .A4(n9860), .ZN(n9864)
         );
  NOR3_X1 U10901 ( .A1(n9866), .A2(n9865), .A3(n9864), .ZN(n9882) );
  AOI22_X1 U10902 ( .A1(n9869), .A2(keyinput3), .B1(keyinput12), .B2(n9868), 
        .ZN(n9867) );
  OAI221_X1 U10903 ( .B1(n9869), .B2(keyinput3), .C1(n9868), .C2(keyinput12), 
        .A(n9867), .ZN(n9880) );
  AOI22_X1 U10904 ( .A1(n9871), .A2(keyinput58), .B1(keyinput23), .B2(n9904), 
        .ZN(n9870) );
  OAI221_X1 U10905 ( .B1(n9871), .B2(keyinput58), .C1(n9904), .C2(keyinput23), 
        .A(n9870), .ZN(n9879) );
  INV_X1 U10906 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9874) );
  AOI22_X1 U10907 ( .A1(n9874), .A2(keyinput52), .B1(n9873), .B2(keyinput63), 
        .ZN(n9872) );
  OAI221_X1 U10908 ( .B1(n9874), .B2(keyinput52), .C1(n9873), .C2(keyinput63), 
        .A(n9872), .ZN(n9878) );
  XNOR2_X1 U10909 ( .A(P1_REG3_REG_1__SCAN_IN), .B(keyinput9), .ZN(n9876) );
  XNOR2_X1 U10910 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput40), .ZN(n9875)
         );
  NAND2_X1 U10911 ( .A1(n9876), .A2(n9875), .ZN(n9877) );
  NOR4_X1 U10912 ( .A1(n9880), .A2(n9879), .A3(n9878), .A4(n9877), .ZN(n9881)
         );
  NAND4_X1 U10913 ( .A1(n9884), .A2(n9883), .A3(n9882), .A4(n9881), .ZN(n9885)
         );
  NOR2_X1 U10914 ( .A1(n9886), .A2(n9885), .ZN(n9889) );
  NAND2_X1 U10915 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9887), .ZN(n9888) );
  XNOR2_X1 U10916 ( .A(n9889), .B(n9888), .ZN(n9918) );
  NAND4_X1 U10917 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9891), .A3(n9890), .A4(
        n6573), .ZN(n9894) );
  NAND4_X1 U10918 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), 
        .A3(P2_IR_REG_26__SCAN_IN), .A4(n9892), .ZN(n9893) );
  NOR4_X1 U10919 ( .A1(n9895), .A2(P2_IR_REG_5__SCAN_IN), .A3(n9894), .A4(
        n9893), .ZN(n9896) );
  NAND3_X1 U10920 ( .A1(n9896), .A2(P1_ADDR_REG_12__SCAN_IN), .A3(
        P1_ADDR_REG_14__SCAN_IN), .ZN(n9899) );
  NAND4_X1 U10921 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .A3(n5181), .A4(n9897), .ZN(n9898) );
  NOR2_X1 U10922 ( .A1(n9899), .A2(n9898), .ZN(n9916) );
  NOR4_X1 U10923 ( .A1(SI_2_), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_IR_REG_29__SCAN_IN), .A4(P2_REG0_REG_22__SCAN_IN), .ZN(n9903) );
  NOR4_X1 U10924 ( .A1(P1_D_REG_26__SCAN_IN), .A2(SI_12_), .A3(
        P2_REG1_REG_9__SCAN_IN), .A4(P2_REG1_REG_1__SCAN_IN), .ZN(n9902) );
  NOR4_X1 U10925 ( .A1(P1_RD_REG_SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), .A3(
        P1_REG0_REG_9__SCAN_IN), .A4(SI_29_), .ZN(n9901) );
  NOR4_X1 U10926 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_REG1_REG_19__SCAN_IN), 
        .A3(P2_REG3_REG_16__SCAN_IN), .A4(P2_REG2_REG_21__SCAN_IN), .ZN(n9900)
         );
  AND4_X1 U10927 ( .A1(n9903), .A2(n9902), .A3(n9901), .A4(n9900), .ZN(n9915)
         );
  NAND4_X1 U10928 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(
        P2_DATAO_REG_25__SCAN_IN), .A3(SI_8_), .A4(n9904), .ZN(n9908) );
  NAND4_X1 U10929 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(P1_DATAO_REG_9__SCAN_IN), .A3(P2_REG3_REG_18__SCAN_IN), .A4(P2_REG3_REG_10__SCAN_IN), .ZN(n9907) );
  NAND4_X1 U10930 ( .A1(SI_11_), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_REG3_REG_8__SCAN_IN), .A4(P2_REG1_REG_4__SCAN_IN), .ZN(n9906) );
  NAND4_X1 U10931 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG2_REG_11__SCAN_IN), .A4(P2_REG3_REG_0__SCAN_IN), .ZN(n9905)
         );
  NOR4_X1 U10932 ( .A1(n9908), .A2(n9907), .A3(n9906), .A4(n9905), .ZN(n9914)
         );
  NAND4_X1 U10933 ( .A1(P1_REG1_REG_27__SCAN_IN), .A2(P1_REG0_REG_25__SCAN_IN), 
        .A3(P1_REG0_REG_24__SCAN_IN), .A4(P1_REG1_REG_31__SCAN_IN), .ZN(n9912)
         );
  NAND4_X1 U10934 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .A3(SI_20_), .A4(P1_REG1_REG_9__SCAN_IN), .ZN(n9911) );
  NAND4_X1 U10935 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_REG0_REG_14__SCAN_IN), 
        .A3(P1_REG3_REG_1__SCAN_IN), .A4(P1_REG2_REG_18__SCAN_IN), .ZN(n9910)
         );
  NAND4_X1 U10936 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG2_REG_26__SCAN_IN), 
        .A3(P1_REG0_REG_16__SCAN_IN), .A4(P2_REG0_REG_14__SCAN_IN), .ZN(n9909)
         );
  NOR4_X1 U10937 ( .A1(n9912), .A2(n9911), .A3(n9910), .A4(n9909), .ZN(n9913)
         );
  NAND4_X1 U10938 ( .A1(n9916), .A2(n9915), .A3(n9914), .A4(n9913), .ZN(n9917)
         );
  XNOR2_X1 U10939 ( .A(n9918), .B(n9917), .ZN(P2_U3319) );
  XOR2_X1 U10940 ( .A(n9919), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  XOR2_X1 U10941 ( .A(n9920), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  XOR2_X1 U10942 ( .A(n9921), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1071_U48) );
  NOR2_X1 U10943 ( .A1(n9923), .A2(n9922), .ZN(n9924) );
  XOR2_X1 U10944 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n9924), .Z(ADD_1071_U51) );
  OAI21_X1 U10945 ( .B1(n9927), .B2(n9926), .A(n9925), .ZN(n9928) );
  XNOR2_X1 U10946 ( .A(n9928), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U10947 ( .B1(n5350), .B2(n9930), .A(n9929), .ZN(ADD_1071_U47) );
  XOR2_X1 U10948 ( .A(n9932), .B(n9931), .Z(ADD_1071_U54) );
  XOR2_X1 U10949 ( .A(n9934), .B(n9933), .Z(ADD_1071_U53) );
  XNOR2_X1 U10950 ( .A(n9936), .B(n9935), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U5142 ( .A(n5669), .Z(n6976) );
endmodule

