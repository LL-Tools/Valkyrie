

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput63, keyinput62, keyinput61, keyinput60, keyinput59, 
        keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, keyinput53, 
        keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, keyinput47, 
        keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, keyinput41, 
        keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, keyinput35, 
        keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, keyinput29, 
        keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, keyinput23, 
        keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, keyinput17, 
        keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, keyinput11, 
        keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5, 
        keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670;

  CLKBUF_X2 U2246 ( .A(n3550), .Z(n3546) );
  CLKBUF_X2 U2247 ( .A(n2913), .Z(n2005) );
  CLKBUF_X2 U2248 ( .A(n2958), .Z(n3538) );
  CLKBUF_X2 U2249 ( .A(n2952), .Z(n3550) );
  INV_X1 U2250 ( .A(n2611), .ZN(n2838) );
  NAND2_X1 U2251 ( .A1(n2737), .A2(n2736), .ZN(n2739) );
  AND2_X1 U2252 ( .A1(n3577), .A2(n3511), .ZN(n3524) );
  INV_X1 U2253 ( .A(n2585), .ZN(n2641) );
  INV_X2 U2254 ( .A(n2369), .ZN(n2352) );
  INV_X1 U2255 ( .A(n4453), .ZN(n4211) );
  NAND2_X1 U2256 ( .A1(n2299), .A2(n2298), .ZN(n2379) );
  NAND2_X1 U2257 ( .A1(n2032), .A2(IR_REG_31__SCAN_IN), .ZN(n2140) );
  INV_X1 U2259 ( .A(n4458), .ZN(n4136) );
  INV_X4 U2260 ( .A(n2354), .ZN(n2370) );
  INV_X1 U2261 ( .A(n2005), .ZN(n2004) );
  AND2_X1 U2262 ( .A1(n3495), .A2(n4510), .ZN(n2913) );
  NAND2_X4 U2263 ( .A1(n2857), .A2(n2856), .ZN(n3547) );
  OAI21_X2 U2264 ( .B1(n2811), .B2(n2769), .A(n2771), .ZN(n3912) );
  XNOR2_X2 U2265 ( .A(n2739), .B(n2779), .ZN(n2778) );
  XNOR2_X2 U2266 ( .A(n2140), .B(n2350), .ZN(n3897) );
  OAI21_X1 U2267 ( .B1(n4377), .B2(n2129), .A(n2128), .ZN(n4385) );
  NAND2_X1 U2268 ( .A1(n2820), .A2(n2688), .ZN(n4510) );
  NAND2_X1 U2269 ( .A1(n2665), .A2(n2664), .ZN(n2787) );
  AND2_X1 U2270 ( .A1(n3858), .A2(n2647), .ZN(n2820) );
  XNOR2_X1 U2271 ( .A(n2658), .B(IR_REG_24__SCAN_IN), .ZN(n2665) );
  NAND4_X1 U2272 ( .A1(n2340), .A2(n2339), .A3(n2338), .A4(n2337), .ZN(n3884)
         );
  NAND2_X1 U2273 ( .A1(n2688), .A2(n2636), .ZN(n2857) );
  NAND2_X1 U2274 ( .A1(n2657), .A2(IR_REG_31__SCAN_IN), .ZN(n2658) );
  NAND4_X2 U2275 ( .A1(n2358), .A2(n2357), .A3(n2356), .A4(n2355), .ZN(n3881)
         );
  NAND4_X2 U2276 ( .A1(n2142), .A2(n2329), .A3(n2331), .A4(n2330), .ZN(n2854)
         );
  XNOR2_X1 U2277 ( .A(n2609), .B(IR_REG_22__SCAN_IN), .ZN(n4328) );
  INV_X2 U2278 ( .A(n2704), .ZN(n2549) );
  NAND2_X1 U2279 ( .A1(n2291), .A2(n2289), .ZN(n2369) );
  NAND2_X1 U2280 ( .A1(n2604), .A2(IR_REG_31__SCAN_IN), .ZN(n2599) );
  NAND2_X2 U2281 ( .A1(n2291), .A2(n4324), .ZN(n2371) );
  AND2_X1 U2282 ( .A1(n2188), .A2(n2324), .ZN(n2651) );
  NAND2_X1 U2283 ( .A1(n2715), .A2(n2714), .ZN(n3899) );
  INV_X1 U2284 ( .A(IR_REG_4__SCAN_IN), .ZN(n2377) );
  INV_X1 U2285 ( .A(IR_REG_2__SCAN_IN), .ZN(n2350) );
  NOR2_X1 U2286 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2065)
         );
  NOR2_X1 U2287 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2066)
         );
  NOR2_X1 U2288 ( .A1(IR_REG_5__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2067)
         );
  NOR2_X1 U2289 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2068)
         );
  NOR2_X2 U2290 ( .A1(n3915), .A2(n4355), .ZN(n4367) );
  NOR3_X2 U2291 ( .A1(n3658), .A2(n3575), .A3(n3574), .ZN(n3508) );
  NAND2_X1 U2292 ( .A1(n2186), .A2(n4107), .ZN(n2184) );
  INV_X1 U2293 ( .A(n3722), .ZN(n2081) );
  NOR2_X1 U2294 ( .A1(n2228), .A2(n3607), .ZN(n2227) );
  INV_X1 U2295 ( .A(n3677), .ZN(n2228) );
  INV_X1 U2296 ( .A(n4324), .ZN(n2289) );
  NAND2_X1 U2297 ( .A1(n4131), .A2(n4160), .ZN(n2536) );
  INV_X1 U2298 ( .A(n2857), .ZN(n3026) );
  INV_X1 U2299 ( .A(n2830), .ZN(n2705) );
  NAND2_X1 U2300 ( .A1(n2711), .A2(IR_REG_28__SCAN_IN), .ZN(n2298) );
  AND2_X1 U2301 ( .A1(n2829), .A2(n3023), .ZN(n2851) );
  INV_X1 U2302 ( .A(n2371), .ZN(n2594) );
  NAND2_X1 U2303 ( .A1(n4325), .A2(n2289), .ZN(n2354) );
  NAND2_X1 U2304 ( .A1(n2290), .A2(n2288), .ZN(n2291) );
  XNOR2_X1 U2305 ( .A(n2122), .B(n4468), .ZN(n4400) );
  INV_X1 U2306 ( .A(n3938), .ZN(n2122) );
  OR2_X1 U2307 ( .A1(n3986), .A2(n3985), .ZN(n4225) );
  AND2_X1 U2308 ( .A1(n2571), .A2(n2563), .ZN(n4059) );
  AND2_X1 U2309 ( .A1(n2184), .A2(n2042), .ZN(n2180) );
  INV_X1 U2310 ( .A(n2187), .ZN(n2181) );
  NOR2_X1 U2311 ( .A1(n2186), .A2(n4107), .ZN(n2185) );
  INV_X1 U2312 ( .A(n4154), .ZN(n4108) );
  AND2_X1 U2313 ( .A1(n2820), .A2(n4330), .ZN(n4227) );
  AND2_X1 U2314 ( .A1(n2651), .A2(n2007), .ZN(n2294) );
  NAND2_X1 U2315 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2332)
         );
  AOI21_X1 U2316 ( .B1(n2241), .B2(n3223), .A(n2240), .ZN(n2239) );
  INV_X1 U2317 ( .A(n3243), .ZN(n2240) );
  AOI21_X1 U2318 ( .B1(n3223), .B2(n3208), .A(n2242), .ZN(n2238) );
  NOR2_X1 U2319 ( .A1(n2800), .A2(n2115), .ZN(n2114) );
  INV_X1 U2320 ( .A(n2379), .ZN(n2704) );
  INV_X1 U2321 ( .A(n3792), .ZN(n2076) );
  NAND2_X1 U2322 ( .A1(n4054), .A2(n2686), .ZN(n2173) );
  NAND2_X1 U2323 ( .A1(n2081), .A2(n2079), .ZN(n2078) );
  INV_X1 U2324 ( .A(n3790), .ZN(n2079) );
  NAND2_X1 U2325 ( .A1(n2631), .A2(n2025), .ZN(n2077) );
  INV_X1 U2326 ( .A(n2513), .ZN(n2146) );
  INV_X1 U2327 ( .A(n2502), .ZN(n2145) );
  AND2_X1 U2328 ( .A1(n3430), .A2(n3459), .ZN(n2512) );
  NAND2_X1 U2329 ( .A1(n3328), .A2(n2148), .ZN(n2147) );
  AOI21_X1 U2330 ( .B1(n3838), .B2(n2474), .A(n2028), .ZN(n2162) );
  INV_X1 U2331 ( .A(n2474), .ZN(n2160) );
  NAND2_X1 U2332 ( .A1(n3091), .A2(n3769), .ZN(n2097) );
  NOR2_X1 U2333 ( .A1(n2446), .A2(n2153), .ZN(n2152) );
  INV_X1 U2334 ( .A(n2155), .ZN(n2153) );
  OR2_X1 U2335 ( .A1(n3099), .A2(n2451), .ZN(n2446) );
  NAND2_X1 U2336 ( .A1(n2395), .A2(n2157), .ZN(n2154) );
  NOR2_X1 U2337 ( .A1(n2408), .A2(n2158), .ZN(n2157) );
  INV_X1 U2338 ( .A(n2394), .ZN(n2158) );
  OR2_X1 U2339 ( .A1(n3878), .A2(n3151), .ZN(n3763) );
  NAND2_X1 U2340 ( .A1(n3763), .A2(n3765), .ZN(n3125) );
  OR2_X1 U2341 ( .A1(n3882), .A2(n2899), .ZN(n3748) );
  NAND2_X1 U2342 ( .A1(n4208), .A2(n4137), .ZN(n2106) );
  OR2_X1 U2343 ( .A1(n3423), .A2(n3617), .ZN(n3422) );
  INV_X1 U2344 ( .A(IR_REG_26__SCAN_IN), .ZN(n2254) );
  INV_X1 U2345 ( .A(n2294), .ZN(n2662) );
  INV_X1 U2346 ( .A(IR_REG_25__SCAN_IN), .ZN(n4654) );
  INV_X1 U2347 ( .A(n2227), .ZN(n2226) );
  NAND2_X1 U2348 ( .A1(n2227), .A2(n2225), .ZN(n2224) );
  AOI22_X1 U2349 ( .A1(n2239), .A2(n2235), .B1(n2238), .B2(n2234), .ZN(n2233)
         );
  INV_X1 U2350 ( .A(n3208), .ZN(n2234) );
  INV_X1 U2351 ( .A(n2241), .ZN(n2235) );
  INV_X1 U2352 ( .A(n2248), .ZN(n2246) );
  OAI21_X1 U2353 ( .B1(n3615), .B2(n2249), .A(n3462), .ZN(n2248) );
  NAND2_X1 U2354 ( .A1(n3458), .A2(n2252), .ZN(n2249) );
  NAND2_X1 U2355 ( .A1(n2250), .A2(n2245), .ZN(n2244) );
  INV_X1 U2356 ( .A(n3445), .ZN(n2245) );
  NOR2_X1 U2357 ( .A1(n3615), .A2(n2251), .ZN(n2250) );
  NOR2_X1 U2358 ( .A1(n3458), .A2(n2252), .ZN(n2251) );
  NOR2_X1 U2359 ( .A1(n3509), .A2(n3510), .ZN(n3511) );
  NAND2_X1 U2360 ( .A1(n2914), .A2(n2917), .ZN(n2919) );
  XNOR2_X1 U2361 ( .A(n2905), .B(n3533), .ZN(n2943) );
  NAND2_X1 U2362 ( .A1(n2208), .A2(n3002), .ZN(n2207) );
  INV_X1 U2363 ( .A(n2997), .ZN(n2208) );
  AOI22_X1 U2364 ( .A1(n2791), .A2(IR_REG_0__SCAN_IN), .B1(n3062), .B2(n2902), 
        .ZN(n2792) );
  NOR2_X1 U2365 ( .A1(n2239), .A2(n2238), .ZN(n2236) );
  AOI21_X1 U2366 ( .B1(n2200), .B2(n2199), .A(n2198), .ZN(n2197) );
  INV_X1 U2367 ( .A(n3594), .ZN(n2198) );
  INV_X1 U2368 ( .A(n4328), .ZN(n3858) );
  OR2_X1 U2369 ( .A1(n2354), .A2(n2716), .ZN(n2329) );
  NAND2_X1 U2370 ( .A1(n2370), .A2(REG1_REG_0__SCAN_IN), .ZN(n2337) );
  XNOR2_X1 U2371 ( .A(n2732), .B(n2731), .ZN(n2782) );
  OAI21_X1 U2372 ( .B1(n2778), .B2(n2738), .A(n2740), .ZN(n2803) );
  NAND2_X1 U2373 ( .A1(n2132), .A2(REG1_REG_12__SCAN_IN), .ZN(n2129) );
  INV_X1 U2374 ( .A(n4386), .ZN(n2132) );
  OR2_X1 U2375 ( .A1(n4377), .A2(n4378), .ZN(n2131) );
  NAND2_X1 U2376 ( .A1(n4370), .A2(n3932), .ZN(n3934) );
  NAND2_X1 U2377 ( .A1(n2124), .A2(REG2_REG_14__SCAN_IN), .ZN(n2126) );
  INV_X1 U2378 ( .A(n4400), .ZN(n2124) );
  XNOR2_X1 U2379 ( .A(n3957), .B(n2108), .ZN(n3941) );
  INV_X1 U2380 ( .A(n3956), .ZN(n2108) );
  NAND2_X1 U2381 ( .A1(n3941), .A2(n3424), .ZN(n3958) );
  NAND2_X1 U2382 ( .A1(n4419), .A2(n2139), .ZN(n2138) );
  OR2_X1 U2383 ( .A1(n3960), .A2(REG1_REG_17__SCAN_IN), .ZN(n2139) );
  NOR2_X1 U2384 ( .A1(n2138), .A2(n4432), .ZN(n4431) );
  NAND2_X1 U2385 ( .A1(n2379), .A2(DATAI_27_), .ZN(n3998) );
  OAI22_X1 U2386 ( .A1(n4047), .A2(n2569), .B1(n3441), .B2(n4073), .ZN(n4029)
         );
  NAND2_X1 U2387 ( .A1(n2551), .A2(REG3_REG_23__SCAN_IN), .ZN(n2562) );
  NAND2_X1 U2388 ( .A1(n2174), .A2(n2176), .ZN(n4094) );
  AND2_X1 U2389 ( .A1(n4095), .A2(n2177), .ZN(n2176) );
  NAND2_X1 U2390 ( .A1(n2178), .A2(n2179), .ZN(n2177) );
  OR2_X1 U2391 ( .A1(n4108), .A2(n4137), .ZN(n2187) );
  OR2_X1 U2392 ( .A1(n2514), .A2(n3639), .ZN(n2516) );
  NAND2_X1 U2393 ( .A1(n2501), .A2(n3390), .ZN(n2502) );
  INV_X1 U2394 ( .A(n3871), .ZN(n2501) );
  OR2_X1 U2395 ( .A1(n2489), .A2(n2147), .ZN(n3327) );
  NAND2_X1 U2396 ( .A1(n2163), .A2(n3264), .ZN(n3263) );
  AND2_X1 U2397 ( .A1(n2828), .A2(n2827), .ZN(n3023) );
  AND2_X1 U2398 ( .A1(n2089), .A2(n2088), .ZN(n4232) );
  INV_X1 U2399 ( .A(n3983), .ZN(n2088) );
  NAND2_X1 U2400 ( .A1(n2090), .A2(n4196), .ZN(n2089) );
  NAND2_X1 U2401 ( .A1(n2549), .A2(DATAI_20_), .ZN(n4137) );
  AND3_X1 U2402 ( .A1(n2680), .A2(n2679), .A3(n2678), .ZN(n2690) );
  AND2_X1 U2403 ( .A1(n2931), .A2(n4461), .ZN(n2836) );
  AND2_X1 U2404 ( .A1(n2286), .A2(n2283), .ZN(n2287) );
  AND2_X1 U2405 ( .A1(n2285), .A2(n2297), .ZN(n2286) );
  INV_X1 U2406 ( .A(IR_REG_29__SCAN_IN), .ZN(n2285) );
  MUX2_X1 U2407 ( .A(IR_REG_31__SCAN_IN), .B(n2284), .S(IR_REG_29__SCAN_IN), 
        .Z(n2290) );
  AND2_X1 U2408 ( .A1(n2022), .A2(n2189), .ZN(n2188) );
  XNOR2_X1 U2409 ( .A(n2666), .B(n2667), .ZN(n2930) );
  INV_X1 U2410 ( .A(IR_REG_16__SCAN_IN), .ZN(n2317) );
  INV_X1 U2411 ( .A(n3882), .ZN(n3173) );
  INV_X1 U2412 ( .A(n4059), .ZN(n2064) );
  NAND2_X1 U2413 ( .A1(n3583), .A2(n3482), .ZN(n3648) );
  NAND2_X1 U2414 ( .A1(n2588), .A2(n2014), .ZN(n4019) );
  OR2_X1 U2415 ( .A1(n2544), .A2(n2543), .ZN(n4154) );
  NAND2_X1 U2416 ( .A1(n2542), .A2(n2044), .ZN(n2543) );
  AND2_X1 U2417 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n2714)
         );
  XNOR2_X1 U2418 ( .A(n3934), .B(n4472), .ZN(n4382) );
  NAND2_X1 U2419 ( .A1(n4382), .A2(REG2_REG_12__SCAN_IN), .ZN(n4381) );
  INV_X1 U2420 ( .A(n4470), .ZN(n4394) );
  OR2_X1 U2421 ( .A1(n4413), .A2(n3337), .ZN(n2123) );
  NAND2_X1 U2422 ( .A1(n3939), .A2(n2127), .ZN(n2121) );
  NAND2_X1 U2423 ( .A1(n4423), .A2(n4424), .ZN(n4422) );
  INV_X1 U2424 ( .A(n4431), .ZN(n2137) );
  AOI21_X1 U2425 ( .B1(n2138), .B2(n4432), .A(n4430), .ZN(n2136) );
  INV_X1 U2426 ( .A(n2135), .ZN(n2134) );
  AOI21_X1 U2427 ( .B1(n4434), .B2(ADDR_REG_18__SCAN_IN), .A(n4433), .ZN(n2135) );
  AND2_X1 U2428 ( .A1(n2749), .A2(n3857), .ZN(n4439) );
  NAND2_X1 U2429 ( .A1(n4225), .A2(n2107), .ZN(n4231) );
  OR2_X1 U2430 ( .A1(n3988), .A2(n3987), .ZN(n2107) );
  NAND2_X1 U2431 ( .A1(n2294), .A2(n2287), .ZN(n2288) );
  AND2_X1 U2432 ( .A1(n3208), .A2(n2242), .ZN(n2241) );
  INV_X1 U2433 ( .A(n3693), .ZN(n2252) );
  OAI21_X1 U2434 ( .B1(n3447), .B2(n3446), .A(n3445), .ZN(n2253) );
  AOI21_X1 U2435 ( .B1(REG2_REG_2__SCAN_IN), .B2(n4335), .A(n3903), .ZN(n2729)
         );
  NOR2_X1 U2436 ( .A1(n4407), .A2(n3921), .ZN(n3949) );
  NAND2_X1 U2437 ( .A1(n2582), .A2(n2171), .ZN(n2169) );
  OR2_X1 U2438 ( .A1(n3744), .A2(n3998), .ZN(n2170) );
  INV_X1 U2439 ( .A(n2173), .ZN(n2165) );
  NAND2_X1 U2440 ( .A1(n2077), .A2(n2074), .ZN(n4031) );
  OR2_X1 U2441 ( .A1(n2562), .A2(n3444), .ZN(n2571) );
  INV_X1 U2442 ( .A(n2180), .ZN(n2178) );
  AND2_X1 U2443 ( .A1(n2630), .A2(n2629), .ZN(n3786) );
  NAND2_X1 U2444 ( .A1(n4193), .A2(n3718), .ZN(n4147) );
  NAND2_X1 U2445 ( .A1(n2962), .A2(n2156), .ZN(n2155) );
  INV_X1 U2446 ( .A(n3879), .ZN(n2156) );
  AND2_X1 U2447 ( .A1(n2342), .A2(n2366), .ZN(n2150) );
  INV_X1 U2448 ( .A(n3753), .ZN(n2083) );
  NAND2_X1 U2449 ( .A1(n2891), .A2(n3835), .ZN(n2890) );
  XNOR2_X1 U2450 ( .A(n3978), .B(n2091), .ZN(n2090) );
  INV_X1 U2451 ( .A(n3979), .ZN(n2091) );
  NOR2_X1 U2452 ( .A1(n2686), .A2(n3441), .ZN(n2099) );
  NAND2_X1 U2453 ( .A1(n3273), .A2(n3297), .ZN(n2102) );
  XNOR2_X1 U2454 ( .A(n2603), .B(IR_REG_21__SCAN_IN), .ZN(n2636) );
  AND2_X1 U2455 ( .A1(n2599), .A2(n2602), .ZN(n2603) );
  INV_X1 U2456 ( .A(IR_REG_19__SCAN_IN), .ZN(n2606) );
  NAND2_X1 U2457 ( .A1(n2300), .A2(n2261), .ZN(n2522) );
  INV_X1 U2458 ( .A(n2314), .ZN(n2300) );
  NOR2_X1 U2459 ( .A1(IR_REG_13__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2189)
         );
  INV_X1 U2460 ( .A(IR_REG_10__SCAN_IN), .ZN(n4655) );
  INV_X1 U2461 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4601) );
  INV_X1 U2462 ( .A(n2019), .ZN(n2216) );
  AOI21_X1 U2463 ( .B1(n2221), .B2(n2226), .A(n2029), .ZN(n2217) );
  INV_X1 U2464 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3444) );
  NAND2_X1 U2465 ( .A1(n2274), .A2(REG3_REG_19__SCAN_IN), .ZN(n2538) );
  OR2_X1 U2466 ( .A1(n2538), .A2(n3651), .ZN(n2540) );
  INV_X1 U2467 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3651) );
  INV_X1 U2468 ( .A(n3358), .ZN(n3351) );
  NOR2_X1 U2469 ( .A1(n2253), .A2(n3458), .ZN(n3690) );
  NAND2_X1 U2470 ( .A1(n2253), .A2(n3458), .ZN(n3691) );
  AND2_X1 U2471 ( .A1(n2598), .A2(n2016), .ZN(n3982) );
  OR2_X1 U2472 ( .A1(n3560), .A2(n2641), .ZN(n2598) );
  NOR2_X1 U2473 ( .A1(n2050), .A2(n2070), .ZN(n2069) );
  NOR2_X1 U2474 ( .A1(n2354), .A2(n4546), .ZN(n2070) );
  NAND2_X1 U2475 ( .A1(n2370), .A2(REG1_REG_14__SCAN_IN), .ZN(n2495) );
  NAND2_X1 U2476 ( .A1(n2370), .A2(REG1_REG_13__SCAN_IN), .ZN(n2322) );
  AND2_X1 U2477 ( .A1(n3888), .A2(n2038), .ZN(n3885) );
  AOI21_X1 U2478 ( .B1(n4336), .B2(REG2_REG_1__SCAN_IN), .A(n3885), .ZN(n3905)
         );
  CLKBUF_X1 U2479 ( .A(n2359), .Z(n2360) );
  NOR2_X1 U2480 ( .A1(n2113), .A2(n2116), .ZN(n2760) );
  OAI21_X1 U2481 ( .B1(n2120), .B2(n2800), .A(n2030), .ZN(n2116) );
  AND2_X1 U2482 ( .A1(n2782), .A2(n2114), .ZN(n2113) );
  NAND2_X1 U2483 ( .A1(n4350), .A2(n2109), .ZN(n3930) );
  NAND2_X1 U2484 ( .A1(n3925), .A2(REG2_REG_9__SCAN_IN), .ZN(n2109) );
  NOR2_X1 U2485 ( .A1(n4345), .A2(n2047), .ZN(n3914) );
  NOR2_X1 U2486 ( .A1(n3919), .A2(n4395), .ZN(n4409) );
  AND2_X1 U2487 ( .A1(n2710), .A2(n2709), .ZN(n2749) );
  NOR2_X1 U2488 ( .A1(n4225), .A2(n4228), .ZN(n4224) );
  OAI21_X1 U2489 ( .B1(n4029), .B2(n2166), .A(n2164), .ZN(n3972) );
  INV_X1 U2490 ( .A(n2167), .ZN(n2166) );
  AOI21_X1 U2491 ( .B1(n2167), .B2(n2165), .A(n2168), .ZN(n2164) );
  AOI21_X1 U2492 ( .B1(n2173), .B2(n2043), .A(n2009), .ZN(n2167) );
  NAND2_X1 U2493 ( .A1(n2080), .A2(n2635), .ZN(n3996) );
  NAND2_X1 U2494 ( .A1(n2077), .A2(n2073), .ZN(n2080) );
  NOR2_X1 U2495 ( .A1(n3791), .A2(n2075), .ZN(n2073) );
  NAND2_X1 U2496 ( .A1(n2077), .A2(n2078), .ZN(n4050) );
  OR2_X1 U2497 ( .A1(n2545), .A2(n3661), .ZN(n2553) );
  AND2_X1 U2498 ( .A1(n2559), .A2(n2558), .ZN(n4091) );
  NAND2_X1 U2499 ( .A1(n2631), .A2(n3786), .ZN(n4105) );
  INV_X1 U2500 ( .A(n2505), .ZN(n2272) );
  NAND2_X1 U2501 ( .A1(n3426), .A2(n3828), .ZN(n4193) );
  NAND2_X1 U2502 ( .A1(n3406), .A2(n3713), .ZN(n3426) );
  INV_X1 U2503 ( .A(n2143), .ZN(n3421) );
  NOR2_X1 U2504 ( .A1(n2512), .A2(n2026), .ZN(n2144) );
  OR2_X1 U2505 ( .A1(n2503), .A2(n3695), .ZN(n2505) );
  OR2_X1 U2506 ( .A1(n3408), .A2(n3822), .ZN(n3406) );
  AOI21_X1 U2507 ( .B1(n2162), .B2(n2160), .A(n2027), .ZN(n2159) );
  INV_X1 U2508 ( .A(n2162), .ZN(n2161) );
  OR2_X1 U2509 ( .A1(n2478), .A2(n3314), .ZN(n2491) );
  AOI21_X1 U2510 ( .B1(n2095), .B2(n2094), .A(n2093), .ZN(n2092) );
  INV_X1 U2511 ( .A(n3769), .ZN(n2094) );
  AND2_X1 U2512 ( .A1(n2151), .A2(n2034), .ZN(n3238) );
  NAND2_X1 U2513 ( .A1(n3125), .A2(n2431), .ZN(n3099) );
  NAND2_X1 U2514 ( .A1(n3150), .A2(n3763), .ZN(n2616) );
  AND2_X1 U2515 ( .A1(n2072), .A2(n2071), .ZN(n3150) );
  NAND2_X1 U2516 ( .A1(n3048), .A2(n3045), .ZN(n2072) );
  INV_X1 U2517 ( .A(n3125), .ZN(n3837) );
  OAI21_X1 U2518 ( .B1(n3113), .B2(n3112), .A(n3760), .ZN(n3048) );
  AND2_X1 U2519 ( .A1(n3177), .A2(n3037), .ZN(n3121) );
  OAI21_X1 U2520 ( .B1(n2890), .B2(n2085), .A(n2082), .ZN(n3029) );
  AOI21_X1 U2521 ( .B1(n2264), .B2(n2084), .A(n2083), .ZN(n2082) );
  INV_X1 U2522 ( .A(n2264), .ZN(n2085) );
  INV_X1 U2523 ( .A(n3748), .ZN(n2084) );
  INV_X1 U2524 ( .A(n4090), .ZN(n4200) );
  AND2_X1 U2525 ( .A1(n3753), .A2(n3750), .ZN(n2264) );
  NAND2_X1 U2526 ( .A1(n2890), .A2(n3748), .ZN(n3171) );
  NAND2_X1 U2527 ( .A1(n2610), .A2(n2838), .ZN(n4135) );
  NAND2_X1 U2528 ( .A1(n3748), .A2(n3751), .ZN(n2888) );
  AND2_X1 U2529 ( .A1(n3069), .A2(n2342), .ZN(n2889) );
  INV_X1 U2530 ( .A(n4227), .ZN(n4198) );
  NOR2_X1 U2531 ( .A1(n4484), .A2(n4329), .ZN(n2835) );
  INV_X1 U2532 ( .A(n4219), .ZN(n4228) );
  AND2_X1 U2533 ( .A1(n4076), .A2(n2058), .ZN(n4004) );
  NAND2_X1 U2534 ( .A1(n4076), .A2(n2099), .ZN(n4039) );
  NAND2_X1 U2535 ( .A1(n4076), .A2(n4058), .ZN(n4057) );
  NOR2_X1 U2536 ( .A1(n4253), .A2(n3578), .ZN(n4076) );
  NAND2_X1 U2537 ( .A1(n2549), .A2(DATAI_23_), .ZN(n4078) );
  INV_X1 U2538 ( .A(n2106), .ZN(n2105) );
  INV_X1 U2539 ( .A(n2048), .ZN(n2104) );
  INV_X1 U2540 ( .A(n4181), .ZN(n4161) );
  NOR3_X1 U2541 ( .A1(n3422), .A2(n2048), .A3(n3641), .ZN(n4163) );
  NOR2_X1 U2542 ( .A1(n3422), .A2(n3641), .ZN(n4206) );
  NOR3_X1 U2543 ( .A1(n3271), .A2(n2100), .A3(n2102), .ZN(n3413) );
  OR2_X1 U2544 ( .A1(n3351), .A2(n3399), .ZN(n2100) );
  NOR2_X1 U2545 ( .A1(n3271), .A2(n3216), .ZN(n3298) );
  OR2_X1 U2546 ( .A1(n3105), .A2(n3085), .ZN(n3234) );
  OR2_X1 U2547 ( .A1(n3234), .A2(n3233), .ZN(n3271) );
  NOR2_X1 U2548 ( .A1(n3157), .A2(n3156), .ZN(n3160) );
  NAND2_X1 U2549 ( .A1(n3121), .A2(n3120), .ZN(n3119) );
  NAND2_X1 U2550 ( .A1(n2098), .A2(n2962), .ZN(n3157) );
  INV_X1 U2551 ( .A(n3119), .ZN(n2098) );
  INV_X1 U2552 ( .A(n4510), .ZN(n4489) );
  NAND2_X1 U2553 ( .A1(n2663), .A2(n4327), .ZN(n2826) );
  AND2_X1 U2554 ( .A1(IR_REG_27__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2296)
         );
  OR2_X1 U2555 ( .A1(n2294), .A2(n2349), .ZN(n2295) );
  NAND2_X1 U2556 ( .A1(n2662), .A2(n2661), .ZN(n2681) );
  INV_X1 U2557 ( .A(IR_REG_23__SCAN_IN), .ZN(n2667) );
  INV_X1 U2558 ( .A(n2636), .ZN(n2647) );
  INV_X1 U2559 ( .A(IR_REG_15__SCAN_IN), .ZN(n2315) );
  OR3_X1 U2560 ( .A1(n2441), .A2(IR_REG_7__SCAN_IN), .A3(IR_REG_8__SCAN_IN), 
        .ZN(n2443) );
  NOR2_X1 U2561 ( .A1(n2443), .A2(IR_REG_9__SCAN_IN), .ZN(n2470) );
  INV_X1 U2562 ( .A(IR_REG_7__SCAN_IN), .ZN(n2419) );
  INV_X1 U2563 ( .A(IR_REG_6__SCAN_IN), .ZN(n2417) );
  NAND2_X1 U2564 ( .A1(n2977), .A2(n2976), .ZN(n2998) );
  NAND2_X1 U2565 ( .A1(n2226), .A2(n2223), .ZN(n2218) );
  NOR2_X1 U2566 ( .A1(n2012), .A2(n2225), .ZN(n2220) );
  INV_X1 U2567 ( .A(n4078), .ZN(n3578) );
  INV_X1 U2568 ( .A(n3202), .ZN(n3233) );
  AND2_X1 U2569 ( .A1(n2019), .A2(n2221), .ZN(n2211) );
  OAI21_X1 U2570 ( .B1(n2019), .B2(n2217), .A(n2213), .ZN(n2212) );
  NAND2_X1 U2571 ( .A1(n2217), .A2(n2214), .ZN(n2213) );
  NAND2_X1 U2572 ( .A1(n2222), .A2(n2216), .ZN(n2214) );
  NAND2_X1 U2573 ( .A1(n2217), .A2(n2216), .ZN(n2215) );
  NAND2_X1 U2574 ( .A1(n2204), .A2(n3002), .ZN(n3080) );
  NAND2_X1 U2575 ( .A1(n2998), .A2(n2997), .ZN(n2204) );
  INV_X1 U2576 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3600) );
  INV_X1 U2577 ( .A(n3696), .ZN(n3683) );
  NAND2_X1 U2578 ( .A1(n3650), .A2(n3596), .ZN(n3599) );
  NAND2_X1 U2579 ( .A1(n2232), .A2(n2233), .ZN(n3308) );
  OR2_X1 U2580 ( .A1(n3222), .A2(n2236), .ZN(n2232) );
  INV_X1 U2581 ( .A(n4073), .ZN(n4034) );
  NAND3_X1 U2582 ( .A1(n2948), .A2(n2947), .A3(n2255), .ZN(n3626) );
  AOI21_X1 U2583 ( .B1(n2243), .B2(n2008), .A(n2031), .ZN(n3638) );
  INV_X1 U2584 ( .A(n2206), .ZN(n2205) );
  OAI21_X1 U2585 ( .B1(n3079), .B2(n2207), .A(n3078), .ZN(n2206) );
  AND2_X1 U2586 ( .A1(n2851), .A2(n2839), .ZN(n3696) );
  NAND2_X1 U2587 ( .A1(n2837), .A2(n4211), .ZN(n3640) );
  NAND2_X1 U2588 ( .A1(n3648), .A2(n3647), .ZN(n3650) );
  NAND2_X1 U2589 ( .A1(n2230), .A2(n2229), .ZN(n3384) );
  AOI21_X1 U2590 ( .B1(n2006), .B2(n2236), .A(n2231), .ZN(n2230) );
  INV_X1 U2591 ( .A(n3307), .ZN(n2231) );
  AND2_X1 U2592 ( .A1(n2195), .A2(n2197), .ZN(n2194) );
  INV_X1 U2593 ( .A(n3660), .ZN(n2195) );
  NAND2_X1 U2594 ( .A1(n2196), .A2(n2197), .ZN(n3659) );
  NAND2_X1 U2595 ( .A1(n2237), .A2(n3208), .ZN(n3245) );
  OR2_X1 U2596 ( .A1(n3222), .A2(n3223), .ZN(n2237) );
  OAI21_X1 U2597 ( .B1(n3638), .B2(n3634), .A(n3635), .ZN(n3671) );
  INV_X1 U2598 ( .A(n3697), .ZN(n3681) );
  INV_X1 U2599 ( .A(n3640), .ZN(n3680) );
  AND2_X1 U2600 ( .A1(n2583), .A2(n2579), .ZN(n4024) );
  INV_X1 U2601 ( .A(n3688), .ZN(n3704) );
  NAND2_X1 U2602 ( .A1(n2370), .A2(REG1_REG_31__SCAN_IN), .ZN(n3708) );
  NAND2_X1 U2603 ( .A1(n2370), .A2(REG1_REG_30__SCAN_IN), .ZN(n2725) );
  INV_X1 U2604 ( .A(n3982), .ZN(n4001) );
  INV_X1 U2605 ( .A(n4091), .ZN(n3867) );
  NAND2_X1 U2606 ( .A1(n2370), .A2(REG1_REG_19__SCAN_IN), .ZN(n2530) );
  NAND2_X1 U2607 ( .A1(n2370), .A2(REG1_REG_18__SCAN_IN), .ZN(n2306) );
  NAND2_X1 U2608 ( .A1(n2370), .A2(REG1_REG_17__SCAN_IN), .ZN(n2520) );
  NAND2_X1 U2609 ( .A1(n2370), .A2(REG1_REG_16__SCAN_IN), .ZN(n2312) );
  NAND2_X1 U2610 ( .A1(n2370), .A2(REG1_REG_15__SCAN_IN), .ZN(n2508) );
  NAND2_X1 U2611 ( .A1(n2370), .A2(REG1_REG_12__SCAN_IN), .ZN(n2481) );
  NAND2_X1 U2612 ( .A1(n2370), .A2(REG1_REG_11__SCAN_IN), .ZN(n2468) );
  NAND2_X1 U2613 ( .A1(n2370), .A2(REG1_REG_9__SCAN_IN), .ZN(n2439) );
  NAND4_X1 U2614 ( .A1(n2416), .A2(n2415), .A3(n2414), .A4(n2413), .ZN(n3878)
         );
  NAND2_X1 U2615 ( .A1(n2370), .A2(REG1_REG_7__SCAN_IN), .ZN(n2415) );
  OR2_X1 U2616 ( .A1(n2371), .A2(n3180), .ZN(n2356) );
  NAND4_X1 U2617 ( .A1(n2348), .A2(n2347), .A3(n2346), .A4(n2345), .ZN(n3882)
         );
  OR2_X1 U2618 ( .A1(n2371), .A2(n2344), .ZN(n2346) );
  OR2_X1 U2619 ( .A1(n2517), .A2(n2328), .ZN(n2142) );
  OR2_X1 U2620 ( .A1(n2371), .A2(n2327), .ZN(n2330) );
  OR2_X1 U2621 ( .A1(n2369), .A2(n2336), .ZN(n2338) );
  NAND2_X1 U2622 ( .A1(n2717), .A2(n2718), .ZN(n3902) );
  XNOR2_X1 U2623 ( .A(n2735), .B(n2734), .ZN(n2733) );
  NAND2_X1 U2624 ( .A1(n2119), .A2(n2120), .ZN(n2118) );
  NAND2_X1 U2625 ( .A1(n2782), .A2(REG2_REG_4__SCAN_IN), .ZN(n2119) );
  INV_X1 U2626 ( .A(n2800), .ZN(n2117) );
  XNOR2_X1 U2627 ( .A(n2766), .B(n2759), .ZN(n2764) );
  OR2_X1 U2628 ( .A1(n2813), .A2(n2812), .ZN(n2816) );
  OR2_X1 U2629 ( .A1(n2773), .A2(n2772), .ZN(n3911) );
  NAND2_X1 U2630 ( .A1(n2112), .A2(n2110), .ZN(n4351) );
  NAND2_X1 U2631 ( .A1(n3927), .A2(n2111), .ZN(n2110) );
  NAND2_X1 U2632 ( .A1(n3926), .A2(REG2_REG_8__SCAN_IN), .ZN(n2112) );
  INV_X1 U2633 ( .A(n3928), .ZN(n2111) );
  NAND2_X1 U2634 ( .A1(n4351), .A2(n4352), .ZN(n4350) );
  AND2_X1 U2635 ( .A1(n3913), .A2(n2133), .ZN(n4345) );
  INV_X1 U2636 ( .A(n4346), .ZN(n2133) );
  INV_X1 U2637 ( .A(n3913), .ZN(n4347) );
  XNOR2_X1 U2638 ( .A(n3914), .B(n4364), .ZN(n4356) );
  INV_X1 U2639 ( .A(n4473), .ZN(n4375) );
  INV_X1 U2640 ( .A(n2131), .ZN(n4376) );
  INV_X1 U2641 ( .A(n3917), .ZN(n2130) );
  NAND2_X1 U2642 ( .A1(n4381), .A2(n3935), .ZN(n4390) );
  INV_X1 U2643 ( .A(n2126), .ZN(n4399) );
  INV_X1 U2644 ( .A(n3939), .ZN(n2125) );
  NAND2_X1 U2645 ( .A1(n3958), .A2(n3959), .ZN(n4423) );
  AND2_X1 U2646 ( .A1(n2710), .A2(n2706), .ZN(n4434) );
  AND2_X1 U2647 ( .A1(n2749), .A2(n2794), .ZN(n4427) );
  INV_X1 U2648 ( .A(n4427), .ZN(n4430) );
  AOI21_X1 U2649 ( .B1(n3961), .B2(REG1_REG_18__SCAN_IN), .A(n4431), .ZN(n3953) );
  XNOR2_X1 U2650 ( .A(n3972), .B(n3971), .ZN(n3566) );
  AND2_X1 U2651 ( .A1(n2592), .A2(n2584), .ZN(n4006) );
  OAI21_X1 U2652 ( .B1(n4011), .B2(n2582), .A(n2171), .ZN(n3994) );
  OR2_X1 U2653 ( .A1(n2018), .A2(n4097), .ZN(n4253) );
  NAND2_X1 U2654 ( .A1(n2175), .A2(n2179), .ZN(n4096) );
  NAND2_X1 U2655 ( .A1(n2183), .A2(n2180), .ZN(n2175) );
  NAND2_X1 U2656 ( .A1(n2182), .A2(n2187), .ZN(n4104) );
  NAND2_X1 U2657 ( .A1(n2183), .A2(n2042), .ZN(n2182) );
  NAND2_X1 U2658 ( .A1(n3327), .A2(n2502), .ZN(n3411) );
  NAND2_X1 U2659 ( .A1(n3263), .A2(n2474), .ZN(n3304) );
  NAND2_X1 U2660 ( .A1(n2395), .A2(n2394), .ZN(n3046) );
  XNOR2_X1 U2661 ( .A(n2599), .B(IR_REG_19__SCAN_IN), .ZN(n2611) );
  INV_X1 U2662 ( .A(n4210), .ZN(n4446) );
  INV_X1 U2663 ( .A(n4524), .ZN(n4522) );
  NAND2_X1 U2664 ( .A1(n4232), .A2(n2086), .ZN(n4288) );
  NOR2_X1 U2665 ( .A1(n2020), .A2(n2087), .ZN(n2086) );
  NOR2_X1 U2666 ( .A1(n4231), .A2(n4510), .ZN(n2087) );
  INV_X2 U2667 ( .A(n4514), .ZN(n4516) );
  NAND2_X1 U2668 ( .A1(n2191), .A2(n2190), .ZN(n4324) );
  NAND2_X1 U2669 ( .A1(n2288), .A2(n2023), .ZN(n2190) );
  NOR2_X1 U2670 ( .A1(IR_REG_31__SCAN_IN), .A2(n3519), .ZN(n2192) );
  AND2_X1 U2671 ( .A1(n2290), .A2(n2288), .ZN(n4325) );
  INV_X1 U2672 ( .A(n2849), .ZN(n4337) );
  INV_X1 U2673 ( .A(n2681), .ZN(n4327) );
  AND2_X1 U2674 ( .A1(n2930), .A2(STATE_REG_SCAN_IN), .ZN(n4461) );
  INV_X1 U2675 ( .A(n2647), .ZN(n4329) );
  XNOR2_X1 U2676 ( .A(n2484), .B(IR_REG_11__SCAN_IN), .ZN(n4473) );
  INV_X1 U2677 ( .A(IR_REG_0__SCAN_IN), .ZN(n2795) );
  INV_X2 U2678 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NAND2_X1 U2679 ( .A1(n2021), .A2(n2062), .ZN(U3226) );
  NOR2_X1 U2680 ( .A1(n3515), .A2(n2063), .ZN(n2062) );
  NOR2_X1 U2681 ( .A1(n3702), .A2(n2064), .ZN(n2063) );
  INV_X1 U2682 ( .A(n2118), .ZN(n2801) );
  AOI21_X1 U2683 ( .B1(n2137), .B2(n2136), .A(n2134), .ZN(n4441) );
  INV_X1 U2684 ( .A(IR_REG_30__SCAN_IN), .ZN(n3519) );
  AND2_X1 U2685 ( .A1(n2233), .A2(n2054), .ZN(n2006) );
  AND2_X1 U2686 ( .A1(n4654), .A2(n2254), .ZN(n2007) );
  AND2_X1 U2687 ( .A1(n2250), .A2(n2247), .ZN(n2008) );
  OR2_X1 U2688 ( .A1(n2589), .A2(n2172), .ZN(n2009) );
  AND2_X1 U2689 ( .A1(n2007), .A2(n2283), .ZN(n2010) );
  AND2_X1 U2690 ( .A1(n2209), .A2(n3002), .ZN(n2011) );
  NAND2_X1 U2691 ( .A1(n2033), .A2(n2184), .ZN(n2179) );
  INV_X1 U2692 ( .A(n4129), .ZN(n2186) );
  AND2_X1 U2693 ( .A1(n3537), .A2(n3536), .ZN(n2012) );
  OAI22_X1 U2694 ( .A1(n3238), .A2(n2462), .B1(n2461), .B2(n3202), .ZN(n3262)
         );
  INV_X1 U2695 ( .A(n3262), .ZN(n2163) );
  OR3_X1 U2696 ( .A1(n3422), .A2(n2048), .A3(n2106), .ZN(n2013) );
  INV_X1 U2697 ( .A(n4054), .ZN(n4017) );
  NAND2_X1 U2698 ( .A1(n2577), .A2(n2576), .ZN(n4054) );
  AND2_X1 U2699 ( .A1(n2056), .A2(n2586), .ZN(n2014) );
  OR3_X1 U2700 ( .A1(n3271), .A2(n2102), .A3(n3351), .ZN(n2015) );
  AND2_X1 U2701 ( .A1(n2057), .A2(n2595), .ZN(n2016) );
  AND2_X1 U2702 ( .A1(n2099), .A2(n4022), .ZN(n2017) );
  NAND2_X1 U2703 ( .A1(n4325), .A2(n4324), .ZN(n2517) );
  OR2_X1 U2704 ( .A1(n3422), .A2(n2103), .ZN(n2018) );
  XOR2_X1 U2705 ( .A(n3552), .B(n3551), .Z(n2019) );
  NAND2_X1 U2706 ( .A1(n2219), .A2(n2218), .ZN(n3567) );
  AND2_X1 U2707 ( .A1(n4230), .A2(n4512), .ZN(n2020) );
  OR2_X1 U2708 ( .A1(n3514), .A2(n3688), .ZN(n2021) );
  AND4_X1 U2709 ( .A1(n2258), .A2(n2282), .A3(n2281), .A4(n4653), .ZN(n2022)
         );
  AND2_X1 U2710 ( .A1(IR_REG_31__SCAN_IN), .A2(n3519), .ZN(n2023) );
  AND2_X1 U2711 ( .A1(n2924), .A2(n2923), .ZN(n2024) );
  AND2_X1 U2712 ( .A1(n2081), .A2(n3786), .ZN(n2025) );
  AND2_X1 U2713 ( .A1(n2145), .A2(n2513), .ZN(n2026) );
  INV_X1 U2714 ( .A(IR_REG_27__SCAN_IN), .ZN(n2283) );
  AND2_X1 U2715 ( .A1(n3353), .A2(n3297), .ZN(n2027) );
  INV_X1 U2716 ( .A(IR_REG_13__SCAN_IN), .ZN(n2278) );
  NOR2_X1 U2717 ( .A1(n3353), .A2(n3297), .ZN(n2028) );
  INV_X1 U2718 ( .A(n2075), .ZN(n2074) );
  NAND2_X1 U2719 ( .A1(n2078), .A2(n2076), .ZN(n2075) );
  NOR2_X1 U2720 ( .A1(n3545), .A2(n3544), .ZN(n2029) );
  INV_X1 U2721 ( .A(n3244), .ZN(n2242) );
  OAI21_X1 U2722 ( .B1(n2589), .B2(n2169), .A(n2170), .ZN(n2168) );
  OR2_X1 U2723 ( .A1(n2807), .A2(n2383), .ZN(n2030) );
  NAND2_X1 U2724 ( .A1(n2246), .A2(n2244), .ZN(n2031) );
  INV_X1 U2725 ( .A(n2222), .ZN(n2221) );
  AND2_X1 U2726 ( .A1(n2787), .A2(n2857), .ZN(n3495) );
  INV_X1 U2727 ( .A(n3495), .ZN(n2958) );
  OR2_X1 U2728 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2032) );
  OR2_X1 U2729 ( .A1(n2185), .A2(n2181), .ZN(n2033) );
  OR2_X1 U2730 ( .A1(n2451), .A2(n2450), .ZN(n2034) );
  NAND2_X1 U2731 ( .A1(n3876), .A2(n3085), .ZN(n2035) );
  AND2_X1 U2732 ( .A1(n2289), .A2(REG0_REG_1__SCAN_IN), .ZN(n2036) );
  INV_X1 U2733 ( .A(n2172), .ZN(n2171) );
  NOR2_X1 U2734 ( .A1(n4036), .A2(n2687), .ZN(n2172) );
  INV_X1 U2735 ( .A(IR_REG_31__SCAN_IN), .ZN(n2349) );
  AND2_X1 U2736 ( .A1(n2287), .A2(IR_REG_30__SCAN_IN), .ZN(n2037) );
  AND2_X1 U2737 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n2038)
         );
  AND2_X1 U2738 ( .A1(n2010), .A2(n2297), .ZN(n2039) );
  INV_X1 U2739 ( .A(n2201), .ZN(n2200) );
  OR2_X1 U2740 ( .A1(n3593), .A2(n2202), .ZN(n2201) );
  INV_X1 U2741 ( .A(n2096), .ZN(n2095) );
  NAND2_X1 U2742 ( .A1(n2097), .A2(n3774), .ZN(n2096) );
  OR2_X1 U2743 ( .A1(n2147), .A2(n2146), .ZN(n2040) );
  NAND2_X1 U2744 ( .A1(n4076), .A2(n2017), .ZN(n2041) );
  INV_X1 U2745 ( .A(IR_REG_28__SCAN_IN), .ZN(n2297) );
  NAND2_X1 U2746 ( .A1(n2324), .A2(n2189), .ZN(n2314) );
  INV_X1 U2747 ( .A(n3762), .ZN(n2071) );
  OR2_X1 U2748 ( .A1(n4154), .A2(n4128), .ZN(n2042) );
  NOR2_X1 U2749 ( .A1(n4054), .A2(n2686), .ZN(n2043) );
  INV_X1 U2750 ( .A(n3606), .ZN(n2225) );
  INV_X1 U2751 ( .A(n2962), .ZN(n3053) );
  NAND2_X1 U2752 ( .A1(n2324), .A2(n2278), .ZN(n2497) );
  OR2_X1 U2753 ( .A1(n2354), .A2(n4263), .ZN(n2044) );
  INV_X1 U2754 ( .A(n2012), .ZN(n2223) );
  AND2_X1 U2755 ( .A1(n2126), .A2(n2125), .ZN(n2045) );
  AND2_X1 U2756 ( .A1(n2131), .A2(n2130), .ZN(n2046) );
  AND2_X1 U2757 ( .A1(n3925), .A2(REG1_REG_9__SCAN_IN), .ZN(n2047) );
  INV_X1 U2758 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2115) );
  NAND2_X1 U2759 ( .A1(n4161), .A2(n4160), .ZN(n2048) );
  INV_X2 U2760 ( .A(n4188), .ZN(n4458) );
  NAND2_X1 U2761 ( .A1(n3025), .A2(n4211), .ZN(n4188) );
  INV_X1 U2762 ( .A(n3596), .ZN(n2202) );
  INV_X1 U2763 ( .A(n3933), .ZN(n4472) );
  NAND2_X1 U2764 ( .A1(n2154), .A2(n2155), .ZN(n3098) );
  NAND2_X1 U2765 ( .A1(n2379), .A2(DATAI_24_), .ZN(n4058) );
  INV_X1 U2766 ( .A(n3647), .ZN(n2199) );
  INV_X1 U2767 ( .A(n3771), .ZN(n2093) );
  INV_X1 U2768 ( .A(n4208), .ZN(n3641) );
  NOR2_X1 U2769 ( .A1(n3222), .A2(n3223), .ZN(n2049) );
  NAND2_X1 U2770 ( .A1(n2549), .A2(DATAI_26_), .ZN(n4022) );
  NOR2_X1 U2771 ( .A1(n2369), .A2(n4529), .ZN(n2050) );
  OR2_X1 U2772 ( .A1(n2354), .A2(n4545), .ZN(n2051) );
  OR2_X1 U2773 ( .A1(n2354), .A2(n2597), .ZN(n2052) );
  INV_X1 U2774 ( .A(n3446), .ZN(n2247) );
  INV_X1 U2775 ( .A(n2101), .ZN(n3357) );
  NOR2_X1 U2776 ( .A1(n3271), .A2(n2102), .ZN(n2101) );
  INV_X1 U2777 ( .A(n3079), .ZN(n2209) );
  AND2_X1 U2778 ( .A1(n2580), .A2(n2069), .ZN(n2053) );
  NAND2_X1 U2779 ( .A1(n3251), .A2(n3252), .ZN(n2054) );
  NAND2_X1 U2780 ( .A1(n2651), .A2(n2010), .ZN(n2055) );
  AND2_X1 U2781 ( .A1(n2587), .A2(n2051), .ZN(n2056) );
  AND2_X1 U2782 ( .A1(n2596), .A2(n2052), .ZN(n2057) );
  NAND2_X1 U2783 ( .A1(n2549), .A2(DATAI_21_), .ZN(n4107) );
  AND2_X1 U2784 ( .A1(n2017), .A2(n3998), .ZN(n2058) );
  NOR2_X2 U2785 ( .A1(n3516), .A2(n2931), .ZN(U4043) );
  NAND2_X1 U2786 ( .A1(n2379), .A2(DATAI_25_), .ZN(n4040) );
  INV_X1 U2787 ( .A(n4040), .ZN(n2686) );
  INV_X1 U2788 ( .A(n2854), .ZN(n2141) );
  AND2_X1 U2789 ( .A1(n2118), .A2(n2117), .ZN(n2060) );
  INV_X1 U2790 ( .A(IR_REG_20__SCAN_IN), .ZN(n2607) );
  AOI21_X2 U2791 ( .B1(n4470), .B2(REG1_REG_13__SCAN_IN), .A(n4385), .ZN(n3918) );
  AOI21_X2 U2792 ( .B1(n4473), .B2(REG1_REG_11__SCAN_IN), .A(n4365), .ZN(n3916) );
  XOR2_X1 U2793 ( .A(n4468), .B(n3918), .Z(n4396) );
  NAND2_X1 U2794 ( .A1(n3923), .A2(n3922), .ZN(n3950) );
  NAND2_X1 U2795 ( .A1(n4420), .A2(n4421), .ZN(n4419) );
  NAND2_X1 U2796 ( .A1(n2802), .A2(n2742), .ZN(n2766) );
  XNOR2_X1 U2797 ( .A(n3912), .B(n3928), .ZN(n2773) );
  NAND2_X1 U2798 ( .A1(n2768), .A2(n2767), .ZN(n2811) );
  NAND2_X1 U2799 ( .A1(n2061), .A2(n3522), .ZN(n3513) );
  INV_X1 U2800 ( .A(n3524), .ZN(n2061) );
  NAND2_X1 U2801 ( .A1(n3222), .A2(n2006), .ZN(n2229) );
  INV_X4 U2802 ( .A(n3550), .ZN(n2978) );
  NAND4_X1 U2803 ( .A1(n2068), .A2(n2067), .A3(n2066), .A4(n2065), .ZN(n2277)
         );
  OAI21_X1 U2804 ( .B1(n3093), .B2(n2096), .A(n2092), .ZN(n3292) );
  OAI21_X1 U2805 ( .B1(n3093), .B2(n3091), .A(n3769), .ZN(n3228) );
  NAND3_X1 U2806 ( .A1(n2105), .A2(n2104), .A3(n4107), .ZN(n2103) );
  NAND2_X1 U2807 ( .A1(n2732), .A2(n2779), .ZN(n2120) );
  OAI21_X1 U2808 ( .B1(n4400), .B2(n2123), .A(n2121), .ZN(n4412) );
  INV_X1 U2809 ( .A(n4413), .ZN(n2127) );
  NAND2_X1 U2810 ( .A1(n3917), .A2(n2132), .ZN(n2128) );
  XNOR2_X2 U2811 ( .A(n3916), .B(n4472), .ZN(n4377) );
  NAND2_X1 U2812 ( .A1(n2141), .A2(n3063), .ZN(n2613) );
  OAI21_X1 U2813 ( .B1(n2489), .B2(n2040), .A(n2144), .ZN(n2143) );
  NOR2_X1 U2814 ( .A1(n2489), .A2(n2488), .ZN(n3329) );
  INV_X1 U2815 ( .A(n2488), .ZN(n2148) );
  NAND2_X1 U2816 ( .A1(n3070), .A2(n2612), .ZN(n3069) );
  NAND2_X1 U2817 ( .A1(n2149), .A2(n2367), .ZN(n3019) );
  NAND3_X1 U2818 ( .A1(n2150), .A2(n2888), .A3(n3069), .ZN(n2149) );
  NAND2_X1 U2819 ( .A1(n2154), .A2(n2152), .ZN(n2151) );
  OAI21_X1 U2820 ( .B1(n3262), .B2(n2161), .A(n2159), .ZN(n3345) );
  OAI21_X1 U2821 ( .B1(n4029), .B2(n2043), .A(n2173), .ZN(n4011) );
  INV_X1 U2822 ( .A(n4121), .ZN(n2183) );
  NAND2_X1 U2823 ( .A1(n4121), .A2(n2179), .ZN(n2174) );
  AOI21_X1 U2824 ( .B1(n2294), .B2(n2037), .A(n2192), .ZN(n2191) );
  NAND2_X1 U2825 ( .A1(n2291), .A2(n2036), .ZN(n2331) );
  INV_X1 U2826 ( .A(IR_REG_0__SCAN_IN), .ZN(n2193) );
  NAND3_X1 U2827 ( .A1(n2350), .A2(n2193), .A3(n2333), .ZN(n2359) );
  AND2_X2 U2828 ( .A1(n2196), .A2(n2194), .ZN(n3658) );
  OR2_X2 U2829 ( .A1(n3648), .A2(n2201), .ZN(n2196) );
  NAND2_X1 U2830 ( .A1(n2203), .A2(n2205), .ZN(n3193) );
  NAND3_X1 U2831 ( .A1(n2977), .A2(n2976), .A3(n2011), .ZN(n2203) );
  NAND2_X1 U2832 ( .A1(n3605), .A2(n2211), .ZN(n2210) );
  OAI211_X1 U2833 ( .C1(n3605), .C2(n2215), .A(n2212), .B(n2210), .ZN(n3557)
         );
  NAND2_X1 U2834 ( .A1(n3605), .A2(n2220), .ZN(n2219) );
  AOI21_X1 U2835 ( .B1(n3605), .B2(n3606), .A(n3607), .ZN(n3679) );
  NAND3_X1 U2836 ( .A1(n3568), .A2(n2224), .A3(n2223), .ZN(n2222) );
  INV_X1 U2837 ( .A(n3447), .ZN(n2243) );
  NAND2_X1 U2838 ( .A1(n2651), .A2(n4654), .ZN(n2654) );
  NAND2_X1 U2839 ( .A1(n2651), .A2(n2039), .ZN(n2639) );
  XNOR2_X2 U2840 ( .A(n2332), .B(n2333), .ZN(n3889) );
  NAND2_X1 U2841 ( .A1(n4094), .A2(n2550), .ZN(n4064) );
  OR2_X1 U2842 ( .A1(n2517), .A2(n3038), .ZN(n2375) );
  INV_X1 U2843 ( .A(n2517), .ZN(n2585) );
  OAI21_X2 U2844 ( .B1(n3524), .B2(n3523), .A(n3522), .ZN(n3605) );
  NAND2_X1 U2845 ( .A1(n2946), .A2(n2945), .ZN(n2255) );
  AND2_X1 U2846 ( .A1(n2361), .A2(n2377), .ZN(n2256) );
  AND3_X1 U2847 ( .A1(n2607), .A2(n2606), .A3(n2605), .ZN(n2257) );
  AND4_X1 U2848 ( .A1(n2315), .A2(n2667), .A3(n2606), .A4(n2280), .ZN(n2258)
         );
  NAND2_X1 U2849 ( .A1(n3168), .A2(n2365), .ZN(n2259) );
  OR2_X1 U2850 ( .A1(n3867), .A2(n3578), .ZN(n2260) );
  INV_X1 U2851 ( .A(n4097), .ZN(n3662) );
  AND2_X1 U2852 ( .A1(n2549), .A2(DATAI_22_), .ZN(n4097) );
  INV_X1 U2853 ( .A(IR_REG_14__SCAN_IN), .ZN(n2279) );
  AND2_X1 U2854 ( .A1(n2315), .A2(n2317), .ZN(n2261) );
  INV_X1 U2855 ( .A(n3390), .ZN(n3399) );
  OR2_X1 U2856 ( .A1(n3558), .A2(n4320), .ZN(n2262) );
  OR2_X1 U2857 ( .A1(n3558), .A2(n4275), .ZN(n2263) );
  OAI211_X1 U2858 ( .C1(n4098), .C2(n2641), .A(n2548), .B(n2547), .ZN(n4110)
         );
  INV_X1 U2859 ( .A(IR_REG_22__SCAN_IN), .ZN(n2280) );
  INV_X1 U2860 ( .A(IR_REG_18__SCAN_IN), .ZN(n2532) );
  NOR2_X1 U2861 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n4653)
         );
  NOR2_X1 U2862 ( .A1(n4091), .A2(n4078), .ZN(n2560) );
  INV_X1 U2863 ( .A(n2516), .ZN(n2273) );
  INV_X1 U2864 ( .A(n4468), .ZN(n3937) );
  OR2_X1 U2865 ( .A1(n3880), .A2(n3037), .ZN(n3754) );
  NAND2_X1 U2866 ( .A1(n2712), .A2(n2297), .ZN(n2299) );
  OR2_X1 U2867 ( .A1(n3384), .A2(n3383), .ZN(n3385) );
  OAI21_X1 U2868 ( .B1(n2958), .B2(n3068), .A(n2855), .ZN(n2858) );
  OR2_X1 U2869 ( .A1(n2826), .A2(n2825), .ZN(n2828) );
  AOI21_X1 U2870 ( .B1(n4064), .B2(n2260), .A(n2560), .ZN(n2561) );
  NAND2_X1 U2871 ( .A1(n4110), .A2(n4097), .ZN(n2550) );
  NAND2_X1 U2872 ( .A1(n2273), .A2(REG3_REG_18__SCAN_IN), .ZN(n2526) );
  NAND2_X1 U2873 ( .A1(n2272), .A2(REG3_REG_16__SCAN_IN), .ZN(n2514) );
  AND2_X1 U2874 ( .A1(n3872), .A2(n3351), .ZN(n2488) );
  OR2_X1 U2875 ( .A1(n2435), .A2(n2268), .ZN(n2453) );
  INV_X1 U2876 ( .A(n3151), .ZN(n3156) );
  AND2_X1 U2877 ( .A1(n3884), .A2(n3062), .ZN(n3070) );
  OR2_X1 U2878 ( .A1(n2583), .A2(n3569), .ZN(n2592) );
  OR2_X1 U2879 ( .A1(n2453), .A2(n4601), .ZN(n2464) );
  XNOR2_X1 U2880 ( .A(n2858), .B(n3547), .ZN(n2876) );
  INV_X1 U2881 ( .A(n4036), .ZN(n3999) );
  NAND2_X1 U2882 ( .A1(n2920), .A2(n2919), .ZN(n2926) );
  INV_X1 U2883 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3661) );
  NAND2_X1 U2884 ( .A1(n3624), .A2(n2957), .ZN(n2975) );
  OR2_X1 U2885 ( .A1(n2578), .A2(n3682), .ZN(n2583) );
  INV_X1 U2886 ( .A(IR_REG_3__SCAN_IN), .ZN(n2361) );
  INV_X1 U2887 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3314) );
  INV_X1 U2888 ( .A(REG3_REG_15__SCAN_IN), .ZN(n3695) );
  INV_X1 U2889 ( .A(REG3_REG_17__SCAN_IN), .ZN(n3639) );
  INV_X1 U2890 ( .A(n4326), .ZN(n2794) );
  INV_X1 U2891 ( .A(n4022), .ZN(n2687) );
  INV_X1 U2892 ( .A(n2561), .ZN(n4047) );
  INV_X1 U2893 ( .A(n3454), .ZN(n3617) );
  NAND2_X1 U2894 ( .A1(n2705), .A2(n4337), .ZN(n4204) );
  OR2_X1 U2895 ( .A1(n2826), .A2(D_REG_0__SCAN_IN), .ZN(n2684) );
  INV_X1 U2896 ( .A(n4107), .ZN(n4113) );
  AND2_X1 U2897 ( .A1(n3768), .A2(n3764), .ZN(n3815) );
  AND2_X1 U2898 ( .A1(n3756), .A2(n3760), .ZN(n3833) );
  INV_X1 U2899 ( .A(n4196), .ZN(n4158) );
  INV_X1 U2900 ( .A(n2911), .ZN(n3179) );
  OR2_X1 U2901 ( .A1(n2540), .A2(n3600), .ZN(n2545) );
  AND2_X1 U2902 ( .A1(n2851), .A2(n2850), .ZN(n3697) );
  INV_X1 U2903 ( .A(n3702), .ZN(n3686) );
  OR3_X1 U2904 ( .A1(n3546), .A2(n3516), .A3(n2856), .ZN(n3862) );
  NAND2_X1 U2905 ( .A1(n2581), .A2(n2053), .ZN(n4036) );
  OR2_X1 U2906 ( .A1(n2369), .A2(n2368), .ZN(n2374) );
  OR2_X1 U2907 ( .A1(n2371), .A2(n2335), .ZN(n2340) );
  AND2_X1 U2908 ( .A1(n2749), .A2(n2849), .ZN(n4403) );
  INV_X1 U2909 ( .A(n4204), .ZN(n4155) );
  NAND2_X1 U2910 ( .A1(n3741), .A2(n2637), .ZN(n4196) );
  AND2_X1 U2911 ( .A1(n2836), .A2(n2835), .ZN(n4453) );
  AND2_X1 U2912 ( .A1(n2684), .A2(n2683), .ZN(n2829) );
  INV_X1 U2913 ( .A(n4512), .ZN(n4501) );
  NAND2_X1 U2914 ( .A1(n4135), .A2(n4484), .ZN(n4512) );
  INV_X1 U2915 ( .A(n2829), .ZN(n3024) );
  INV_X1 U2916 ( .A(n4461), .ZN(n3516) );
  INV_X1 U2917 ( .A(n2665), .ZN(n2682) );
  AND2_X1 U2918 ( .A1(n2935), .A2(n2934), .ZN(n3702) );
  NAND2_X1 U2919 ( .A1(n2851), .A2(n2833), .ZN(n3688) );
  NAND2_X1 U2920 ( .A1(n2568), .A2(n2567), .ZN(n4073) );
  INV_X1 U2921 ( .A(n4439), .ZN(n4398) );
  INV_X1 U2922 ( .A(n4475), .ZN(n4364) );
  INV_X1 U2923 ( .A(n4466), .ZN(n4417) );
  NAND2_X1 U2924 ( .A1(n4188), .A2(n3104), .ZN(n4217) );
  OR2_X1 U2925 ( .A1(n4183), .A2(n4510), .ZN(n4210) );
  NAND2_X1 U2926 ( .A1(n4524), .A2(n4489), .ZN(n4275) );
  AND2_X2 U2927 ( .A1(n2690), .A2(n2829), .ZN(n4524) );
  NAND2_X1 U2928 ( .A1(n4516), .A2(n4489), .ZN(n4320) );
  NAND2_X1 U2929 ( .A1(n2690), .A2(n3024), .ZN(n4514) );
  INV_X1 U2930 ( .A(n4460), .ZN(n4459) );
  NAND2_X1 U2931 ( .A1(n2826), .A2(n2836), .ZN(n4460) );
  INV_X1 U2932 ( .A(n3960), .ZN(n4465) );
  NAND2_X1 U2933 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2399) );
  INV_X1 U2934 ( .A(n2399), .ZN(n2266) );
  AND2_X1 U2935 ( .A1(REG3_REG_5__SCAN_IN), .A2(REG3_REG_6__SCAN_IN), .ZN(
        n2265) );
  NAND2_X1 U2936 ( .A1(n2266), .A2(n2265), .ZN(n2411) );
  INV_X1 U2937 ( .A(n2411), .ZN(n2267) );
  NAND2_X1 U2938 ( .A1(n2267), .A2(REG3_REG_7__SCAN_IN), .ZN(n2435) );
  NAND2_X1 U2939 ( .A1(REG3_REG_8__SCAN_IN), .A2(REG3_REG_9__SCAN_IN), .ZN(
        n2268) );
  INV_X1 U2940 ( .A(n2464), .ZN(n2269) );
  NAND2_X1 U2941 ( .A1(n2269), .A2(REG3_REG_11__SCAN_IN), .ZN(n2476) );
  INV_X1 U2942 ( .A(n2476), .ZN(n2270) );
  NAND2_X1 U2943 ( .A1(n2270), .A2(REG3_REG_12__SCAN_IN), .ZN(n2478) );
  INV_X1 U2944 ( .A(n2491), .ZN(n2271) );
  NAND2_X1 U2945 ( .A1(n2271), .A2(REG3_REG_14__SCAN_IN), .ZN(n2503) );
  INV_X1 U2946 ( .A(n2526), .ZN(n2274) );
  NAND2_X1 U2947 ( .A1(n2540), .A2(n3600), .ZN(n2275) );
  NAND2_X1 U2948 ( .A1(n2545), .A2(n2275), .ZN(n4115) );
  INV_X1 U2949 ( .A(n2359), .ZN(n2276) );
  NAND2_X1 U2950 ( .A1(n2276), .A2(n2256), .ZN(n2388) );
  NOR2_X2 U2951 ( .A1(n2388), .A2(n2277), .ZN(n2324) );
  NOR2_X1 U2952 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(n2282)
         );
  NOR2_X1 U2953 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2281)
         );
  NAND2_X1 U2954 ( .A1(n2639), .A2(IR_REG_31__SCAN_IN), .ZN(n2284) );
  AOI22_X1 U2955 ( .A1(n2370), .A2(REG1_REG_21__SCAN_IN), .B1(n2352), .B2(
        REG0_REG_21__SCAN_IN), .ZN(n2293) );
  NAND2_X1 U2956 ( .A1(n2594), .A2(REG2_REG_21__SCAN_IN), .ZN(n2292) );
  OAI211_X1 U2957 ( .C1(n4115), .C2(n2641), .A(n2293), .B(n2292), .ZN(n4129)
         );
  NAND2_X1 U2958 ( .A1(n2295), .A2(n2283), .ZN(n2712) );
  NAND2_X1 U2959 ( .A1(n2662), .A2(n2296), .ZN(n2711) );
  NOR2_X2 U2960 ( .A1(n2522), .A2(IR_REG_17__SCAN_IN), .ZN(n2533) );
  INV_X1 U2961 ( .A(n2533), .ZN(n2301) );
  NAND2_X1 U2962 ( .A1(n2301), .A2(IR_REG_31__SCAN_IN), .ZN(n2302) );
  XNOR2_X1 U2963 ( .A(n2302), .B(IR_REG_18__SCAN_IN), .ZN(n3961) );
  MUX2_X1 U2964 ( .A(n3961), .B(DATAI_18_), .S(n2549), .Z(n4181) );
  NAND2_X1 U2965 ( .A1(n2594), .A2(REG2_REG_18__SCAN_IN), .ZN(n2307) );
  INV_X1 U2966 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3948) );
  INV_X1 U2967 ( .A(REG0_REG_18__SCAN_IN), .ZN(n4527) );
  OR2_X1 U2968 ( .A1(n2369), .A2(n4527), .ZN(n2305) );
  INV_X1 U2969 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4575) );
  NAND2_X1 U2970 ( .A1(n2516), .A2(n4575), .ZN(n2303) );
  NAND2_X1 U2971 ( .A1(n2526), .A2(n2303), .ZN(n4184) );
  OR2_X1 U2972 ( .A1(n2641), .A2(n4184), .ZN(n2304) );
  NAND4_X1 U2973 ( .A1(n2307), .A2(n2306), .A3(n2305), .A4(n2304), .ZN(n4201)
         );
  NAND2_X1 U2974 ( .A1(n2352), .A2(REG0_REG_16__SCAN_IN), .ZN(n2313) );
  INV_X1 U2975 ( .A(REG1_REG_16__SCAN_IN), .ZN(n3922) );
  INV_X1 U2976 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2308) );
  NAND2_X1 U2977 ( .A1(n2505), .A2(n2308), .ZN(n2309) );
  NAND2_X1 U2978 ( .A1(n2514), .A2(n2309), .ZN(n3620) );
  OR2_X1 U2979 ( .A1(n2641), .A2(n3620), .ZN(n2311) );
  INV_X1 U2980 ( .A(REG2_REG_16__SCAN_IN), .ZN(n3424) );
  OR2_X1 U2981 ( .A1(n2371), .A2(n3424), .ZN(n2310) );
  NAND4_X1 U2982 ( .A1(n2313), .A2(n2312), .A3(n2311), .A4(n2310), .ZN(n3869)
         );
  INV_X1 U2983 ( .A(n3869), .ZN(n4205) );
  NAND2_X1 U2984 ( .A1(n2314), .A2(IR_REG_31__SCAN_IN), .ZN(n2510) );
  NAND2_X1 U2985 ( .A1(n2510), .A2(n2315), .ZN(n2316) );
  NAND2_X1 U2986 ( .A1(n2316), .A2(IR_REG_31__SCAN_IN), .ZN(n2318) );
  XNOR2_X1 U2987 ( .A(n2318), .B(n2317), .ZN(n3956) );
  INV_X1 U2988 ( .A(DATAI_16_), .ZN(n4591) );
  MUX2_X1 U2989 ( .A(n3956), .B(n4591), .S(n2549), .Z(n3454) );
  NAND2_X1 U2990 ( .A1(n2352), .A2(REG0_REG_13__SCAN_IN), .ZN(n2323) );
  INV_X1 U2991 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4535) );
  NAND2_X1 U2992 ( .A1(n2478), .A2(n3314), .ZN(n2319) );
  NAND2_X1 U2993 ( .A1(n2491), .A2(n2319), .ZN(n3359) );
  OR2_X1 U2994 ( .A1(n2517), .A2(n3359), .ZN(n2321) );
  INV_X1 U2995 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3360) );
  OR2_X1 U2996 ( .A1(n2371), .A2(n3360), .ZN(n2320) );
  NAND4_X1 U2997 ( .A1(n2323), .A2(n2322), .A3(n2321), .A4(n2320), .ZN(n3872)
         );
  INV_X1 U2998 ( .A(n3872), .ZN(n3334) );
  OR2_X1 U2999 ( .A1(n2324), .A2(n2349), .ZN(n2325) );
  XNOR2_X1 U3000 ( .A(n2325), .B(IR_REG_13__SCAN_IN), .ZN(n4470) );
  INV_X1 U3001 ( .A(DATAI_13_), .ZN(n2326) );
  MUX2_X1 U3002 ( .A(n4394), .B(n2326), .S(n2549), .Z(n3358) );
  INV_X1 U3003 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2327) );
  INV_X1 U3004 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2328) );
  INV_X1 U3005 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2716) );
  INV_X1 U3006 ( .A(IR_REG_1__SCAN_IN), .ZN(n2333) );
  INV_X1 U3007 ( .A(DATAI_1_), .ZN(n2334) );
  MUX2_X1 U3008 ( .A(n3889), .B(n2334), .S(n2379), .Z(n3068) );
  NAND2_X1 U3009 ( .A1(n2854), .A2(n3068), .ZN(n3746) );
  NAND2_X1 U3010 ( .A1(n2613), .A2(n3746), .ZN(n2612) );
  INV_X1 U3011 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2335) );
  INV_X1 U3012 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2752) );
  OR2_X1 U3013 ( .A1(n2517), .A2(n2752), .ZN(n2339) );
  INV_X1 U3014 ( .A(REG0_REG_0__SCAN_IN), .ZN(n2336) );
  INV_X1 U3015 ( .A(REG1_REG_0__SCAN_IN), .ZN(n3891) );
  INV_X1 U3016 ( .A(DATAI_0_), .ZN(n2341) );
  MUX2_X1 U3017 ( .A(n2795), .B(n2341), .S(n2379), .Z(n2821) );
  INV_X1 U3018 ( .A(n2821), .ZN(n3062) );
  INV_X1 U3019 ( .A(n3068), .ZN(n3063) );
  NAND2_X1 U3020 ( .A1(n2854), .A2(n3063), .ZN(n2342) );
  NAND2_X1 U3021 ( .A1(n2585), .A2(REG3_REG_2__SCAN_IN), .ZN(n2348) );
  INV_X1 U3022 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2343) );
  OR2_X1 U3023 ( .A1(n2369), .A2(n2343), .ZN(n2347) );
  INV_X1 U3024 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2344) );
  INV_X1 U3025 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2713) );
  OR2_X1 U3026 ( .A1(n2354), .A2(n2713), .ZN(n2345) );
  INV_X1 U3027 ( .A(DATAI_2_), .ZN(n2351) );
  MUX2_X1 U3028 ( .A(n3897), .B(n2351), .S(n2379), .Z(n2899) );
  NAND2_X1 U3029 ( .A1(n3882), .A2(n2899), .ZN(n3751) );
  NAND2_X1 U3030 ( .A1(n2352), .A2(REG0_REG_3__SCAN_IN), .ZN(n2358) );
  OR2_X1 U3031 ( .A1(n2517), .A2(REG3_REG_3__SCAN_IN), .ZN(n2357) );
  INV_X1 U3032 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3180) );
  INV_X1 U3033 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2353) );
  OR2_X1 U3034 ( .A1(n2354), .A2(n2353), .ZN(n2355) );
  NAND2_X1 U3035 ( .A1(n2360), .A2(IR_REG_31__SCAN_IN), .ZN(n2362) );
  NAND2_X1 U3036 ( .A1(n2362), .A2(n2361), .ZN(n2376) );
  OR2_X1 U3037 ( .A1(n2362), .A2(n2361), .ZN(n2363) );
  NAND2_X1 U3038 ( .A1(n2376), .A2(n2363), .ZN(n2734) );
  INV_X1 U3039 ( .A(DATAI_3_), .ZN(n2364) );
  MUX2_X1 U3040 ( .A(n2734), .B(n2364), .S(n2379), .Z(n2911) );
  NAND2_X1 U3041 ( .A1(n3881), .A2(n3179), .ZN(n2366) );
  NAND2_X1 U3042 ( .A1(n3173), .A2(n2899), .ZN(n3168) );
  INV_X1 U3043 ( .A(n3881), .ZN(n2896) );
  NAND2_X1 U3044 ( .A1(n2896), .A2(n2911), .ZN(n2365) );
  NAND2_X1 U3045 ( .A1(n2366), .A2(n2259), .ZN(n2367) );
  INV_X1 U3046 ( .A(n3019), .ZN(n2380) );
  OAI21_X1 U3047 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        n2399), .ZN(n3038) );
  INV_X1 U3048 ( .A(REG0_REG_4__SCAN_IN), .ZN(n2368) );
  NAND2_X1 U3049 ( .A1(n2370), .A2(REG1_REG_4__SCAN_IN), .ZN(n2373) );
  OR2_X1 U3050 ( .A1(n2371), .A2(n2115), .ZN(n2372) );
  NAND4_X2 U3051 ( .A1(n2375), .A2(n2374), .A3(n2373), .A4(n2372), .ZN(n3880)
         );
  NAND2_X1 U3052 ( .A1(n2376), .A2(IR_REG_31__SCAN_IN), .ZN(n2378) );
  XNOR2_X1 U3053 ( .A(n2378), .B(n2377), .ZN(n2731) );
  INV_X1 U3054 ( .A(DATAI_4_), .ZN(n2694) );
  MUX2_X1 U3055 ( .A(n2731), .B(n2694), .S(n2379), .Z(n3037) );
  NAND2_X1 U3056 ( .A1(n3880), .A2(n3037), .ZN(n3757) );
  NAND2_X1 U3057 ( .A1(n3754), .A2(n3757), .ZN(n3028) );
  INV_X1 U3058 ( .A(n3028), .ZN(n3836) );
  NAND2_X1 U3059 ( .A1(n2380), .A2(n3028), .ZN(n3021) );
  INV_X1 U3060 ( .A(n3037), .ZN(n2938) );
  NAND2_X1 U3061 ( .A1(n3880), .A2(n2938), .ZN(n2381) );
  NAND2_X1 U3062 ( .A1(n3021), .A2(n2381), .ZN(n3118) );
  NAND2_X1 U3063 ( .A1(n2370), .A2(REG1_REG_5__SCAN_IN), .ZN(n2387) );
  INV_X1 U3064 ( .A(REG0_REG_5__SCAN_IN), .ZN(n2382) );
  OR2_X1 U3065 ( .A1(n2369), .A2(n2382), .ZN(n2386) );
  INV_X1 U3066 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2398) );
  XNOR2_X1 U3067 ( .A(n2399), .B(n2398), .ZN(n3629) );
  OR2_X1 U3068 ( .A1(n2517), .A2(n3629), .ZN(n2385) );
  INV_X1 U3069 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2383) );
  OR2_X1 U3070 ( .A1(n2371), .A2(n2383), .ZN(n2384) );
  NAND4_X1 U3071 ( .A1(n2387), .A2(n2386), .A3(n2385), .A4(n2384), .ZN(n3033)
         );
  INV_X1 U3072 ( .A(n3033), .ZN(n3050) );
  NAND2_X1 U3073 ( .A1(n2388), .A2(IR_REG_31__SCAN_IN), .ZN(n2389) );
  MUX2_X1 U3074 ( .A(IR_REG_31__SCAN_IN), .B(n2389), .S(IR_REG_5__SCAN_IN), 
        .Z(n2391) );
  NOR2_X1 U3075 ( .A1(n2388), .A2(IR_REG_5__SCAN_IN), .ZN(n2418) );
  INV_X1 U3076 ( .A(n2418), .ZN(n2390) );
  NAND2_X1 U3077 ( .A1(n2391), .A2(n2390), .ZN(n2807) );
  INV_X1 U3078 ( .A(DATAI_5_), .ZN(n2392) );
  MUX2_X1 U3079 ( .A(n2807), .B(n2392), .S(n2549), .Z(n3120) );
  NAND2_X1 U3080 ( .A1(n3050), .A2(n3120), .ZN(n2393) );
  NAND2_X1 U3081 ( .A1(n3118), .A2(n2393), .ZN(n2395) );
  INV_X1 U3082 ( .A(n3120), .ZN(n3628) );
  NAND2_X1 U3083 ( .A1(n3033), .A2(n3628), .ZN(n2394) );
  NAND2_X1 U3084 ( .A1(n2370), .A2(REG1_REG_6__SCAN_IN), .ZN(n2405) );
  INV_X1 U3085 ( .A(REG0_REG_6__SCAN_IN), .ZN(n2396) );
  OR2_X1 U3086 ( .A1(n2369), .A2(n2396), .ZN(n2404) );
  INV_X1 U3087 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2397) );
  OAI21_X1 U3088 ( .B1(n2399), .B2(n2398), .A(n2397), .ZN(n2400) );
  NAND2_X1 U3089 ( .A1(n2400), .A2(n2411), .ZN(n3143) );
  OR2_X1 U3090 ( .A1(n2641), .A2(n3143), .ZN(n2403) );
  INV_X1 U3091 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2401) );
  OR2_X1 U3092 ( .A1(n2371), .A2(n2401), .ZN(n2402) );
  NAND4_X1 U3093 ( .A1(n2405), .A2(n2404), .A3(n2403), .A4(n2402), .ZN(n3879)
         );
  OR2_X1 U3094 ( .A1(n2418), .A2(n2349), .ZN(n2406) );
  XNOR2_X1 U3095 ( .A(n2406), .B(n2417), .ZN(n2759) );
  INV_X1 U3096 ( .A(DATAI_6_), .ZN(n2407) );
  MUX2_X1 U3097 ( .A(n2759), .B(n2407), .S(n2549), .Z(n2962) );
  AND2_X1 U3098 ( .A1(n3879), .A2(n3053), .ZN(n2408) );
  NAND2_X1 U3099 ( .A1(n2352), .A2(REG0_REG_7__SCAN_IN), .ZN(n2416) );
  INV_X1 U3100 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2770) );
  INV_X1 U3101 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2409) );
  OR2_X1 U3102 ( .A1(n2371), .A2(n2409), .ZN(n2414) );
  INV_X1 U3103 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2410) );
  NAND2_X1 U3104 ( .A1(n2411), .A2(n2410), .ZN(n2412) );
  NAND2_X1 U3105 ( .A1(n2435), .A2(n2412), .ZN(n3161) );
  OR2_X1 U3106 ( .A1(n2641), .A2(n3161), .ZN(n2413) );
  NAND2_X1 U3107 ( .A1(n2418), .A2(n2417), .ZN(n2441) );
  NAND2_X1 U3108 ( .A1(n2441), .A2(IR_REG_31__SCAN_IN), .ZN(n2420) );
  NAND2_X1 U3109 ( .A1(n2420), .A2(n2419), .ZN(n2427) );
  OR2_X1 U3110 ( .A1(n2420), .A2(n2419), .ZN(n2421) );
  NAND2_X1 U3111 ( .A1(n2427), .A2(n2421), .ZN(n4331) );
  INV_X1 U3112 ( .A(DATAI_7_), .ZN(n4594) );
  MUX2_X1 U3113 ( .A(n4331), .B(n4594), .S(n2549), .Z(n3151) );
  NAND2_X1 U3114 ( .A1(n3878), .A2(n3151), .ZN(n3765) );
  NAND2_X1 U3115 ( .A1(n2370), .A2(REG1_REG_8__SCAN_IN), .ZN(n2426) );
  INV_X1 U3116 ( .A(REG0_REG_8__SCAN_IN), .ZN(n2422) );
  OR2_X1 U3117 ( .A1(n2369), .A2(n2422), .ZN(n2425) );
  INV_X1 U3118 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2434) );
  XNOR2_X1 U3119 ( .A(n2435), .B(n2434), .ZN(n3186) );
  OR2_X1 U3120 ( .A1(n2641), .A2(n3186), .ZN(n2424) );
  INV_X1 U3121 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3929) );
  OR2_X1 U3122 ( .A1(n2371), .A2(n3929), .ZN(n2423) );
  NAND4_X1 U3123 ( .A1(n2426), .A2(n2425), .A3(n2424), .A4(n2423), .ZN(n3877)
         );
  INV_X1 U3124 ( .A(n3877), .ZN(n2430) );
  NAND2_X1 U3125 ( .A1(n2427), .A2(IR_REG_31__SCAN_IN), .ZN(n2429) );
  INV_X1 U3126 ( .A(IR_REG_8__SCAN_IN), .ZN(n2428) );
  XNOR2_X1 U3127 ( .A(n2429), .B(n2428), .ZN(n3928) );
  INV_X1 U3128 ( .A(DATAI_8_), .ZN(n2697) );
  MUX2_X1 U3129 ( .A(n3928), .B(n2697), .S(n2549), .Z(n3129) );
  AND2_X1 U3130 ( .A1(n2430), .A2(n3129), .ZN(n2449) );
  INV_X1 U3131 ( .A(n2449), .ZN(n2431) );
  NAND2_X1 U3132 ( .A1(n2352), .A2(REG0_REG_9__SCAN_IN), .ZN(n2440) );
  INV_X1 U3133 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2432) );
  INV_X1 U3134 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2433) );
  OAI21_X1 U3135 ( .B1(n2435), .B2(n2434), .A(n2433), .ZN(n2436) );
  NAND2_X1 U3136 ( .A1(n2436), .A2(n2453), .ZN(n3107) );
  OR2_X1 U3137 ( .A1(n2641), .A2(n3107), .ZN(n2438) );
  INV_X1 U3138 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3108) );
  OR2_X1 U3139 ( .A1(n2371), .A2(n3108), .ZN(n2437) );
  NAND4_X1 U3140 ( .A1(n2440), .A2(n2439), .A3(n2438), .A4(n2437), .ZN(n3876)
         );
  INV_X1 U3141 ( .A(n3876), .ZN(n3230) );
  NAND2_X1 U3142 ( .A1(n2443), .A2(IR_REG_31__SCAN_IN), .ZN(n2442) );
  MUX2_X1 U3143 ( .A(IR_REG_31__SCAN_IN), .B(n2442), .S(IR_REG_9__SCAN_IN), 
        .Z(n2445) );
  INV_X1 U3144 ( .A(n2470), .ZN(n2444) );
  NAND2_X1 U3145 ( .A1(n2445), .A2(n2444), .ZN(n4477) );
  INV_X1 U3146 ( .A(DATAI_9_), .ZN(n4595) );
  MUX2_X1 U3147 ( .A(n4477), .B(n4595), .S(n2549), .Z(n3106) );
  AND2_X1 U31480 ( .A1(n3230), .A2(n3106), .ZN(n2451) );
  INV_X1 U31490 ( .A(n3106), .ZN(n3085) );
  NAND2_X1 U3150 ( .A1(n3878), .A2(n3156), .ZN(n3126) );
  INV_X1 U3151 ( .A(n3129), .ZN(n3135) );
  NAND2_X1 U3152 ( .A1(n3877), .A2(n3135), .ZN(n2447) );
  AND2_X1 U3153 ( .A1(n3126), .A2(n2447), .ZN(n2448) );
  OR2_X1 U3154 ( .A1(n2449), .A2(n2448), .ZN(n3100) );
  AND2_X1 U3155 ( .A1(n2035), .A2(n3100), .ZN(n2450) );
  NAND2_X1 U3156 ( .A1(n2370), .A2(REG1_REG_10__SCAN_IN), .ZN(n2458) );
  INV_X1 U3157 ( .A(REG0_REG_10__SCAN_IN), .ZN(n2452) );
  OR2_X1 U3158 ( .A1(n2369), .A2(n2452), .ZN(n2457) );
  NAND2_X1 U3159 ( .A1(n2453), .A2(n4601), .ZN(n2454) );
  NAND2_X1 U3160 ( .A1(n2464), .A2(n2454), .ZN(n3236) );
  OR2_X1 U3161 ( .A1(n2641), .A2(n3236), .ZN(n2456) );
  INV_X1 U3162 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3237) );
  OR2_X1 U3163 ( .A1(n2371), .A2(n3237), .ZN(n2455) );
  NAND4_X1 U3164 ( .A1(n2458), .A2(n2457), .A3(n2456), .A4(n2455), .ZN(n3875)
         );
  OR2_X1 U3165 ( .A1(n2470), .A2(n2349), .ZN(n2459) );
  XNOR2_X1 U3166 ( .A(n2459), .B(IR_REG_10__SCAN_IN), .ZN(n4475) );
  INV_X1 U3167 ( .A(DATAI_10_), .ZN(n2460) );
  MUX2_X1 U3168 ( .A(n4364), .B(n2460), .S(n2549), .Z(n3202) );
  NOR2_X1 U3169 ( .A1(n3875), .A2(n3233), .ZN(n2462) );
  INV_X1 U3170 ( .A(n3875), .ZN(n2461) );
  NAND2_X1 U3171 ( .A1(n2352), .A2(REG0_REG_11__SCAN_IN), .ZN(n2469) );
  INV_X1 U3172 ( .A(REG1_REG_11__SCAN_IN), .ZN(n2463) );
  INV_X1 U3173 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3215) );
  NAND2_X1 U3174 ( .A1(n2464), .A2(n3215), .ZN(n2465) );
  NAND2_X1 U3175 ( .A1(n2476), .A2(n2465), .ZN(n3275) );
  OR2_X1 U3176 ( .A1(n2641), .A2(n3275), .ZN(n2467) );
  INV_X1 U3177 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3276) );
  OR2_X1 U3178 ( .A1(n2371), .A2(n3276), .ZN(n2466) );
  NAND4_X1 U3179 ( .A1(n2469), .A2(n2468), .A3(n2467), .A4(n2466), .ZN(n3874)
         );
  NAND2_X1 U3180 ( .A1(n2470), .A2(n4655), .ZN(n2471) );
  NAND2_X1 U3181 ( .A1(n2471), .A2(IR_REG_31__SCAN_IN), .ZN(n2484) );
  INV_X1 U3182 ( .A(DATAI_11_), .ZN(n2472) );
  MUX2_X1 U3183 ( .A(n4375), .B(n2472), .S(n2549), .Z(n3273) );
  OR2_X1 U3184 ( .A1(n3874), .A2(n3273), .ZN(n3289) );
  NAND2_X1 U3185 ( .A1(n3874), .A2(n3273), .ZN(n3291) );
  NAND2_X1 U3186 ( .A1(n3289), .A2(n3291), .ZN(n3264) );
  INV_X1 U3187 ( .A(n3264), .ZN(n3838) );
  INV_X1 U3188 ( .A(n3874), .ZN(n2473) );
  NAND2_X1 U3189 ( .A1(n2473), .A2(n3273), .ZN(n2474) );
  NAND2_X1 U3190 ( .A1(n2352), .A2(REG0_REG_12__SCAN_IN), .ZN(n2482) );
  INV_X1 U3191 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4378) );
  INV_X1 U3192 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2475) );
  NAND2_X1 U3193 ( .A1(n2476), .A2(n2475), .ZN(n2477) );
  NAND2_X1 U3194 ( .A1(n2478), .A2(n2477), .ZN(n3300) );
  OR2_X1 U3195 ( .A1(n2641), .A2(n3300), .ZN(n2480) );
  INV_X1 U3196 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3301) );
  OR2_X1 U3197 ( .A1(n2371), .A2(n3301), .ZN(n2479) );
  NAND4_X1 U3198 ( .A1(n2482), .A2(n2481), .A3(n2480), .A4(n2479), .ZN(n3873)
         );
  INV_X1 U3199 ( .A(n3873), .ZN(n3353) );
  INV_X1 U3200 ( .A(IR_REG_11__SCAN_IN), .ZN(n2483) );
  NAND2_X1 U3201 ( .A1(n2484), .A2(n2483), .ZN(n2485) );
  NAND2_X1 U3202 ( .A1(n2485), .A2(IR_REG_31__SCAN_IN), .ZN(n2486) );
  XNOR2_X1 U3203 ( .A(n2486), .B(IR_REG_12__SCAN_IN), .ZN(n3933) );
  INV_X1 U3204 ( .A(DATAI_12_), .ZN(n2487) );
  MUX2_X1 U3205 ( .A(n4472), .B(n2487), .S(n2549), .Z(n3297) );
  INV_X1 U3206 ( .A(n3297), .ZN(n3256) );
  AOI21_X1 U3207 ( .B1(n3334), .B2(n3358), .A(n3345), .ZN(n2489) );
  NAND2_X1 U3208 ( .A1(n2352), .A2(REG0_REG_14__SCAN_IN), .ZN(n2496) );
  INV_X1 U3209 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4397) );
  INV_X1 U32100 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2490) );
  NAND2_X1 U32110 ( .A1(n2491), .A2(n2490), .ZN(n2492) );
  NAND2_X1 U32120 ( .A1(n2503), .A2(n2492), .ZN(n3402) );
  OR2_X1 U32130 ( .A1(n2517), .A2(n3402), .ZN(n2494) );
  INV_X1 U32140 ( .A(REG2_REG_14__SCAN_IN), .ZN(n3337) );
  OR2_X1 U32150 ( .A1(n2371), .A2(n3337), .ZN(n2493) );
  NAND4_X1 U32160 ( .A1(n2496), .A2(n2495), .A3(n2494), .A4(n2493), .ZN(n3871)
         );
  NAND2_X1 U32170 ( .A1(n2497), .A2(IR_REG_31__SCAN_IN), .ZN(n2498) );
  MUX2_X1 U32180 ( .A(IR_REG_31__SCAN_IN), .B(n2498), .S(IR_REG_14__SCAN_IN), 
        .Z(n2499) );
  AND2_X1 U32190 ( .A1(n2499), .A2(n2314), .ZN(n4468) );
  INV_X1 U32200 ( .A(DATAI_14_), .ZN(n2500) );
  MUX2_X1 U32210 ( .A(n3937), .B(n2500), .S(n2549), .Z(n3390) );
  OR2_X1 U32220 ( .A1(n3871), .A2(n3390), .ZN(n3711) );
  NAND2_X1 U32230 ( .A1(n3871), .A2(n3390), .ZN(n3712) );
  NAND2_X1 U32240 ( .A1(n3711), .A2(n3712), .ZN(n3328) );
  NAND2_X1 U32250 ( .A1(n2352), .A2(REG0_REG_15__SCAN_IN), .ZN(n2509) );
  INV_X1 U32260 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3920) );
  NAND2_X1 U32270 ( .A1(n2503), .A2(n3695), .ZN(n2504) );
  NAND2_X1 U32280 ( .A1(n2505), .A2(n2504), .ZN(n3701) );
  OR2_X1 U32290 ( .A1(n2517), .A2(n3701), .ZN(n2507) );
  INV_X1 U32300 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3414) );
  OR2_X1 U32310 ( .A1(n2371), .A2(n3414), .ZN(n2506) );
  NAND4_X1 U32320 ( .A1(n2509), .A2(n2508), .A3(n2507), .A4(n2506), .ZN(n3870)
         );
  XNOR2_X1 U32330 ( .A(n2510), .B(IR_REG_15__SCAN_IN), .ZN(n4466) );
  INV_X1 U32340 ( .A(DATAI_15_), .ZN(n2511) );
  MUX2_X1 U32350 ( .A(n4417), .B(n2511), .S(n2549), .Z(n3459) );
  INV_X1 U32360 ( .A(n3459), .ZN(n3698) );
  NAND2_X1 U32370 ( .A1(n3870), .A2(n3698), .ZN(n2513) );
  INV_X1 U32380 ( .A(n3870), .ZN(n3430) );
  OR2_X1 U32390 ( .A1(n3869), .A2(n3454), .ZN(n3784) );
  NAND2_X1 U32400 ( .A1(n3869), .A2(n3454), .ZN(n4192) );
  NAND2_X1 U32410 ( .A1(n3784), .A2(n4192), .ZN(n3420) );
  NAND2_X1 U32420 ( .A1(n3421), .A2(n3420), .ZN(n3419) );
  OAI21_X1 U32430 ( .B1(n4205), .B2(n3454), .A(n3419), .ZN(n4191) );
  NAND2_X1 U32440 ( .A1(n2352), .A2(REG0_REG_17__SCAN_IN), .ZN(n2521) );
  INV_X1 U32450 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4273) );
  NAND2_X1 U32460 ( .A1(n2514), .A2(n3639), .ZN(n2515) );
  NAND2_X1 U32470 ( .A1(n2516), .A2(n2515), .ZN(n4212) );
  OR2_X1 U32480 ( .A1(n2517), .A2(n4212), .ZN(n2519) );
  INV_X1 U32490 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4213) );
  OR2_X1 U32500 ( .A1(n2371), .A2(n4213), .ZN(n2518) );
  NAND4_X1 U32510 ( .A1(n2521), .A2(n2520), .A3(n2519), .A4(n2518), .ZN(n3868)
         );
  INV_X1 U32520 ( .A(n3868), .ZN(n4178) );
  NAND2_X1 U32530 ( .A1(n2522), .A2(IR_REG_31__SCAN_IN), .ZN(n2523) );
  XNOR2_X1 U32540 ( .A(n2523), .B(IR_REG_17__SCAN_IN), .ZN(n3960) );
  INV_X1 U32550 ( .A(DATAI_17_), .ZN(n4464) );
  MUX2_X1 U32560 ( .A(n4465), .B(n4464), .S(n2549), .Z(n4208) );
  NAND2_X1 U32570 ( .A1(n4178), .A2(n4208), .ZN(n2524) );
  AOI22_X1 U32580 ( .A1(n4191), .A2(n2524), .B1(n3641), .B2(n3868), .ZN(n4172)
         );
  OR2_X1 U32590 ( .A1(n4201), .A2(n4161), .ZN(n4148) );
  NAND2_X1 U32600 ( .A1(n4201), .A2(n4161), .ZN(n4149) );
  NAND2_X1 U32610 ( .A1(n4148), .A2(n4149), .ZN(n4171) );
  NAND2_X1 U32620 ( .A1(n4172), .A2(n4171), .ZN(n4170) );
  OAI21_X1 U32630 ( .B1(n4181), .B2(n4201), .A(n4170), .ZN(n4145) );
  NAND2_X1 U32640 ( .A1(n2352), .A2(REG0_REG_19__SCAN_IN), .ZN(n2531) );
  INV_X1 U32650 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4543) );
  INV_X1 U32660 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2525) );
  NAND2_X1 U32670 ( .A1(n2526), .A2(n2525), .ZN(n2527) );
  NAND2_X1 U32680 ( .A1(n2538), .A2(n2527), .ZN(n4164) );
  OR2_X1 U32690 ( .A1(n2641), .A2(n4164), .ZN(n2529) );
  INV_X1 U32700 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4165) );
  OR2_X1 U32710 ( .A1(n2371), .A2(n4165), .ZN(n2528) );
  NAND4_X1 U32720 ( .A1(n2531), .A2(n2530), .A3(n2529), .A4(n2528), .ZN(n4176)
         );
  NAND2_X1 U32730 ( .A1(n2533), .A2(n2532), .ZN(n2604) );
  INV_X1 U32740 ( .A(DATAI_19_), .ZN(n2534) );
  MUX2_X1 U32750 ( .A(n2838), .B(n2534), .S(n2549), .Z(n4160) );
  INV_X1 U32760 ( .A(n4160), .ZN(n3587) );
  NAND2_X1 U32770 ( .A1(n4176), .A2(n3587), .ZN(n2535) );
  NAND2_X1 U32780 ( .A1(n4145), .A2(n2535), .ZN(n2537) );
  INV_X1 U32790 ( .A(n4176), .ZN(n4131) );
  NAND2_X1 U32800 ( .A1(n2537), .A2(n2536), .ZN(n4121) );
  NAND2_X1 U32810 ( .A1(n2538), .A2(n3651), .ZN(n2539) );
  NAND2_X1 U32820 ( .A1(n2540), .A2(n2539), .ZN(n4138) );
  NAND2_X1 U32830 ( .A1(n2594), .A2(REG2_REG_20__SCAN_IN), .ZN(n2541) );
  OAI21_X1 U32840 ( .B1(n4138), .B2(n2641), .A(n2541), .ZN(n2544) );
  INV_X1 U32850 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4263) );
  NAND2_X1 U32860 ( .A1(n2352), .A2(REG0_REG_20__SCAN_IN), .ZN(n2542) );
  INV_X1 U32870 ( .A(n4137), .ZN(n4128) );
  NAND2_X1 U32880 ( .A1(n2545), .A2(n3661), .ZN(n2546) );
  NAND2_X1 U32890 ( .A1(n2553), .A2(n2546), .ZN(n4098) );
  AOI22_X1 U32900 ( .A1(n2594), .A2(REG2_REG_22__SCAN_IN), .B1(n2352), .B2(
        REG0_REG_22__SCAN_IN), .ZN(n2548) );
  NAND2_X1 U32910 ( .A1(n2370), .A2(REG1_REG_22__SCAN_IN), .ZN(n2547) );
  OR2_X1 U32920 ( .A1(n4110), .A2(n3662), .ZN(n4068) );
  NAND2_X1 U32930 ( .A1(n4110), .A2(n3662), .ZN(n2632) );
  NAND2_X1 U32940 ( .A1(n4068), .A2(n2632), .ZN(n4095) );
  INV_X1 U32950 ( .A(n4110), .ZN(n4071) );
  INV_X1 U32960 ( .A(n2553), .ZN(n2551) );
  INV_X1 U32970 ( .A(REG3_REG_23__SCAN_IN), .ZN(n2552) );
  NAND2_X1 U32980 ( .A1(n2553), .A2(n2552), .ZN(n2554) );
  NAND2_X1 U32990 ( .A1(n2562), .A2(n2554), .ZN(n4080) );
  OR2_X1 U33000 ( .A1(n4080), .A2(n2641), .ZN(n2559) );
  INV_X1 U33010 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4081) );
  NAND2_X1 U33020 ( .A1(n2370), .A2(REG1_REG_23__SCAN_IN), .ZN(n2556) );
  NAND2_X1 U33030 ( .A1(n2352), .A2(REG0_REG_23__SCAN_IN), .ZN(n2555) );
  OAI211_X1 U33040 ( .C1(n4081), .C2(n2371), .A(n2556), .B(n2555), .ZN(n2557)
         );
  INV_X1 U33050 ( .A(n2557), .ZN(n2558) );
  NAND2_X1 U33060 ( .A1(n2562), .A2(n3444), .ZN(n2563) );
  NAND2_X1 U33070 ( .A1(n4059), .A2(n2585), .ZN(n2568) );
  INV_X1 U33080 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4526) );
  NAND2_X1 U33090 ( .A1(n2370), .A2(REG1_REG_24__SCAN_IN), .ZN(n2565) );
  NAND2_X1 U33100 ( .A1(n2594), .A2(REG2_REG_24__SCAN_IN), .ZN(n2564) );
  OAI211_X1 U33110 ( .C1(n2369), .C2(n4526), .A(n2565), .B(n2564), .ZN(n2566)
         );
  INV_X1 U33120 ( .A(n2566), .ZN(n2567) );
  NOR2_X1 U33130 ( .A1(n4034), .A2(n4058), .ZN(n2569) );
  INV_X1 U33140 ( .A(n4058), .ZN(n3441) );
  INV_X1 U33150 ( .A(n2571), .ZN(n2570) );
  NAND2_X1 U33160 ( .A1(n2570), .A2(REG3_REG_25__SCAN_IN), .ZN(n2578) );
  INV_X1 U33170 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4602) );
  NAND2_X1 U33180 ( .A1(n2571), .A2(n4602), .ZN(n2572) );
  NAND2_X1 U33190 ( .A1(n2578), .A2(n2572), .ZN(n3609) );
  OR2_X1 U33200 ( .A1(n3609), .A2(n2641), .ZN(n2577) );
  INV_X1 U33210 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4530) );
  NAND2_X1 U33220 ( .A1(n2370), .A2(REG1_REG_25__SCAN_IN), .ZN(n2574) );
  NAND2_X1 U33230 ( .A1(n2594), .A2(REG2_REG_25__SCAN_IN), .ZN(n2573) );
  OAI211_X1 U33240 ( .C1(n2369), .C2(n4530), .A(n2574), .B(n2573), .ZN(n2575)
         );
  INV_X1 U33250 ( .A(n2575), .ZN(n2576) );
  INV_X1 U33260 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3682) );
  NAND2_X1 U33270 ( .A1(n2578), .A2(n3682), .ZN(n2579) );
  NAND2_X1 U33280 ( .A1(n4024), .A2(n2585), .ZN(n2581) );
  INV_X1 U33290 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4546) );
  NAND2_X1 U33300 ( .A1(n2594), .A2(REG2_REG_26__SCAN_IN), .ZN(n2580) );
  INV_X1 U33310 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4529) );
  NOR2_X1 U33320 ( .A1(n3999), .A2(n4022), .ZN(n2582) );
  INV_X1 U33330 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3569) );
  NAND2_X1 U33340 ( .A1(n2583), .A2(n3569), .ZN(n2584) );
  NAND2_X1 U33350 ( .A1(n4006), .A2(n2585), .ZN(n2588) );
  INV_X1 U33360 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4545) );
  NAND2_X1 U33370 ( .A1(n2594), .A2(REG2_REG_27__SCAN_IN), .ZN(n2587) );
  NAND2_X1 U33380 ( .A1(n2352), .A2(REG0_REG_27__SCAN_IN), .ZN(n2586) );
  INV_X1 U33390 ( .A(n3998), .ZN(n4005) );
  NOR2_X1 U33400 ( .A1(n4019), .A2(n4005), .ZN(n2589) );
  INV_X1 U33410 ( .A(n4019), .ZN(n3744) );
  INV_X1 U33420 ( .A(n2592), .ZN(n2590) );
  NAND2_X1 U33430 ( .A1(n2590), .A2(REG3_REG_28__SCAN_IN), .ZN(n3984) );
  INV_X1 U33440 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2591) );
  NAND2_X1 U33450 ( .A1(n2592), .A2(n2591), .ZN(n2593) );
  NAND2_X1 U33460 ( .A1(n3984), .A2(n2593), .ZN(n3560) );
  INV_X1 U33470 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2597) );
  NAND2_X1 U33480 ( .A1(n2594), .A2(REG2_REG_28__SCAN_IN), .ZN(n2596) );
  NAND2_X1 U33490 ( .A1(n2352), .A2(REG0_REG_28__SCAN_IN), .ZN(n2595) );
  NAND2_X1 U33500 ( .A1(n2379), .A2(DATAI_28_), .ZN(n3549) );
  NAND2_X1 U33510 ( .A1(n4001), .A2(n3549), .ZN(n3974) );
  INV_X1 U33520 ( .A(n3549), .ZN(n3970) );
  NAND2_X1 U3353 ( .A1(n3982), .A2(n3970), .ZN(n3975) );
  NAND2_X1 U33540 ( .A1(n3974), .A2(n3975), .ZN(n3971) );
  NAND2_X1 U3355 ( .A1(n2599), .A2(n2606), .ZN(n2600) );
  NAND2_X1 U3356 ( .A1(n2600), .A2(IR_REG_31__SCAN_IN), .ZN(n2601) );
  XNOR2_X2 U3357 ( .A(n2601), .B(n2607), .ZN(n2688) );
  OAI21_X1 U3358 ( .B1(IR_REG_20__SCAN_IN), .B2(IR_REG_19__SCAN_IN), .A(
        IR_REG_31__SCAN_IN), .ZN(n2602) );
  INV_X1 U3359 ( .A(n2604), .ZN(n2608) );
  INV_X1 U3360 ( .A(IR_REG_21__SCAN_IN), .ZN(n2605) );
  NAND2_X1 U3361 ( .A1(n2608), .A2(n2257), .ZN(n2656) );
  NAND2_X1 U3362 ( .A1(n2656), .A2(IR_REG_31__SCAN_IN), .ZN(n2609) );
  XNOR2_X1 U3363 ( .A(n3026), .B(n3858), .ZN(n2610) );
  NAND2_X1 U3364 ( .A1(n2688), .A2(n2611), .ZN(n4451) );
  OR2_X1 U3365 ( .A1(n4451), .A2(n4328), .ZN(n4484) );
  OR2_X1 U3366 ( .A1(n3884), .A2(n2821), .ZN(n3066) );
  OAI21_X1 U3367 ( .B1(n2612), .B2(n3066), .A(n2613), .ZN(n2891) );
  INV_X1 U3368 ( .A(n2888), .ZN(n3835) );
  OR2_X1 U3369 ( .A1(n3881), .A2(n2911), .ZN(n3753) );
  NAND2_X1 U3370 ( .A1(n3881), .A2(n2911), .ZN(n3750) );
  INV_X1 U3371 ( .A(n3754), .ZN(n2614) );
  OR2_X1 U3372 ( .A1(n3029), .A2(n2614), .ZN(n2615) );
  NAND2_X1 U3373 ( .A1(n2615), .A2(n3757), .ZN(n3113) );
  AND2_X1 U3374 ( .A1(n3033), .A2(n3120), .ZN(n3112) );
  OR2_X1 U3375 ( .A1(n3033), .A2(n3120), .ZN(n3760) );
  NAND2_X1 U3376 ( .A1(n3879), .A2(n2962), .ZN(n3045) );
  NOR2_X1 U3377 ( .A1(n3879), .A2(n2962), .ZN(n3762) );
  NAND2_X1 U3378 ( .A1(n2616), .A2(n3765), .ZN(n3128) );
  OR2_X1 U3379 ( .A1(n3877), .A2(n3129), .ZN(n3768) );
  NAND2_X1 U3380 ( .A1(n3128), .A2(n3768), .ZN(n2617) );
  NAND2_X1 U3381 ( .A1(n3877), .A2(n3129), .ZN(n3764) );
  NAND2_X1 U3382 ( .A1(n2617), .A2(n3764), .ZN(n3093) );
  AND2_X1 U3383 ( .A1(n3876), .A2(n3106), .ZN(n3091) );
  OR2_X1 U3384 ( .A1(n3876), .A2(n3106), .ZN(n3769) );
  NAND2_X1 U3385 ( .A1(n3875), .A2(n3202), .ZN(n3774) );
  OR2_X1 U3386 ( .A1(n3875), .A2(n3202), .ZN(n3771) );
  NAND2_X1 U3387 ( .A1(n3873), .A2(n3297), .ZN(n3346) );
  NAND2_X1 U3388 ( .A1(n3872), .A2(n3358), .ZN(n3342) );
  NAND2_X1 U3389 ( .A1(n3346), .A2(n3342), .ZN(n2619) );
  INV_X1 U3390 ( .A(n3291), .ZN(n2618) );
  NOR2_X1 U3391 ( .A1(n2619), .A2(n2618), .ZN(n3775) );
  NAND2_X1 U3392 ( .A1(n3292), .A2(n3775), .ZN(n2622) );
  INV_X1 U3393 ( .A(n2619), .ZN(n2621) );
  OR2_X1 U3394 ( .A1(n3873), .A2(n3297), .ZN(n3348) );
  NAND2_X1 U3395 ( .A1(n3289), .A2(n3348), .ZN(n2620) );
  NOR2_X1 U3396 ( .A1(n3872), .A2(n3358), .ZN(n3343) );
  AOI21_X1 U3397 ( .B1(n2621), .B2(n2620), .A(n3343), .ZN(n3777) );
  NAND2_X1 U3398 ( .A1(n2622), .A2(n3777), .ZN(n3717) );
  INV_X1 U3399 ( .A(n3328), .ZN(n3832) );
  NAND2_X1 U3400 ( .A1(n3717), .A2(n3832), .ZN(n2623) );
  NAND2_X1 U3401 ( .A1(n2623), .A2(n3711), .ZN(n3408) );
  OR2_X1 U3402 ( .A1(n3870), .A2(n3459), .ZN(n3715) );
  NAND2_X1 U3403 ( .A1(n3870), .A2(n3459), .ZN(n3713) );
  NAND2_X1 U3404 ( .A1(n3715), .A2(n3713), .ZN(n3822) );
  INV_X1 U3405 ( .A(n3420), .ZN(n3828) );
  NAND2_X1 U3406 ( .A1(n3868), .A2(n4208), .ZN(n3812) );
  AND2_X1 U3407 ( .A1(n4192), .A2(n3812), .ZN(n3718) );
  NAND2_X1 U3408 ( .A1(n4176), .A2(n4160), .ZN(n2624) );
  AND2_X1 U3409 ( .A1(n4149), .A2(n2624), .ZN(n4122) );
  OR2_X1 U3410 ( .A1(n3868), .A2(n4208), .ZN(n4146) );
  NAND2_X1 U3411 ( .A1(n4148), .A2(n4146), .ZN(n2626) );
  NOR2_X1 U3412 ( .A1(n4176), .A2(n4160), .ZN(n2625) );
  AOI21_X1 U3413 ( .B1(n4122), .B2(n2626), .A(n2625), .ZN(n4123) );
  NAND2_X1 U3414 ( .A1(n4108), .A2(n4128), .ZN(n2627) );
  AND2_X1 U3415 ( .A1(n4123), .A2(n2627), .ZN(n2628) );
  NAND2_X1 U3416 ( .A1(n4147), .A2(n2628), .ZN(n2631) );
  INV_X1 U3417 ( .A(n2628), .ZN(n3787) );
  OR2_X1 U3418 ( .A1(n3787), .A2(n4122), .ZN(n2630) );
  NAND2_X1 U3419 ( .A1(n4154), .A2(n4137), .ZN(n2629) );
  OR2_X1 U3420 ( .A1(n4129), .A2(n4107), .ZN(n4066) );
  AND2_X1 U3421 ( .A1(n4068), .A2(n4066), .ZN(n3790) );
  NAND2_X1 U3422 ( .A1(n3867), .A2(n4078), .ZN(n3811) );
  AND2_X1 U3423 ( .A1(n3811), .A2(n2632), .ZN(n3794) );
  AND2_X1 U3424 ( .A1(n4129), .A2(n4107), .ZN(n4065) );
  NAND2_X1 U3425 ( .A1(n4068), .A2(n4065), .ZN(n2633) );
  NAND2_X1 U3426 ( .A1(n3794), .A2(n2633), .ZN(n3722) );
  NAND2_X1 U3427 ( .A1(n4034), .A2(n3441), .ZN(n3820) );
  NAND2_X1 U3428 ( .A1(n4091), .A2(n3578), .ZN(n4048) );
  NAND2_X1 U3429 ( .A1(n3820), .A2(n4048), .ZN(n3792) );
  NAND2_X1 U3430 ( .A1(n3999), .A2(n2687), .ZN(n3808) );
  NAND2_X1 U3431 ( .A1(n4017), .A2(n2686), .ZN(n4012) );
  AND2_X1 U3432 ( .A1(n3808), .A2(n4012), .ZN(n3728) );
  INV_X1 U3433 ( .A(n3728), .ZN(n3791) );
  NAND2_X1 U3434 ( .A1(n4054), .A2(n4040), .ZN(n3810) );
  NAND2_X1 U3435 ( .A1(n4073), .A2(n4058), .ZN(n4030) );
  AND2_X1 U3436 ( .A1(n3810), .A2(n4030), .ZN(n3724) );
  INV_X1 U3437 ( .A(n3724), .ZN(n4013) );
  NAND2_X1 U3438 ( .A1(n3728), .A2(n4013), .ZN(n2634) );
  AND2_X1 U3439 ( .A1(n4036), .A2(n4022), .ZN(n3735) );
  INV_X1 U3440 ( .A(n3735), .ZN(n3809) );
  NAND2_X1 U3441 ( .A1(n2634), .A2(n3809), .ZN(n3796) );
  INV_X1 U3442 ( .A(n3796), .ZN(n2635) );
  XNOR2_X1 U3443 ( .A(n4019), .B(n3998), .ZN(n3997) );
  NOR2_X1 U3444 ( .A1(n3996), .A2(n3997), .ZN(n3995) );
  OR2_X1 U3445 ( .A1(n4019), .A2(n3998), .ZN(n3727) );
  INV_X1 U3446 ( .A(n3727), .ZN(n3730) );
  NOR2_X1 U3447 ( .A1(n3995), .A2(n3730), .ZN(n3977) );
  XNOR2_X1 U3448 ( .A(n3977), .B(n3971), .ZN(n2650) );
  OR2_X1 U3449 ( .A1(n2647), .A2(n2688), .ZN(n3741) );
  NAND2_X1 U3450 ( .A1(n4328), .A2(n2611), .ZN(n2637) );
  NAND2_X1 U3451 ( .A1(n4328), .A2(n4329), .ZN(n2830) );
  NAND2_X1 U3452 ( .A1(n2055), .A2(IR_REG_31__SCAN_IN), .ZN(n2638) );
  MUX2_X1 U3453 ( .A(IR_REG_31__SCAN_IN), .B(n2638), .S(IR_REG_28__SCAN_IN), 
        .Z(n2640) );
  NAND2_X1 U3454 ( .A1(n2640), .A2(n2639), .ZN(n2849) );
  OR2_X1 U3455 ( .A1(n3984), .A2(n2641), .ZN(n2646) );
  INV_X1 U3456 ( .A(REG2_REG_29__SCAN_IN), .ZN(n3989) );
  NAND2_X1 U3457 ( .A1(n2352), .A2(REG0_REG_29__SCAN_IN), .ZN(n2643) );
  NAND2_X1 U34580 ( .A1(n2370), .A2(REG1_REG_29__SCAN_IN), .ZN(n2642) );
  OAI211_X1 U34590 ( .C1(n3989), .C2(n2371), .A(n2643), .B(n2642), .ZN(n2644)
         );
  INV_X1 U3460 ( .A(n2644), .ZN(n2645) );
  NAND2_X1 U3461 ( .A1(n2646), .A2(n2645), .ZN(n3866) );
  NAND2_X1 U3462 ( .A1(n2705), .A2(n2849), .ZN(n4090) );
  INV_X1 U3463 ( .A(n2688), .ZN(n4330) );
  AOI22_X1 U3464 ( .A1(n3866), .A2(n4200), .B1(n3970), .B2(n4227), .ZN(n2648)
         );
  OAI21_X1 U3465 ( .B1(n3744), .B2(n4204), .A(n2648), .ZN(n2649) );
  AOI21_X1 U3466 ( .B1(n2650), .B2(n4196), .A(n2649), .ZN(n3561) );
  OAI21_X1 U34670 ( .B1(n3566), .B2(n4501), .A(n3561), .ZN(n2691) );
  INV_X1 U3468 ( .A(n2651), .ZN(n2652) );
  NAND2_X1 U34690 ( .A1(n2652), .A2(IR_REG_31__SCAN_IN), .ZN(n2653) );
  MUX2_X1 U3470 ( .A(IR_REG_31__SCAN_IN), .B(n2653), .S(IR_REG_25__SCAN_IN), 
        .Z(n2655) );
  NAND2_X1 U34710 ( .A1(n2655), .A2(n2654), .ZN(n2700) );
  NAND2_X1 U3472 ( .A1(n2700), .A2(B_REG_SCAN_IN), .ZN(n2659) );
  OAI21_X2 U34730 ( .B1(n2656), .B2(IR_REG_22__SCAN_IN), .A(IR_REG_31__SCAN_IN), .ZN(n2666) );
  NAND2_X1 U3474 ( .A1(n2666), .A2(n2667), .ZN(n2657) );
  MUX2_X1 U34750 ( .A(n2659), .B(B_REG_SCAN_IN), .S(n2665), .Z(n2663) );
  NAND2_X1 U3476 ( .A1(n2654), .A2(IR_REG_31__SCAN_IN), .ZN(n2660) );
  MUX2_X1 U34770 ( .A(IR_REG_31__SCAN_IN), .B(n2660), .S(IR_REG_26__SCAN_IN), 
        .Z(n2661) );
  NAND2_X1 U3478 ( .A1(n2681), .A2(n2700), .ZN(n2827) );
  OAI21_X1 U34790 ( .B1(n2826), .B2(D_REG_1__SCAN_IN), .A(n2827), .ZN(n2680)
         );
  NOR2_X1 U3480 ( .A1(n2681), .A2(n2700), .ZN(n2664) );
  NAND2_X1 U34810 ( .A1(n2688), .A2(n2838), .ZN(n2668) );
  NAND2_X1 U3482 ( .A1(n2705), .A2(n2668), .ZN(n2929) );
  NAND2_X1 U34830 ( .A1(n2836), .A2(n2929), .ZN(n2844) );
  NOR2_X1 U3484 ( .A1(n2844), .A2(n2835), .ZN(n2679) );
  NOR4_X1 U34850 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_18__SCAN_IN), .A3(
        D_REG_19__SCAN_IN), .A4(D_REG_21__SCAN_IN), .ZN(n2672) );
  NOR4_X1 U3486 ( .A1(D_REG_12__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_17__SCAN_IN), .A4(D_REG_15__SCAN_IN), .ZN(n2671) );
  NOR4_X1 U34870 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_29__SCAN_IN), .ZN(n2670) );
  NOR4_X1 U3488 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_25__SCAN_IN), .A3(
        D_REG_23__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2669) );
  NAND4_X1 U34890 ( .A1(n2672), .A2(n2671), .A3(n2670), .A4(n2669), .ZN(n2677)
         );
  NOR2_X1 U3490 ( .A1(D_REG_5__SCAN_IN), .A2(D_REG_13__SCAN_IN), .ZN(n4651) );
  NOR4_X1 U34910 ( .A1(D_REG_30__SCAN_IN), .A2(D_REG_31__SCAN_IN), .A3(
        D_REG_20__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2675) );
  NOR4_X1 U3492 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_9__SCAN_IN), .A3(
        D_REG_10__SCAN_IN), .A4(D_REG_11__SCAN_IN), .ZN(n2674) );
  NOR4_X1 U34930 ( .A1(D_REG_3__SCAN_IN), .A2(D_REG_2__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_6__SCAN_IN), .ZN(n2673) );
  NAND4_X1 U3494 ( .A1(n4651), .A2(n2675), .A3(n2674), .A4(n2673), .ZN(n2676)
         );
  NOR2_X1 U34950 ( .A1(n2677), .A2(n2676), .ZN(n2824) );
  OR2_X1 U3496 ( .A1(n2826), .A2(n2824), .ZN(n2678) );
  NAND2_X1 U34970 ( .A1(n2682), .A2(n2681), .ZN(n2683) );
  MUX2_X1 U3498 ( .A(REG1_REG_28__SCAN_IN), .B(n2691), .S(n4524), .Z(n2685) );
  INV_X1 U34990 ( .A(n2685), .ZN(n2689) );
  AND2_X1 U3500 ( .A1(n3068), .A2(n2821), .ZN(n3061) );
  NAND2_X1 U35010 ( .A1(n3061), .A2(n2899), .ZN(n3178) );
  NOR2_X1 U3502 ( .A1(n3178), .A2(n3179), .ZN(n3177) );
  NAND2_X1 U35030 ( .A1(n3160), .A2(n3129), .ZN(n3105) );
  INV_X1 U3504 ( .A(n3273), .ZN(n3216) );
  NAND2_X1 U35050 ( .A1(n3413), .A2(n3459), .ZN(n3423) );
  NAND2_X1 U35060 ( .A1(n4004), .A2(n3549), .ZN(n3986) );
  OAI21_X1 U35070 ( .B1(n4004), .B2(n3549), .A(n3986), .ZN(n3558) );
  NAND2_X1 U35080 ( .A1(n2689), .A2(n2263), .ZN(U3546) );
  MUX2_X1 U35090 ( .A(REG0_REG_28__SCAN_IN), .B(n2691), .S(n4516), .Z(n2692)
         );
  INV_X1 U35100 ( .A(n2692), .ZN(n2693) );
  NAND2_X1 U35110 ( .A1(n2693), .A2(n2262), .ZN(U3514) );
  MUX2_X1 U35120 ( .A(n2694), .B(n2731), .S(STATE_REG_SCAN_IN), .Z(n2695) );
  INV_X1 U35130 ( .A(n2695), .ZN(U3348) );
  MUX2_X1 U35140 ( .A(n2759), .B(n2407), .S(U3149), .Z(n2696) );
  INV_X1 U35150 ( .A(n2696), .ZN(U3346) );
  MUX2_X1 U35160 ( .A(n2697), .B(n3928), .S(STATE_REG_SCAN_IN), .Z(n2698) );
  INV_X1 U35170 ( .A(n2698), .ZN(U3344) );
  NAND2_X1 U35180 ( .A1(U3149), .A2(DATAI_16_), .ZN(n2699) );
  OAI21_X1 U35190 ( .B1(n3956), .B2(U3149), .A(n2699), .ZN(U3336) );
  INV_X1 U35200 ( .A(DATAI_25_), .ZN(n4589) );
  INV_X1 U35210 ( .A(n2700), .ZN(n2701) );
  NAND2_X1 U35220 ( .A1(n2701), .A2(STATE_REG_SCAN_IN), .ZN(n2702) );
  OAI21_X1 U35230 ( .B1(STATE_REG_SCAN_IN), .B2(n4589), .A(n2702), .ZN(U3327)
         );
  MUX2_X1 U35240 ( .A(n2534), .B(n2838), .S(STATE_REG_SCAN_IN), .Z(n2703) );
  INV_X1 U35250 ( .A(n2703), .ZN(U3333) );
  NOR2_X1 U35260 ( .A1(n2930), .A2(U3149), .ZN(n3859) );
  OR2_X1 U35270 ( .A1(n2836), .A2(n3859), .ZN(n2710) );
  AOI21_X1 U35280 ( .B1(n2705), .B2(n2930), .A(n2704), .ZN(n2709) );
  INV_X1 U35290 ( .A(n2709), .ZN(n2706) );
  NOR2_X1 U35300 ( .A1(n4434), .A2(U4043), .ZN(U3148) );
  INV_X1 U35310 ( .A(D_REG_1__SCAN_IN), .ZN(n4612) );
  INV_X1 U35320 ( .A(n2827), .ZN(n2707) );
  AOI22_X1 U35330 ( .A1(n4460), .A2(n4612), .B1(n2707), .B2(n4461), .ZN(U3459)
         );
  INV_X1 U35340 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n4566) );
  NAND2_X1 U35350 ( .A1(n3033), .A2(U4043), .ZN(n2708) );
  OAI21_X1 U35360 ( .B1(U4043), .B2(n4566), .A(n2708), .ZN(U3555) );
  INV_X1 U35370 ( .A(n4403), .ZN(n4442) );
  AND2_X1 U35380 ( .A1(n2712), .A2(n2711), .ZN(n4326) );
  MUX2_X1 U35390 ( .A(n2713), .B(REG1_REG_2__SCAN_IN), .S(n3897), .Z(n2718) );
  MUX2_X1 U35400 ( .A(n2716), .B(REG1_REG_1__SCAN_IN), .S(n3889), .Z(n2715) );
  OR2_X1 U35410 ( .A1(n3889), .A2(n2716), .ZN(n3898) );
  NAND2_X1 U35420 ( .A1(n3899), .A2(n3898), .ZN(n2717) );
  INV_X1 U35430 ( .A(n3897), .ZN(n4335) );
  NAND2_X1 U35440 ( .A1(n4335), .A2(REG1_REG_2__SCAN_IN), .ZN(n2719) );
  NAND2_X1 U35450 ( .A1(n3902), .A2(n2719), .ZN(n2735) );
  XOR2_X1 U35460 ( .A(n2733), .B(REG1_REG_3__SCAN_IN), .Z(n2721) );
  NOR2_X1 U35470 ( .A1(n2849), .A2(n2794), .ZN(n3857) );
  INV_X1 U35480 ( .A(n3889), .ZN(n4336) );
  XNOR2_X1 U35490 ( .A(n3889), .B(REG2_REG_1__SCAN_IN), .ZN(n3888) );
  MUX2_X1 U35500 ( .A(REG2_REG_2__SCAN_IN), .B(n2344), .S(n3897), .Z(n3904) );
  NOR2_X1 U35510 ( .A1(n3905), .A2(n3904), .ZN(n3903) );
  XNOR2_X1 U35520 ( .A(n2729), .B(n2734), .ZN(n2730) );
  XNOR2_X1 U35530 ( .A(n2730), .B(REG2_REG_3__SCAN_IN), .ZN(n2720) );
  AOI22_X1 U35540 ( .A1(n4427), .A2(n2721), .B1(n4439), .B2(n2720), .ZN(n2723)
         );
  AOI22_X1 U35550 ( .A1(n4434), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n2722) );
  OAI211_X1 U35560 ( .C1(n2734), .C2(n4442), .A(n2723), .B(n2722), .ZN(U3243)
         );
  INV_X1 U35570 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n4572) );
  INV_X1 U35580 ( .A(REG2_REG_30__SCAN_IN), .ZN(n2727) );
  NAND2_X1 U35590 ( .A1(n2352), .A2(REG0_REG_30__SCAN_IN), .ZN(n2726) );
  INV_X1 U35600 ( .A(REG1_REG_30__SCAN_IN), .ZN(n2724) );
  OAI211_X1 U35610 ( .C1(n2371), .C2(n2727), .A(n2726), .B(n2725), .ZN(n3980)
         );
  NAND2_X1 U35620 ( .A1(n3980), .A2(U4043), .ZN(n2728) );
  OAI21_X1 U35630 ( .B1(U4043), .B2(n4572), .A(n2728), .ZN(U3580) );
  INV_X1 U35640 ( .A(n2807), .ZN(n4333) );
  OAI22_X1 U35650 ( .A1(n2730), .A2(n3180), .B1(n2729), .B2(n2734), .ZN(n2732)
         );
  INV_X1 U35660 ( .A(n2731), .ZN(n2779) );
  MUX2_X1 U35670 ( .A(REG2_REG_5__SCAN_IN), .B(n2383), .S(n2807), .Z(n2800) );
  XOR2_X1 U35680 ( .A(n2759), .B(n2760), .Z(n2762) );
  XNOR2_X1 U35690 ( .A(n2762), .B(REG2_REG_6__SCAN_IN), .ZN(n2747) );
  NAND2_X1 U35700 ( .A1(n2733), .A2(REG1_REG_3__SCAN_IN), .ZN(n2737) );
  INV_X1 U35710 ( .A(n2734), .ZN(n4334) );
  NAND2_X1 U35720 ( .A1(n2735), .A2(n4334), .ZN(n2736) );
  INV_X1 U35730 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2738) );
  NAND2_X1 U35740 ( .A1(n2739), .A2(n2779), .ZN(n2740) );
  INV_X1 U35750 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2741) );
  MUX2_X1 U35760 ( .A(n2741), .B(REG1_REG_5__SCAN_IN), .S(n2807), .Z(n2804) );
  NAND2_X1 U35770 ( .A1(n2803), .A2(n2804), .ZN(n2802) );
  NAND2_X1 U35780 ( .A1(n4333), .A2(REG1_REG_5__SCAN_IN), .ZN(n2742) );
  XOR2_X1 U35790 ( .A(n2764), .B(REG1_REG_6__SCAN_IN), .Z(n2745) );
  NOR2_X1 U35800 ( .A1(STATE_REG_SCAN_IN), .A2(n2397), .ZN(n2966) );
  AOI21_X1 U35810 ( .B1(n4434), .B2(ADDR_REG_6__SCAN_IN), .A(n2966), .ZN(n2743) );
  OAI21_X1 U3582 ( .B1(n4442), .B2(n2759), .A(n2743), .ZN(n2744) );
  AOI21_X1 U3583 ( .B1(n4427), .B2(n2745), .A(n2744), .ZN(n2746) );
  OAI21_X1 U3584 ( .B1(n2747), .B2(n4398), .A(n2746), .ZN(U3246) );
  INV_X1 U3585 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n4567) );
  NAND2_X1 U3586 ( .A1(n2854), .A2(U4043), .ZN(n2748) );
  OAI21_X1 U3587 ( .B1(U4043), .B2(n4567), .A(n2748), .ZN(U3551) );
  INV_X1 U3588 ( .A(n2749), .ZN(n2754) );
  OAI21_X1 U3589 ( .B1(n4326), .B2(REG1_REG_0__SCAN_IN), .A(n2795), .ZN(n2751)
         );
  NAND2_X1 U3590 ( .A1(n4326), .A2(n2335), .ZN(n2750) );
  NAND2_X1 U3591 ( .A1(n4337), .A2(n2750), .ZN(n2796) );
  MUX2_X1 U3592 ( .A(n2751), .B(n2795), .S(n2796), .Z(n2753) );
  OAI22_X1 U3593 ( .A1(n2754), .A2(n2753), .B1(STATE_REG_SCAN_IN), .B2(n2752), 
        .ZN(n2756) );
  NOR3_X1 U3594 ( .A1(n4430), .A2(REG1_REG_0__SCAN_IN), .A3(n2795), .ZN(n2755)
         );
  AOI211_X1 U3595 ( .C1(n4434), .C2(ADDR_REG_0__SCAN_IN), .A(n2756), .B(n2755), 
        .ZN(n2757) );
  INV_X1 U3596 ( .A(n2757), .ZN(U3240) );
  INV_X1 U3597 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n4570) );
  NAND2_X1 U3598 ( .A1(n4110), .A2(U4043), .ZN(n2758) );
  OAI21_X1 U3599 ( .B1(U4043), .B2(n4570), .A(n2758), .ZN(U3572) );
  INV_X1 U3600 ( .A(n2759), .ZN(n2765) );
  INV_X1 U3601 ( .A(n2760), .ZN(n2761) );
  AOI22_X1 U3602 ( .A1(n2762), .A2(REG2_REG_6__SCAN_IN), .B1(n2765), .B2(n2761), .ZN(n2813) );
  MUX2_X1 U3603 ( .A(REG2_REG_7__SCAN_IN), .B(n2409), .S(n4331), .Z(n2812) );
  OAI21_X1 U3604 ( .B1(n2409), .B2(n4331), .A(n2816), .ZN(n3927) );
  XNOR2_X1 U3605 ( .A(n3927), .B(n3928), .ZN(n3926) );
  XNOR2_X1 U3606 ( .A(n3926), .B(REG2_REG_8__SCAN_IN), .ZN(n2777) );
  AND2_X1 U3607 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3013) );
  NOR2_X1 U3608 ( .A1(n4442), .A2(n3928), .ZN(n2763) );
  AOI211_X1 U3609 ( .C1(n4434), .C2(ADDR_REG_8__SCAN_IN), .A(n3013), .B(n2763), 
        .ZN(n2776) );
  NAND2_X1 U3610 ( .A1(n2764), .A2(REG1_REG_6__SCAN_IN), .ZN(n2768) );
  NAND2_X1 U3611 ( .A1(n2766), .A2(n2765), .ZN(n2767) );
  NOR2_X1 U3612 ( .A1(n4331), .A2(n2770), .ZN(n2769) );
  NAND2_X1 U3613 ( .A1(n4331), .A2(n2770), .ZN(n2771) );
  INV_X1 U3614 ( .A(n2773), .ZN(n2774) );
  INV_X1 U3615 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2772) );
  OAI211_X1 U3616 ( .C1(n2774), .C2(REG1_REG_8__SCAN_IN), .A(n3911), .B(n4427), 
        .ZN(n2775) );
  OAI211_X1 U3617 ( .C1(n2777), .C2(n4398), .A(n2776), .B(n2775), .ZN(U3248)
         );
  XNOR2_X1 U3618 ( .A(n2778), .B(REG1_REG_4__SCAN_IN), .ZN(n2786) );
  INV_X1 U3619 ( .A(ADDR_REG_4__SCAN_IN), .ZN(n4560) );
  INV_X1 U3620 ( .A(n4434), .ZN(n2781) );
  NAND2_X1 U3621 ( .A1(n4403), .A2(n2779), .ZN(n2780) );
  NAND2_X1 U3622 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n2936) );
  OAI211_X1 U3623 ( .C1(n4560), .C2(n2781), .A(n2780), .B(n2936), .ZN(n2785)
         );
  XNOR2_X1 U3624 ( .A(n2782), .B(REG2_REG_4__SCAN_IN), .ZN(n2783) );
  NOR2_X1 U3625 ( .A1(n4398), .A2(n2783), .ZN(n2784) );
  AOI211_X1 U3626 ( .C1(n4427), .C2(n2786), .A(n2785), .B(n2784), .ZN(n2799)
         );
  AND2_X2 U3627 ( .A1(n2787), .A2(n3026), .ZN(n2902) );
  NAND2_X1 U3628 ( .A1(n3884), .A2(n2902), .ZN(n2790) );
  OR2_X1 U3629 ( .A1(n2821), .A2(n2958), .ZN(n2862) );
  OR2_X1 U3630 ( .A1(n2931), .A2(n3891), .ZN(n2788) );
  AND2_X1 U3631 ( .A1(n2862), .A2(n2788), .ZN(n2789) );
  NAND2_X1 U3632 ( .A1(n2790), .A2(n2789), .ZN(n2861) );
  NAND2_X1 U3633 ( .A1(n2913), .A2(n3884), .ZN(n2793) );
  INV_X1 U3634 ( .A(n2931), .ZN(n2791) );
  NAND2_X1 U3635 ( .A1(n2793), .A2(n2792), .ZN(n2860) );
  XNOR2_X1 U3636 ( .A(n2861), .B(n2860), .ZN(n2847) );
  NAND3_X1 U3637 ( .A1(n2847), .A2(n4337), .A3(n2794), .ZN(n2798) );
  NOR2_X1 U3638 ( .A1(n2795), .A2(n2335), .ZN(n3887) );
  AOI22_X1 U3639 ( .A1(n3887), .A2(n3857), .B1(n2796), .B2(n2795), .ZN(n2797)
         );
  NAND3_X1 U3640 ( .A1(n2798), .A2(U4043), .A3(n2797), .ZN(n3908) );
  NAND2_X1 U3641 ( .A1(n2799), .A2(n3908), .ZN(U3244) );
  AOI211_X1 U3642 ( .C1(n2801), .C2(n2800), .A(n2060), .B(n4398), .ZN(n2809)
         );
  AND2_X1 U3643 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3627) );
  AOI21_X1 U3644 ( .B1(n4434), .B2(ADDR_REG_5__SCAN_IN), .A(n3627), .ZN(n2806)
         );
  OAI211_X1 U3645 ( .C1(n2804), .C2(n2803), .A(n4427), .B(n2802), .ZN(n2805)
         );
  OAI211_X1 U3646 ( .C1(n4442), .C2(n2807), .A(n2806), .B(n2805), .ZN(n2808)
         );
  OR2_X1 U3647 ( .A1(n2809), .A2(n2808), .ZN(U3245) );
  XOR2_X1 U3648 ( .A(n2770), .B(n4331), .Z(n2810) );
  XNOR2_X1 U3649 ( .A(n2811), .B(n2810), .ZN(n2819) );
  AOI21_X1 U3650 ( .B1(n2813), .B2(n2812), .A(n4398), .ZN(n2817) );
  AND2_X1 U3651 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n2983) );
  AOI21_X1 U3652 ( .B1(n4434), .B2(ADDR_REG_7__SCAN_IN), .A(n2983), .ZN(n2814)
         );
  OAI21_X1 U3653 ( .B1(n4442), .B2(n4331), .A(n2814), .ZN(n2815) );
  AOI21_X1 U3654 ( .B1(n2817), .B2(n2816), .A(n2815), .ZN(n2818) );
  OAI21_X1 U3655 ( .B1(n4430), .B2(n2819), .A(n2818), .ZN(U3247) );
  INV_X1 U3656 ( .A(n4484), .ZN(n4495) );
  NAND2_X1 U3657 ( .A1(n3884), .A2(n2821), .ZN(n3745) );
  NAND2_X1 U3658 ( .A1(n3066), .A2(n3745), .ZN(n4454) );
  INV_X1 U3659 ( .A(n2820), .ZN(n2831) );
  NOR2_X1 U3660 ( .A1(n2821), .A2(n2831), .ZN(n4452) );
  INV_X1 U3661 ( .A(n4135), .ZN(n3268) );
  OAI21_X1 U3662 ( .B1(n3268), .B2(n4196), .A(n4454), .ZN(n2822) );
  OAI21_X1 U3663 ( .B1(n2141), .B2(n4090), .A(n2822), .ZN(n4450) );
  AOI211_X1 U3664 ( .C1(n4495), .C2(n4454), .A(n4452), .B(n4450), .ZN(n4478)
         );
  NAND2_X1 U3665 ( .A1(n4522), .A2(REG1_REG_0__SCAN_IN), .ZN(n2823) );
  OAI21_X1 U3666 ( .B1(n4478), .B2(n4522), .A(n2823), .ZN(U3518) );
  AND2_X1 U3667 ( .A1(n2824), .A2(D_REG_1__SCAN_IN), .ZN(n2825) );
  INV_X1 U3668 ( .A(n2836), .ZN(n2832) );
  OAI211_X1 U3669 ( .C1(n2838), .C2(n2831), .A(n4198), .B(n2830), .ZN(n2841)
         );
  NOR2_X1 U3670 ( .A1(n2832), .A2(n2841), .ZN(n2833) );
  AND2_X1 U3671 ( .A1(n2836), .A2(n4227), .ZN(n2834) );
  NAND2_X1 U3672 ( .A1(n2851), .A2(n2834), .ZN(n2837) );
  INV_X2 U3673 ( .A(n2902), .ZN(n2952) );
  NAND2_X1 U3674 ( .A1(n4328), .A2(n2838), .ZN(n2856) );
  NOR2_X1 U3675 ( .A1(n3862), .A2(n4337), .ZN(n2839) );
  AOI22_X1 U3676 ( .A1(n3062), .A2(n3640), .B1(n3696), .B2(n2854), .ZN(n2846)
         );
  INV_X1 U3677 ( .A(n2851), .ZN(n2843) );
  INV_X1 U3678 ( .A(n3862), .ZN(n2840) );
  NAND2_X1 U3679 ( .A1(n2843), .A2(n2840), .ZN(n2934) );
  NAND2_X1 U3680 ( .A1(n2841), .A2(n4198), .ZN(n2842) );
  NAND2_X1 U3681 ( .A1(n2843), .A2(n2842), .ZN(n2932) );
  INV_X1 U3682 ( .A(n2844), .ZN(n3022) );
  NAND3_X1 U3683 ( .A1(n2934), .A2(n2932), .A3(n3022), .ZN(n2885) );
  INV_X1 U3684 ( .A(n2885), .ZN(n2869) );
  OR2_X1 U3685 ( .A1(n2869), .A2(n2752), .ZN(n2845) );
  OAI211_X1 U3686 ( .C1(n2847), .C2(n3688), .A(n2846), .B(n2845), .ZN(U3229)
         );
  INV_X1 U3687 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n4569) );
  NAND2_X1 U3688 ( .A1(n4036), .A2(U4043), .ZN(n2848) );
  OAI21_X1 U3689 ( .B1(U4043), .B2(n4569), .A(n2848), .ZN(U3576) );
  INV_X1 U3690 ( .A(n3884), .ZN(n2852) );
  NOR2_X1 U3691 ( .A1(n3862), .A2(n2849), .ZN(n2850) );
  OAI22_X1 U3692 ( .A1(n2852), .A2(n3681), .B1(n3683), .B2(n3173), .ZN(n2853)
         );
  AOI21_X1 U3693 ( .B1(n3063), .B2(n3640), .A(n2853), .ZN(n2868) );
  NAND2_X1 U3694 ( .A1(n2854), .A2(n2902), .ZN(n2855) );
  NOR2_X1 U3695 ( .A1(n2952), .A2(n3068), .ZN(n2859) );
  AOI21_X1 U3696 ( .B1(n2913), .B2(n2854), .A(n2859), .ZN(n2874) );
  XNOR2_X1 U3697 ( .A(n2876), .B(n2874), .ZN(n2866) );
  NAND2_X1 U3698 ( .A1(n2861), .A2(n2860), .ZN(n2864) );
  INV_X4 U3699 ( .A(n3547), .ZN(n3533) );
  NAND2_X1 U3700 ( .A1(n2862), .A2(n3533), .ZN(n2863) );
  NAND2_X1 U3701 ( .A1(n2864), .A2(n2863), .ZN(n2865) );
  NAND2_X1 U3702 ( .A1(n2866), .A2(n2865), .ZN(n2878) );
  OAI211_X1 U3703 ( .C1(n2866), .C2(n2865), .A(n2878), .B(n3704), .ZN(n2867)
         );
  OAI211_X1 U3704 ( .C1(n2869), .C2(n2328), .A(n2868), .B(n2867), .ZN(U3219)
         );
  NAND2_X1 U3705 ( .A1(n3882), .A2(n2902), .ZN(n2871) );
  OR2_X1 U3706 ( .A1(n2899), .A2(n2958), .ZN(n2870) );
  NAND2_X1 U3707 ( .A1(n2871), .A2(n2870), .ZN(n2872) );
  XNOR2_X1 U3708 ( .A(n2872), .B(n3533), .ZN(n2916) );
  NOR2_X1 U3709 ( .A1(n2952), .A2(n2899), .ZN(n2873) );
  AOI21_X1 U3710 ( .B1(n2913), .B2(n3882), .A(n2873), .ZN(n2915) );
  XNOR2_X1 U3711 ( .A(n2916), .B(n2915), .ZN(n2882) );
  INV_X1 U3712 ( .A(n2874), .ZN(n2875) );
  NAND2_X1 U3713 ( .A1(n2876), .A2(n2875), .ZN(n2877) );
  NAND2_X1 U3714 ( .A1(n2878), .A2(n2877), .ZN(n2879) );
  INV_X1 U3715 ( .A(n2879), .ZN(n2881) );
  INV_X1 U3716 ( .A(n2882), .ZN(n2880) );
  NAND2_X1 U3717 ( .A1(n2881), .A2(n2880), .ZN(n2925) );
  INV_X1 U3718 ( .A(n2925), .ZN(n2907) );
  AOI21_X1 U3719 ( .B1(n2882), .B2(n2879), .A(n2907), .ZN(n2887) );
  AOI22_X1 U3720 ( .A1(n3696), .A2(n3881), .B1(n3697), .B2(n2854), .ZN(n2883)
         );
  OAI21_X1 U3721 ( .B1(n3680), .B2(n2899), .A(n2883), .ZN(n2884) );
  AOI21_X1 U3722 ( .B1(REG3_REG_2__SCAN_IN), .B2(n2885), .A(n2884), .ZN(n2886)
         );
  OAI21_X1 U3723 ( .B1(n2887), .B2(n3688), .A(n2886), .ZN(U3234) );
  NAND2_X1 U3724 ( .A1(n2889), .A2(n2888), .ZN(n3169) );
  OAI21_X1 U3725 ( .B1(n2889), .B2(n2888), .A(n3169), .ZN(n4444) );
  INV_X1 U3726 ( .A(n4444), .ZN(n2898) );
  OAI21_X1 U3727 ( .B1(n3835), .B2(n2891), .A(n2890), .ZN(n2892) );
  NAND2_X1 U3728 ( .A1(n2892), .A2(n4196), .ZN(n2895) );
  INV_X1 U3729 ( .A(n2899), .ZN(n2893) );
  AOI22_X1 U3730 ( .A1(n2854), .A2(n4155), .B1(n2893), .B2(n4227), .ZN(n2894)
         );
  OAI211_X1 U3731 ( .C1(n2896), .C2(n4090), .A(n2895), .B(n2894), .ZN(n2897)
         );
  AOI21_X1 U3732 ( .B1(n3268), .B2(n4444), .A(n2897), .ZN(n4449) );
  OAI21_X1 U3733 ( .B1(n2898), .B2(n4484), .A(n4449), .ZN(n3043) );
  OAI21_X1 U3734 ( .B1(n3061), .B2(n2899), .A(n3178), .ZN(n4443) );
  OAI22_X1 U3735 ( .A1(n4275), .A2(n4443), .B1(n4524), .B2(n2713), .ZN(n2900)
         );
  AOI21_X1 U3736 ( .B1(n3043), .B2(n4524), .A(n2900), .ZN(n2901) );
  INV_X1 U3737 ( .A(n2901), .ZN(U3520) );
  OR2_X1 U3738 ( .A1(n3037), .A2(n2958), .ZN(n2904) );
  NAND2_X1 U3739 ( .A1(n3880), .A2(n2902), .ZN(n2903) );
  NAND2_X1 U3740 ( .A1(n2904), .A2(n2903), .ZN(n2905) );
  NOR2_X1 U3741 ( .A1(n2952), .A2(n3037), .ZN(n2906) );
  AOI21_X1 U3742 ( .B1(n2913), .B2(n3880), .A(n2906), .ZN(n2944) );
  XNOR2_X1 U3743 ( .A(n2943), .B(n2944), .ZN(n2922) );
  NAND2_X1 U3744 ( .A1(n2902), .A2(n3881), .ZN(n2909) );
  OR2_X1 U3745 ( .A1(n2911), .A2(n2958), .ZN(n2908) );
  NAND2_X1 U3746 ( .A1(n2909), .A2(n2908), .ZN(n2910) );
  XNOR2_X1 U3747 ( .A(n2910), .B(n3547), .ZN(n2918) );
  INV_X1 U3748 ( .A(n2918), .ZN(n2914) );
  NOR2_X1 U3749 ( .A1(n2952), .A2(n2911), .ZN(n2912) );
  AOI21_X1 U3750 ( .B1(n2913), .B2(n3881), .A(n2912), .ZN(n2917) );
  NAND2_X1 U3751 ( .A1(n2916), .A2(n2915), .ZN(n2989) );
  AND2_X1 U3752 ( .A1(n2919), .A2(n2989), .ZN(n2923) );
  NAND2_X1 U3753 ( .A1(n2925), .A2(n2923), .ZN(n2921) );
  XNOR2_X1 U3754 ( .A(n2918), .B(n2917), .ZN(n2991) );
  INV_X1 U3755 ( .A(n2991), .ZN(n2920) );
  AND2_X1 U3756 ( .A1(n2921), .A2(n2926), .ZN(n2928) );
  INV_X1 U3757 ( .A(n2922), .ZN(n2924) );
  NAND2_X1 U3758 ( .A1(n2925), .A2(n2024), .ZN(n2948) );
  OR2_X1 U3759 ( .A1(n2926), .A2(n2922), .ZN(n2947) );
  NAND2_X1 U3760 ( .A1(n2948), .A2(n2947), .ZN(n2927) );
  AOI211_X1 U3761 ( .C1(n2922), .C2(n2928), .A(n3688), .B(n2927), .ZN(n2942)
         );
  NAND4_X1 U3762 ( .A1(n2932), .A2(n2931), .A3(n2930), .A4(n2929), .ZN(n2933)
         );
  NAND2_X1 U3763 ( .A1(n2933), .A2(STATE_REG_SCAN_IN), .ZN(n2935) );
  INV_X1 U3764 ( .A(n2936), .ZN(n2937) );
  AOI21_X1 U3765 ( .B1(n3697), .B2(n3881), .A(n2937), .ZN(n2940) );
  AOI22_X1 U3766 ( .A1(n2938), .A2(n3640), .B1(n3696), .B2(n3033), .ZN(n2939)
         );
  OAI211_X1 U3767 ( .C1(n3702), .C2(n3038), .A(n2940), .B(n2939), .ZN(n2941)
         );
  OR2_X1 U3768 ( .A1(n2942), .A2(n2941), .ZN(U3227) );
  INV_X1 U3769 ( .A(n2943), .ZN(n2946) );
  INV_X1 U3770 ( .A(n2944), .ZN(n2945) );
  NAND2_X1 U3771 ( .A1(n3033), .A2(n2978), .ZN(n2950) );
  OR2_X1 U3772 ( .A1(n3120), .A2(n3538), .ZN(n2949) );
  NAND2_X1 U3773 ( .A1(n2950), .A2(n2949), .ZN(n2951) );
  XNOR2_X1 U3774 ( .A(n2951), .B(n3547), .ZN(n2956) );
  NOR2_X1 U3775 ( .A1(n3550), .A2(n3120), .ZN(n2953) );
  AOI21_X1 U3776 ( .B1(n2005), .B2(n3033), .A(n2953), .ZN(n2954) );
  XNOR2_X1 U3777 ( .A(n2956), .B(n2954), .ZN(n3625) );
  NAND2_X1 U3778 ( .A1(n3626), .A2(n3625), .ZN(n3624) );
  INV_X1 U3779 ( .A(n2954), .ZN(n2955) );
  NAND2_X1 U3780 ( .A1(n2956), .A2(n2955), .ZN(n2957) );
  NAND2_X1 U3781 ( .A1(n3879), .A2(n2978), .ZN(n2960) );
  OR2_X1 U3782 ( .A1(n2962), .A2(n3538), .ZN(n2959) );
  NAND2_X1 U3783 ( .A1(n2960), .A2(n2959), .ZN(n2961) );
  XNOR2_X1 U3784 ( .A(n2961), .B(n3547), .ZN(n2973) );
  NAND2_X1 U3785 ( .A1(n2005), .A2(n3879), .ZN(n2964) );
  OR2_X1 U3786 ( .A1(n2962), .A2(n3546), .ZN(n2963) );
  NAND2_X1 U3787 ( .A1(n2964), .A2(n2963), .ZN(n2974) );
  XNOR2_X1 U3788 ( .A(n2973), .B(n2974), .ZN(n2965) );
  XNOR2_X1 U3789 ( .A(n2975), .B(n2965), .ZN(n2970) );
  AOI21_X1 U3790 ( .B1(n3697), .B2(n3033), .A(n2966), .ZN(n2968) );
  AOI22_X1 U3791 ( .A1(n3053), .A2(n3640), .B1(n3696), .B2(n3878), .ZN(n2967)
         );
  OAI211_X1 U3792 ( .C1(n3702), .C2(n3143), .A(n2968), .B(n2967), .ZN(n2969)
         );
  AOI21_X1 U3793 ( .B1(n2970), .B2(n3704), .A(n2969), .ZN(n2971) );
  INV_X1 U3794 ( .A(n2971), .ZN(U3236) );
  INV_X1 U3795 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n4573) );
  NAND2_X1 U3796 ( .A1(n4019), .A2(U4043), .ZN(n2972) );
  OAI21_X1 U3797 ( .B1(U4043), .B2(n4573), .A(n2972), .ZN(U3577) );
  OAI21_X1 U3798 ( .B1(n2975), .B2(n2974), .A(n2973), .ZN(n2977) );
  NAND2_X1 U3799 ( .A1(n2975), .A2(n2974), .ZN(n2976) );
  NAND2_X1 U3800 ( .A1(n3878), .A2(n2978), .ZN(n2980) );
  OR2_X1 U3801 ( .A1(n3151), .A2(n3538), .ZN(n2979) );
  NAND2_X1 U3802 ( .A1(n2980), .A2(n2979), .ZN(n2981) );
  XNOR2_X1 U3803 ( .A(n2981), .B(n3547), .ZN(n3001) );
  NOR2_X1 U3804 ( .A1(n3550), .A2(n3151), .ZN(n2982) );
  AOI21_X1 U3805 ( .B1(n2005), .B2(n3878), .A(n2982), .ZN(n2999) );
  XNOR2_X1 U3806 ( .A(n3001), .B(n2999), .ZN(n2997) );
  XOR2_X1 U3807 ( .A(n2998), .B(n2997), .Z(n2987) );
  AOI21_X1 U3808 ( .B1(n3696), .B2(n3877), .A(n2983), .ZN(n2985) );
  AOI22_X1 U3809 ( .A1(n3156), .A2(n3640), .B1(n3697), .B2(n3879), .ZN(n2984)
         );
  OAI211_X1 U3810 ( .C1(n3702), .C2(n3161), .A(n2985), .B(n2984), .ZN(n2986)
         );
  AOI21_X1 U3811 ( .B1(n2987), .B2(n3704), .A(n2986), .ZN(n2988) );
  INV_X1 U3812 ( .A(n2988), .ZN(U3210) );
  NAND2_X1 U3813 ( .A1(n2925), .A2(n2989), .ZN(n2990) );
  XOR2_X1 U3814 ( .A(n2991), .B(n2990), .Z(n2996) );
  INV_X1 U3815 ( .A(n3880), .ZN(n2992) );
  OAI22_X1 U3816 ( .A1(n3173), .A2(n3681), .B1(n3683), .B2(n2992), .ZN(n2994)
         );
  MUX2_X1 U3817 ( .A(n3686), .B(U3149), .S(REG3_REG_3__SCAN_IN), .Z(n2993) );
  AOI211_X1 U3818 ( .C1(n3179), .C2(n3640), .A(n2994), .B(n2993), .ZN(n2995)
         );
  OAI21_X1 U3819 ( .B1(n3688), .B2(n2996), .A(n2995), .ZN(U3215) );
  INV_X1 U3820 ( .A(n2999), .ZN(n3000) );
  NAND2_X1 U3821 ( .A1(n3001), .A2(n3000), .ZN(n3002) );
  NAND2_X1 U3822 ( .A1(n3877), .A2(n2978), .ZN(n3004) );
  OR2_X1 U3823 ( .A1(n3129), .A2(n3538), .ZN(n3003) );
  NAND2_X1 U3824 ( .A1(n3004), .A2(n3003), .ZN(n3005) );
  XNOR2_X1 U3825 ( .A(n3005), .B(n3547), .ZN(n3008) );
  NAND2_X1 U3826 ( .A1(n2005), .A2(n3877), .ZN(n3007) );
  OR2_X1 U3827 ( .A1(n3129), .A2(n3550), .ZN(n3006) );
  NAND2_X1 U3828 ( .A1(n3007), .A2(n3006), .ZN(n3009) );
  AND2_X1 U3829 ( .A1(n3008), .A2(n3009), .ZN(n3079) );
  INV_X1 U3830 ( .A(n3008), .ZN(n3011) );
  INV_X1 U3831 ( .A(n3009), .ZN(n3010) );
  NAND2_X1 U3832 ( .A1(n3011), .A2(n3010), .ZN(n3078) );
  NAND2_X1 U3833 ( .A1(n2209), .A2(n3078), .ZN(n3012) );
  XNOR2_X1 U3834 ( .A(n3080), .B(n3012), .ZN(n3017) );
  AOI21_X1 U3835 ( .B1(n3697), .B2(n3878), .A(n3013), .ZN(n3015) );
  AOI22_X1 U3836 ( .A1(n3135), .A2(n3640), .B1(n3696), .B2(n3876), .ZN(n3014)
         );
  OAI211_X1 U3837 ( .C1(n3702), .C2(n3186), .A(n3015), .B(n3014), .ZN(n3016)
         );
  AOI21_X1 U3838 ( .B1(n3017), .B2(n3704), .A(n3016), .ZN(n3018) );
  INV_X1 U3839 ( .A(n3018), .ZN(U3218) );
  NAND2_X1 U3840 ( .A1(n3019), .A2(n3836), .ZN(n3020) );
  NAND2_X1 U3841 ( .A1(n3021), .A2(n3020), .ZN(n4491) );
  NAND3_X1 U3842 ( .A1(n3024), .A2(n3023), .A3(n3022), .ZN(n3025) );
  NAND2_X1 U3843 ( .A1(n3026), .A2(n2611), .ZN(n3103) );
  INV_X1 U3844 ( .A(n3103), .ZN(n3027) );
  NAND2_X1 U3845 ( .A1(n4188), .A2(n3027), .ZN(n4144) );
  XNOR2_X1 U3846 ( .A(n3029), .B(n3028), .ZN(n3035) );
  NAND2_X1 U3847 ( .A1(n3881), .A2(n4155), .ZN(n3030) );
  OAI21_X1 U3848 ( .B1(n4198), .B2(n3037), .A(n3030), .ZN(n3032) );
  NOR2_X1 U3849 ( .A1(n4491), .A2(n4135), .ZN(n3031) );
  AOI211_X1 U3850 ( .C1(n4200), .C2(n3033), .A(n3032), .B(n3031), .ZN(n3034)
         );
  OAI21_X1 U3851 ( .B1(n4158), .B2(n3035), .A(n3034), .ZN(n4493) );
  INV_X1 U3852 ( .A(n3121), .ZN(n3036) );
  OAI211_X1 U3853 ( .C1(n3177), .C2(n3037), .A(n3036), .B(n4489), .ZN(n4492)
         );
  OAI22_X1 U3854 ( .A1(n4492), .A2(n2611), .B1(n4211), .B2(n3038), .ZN(n3039)
         );
  OAI21_X1 U3855 ( .B1(n4493), .B2(n3039), .A(n4136), .ZN(n3041) );
  NAND2_X1 U3856 ( .A1(n4458), .A2(REG2_REG_4__SCAN_IN), .ZN(n3040) );
  OAI211_X1 U3857 ( .C1(n4491), .C2(n4144), .A(n3041), .B(n3040), .ZN(U3286)
         );
  OAI22_X1 U3858 ( .A1(n4320), .A2(n4443), .B1(n4516), .B2(n2343), .ZN(n3042)
         );
  AOI21_X1 U3859 ( .B1(n3043), .B2(n4516), .A(n3042), .ZN(n3044) );
  INV_X1 U3860 ( .A(n3044), .ZN(U3471) );
  INV_X1 U3861 ( .A(n3045), .ZN(n3759) );
  OR2_X1 U3862 ( .A1(n3759), .A2(n3762), .ZN(n3047) );
  XNOR2_X1 U3863 ( .A(n3046), .B(n3047), .ZN(n3144) );
  INV_X1 U3864 ( .A(n3047), .ZN(n3834) );
  XNOR2_X1 U3865 ( .A(n3048), .B(n3834), .ZN(n3052) );
  AOI22_X1 U3866 ( .A1(n3878), .A2(n4200), .B1(n3053), .B2(n4227), .ZN(n3049)
         );
  OAI21_X1 U3867 ( .B1(n3050), .B2(n4204), .A(n3049), .ZN(n3051) );
  AOI21_X1 U3868 ( .B1(n3052), .B2(n4196), .A(n3051), .ZN(n3149) );
  OAI21_X1 U3869 ( .B1(n4501), .B2(n3144), .A(n3149), .ZN(n3059) );
  NAND2_X1 U3870 ( .A1(n3119), .A2(n3053), .ZN(n3054) );
  NAND2_X1 U3871 ( .A1(n3157), .A2(n3054), .ZN(n3142) );
  INV_X1 U3872 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3055) );
  OAI22_X1 U3873 ( .A1(n4275), .A2(n3142), .B1(n4524), .B2(n3055), .ZN(n3056)
         );
  AOI21_X1 U3874 ( .B1(n3059), .B2(n4524), .A(n3056), .ZN(n3057) );
  INV_X1 U3875 ( .A(n3057), .ZN(U3524) );
  OAI22_X1 U3876 ( .A1(n4320), .A2(n3142), .B1(n4516), .B2(n2396), .ZN(n3058)
         );
  AOI21_X1 U3877 ( .B1(n3059), .B2(n4516), .A(n3058), .ZN(n3060) );
  INV_X1 U3878 ( .A(n3060), .ZN(U3479) );
  NAND2_X1 U3879 ( .A1(n4188), .A2(n2838), .ZN(n4183) );
  INV_X1 U3880 ( .A(n3061), .ZN(n3065) );
  NAND2_X1 U3881 ( .A1(n3063), .A2(n3062), .ZN(n3064) );
  NAND2_X1 U3882 ( .A1(n3065), .A2(n3064), .ZN(n4479) );
  INV_X1 U3883 ( .A(n3066), .ZN(n3747) );
  XNOR2_X1 U3884 ( .A(n2612), .B(n3747), .ZN(n3074) );
  NAND2_X1 U3885 ( .A1(n3882), .A2(n4200), .ZN(n3067) );
  OAI21_X1 U3886 ( .B1(n4198), .B2(n3068), .A(n3067), .ZN(n3072) );
  OAI21_X1 U3887 ( .B1(n2612), .B2(n3070), .A(n3069), .ZN(n4480) );
  NOR2_X1 U3888 ( .A1(n4480), .A2(n4135), .ZN(n3071) );
  AOI211_X1 U3889 ( .C1(n4155), .C2(n3884), .A(n3072), .B(n3071), .ZN(n3073)
         );
  OAI21_X1 U3890 ( .B1(n4158), .B2(n3074), .A(n3073), .ZN(n4482) );
  AOI22_X1 U3891 ( .A1(n4458), .A2(REG2_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(n4453), .ZN(n3075) );
  OAI21_X1 U3892 ( .B1(n4144), .B2(n4480), .A(n3075), .ZN(n3076) );
  AOI21_X1 U3893 ( .B1(n4482), .B2(n4188), .A(n3076), .ZN(n3077) );
  OAI21_X1 U3894 ( .B1(n4210), .B2(n4479), .A(n3077), .ZN(U3289) );
  NAND2_X1 U3895 ( .A1(n3876), .A2(n2978), .ZN(n3082) );
  OR2_X1 U3896 ( .A1(n3106), .A2(n3538), .ZN(n3081) );
  NAND2_X1 U3897 ( .A1(n3082), .A2(n3081), .ZN(n3083) );
  XNOR2_X1 U3898 ( .A(n3083), .B(n3547), .ZN(n3194) );
  NOR2_X1 U3899 ( .A1(n3550), .A2(n3106), .ZN(n3084) );
  AOI21_X1 U3900 ( .B1(n2005), .B2(n3876), .A(n3084), .ZN(n3195) );
  XNOR2_X1 U3901 ( .A(n3194), .B(n3195), .ZN(n3192) );
  XNOR2_X1 U3902 ( .A(n3193), .B(n3192), .ZN(n3089) );
  AND2_X1 U3903 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4348) );
  AOI21_X1 U3904 ( .B1(n3696), .B2(n3875), .A(n4348), .ZN(n3087) );
  AOI22_X1 U3905 ( .A1(n3085), .A2(n3640), .B1(n3697), .B2(n3877), .ZN(n3086)
         );
  OAI211_X1 U3906 ( .C1(n3702), .C2(n3107), .A(n3087), .B(n3086), .ZN(n3088)
         );
  AOI21_X1 U3907 ( .B1(n3089), .B2(n3704), .A(n3088), .ZN(n3090) );
  INV_X1 U3908 ( .A(n3090), .ZN(U3228) );
  INV_X1 U3909 ( .A(n3091), .ZN(n3772) );
  AND2_X1 U3910 ( .A1(n3772), .A2(n3769), .ZN(n3817) );
  INV_X1 U3911 ( .A(n3817), .ZN(n3092) );
  XNOR2_X1 U3912 ( .A(n3093), .B(n3092), .ZN(n3097) );
  NAND2_X1 U3913 ( .A1(n3877), .A2(n4155), .ZN(n3095) );
  NAND2_X1 U3914 ( .A1(n3875), .A2(n4200), .ZN(n3094) );
  OAI211_X1 U3915 ( .C1(n4198), .C2(n3106), .A(n3095), .B(n3094), .ZN(n3096)
         );
  AOI21_X1 U3916 ( .B1(n3097), .B2(n4196), .A(n3096), .ZN(n4508) );
  OR2_X1 U3917 ( .A1(n3098), .A2(n3099), .ZN(n3101) );
  NAND2_X1 U3918 ( .A1(n3101), .A2(n3100), .ZN(n3102) );
  XNOR2_X1 U3919 ( .A(n3102), .B(n3817), .ZN(n4513) );
  NAND2_X1 U3920 ( .A1(n4135), .A2(n3103), .ZN(n3104) );
  INV_X1 U3921 ( .A(n4217), .ZN(n3412) );
  INV_X1 U3922 ( .A(n3105), .ZN(n3133) );
  OAI21_X1 U3923 ( .B1(n3133), .B2(n3106), .A(n3234), .ZN(n4509) );
  NOR2_X1 U3924 ( .A1(n4509), .A2(n4210), .ZN(n3110) );
  OAI22_X1 U3925 ( .A1(n4188), .A2(n3108), .B1(n3107), .B2(n4211), .ZN(n3109)
         );
  AOI211_X1 U3926 ( .C1(n4513), .C2(n3412), .A(n3110), .B(n3109), .ZN(n3111)
         );
  OAI21_X1 U3927 ( .B1(n4458), .B2(n4508), .A(n3111), .ZN(U3281) );
  INV_X1 U3928 ( .A(n3112), .ZN(n3756) );
  XOR2_X1 U3929 ( .A(n3833), .B(n3113), .Z(n3117) );
  NAND2_X1 U3930 ( .A1(n3880), .A2(n4155), .ZN(n3115) );
  NAND2_X1 U3931 ( .A1(n3879), .A2(n4200), .ZN(n3114) );
  OAI211_X1 U3932 ( .C1(n4198), .C2(n3120), .A(n3115), .B(n3114), .ZN(n3116)
         );
  AOI21_X1 U3933 ( .B1(n3117), .B2(n4196), .A(n3116), .ZN(n4497) );
  XNOR2_X1 U3934 ( .A(n3118), .B(n3833), .ZN(n4500) );
  OAI21_X1 U3935 ( .B1(n3121), .B2(n3120), .A(n3119), .ZN(n4498) );
  NOR2_X1 U3936 ( .A1(n4210), .A2(n4498), .ZN(n3123) );
  OAI22_X1 U3937 ( .A1(n4136), .A2(n2383), .B1(n3629), .B2(n4211), .ZN(n3122)
         );
  AOI211_X1 U3938 ( .C1(n4500), .C2(n3412), .A(n3123), .B(n3122), .ZN(n3124)
         );
  OAI21_X1 U3939 ( .B1(n4497), .B2(n4458), .A(n3124), .ZN(U3285) );
  OR2_X1 U3940 ( .A1(n3098), .A2(n3837), .ZN(n4505) );
  NAND2_X1 U3941 ( .A1(n4505), .A2(n3126), .ZN(n3127) );
  XNOR2_X1 U3942 ( .A(n3127), .B(n3815), .ZN(n3184) );
  XNOR2_X1 U3943 ( .A(n3128), .B(n3815), .ZN(n3132) );
  OAI22_X1 U3944 ( .A1(n3230), .A2(n4090), .B1(n3129), .B2(n4198), .ZN(n3130)
         );
  AOI21_X1 U3945 ( .B1(n4155), .B2(n3878), .A(n3130), .ZN(n3131) );
  OAI21_X1 U3946 ( .B1(n3132), .B2(n4158), .A(n3131), .ZN(n3185) );
  AOI21_X1 U3947 ( .B1(n3184), .B2(n4512), .A(n3185), .ZN(n3141) );
  INV_X1 U3948 ( .A(n3160), .ZN(n3134) );
  AOI21_X1 U3949 ( .B1(n3135), .B2(n3134), .A(n3133), .ZN(n3188) );
  INV_X1 U3950 ( .A(n4320), .ZN(n3137) );
  NOR2_X1 U3951 ( .A1(n4516), .A2(n2422), .ZN(n3136) );
  AOI21_X1 U3952 ( .B1(n3188), .B2(n3137), .A(n3136), .ZN(n3138) );
  OAI21_X1 U3953 ( .B1(n3141), .B2(n4514), .A(n3138), .ZN(U3483) );
  INV_X1 U3954 ( .A(n4275), .ZN(n3139) );
  AOI22_X1 U3955 ( .A1(n3188), .A2(n3139), .B1(n4522), .B2(REG1_REG_8__SCAN_IN), .ZN(n3140) );
  OAI21_X1 U3956 ( .B1(n3141), .B2(n4522), .A(n3140), .ZN(U3526) );
  INV_X1 U3957 ( .A(n3142), .ZN(n3147) );
  OAI22_X1 U3958 ( .A1(n4136), .A2(n2401), .B1(n3143), .B2(n4211), .ZN(n3146)
         );
  NOR2_X1 U3959 ( .A1(n3144), .A2(n4217), .ZN(n3145) );
  AOI211_X1 U3960 ( .C1(n3147), .C2(n4446), .A(n3146), .B(n3145), .ZN(n3148)
         );
  OAI21_X1 U3961 ( .B1(n4458), .B2(n3149), .A(n3148), .ZN(U3284) );
  XNOR2_X1 U3962 ( .A(n3150), .B(n3837), .ZN(n3155) );
  NOR2_X1 U3963 ( .A1(n4198), .A2(n3151), .ZN(n3152) );
  AOI21_X1 U3964 ( .B1(n3877), .B2(n4200), .A(n3152), .ZN(n3154) );
  NAND2_X1 U3965 ( .A1(n3879), .A2(n4155), .ZN(n3153) );
  OAI211_X1 U3966 ( .C1(n3155), .C2(n4158), .A(n3154), .B(n3153), .ZN(n4503)
         );
  INV_X1 U3967 ( .A(n4503), .ZN(n3167) );
  INV_X1 U3968 ( .A(n4183), .ZN(n3165) );
  NAND2_X1 U3969 ( .A1(n3157), .A2(n3156), .ZN(n3158) );
  NAND2_X1 U3970 ( .A1(n3158), .A2(n4489), .ZN(n3159) );
  NOR2_X1 U3971 ( .A1(n3160), .A2(n3159), .ZN(n4504) );
  OAI22_X1 U3972 ( .A1(n4188), .A2(n2409), .B1(n3161), .B2(n4211), .ZN(n3164)
         );
  INV_X1 U3973 ( .A(n4505), .ZN(n3162) );
  AND2_X1 U3974 ( .A1(n3098), .A2(n3837), .ZN(n4502) );
  NOR3_X1 U3975 ( .A1(n3162), .A2(n4502), .A3(n4217), .ZN(n3163) );
  AOI211_X1 U3976 ( .C1(n3165), .C2(n4504), .A(n3164), .B(n3163), .ZN(n3166)
         );
  OAI21_X1 U3977 ( .B1(n4458), .B2(n3167), .A(n3166), .ZN(U3283) );
  NAND2_X1 U3978 ( .A1(n3169), .A2(n3168), .ZN(n3170) );
  XNOR2_X1 U3979 ( .A(n3170), .B(n2264), .ZN(n4485) );
  XNOR2_X1 U3980 ( .A(n3171), .B(n2264), .ZN(n3175) );
  AOI22_X1 U3981 ( .A1(n3880), .A2(n4200), .B1(n4227), .B2(n3179), .ZN(n3172)
         );
  OAI21_X1 U3982 ( .B1(n3173), .B2(n4204), .A(n3172), .ZN(n3174) );
  AOI21_X1 U3983 ( .B1(n3175), .B2(n4196), .A(n3174), .ZN(n3176) );
  OAI21_X1 U3984 ( .B1(n4485), .B2(n4135), .A(n3176), .ZN(n4486) );
  NAND2_X1 U3985 ( .A1(n4486), .A2(n4136), .ZN(n3183) );
  AOI21_X1 U3986 ( .B1(n3179), .B2(n3178), .A(n3177), .ZN(n4488) );
  OAI22_X1 U3987 ( .A1(n4136), .A2(n3180), .B1(REG3_REG_3__SCAN_IN), .B2(n4211), .ZN(n3181) );
  AOI21_X1 U3988 ( .B1(n4446), .B2(n4488), .A(n3181), .ZN(n3182) );
  OAI211_X1 U3989 ( .C1(n4485), .C2(n4144), .A(n3183), .B(n3182), .ZN(U3287)
         );
  INV_X1 U3990 ( .A(n3184), .ZN(n3191) );
  NAND2_X1 U3991 ( .A1(n3185), .A2(n4136), .ZN(n3190) );
  OAI22_X1 U3992 ( .A1(n4188), .A2(n3929), .B1(n3186), .B2(n4211), .ZN(n3187)
         );
  AOI21_X1 U3993 ( .B1(n3188), .B2(n4446), .A(n3187), .ZN(n3189) );
  OAI211_X1 U3994 ( .C1(n3191), .C2(n4217), .A(n3190), .B(n3189), .ZN(U3282)
         );
  NAND2_X1 U3995 ( .A1(n3193), .A2(n3192), .ZN(n3198) );
  INV_X1 U3996 ( .A(n3194), .ZN(n3196) );
  NAND2_X1 U3997 ( .A1(n3196), .A2(n3195), .ZN(n3197) );
  NAND2_X1 U3998 ( .A1(n3198), .A2(n3197), .ZN(n3222) );
  NAND2_X1 U3999 ( .A1(n3875), .A2(n2978), .ZN(n3200) );
  OR2_X1 U4000 ( .A1(n3202), .A2(n3538), .ZN(n3199) );
  NAND2_X1 U4001 ( .A1(n3200), .A2(n3199), .ZN(n3201) );
  XNOR2_X1 U4002 ( .A(n3201), .B(n3533), .ZN(n3204) );
  NOR2_X1 U4003 ( .A1(n3546), .A2(n3202), .ZN(n3203) );
  AOI21_X1 U4004 ( .B1(n2005), .B2(n3875), .A(n3203), .ZN(n3205) );
  XNOR2_X1 U4005 ( .A(n3204), .B(n3205), .ZN(n3223) );
  INV_X1 U4006 ( .A(n3204), .ZN(n3207) );
  INV_X1 U4007 ( .A(n3205), .ZN(n3206) );
  NAND2_X1 U4008 ( .A1(n3207), .A2(n3206), .ZN(n3208) );
  NAND2_X1 U4009 ( .A1(n3874), .A2(n2978), .ZN(n3210) );
  OR2_X1 U4010 ( .A1(n3273), .A2(n3538), .ZN(n3209) );
  NAND2_X1 U4011 ( .A1(n3210), .A2(n3209), .ZN(n3211) );
  XNOR2_X1 U4012 ( .A(n3211), .B(n3547), .ZN(n3243) );
  NAND2_X1 U4013 ( .A1(n2005), .A2(n3874), .ZN(n3213) );
  OR2_X1 U4014 ( .A1(n3273), .A2(n3546), .ZN(n3212) );
  NAND2_X1 U4015 ( .A1(n3213), .A2(n3212), .ZN(n3244) );
  XNOR2_X1 U4016 ( .A(n3243), .B(n3244), .ZN(n3214) );
  XNOR2_X1 U4017 ( .A(n3245), .B(n3214), .ZN(n3220) );
  NOR2_X1 U4018 ( .A1(STATE_REG_SCAN_IN), .A2(n3215), .ZN(n4368) );
  AOI21_X1 U4019 ( .B1(n3696), .B2(n3873), .A(n4368), .ZN(n3218) );
  AOI22_X1 U4020 ( .A1(n3216), .A2(n3640), .B1(n3697), .B2(n3875), .ZN(n3217)
         );
  OAI211_X1 U4021 ( .C1(n3702), .C2(n3275), .A(n3218), .B(n3217), .ZN(n3219)
         );
  AOI21_X1 U4022 ( .B1(n3220), .B2(n3704), .A(n3219), .ZN(n3221) );
  INV_X1 U4023 ( .A(n3221), .ZN(U3233) );
  AOI211_X1 U4024 ( .C1(n3223), .C2(n3222), .A(n3688), .B(n2049), .ZN(n3227)
         );
  AND2_X1 U4025 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4358) );
  AOI21_X1 U4026 ( .B1(n3697), .B2(n3876), .A(n4358), .ZN(n3225) );
  AOI22_X1 U4027 ( .A1(n3233), .A2(n3640), .B1(n3696), .B2(n3874), .ZN(n3224)
         );
  OAI211_X1 U4028 ( .C1(n3702), .C2(n3236), .A(n3225), .B(n3224), .ZN(n3226)
         );
  OR2_X1 U4029 ( .A1(n3227), .A2(n3226), .ZN(U3214) );
  NAND2_X1 U4030 ( .A1(n3771), .A2(n3774), .ZN(n3813) );
  XOR2_X1 U4031 ( .A(n3813), .B(n3228), .Z(n3232) );
  AOI22_X1 U4032 ( .A1(n3874), .A2(n4200), .B1(n4227), .B2(n3233), .ZN(n3229)
         );
  OAI21_X1 U4033 ( .B1(n3230), .B2(n4204), .A(n3229), .ZN(n3231) );
  AOI21_X1 U4034 ( .B1(n3232), .B2(n4196), .A(n3231), .ZN(n3281) );
  NAND2_X1 U4035 ( .A1(n3234), .A2(n3233), .ZN(n3235) );
  NAND2_X1 U4036 ( .A1(n3271), .A2(n3235), .ZN(n3285) );
  INV_X1 U4037 ( .A(n3285), .ZN(n3241) );
  OAI22_X1 U4038 ( .A1(n4136), .A2(n3237), .B1(n3236), .B2(n4211), .ZN(n3240)
         );
  XOR2_X1 U4039 ( .A(n3813), .B(n3238), .Z(n3282) );
  NOR2_X1 U4040 ( .A1(n3282), .A2(n4217), .ZN(n3239) );
  AOI211_X1 U4041 ( .C1(n3241), .C2(n4446), .A(n3240), .B(n3239), .ZN(n3242)
         );
  OAI21_X1 U4042 ( .B1(n4458), .B2(n3281), .A(n3242), .ZN(U3280) );
  NAND2_X1 U40430 ( .A1(n3873), .A2(n2978), .ZN(n3247) );
  OR2_X1 U4044 ( .A1(n3297), .A2(n3538), .ZN(n3246) );
  NAND2_X1 U4045 ( .A1(n3247), .A2(n3246), .ZN(n3248) );
  XNOR2_X1 U4046 ( .A(n3248), .B(n3547), .ZN(n3251) );
  NAND2_X1 U4047 ( .A1(n2005), .A2(n3873), .ZN(n3250) );
  OR2_X1 U4048 ( .A1(n3297), .A2(n3546), .ZN(n3249) );
  NAND2_X1 U4049 ( .A1(n3250), .A2(n3249), .ZN(n3252) );
  INV_X1 U4050 ( .A(n3251), .ZN(n3254) );
  INV_X1 U4051 ( .A(n3252), .ZN(n3253) );
  NAND2_X1 U4052 ( .A1(n3254), .A2(n3253), .ZN(n3307) );
  NAND2_X1 U4053 ( .A1(n2054), .A2(n3307), .ZN(n3255) );
  XNOR2_X1 U4054 ( .A(n3308), .B(n3255), .ZN(n3260) );
  AND2_X1 U4055 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4379) );
  AOI21_X1 U4056 ( .B1(n3697), .B2(n3874), .A(n4379), .ZN(n3258) );
  AOI22_X1 U4057 ( .A1(n3256), .A2(n3640), .B1(n3696), .B2(n3872), .ZN(n3257)
         );
  OAI211_X1 U4058 ( .C1(n3702), .C2(n3300), .A(n3258), .B(n3257), .ZN(n3259)
         );
  AOI21_X1 U4059 ( .B1(n3260), .B2(n3704), .A(n3259), .ZN(n3261) );
  INV_X1 U4060 ( .A(n3261), .ZN(U3221) );
  XNOR2_X1 U4061 ( .A(n3292), .B(n3264), .ZN(n3270) );
  OAI21_X1 U4062 ( .B1(n2163), .B2(n3264), .A(n3263), .ZN(n3321) );
  NAND2_X1 U4063 ( .A1(n3875), .A2(n4155), .ZN(n3266) );
  NAND2_X1 U4064 ( .A1(n3873), .A2(n4200), .ZN(n3265) );
  OAI211_X1 U4065 ( .C1(n4198), .C2(n3273), .A(n3266), .B(n3265), .ZN(n3267)
         );
  AOI21_X1 U4066 ( .B1(n3321), .B2(n3268), .A(n3267), .ZN(n3269) );
  OAI21_X1 U4067 ( .B1(n4158), .B2(n3270), .A(n3269), .ZN(n3320) );
  INV_X1 U4068 ( .A(n3320), .ZN(n3280) );
  INV_X1 U4069 ( .A(n4144), .ZN(n4455) );
  INV_X1 U4070 ( .A(n3271), .ZN(n3274) );
  INV_X1 U4071 ( .A(n3298), .ZN(n3272) );
  OAI21_X1 U4072 ( .B1(n3274), .B2(n3273), .A(n3272), .ZN(n3326) );
  NOR2_X1 U4073 ( .A1(n3326), .A2(n4210), .ZN(n3278) );
  OAI22_X1 U4074 ( .A1(n4188), .A2(n3276), .B1(n3275), .B2(n4211), .ZN(n3277)
         );
  AOI211_X1 U4075 ( .C1(n3321), .C2(n4455), .A(n3278), .B(n3277), .ZN(n3279)
         );
  OAI21_X1 U4076 ( .B1(n3280), .B2(n4458), .A(n3279), .ZN(U3279) );
  OAI21_X1 U4077 ( .B1(n3282), .B2(n4501), .A(n3281), .ZN(n3287) );
  INV_X1 U4078 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4357) );
  OAI22_X1 U4079 ( .A1(n3285), .A2(n4275), .B1(n4524), .B2(n4357), .ZN(n3283)
         );
  AOI21_X1 U4080 ( .B1(n3287), .B2(n4524), .A(n3283), .ZN(n3284) );
  INV_X1 U4081 ( .A(n3284), .ZN(U3528) );
  OAI22_X1 U4082 ( .A1(n3285), .A2(n4320), .B1(n4516), .B2(n2452), .ZN(n3286)
         );
  AOI21_X1 U4083 ( .B1(n3287), .B2(n4516), .A(n3286), .ZN(n3288) );
  INV_X1 U4084 ( .A(n3288), .ZN(U3487) );
  INV_X1 U4085 ( .A(n3289), .ZN(n3290) );
  AOI21_X1 U4086 ( .B1(n3292), .B2(n3291), .A(n3290), .ZN(n3349) );
  NAND2_X1 U4087 ( .A1(n3348), .A2(n3346), .ZN(n3814) );
  XNOR2_X1 U4088 ( .A(n3349), .B(n3814), .ZN(n3296) );
  NAND2_X1 U4089 ( .A1(n3874), .A2(n4155), .ZN(n3294) );
  NAND2_X1 U4090 ( .A1(n3872), .A2(n4200), .ZN(n3293) );
  OAI211_X1 U4091 ( .C1(n4198), .C2(n3297), .A(n3294), .B(n3293), .ZN(n3295)
         );
  AOI21_X1 U4092 ( .B1(n3296), .B2(n4196), .A(n3295), .ZN(n3366) );
  OR2_X1 U4093 ( .A1(n3298), .A2(n3297), .ZN(n3299) );
  NAND2_X1 U4094 ( .A1(n3357), .A2(n3299), .ZN(n3373) );
  INV_X1 U4095 ( .A(n3373), .ZN(n3303) );
  OAI22_X1 U4096 ( .A1(n4188), .A2(n3301), .B1(n3300), .B2(n4211), .ZN(n3302)
         );
  AOI21_X1 U4097 ( .B1(n3303), .B2(n4446), .A(n3302), .ZN(n3306) );
  XNOR2_X1 U4098 ( .A(n3304), .B(n3814), .ZN(n3365) );
  NAND2_X1 U4099 ( .A1(n3365), .A2(n3412), .ZN(n3305) );
  OAI211_X1 U4100 ( .C1(n3366), .C2(n4458), .A(n3306), .B(n3305), .ZN(U3278)
         );
  NOR2_X1 U4101 ( .A1(n3546), .A2(n3358), .ZN(n3309) );
  AOI21_X1 U4102 ( .B1(n2005), .B2(n3872), .A(n3309), .ZN(n3381) );
  NAND2_X1 U4103 ( .A1(n3872), .A2(n2978), .ZN(n3311) );
  OR2_X1 U4104 ( .A1(n3358), .A2(n3538), .ZN(n3310) );
  NAND2_X1 U4105 ( .A1(n3311), .A2(n3310), .ZN(n3312) );
  XNOR2_X1 U4106 ( .A(n3312), .B(n3533), .ZN(n3383) );
  XOR2_X1 U4107 ( .A(n3381), .B(n3383), .Z(n3313) );
  XNOR2_X1 U4108 ( .A(n3384), .B(n3313), .ZN(n3318) );
  NOR2_X1 U4109 ( .A1(STATE_REG_SCAN_IN), .A2(n3314), .ZN(n4387) );
  AOI21_X1 U4110 ( .B1(n3696), .B2(n3871), .A(n4387), .ZN(n3316) );
  AOI22_X1 U4111 ( .A1(n3351), .A2(n3640), .B1(n3697), .B2(n3873), .ZN(n3315)
         );
  OAI211_X1 U4112 ( .C1(n3702), .C2(n3359), .A(n3316), .B(n3315), .ZN(n3317)
         );
  AOI21_X1 U4113 ( .B1(n3318), .B2(n3704), .A(n3317), .ZN(n3319) );
  INV_X1 U4114 ( .A(n3319), .ZN(U3231) );
  INV_X1 U4115 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3322) );
  AOI21_X1 U4116 ( .B1(n4495), .B2(n3321), .A(n3320), .ZN(n3324) );
  MUX2_X1 U4117 ( .A(n3322), .B(n3324), .S(n4516), .Z(n3323) );
  OAI21_X1 U4118 ( .B1(n3326), .B2(n4320), .A(n3323), .ZN(U3489) );
  MUX2_X1 U4119 ( .A(n2463), .B(n3324), .S(n4524), .Z(n3325) );
  OAI21_X1 U4120 ( .B1(n3326), .B2(n4275), .A(n3325), .ZN(U3529) );
  OAI21_X1 U4121 ( .B1(n3329), .B2(n3328), .A(n3327), .ZN(n3375) );
  INV_X1 U4122 ( .A(n3375), .ZN(n3341) );
  XNOR2_X1 U4123 ( .A(n3717), .B(n3832), .ZN(n3330) );
  NAND2_X1 U4124 ( .A1(n3330), .A2(n4196), .ZN(n3333) );
  NOR2_X1 U4125 ( .A1(n4198), .A2(n3390), .ZN(n3331) );
  AOI21_X1 U4126 ( .B1(n3870), .B2(n4200), .A(n3331), .ZN(n3332) );
  OAI211_X1 U4127 ( .C1(n3334), .C2(n4204), .A(n3333), .B(n3332), .ZN(n3374)
         );
  INV_X1 U4128 ( .A(n3413), .ZN(n3336) );
  NAND2_X1 U4129 ( .A1(n2015), .A2(n3399), .ZN(n3335) );
  NAND2_X1 U4130 ( .A1(n3336), .A2(n3335), .ZN(n3380) );
  NOR2_X1 U4131 ( .A1(n3380), .A2(n4210), .ZN(n3339) );
  OAI22_X1 U4132 ( .A1(n4188), .A2(n3337), .B1(n3402), .B2(n4211), .ZN(n3338)
         );
  AOI211_X1 U4133 ( .C1(n3374), .C2(n4136), .A(n3339), .B(n3338), .ZN(n3340)
         );
  OAI21_X1 U4134 ( .B1(n3341), .B2(n4217), .A(n3340), .ZN(U3276) );
  INV_X1 U4135 ( .A(n3342), .ZN(n3344) );
  OR2_X1 U4136 ( .A1(n3344), .A2(n3343), .ZN(n3818) );
  XOR2_X1 U4137 ( .A(n3818), .B(n3345), .Z(n3433) );
  INV_X1 U4138 ( .A(n3346), .ZN(n3347) );
  AOI21_X1 U4139 ( .B1(n3349), .B2(n3348), .A(n3347), .ZN(n3350) );
  XOR2_X1 U4140 ( .A(n3818), .B(n3350), .Z(n3355) );
  AOI22_X1 U4141 ( .A1(n3871), .A2(n4200), .B1(n4227), .B2(n3351), .ZN(n3352)
         );
  OAI21_X1 U4142 ( .B1(n3353), .B2(n4204), .A(n3352), .ZN(n3354) );
  AOI21_X1 U4143 ( .B1(n3355), .B2(n4196), .A(n3354), .ZN(n3356) );
  OAI21_X1 U4144 ( .B1(n3433), .B2(n4135), .A(n3356), .ZN(n3434) );
  NAND2_X1 U4145 ( .A1(n3434), .A2(n4136), .ZN(n3364) );
  OAI21_X1 U4146 ( .B1(n2101), .B2(n3358), .A(n2015), .ZN(n3440) );
  INV_X1 U4147 ( .A(n3440), .ZN(n3362) );
  OAI22_X1 U4148 ( .A1(n4188), .A2(n3360), .B1(n3359), .B2(n4211), .ZN(n3361)
         );
  AOI21_X1 U4149 ( .B1(n3362), .B2(n4446), .A(n3361), .ZN(n3363) );
  OAI211_X1 U4150 ( .C1(n3433), .C2(n4144), .A(n3364), .B(n3363), .ZN(U3277)
         );
  NAND2_X1 U4151 ( .A1(n3365), .A2(n4512), .ZN(n3367) );
  NAND2_X1 U4152 ( .A1(n3367), .A2(n3366), .ZN(n3370) );
  MUX2_X1 U4153 ( .A(REG1_REG_12__SCAN_IN), .B(n3370), .S(n4524), .Z(n3368) );
  INV_X1 U4154 ( .A(n3368), .ZN(n3369) );
  OAI21_X1 U4155 ( .B1(n4275), .B2(n3373), .A(n3369), .ZN(U3530) );
  MUX2_X1 U4156 ( .A(REG0_REG_12__SCAN_IN), .B(n3370), .S(n4516), .Z(n3371) );
  INV_X1 U4157 ( .A(n3371), .ZN(n3372) );
  OAI21_X1 U4158 ( .B1(n3373), .B2(n4320), .A(n3372), .ZN(U3491) );
  AOI21_X1 U4159 ( .B1(n3375), .B2(n4512), .A(n3374), .ZN(n3377) );
  MUX2_X1 U4160 ( .A(n4397), .B(n3377), .S(n4524), .Z(n3376) );
  OAI21_X1 U4161 ( .B1(n4275), .B2(n3380), .A(n3376), .ZN(U3532) );
  INV_X1 U4162 ( .A(REG0_REG_14__SCAN_IN), .ZN(n3378) );
  MUX2_X1 U4163 ( .A(n3378), .B(n3377), .S(n4516), .Z(n3379) );
  OAI21_X1 U4164 ( .B1(n3380), .B2(n4320), .A(n3379), .ZN(U3495) );
  AOI21_X1 U4165 ( .B1(n3384), .B2(n3383), .A(n3381), .ZN(n3382) );
  INV_X1 U4166 ( .A(n3382), .ZN(n3386) );
  NAND2_X2 U4167 ( .A1(n3386), .A2(n3385), .ZN(n3447) );
  NAND2_X1 U4168 ( .A1(n3871), .A2(n2978), .ZN(n3388) );
  OR2_X1 U4169 ( .A1(n3390), .A2(n3538), .ZN(n3387) );
  NAND2_X1 U4170 ( .A1(n3388), .A2(n3387), .ZN(n3389) );
  XNOR2_X1 U4171 ( .A(n3389), .B(n3547), .ZN(n3393) );
  NAND2_X1 U4172 ( .A1(n2005), .A2(n3871), .ZN(n3392) );
  OR2_X1 U4173 ( .A1(n3390), .A2(n3546), .ZN(n3391) );
  NAND2_X1 U4174 ( .A1(n3392), .A2(n3391), .ZN(n3394) );
  AND2_X1 U4175 ( .A1(n3393), .A2(n3394), .ZN(n3446) );
  INV_X1 U4176 ( .A(n3393), .ZN(n3396) );
  INV_X1 U4177 ( .A(n3394), .ZN(n3395) );
  NAND2_X1 U4178 ( .A1(n3396), .A2(n3395), .ZN(n3445) );
  NAND2_X1 U4179 ( .A1(n2247), .A2(n3445), .ZN(n3397) );
  XNOR2_X1 U4180 ( .A(n3447), .B(n3397), .ZN(n3404) );
  NAND2_X1 U4181 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4404) );
  INV_X1 U4182 ( .A(n4404), .ZN(n3398) );
  AOI21_X1 U4183 ( .B1(n3697), .B2(n3872), .A(n3398), .ZN(n3401) );
  AOI22_X1 U4184 ( .A1(n3399), .A2(n3640), .B1(n3696), .B2(n3870), .ZN(n3400)
         );
  OAI211_X1 U4185 ( .C1(n3702), .C2(n3402), .A(n3401), .B(n3400), .ZN(n3403)
         );
  AOI21_X1 U4186 ( .B1(n3404), .B2(n3704), .A(n3403), .ZN(n3405) );
  INV_X1 U4187 ( .A(n3405), .ZN(U3212) );
  OAI22_X1 U4188 ( .A1(n4205), .A2(n4090), .B1(n4198), .B2(n3459), .ZN(n3410)
         );
  INV_X1 U4189 ( .A(n3406), .ZN(n3407) );
  AOI211_X1 U4190 ( .C1(n3408), .C2(n3822), .A(n4158), .B(n3407), .ZN(n3409)
         );
  AOI211_X1 U4191 ( .C1(n4155), .C2(n3871), .A(n3410), .B(n3409), .ZN(n4281)
         );
  XNOR2_X1 U4192 ( .A(n3411), .B(n3822), .ZN(n4280) );
  NAND2_X1 U4193 ( .A1(n4280), .A2(n3412), .ZN(n3418) );
  XNOR2_X1 U4194 ( .A(n3413), .B(n3459), .ZN(n4283) );
  INV_X1 U4195 ( .A(n4283), .ZN(n3416) );
  OAI22_X1 U4196 ( .A1(n4188), .A2(n3414), .B1(n3701), .B2(n4211), .ZN(n3415)
         );
  AOI21_X1 U4197 ( .B1(n3416), .B2(n4446), .A(n3415), .ZN(n3417) );
  OAI211_X1 U4198 ( .C1(n4458), .C2(n4281), .A(n3418), .B(n3417), .ZN(U3275)
         );
  OAI21_X1 U4199 ( .B1(n3421), .B2(n3420), .A(n3419), .ZN(n4279) );
  INV_X1 U4200 ( .A(n3422), .ZN(n4209) );
  AOI21_X1 U4201 ( .B1(n3617), .B2(n3423), .A(n4209), .ZN(n4277) );
  OAI22_X1 U4202 ( .A1(n4188), .A2(n3424), .B1(n3620), .B2(n4211), .ZN(n3425)
         );
  AOI21_X1 U4203 ( .B1(n4277), .B2(n4446), .A(n3425), .ZN(n3432) );
  OAI211_X1 U4204 ( .C1(n3828), .C2(n3426), .A(n4193), .B(n4196), .ZN(n3429)
         );
  NOR2_X1 U4205 ( .A1(n4198), .A2(n3454), .ZN(n3427) );
  AOI21_X1 U4206 ( .B1(n3868), .B2(n4200), .A(n3427), .ZN(n3428) );
  OAI211_X1 U4207 ( .C1(n3430), .C2(n4204), .A(n3429), .B(n3428), .ZN(n4276)
         );
  NAND2_X1 U4208 ( .A1(n4276), .A2(n4136), .ZN(n3431) );
  OAI211_X1 U4209 ( .C1(n4279), .C2(n4217), .A(n3432), .B(n3431), .ZN(U3274)
         );
  INV_X1 U4210 ( .A(n3433), .ZN(n3435) );
  AOI21_X1 U4211 ( .B1(n4495), .B2(n3435), .A(n3434), .ZN(n3437) );
  MUX2_X1 U4212 ( .A(n4535), .B(n3437), .S(n4524), .Z(n3436) );
  OAI21_X1 U4213 ( .B1(n4275), .B2(n3440), .A(n3436), .ZN(U3531) );
  INV_X1 U4214 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3438) );
  MUX2_X1 U4215 ( .A(n3438), .B(n3437), .S(n4516), .Z(n3439) );
  OAI21_X1 U4216 ( .B1(n3440), .B2(n4320), .A(n3439), .ZN(U3493) );
  AOI22_X1 U4217 ( .A1(n3697), .A2(n3867), .B1(n3640), .B2(n3441), .ZN(n3443)
         );
  NAND2_X1 U4218 ( .A1(n4054), .A2(n3696), .ZN(n3442) );
  OAI211_X1 U4219 ( .C1(STATE_REG_SCAN_IN), .C2(n3444), .A(n3443), .B(n3442), 
        .ZN(n3515) );
  NAND2_X1 U4220 ( .A1(n3870), .A2(n2978), .ZN(n3449) );
  OR2_X1 U4221 ( .A1(n3459), .A2(n3538), .ZN(n3448) );
  NAND2_X1 U4222 ( .A1(n3449), .A2(n3448), .ZN(n3450) );
  XNOR2_X1 U4223 ( .A(n3450), .B(n3533), .ZN(n3458) );
  NAND2_X1 U4224 ( .A1(n3869), .A2(n2978), .ZN(n3452) );
  OR2_X1 U4225 ( .A1(n3454), .A2(n3538), .ZN(n3451) );
  NAND2_X1 U4226 ( .A1(n3452), .A2(n3451), .ZN(n3453) );
  XNOR2_X1 U4227 ( .A(n3453), .B(n3533), .ZN(n3457) );
  NOR2_X1 U4228 ( .A1(n3546), .A2(n3454), .ZN(n3455) );
  AOI21_X1 U4229 ( .B1(n2005), .B2(n3869), .A(n3455), .ZN(n3456) );
  NAND2_X1 U4230 ( .A1(n3457), .A2(n3456), .ZN(n3462) );
  OAI21_X1 U4231 ( .B1(n3457), .B2(n3456), .A(n3462), .ZN(n3615) );
  NAND2_X1 U4232 ( .A1(n2005), .A2(n3870), .ZN(n3461) );
  OR2_X1 U4233 ( .A1(n3459), .A2(n3546), .ZN(n3460) );
  NAND2_X1 U4234 ( .A1(n3461), .A2(n3460), .ZN(n3693) );
  NAND2_X1 U4235 ( .A1(n3868), .A2(n2978), .ZN(n3464) );
  OR2_X1 U4236 ( .A1(n4208), .A2(n3538), .ZN(n3463) );
  NAND2_X1 U4237 ( .A1(n3464), .A2(n3463), .ZN(n3465) );
  XNOR2_X1 U4238 ( .A(n3465), .B(n3533), .ZN(n3468) );
  NOR2_X1 U4239 ( .A1(n3546), .A2(n4208), .ZN(n3466) );
  AOI21_X1 U4240 ( .B1(n2005), .B2(n3868), .A(n3466), .ZN(n3467) );
  NOR2_X1 U4241 ( .A1(n3468), .A2(n3467), .ZN(n3634) );
  NAND2_X1 U4242 ( .A1(n3468), .A2(n3467), .ZN(n3635) );
  INV_X1 U4243 ( .A(n3671), .ZN(n3472) );
  AOI22_X1 U4244 ( .A1(n2005), .A2(n4201), .B1(n2978), .B2(n4181), .ZN(n3470)
         );
  INV_X1 U4245 ( .A(n3470), .ZN(n3668) );
  AOI22_X1 U4246 ( .A1(n4201), .A2(n2978), .B1(n3495), .B2(n4181), .ZN(n3469)
         );
  XNOR2_X1 U4247 ( .A(n3469), .B(n3547), .ZN(n3669) );
  AOI21_X1 U4248 ( .B1(n3671), .B2(n3470), .A(n3669), .ZN(n3471) );
  AOI21_X1 U4249 ( .B1(n3472), .B2(n3668), .A(n3471), .ZN(n3584) );
  NAND2_X1 U4250 ( .A1(n4176), .A2(n2978), .ZN(n3474) );
  OR2_X1 U4251 ( .A1(n4160), .A2(n3538), .ZN(n3473) );
  NAND2_X1 U4252 ( .A1(n3474), .A2(n3473), .ZN(n3475) );
  XNOR2_X1 U4253 ( .A(n3475), .B(n3533), .ZN(n3478) );
  INV_X1 U4254 ( .A(n3478), .ZN(n3480) );
  NOR2_X1 U4255 ( .A1(n3546), .A2(n4160), .ZN(n3476) );
  AOI21_X1 U4256 ( .B1(n2005), .B2(n4176), .A(n3476), .ZN(n3477) );
  INV_X1 U4257 ( .A(n3477), .ZN(n3479) );
  AND2_X1 U4258 ( .A1(n3478), .A2(n3477), .ZN(n3481) );
  AOI21_X1 U4259 ( .B1(n3480), .B2(n3479), .A(n3481), .ZN(n3585) );
  NAND2_X1 U4260 ( .A1(n3584), .A2(n3585), .ZN(n3583) );
  INV_X1 U4261 ( .A(n3481), .ZN(n3482) );
  NAND2_X1 U4262 ( .A1(n4154), .A2(n2978), .ZN(n3484) );
  OR2_X1 U4263 ( .A1(n3538), .A2(n4137), .ZN(n3483) );
  NAND2_X1 U4264 ( .A1(n3484), .A2(n3483), .ZN(n3485) );
  XNOR2_X1 U4265 ( .A(n3485), .B(n3533), .ZN(n3488) );
  NOR2_X1 U4266 ( .A1(n3546), .A2(n4137), .ZN(n3486) );
  AOI21_X1 U4267 ( .B1(n4154), .B2(n2005), .A(n3486), .ZN(n3487) );
  OR2_X1 U4268 ( .A1(n3488), .A2(n3487), .ZN(n3647) );
  NAND2_X1 U4269 ( .A1(n3488), .A2(n3487), .ZN(n3596) );
  NAND2_X1 U4270 ( .A1(n4129), .A2(n2978), .ZN(n3490) );
  OR2_X1 U4271 ( .A1(n3538), .A2(n4107), .ZN(n3489) );
  NAND2_X1 U4272 ( .A1(n3490), .A2(n3489), .ZN(n3491) );
  XNOR2_X1 U4273 ( .A(n3491), .B(n3533), .ZN(n3494) );
  NOR2_X1 U4274 ( .A1(n3546), .A2(n4107), .ZN(n3492) );
  AOI21_X1 U4275 ( .B1(n4129), .B2(n2005), .A(n3492), .ZN(n3493) );
  AND2_X1 U4276 ( .A1(n3494), .A2(n3493), .ZN(n3593) );
  OR2_X1 U4277 ( .A1(n3494), .A2(n3493), .ZN(n3594) );
  AOI22_X1 U4278 ( .A1(n4110), .A2(n2978), .B1(n3495), .B2(n4097), .ZN(n3496)
         );
  XNOR2_X1 U4279 ( .A(n3496), .B(n3547), .ZN(n3497) );
  AOI22_X1 U4280 ( .A1(n4110), .A2(n2005), .B1(n2978), .B2(n4097), .ZN(n3498)
         );
  XNOR2_X1 U4281 ( .A(n3497), .B(n3498), .ZN(n3660) );
  INV_X1 U4282 ( .A(n3497), .ZN(n3500) );
  INV_X1 U4283 ( .A(n3498), .ZN(n3499) );
  NOR2_X1 U4284 ( .A1(n3500), .A2(n3499), .ZN(n3575) );
  NOR2_X1 U4285 ( .A1(n3546), .A2(n4078), .ZN(n3501) );
  AOI21_X1 U4286 ( .B1(n3867), .B2(n2005), .A(n3501), .ZN(n3504) );
  OAI22_X1 U4287 ( .A1(n4091), .A2(n3546), .B1(n3538), .B2(n4078), .ZN(n3502)
         );
  XNOR2_X1 U4288 ( .A(n3502), .B(n3547), .ZN(n3503) );
  XOR2_X1 U4289 ( .A(n3504), .B(n3503), .Z(n3574) );
  INV_X1 U4290 ( .A(n3503), .ZN(n3505) );
  NOR2_X1 U4291 ( .A1(n3505), .A2(n3504), .ZN(n3509) );
  NAND2_X1 U4292 ( .A1(n4073), .A2(n2005), .ZN(n3507) );
  OR2_X1 U4293 ( .A1(n3546), .A2(n4058), .ZN(n3506) );
  NAND2_X1 U4294 ( .A1(n3507), .A2(n3506), .ZN(n3510) );
  OAI21_X1 U4295 ( .B1(n3508), .B2(n3509), .A(n3510), .ZN(n3522) );
  INV_X1 U4296 ( .A(n3508), .ZN(n3577) );
  OAI22_X1 U4297 ( .A1(n4034), .A2(n3550), .B1(n3538), .B2(n4058), .ZN(n3512)
         );
  XOR2_X1 U4298 ( .A(n3547), .B(n3512), .Z(n3523) );
  XNOR2_X1 U4299 ( .A(n3513), .B(n3523), .ZN(n3514) );
  INV_X1 U4300 ( .A(D_REG_0__SCAN_IN), .ZN(n3518) );
  NOR3_X1 U4301 ( .A1(n3516), .A2(n2665), .A3(n4327), .ZN(n3517) );
  AOI21_X1 U4302 ( .B1(n4460), .B2(n3518), .A(n3517), .ZN(U3458) );
  NAND3_X1 U4303 ( .A1(n3519), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3521) );
  INV_X1 U4304 ( .A(DATAI_31_), .ZN(n3520) );
  OAI22_X1 U4305 ( .A1(n2288), .A2(n3521), .B1(STATE_REG_SCAN_IN), .B2(n3520), 
        .ZN(U3321) );
  NAND2_X1 U4306 ( .A1(n4054), .A2(n2978), .ZN(n3526) );
  OR2_X1 U4307 ( .A1(n3538), .A2(n4040), .ZN(n3525) );
  NAND2_X1 U4308 ( .A1(n3526), .A2(n3525), .ZN(n3527) );
  XNOR2_X1 U4309 ( .A(n3527), .B(n3533), .ZN(n3530) );
  NOR2_X1 U4310 ( .A1(n3550), .A2(n4040), .ZN(n3528) );
  AOI21_X1 U4311 ( .B1(n4054), .B2(n2005), .A(n3528), .ZN(n3529) );
  NAND2_X1 U4312 ( .A1(n3530), .A2(n3529), .ZN(n3606) );
  NOR2_X1 U4313 ( .A1(n3530), .A2(n3529), .ZN(n3607) );
  NAND2_X1 U4314 ( .A1(n4036), .A2(n2978), .ZN(n3532) );
  OR2_X1 U4315 ( .A1(n3538), .A2(n4022), .ZN(n3531) );
  NAND2_X1 U4316 ( .A1(n3532), .A2(n3531), .ZN(n3534) );
  XNOR2_X1 U4317 ( .A(n3534), .B(n3533), .ZN(n3537) );
  NOR2_X1 U4318 ( .A1(n3546), .A2(n4022), .ZN(n3535) );
  AOI21_X1 U4319 ( .B1(n4036), .B2(n2005), .A(n3535), .ZN(n3536) );
  OR2_X1 U4320 ( .A1(n3537), .A2(n3536), .ZN(n3677) );
  NAND2_X1 U4321 ( .A1(n4019), .A2(n2978), .ZN(n3540) );
  OR2_X1 U4322 ( .A1(n3538), .A2(n3998), .ZN(n3539) );
  NAND2_X1 U4323 ( .A1(n3540), .A2(n3539), .ZN(n3541) );
  XNOR2_X1 U4324 ( .A(n3541), .B(n3547), .ZN(n3543) );
  NOR2_X1 U4325 ( .A1(n3550), .A2(n3998), .ZN(n3542) );
  AOI21_X1 U4326 ( .B1(n4019), .B2(n2005), .A(n3542), .ZN(n3544) );
  XNOR2_X1 U4327 ( .A(n3543), .B(n3544), .ZN(n3568) );
  INV_X1 U4328 ( .A(n3543), .ZN(n3545) );
  OAI22_X1 U4329 ( .A1(n3982), .A2(n3546), .B1(n3538), .B2(n3549), .ZN(n3548)
         );
  XNOR2_X1 U4330 ( .A(n3548), .B(n3547), .ZN(n3552) );
  OAI22_X1 U4331 ( .A1(n3982), .A2(n2004), .B1(n3550), .B2(n3549), .ZN(n3551)
         );
  AOI22_X1 U4332 ( .A1(n3866), .A2(n3696), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3554) );
  AOI22_X1 U4333 ( .A1(n4019), .A2(n3697), .B1(n3970), .B2(n3640), .ZN(n3553)
         );
  OAI211_X1 U4334 ( .C1(n3702), .C2(n3560), .A(n3554), .B(n3553), .ZN(n3555)
         );
  INV_X1 U4335 ( .A(n3555), .ZN(n3556) );
  OAI21_X1 U4336 ( .B1(n3557), .B2(n3688), .A(n3556), .ZN(U3217) );
  INV_X1 U4337 ( .A(n3558), .ZN(n3564) );
  INV_X1 U4338 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3559) );
  OAI22_X1 U4339 ( .A1(n3560), .A2(n4211), .B1(n3559), .B2(n4136), .ZN(n3563)
         );
  NOR2_X1 U4340 ( .A1(n3561), .A2(n4458), .ZN(n3562) );
  AOI211_X1 U4341 ( .C1(n4446), .C2(n3564), .A(n3563), .B(n3562), .ZN(n3565)
         );
  OAI21_X1 U4342 ( .B1(n3566), .B2(n4217), .A(n3565), .ZN(U3262) );
  XNOR2_X1 U4343 ( .A(n3567), .B(n3568), .ZN(n3573) );
  OAI22_X1 U4344 ( .A1(n3999), .A2(n3681), .B1(STATE_REG_SCAN_IN), .B2(n3569), 
        .ZN(n3571) );
  OAI22_X1 U4345 ( .A1(n3982), .A2(n3683), .B1(n3680), .B2(n3998), .ZN(n3570)
         );
  AOI211_X1 U4346 ( .C1(n4006), .C2(n3686), .A(n3571), .B(n3570), .ZN(n3572)
         );
  OAI21_X1 U4347 ( .B1(n3573), .B2(n3688), .A(n3572), .ZN(U3211) );
  OAI21_X1 U4348 ( .B1(n3658), .B2(n3575), .A(n3574), .ZN(n3576) );
  NAND3_X1 U4349 ( .A1(n3577), .A2(n3704), .A3(n3576), .ZN(n3582) );
  AOI22_X1 U4350 ( .A1(n4073), .A2(n3696), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3581) );
  AOI22_X1 U4351 ( .A1(n3578), .A2(n3640), .B1(n3697), .B2(n4110), .ZN(n3580)
         );
  OR2_X1 U4352 ( .A1(n3702), .A2(n4080), .ZN(n3579) );
  NAND4_X1 U4353 ( .A1(n3582), .A2(n3581), .A3(n3580), .A4(n3579), .ZN(U3213)
         );
  OAI21_X1 U4354 ( .B1(n3585), .B2(n3584), .A(n3583), .ZN(n3591) );
  NAND2_X1 U4355 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3965) );
  INV_X1 U4356 ( .A(n3965), .ZN(n3586) );
  AOI21_X1 U4357 ( .B1(n3696), .B2(n4154), .A(n3586), .ZN(n3589) );
  AOI22_X1 U4358 ( .A1(n3587), .A2(n3640), .B1(n3697), .B2(n4201), .ZN(n3588)
         );
  OAI211_X1 U4359 ( .C1(n3702), .C2(n4164), .A(n3589), .B(n3588), .ZN(n3590)
         );
  AOI21_X1 U4360 ( .B1(n3591), .B2(n3704), .A(n3590), .ZN(n3592) );
  INV_X1 U4361 ( .A(n3592), .ZN(U3216) );
  INV_X1 U4362 ( .A(n3593), .ZN(n3595) );
  NAND2_X1 U4363 ( .A1(n3595), .A2(n3594), .ZN(n3598) );
  OAI211_X1 U4364 ( .C1(n3648), .C2(n2202), .A(n3647), .B(n3598), .ZN(n3597)
         );
  OAI211_X1 U4365 ( .C1(n3599), .C2(n3598), .A(n3704), .B(n3597), .ZN(n3604)
         );
  OAI22_X1 U4366 ( .A1(n3680), .A2(n4107), .B1(n3681), .B2(n4108), .ZN(n3602)
         );
  OAI22_X1 U4367 ( .A1(n3683), .A2(n4071), .B1(STATE_REG_SCAN_IN), .B2(n3600), 
        .ZN(n3601) );
  NOR2_X1 U4368 ( .A1(n3602), .A2(n3601), .ZN(n3603) );
  OAI211_X1 U4369 ( .C1(n3702), .C2(n4115), .A(n3604), .B(n3603), .ZN(U3220)
         );
  NOR2_X1 U4370 ( .A1(n3607), .A2(n2225), .ZN(n3608) );
  XNOR2_X1 U4371 ( .A(n3605), .B(n3608), .ZN(n3613) );
  INV_X1 U4372 ( .A(n3609), .ZN(n4042) );
  OAI22_X1 U4373 ( .A1(n4034), .A2(n3681), .B1(n3680), .B2(n4040), .ZN(n3611)
         );
  OAI22_X1 U4374 ( .A1(n3999), .A2(n3683), .B1(STATE_REG_SCAN_IN), .B2(n4602), 
        .ZN(n3610) );
  AOI211_X1 U4375 ( .C1(n4042), .C2(n3686), .A(n3611), .B(n3610), .ZN(n3612)
         );
  OAI21_X1 U4376 ( .B1(n3613), .B2(n3688), .A(n3612), .ZN(U3222) );
  OAI21_X1 U4377 ( .B1(n3690), .B2(n3693), .A(n3691), .ZN(n3614) );
  XOR2_X1 U4378 ( .A(n3615), .B(n3614), .Z(n3622) );
  NAND2_X1 U4379 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n3943) );
  INV_X1 U4380 ( .A(n3943), .ZN(n3616) );
  AOI21_X1 U4381 ( .B1(n3696), .B2(n3868), .A(n3616), .ZN(n3619) );
  AOI22_X1 U4382 ( .A1(n3617), .A2(n3640), .B1(n3697), .B2(n3870), .ZN(n3618)
         );
  OAI211_X1 U4383 ( .C1(n3702), .C2(n3620), .A(n3619), .B(n3618), .ZN(n3621)
         );
  AOI21_X1 U4384 ( .B1(n3622), .B2(n3704), .A(n3621), .ZN(n3623) );
  INV_X1 U4385 ( .A(n3623), .ZN(U3223) );
  OAI211_X1 U4386 ( .C1(n3626), .C2(n3625), .A(n3624), .B(n3704), .ZN(n3633)
         );
  AOI21_X1 U4387 ( .B1(n3697), .B2(n3880), .A(n3627), .ZN(n3632) );
  AOI22_X1 U4388 ( .A1(n3628), .A2(n3640), .B1(n3696), .B2(n3879), .ZN(n3631)
         );
  OR2_X1 U4389 ( .A1(n3702), .A2(n3629), .ZN(n3630) );
  NAND4_X1 U4390 ( .A1(n3633), .A2(n3632), .A3(n3631), .A4(n3630), .ZN(U3224)
         );
  INV_X1 U4391 ( .A(n3634), .ZN(n3636) );
  NAND2_X1 U4392 ( .A1(n3636), .A2(n3635), .ZN(n3637) );
  XNOR2_X1 U4393 ( .A(n3638), .B(n3637), .ZN(n3645) );
  NOR2_X1 U4394 ( .A1(STATE_REG_SCAN_IN), .A2(n3639), .ZN(n4418) );
  AOI21_X1 U4395 ( .B1(n3696), .B2(n4201), .A(n4418), .ZN(n3643) );
  AOI22_X1 U4396 ( .A1(n3641), .A2(n3640), .B1(n3697), .B2(n3869), .ZN(n3642)
         );
  OAI211_X1 U4397 ( .C1(n3702), .C2(n4212), .A(n3643), .B(n3642), .ZN(n3644)
         );
  AOI21_X1 U4398 ( .B1(n3645), .B2(n3704), .A(n3644), .ZN(n3646) );
  INV_X1 U4399 ( .A(n3646), .ZN(U3225) );
  NOR2_X1 U4400 ( .A1(n2202), .A2(n2199), .ZN(n3649) );
  OAI22_X1 U4401 ( .A1(n3650), .A2(n2202), .B1(n3649), .B2(n3648), .ZN(n3656)
         );
  NOR2_X1 U4402 ( .A1(n3651), .A2(STATE_REG_SCAN_IN), .ZN(n3652) );
  AOI21_X1 U4403 ( .B1(n3696), .B2(n4129), .A(n3652), .ZN(n3654) );
  AOI22_X1 U4404 ( .A1(n4128), .A2(n3640), .B1(n3697), .B2(n4176), .ZN(n3653)
         );
  OAI211_X1 U4405 ( .C1(n3702), .C2(n4138), .A(n3654), .B(n3653), .ZN(n3655)
         );
  AOI21_X1 U4406 ( .B1(n3656), .B2(n3704), .A(n3655), .ZN(n3657) );
  INV_X1 U4407 ( .A(n3657), .ZN(U3230) );
  AOI21_X1 U4408 ( .B1(n3660), .B2(n3659), .A(n3658), .ZN(n3667) );
  INV_X1 U4409 ( .A(n4098), .ZN(n3665) );
  OAI22_X1 U4410 ( .A1(n3683), .A2(n4091), .B1(STATE_REG_SCAN_IN), .B2(n3661), 
        .ZN(n3664) );
  OAI22_X1 U4411 ( .A1(n3680), .A2(n3662), .B1(n3681), .B2(n2186), .ZN(n3663)
         );
  AOI211_X1 U4412 ( .C1(n3665), .C2(n3686), .A(n3664), .B(n3663), .ZN(n3666)
         );
  OAI21_X1 U4413 ( .B1(n3667), .B2(n3688), .A(n3666), .ZN(U3232) );
  XNOR2_X1 U4414 ( .A(n3669), .B(n3668), .ZN(n3670) );
  XNOR2_X1 U4415 ( .A(n3671), .B(n3670), .ZN(n3675) );
  AND2_X1 U4416 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4433) );
  AOI21_X1 U4417 ( .B1(n3696), .B2(n4176), .A(n4433), .ZN(n3673) );
  AOI22_X1 U4418 ( .A1(n4181), .A2(n3640), .B1(n3697), .B2(n3868), .ZN(n3672)
         );
  OAI211_X1 U4419 ( .C1(n3702), .C2(n4184), .A(n3673), .B(n3672), .ZN(n3674)
         );
  AOI21_X1 U4420 ( .B1(n3675), .B2(n3704), .A(n3674), .ZN(n3676) );
  INV_X1 U4421 ( .A(n3676), .ZN(U3235) );
  NAND2_X1 U4422 ( .A1(n3677), .A2(n2223), .ZN(n3678) );
  XNOR2_X1 U4423 ( .A(n3679), .B(n3678), .ZN(n3689) );
  OAI22_X1 U4424 ( .A1(n4017), .A2(n3681), .B1(n3680), .B2(n4022), .ZN(n3685)
         );
  OAI22_X1 U4425 ( .A1(n3744), .A2(n3683), .B1(STATE_REG_SCAN_IN), .B2(n3682), 
        .ZN(n3684) );
  AOI211_X1 U4426 ( .C1(n4024), .C2(n3686), .A(n3685), .B(n3684), .ZN(n3687)
         );
  OAI21_X1 U4427 ( .B1(n3689), .B2(n3688), .A(n3687), .ZN(U3237) );
  INV_X1 U4428 ( .A(n3690), .ZN(n3692) );
  NAND2_X1 U4429 ( .A1(n3692), .A2(n3691), .ZN(n3694) );
  XNOR2_X1 U4430 ( .A(n3694), .B(n3693), .ZN(n3705) );
  NOR2_X1 U4431 ( .A1(STATE_REG_SCAN_IN), .A2(n3695), .ZN(n4411) );
  AOI21_X1 U4432 ( .B1(n3696), .B2(n3869), .A(n4411), .ZN(n3700) );
  AOI22_X1 U4433 ( .A1(n3698), .A2(n3640), .B1(n3697), .B2(n3871), .ZN(n3699)
         );
  OAI211_X1 U4434 ( .C1(n3702), .C2(n3701), .A(n3700), .B(n3699), .ZN(n3703)
         );
  AOI21_X1 U4435 ( .B1(n3705), .B2(n3704), .A(n3703), .ZN(n3706) );
  INV_X1 U4436 ( .A(n3706), .ZN(U3238) );
  NAND2_X1 U4437 ( .A1(n2379), .A2(DATAI_30_), .ZN(n4219) );
  INV_X1 U4438 ( .A(REG2_REG_31__SCAN_IN), .ZN(n3710) );
  NAND2_X1 U4439 ( .A1(n2352), .A2(REG0_REG_31__SCAN_IN), .ZN(n3709) );
  INV_X1 U4440 ( .A(REG1_REG_31__SCAN_IN), .ZN(n3707) );
  OAI211_X1 U4441 ( .C1(n2371), .C2(n3710), .A(n3709), .B(n3708), .ZN(n4221)
         );
  NAND2_X1 U4442 ( .A1(n3711), .A2(n3715), .ZN(n3776) );
  INV_X1 U4443 ( .A(n3712), .ZN(n3716) );
  INV_X1 U4444 ( .A(n3713), .ZN(n3714) );
  AOI21_X1 U4445 ( .B1(n3716), .B2(n3715), .A(n3714), .ZN(n3781) );
  OAI21_X1 U4446 ( .B1(n3717), .B2(n3776), .A(n3781), .ZN(n3720) );
  INV_X1 U4447 ( .A(n3718), .ZN(n3719) );
  AOI21_X1 U4448 ( .B1(n3720), .B2(n3784), .A(n3719), .ZN(n3721) );
  OAI21_X1 U4449 ( .B1(n3721), .B2(n3787), .A(n3786), .ZN(n3723) );
  AOI21_X1 U4450 ( .B1(n3790), .B2(n3723), .A(n3722), .ZN(n3725) );
  OAI21_X1 U4451 ( .B1(n3725), .B2(n3792), .A(n3724), .ZN(n3726) );
  NAND4_X1 U4452 ( .A1(n3728), .A2(n3975), .A3(n3727), .A4(n3726), .ZN(n3738)
         );
  INV_X1 U4453 ( .A(n3866), .ZN(n3732) );
  NAND2_X1 U4454 ( .A1(n2379), .A2(DATAI_29_), .ZN(n3987) );
  INV_X1 U4455 ( .A(n3987), .ZN(n3985) );
  NAND2_X1 U4456 ( .A1(n2379), .A2(DATAI_31_), .ZN(n3802) );
  NAND2_X1 U4457 ( .A1(n4221), .A2(n3802), .ZN(n3805) );
  OR2_X1 U4458 ( .A1(n3980), .A2(n4219), .ZN(n3729) );
  NAND2_X1 U4459 ( .A1(n3805), .A2(n3729), .ZN(n3830) );
  AOI21_X1 U4460 ( .B1(n3732), .B2(n3985), .A(n3830), .ZN(n3733) );
  INV_X1 U4461 ( .A(n3733), .ZN(n3737) );
  INV_X1 U4462 ( .A(n3975), .ZN(n3731) );
  NOR2_X1 U4463 ( .A1(n3731), .A2(n3730), .ZN(n3734) );
  OAI21_X1 U4464 ( .B1(n3732), .B2(n3985), .A(n3974), .ZN(n3795) );
  OAI21_X1 U4465 ( .B1(n3734), .B2(n3795), .A(n3733), .ZN(n3799) );
  NOR3_X1 U4466 ( .A1(n3735), .A2(n3997), .A3(n3795), .ZN(n3736) );
  OAI22_X1 U4467 ( .A1(n3738), .A2(n3737), .B1(n3799), .B2(n3736), .ZN(n3739)
         );
  OAI21_X1 U4468 ( .B1(n4219), .B2(n4221), .A(n3739), .ZN(n3743) );
  AND2_X1 U4469 ( .A1(n3980), .A2(n4219), .ZN(n3801) );
  INV_X1 U4470 ( .A(n4221), .ZN(n3740) );
  INV_X1 U4471 ( .A(n3802), .ZN(n4222) );
  OAI21_X1 U4472 ( .B1(n3801), .B2(n3740), .A(n4222), .ZN(n3742) );
  AOI21_X1 U4473 ( .B1(n3743), .B2(n3742), .A(n3741), .ZN(n3855) );
  NOR2_X1 U4474 ( .A1(n3744), .A2(n4005), .ZN(n3798) );
  OAI211_X1 U4475 ( .C1(n3747), .C2(n4329), .A(n3746), .B(n3745), .ZN(n3749)
         );
  NAND3_X1 U4476 ( .A1(n3749), .A2(n3748), .A3(n2613), .ZN(n3752) );
  NAND3_X1 U4477 ( .A1(n3752), .A2(n3751), .A3(n3750), .ZN(n3755) );
  NAND3_X1 U4478 ( .A1(n3755), .A2(n3754), .A3(n3753), .ZN(n3758) );
  NAND3_X1 U4479 ( .A1(n3758), .A2(n3757), .A3(n3756), .ZN(n3761) );
  AOI21_X1 U4480 ( .B1(n3761), .B2(n3760), .A(n3759), .ZN(n3767) );
  NAND2_X1 U4481 ( .A1(n2071), .A2(n3763), .ZN(n3766) );
  OAI211_X1 U4482 ( .C1(n3767), .C2(n3766), .A(n3765), .B(n3764), .ZN(n3770)
         );
  NAND3_X1 U4483 ( .A1(n3770), .A2(n3769), .A3(n3768), .ZN(n3773) );
  AOI21_X1 U4484 ( .B1(n3773), .B2(n3772), .A(n2093), .ZN(n3780) );
  NAND2_X1 U4485 ( .A1(n3775), .A2(n3774), .ZN(n3779) );
  INV_X1 U4486 ( .A(n3776), .ZN(n3778) );
  OAI211_X1 U4487 ( .C1(n3780), .C2(n3779), .A(n3778), .B(n3777), .ZN(n3782)
         );
  NAND3_X1 U4488 ( .A1(n3782), .A2(n3781), .A3(n4192), .ZN(n3785) );
  INV_X1 U4489 ( .A(n3812), .ZN(n3783) );
  AOI21_X1 U4490 ( .B1(n3785), .B2(n3784), .A(n3783), .ZN(n3788) );
  INV_X1 U4491 ( .A(n4065), .ZN(n3821) );
  OAI211_X1 U4492 ( .C1(n3788), .C2(n3787), .A(n3786), .B(n3821), .ZN(n3789)
         );
  NAND2_X1 U4493 ( .A1(n3790), .A2(n3789), .ZN(n3793) );
  AOI211_X1 U4494 ( .C1(n3794), .C2(n3793), .A(n3792), .B(n3791), .ZN(n3797)
         );
  NOR4_X1 U4495 ( .A1(n3798), .A2(n3797), .A3(n3796), .A4(n3795), .ZN(n3800)
         );
  OR2_X1 U4496 ( .A1(n3800), .A2(n3799), .ZN(n3807) );
  INV_X1 U4497 ( .A(n3801), .ZN(n3804) );
  OR2_X1 U4498 ( .A1(n4221), .A2(n3802), .ZN(n3803) );
  NAND2_X1 U4499 ( .A1(n3804), .A2(n3803), .ZN(n3829) );
  NAND2_X1 U4500 ( .A1(n3829), .A2(n3805), .ZN(n3806) );
  NAND2_X1 U4501 ( .A1(n3807), .A2(n3806), .ZN(n3853) );
  NAND2_X1 U4502 ( .A1(n3809), .A2(n3808), .ZN(n4015) );
  INV_X1 U4503 ( .A(n4015), .ZN(n3848) );
  NAND2_X1 U4504 ( .A1(n4012), .A2(n3810), .ZN(n4033) );
  INV_X1 U4505 ( .A(n4033), .ZN(n3847) );
  NAND2_X1 U4506 ( .A1(n3811), .A2(n4048), .ZN(n4069) );
  NAND2_X1 U4507 ( .A1(n4146), .A2(n3812), .ZN(n4194) );
  NOR2_X1 U4508 ( .A1(n3814), .A2(n3813), .ZN(n3816) );
  NAND3_X1 U4509 ( .A1(n3817), .A2(n3816), .A3(n3815), .ZN(n3819) );
  NOR4_X1 U4510 ( .A1(n4069), .A2(n4194), .A3(n3819), .A4(n3818), .ZN(n3844)
         );
  NAND2_X1 U4511 ( .A1(n3820), .A2(n4030), .ZN(n4052) );
  NAND2_X1 U4512 ( .A1(n3821), .A2(n4066), .ZN(n4106) );
  INV_X1 U4513 ( .A(n4106), .ZN(n3825) );
  INV_X1 U4514 ( .A(n2612), .ZN(n3824) );
  INV_X1 U4515 ( .A(n3822), .ZN(n3823) );
  NAND4_X1 U4516 ( .A1(n3825), .A2(n3824), .A3(n2264), .A4(n3823), .ZN(n3826)
         );
  NOR2_X1 U4517 ( .A1(n4052), .A2(n3826), .ZN(n3843) );
  INV_X1 U4518 ( .A(n4454), .ZN(n3827) );
  NAND2_X1 U4519 ( .A1(n3828), .A2(n3827), .ZN(n3831) );
  NOR4_X1 U4520 ( .A1(n4095), .A2(n3831), .A3(n3830), .A4(n3829), .ZN(n3842)
         );
  INV_X1 U4521 ( .A(n4171), .ZN(n4174) );
  NAND4_X1 U4522 ( .A1(n3834), .A2(n3833), .A3(n4174), .A4(n3832), .ZN(n3840)
         );
  NAND4_X1 U4523 ( .A1(n3838), .A2(n3837), .A3(n3836), .A4(n3835), .ZN(n3839)
         );
  NOR2_X1 U4524 ( .A1(n3840), .A2(n3839), .ZN(n3841) );
  AND4_X1 U4525 ( .A1(n3844), .A2(n3843), .A3(n3842), .A4(n3841), .ZN(n3846)
         );
  XNOR2_X1 U4526 ( .A(n4154), .B(n4137), .ZN(n4125) );
  XNOR2_X1 U4527 ( .A(n4176), .B(n4160), .ZN(n4152) );
  NOR2_X1 U4528 ( .A1(n4125), .A2(n4152), .ZN(n3845) );
  NAND4_X1 U4529 ( .A1(n3848), .A2(n3847), .A3(n3846), .A4(n3845), .ZN(n3849)
         );
  XNOR2_X1 U4530 ( .A(n3866), .B(n3987), .ZN(n3979) );
  NOR3_X1 U4531 ( .A1(n3971), .A2(n3849), .A3(n3979), .ZN(n3851) );
  INV_X1 U4532 ( .A(n3997), .ZN(n3850) );
  AOI21_X1 U4533 ( .B1(n3851), .B2(n3850), .A(n4329), .ZN(n3852) );
  MUX2_X1 U4534 ( .A(n3853), .B(n3852), .S(n4330), .Z(n3854) );
  NOR2_X1 U4535 ( .A1(n3855), .A2(n3854), .ZN(n3856) );
  XNOR2_X1 U4536 ( .A(n3856), .B(n2611), .ZN(n3865) );
  INV_X1 U4537 ( .A(n3859), .ZN(n3864) );
  INV_X1 U4538 ( .A(n3857), .ZN(n3861) );
  NAND2_X1 U4539 ( .A1(n3859), .A2(n3858), .ZN(n3860) );
  OAI211_X1 U4540 ( .C1(n3862), .C2(n3861), .A(B_REG_SCAN_IN), .B(n3860), .ZN(
        n3863) );
  OAI21_X1 U4541 ( .B1(n3865), .B2(n3864), .A(n3863), .ZN(U3239) );
  MUX2_X1 U4542 ( .A(n4221), .B(DATAO_REG_31__SCAN_IN), .S(n3883), .Z(U3581)
         );
  INV_X2 U4543 ( .A(U4043), .ZN(n3883) );
  MUX2_X1 U4544 ( .A(n3866), .B(DATAO_REG_29__SCAN_IN), .S(n3883), .Z(U3579)
         );
  MUX2_X1 U4545 ( .A(n4001), .B(DATAO_REG_28__SCAN_IN), .S(n3883), .Z(U3578)
         );
  MUX2_X1 U4546 ( .A(n4054), .B(DATAO_REG_25__SCAN_IN), .S(n3883), .Z(U3575)
         );
  MUX2_X1 U4547 ( .A(n4073), .B(DATAO_REG_24__SCAN_IN), .S(n3883), .Z(U3574)
         );
  MUX2_X1 U4548 ( .A(n3867), .B(DATAO_REG_23__SCAN_IN), .S(n3883), .Z(U3573)
         );
  MUX2_X1 U4549 ( .A(n4154), .B(DATAO_REG_20__SCAN_IN), .S(n3883), .Z(U3570)
         );
  MUX2_X1 U4550 ( .A(n4176), .B(DATAO_REG_19__SCAN_IN), .S(n3883), .Z(U3569)
         );
  MUX2_X1 U4551 ( .A(n4201), .B(DATAO_REG_18__SCAN_IN), .S(n3883), .Z(U3568)
         );
  MUX2_X1 U4552 ( .A(n3868), .B(DATAO_REG_17__SCAN_IN), .S(n3883), .Z(U3567)
         );
  MUX2_X1 U4553 ( .A(n3869), .B(DATAO_REG_16__SCAN_IN), .S(n3883), .Z(U3566)
         );
  MUX2_X1 U4554 ( .A(n3870), .B(DATAO_REG_15__SCAN_IN), .S(n3883), .Z(U3565)
         );
  MUX2_X1 U4555 ( .A(n3871), .B(DATAO_REG_14__SCAN_IN), .S(n3883), .Z(U3564)
         );
  MUX2_X1 U4556 ( .A(n3872), .B(DATAO_REG_13__SCAN_IN), .S(n3883), .Z(U3563)
         );
  MUX2_X1 U4557 ( .A(n3873), .B(DATAO_REG_12__SCAN_IN), .S(n3883), .Z(U3562)
         );
  MUX2_X1 U4558 ( .A(n3874), .B(DATAO_REG_11__SCAN_IN), .S(n3883), .Z(U3561)
         );
  MUX2_X1 U4559 ( .A(n3875), .B(DATAO_REG_10__SCAN_IN), .S(n3883), .Z(U3560)
         );
  MUX2_X1 U4560 ( .A(n3876), .B(DATAO_REG_9__SCAN_IN), .S(n3883), .Z(U3559) );
  MUX2_X1 U4561 ( .A(n3877), .B(DATAO_REG_8__SCAN_IN), .S(n3883), .Z(U3558) );
  MUX2_X1 U4562 ( .A(n3878), .B(DATAO_REG_7__SCAN_IN), .S(n3883), .Z(U3557) );
  MUX2_X1 U4563 ( .A(n3879), .B(DATAO_REG_6__SCAN_IN), .S(n3883), .Z(U3556) );
  MUX2_X1 U4564 ( .A(n3880), .B(DATAO_REG_4__SCAN_IN), .S(n3883), .Z(U3554) );
  MUX2_X1 U4565 ( .A(n3881), .B(DATAO_REG_3__SCAN_IN), .S(n3883), .Z(U3553) );
  MUX2_X1 U4566 ( .A(n3882), .B(DATAO_REG_2__SCAN_IN), .S(n3883), .Z(U3552) );
  MUX2_X1 U4567 ( .A(n3884), .B(DATAO_REG_0__SCAN_IN), .S(n3883), .Z(U3550) );
  INV_X1 U4568 ( .A(n3885), .ZN(n3886) );
  OAI211_X1 U4569 ( .C1(n3888), .C2(n3887), .A(n4439), .B(n3886), .ZN(n3896)
         );
  MUX2_X1 U4570 ( .A(REG1_REG_1__SCAN_IN), .B(n2716), .S(n3889), .Z(n3890) );
  OAI21_X1 U4571 ( .B1(n2795), .B2(n3891), .A(n3890), .ZN(n3892) );
  NAND3_X1 U4572 ( .A1(n4427), .A2(n3899), .A3(n3892), .ZN(n3895) );
  NAND2_X1 U4573 ( .A1(n4403), .A2(n4336), .ZN(n3894) );
  AOI22_X1 U4574 ( .A1(n4434), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3893) );
  NAND4_X1 U4575 ( .A1(n3896), .A2(n3895), .A3(n3894), .A4(n3893), .ZN(U3241)
         );
  MUX2_X1 U4576 ( .A(REG1_REG_2__SCAN_IN), .B(n2713), .S(n3897), .Z(n3900) );
  NAND3_X1 U4577 ( .A1(n3900), .A2(n3899), .A3(n3898), .ZN(n3901) );
  AND3_X1 U4578 ( .A1(n3902), .A2(n4427), .A3(n3901), .ZN(n3907) );
  AOI211_X1 U4579 ( .C1(n3905), .C2(n3904), .A(n3903), .B(n4398), .ZN(n3906)
         );
  AOI211_X1 U4580 ( .C1(n4403), .C2(n4335), .A(n3907), .B(n3906), .ZN(n3910)
         );
  AOI22_X1 U4581 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4434), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3909) );
  NAND3_X1 U4582 ( .A1(n3910), .A2(n3909), .A3(n3908), .ZN(U3242) );
  INV_X1 U4583 ( .A(n4477), .ZN(n3925) );
  OAI21_X1 U4584 ( .B1(n3912), .B2(n3928), .A(n3911), .ZN(n3913) );
  AOI22_X1 U4585 ( .A1(n3925), .A2(n2432), .B1(REG1_REG_9__SCAN_IN), .B2(n4477), .ZN(n4346) );
  NOR2_X1 U4586 ( .A1(n3914), .A2(n4364), .ZN(n3915) );
  NOR2_X1 U4587 ( .A1(n4357), .A2(n4356), .ZN(n4355) );
  AOI22_X1 U4588 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4375), .B1(n4473), .B2(
        n2463), .ZN(n4366) );
  NOR2_X1 U4589 ( .A1(n4367), .A2(n4366), .ZN(n4365) );
  NOR2_X1 U4590 ( .A1(n3916), .A2(n4472), .ZN(n3917) );
  AOI22_X1 U4591 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4394), .B1(n4470), .B2(
        n4535), .ZN(n4386) );
  NOR2_X1 U4592 ( .A1(n3918), .A2(n3937), .ZN(n3919) );
  NOR2_X1 U4593 ( .A1(n4397), .A2(n4396), .ZN(n4395) );
  AOI22_X1 U4594 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4417), .B1(n4466), .B2(
        n3920), .ZN(n4408) );
  NOR2_X1 U4595 ( .A1(n4409), .A2(n4408), .ZN(n4407) );
  AND2_X1 U4596 ( .A1(n4466), .A2(REG1_REG_15__SCAN_IN), .ZN(n3921) );
  XOR2_X1 U4597 ( .A(n3956), .B(n3949), .Z(n3923) );
  OAI21_X1 U4598 ( .B1(n3923), .B2(n3922), .A(n3950), .ZN(n3924) );
  NAND2_X1 U4599 ( .A1(n3924), .A2(n4427), .ZN(n3947) );
  NAND2_X1 U4600 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4473), .ZN(n3932) );
  AOI22_X1 U4601 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4473), .B1(n4375), .B2(
        n3276), .ZN(n4372) );
  AOI22_X1 U4602 ( .A1(n3925), .A2(REG2_REG_9__SCAN_IN), .B1(n3108), .B2(n4477), .ZN(n4352) );
  NAND2_X1 U4603 ( .A1(n4475), .A2(n3930), .ZN(n3931) );
  XNOR2_X1 U4604 ( .A(n4364), .B(n3930), .ZN(n4361) );
  NAND2_X1 U4605 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4361), .ZN(n4360) );
  NAND2_X1 U4606 ( .A1(n3931), .A2(n4360), .ZN(n4371) );
  NAND2_X1 U4607 ( .A1(n4372), .A2(n4371), .ZN(n4370) );
  NAND2_X1 U4608 ( .A1(n3933), .A2(n3934), .ZN(n3935) );
  NAND2_X1 U4609 ( .A1(n3360), .A2(n4394), .ZN(n3936) );
  AOI22_X1 U4610 ( .A1(REG2_REG_13__SCAN_IN), .A2(n4470), .B1(n4390), .B2(
        n3936), .ZN(n3938) );
  NOR2_X1 U4611 ( .A1(n3938), .A2(n3937), .ZN(n3939) );
  AOI22_X1 U4612 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4417), .B1(n4466), .B2(
        n3414), .ZN(n4413) );
  AND2_X1 U4613 ( .A1(n4466), .A2(REG2_REG_15__SCAN_IN), .ZN(n3940) );
  NOR2_X1 U4614 ( .A1(n4412), .A2(n3940), .ZN(n3957) );
  OAI21_X1 U4615 ( .B1(n3941), .B2(n3424), .A(n3958), .ZN(n3945) );
  NAND2_X1 U4616 ( .A1(n4434), .A2(ADDR_REG_16__SCAN_IN), .ZN(n3942) );
  OAI211_X1 U4617 ( .C1(n4442), .C2(n3956), .A(n3943), .B(n3942), .ZN(n3944)
         );
  AOI21_X1 U4618 ( .B1(n3945), .B2(n4439), .A(n3944), .ZN(n3946) );
  NAND2_X1 U4619 ( .A1(n3947), .A2(n3946), .ZN(U3256) );
  INV_X1 U4620 ( .A(n3961), .ZN(n4463) );
  AOI22_X1 U4621 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4463), .B1(n3961), .B2(
        n3948), .ZN(n4432) );
  AOI22_X1 U4622 ( .A1(n3960), .A2(REG1_REG_17__SCAN_IN), .B1(n4273), .B2(
        n4465), .ZN(n4421) );
  NAND2_X1 U4623 ( .A1(n3949), .A2(n3956), .ZN(n3951) );
  NAND2_X1 U4624 ( .A1(n3951), .A2(n3950), .ZN(n4420) );
  XNOR2_X1 U4625 ( .A(n2611), .B(REG1_REG_19__SCAN_IN), .ZN(n3952) );
  XNOR2_X1 U4626 ( .A(n3953), .B(n3952), .ZN(n3969) );
  NAND2_X1 U4627 ( .A1(REG2_REG_18__SCAN_IN), .A2(n3961), .ZN(n3954) );
  OAI21_X1 U4628 ( .B1(REG2_REG_18__SCAN_IN), .B2(n3961), .A(n3954), .ZN(n4437) );
  NOR2_X1 U4629 ( .A1(n3960), .A2(REG2_REG_17__SCAN_IN), .ZN(n3955) );
  AOI21_X1 U4630 ( .B1(REG2_REG_17__SCAN_IN), .B2(n3960), .A(n3955), .ZN(n4424) );
  NAND2_X1 U4631 ( .A1(n3957), .A2(n3956), .ZN(n3959) );
  OAI21_X1 U4632 ( .B1(n3960), .B2(REG2_REG_17__SCAN_IN), .A(n4422), .ZN(n4436) );
  NOR2_X1 U4633 ( .A1(n4437), .A2(n4436), .ZN(n4435) );
  AOI21_X1 U4634 ( .B1(n3961), .B2(REG2_REG_18__SCAN_IN), .A(n4435), .ZN(n3963) );
  MUX2_X1 U4635 ( .A(REG2_REG_19__SCAN_IN), .B(n4165), .S(n2611), .Z(n3962) );
  XNOR2_X1 U4636 ( .A(n3963), .B(n3962), .ZN(n3967) );
  NAND2_X1 U4637 ( .A1(n4434), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3964) );
  OAI211_X1 U4638 ( .C1(n4442), .C2(n2838), .A(n3965), .B(n3964), .ZN(n3966)
         );
  AOI21_X1 U4639 ( .B1(n3967), .B2(n4439), .A(n3966), .ZN(n3968) );
  OAI21_X1 U4640 ( .B1(n3969), .B2(n4430), .A(n3968), .ZN(U3259) );
  AOI22_X1 U4641 ( .A1(n3972), .A2(n3971), .B1(n3970), .B2(n4001), .ZN(n3973)
         );
  XNOR2_X1 U4642 ( .A(n3973), .B(n3979), .ZN(n4230) );
  INV_X1 U4643 ( .A(n4230), .ZN(n3993) );
  INV_X1 U4644 ( .A(n3974), .ZN(n3976) );
  OAI21_X1 U4645 ( .B1(n3977), .B2(n3976), .A(n3975), .ZN(n3978) );
  AOI21_X1 U4646 ( .B1(B_REG_SCAN_IN), .B2(n4326), .A(n4090), .ZN(n4220) );
  AOI22_X1 U4647 ( .A1(n3980), .A2(n4220), .B1(n4227), .B2(n3985), .ZN(n3981)
         );
  OAI21_X1 U4648 ( .B1(n3982), .B2(n4204), .A(n3981), .ZN(n3983) );
  OAI21_X1 U4649 ( .B1(n3984), .B2(n4211), .A(n4232), .ZN(n3991) );
  INV_X1 U4650 ( .A(n3986), .ZN(n3988) );
  OAI22_X1 U4651 ( .A1(n4231), .A2(n4210), .B1(n3989), .B2(n4136), .ZN(n3990)
         );
  AOI21_X1 U4652 ( .B1(n3991), .B2(n4188), .A(n3990), .ZN(n3992) );
  OAI21_X1 U4653 ( .B1(n3993), .B2(n4217), .A(n3992), .ZN(U3354) );
  XOR2_X1 U4654 ( .A(n3997), .B(n3994), .Z(n4236) );
  AOI21_X1 U4655 ( .B1(n3997), .B2(n3996), .A(n3995), .ZN(n4003) );
  OAI22_X1 U4656 ( .A1(n3999), .A2(n4204), .B1(n3998), .B2(n4198), .ZN(n4000)
         );
  AOI21_X1 U4657 ( .B1(n4001), .B2(n4200), .A(n4000), .ZN(n4002) );
  OAI21_X1 U4658 ( .B1(n4003), .B2(n4158), .A(n4002), .ZN(n4233) );
  AOI21_X1 U4659 ( .B1(n4005), .B2(n2041), .A(n4004), .ZN(n4234) );
  INV_X1 U4660 ( .A(n4234), .ZN(n4008) );
  AOI22_X1 U4661 ( .A1(n4006), .A2(n4453), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4458), .ZN(n4007) );
  OAI21_X1 U4662 ( .B1(n4008), .B2(n4210), .A(n4007), .ZN(n4009) );
  AOI21_X1 U4663 ( .B1(n4233), .B2(n4188), .A(n4009), .ZN(n4010) );
  OAI21_X1 U4664 ( .B1(n4236), .B2(n4217), .A(n4010), .ZN(U3263) );
  XOR2_X1 U4665 ( .A(n4015), .B(n4011), .Z(n4238) );
  INV_X1 U4666 ( .A(n4238), .ZN(n4028) );
  INV_X1 U4667 ( .A(n4031), .ZN(n4014) );
  OAI21_X1 U4668 ( .B1(n4014), .B2(n4013), .A(n4012), .ZN(n4016) );
  XNOR2_X1 U4669 ( .A(n4016), .B(n4015), .ZN(n4021) );
  OAI22_X1 U4670 ( .A1(n4017), .A2(n4204), .B1(n4022), .B2(n4198), .ZN(n4018)
         );
  AOI21_X1 U4671 ( .B1(n4200), .B2(n4019), .A(n4018), .ZN(n4020) );
  OAI21_X1 U4672 ( .B1(n4021), .B2(n4158), .A(n4020), .ZN(n4237) );
  INV_X1 U4673 ( .A(n4039), .ZN(n4023) );
  OAI21_X1 U4674 ( .B1(n4023), .B2(n4022), .A(n2041), .ZN(n4292) );
  AOI22_X1 U4675 ( .A1(n4024), .A2(n4453), .B1(n4458), .B2(
        REG2_REG_26__SCAN_IN), .ZN(n4025) );
  OAI21_X1 U4676 ( .B1(n4292), .B2(n4210), .A(n4025), .ZN(n4026) );
  AOI21_X1 U4677 ( .B1(n4237), .B2(n4136), .A(n4026), .ZN(n4027) );
  OAI21_X1 U4678 ( .B1(n4028), .B2(n4217), .A(n4027), .ZN(U3264) );
  XNOR2_X1 U4679 ( .A(n4029), .B(n4033), .ZN(n4241) );
  INV_X1 U4680 ( .A(n4241), .ZN(n4046) );
  NAND2_X1 U4681 ( .A1(n4031), .A2(n4030), .ZN(n4032) );
  XOR2_X1 U4682 ( .A(n4033), .B(n4032), .Z(n4038) );
  OAI22_X1 U4683 ( .A1(n4034), .A2(n4204), .B1(n4040), .B2(n4198), .ZN(n4035)
         );
  AOI21_X1 U4684 ( .B1(n4200), .B2(n4036), .A(n4035), .ZN(n4037) );
  OAI21_X1 U4685 ( .B1(n4038), .B2(n4158), .A(n4037), .ZN(n4240) );
  INV_X1 U4686 ( .A(n4057), .ZN(n4041) );
  OAI21_X1 U4687 ( .B1(n4041), .B2(n4040), .A(n4039), .ZN(n4295) );
  AOI22_X1 U4688 ( .A1(REG2_REG_25__SCAN_IN), .A2(n4458), .B1(n4042), .B2(
        n4453), .ZN(n4043) );
  OAI21_X1 U4689 ( .B1(n4295), .B2(n4210), .A(n4043), .ZN(n4044) );
  AOI21_X1 U4690 ( .B1(n4240), .B2(n4188), .A(n4044), .ZN(n4045) );
  OAI21_X1 U4691 ( .B1(n4046), .B2(n4217), .A(n4045), .ZN(U3265) );
  XOR2_X1 U4692 ( .A(n4052), .B(n4047), .Z(n4245) );
  INV_X1 U4693 ( .A(n4245), .ZN(n4063) );
  INV_X1 U4694 ( .A(n4048), .ZN(n4049) );
  NOR2_X1 U4695 ( .A1(n4050), .A2(n4049), .ZN(n4051) );
  XOR2_X1 U4696 ( .A(n4052), .B(n4051), .Z(n4056) );
  OAI22_X1 U4697 ( .A1(n4091), .A2(n4204), .B1(n4198), .B2(n4058), .ZN(n4053)
         );
  AOI21_X1 U4698 ( .B1(n4054), .B2(n4200), .A(n4053), .ZN(n4055) );
  OAI21_X1 U4699 ( .B1(n4056), .B2(n4158), .A(n4055), .ZN(n4244) );
  OAI21_X1 U4700 ( .B1(n4076), .B2(n4058), .A(n4057), .ZN(n4298) );
  AOI22_X1 U4701 ( .A1(n4458), .A2(REG2_REG_24__SCAN_IN), .B1(n4059), .B2(
        n4453), .ZN(n4060) );
  OAI21_X1 U4702 ( .B1(n4298), .B2(n4210), .A(n4060), .ZN(n4061) );
  AOI21_X1 U4703 ( .B1(n4244), .B2(n4188), .A(n4061), .ZN(n4062) );
  OAI21_X1 U4704 ( .B1(n4063), .B2(n4217), .A(n4062), .ZN(U3266) );
  XOR2_X1 U4705 ( .A(n4069), .B(n4064), .Z(n4249) );
  INV_X1 U4706 ( .A(n4249), .ZN(n4085) );
  OR2_X1 U4707 ( .A1(n4105), .A2(n4065), .ZN(n4067) );
  NAND2_X1 U4708 ( .A1(n4067), .A2(n4066), .ZN(n4087) );
  INV_X1 U4709 ( .A(n4095), .ZN(n4088) );
  NAND2_X1 U4710 ( .A1(n4087), .A2(n4088), .ZN(n4086) );
  NAND2_X1 U4711 ( .A1(n4086), .A2(n4068), .ZN(n4070) );
  XNOR2_X1 U4712 ( .A(n4070), .B(n4069), .ZN(n4075) );
  OAI22_X1 U4713 ( .A1(n4071), .A2(n4204), .B1(n4198), .B2(n4078), .ZN(n4072)
         );
  AOI21_X1 U4714 ( .B1(n4200), .B2(n4073), .A(n4072), .ZN(n4074) );
  OAI21_X1 U4715 ( .B1(n4075), .B2(n4158), .A(n4074), .ZN(n4248) );
  INV_X1 U4716 ( .A(n4253), .ZN(n4079) );
  INV_X1 U4717 ( .A(n4076), .ZN(n4077) );
  OAI21_X1 U4718 ( .B1(n4079), .B2(n4078), .A(n4077), .ZN(n4302) );
  NOR2_X1 U4719 ( .A1(n4302), .A2(n4210), .ZN(n4083) );
  OAI22_X1 U4720 ( .A1(n4136), .A2(n4081), .B1(n4080), .B2(n4211), .ZN(n4082)
         );
  AOI211_X1 U4721 ( .C1(n4248), .C2(n4188), .A(n4083), .B(n4082), .ZN(n4084)
         );
  OAI21_X1 U4722 ( .B1(n4085), .B2(n4217), .A(n4084), .ZN(U3267) );
  OAI21_X1 U4723 ( .B1(n4088), .B2(n4087), .A(n4086), .ZN(n4093) );
  AOI22_X1 U4724 ( .A1(n4129), .A2(n4155), .B1(n4097), .B2(n4227), .ZN(n4089)
         );
  OAI21_X1 U4725 ( .B1(n4091), .B2(n4090), .A(n4089), .ZN(n4092) );
  AOI21_X1 U4726 ( .B1(n4093), .B2(n4196), .A(n4092), .ZN(n4255) );
  OAI21_X1 U4727 ( .B1(n4096), .B2(n4095), .A(n4094), .ZN(n4256) );
  OR2_X1 U4728 ( .A1(n4256), .A2(n4217), .ZN(n4103) );
  NAND2_X1 U4729 ( .A1(n2018), .A2(n4097), .ZN(n4252) );
  AND2_X1 U4730 ( .A1(n4252), .A2(n4446), .ZN(n4101) );
  INV_X1 U4731 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4099) );
  OAI22_X1 U4732 ( .A1(n4136), .A2(n4099), .B1(n4098), .B2(n4211), .ZN(n4100)
         );
  AOI21_X1 U4733 ( .B1(n4101), .B2(n4253), .A(n4100), .ZN(n4102) );
  OAI211_X1 U4734 ( .C1(n4458), .C2(n4255), .A(n4103), .B(n4102), .ZN(U3268)
         );
  XOR2_X1 U4735 ( .A(n4106), .B(n4104), .Z(n4258) );
  INV_X1 U4736 ( .A(n4258), .ZN(n4120) );
  XOR2_X1 U4737 ( .A(n4106), .B(n4105), .Z(n4112) );
  OAI22_X1 U4738 ( .A1(n4108), .A2(n4204), .B1(n4107), .B2(n4198), .ZN(n4109)
         );
  AOI21_X1 U4739 ( .B1(n4200), .B2(n4110), .A(n4109), .ZN(n4111) );
  OAI21_X1 U4740 ( .B1(n4112), .B2(n4158), .A(n4111), .ZN(n4257) );
  NAND2_X1 U4741 ( .A1(n2013), .A2(n4113), .ZN(n4114) );
  NAND2_X1 U4742 ( .A1(n2018), .A2(n4114), .ZN(n4307) );
  INV_X1 U4743 ( .A(n4115), .ZN(n4116) );
  AOI22_X1 U4744 ( .A1(n4458), .A2(REG2_REG_21__SCAN_IN), .B1(n4116), .B2(
        n4453), .ZN(n4117) );
  OAI21_X1 U4745 ( .B1(n4307), .B2(n4210), .A(n4117), .ZN(n4118) );
  AOI21_X1 U4746 ( .B1(n4257), .B2(n4188), .A(n4118), .ZN(n4119) );
  OAI21_X1 U4747 ( .B1(n4120), .B2(n4217), .A(n4119), .ZN(U3269) );
  XNOR2_X1 U4748 ( .A(n2183), .B(n4125), .ZN(n4260) );
  INV_X1 U4749 ( .A(n4122), .ZN(n4124) );
  OAI21_X1 U4750 ( .B1(n4147), .B2(n4124), .A(n4123), .ZN(n4127) );
  INV_X1 U4751 ( .A(n4125), .ZN(n4126) );
  XNOR2_X1 U4752 ( .A(n4127), .B(n4126), .ZN(n4133) );
  AOI22_X1 U4753 ( .A1(n4129), .A2(n4200), .B1(n4227), .B2(n4128), .ZN(n4130)
         );
  OAI21_X1 U4754 ( .B1(n4131), .B2(n4204), .A(n4130), .ZN(n4132) );
  AOI21_X1 U4755 ( .B1(n4133), .B2(n4196), .A(n4132), .ZN(n4134) );
  OAI21_X1 U4756 ( .B1(n4260), .B2(n4135), .A(n4134), .ZN(n4261) );
  NAND2_X1 U4757 ( .A1(n4261), .A2(n4136), .ZN(n4143) );
  OAI21_X1 U4758 ( .B1(n4163), .B2(n4137), .A(n2013), .ZN(n4311) );
  INV_X1 U4759 ( .A(n4311), .ZN(n4141) );
  INV_X1 U4760 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4139) );
  OAI22_X1 U4761 ( .A1(n4136), .A2(n4139), .B1(n4138), .B2(n4211), .ZN(n4140)
         );
  AOI21_X1 U4762 ( .B1(n4141), .B2(n4446), .A(n4140), .ZN(n4142) );
  OAI211_X1 U4763 ( .C1(n4260), .C2(n4144), .A(n4143), .B(n4142), .ZN(U3270)
         );
  XNOR2_X1 U4764 ( .A(n4145), .B(n4152), .ZN(n4266) );
  INV_X1 U4765 ( .A(n4266), .ZN(n4169) );
  NAND2_X1 U4766 ( .A1(n4147), .A2(n4146), .ZN(n4175) );
  INV_X1 U4767 ( .A(n4148), .ZN(n4150) );
  OAI21_X1 U4768 ( .B1(n4175), .B2(n4150), .A(n4149), .ZN(n4151) );
  XOR2_X1 U4769 ( .A(n4152), .B(n4151), .Z(n4159) );
  NOR2_X1 U4770 ( .A1(n4198), .A2(n4160), .ZN(n4153) );
  AOI21_X1 U4771 ( .B1(n4154), .B2(n4200), .A(n4153), .ZN(n4157) );
  NAND2_X1 U4772 ( .A1(n4201), .A2(n4155), .ZN(n4156) );
  OAI211_X1 U4773 ( .C1(n4159), .C2(n4158), .A(n4157), .B(n4156), .ZN(n4265)
         );
  AOI21_X1 U4774 ( .B1(n4206), .B2(n4161), .A(n4160), .ZN(n4162) );
  OR2_X1 U4775 ( .A1(n4163), .A2(n4162), .ZN(n4315) );
  NOR2_X1 U4776 ( .A1(n4315), .A2(n4210), .ZN(n4167) );
  OAI22_X1 U4777 ( .A1(n4136), .A2(n4165), .B1(n4164), .B2(n4211), .ZN(n4166)
         );
  AOI211_X1 U4778 ( .C1(n4265), .C2(n4188), .A(n4167), .B(n4166), .ZN(n4168)
         );
  OAI21_X1 U4779 ( .B1(n4169), .B2(n4217), .A(n4168), .ZN(U3271) );
  OAI21_X1 U4780 ( .B1(n4172), .B2(n4171), .A(n4170), .ZN(n4173) );
  INV_X1 U4781 ( .A(n4173), .ZN(n4270) );
  XNOR2_X1 U4782 ( .A(n4175), .B(n4174), .ZN(n4180) );
  AOI22_X1 U4783 ( .A1(n4176), .A2(n4200), .B1(n4227), .B2(n4181), .ZN(n4177)
         );
  OAI21_X1 U4784 ( .B1(n4178), .B2(n4204), .A(n4177), .ZN(n4179) );
  AOI21_X1 U4785 ( .B1(n4180), .B2(n4196), .A(n4179), .ZN(n4269) );
  INV_X1 U4786 ( .A(n4269), .ZN(n4189) );
  XNOR2_X1 U4787 ( .A(n4206), .B(n4181), .ZN(n4182) );
  NAND2_X1 U4788 ( .A1(n4182), .A2(n4489), .ZN(n4268) );
  NOR2_X1 U4789 ( .A1(n4268), .A2(n4183), .ZN(n4187) );
  INV_X1 U4790 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4185) );
  OAI22_X1 U4791 ( .A1(n4188), .A2(n4185), .B1(n4184), .B2(n4211), .ZN(n4186)
         );
  AOI211_X1 U4792 ( .C1(n4189), .C2(n4188), .A(n4187), .B(n4186), .ZN(n4190)
         );
  OAI21_X1 U4793 ( .B1(n4270), .B2(n4217), .A(n4190), .ZN(U3272) );
  XOR2_X1 U4794 ( .A(n4194), .B(n4191), .Z(n4272) );
  INV_X1 U4795 ( .A(n4272), .ZN(n4218) );
  NAND2_X1 U4796 ( .A1(n4193), .A2(n4192), .ZN(n4195) );
  XNOR2_X1 U4797 ( .A(n4195), .B(n4194), .ZN(n4197) );
  NAND2_X1 U4798 ( .A1(n4197), .A2(n4196), .ZN(n4203) );
  NOR2_X1 U4799 ( .A1(n4198), .A2(n4208), .ZN(n4199) );
  AOI21_X1 U4800 ( .B1(n4201), .B2(n4200), .A(n4199), .ZN(n4202) );
  OAI211_X1 U4801 ( .C1(n4205), .C2(n4204), .A(n4203), .B(n4202), .ZN(n4271)
         );
  INV_X1 U4802 ( .A(n4206), .ZN(n4207) );
  OAI21_X1 U4803 ( .B1(n4209), .B2(n4208), .A(n4207), .ZN(n4321) );
  NOR2_X1 U4804 ( .A1(n4321), .A2(n4210), .ZN(n4215) );
  OAI22_X1 U4805 ( .A1(n4136), .A2(n4213), .B1(n4212), .B2(n4211), .ZN(n4214)
         );
  AOI211_X1 U4806 ( .C1(n4271), .C2(n4136), .A(n4215), .B(n4214), .ZN(n4216)
         );
  OAI21_X1 U4807 ( .B1(n4218), .B2(n4217), .A(n4216), .ZN(U3273) );
  XNOR2_X1 U4808 ( .A(n4224), .B(n4222), .ZN(n4339) );
  INV_X1 U4809 ( .A(n4339), .ZN(n4285) );
  AND2_X1 U4810 ( .A1(n4221), .A2(n4220), .ZN(n4226) );
  AOI21_X1 U4811 ( .B1(n4222), .B2(n4227), .A(n4226), .ZN(n4341) );
  MUX2_X1 U4812 ( .A(n3707), .B(n4341), .S(n4524), .Z(n4223) );
  OAI21_X1 U4813 ( .B1(n4285), .B2(n4275), .A(n4223), .ZN(U3549) );
  AOI21_X1 U4814 ( .B1(n4228), .B2(n4225), .A(n4224), .ZN(n4342) );
  INV_X1 U4815 ( .A(n4342), .ZN(n4287) );
  AOI21_X1 U4816 ( .B1(n4228), .B2(n4227), .A(n4226), .ZN(n4344) );
  MUX2_X1 U4817 ( .A(n2724), .B(n4344), .S(n4524), .Z(n4229) );
  OAI21_X1 U4818 ( .B1(n4287), .B2(n4275), .A(n4229), .ZN(U3548) );
  MUX2_X1 U4819 ( .A(REG1_REG_29__SCAN_IN), .B(n4288), .S(n4524), .Z(U3547) );
  AOI21_X1 U4820 ( .B1(n4489), .B2(n4234), .A(n4233), .ZN(n4235) );
  OAI21_X1 U4821 ( .B1(n4236), .B2(n4501), .A(n4235), .ZN(n4289) );
  MUX2_X1 U4822 ( .A(REG1_REG_27__SCAN_IN), .B(n4289), .S(n4524), .Z(U3545) );
  AOI21_X1 U4823 ( .B1(n4238), .B2(n4512), .A(n4237), .ZN(n4290) );
  MUX2_X1 U4824 ( .A(n4546), .B(n4290), .S(n4524), .Z(n4239) );
  OAI21_X1 U4825 ( .B1(n4275), .B2(n4292), .A(n4239), .ZN(U3544) );
  INV_X1 U4826 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4242) );
  AOI21_X1 U4827 ( .B1(n4241), .B2(n4512), .A(n4240), .ZN(n4293) );
  MUX2_X1 U4828 ( .A(n4242), .B(n4293), .S(n4524), .Z(n4243) );
  OAI21_X1 U4829 ( .B1(n4275), .B2(n4295), .A(n4243), .ZN(U3543) );
  INV_X1 U4830 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4246) );
  AOI21_X1 U4831 ( .B1(n4245), .B2(n4512), .A(n4244), .ZN(n4296) );
  MUX2_X1 U4832 ( .A(n4246), .B(n4296), .S(n4524), .Z(n4247) );
  OAI21_X1 U4833 ( .B1(n4275), .B2(n4298), .A(n4247), .ZN(U3542) );
  INV_X1 U4834 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4250) );
  AOI21_X1 U4835 ( .B1(n4249), .B2(n4512), .A(n4248), .ZN(n4299) );
  MUX2_X1 U4836 ( .A(n4250), .B(n4299), .S(n4524), .Z(n4251) );
  OAI21_X1 U4837 ( .B1(n4275), .B2(n4302), .A(n4251), .ZN(U3541) );
  NAND3_X1 U4838 ( .A1(n4253), .A2(n4489), .A3(n4252), .ZN(n4254) );
  OAI211_X1 U4839 ( .C1(n4256), .C2(n4501), .A(n4255), .B(n4254), .ZN(n4303)
         );
  MUX2_X1 U4840 ( .A(REG1_REG_22__SCAN_IN), .B(n4303), .S(n4524), .Z(U3540) );
  INV_X1 U4841 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4542) );
  AOI21_X1 U4842 ( .B1(n4258), .B2(n4512), .A(n4257), .ZN(n4304) );
  MUX2_X1 U4843 ( .A(n4542), .B(n4304), .S(n4524), .Z(n4259) );
  OAI21_X1 U4844 ( .B1(n4275), .B2(n4307), .A(n4259), .ZN(U3539) );
  INV_X1 U4845 ( .A(n4260), .ZN(n4262) );
  AOI21_X1 U4846 ( .B1(n4495), .B2(n4262), .A(n4261), .ZN(n4308) );
  MUX2_X1 U4847 ( .A(n4263), .B(n4308), .S(n4524), .Z(n4264) );
  OAI21_X1 U4848 ( .B1(n4275), .B2(n4311), .A(n4264), .ZN(U3538) );
  AOI21_X1 U4849 ( .B1(n4266), .B2(n4512), .A(n4265), .ZN(n4312) );
  MUX2_X1 U4850 ( .A(n4543), .B(n4312), .S(n4524), .Z(n4267) );
  OAI21_X1 U4851 ( .B1(n4275), .B2(n4315), .A(n4267), .ZN(U3537) );
  OAI211_X1 U4852 ( .C1(n4270), .C2(n4501), .A(n4269), .B(n4268), .ZN(n4316)
         );
  MUX2_X1 U4853 ( .A(REG1_REG_18__SCAN_IN), .B(n4316), .S(n4524), .Z(U3536) );
  AOI21_X1 U4854 ( .B1(n4272), .B2(n4512), .A(n4271), .ZN(n4317) );
  MUX2_X1 U4855 ( .A(n4273), .B(n4317), .S(n4524), .Z(n4274) );
  OAI21_X1 U4856 ( .B1(n4275), .B2(n4321), .A(n4274), .ZN(U3535) );
  AOI21_X1 U4857 ( .B1(n4489), .B2(n4277), .A(n4276), .ZN(n4278) );
  OAI21_X1 U4858 ( .B1(n4279), .B2(n4501), .A(n4278), .ZN(n4322) );
  MUX2_X1 U4859 ( .A(REG1_REG_16__SCAN_IN), .B(n4322), .S(n4524), .Z(U3534) );
  NAND2_X1 U4860 ( .A1(n4280), .A2(n4512), .ZN(n4282) );
  OAI211_X1 U4861 ( .C1(n4283), .C2(n4510), .A(n4282), .B(n4281), .ZN(n4323)
         );
  MUX2_X1 U4862 ( .A(REG1_REG_15__SCAN_IN), .B(n4323), .S(n4524), .Z(U3533) );
  INV_X1 U4863 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4532) );
  MUX2_X1 U4864 ( .A(n4532), .B(n4341), .S(n4516), .Z(n4284) );
  OAI21_X1 U4865 ( .B1(n4285), .B2(n4320), .A(n4284), .ZN(U3517) );
  INV_X1 U4866 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4533) );
  MUX2_X1 U4867 ( .A(n4533), .B(n4344), .S(n4516), .Z(n4286) );
  OAI21_X1 U4868 ( .B1(n4287), .B2(n4320), .A(n4286), .ZN(U3516) );
  MUX2_X1 U4869 ( .A(REG0_REG_29__SCAN_IN), .B(n4288), .S(n4516), .Z(U3515) );
  MUX2_X1 U4870 ( .A(REG0_REG_27__SCAN_IN), .B(n4289), .S(n4516), .Z(U3513) );
  MUX2_X1 U4871 ( .A(n4529), .B(n4290), .S(n4516), .Z(n4291) );
  OAI21_X1 U4872 ( .B1(n4292), .B2(n4320), .A(n4291), .ZN(U3512) );
  MUX2_X1 U4873 ( .A(n4530), .B(n4293), .S(n4516), .Z(n4294) );
  OAI21_X1 U4874 ( .B1(n4295), .B2(n4320), .A(n4294), .ZN(U3511) );
  MUX2_X1 U4875 ( .A(n4526), .B(n4296), .S(n4516), .Z(n4297) );
  OAI21_X1 U4876 ( .B1(n4298), .B2(n4320), .A(n4297), .ZN(U3510) );
  INV_X1 U4877 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4300) );
  MUX2_X1 U4878 ( .A(n4300), .B(n4299), .S(n4516), .Z(n4301) );
  OAI21_X1 U4879 ( .B1(n4302), .B2(n4320), .A(n4301), .ZN(U3509) );
  MUX2_X1 U4880 ( .A(REG0_REG_22__SCAN_IN), .B(n4303), .S(n4516), .Z(U3508) );
  INV_X1 U4881 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4305) );
  MUX2_X1 U4882 ( .A(n4305), .B(n4304), .S(n4516), .Z(n4306) );
  OAI21_X1 U4883 ( .B1(n4307), .B2(n4320), .A(n4306), .ZN(U3507) );
  INV_X1 U4884 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4309) );
  MUX2_X1 U4885 ( .A(n4309), .B(n4308), .S(n4516), .Z(n4310) );
  OAI21_X1 U4886 ( .B1(n4311), .B2(n4320), .A(n4310), .ZN(U3506) );
  INV_X1 U4887 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4313) );
  MUX2_X1 U4888 ( .A(n4313), .B(n4312), .S(n4516), .Z(n4314) );
  OAI21_X1 U4889 ( .B1(n4315), .B2(n4320), .A(n4314), .ZN(U3505) );
  MUX2_X1 U4890 ( .A(REG0_REG_18__SCAN_IN), .B(n4316), .S(n4516), .Z(U3503) );
  INV_X1 U4891 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4318) );
  MUX2_X1 U4892 ( .A(n4318), .B(n4317), .S(n4516), .Z(n4319) );
  OAI21_X1 U4893 ( .B1(n4321), .B2(n4320), .A(n4319), .ZN(U3501) );
  MUX2_X1 U4894 ( .A(REG0_REG_16__SCAN_IN), .B(n4322), .S(n4516), .Z(U3499) );
  MUX2_X1 U4895 ( .A(REG0_REG_15__SCAN_IN), .B(n4323), .S(n4516), .Z(U3497) );
  MUX2_X1 U4896 ( .A(DATAI_30_), .B(n4324), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U4897 ( .A(DATAI_29_), .B(n4325), .S(STATE_REG_SCAN_IN), .Z(U3323)
         );
  MUX2_X1 U4898 ( .A(DATAI_27_), .B(n4326), .S(STATE_REG_SCAN_IN), .Z(U3325)
         );
  MUX2_X1 U4899 ( .A(DATAI_26_), .B(n4327), .S(STATE_REG_SCAN_IN), .Z(U3326)
         );
  MUX2_X1 U4900 ( .A(n2665), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U4901 ( .A(n4328), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U4902 ( .A(n4329), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U4903 ( .A(DATAI_20_), .B(n4330), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  INV_X1 U4904 ( .A(n4331), .ZN(n4332) );
  MUX2_X1 U4905 ( .A(DATAI_7_), .B(n4332), .S(STATE_REG_SCAN_IN), .Z(U3345) );
  MUX2_X1 U4906 ( .A(n4333), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U4907 ( .A(DATAI_3_), .B(n4334), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U4908 ( .A(n4335), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U4909 ( .A(n4336), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  OAI22_X1 U4910 ( .A1(U3149), .A2(n4337), .B1(DATAI_28_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4338) );
  INV_X1 U4911 ( .A(n4338), .ZN(U3324) );
  AOI22_X1 U4912 ( .A1(n4339), .A2(n4446), .B1(n4458), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n4340) );
  OAI21_X1 U4913 ( .B1(n4458), .B2(n4341), .A(n4340), .ZN(U3260) );
  AOI22_X1 U4914 ( .A1(n4342), .A2(n4446), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4458), .ZN(n4343) );
  OAI21_X1 U4915 ( .B1(n4458), .B2(n4344), .A(n4343), .ZN(U3261) );
  AOI211_X1 U4916 ( .C1(n4347), .C2(n4346), .A(n4345), .B(n4430), .ZN(n4349)
         );
  AOI211_X1 U4917 ( .C1(n4434), .C2(ADDR_REG_9__SCAN_IN), .A(n4349), .B(n4348), 
        .ZN(n4354) );
  OAI211_X1 U4918 ( .C1(n4352), .C2(n4351), .A(n4439), .B(n4350), .ZN(n4353)
         );
  OAI211_X1 U4919 ( .C1(n4442), .C2(n4477), .A(n4354), .B(n4353), .ZN(U3249)
         );
  AOI211_X1 U4920 ( .C1(n4357), .C2(n4356), .A(n4355), .B(n4430), .ZN(n4359)
         );
  AOI211_X1 U4921 ( .C1(n4434), .C2(ADDR_REG_10__SCAN_IN), .A(n4359), .B(n4358), .ZN(n4363) );
  OAI211_X1 U4922 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4361), .A(n4439), .B(n4360), .ZN(n4362) );
  OAI211_X1 U4923 ( .C1(n4442), .C2(n4364), .A(n4363), .B(n4362), .ZN(U3250)
         );
  AOI211_X1 U4924 ( .C1(n4367), .C2(n4366), .A(n4365), .B(n4430), .ZN(n4369)
         );
  AOI211_X1 U4925 ( .C1(n4434), .C2(ADDR_REG_11__SCAN_IN), .A(n4369), .B(n4368), .ZN(n4374) );
  OAI211_X1 U4926 ( .C1(n4372), .C2(n4371), .A(n4439), .B(n4370), .ZN(n4373)
         );
  OAI211_X1 U4927 ( .C1(n4442), .C2(n4375), .A(n4374), .B(n4373), .ZN(U3251)
         );
  AOI211_X1 U4928 ( .C1(n4378), .C2(n4377), .A(n4376), .B(n4430), .ZN(n4380)
         );
  AOI211_X1 U4929 ( .C1(n4434), .C2(ADDR_REG_12__SCAN_IN), .A(n4380), .B(n4379), .ZN(n4384) );
  OAI211_X1 U4930 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4382), .A(n4439), .B(n4381), .ZN(n4383) );
  OAI211_X1 U4931 ( .C1(n4442), .C2(n4472), .A(n4384), .B(n4383), .ZN(U3252)
         );
  AOI211_X1 U4932 ( .C1(n2046), .C2(n4386), .A(n4385), .B(n4430), .ZN(n4388)
         );
  AOI211_X1 U4933 ( .C1(n4434), .C2(ADDR_REG_13__SCAN_IN), .A(n4388), .B(n4387), .ZN(n4393) );
  AOI22_X1 U4934 ( .A1(REG2_REG_13__SCAN_IN), .A2(n4470), .B1(n4394), .B2(
        n3360), .ZN(n4391) );
  AOI21_X1 U4935 ( .B1(n4391), .B2(n4390), .A(n4398), .ZN(n4389) );
  OAI21_X1 U4936 ( .B1(n4391), .B2(n4390), .A(n4389), .ZN(n4392) );
  OAI211_X1 U4937 ( .C1(n4442), .C2(n4394), .A(n4393), .B(n4392), .ZN(U3253)
         );
  NAND2_X1 U4938 ( .A1(ADDR_REG_14__SCAN_IN), .A2(n4434), .ZN(n4406) );
  AOI211_X1 U4939 ( .C1(n4397), .C2(n4396), .A(n4395), .B(n4430), .ZN(n4402)
         );
  AOI211_X1 U4940 ( .C1(n3337), .C2(n4400), .A(n4399), .B(n4398), .ZN(n4401)
         );
  AOI211_X1 U4941 ( .C1(n4403), .C2(n4468), .A(n4402), .B(n4401), .ZN(n4405)
         );
  NAND3_X1 U4942 ( .A1(n4406), .A2(n4405), .A3(n4404), .ZN(U3254) );
  AOI211_X1 U4943 ( .C1(n4409), .C2(n4408), .A(n4407), .B(n4430), .ZN(n4410)
         );
  AOI211_X1 U4944 ( .C1(n4434), .C2(ADDR_REG_15__SCAN_IN), .A(n4411), .B(n4410), .ZN(n4416) );
  AOI21_X1 U4945 ( .B1(n4413), .B2(n2045), .A(n4412), .ZN(n4414) );
  NAND2_X1 U4946 ( .A1(n4439), .A2(n4414), .ZN(n4415) );
  OAI211_X1 U4947 ( .C1(n4442), .C2(n4417), .A(n4416), .B(n4415), .ZN(U3255)
         );
  AOI21_X1 U4948 ( .B1(n4434), .B2(ADDR_REG_17__SCAN_IN), .A(n4418), .ZN(n4429) );
  OAI21_X1 U4949 ( .B1(n4421), .B2(n4420), .A(n4419), .ZN(n4426) );
  OAI21_X1 U4950 ( .B1(n4424), .B2(n4423), .A(n4422), .ZN(n4425) );
  AOI22_X1 U4951 ( .A1(n4427), .A2(n4426), .B1(n4439), .B2(n4425), .ZN(n4428)
         );
  OAI211_X1 U4952 ( .C1(n4465), .C2(n4442), .A(n4429), .B(n4428), .ZN(U3257)
         );
  AOI21_X1 U4953 ( .B1(n4437), .B2(n4436), .A(n4435), .ZN(n4438) );
  NAND2_X1 U4954 ( .A1(n4439), .A2(n4438), .ZN(n4440) );
  OAI211_X1 U4955 ( .C1(n4442), .C2(n4463), .A(n4441), .B(n4440), .ZN(U3258)
         );
  AOI22_X1 U4956 ( .A1(REG3_REG_2__SCAN_IN), .A2(n4453), .B1(
        REG2_REG_2__SCAN_IN), .B2(n4458), .ZN(n4448) );
  INV_X1 U4957 ( .A(n4443), .ZN(n4445) );
  AOI22_X1 U4958 ( .A1(n4446), .A2(n4445), .B1(n4455), .B2(n4444), .ZN(n4447)
         );
  OAI211_X1 U4959 ( .C1(n4458), .C2(n4449), .A(n4448), .B(n4447), .ZN(U3288)
         );
  AOI21_X1 U4960 ( .B1(n4452), .B2(n4451), .A(n4450), .ZN(n4457) );
  AOI22_X1 U4961 ( .A1(n4455), .A2(n4454), .B1(REG3_REG_0__SCAN_IN), .B2(n4453), .ZN(n4456) );
  OAI221_X1 U4962 ( .B1(n4458), .B2(n4457), .C1(n4136), .C2(n2335), .A(n4456), 
        .ZN(U3290) );
  AND2_X1 U4963 ( .A1(D_REG_31__SCAN_IN), .A2(n4460), .ZN(U3291) );
  AND2_X1 U4964 ( .A1(D_REG_30__SCAN_IN), .A2(n4460), .ZN(U3292) );
  AND2_X1 U4965 ( .A1(D_REG_29__SCAN_IN), .A2(n4460), .ZN(U3293) );
  AND2_X1 U4966 ( .A1(D_REG_28__SCAN_IN), .A2(n4460), .ZN(U3294) );
  AND2_X1 U4967 ( .A1(D_REG_27__SCAN_IN), .A2(n4460), .ZN(U3295) );
  AND2_X1 U4968 ( .A1(D_REG_26__SCAN_IN), .A2(n4460), .ZN(U3296) );
  AND2_X1 U4969 ( .A1(D_REG_25__SCAN_IN), .A2(n4460), .ZN(U3297) );
  AND2_X1 U4970 ( .A1(D_REG_24__SCAN_IN), .A2(n4460), .ZN(U3298) );
  AND2_X1 U4971 ( .A1(D_REG_23__SCAN_IN), .A2(n4460), .ZN(U3299) );
  AND2_X1 U4972 ( .A1(D_REG_22__SCAN_IN), .A2(n4460), .ZN(U3300) );
  AND2_X1 U4973 ( .A1(D_REG_21__SCAN_IN), .A2(n4460), .ZN(U3301) );
  INV_X1 U4974 ( .A(D_REG_20__SCAN_IN), .ZN(n4626) );
  NOR2_X1 U4975 ( .A1(n4459), .A2(n4626), .ZN(U3302) );
  AND2_X1 U4976 ( .A1(D_REG_19__SCAN_IN), .A2(n4460), .ZN(U3303) );
  AND2_X1 U4977 ( .A1(D_REG_18__SCAN_IN), .A2(n4460), .ZN(U3304) );
  AND2_X1 U4978 ( .A1(D_REG_17__SCAN_IN), .A2(n4460), .ZN(U3305) );
  AND2_X1 U4979 ( .A1(D_REG_16__SCAN_IN), .A2(n4460), .ZN(U3306) );
  AND2_X1 U4980 ( .A1(D_REG_15__SCAN_IN), .A2(n4460), .ZN(U3307) );
  AND2_X1 U4981 ( .A1(D_REG_14__SCAN_IN), .A2(n4460), .ZN(U3308) );
  INV_X1 U4982 ( .A(D_REG_13__SCAN_IN), .ZN(n4627) );
  NOR2_X1 U4983 ( .A1(n4459), .A2(n4627), .ZN(U3309) );
  AND2_X1 U4984 ( .A1(D_REG_12__SCAN_IN), .A2(n4460), .ZN(U3310) );
  AND2_X1 U4985 ( .A1(D_REG_11__SCAN_IN), .A2(n4460), .ZN(U3311) );
  AND2_X1 U4986 ( .A1(D_REG_10__SCAN_IN), .A2(n4460), .ZN(U3312) );
  AND2_X1 U4987 ( .A1(D_REG_9__SCAN_IN), .A2(n4460), .ZN(U3313) );
  INV_X1 U4988 ( .A(D_REG_8__SCAN_IN), .ZN(n4624) );
  NOR2_X1 U4989 ( .A1(n4459), .A2(n4624), .ZN(U3314) );
  AND2_X1 U4990 ( .A1(D_REG_7__SCAN_IN), .A2(n4460), .ZN(U3315) );
  AND2_X1 U4991 ( .A1(D_REG_6__SCAN_IN), .A2(n4460), .ZN(U3316) );
  INV_X1 U4992 ( .A(D_REG_5__SCAN_IN), .ZN(n4623) );
  NOR2_X1 U4993 ( .A1(n4459), .A2(n4623), .ZN(U3317) );
  AND2_X1 U4994 ( .A1(D_REG_4__SCAN_IN), .A2(n4460), .ZN(U3318) );
  INV_X1 U4995 ( .A(D_REG_3__SCAN_IN), .ZN(n4613) );
  NOR2_X1 U4996 ( .A1(n4459), .A2(n4613), .ZN(U3319) );
  AND2_X1 U4997 ( .A1(D_REG_2__SCAN_IN), .A2(n4460), .ZN(U3320) );
  INV_X1 U4998 ( .A(DATAI_23_), .ZN(n4462) );
  AOI21_X1 U4999 ( .B1(U3149), .B2(n4462), .A(n4461), .ZN(U3329) );
  INV_X1 U5000 ( .A(DATAI_18_), .ZN(n4592) );
  AOI22_X1 U5001 ( .A1(STATE_REG_SCAN_IN), .A2(n4463), .B1(n4592), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U5002 ( .A1(STATE_REG_SCAN_IN), .A2(n4465), .B1(n4464), .B2(U3149), 
        .ZN(U3335) );
  OAI22_X1 U5003 ( .A1(U3149), .A2(n4466), .B1(DATAI_15_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4467) );
  INV_X1 U5004 ( .A(n4467), .ZN(U3337) );
  OAI22_X1 U5005 ( .A1(U3149), .A2(n4468), .B1(DATAI_14_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4469) );
  INV_X1 U5006 ( .A(n4469), .ZN(U3338) );
  OAI22_X1 U5007 ( .A1(U3149), .A2(n4470), .B1(DATAI_13_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4471) );
  INV_X1 U5008 ( .A(n4471), .ZN(U3339) );
  AOI22_X1 U5009 ( .A1(STATE_REG_SCAN_IN), .A2(n4472), .B1(n2487), .B2(U3149), 
        .ZN(U3340) );
  OAI22_X1 U5010 ( .A1(U3149), .A2(n4473), .B1(DATAI_11_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4474) );
  INV_X1 U5011 ( .A(n4474), .ZN(U3341) );
  OAI22_X1 U5012 ( .A1(U3149), .A2(n4475), .B1(DATAI_10_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4476) );
  INV_X1 U5013 ( .A(n4476), .ZN(U3342) );
  AOI22_X1 U5014 ( .A1(STATE_REG_SCAN_IN), .A2(n4477), .B1(n4595), .B2(U3149), 
        .ZN(U3343) );
  AOI22_X1 U5015 ( .A1(STATE_REG_SCAN_IN), .A2(n2795), .B1(n2341), .B2(U3149), 
        .ZN(U3352) );
  AOI22_X1 U5016 ( .A1(n4516), .A2(n4478), .B1(n2336), .B2(n4514), .ZN(U3467)
         );
  OAI22_X1 U5017 ( .A1(n4480), .A2(n4484), .B1(n4510), .B2(n4479), .ZN(n4481)
         );
  NOR2_X1 U5018 ( .A1(n4482), .A2(n4481), .ZN(n4517) );
  INV_X1 U5019 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4483) );
  AOI22_X1 U5020 ( .A1(n4516), .A2(n4517), .B1(n4483), .B2(n4514), .ZN(U3469)
         );
  NOR2_X1 U5021 ( .A1(n4485), .A2(n4484), .ZN(n4487) );
  AOI211_X1 U5022 ( .C1(n4489), .C2(n4488), .A(n4487), .B(n4486), .ZN(n4518)
         );
  INV_X1 U5023 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4490) );
  AOI22_X1 U5024 ( .A1(n4516), .A2(n4518), .B1(n4490), .B2(n4514), .ZN(U3473)
         );
  INV_X1 U5025 ( .A(n4491), .ZN(n4496) );
  INV_X1 U5026 ( .A(n4492), .ZN(n4494) );
  AOI211_X1 U5027 ( .C1(n4496), .C2(n4495), .A(n4494), .B(n4493), .ZN(n4519)
         );
  AOI22_X1 U5028 ( .A1(n4516), .A2(n4519), .B1(n2368), .B2(n4514), .ZN(U3475)
         );
  OAI21_X1 U5029 ( .B1(n4510), .B2(n4498), .A(n4497), .ZN(n4499) );
  AOI21_X1 U5030 ( .B1(n4500), .B2(n4512), .A(n4499), .ZN(n4520) );
  AOI22_X1 U5031 ( .A1(n4516), .A2(n4520), .B1(n2382), .B2(n4514), .ZN(U3477)
         );
  NOR2_X1 U5032 ( .A1(n4502), .A2(n4501), .ZN(n4506) );
  AOI211_X1 U5033 ( .C1(n4506), .C2(n4505), .A(n4504), .B(n4503), .ZN(n4521)
         );
  INV_X1 U5034 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4507) );
  AOI22_X1 U5035 ( .A1(n4516), .A2(n4521), .B1(n4507), .B2(n4514), .ZN(U3481)
         );
  OAI21_X1 U5036 ( .B1(n4510), .B2(n4509), .A(n4508), .ZN(n4511) );
  AOI21_X1 U5037 ( .B1(n4513), .B2(n4512), .A(n4511), .ZN(n4523) );
  INV_X1 U5038 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4515) );
  AOI22_X1 U5039 ( .A1(n4516), .A2(n4523), .B1(n4515), .B2(n4514), .ZN(U3485)
         );
  AOI22_X1 U5040 ( .A1(n4524), .A2(n4517), .B1(n2716), .B2(n4522), .ZN(U3519)
         );
  AOI22_X1 U5041 ( .A1(n4524), .A2(n4518), .B1(n2353), .B2(n4522), .ZN(U3521)
         );
  AOI22_X1 U5042 ( .A1(n4524), .A2(n4519), .B1(n2738), .B2(n4522), .ZN(U3522)
         );
  AOI22_X1 U5043 ( .A1(n4524), .A2(n4520), .B1(n2741), .B2(n4522), .ZN(U3523)
         );
  AOI22_X1 U5044 ( .A1(n4524), .A2(n4521), .B1(n2770), .B2(n4522), .ZN(U3525)
         );
  AOI22_X1 U5045 ( .A1(n4524), .A2(n4523), .B1(n2432), .B2(n4522), .ZN(U3527)
         );
  AOI22_X1 U5046 ( .A1(n4527), .A2(keyinput24), .B1(keyinput5), .B2(n4526), 
        .ZN(n4525) );
  OAI221_X1 U5047 ( .B1(n4527), .B2(keyinput24), .C1(n4526), .C2(keyinput5), 
        .A(n4525), .ZN(n4539) );
  AOI22_X1 U5048 ( .A1(n4530), .A2(keyinput8), .B1(n4529), .B2(keyinput12), 
        .ZN(n4528) );
  OAI221_X1 U5049 ( .B1(n4530), .B2(keyinput8), .C1(n4529), .C2(keyinput12), 
        .A(n4528), .ZN(n4538) );
  AOI22_X1 U5050 ( .A1(n4533), .A2(keyinput60), .B1(keyinput44), .B2(n4532), 
        .ZN(n4531) );
  OAI221_X1 U5051 ( .B1(n4533), .B2(keyinput60), .C1(n4532), .C2(keyinput44), 
        .A(n4531), .ZN(n4537) );
  AOI22_X1 U5052 ( .A1(n2738), .A2(keyinput37), .B1(n4535), .B2(keyinput19), 
        .ZN(n4534) );
  OAI221_X1 U5053 ( .B1(n2738), .B2(keyinput37), .C1(n4535), .C2(keyinput19), 
        .A(n4534), .ZN(n4536) );
  NOR4_X1 U5054 ( .A1(n4539), .A2(n4538), .A3(n4537), .A4(n4536), .ZN(n4583)
         );
  AOI22_X1 U5055 ( .A1(n3180), .A2(keyinput31), .B1(n2401), .B2(keyinput50), 
        .ZN(n4540) );
  OAI221_X1 U5056 ( .B1(n3180), .B2(keyinput31), .C1(n2401), .C2(keyinput50), 
        .A(n4540), .ZN(n4552) );
  AOI22_X1 U5057 ( .A1(n4543), .A2(keyinput53), .B1(n4542), .B2(keyinput43), 
        .ZN(n4541) );
  OAI221_X1 U5058 ( .B1(n4543), .B2(keyinput53), .C1(n4542), .C2(keyinput43), 
        .A(n4541), .ZN(n4551) );
  AOI22_X1 U5059 ( .A1(n4546), .A2(keyinput41), .B1(n4545), .B2(keyinput33), 
        .ZN(n4544) );
  OAI221_X1 U5060 ( .B1(n4546), .B2(keyinput41), .C1(n4545), .C2(keyinput33), 
        .A(n4544), .ZN(n4550) );
  XNOR2_X1 U5061 ( .A(REG2_REG_1__SCAN_IN), .B(keyinput21), .ZN(n4548) );
  XNOR2_X1 U5062 ( .A(REG1_REG_28__SCAN_IN), .B(keyinput1), .ZN(n4547) );
  NAND2_X1 U5063 ( .A1(n4548), .A2(n4547), .ZN(n4549) );
  NOR4_X1 U5064 ( .A1(n4552), .A2(n4551), .A3(n4550), .A4(n4549), .ZN(n4582)
         );
  AOI22_X1 U5065 ( .A1(n3929), .A2(keyinput57), .B1(n3237), .B2(keyinput46), 
        .ZN(n4553) );
  OAI221_X1 U5066 ( .B1(n3929), .B2(keyinput57), .C1(n3237), .C2(keyinput46), 
        .A(n4553), .ZN(n4564) );
  AOI22_X1 U5067 ( .A1(n4185), .A2(keyinput2), .B1(n4099), .B2(keyinput6), 
        .ZN(n4554) );
  OAI221_X1 U5068 ( .B1(n4185), .B2(keyinput2), .C1(n4099), .C2(keyinput6), 
        .A(n4554), .ZN(n4563) );
  INV_X1 U5069 ( .A(ADDR_REG_8__SCAN_IN), .ZN(n4557) );
  INV_X1 U5070 ( .A(ADDR_REG_13__SCAN_IN), .ZN(n4556) );
  AOI22_X1 U5071 ( .A1(n4557), .A2(keyinput0), .B1(n4556), .B2(keyinput35), 
        .ZN(n4555) );
  OAI221_X1 U5072 ( .B1(n4557), .B2(keyinput0), .C1(n4556), .C2(keyinput35), 
        .A(n4555), .ZN(n4562) );
  INV_X1 U5073 ( .A(ADDR_REG_7__SCAN_IN), .ZN(n4559) );
  AOI22_X1 U5074 ( .A1(n4560), .A2(keyinput18), .B1(keyinput14), .B2(n4559), 
        .ZN(n4558) );
  OAI221_X1 U5075 ( .B1(n4560), .B2(keyinput18), .C1(n4559), .C2(keyinput14), 
        .A(n4558), .ZN(n4561) );
  NOR4_X1 U5076 ( .A1(n4564), .A2(n4563), .A3(n4562), .A4(n4561), .ZN(n4581)
         );
  AOI22_X1 U5077 ( .A1(n4567), .A2(keyinput4), .B1(keyinput39), .B2(n4566), 
        .ZN(n4565) );
  OAI221_X1 U5078 ( .B1(n4567), .B2(keyinput4), .C1(n4566), .C2(keyinput39), 
        .A(n4565), .ZN(n4579) );
  AOI22_X1 U5079 ( .A1(n4570), .A2(keyinput42), .B1(n4569), .B2(keyinput61), 
        .ZN(n4568) );
  OAI221_X1 U5080 ( .B1(n4570), .B2(keyinput42), .C1(n4569), .C2(keyinput61), 
        .A(n4568), .ZN(n4578) );
  AOI22_X1 U5081 ( .A1(n4573), .A2(keyinput32), .B1(keyinput49), .B2(n4572), 
        .ZN(n4571) );
  OAI221_X1 U5082 ( .B1(n4573), .B2(keyinput32), .C1(n4572), .C2(keyinput49), 
        .A(n4571), .ZN(n4577) );
  AOI22_X1 U5083 ( .A1(n4575), .A2(keyinput7), .B1(keyinput58), .B2(n2397), 
        .ZN(n4574) );
  OAI221_X1 U5084 ( .B1(n4575), .B2(keyinput7), .C1(n2397), .C2(keyinput58), 
        .A(n4574), .ZN(n4576) );
  NOR4_X1 U5085 ( .A1(n4579), .A2(n4578), .A3(n4577), .A4(n4576), .ZN(n4580)
         );
  NAND4_X1 U5086 ( .A1(n4583), .A2(n4582), .A3(n4581), .A4(n4580), .ZN(n4639)
         );
  INV_X1 U5087 ( .A(DATAI_30_), .ZN(n4586) );
  INV_X1 U5088 ( .A(DATAI_26_), .ZN(n4585) );
  AOI22_X1 U5089 ( .A1(n4586), .A2(keyinput28), .B1(n4585), .B2(keyinput23), 
        .ZN(n4584) );
  OAI221_X1 U5090 ( .B1(n4586), .B2(keyinput28), .C1(n4585), .C2(keyinput23), 
        .A(n4584), .ZN(n4599) );
  INV_X1 U5091 ( .A(DATAI_24_), .ZN(n4588) );
  AOI22_X1 U5092 ( .A1(n4589), .A2(keyinput30), .B1(keyinput40), .B2(n4588), 
        .ZN(n4587) );
  OAI221_X1 U5093 ( .B1(n4589), .B2(keyinput30), .C1(n4588), .C2(keyinput40), 
        .A(n4587), .ZN(n4598) );
  AOI22_X1 U5094 ( .A1(n4592), .A2(keyinput54), .B1(n4591), .B2(keyinput3), 
        .ZN(n4590) );
  OAI221_X1 U5095 ( .B1(n4592), .B2(keyinput54), .C1(n4591), .C2(keyinput3), 
        .A(n4590), .ZN(n4597) );
  AOI22_X1 U5096 ( .A1(n4595), .A2(keyinput17), .B1(keyinput45), .B2(n4594), 
        .ZN(n4593) );
  OAI221_X1 U5097 ( .B1(n4595), .B2(keyinput17), .C1(n4594), .C2(keyinput45), 
        .A(n4593), .ZN(n4596) );
  NOR4_X1 U5098 ( .A1(n4599), .A2(n4598), .A3(n4597), .A4(n4596), .ZN(n4637)
         );
  AOI22_X1 U5099 ( .A1(n4602), .A2(keyinput48), .B1(keyinput29), .B2(n4601), 
        .ZN(n4600) );
  OAI221_X1 U5100 ( .B1(n4602), .B2(keyinput48), .C1(n4601), .C2(keyinput29), 
        .A(n4600), .ZN(n4610) );
  XNOR2_X1 U5101 ( .A(REG3_REG_17__SCAN_IN), .B(keyinput34), .ZN(n4606) );
  XNOR2_X1 U5102 ( .A(DATAI_3_), .B(keyinput62), .ZN(n4605) );
  XNOR2_X1 U5103 ( .A(IR_REG_10__SCAN_IN), .B(keyinput16), .ZN(n4604) );
  XNOR2_X1 U5104 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput59), .ZN(n4603) );
  NAND4_X1 U5105 ( .A1(n4606), .A2(n4605), .A3(n4604), .A4(n4603), .ZN(n4609)
         );
  XNOR2_X1 U5106 ( .A(keyinput51), .B(n2341), .ZN(n4608) );
  XNOR2_X1 U5107 ( .A(keyinput25), .B(n2483), .ZN(n4607) );
  NOR4_X1 U5108 ( .A1(n4610), .A2(n4609), .A3(n4608), .A4(n4607), .ZN(n4636)
         );
  AOI22_X1 U5109 ( .A1(n4613), .A2(keyinput15), .B1(n4612), .B2(keyinput26), 
        .ZN(n4611) );
  OAI221_X1 U5110 ( .B1(n4613), .B2(keyinput15), .C1(n4612), .C2(keyinput26), 
        .A(n4611), .ZN(n4621) );
  XNOR2_X1 U5111 ( .A(keyinput20), .B(n2279), .ZN(n4620) );
  XNOR2_X1 U5112 ( .A(keyinput47), .B(n2607), .ZN(n4619) );
  XNOR2_X1 U5113 ( .A(IR_REG_15__SCAN_IN), .B(keyinput38), .ZN(n4617) );
  XNOR2_X1 U5114 ( .A(IR_REG_13__SCAN_IN), .B(keyinput63), .ZN(n4616) );
  XNOR2_X1 U5115 ( .A(IR_REG_25__SCAN_IN), .B(keyinput13), .ZN(n4615) );
  XNOR2_X1 U5116 ( .A(IR_REG_18__SCAN_IN), .B(keyinput27), .ZN(n4614) );
  NAND4_X1 U5117 ( .A1(n4617), .A2(n4616), .A3(n4615), .A4(n4614), .ZN(n4618)
         );
  NOR4_X1 U5118 ( .A1(n4621), .A2(n4620), .A3(n4619), .A4(n4618), .ZN(n4635)
         );
  AOI22_X1 U5119 ( .A1(n4624), .A2(keyinput10), .B1(n4623), .B2(keyinput11), 
        .ZN(n4622) );
  OAI221_X1 U5120 ( .B1(n4624), .B2(keyinput10), .C1(n4623), .C2(keyinput11), 
        .A(n4622), .ZN(n4633) );
  AOI22_X1 U5121 ( .A1(n4627), .A2(keyinput9), .B1(keyinput22), .B2(n4626), 
        .ZN(n4625) );
  OAI221_X1 U5122 ( .B1(n4627), .B2(keyinput9), .C1(n4626), .C2(keyinput22), 
        .A(n4625), .ZN(n4632) );
  AOI22_X1 U5123 ( .A1(n2336), .A2(keyinput52), .B1(keyinput56), .B2(n2368), 
        .ZN(n4628) );
  OAI221_X1 U5124 ( .B1(n2336), .B2(keyinput52), .C1(n2368), .C2(keyinput56), 
        .A(n4628), .ZN(n4631) );
  AOI22_X1 U5125 ( .A1(n2382), .A2(keyinput55), .B1(n2396), .B2(keyinput36), 
        .ZN(n4629) );
  OAI221_X1 U5126 ( .B1(n2382), .B2(keyinput55), .C1(n2396), .C2(keyinput36), 
        .A(n4629), .ZN(n4630) );
  NOR4_X1 U5127 ( .A1(n4633), .A2(n4632), .A3(n4631), .A4(n4630), .ZN(n4634)
         );
  NAND4_X1 U5128 ( .A1(n4637), .A2(n4636), .A3(n4635), .A4(n4634), .ZN(n4638)
         );
  NOR2_X1 U5129 ( .A1(n4639), .A2(n4638), .ZN(n4667) );
  NOR4_X1 U5130 ( .A1(REG2_REG_10__SCAN_IN), .A2(REG2_REG_1__SCAN_IN), .A3(
        REG0_REG_0__SCAN_IN), .A4(ADDR_REG_8__SCAN_IN), .ZN(n4665) );
  NAND3_X1 U5131 ( .A1(ADDR_REG_13__SCAN_IN), .A2(DATAO_REG_26__SCAN_IN), .A3(
        n2401), .ZN(n4642) );
  NAND4_X1 U5132 ( .A1(DATAI_26_), .A2(DATAO_REG_22__SCAN_IN), .A3(
        DATAO_REG_30__SCAN_IN), .A4(DATAO_REG_5__SCAN_IN), .ZN(n4641) );
  NAND4_X1 U5133 ( .A1(REG1_REG_27__SCAN_IN), .A2(DATAI_16_), .A3(DATAI_0_), 
        .A4(REG0_REG_30__SCAN_IN), .ZN(n4640) );
  NOR4_X1 U5134 ( .A1(ADDR_REG_7__SCAN_IN), .A2(n4642), .A3(n4641), .A4(n4640), 
        .ZN(n4664) );
  NAND4_X1 U5135 ( .A1(D_REG_20__SCAN_IN), .A2(D_REG_8__SCAN_IN), .A3(
        D_REG_3__SCAN_IN), .A4(REG0_REG_26__SCAN_IN), .ZN(n4646) );
  NAND4_X1 U5136 ( .A1(REG1_REG_13__SCAN_IN), .A2(REG0_REG_6__SCAN_IN), .A3(
        REG0_REG_4__SCAN_IN), .A4(ADDR_REG_4__SCAN_IN), .ZN(n4645) );
  NAND4_X1 U5137 ( .A1(REG2_REG_8__SCAN_IN), .A2(REG2_REG_3__SCAN_IN), .A3(
        REG1_REG_4__SCAN_IN), .A4(DATAI_30_), .ZN(n4644) );
  NAND4_X1 U5138 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG2_REG_22__SCAN_IN), .A3(
        REG1_REG_19__SCAN_IN), .A4(REG2_REG_18__SCAN_IN), .ZN(n4643) );
  NOR4_X1 U5139 ( .A1(n4646), .A2(n4645), .A3(n4644), .A4(n4643), .ZN(n4663)
         );
  NOR4_X1 U5140 ( .A1(DATAI_25_), .A2(DATAI_24_), .A3(DATAO_REG_27__SCAN_IN), 
        .A4(DATAO_REG_1__SCAN_IN), .ZN(n4650) );
  NOR4_X1 U5141 ( .A1(D_REG_1__SCAN_IN), .A2(DATAI_7_), .A3(DATAI_18_), .A4(
        REG0_REG_31__SCAN_IN), .ZN(n4649) );
  NOR4_X1 U5142 ( .A1(REG1_REG_28__SCAN_IN), .A2(REG1_REG_26__SCAN_IN), .A3(
        REG0_REG_25__SCAN_IN), .A4(REG0_REG_24__SCAN_IN), .ZN(n4648) );
  NOR4_X1 U5143 ( .A1(DATAI_9_), .A2(REG0_REG_5__SCAN_IN), .A3(DATAI_3_), .A4(
        REG0_REG_18__SCAN_IN), .ZN(n4647) );
  NAND4_X1 U5144 ( .A1(n4650), .A2(n4649), .A3(n4648), .A4(n4647), .ZN(n4661)
         );
  INV_X1 U5145 ( .A(n4651), .ZN(n4660) );
  INV_X1 U5146 ( .A(REG3_REG_4__SCAN_IN), .ZN(n4652) );
  NAND4_X1 U5147 ( .A1(n4653), .A2(REG3_REG_10__SCAN_IN), .A3(
        REG1_REG_21__SCAN_IN), .A4(n4652), .ZN(n4659) );
  NAND4_X1 U5148 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .A3(
        REG3_REG_18__SCAN_IN), .A4(REG3_REG_17__SCAN_IN), .ZN(n4657) );
  NAND3_X1 U5149 ( .A1(n4654), .A2(n2279), .A3(n2397), .ZN(n4656) );
  OR4_X1 U5150 ( .A1(n4657), .A2(n4656), .A3(IR_REG_13__SCAN_IN), .A4(n4655), 
        .ZN(n4658) );
  NOR4_X1 U5151 ( .A1(n4661), .A2(n4660), .A3(n4659), .A4(n4658), .ZN(n4662)
         );
  NAND4_X1 U5152 ( .A1(n4665), .A2(n4664), .A3(n4663), .A4(n4662), .ZN(n4666)
         );
  XNOR2_X1 U5153 ( .A(n4667), .B(n4666), .ZN(n4670) );
  NAND2_X1 U5154 ( .A1(n2186), .A2(U4043), .ZN(n4668) );
  OAI21_X1 U5155 ( .B1(U4043), .B2(DATAO_REG_21__SCAN_IN), .A(n4668), .ZN(
        n4669) );
  XNOR2_X1 U5156 ( .A(n4670), .B(n4669), .ZN(U3571) );
  CLKBUF_X1 U2258 ( .A(n2787), .Z(n2931) );
endmodule

