

module b17_C_AntiSAT_k_256_5 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, 
        keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, 
        keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, 
        keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, 
        keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, 
        keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, 
        keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, 
        keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, 
        keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, 
        keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, 
        keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, 
        keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, 
        keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, 
        keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, 
        keyinput196, keyinput197, keyinput198, keyinput199, keyinput200, 
        keyinput201, keyinput202, keyinput203, keyinput204, keyinput205, 
        keyinput206, keyinput207, keyinput208, keyinput209, keyinput210, 
        keyinput211, keyinput212, keyinput213, keyinput214, keyinput215, 
        keyinput216, keyinput217, keyinput218, keyinput219, keyinput220, 
        keyinput221, keyinput222, keyinput223, keyinput224, keyinput225, 
        keyinput226, keyinput227, keyinput228, keyinput229, keyinput230, 
        keyinput231, keyinput232, keyinput233, keyinput234, keyinput235, 
        keyinput236, keyinput237, keyinput238, keyinput239, keyinput240, 
        keyinput241, keyinput242, keyinput243, keyinput244, keyinput245, 
        keyinput246, keyinput247, keyinput248, keyinput249, keyinput250, 
        keyinput251, keyinput252, keyinput253, keyinput254, keyinput255, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9822, n9823, n9824, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,
         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
         n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
         n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626,
         n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
         n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
         n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650,
         n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
         n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666,
         n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674,
         n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
         n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
         n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,
         n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706,
         n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
         n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722,
         n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,
         n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738,
         n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746,
         n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,
         n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762,
         n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770,
         n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778,
         n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786,
         n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794,
         n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802,
         n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810,
         n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818,
         n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826,
         n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834,
         n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842,
         n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850,
         n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858,
         n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866,
         n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874,
         n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882,
         n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890,
         n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898,
         n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906,
         n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914,
         n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922,
         n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930,
         n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938,
         n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946,
         n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954,
         n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962,
         n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970,
         n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978,
         n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986,
         n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994,
         n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002,
         n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010,
         n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,
         n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026,
         n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034,
         n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042,
         n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050,
         n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058,
         n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066,
         n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,
         n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082,
         n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090,
         n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098,
         n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106,
         n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114,
         n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122,
         n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130,
         n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,
         n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146,
         n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154,
         n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162,
         n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170,
         n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178,
         n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186,
         n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194,
         n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202,
         n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210,
         n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218,
         n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226,
         n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,
         n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242,
         n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250,
         n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258,
         n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266,
         n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274,
         n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282,
         n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290,
         n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298,
         n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
         n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314,
         n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322,
         n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330,
         n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,
         n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346,
         n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354,
         n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362,
         n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370,
         n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
         n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386,
         n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394,
         n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402,
         n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,
         n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418,
         n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426,
         n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434,
         n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442,
         n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
         n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458,
         n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466,
         n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474,
         n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
         n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490,
         n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
         n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
         n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
         n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
         n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
         n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538,
         n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546,
         n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,
         n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562,
         n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570,
         n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,
         n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586,
         n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
         n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602,
         n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610,
         n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618,
         n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626,
         n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634,
         n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642,
         n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650,
         n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658,
         n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,
         n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674,
         n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682,
         n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690,
         n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,
         n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706,
         n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714,
         n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722,
         n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730,
         n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738,
         n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746,
         n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754,
         n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762,
         n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770,
         n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778,
         n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786,
         n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794,
         n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802,
         n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810,
         n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818,
         n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826,
         n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834,
         n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842,
         n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850,
         n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858,
         n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866,
         n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874,
         n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882,
         n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890,
         n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898,
         n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906,
         n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914,
         n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922,
         n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930,
         n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938,
         n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946,
         n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954,
         n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962,
         n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970,
         n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978,
         n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986,
         n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994,
         n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002,
         n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010,
         n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018,
         n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
         n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034,
         n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042,
         n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050,
         n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058,
         n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,
         n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074,
         n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082,
         n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090,
         n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
         n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106,
         n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114,
         n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122,
         n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130,
         n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138,
         n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146,
         n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
         n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
         n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
         n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178,
         n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186,
         n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194,
         n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202,
         n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210,
         n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218,
         n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
         n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234,
         n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,
         n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250,
         n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258,
         n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266,
         n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,
         n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282,
         n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290,
         n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
         n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306,
         n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314,
         n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322,
         n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330,
         n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338,
         n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346,
         n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354,
         n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362,
         n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370,
         n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378,
         n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386,
         n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394,
         n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402,
         n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410,
         n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418,
         n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426,
         n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434,
         n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442,
         n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450,
         n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458,
         n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466,
         n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474,
         n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482,
         n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490,
         n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498,
         n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506,
         n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514,
         n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522,
         n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530,
         n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538,
         n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546,
         n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554,
         n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562,
         n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570,
         n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578,
         n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586,
         n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594,
         n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602,
         n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610,
         n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618,
         n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626,
         n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634,
         n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642,
         n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650,
         n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658,
         n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666,
         n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674,
         n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682,
         n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690,
         n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698,
         n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706,
         n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714,
         n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722,
         n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730,
         n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738,
         n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746,
         n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754,
         n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762,
         n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770,
         n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778,
         n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786,
         n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794,
         n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802,
         n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810,
         n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818,
         n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826,
         n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834,
         n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842,
         n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850,
         n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858,
         n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866,
         n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874,
         n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882,
         n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890,
         n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898,
         n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906,
         n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914,
         n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922,
         n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930,
         n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938,
         n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946,
         n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954,
         n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962,
         n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970,
         n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978,
         n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986,
         n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994,
         n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002,
         n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010,
         n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018,
         n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026,
         n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034,
         n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042,
         n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050,
         n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058,
         n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066,
         n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074,
         n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082,
         n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090,
         n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098,
         n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106,
         n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114,
         n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122,
         n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130,
         n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138,
         n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146,
         n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154,
         n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162,
         n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170,
         n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178,
         n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186,
         n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194,
         n19195, n19197, n19198, n19199, n19200, n19201, n19202, n19203,
         n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211,
         n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219,
         n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227,
         n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235,
         n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
         n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251,
         n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
         n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267,
         n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275,
         n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283,
         n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291,
         n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299,
         n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307,
         n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
         n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323,
         n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331,
         n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339,
         n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347,
         n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355,
         n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363,
         n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371,
         n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
         n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
         n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395,
         n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403,
         n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411,
         n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419,
         n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427,
         n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
         n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443,
         n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451,
         n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459,
         n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467,
         n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475,
         n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483,
         n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491,
         n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499,
         n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507,
         n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515,
         n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523,
         n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531,
         n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539,
         n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547,
         n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555,
         n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563,
         n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571,
         n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579,
         n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587,
         n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595,
         n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603,
         n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611,
         n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619,
         n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627,
         n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635,
         n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643,
         n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651,
         n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659,
         n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667,
         n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675,
         n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683,
         n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691,
         n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699,
         n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707,
         n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715,
         n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
         n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731,
         n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739,
         n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747,
         n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755,
         n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763,
         n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771,
         n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779,
         n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787,
         n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
         n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803,
         n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811,
         n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819,
         n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827,
         n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835,
         n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843,
         n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851,
         n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859,
         n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867,
         n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875,
         n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883,
         n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891,
         n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899,
         n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907,
         n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915,
         n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923,
         n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931,
         n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939,
         n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947,
         n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955,
         n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963,
         n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971,
         n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979,
         n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987,
         n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995,
         n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003,
         n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011,
         n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019,
         n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027,
         n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035,
         n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043,
         n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051,
         n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059,
         n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067,
         n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075,
         n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083,
         n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091,
         n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099,
         n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107,
         n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115,
         n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123,
         n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131,
         n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139,
         n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147,
         n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155,
         n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163,
         n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171,
         n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179,
         n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187,
         n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195,
         n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203,
         n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211,
         n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219,
         n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227,
         n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235,
         n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243,
         n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251,
         n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259,
         n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267,
         n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275,
         n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283,
         n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291,
         n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299,
         n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307,
         n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315,
         n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323,
         n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331,
         n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339,
         n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347,
         n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355,
         n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363,
         n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371,
         n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379,
         n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387,
         n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395,
         n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403,
         n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411,
         n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419,
         n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427,
         n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435,
         n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443,
         n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451,
         n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459,
         n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467,
         n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475,
         n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483,
         n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491,
         n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499,
         n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507,
         n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515,
         n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523,
         n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531,
         n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539,
         n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547,
         n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555,
         n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563,
         n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571,
         n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579,
         n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587,
         n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595,
         n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603,
         n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611,
         n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619,
         n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627,
         n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635,
         n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643,
         n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651,
         n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659,
         n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667,
         n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675,
         n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683,
         n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691,
         n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699,
         n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707,
         n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715,
         n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723,
         n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731,
         n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739,
         n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747,
         n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755,
         n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763,
         n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771,
         n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779,
         n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787,
         n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795,
         n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803,
         n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811,
         n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819,
         n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827,
         n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835,
         n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843,
         n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851,
         n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859,
         n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867,
         n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875,
         n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883,
         n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891,
         n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899,
         n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907,
         n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915,
         n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923,
         n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931,
         n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939,
         n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947,
         n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955,
         n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963,
         n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971,
         n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979,
         n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987,
         n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995,
         n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003,
         n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011,
         n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019,
         n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027,
         n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035,
         n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043,
         n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051,
         n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059,
         n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067,
         n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075,
         n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083,
         n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091,
         n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099,
         n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107,
         n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115,
         n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123,
         n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131,
         n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139,
         n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147,
         n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155,
         n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163,
         n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171,
         n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179,
         n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187,
         n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195,
         n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203,
         n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211,
         n21212, n21213, n21214, n21215, n21216, n21217;

  INV_X1 U11266 ( .A(n19971), .ZN(n19959) );
  INV_X2 U11267 ( .A(n13225), .ZN(n15895) );
  INV_X1 U11268 ( .A(n13570), .ZN(n14441) );
  NOR2_X1 U11269 ( .A1(n11661), .A2(n11660), .ZN(n18167) );
  OR2_X1 U11270 ( .A1(n10522), .A2(n10502), .ZN(n10528) );
  CLKBUF_X2 U11271 ( .A(n12595), .Z(n12871) );
  CLKBUF_X1 U11272 ( .A(n12853), .Z(n13049) );
  CLKBUF_X3 U11273 ( .A(n11545), .Z(n9832) );
  AND2_X1 U11274 ( .A1(n14169), .A2(n12095), .ZN(n12085) );
  CLKBUF_X1 U11275 ( .A(n12225), .Z(n14542) );
  INV_X1 U11276 ( .A(n11684), .ZN(n17139) );
  CLKBUF_X3 U11277 ( .A(n11672), .Z(n9831) );
  INV_X2 U11278 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18762) );
  AND2_X1 U11279 ( .A1(n12271), .A2(n12273), .ZN(n12424) );
  AND2_X1 U11280 ( .A1(n12272), .A2(n12265), .ZN(n12594) );
  INV_X1 U11281 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19859) );
  INV_X1 U11282 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10190) );
  INV_X1 U11283 ( .A(n19180), .ZN(n11197) );
  OR2_X1 U11284 ( .A1(n19158), .A2(n19157), .ZN(n19202) );
  INV_X1 U11285 ( .A(n19202), .ZN(n9822) );
  INV_X1 U11286 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10108) );
  AND2_X2 U11287 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13743) );
  NAND2_X1 U11288 ( .A1(n12542), .A2(n12541), .ZN(n13079) );
  CLKBUF_X3 U11289 ( .A(n10553), .Z(n12093) );
  INV_X1 U11290 ( .A(n12099), .ZN(n10557) );
  AOI22_X1 U11291 ( .A1(n20924), .A2(keyinput168), .B1(n20923), .B2(
        keyinput203), .ZN(n20922) );
  INV_X1 U11292 ( .A(n12402), .ZN(n13141) );
  NAND2_X1 U11293 ( .A1(n11197), .A2(n19174), .ZN(n10465) );
  INV_X1 U11294 ( .A(n19174), .ZN(n11161) );
  NOR2_X1 U11295 ( .A1(n11749), .A2(n15671), .ZN(n18588) );
  NAND4_X1 U11296 ( .A1(n10110), .A2(n12412), .A3(n12509), .A4(n10109), .ZN(
        n12401) );
  AND2_X1 U11297 ( .A1(n14532), .A2(n16293), .ZN(n12064) );
  NOR2_X1 U11298 ( .A1(n10438), .A2(n19169), .ZN(n10445) );
  INV_X1 U11299 ( .A(n11684), .ZN(n9824) );
  INV_X2 U11300 ( .A(n10288), .ZN(n17146) );
  NOR2_X2 U11301 ( .A1(n12401), .A2(n12400), .ZN(n13375) );
  INV_X1 U11302 ( .A(n19945), .ZN(n19934) );
  AND4_X2 U11303 ( .A1(n12363), .A2(n12362), .A3(n12361), .A4(n12360), .ZN(
        n20139) );
  BUF_X1 U11305 ( .A(n10478), .Z(n11117) );
  NOR2_X1 U11306 ( .A1(n19169), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11220) );
  NAND2_X2 U11307 ( .A1(n10438), .A2(n19169), .ZN(n13299) );
  AOI21_X1 U11308 ( .B1(n17614), .B2(n10101), .A(n10091), .ZN(n17609) );
  INV_X1 U11309 ( .A(n17352), .ZN(n18160) );
  AND2_X1 U11310 ( .A1(n14681), .A2(n14682), .ZN(n14680) );
  NAND2_X1 U11311 ( .A1(n11143), .A2(n13299), .ZN(n11199) );
  XNOR2_X1 U11312 ( .A(n10130), .B(n10970), .ZN(n11184) );
  NAND2_X1 U11313 ( .A1(n10000), .A2(n9999), .ZN(n15371) );
  INV_X1 U11314 ( .A(n18878), .ZN(n16261) );
  INV_X1 U11315 ( .A(n17726), .ZN(n17697) );
  INV_X1 U11316 ( .A(n17800), .ZN(n17808) );
  INV_X1 U11317 ( .A(n19928), .ZN(n15867) );
  AND2_X1 U11318 ( .A1(n10522), .A2(n15646), .ZN(n9823) );
  INV_X2 U11319 ( .A(n12078), .ZN(n12050) );
  XNOR2_X2 U11321 ( .A(n13185), .B(n20092), .ZN(n13789) );
  OR2_X4 U11322 ( .A1(n20139), .A2(n20124), .ZN(n13570) );
  AND4_X4 U11323 ( .A1(n12386), .A2(n12385), .A3(n12384), .A4(n12383), .ZN(
        n20124) );
  NAND2_X2 U11325 ( .A1(n13700), .A2(n13178), .ZN(n13185) );
  NOR2_X2 U11326 ( .A1(n13644), .A2(n10222), .ZN(n13696) );
  OAI21_X4 U11327 ( .B1(n13977), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n12437), 
        .ZN(n13170) );
  XNOR2_X2 U11328 ( .A(n13177), .B(n20113), .ZN(n13702) );
  NAND2_X2 U11329 ( .A1(n13633), .A2(n13173), .ZN(n13177) );
  NAND2_X2 U11330 ( .A1(n12470), .A2(n12469), .ZN(n12522) );
  AND3_X4 U11331 ( .A1(n16296), .A2(n10287), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10347) );
  AOI211_X2 U11332 ( .C1(n14854), .C2(n14853), .A(n14852), .B(n14861), .ZN(
        n14855) );
  NOR2_X2 U11333 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11495), .ZN(
        n11630) );
  NAND3_X1 U11334 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(n18769), .ZN(n11495) );
  CLKBUF_X1 U11335 ( .A(n10672), .Z(n9826) );
  BUF_X1 U11336 ( .A(n10672), .Z(n9827) );
  BUF_X2 U11337 ( .A(n18111), .Z(n9828) );
  NAND2_X1 U11338 ( .A1(n14181), .A2(n14180), .ZN(n9976) );
  AOI211_X1 U11340 ( .C1(n16280), .C2(n18997), .A(n11486), .B(n11485), .ZN(
        n11487) );
  NAND2_X1 U11341 ( .A1(n10026), .A2(n15929), .ZN(n14101) );
  OR2_X1 U11342 ( .A1(n10949), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10255) );
  NOR2_X1 U11343 ( .A1(n16077), .A2(n10960), .ZN(n10949) );
  NAND2_X1 U11344 ( .A1(n10200), .A2(n10199), .ZN(n14077) );
  NAND2_X1 U11345 ( .A1(n10648), .A2(n10647), .ZN(n11006) );
  AOI21_X1 U11346 ( .B1(n14913), .B2(n13239), .A(n13238), .ZN(n15891) );
  AND2_X1 U11347 ( .A1(n9971), .A2(n17472), .ZN(n16555) );
  INV_X1 U11348 ( .A(n13865), .ZN(n10200) );
  OR3_X1 U11349 ( .A1(n14669), .A2(n14655), .A3(n10157), .ZN(n14639) );
  NAND2_X1 U11350 ( .A1(n10965), .A2(n16091), .ZN(n16089) );
  OAI21_X1 U11351 ( .B1(n15895), .B2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n13234), .ZN(n14939) );
  NAND3_X1 U11352 ( .A1(n11947), .A2(n9866), .A3(n11948), .ZN(n13680) );
  NAND2_X1 U11353 ( .A1(n12577), .A2(n13776), .ZN(n20122) );
  AND2_X1 U11354 ( .A1(n12514), .A2(n12531), .ZN(n9932) );
  AND2_X1 U11355 ( .A1(n13691), .A2(n10511), .ZN(n19388) );
  NAND2_X1 U11356 ( .A1(n13691), .A2(n10505), .ZN(n10791) );
  NOR2_X1 U11357 ( .A1(n11757), .A2(n18651), .ZN(n11794) );
  INV_X1 U11358 ( .A(n14043), .ZN(n10520) );
  NAND2_X1 U11359 ( .A1(n10493), .A2(n10494), .ZN(n10039) );
  NOR2_X1 U11360 ( .A1(n18163), .A2(n17454), .ZN(n17447) );
  CLKBUF_X3 U11361 ( .A(n16529), .Z(n16853) );
  NAND2_X1 U11362 ( .A1(n13139), .A2(n13123), .ZN(n13604) );
  INV_X2 U11363 ( .A(n13299), .ZN(n19845) );
  INV_X2 U11364 ( .A(n14609), .ZN(n13131) );
  NOR2_X1 U11365 ( .A1(n11576), .A2(n11575), .ZN(n17321) );
  INV_X1 U11366 ( .A(n20124), .ZN(n13620) );
  OR2_X2 U11368 ( .A1(n12293), .A2(n12292), .ZN(n12509) );
  CLKBUF_X2 U11369 ( .A(n20005), .Z(n20819) );
  CLKBUF_X3 U11370 ( .A(n11655), .Z(n9834) );
  BUF_X2 U11371 ( .A(n12424), .Z(n13040) );
  BUF_X2 U11372 ( .A(n12489), .Z(n13039) );
  BUF_X2 U11373 ( .A(n12438), .Z(n13038) );
  CLKBUF_X2 U11374 ( .A(n12496), .Z(n13022) );
  BUF_X2 U11375 ( .A(n12364), .Z(n13047) );
  CLKBUF_X2 U11376 ( .A(n12425), .Z(n13046) );
  BUF_X2 U11377 ( .A(n12594), .Z(n9829) );
  CLKBUF_X2 U11378 ( .A(n12984), .Z(n13048) );
  BUF_X4 U11379 ( .A(n11630), .Z(n9830) );
  NAND2_X4 U11380 ( .A1(n18774), .A2(n18769), .ZN(n16880) );
  INV_X4 U11381 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18769) );
  AND2_X2 U11382 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10549) );
  INV_X2 U11383 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16296) );
  NOR2_X1 U11384 ( .A1(n15408), .A2(n11811), .ZN(n11815) );
  OR2_X1 U11385 ( .A1(n15351), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15446) );
  AND2_X1 U11386 ( .A1(n11877), .A2(n11878), .ZN(n15351) );
  AND2_X1 U11387 ( .A1(n10050), .A2(n9924), .ZN(n15408) );
  AND2_X1 U11388 ( .A1(n11492), .A2(n11491), .ZN(n11493) );
  AND2_X1 U11389 ( .A1(n11158), .A2(n11157), .ZN(n11159) );
  AOI21_X1 U11390 ( .B1(n15553), .B2(n15551), .A(n15549), .ZN(n15535) );
  NAND2_X1 U11391 ( .A1(n9980), .A2(n9910), .ZN(n15553) );
  NOR2_X1 U11392 ( .A1(n15589), .A2(n15695), .ZN(n15571) );
  NAND2_X1 U11393 ( .A1(n10025), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15589) );
  INV_X1 U11394 ( .A(n15423), .ZN(n10025) );
  OAI21_X1 U11395 ( .B1(n14844), .B2(n9922), .A(n10027), .ZN(n9991) );
  AOI211_X1 U11396 ( .C1(n15917), .C2(n14874), .A(n14873), .B(n14872), .ZN(
        n14875) );
  OAI21_X1 U11397 ( .B1(n15188), .B2(n15189), .A(n12201), .ZN(n12217) );
  XNOR2_X1 U11398 ( .A(n9874), .B(n13070), .ZN(n14625) );
  AOI21_X1 U11399 ( .B1(n14637), .B2(n14635), .A(n14636), .ZN(n14848) );
  AND2_X1 U11400 ( .A1(n14870), .A2(n10017), .ZN(n14833) );
  AOI21_X1 U11401 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n14888), .A(
        n14881), .ZN(n14883) );
  OR2_X2 U11402 ( .A1(n14653), .A2(n10127), .ZN(n14635) );
  NOR2_X1 U11403 ( .A1(n12200), .A2(n12199), .ZN(n15181) );
  NAND2_X2 U11404 ( .A1(n14667), .A2(n14668), .ZN(n14653) );
  AND2_X1 U11405 ( .A1(n12177), .A2(n10321), .ZN(n12178) );
  OR2_X1 U11406 ( .A1(n13246), .A2(n15746), .ZN(n10182) );
  NAND2_X1 U11407 ( .A1(n15754), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15753) );
  NOR2_X1 U11408 ( .A1(n14733), .A2(n14734), .ZN(n9844) );
  NOR2_X1 U11409 ( .A1(n10275), .A2(n14186), .ZN(n10018) );
  XNOR2_X1 U11410 ( .A(n11019), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16222) );
  NOR2_X1 U11411 ( .A1(n10277), .A2(n14108), .ZN(n10276) );
  AND2_X1 U11412 ( .A1(n11018), .A2(n10830), .ZN(n11015) );
  XNOR2_X1 U11413 ( .A(n11018), .B(n11020), .ZN(n14214) );
  NAND2_X1 U11414 ( .A1(n14101), .A2(n13229), .ZN(n9990) );
  AOI211_X1 U11415 ( .C1(n19961), .C2(P1_EBX_REG_30__SCAN_IN), .A(n14629), .B(
        n14628), .ZN(n14634) );
  OR2_X1 U11416 ( .A1(n12119), .A2(n12138), .ZN(n10293) );
  OR2_X1 U11417 ( .A1(n15212), .A2(n15211), .ZN(n15214) );
  NAND2_X1 U11418 ( .A1(n9975), .A2(n10828), .ZN(n11018) );
  OR2_X1 U11419 ( .A1(n11009), .A2(n11008), .ZN(n11010) );
  OAI21_X1 U11420 ( .B1(n11011), .B2(n11020), .A(n18949), .ZN(n10785) );
  AND2_X1 U11421 ( .A1(n11011), .A2(n21044), .ZN(n14108) );
  OR2_X1 U11422 ( .A1(n11011), .A2(n21044), .ZN(n14109) );
  XNOR2_X1 U11423 ( .A(n11854), .B(n11480), .ZN(n18997) );
  NAND2_X1 U11424 ( .A1(n10183), .A2(n10186), .ZN(n15932) );
  XNOR2_X1 U11425 ( .A(n11006), .B(n11257), .ZN(n11007) );
  XNOR2_X1 U11426 ( .A(n10778), .B(n9998), .ZN(n11011) );
  AND3_X1 U11427 ( .A1(n10648), .A2(n10647), .A3(n10726), .ZN(n9998) );
  AND2_X1 U11428 ( .A1(n10777), .A2(n10776), .ZN(n10778) );
  NOR2_X1 U11429 ( .A1(n10185), .A2(n10189), .ZN(n10184) );
  AND2_X1 U11430 ( .A1(n13211), .A2(n10187), .ZN(n10186) );
  INV_X1 U11431 ( .A(n10646), .ZN(n10647) );
  NOR2_X1 U11432 ( .A1(n14669), .A2(n14655), .ZN(n14657) );
  NOR2_X1 U11433 ( .A1(n15285), .A2(n15276), .ZN(n15275) );
  OR2_X1 U11434 ( .A1(n14914), .A2(n13243), .ZN(n13244) );
  NAND2_X1 U11435 ( .A1(n14713), .A2(n14670), .ZN(n14669) );
  AND2_X1 U11436 ( .A1(n13208), .A2(n13207), .ZN(n15936) );
  AND2_X1 U11437 ( .A1(n14714), .A2(n14426), .ZN(n14713) );
  INV_X1 U11438 ( .A(n10602), .ZN(n19358) );
  AND2_X1 U11439 ( .A1(n9970), .A2(n9969), .ZN(n16576) );
  OR2_X1 U11440 ( .A1(n13225), .A2(n15970), .ZN(n13234) );
  NAND2_X1 U11441 ( .A1(n13689), .A2(n11942), .ZN(n11948) );
  AOI211_X1 U11442 ( .C1(n10603), .C2(n20990), .A(n19317), .B(n19813), .ZN(
        n19298) );
  XNOR2_X1 U11443 ( .A(n13224), .B(n12636), .ZN(n13212) );
  OR2_X1 U11444 ( .A1(n11946), .A2(n13687), .ZN(n11947) );
  OAI21_X2 U11445 ( .B1(n20122), .B2(n12748), .A(n12565), .ZN(n13721) );
  NAND2_X1 U11446 ( .A1(n12603), .A2(n10192), .ZN(n13224) );
  INV_X1 U11447 ( .A(n10791), .ZN(n19269) );
  NAND2_X1 U11448 ( .A1(n9823), .A2(n10499), .ZN(n19154) );
  AND2_X2 U11449 ( .A1(n13933), .A2(n13931), .ZN(n19945) );
  NAND2_X1 U11450 ( .A1(n9823), .A2(n10500), .ZN(n19240) );
  INV_X1 U11451 ( .A(n19451), .ZN(n19456) );
  NAND2_X1 U11452 ( .A1(n9823), .A2(n10502), .ZN(n10519) );
  NOR2_X1 U11453 ( .A1(n21079), .A2(n17238), .ZN(n17237) );
  NOR2_X1 U11454 ( .A1(n11609), .A2(n17524), .ZN(n17860) );
  OR2_X1 U11455 ( .A1(n10532), .A2(n10527), .ZN(n19580) );
  OR2_X1 U11456 ( .A1(n10528), .A2(n10531), .ZN(n10754) );
  OR2_X1 U11457 ( .A1(n10532), .A2(n10530), .ZN(n19547) );
  OR2_X1 U11458 ( .A1(n10528), .A2(n10526), .ZN(n10752) );
  AND2_X1 U11459 ( .A1(n13575), .A2(n11929), .ZN(n13587) );
  OAI21_X1 U11460 ( .B1(n13691), .B2(n11938), .A(n11937), .ZN(n11945) );
  OR2_X1 U11461 ( .A1(n10532), .A2(n10531), .ZN(n19664) );
  OR2_X1 U11462 ( .A1(n10532), .A2(n10526), .ZN(n19630) );
  NOR2_X1 U11463 ( .A1(n17692), .A2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17678) );
  AND2_X1 U11464 ( .A1(n13811), .A2(n9926), .ZN(n14131) );
  OR2_X1 U11465 ( .A1(n10528), .A2(n10530), .ZN(n10601) );
  NAND2_X1 U11466 ( .A1(n18011), .A2(n17613), .ZN(n11609) );
  BUF_X2 U11467 ( .A(n10522), .Z(n13691) );
  OR2_X1 U11468 ( .A1(n10522), .A2(n14598), .ZN(n10532) );
  OR2_X2 U11469 ( .A1(n12505), .A2(n12506), .ZN(n12558) );
  NAND2_X2 U11470 ( .A1(n14774), .A2(n12509), .ZN(n14773) );
  OR2_X1 U11471 ( .A1(n11607), .A2(n10099), .ZN(n10098) );
  NAND2_X1 U11472 ( .A1(n18129), .A2(n18593), .ZN(n18091) );
  NAND2_X1 U11473 ( .A1(n9985), .A2(n12477), .ZN(n12505) );
  NAND2_X1 U11474 ( .A1(n12555), .A2(n12554), .ZN(n12557) );
  CLKBUF_X1 U11475 ( .A(n13764), .Z(n20197) );
  CLKBUF_X2 U11476 ( .A(n10504), .Z(n14598) );
  NAND2_X1 U11477 ( .A1(n11927), .A2(n11926), .ZN(n15648) );
  AND2_X1 U11478 ( .A1(n18985), .A2(n10501), .ZN(n10523) );
  AND2_X1 U11479 ( .A1(n13603), .A2(n13602), .ZN(n13628) );
  OAI22_X1 U11480 ( .A1(n13752), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n13179), 
        .B2(n12542), .ZN(n9984) );
  CLKBUF_X1 U11481 ( .A(n13752), .Z(n20534) );
  NOR2_X2 U11482 ( .A1(n13356), .A2(n10512), .ZN(n10996) );
  XNOR2_X1 U11483 ( .A(n13513), .B(n20277), .ZN(n20397) );
  NAND2_X1 U11484 ( .A1(n10497), .A2(n10039), .ZN(n15646) );
  AND2_X1 U11485 ( .A1(n9963), .A2(n9962), .ZN(n16629) );
  NAND2_X1 U11486 ( .A1(n10477), .A2(n10476), .ZN(n10269) );
  CLKBUF_X1 U11487 ( .A(n13977), .Z(n20535) );
  NOR2_X1 U11488 ( .A1(n19156), .A2(n19157), .ZN(n19203) );
  OAI21_X1 U11489 ( .B1(n17760), .B2(n10106), .A(n10105), .ZN(n17752) );
  XNOR2_X1 U11490 ( .A(n10482), .B(n10483), .ZN(n10490) );
  OR2_X1 U11491 ( .A1(n10484), .A2(n10483), .ZN(n10485) );
  XNOR2_X1 U11492 ( .A(n11041), .B(n11042), .ZN(n11038) );
  INV_X2 U11493 ( .A(n15201), .ZN(n15259) );
  NOR2_X1 U11494 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n10856), .ZN(n10866) );
  NOR3_X2 U11495 ( .A1(n15672), .A2(n18600), .A3(n15671), .ZN(n18608) );
  OR2_X1 U11496 ( .A1(n10475), .A2(n10474), .ZN(n10476) );
  NAND2_X1 U11497 ( .A1(n9981), .A2(n20238), .ZN(n12483) );
  NAND2_X1 U11498 ( .A1(n12423), .A2(n12422), .ZN(n20170) );
  NAND2_X1 U11499 ( .A1(n10456), .A2(n10455), .ZN(n10474) );
  NAND2_X1 U11500 ( .A1(n10195), .A2(n10481), .ZN(n10483) );
  XNOR2_X1 U11501 ( .A(n11599), .B(n11598), .ZN(n17760) );
  INV_X2 U11502 ( .A(n19062), .ZN(n13451) );
  NAND2_X1 U11503 ( .A1(n10461), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10456) );
  OAI211_X1 U11504 ( .C1(n11117), .C2(n14023), .A(n10489), .B(n10488), .ZN(
        n11042) );
  NAND2_X1 U11505 ( .A1(n10461), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10195) );
  NOR2_X1 U11506 ( .A1(n11250), .A2(n10234), .ZN(n10233) );
  BUF_X2 U11507 ( .A(n11117), .Z(n11128) );
  NAND2_X2 U11508 ( .A1(n18163), .A2(n17393), .ZN(n17457) );
  INV_X1 U11509 ( .A(n10461), .ZN(n10487) );
  NAND2_X1 U11510 ( .A1(n12540), .A2(n12539), .ZN(n20277) );
  OAI21_X1 U11511 ( .B1(n17787), .B2(n10096), .A(n10095), .ZN(n17772) );
  AND2_X1 U11512 ( .A1(n10784), .A2(n10140), .ZN(n10850) );
  INV_X2 U11513 ( .A(n13293), .ZN(n18966) );
  NOR2_X1 U11514 ( .A1(n11242), .A2(n11241), .ZN(n11249) );
  NAND2_X1 U11515 ( .A1(n11739), .A2(n11730), .ZN(n18644) );
  AND2_X1 U11516 ( .A1(n10780), .A2(n10779), .ZN(n10784) );
  INV_X1 U11517 ( .A(n11124), .ZN(n11066) );
  INV_X1 U11518 ( .A(n11726), .ZN(n11730) );
  XNOR2_X1 U11519 ( .A(n11592), .B(n11591), .ZN(n17787) );
  NOR2_X1 U11520 ( .A1(n10683), .A2(n10699), .ZN(n10780) );
  NOR2_X1 U11521 ( .A1(n11726), .A2(n14315), .ZN(n17390) );
  AOI22_X1 U11522 ( .A1(n14166), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n16331), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10455) );
  NAND2_X1 U11523 ( .A1(n9979), .A2(n9978), .ZN(n10462) );
  NOR2_X1 U11524 ( .A1(n10165), .A2(n13725), .ZN(n10164) );
  NOR2_X2 U11525 ( .A1(n14315), .A2(n15765), .ZN(n17190) );
  NOR2_X1 U11526 ( .A1(n18167), .A2(n15672), .ZN(n11898) );
  NOR2_X1 U11527 ( .A1(n11590), .A2(n9893), .ZN(n11592) );
  CLKBUF_X2 U11528 ( .A(n10454), .Z(n14166) );
  OAI21_X1 U11529 ( .B1(n15676), .B2(n14314), .A(n18643), .ZN(n15765) );
  INV_X1 U11530 ( .A(n11207), .ZN(n10429) );
  NAND2_X1 U11531 ( .A1(n12395), .A2(n13620), .ZN(n13544) );
  OR2_X1 U11532 ( .A1(n11215), .A2(n10418), .ZN(n10454) );
  XNOR2_X1 U11533 ( .A(n13610), .B(n13651), .ZN(n13652) );
  AND2_X1 U11534 ( .A1(n13475), .A2(n13474), .ZN(n13477) );
  OAI21_X1 U11535 ( .B1(n10449), .B2(n10453), .A(n10452), .ZN(n11202) );
  OR2_X1 U11536 ( .A1(n11900), .A2(n11728), .ZN(n11748) );
  NOR3_X1 U11537 ( .A1(n18587), .A2(n11733), .A3(n11701), .ZN(n11728) );
  INV_X1 U11538 ( .A(n12909), .ZN(n13068) );
  AOI211_X2 U11539 ( .C1(n11756), .C2(n11755), .A(n11754), .B(n11753), .ZN(
        n18788) );
  NOR2_X1 U11540 ( .A1(n18188), .A2(n18171), .ZN(n11738) );
  MUX2_X1 U11541 ( .A(n11224), .B(n10420), .S(n11197), .Z(n10422) );
  AOI211_X1 U11542 ( .C1(n10434), .C2(n16332), .A(n16331), .B(n21095), .ZN(
        n16336) );
  NOR2_X2 U11543 ( .A1(n17548), .A2(n17549), .ZN(n17532) );
  NOR2_X1 U11544 ( .A1(n17334), .A2(n11773), .ZN(n11594) );
  OR2_X1 U11545 ( .A1(n13547), .A2(n13599), .ZN(n13614) );
  INV_X1 U11546 ( .A(n10465), .ZN(n11194) );
  OR2_X1 U11547 ( .A1(n11169), .A2(n10424), .ZN(n11165) );
  NAND2_X1 U11548 ( .A1(n11776), .A2(n11765), .ZN(n11773) );
  AND2_X2 U11549 ( .A1(n10669), .A2(n10668), .ZN(n10960) );
  NAND2_X1 U11550 ( .A1(n17569), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17548) );
  CLKBUF_X1 U11551 ( .A(n10992), .Z(n16321) );
  NAND2_X1 U11552 ( .A1(n12399), .A2(n12398), .ZN(n15156) );
  AND2_X1 U11553 ( .A1(n18178), .A2(n17193), .ZN(n11733) );
  NAND2_X1 U11554 ( .A1(n11220), .A2(n9826), .ZN(n11440) );
  NAND2_X2 U11555 ( .A1(n12239), .A2(n11220), .ZN(n11233) );
  OR2_X1 U11556 ( .A1(n10992), .A2(n10435), .ZN(n10436) );
  NAND2_X1 U11557 ( .A1(n13131), .A2(n13562), .ZN(n13547) );
  INV_X1 U11558 ( .A(n11772), .ZN(n15768) );
  INV_X1 U11559 ( .A(n18178), .ZN(n17201) );
  AND2_X1 U11560 ( .A1(n10689), .A2(n19199), .ZN(n12239) );
  CLKBUF_X1 U11561 ( .A(n10445), .Z(n13389) );
  NAND3_X1 U11562 ( .A1(n11556), .A2(n11555), .A3(n11554), .ZN(n11765) );
  NAND2_X1 U11563 ( .A1(n13621), .A2(n20146), .ZN(n13128) );
  OR2_X1 U11564 ( .A1(n12388), .A2(n20139), .ZN(n13565) );
  INV_X1 U11565 ( .A(n11589), .ZN(n11776) );
  AND2_X1 U11566 ( .A1(n12404), .A2(n13165), .ZN(n13562) );
  INV_X4 U11567 ( .A(n10672), .ZN(n10689) );
  AND2_X1 U11568 ( .A1(n20150), .A2(n13080), .ZN(n13509) );
  INV_X1 U11569 ( .A(n12396), .ZN(n13621) );
  INV_X1 U11570 ( .A(n10441), .ZN(n10424) );
  NOR2_X2 U11571 ( .A1(n11636), .A2(n11635), .ZN(n18163) );
  NAND2_X1 U11572 ( .A1(n10425), .A2(n10672), .ZN(n10439) );
  AND2_X1 U11573 ( .A1(n9896), .A2(n10170), .ZN(n18178) );
  AND3_X1 U11574 ( .A1(n11553), .A2(n11552), .A3(n11551), .ZN(n11556) );
  INV_X1 U11575 ( .A(n13867), .ZN(n9833) );
  AND2_X1 U11576 ( .A1(n12393), .A2(n20146), .ZN(n9840) );
  CLKBUF_X1 U11577 ( .A(n13080), .Z(n20154) );
  INV_X1 U11578 ( .A(n20139), .ZN(n13538) );
  AND4_X2 U11579 ( .A1(n12313), .A2(n12312), .A3(n12311), .A4(n12310), .ZN(
        n20150) );
  NAND2_X1 U11580 ( .A1(n10369), .A2(n10368), .ZN(n19180) );
  INV_X2 U11581 ( .A(U212), .ZN(n16436) );
  AND4_X1 U11582 ( .A1(n12297), .A2(n12296), .A3(n12295), .A4(n12294), .ZN(
        n12313) );
  NAND2_X1 U11583 ( .A1(n10334), .A2(n16293), .ZN(n10335) );
  AND4_X1 U11584 ( .A1(n12326), .A2(n12325), .A3(n12324), .A4(n12323), .ZN(
        n12331) );
  AND4_X2 U11585 ( .A1(n12283), .A2(n12282), .A3(n12281), .A4(n12280), .ZN(
        n12402) );
  NAND2_X1 U11586 ( .A1(n11691), .A2(n10168), .ZN(n10167) );
  NOR2_X2 U11587 ( .A1(n20117), .A2(n20120), .ZN(n20118) );
  AND4_X1 U11588 ( .A1(n12374), .A2(n12373), .A3(n12372), .A4(n12371), .ZN(
        n12385) );
  AND4_X1 U11589 ( .A1(n12270), .A2(n12269), .A3(n12268), .A4(n12267), .ZN(
        n12281) );
  AND4_X1 U11590 ( .A1(n12263), .A2(n12264), .A3(n12262), .A4(n12261), .ZN(
        n12282) );
  AND4_X1 U11591 ( .A1(n12305), .A2(n12304), .A3(n12303), .A4(n12302), .ZN(
        n12311) );
  AND4_X1 U11592 ( .A1(n12359), .A2(n12358), .A3(n12357), .A4(n12356), .ZN(
        n12360) );
  AND4_X1 U11593 ( .A1(n12321), .A2(n12320), .A3(n12319), .A4(n12318), .ZN(
        n9878) );
  AND4_X1 U11594 ( .A1(n12347), .A2(n12346), .A3(n12345), .A4(n12344), .ZN(
        n12363) );
  AND4_X1 U11595 ( .A1(n12301), .A2(n12300), .A3(n12299), .A4(n12298), .ZN(
        n12312) );
  AND4_X1 U11596 ( .A1(n12309), .A2(n12308), .A3(n12307), .A4(n12306), .ZN(
        n12310) );
  AND4_X1 U11597 ( .A1(n12351), .A2(n12350), .A3(n12349), .A4(n12348), .ZN(
        n12362) );
  AND4_X1 U11598 ( .A1(n12279), .A2(n12278), .A3(n12277), .A4(n12276), .ZN(
        n12280) );
  AND4_X1 U11599 ( .A1(n12355), .A2(n12354), .A3(n12353), .A4(n12352), .ZN(
        n12361) );
  AND4_X1 U11600 ( .A1(n12259), .A2(n12258), .A3(n12257), .A4(n12256), .ZN(
        n12283) );
  AND4_X1 U11601 ( .A1(n12382), .A2(n12381), .A3(n12380), .A4(n12379), .ZN(
        n12383) );
  INV_X2 U11602 ( .A(n17142), .ZN(n17107) );
  AND4_X1 U11603 ( .A1(n12378), .A2(n12377), .A3(n12376), .A4(n12375), .ZN(
        n12384) );
  INV_X2 U11604 ( .A(n11715), .ZN(n17140) );
  INV_X2 U11605 ( .A(n14536), .ZN(n10129) );
  NOR2_X1 U11606 ( .A1(n17742), .A2(n17757), .ZN(n17716) );
  CLKBUF_X3 U11607 ( .A(n15657), .Z(n17143) );
  NAND2_X2 U11608 ( .A1(n18739), .A2(n18677), .ZN(n18720) );
  INV_X4 U11609 ( .A(n10310), .ZN(n17153) );
  INV_X2 U11610 ( .A(n20102), .ZN(n13703) );
  AND3_X1 U11611 ( .A1(n9994), .A2(n9993), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10343) );
  AND3_X1 U11612 ( .A1(n9974), .A2(n9973), .A3(n16293), .ZN(n10303) );
  AND2_X1 U11614 ( .A1(n10394), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10398) );
  OR2_X1 U11615 ( .A1(n11500), .A2(n11499), .ZN(n10310) );
  NOR2_X1 U11616 ( .A1(n18601), .A2(n11500), .ZN(n11544) );
  OAI21_X2 U11617 ( .B1(n12248), .B2(n12247), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n19158) );
  AND2_X2 U11618 ( .A1(n12272), .A2(n13739), .ZN(n12496) );
  NOR2_X1 U11619 ( .A1(n18601), .A2(n11498), .ZN(n11545) );
  AND2_X2 U11620 ( .A1(n12274), .A2(n13745), .ZN(n12491) );
  OR3_X1 U11621 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n11499), .ZN(n11684) );
  NOR3_X2 U11622 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n16880), .ZN(n11581) );
  OR2_X1 U11623 ( .A1(n16880), .A2(n11500), .ZN(n16974) );
  INV_X2 U11624 ( .A(n16477), .ZN(n16479) );
  OAI221_X1 U11625 ( .B1(n20924), .B2(keyinput168), .C1(n20923), .C2(
        keyinput203), .A(n20922), .ZN(n20932) );
  NOR2_X1 U11626 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n13071), .ZN(
        n12265) );
  NOR2_X1 U11627 ( .A1(n10190), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12273) );
  AND2_X1 U11628 ( .A1(n13554), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12274) );
  AND2_X2 U11629 ( .A1(n12260), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12271) );
  AND2_X1 U11630 ( .A1(n10108), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12272) );
  AND2_X2 U11631 ( .A1(n13740), .A2(n13739), .ZN(n12984) );
  NAND2_X1 U11632 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18774), .ZN(
        n11499) );
  NAND3_X2 U11633 ( .A1(n18810), .A2(n18799), .A3(n18809), .ZN(n18138) );
  NAND2_X1 U11634 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18762), .ZN(
        n11498) );
  OR2_X1 U11635 ( .A1(n18601), .A2(n14306), .ZN(n11702) );
  AOI22_X1 U11636 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n20915), .B2(n18769), .ZN(
        n11752) );
  INV_X1 U11637 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10469) );
  NOR2_X2 U11638 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14088) );
  INV_X1 U11639 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13554) );
  AND2_X2 U11640 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13739) );
  NOR2_X2 U11641 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12266) );
  INV_X1 U11642 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12260) );
  AND2_X1 U11643 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13745) );
  NOR2_X1 U11644 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12275) );
  NOR2_X2 U11645 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20570) );
  NAND2_X2 U11646 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18601) );
  NAND3_X1 U11647 ( .A1(n10302), .A2(n10355), .A3(n10354), .ZN(n10356) );
  INV_X1 U11648 ( .A(n11010), .ZN(n10277) );
  XNOR2_X1 U11649 ( .A(n11815), .B(n11814), .ZN(n11828) );
  OAI21_X2 U11650 ( .B1(n10472), .B2(n10471), .A(n10470), .ZN(n10494) );
  NAND2_X1 U11651 ( .A1(n15429), .A2(n15428), .ZN(n15427) );
  OAI21_X1 U11652 ( .B1(n12484), .B2(n13071), .A(n12408), .ZN(n12410) );
  OR2_X1 U11653 ( .A1(n15050), .A2(n9945), .ZN(n13249) );
  OR2_X1 U11654 ( .A1(n15050), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14880) );
  NAND2_X1 U11655 ( .A1(n10276), .A2(n14017), .ZN(n11014) );
  AND2_X1 U11656 ( .A1(n10434), .A2(n10423), .ZN(n11050) );
  AND2_X2 U11657 ( .A1(n10428), .A2(n10270), .ZN(n11192) );
  NAND2_X1 U11658 ( .A1(n12454), .A2(n12455), .ZN(n12422) );
  AND2_X1 U11659 ( .A1(n13691), .A2(n10513), .ZN(n19210) );
  NAND2_X1 U11660 ( .A1(n13691), .A2(n10503), .ZN(n10792) );
  INV_X1 U11661 ( .A(n9891), .ZN(n9835) );
  NAND2_X1 U11662 ( .A1(n9836), .A2(n11873), .ZN(n11877) );
  NOR2_X1 U11663 ( .A1(n11874), .A2(n9835), .ZN(n9836) );
  NAND2_X1 U11664 ( .A1(n10263), .A2(n9888), .ZN(n11873) );
  NAND2_X1 U11665 ( .A1(n10271), .A2(n10019), .ZN(n9837) );
  NAND2_X1 U11666 ( .A1(n9995), .A2(n9996), .ZN(n9838) );
  NAND2_X1 U11667 ( .A1(n10271), .A2(n10019), .ZN(n16221) );
  NAND2_X1 U11668 ( .A1(n9995), .A2(n9996), .ZN(n14178) );
  NAND2_X1 U11669 ( .A1(n14681), .A2(n9839), .ZN(n14733) );
  AND2_X1 U11670 ( .A1(n14682), .A2(n10116), .ZN(n9839) );
  INV_X1 U11671 ( .A(n9847), .ZN(n14725) );
  NAND2_X1 U11672 ( .A1(n13727), .A2(n11950), .ZN(n9841) );
  OR2_X2 U11673 ( .A1(n9841), .A2(n9842), .ZN(n13865) );
  OR2_X1 U11674 ( .A1(n9833), .A2(n11951), .ZN(n9842) );
  NOR2_X2 U11675 ( .A1(n14770), .A2(n14771), .ZN(n14769) );
  NAND2_X2 U11676 ( .A1(n10942), .A2(n10855), .ZN(n10865) );
  NOR2_X2 U11677 ( .A1(n10938), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10941) );
  OAI21_X2 U11678 ( .B1(n10254), .B2(n10255), .A(n14470), .ZN(n10253) );
  NOR2_X2 U11679 ( .A1(n10889), .A2(n10884), .ZN(n10885) );
  NOR2_X2 U11680 ( .A1(n16597), .A2(n16853), .ZN(n16585) );
  NOR2_X2 U11681 ( .A1(n16629), .A2(n16853), .ZN(n16618) );
  NOR2_X2 U11682 ( .A1(n16529), .A2(n9964), .ZN(n16647) );
  XOR2_X2 U11683 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n16349), .Z(
        n16529) );
  NAND2_X1 U11684 ( .A1(n14131), .A2(n13316), .ZN(n15166) );
  NOR2_X2 U11685 ( .A1(n13766), .A2(n13767), .ZN(n13811) );
  INV_X2 U11686 ( .A(n19199), .ZN(n12237) );
  NOR2_X2 U11687 ( .A1(n17416), .A2(n17222), .ZN(n17218) );
  NOR4_X4 U11688 ( .A1(n17315), .A2(n17444), .A3(n17287), .A4(n17196), .ZN(
        n17288) );
  NAND2_X1 U11689 ( .A1(n10038), .A2(n13245), .ZN(n13246) );
  OAI21_X2 U11690 ( .B1(n13164), .B2(n13199), .A(n13163), .ZN(n13487) );
  XNOR2_X2 U11691 ( .A(n12522), .B(n12521), .ZN(n13164) );
  AND2_X1 U11692 ( .A1(n15598), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16212) );
  NAND2_X2 U11693 ( .A1(n10357), .A2(n10356), .ZN(n10441) );
  INV_X2 U11694 ( .A(n11816), .ZN(n10000) );
  NOR2_X2 U11695 ( .A1(n15196), .A2(n15195), .ZN(n15194) );
  NOR2_X4 U11696 ( .A1(n14077), .A2(n14129), .ZN(n14128) );
  NOR2_X2 U11697 ( .A1(n16759), .A2(n17119), .ZN(n17106) );
  NOR2_X2 U11698 ( .A1(n16985), .A2(n16986), .ZN(n16960) );
  NOR3_X2 U11699 ( .A1(n15664), .A2(n16714), .A3(n16733), .ZN(n17065) );
  AND2_X2 U11700 ( .A1(n9844), .A2(n9845), .ZN(n14710) );
  AND2_X1 U11701 ( .A1(n9846), .A2(n12912), .ZN(n9845) );
  INV_X1 U11702 ( .A(n14720), .ZN(n9846) );
  OR2_X1 U11703 ( .A1(n14733), .A2(n14734), .ZN(n9847) );
  NAND2_X1 U11704 ( .A1(n12558), .A2(n13774), .ZN(n20121) );
  NAND2_X1 U11705 ( .A1(n12483), .A2(n20170), .ZN(n13977) );
  NOR2_X2 U11706 ( .A1(n15530), .A2(n15543), .ZN(n15406) );
  NOR2_X1 U11707 ( .A1(n11499), .A2(n11498), .ZN(n11672) );
  NAND2_X1 U11708 ( .A1(n12393), .A2(n20146), .ZN(n12412) );
  AND2_X2 U11709 ( .A1(n12686), .A2(n10122), .ZN(n14239) );
  CLKBUF_X3 U11710 ( .A(n17809), .Z(n9848) );
  AND2_X2 U11712 ( .A1(n14301), .A2(n12783), .ZN(n14681) );
  NAND2_X2 U11713 ( .A1(n13722), .A2(n13721), .ZN(n13720) );
  NAND2_X2 U11714 ( .A1(n13650), .A2(n12531), .ZN(n13722) );
  OAI21_X2 U11715 ( .B1(n18589), .B2(n18600), .A(n18588), .ZN(n18615) );
  NAND2_X1 U11716 ( .A1(n11737), .A2(n11736), .ZN(n18600) );
  AND2_X2 U11717 ( .A1(n14710), .A2(n14711), .ZN(n14667) );
  NOR2_X2 U11718 ( .A1(n12403), .A2(n13128), .ZN(n13501) );
  OAI21_X2 U11719 ( .B1(n12406), .B2(n12409), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12484) );
  OR2_X2 U11720 ( .A1(n13604), .A2(n12405), .ZN(n12409) );
  AND3_X1 U11721 ( .A1(n13620), .A2(n12392), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n13108) );
  NOR2_X1 U11722 ( .A1(n19240), .A2(n10619), .ZN(n10621) );
  NAND2_X1 U11723 ( .A1(n14450), .A2(n10128), .ZN(n10127) );
  INV_X1 U11724 ( .A(n14654), .ZN(n10128) );
  NAND2_X1 U11725 ( .A1(n10256), .A2(n11202), .ZN(n10466) );
  NAND2_X1 U11726 ( .A1(n14599), .A2(n14611), .ZN(n20013) );
  INV_X1 U11727 ( .A(n10960), .ZN(n11020) );
  NAND2_X1 U11728 ( .A1(n9900), .A2(n12556), .ZN(n12605) );
  NAND2_X1 U11729 ( .A1(n10827), .A2(n10826), .ZN(n11012) );
  OR2_X1 U11730 ( .A1(n10810), .A2(n10809), .ZN(n10827) );
  OAI21_X1 U11731 ( .B1(n10792), .B2(n10612), .A(n10611), .ZN(n10615) );
  NAND2_X1 U11732 ( .A1(n19210), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n10611) );
  NOR2_X2 U11733 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10538) );
  INV_X1 U11734 ( .A(n13080), .ZN(n13165) );
  OR2_X1 U11735 ( .A1(n15156), .A2(n20706), .ZN(n13033) );
  OR2_X1 U11736 ( .A1(n10017), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10014) );
  NOR2_X1 U11737 ( .A1(n14841), .A2(n10179), .ZN(n10017) );
  OR2_X1 U11738 ( .A1(n12466), .A2(n12465), .ZN(n13166) );
  AOI21_X1 U11739 ( .B1(n12522), .B2(n12521), .A(n13222), .ZN(n12516) );
  XNOR2_X1 U11740 ( .A(n9984), .B(n12504), .ZN(n12506) );
  INV_X1 U11741 ( .A(n12422), .ZN(n9981) );
  OAI22_X1 U11742 ( .A1(n15149), .A2(n20813), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n20794), .ZN(n20172) );
  NAND2_X1 U11743 ( .A1(n10854), .A2(n13951), .ZN(n10856) );
  NOR2_X1 U11744 ( .A1(n10144), .A2(n10143), .ZN(n10142) );
  INV_X1 U11745 ( .A(n10783), .ZN(n10144) );
  NAND2_X1 U11746 ( .A1(n14542), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12081) );
  NAND2_X1 U11747 ( .A1(n10307), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10060) );
  NAND2_X1 U11748 ( .A1(n10949), .A2(n10950), .ZN(n10246) );
  NOR2_X1 U11749 ( .A1(n10660), .A2(n10659), .ZN(n10669) );
  INV_X1 U11750 ( .A(n14025), .ZN(n10232) );
  NAND2_X1 U11751 ( .A1(n18178), .A2(n9882), .ZN(n11726) );
  NOR2_X2 U11752 ( .A1(n17468), .A2(n17812), .ZN(n16520) );
  NOR2_X1 U11753 ( .A1(n18175), .A2(n17193), .ZN(n18587) );
  INV_X1 U11754 ( .A(n10126), .ZN(n10124) );
  OR2_X1 U11755 ( .A1(n12997), .A2(n20977), .ZN(n13016) );
  NAND2_X1 U11756 ( .A1(n12955), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12976) );
  NAND2_X1 U11757 ( .A1(n15050), .A2(n9918), .ZN(n9986) );
  INV_X1 U11758 ( .A(n14977), .ZN(n9987) );
  NOR2_X1 U11759 ( .A1(n9879), .A2(n9989), .ZN(n9988) );
  INV_X1 U11760 ( .A(n13230), .ZN(n9989) );
  OR3_X1 U11761 ( .A1(n20013), .A2(n13601), .A3(n12396), .ZN(n13602) );
  AOI21_X1 U11762 ( .B1(n10981), .B2(n10980), .A(n10979), .ZN(n11150) );
  AND2_X1 U11763 ( .A1(n16325), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10979) );
  INV_X1 U11764 ( .A(n10978), .ZN(n10981) );
  AND2_X1 U11765 ( .A1(n10940), .A2(n10942), .ZN(n16117) );
  NAND2_X1 U11766 ( .A1(n10852), .A2(n11269), .ZN(n10942) );
  INV_X1 U11767 ( .A(n11132), .ZN(n10219) );
  AND2_X1 U11768 ( .A1(n11875), .A2(n11210), .ZN(n10946) );
  AND2_X1 U11769 ( .A1(n15200), .A2(n15190), .ZN(n11882) );
  NOR2_X2 U11770 ( .A1(n15208), .A2(n15198), .ZN(n15200) );
  AND2_X1 U11771 ( .A1(n10052), .A2(n11809), .ZN(n10051) );
  OR2_X1 U11772 ( .A1(n11810), .A2(n9910), .ZN(n10052) );
  INV_X1 U11773 ( .A(n11810), .ZN(n10053) );
  AND2_X1 U11774 ( .A1(n14089), .A2(n10469), .ZN(n10471) );
  NAND3_X1 U11775 ( .A1(n10464), .A2(n10487), .A3(n10463), .ZN(n10493) );
  AND2_X1 U11776 ( .A1(n10460), .A2(n10459), .ZN(n10464) );
  AOI21_X1 U11777 ( .B1(n11050), .B2(P2_REIP_REG_0__SCAN_IN), .A(n10458), .ZN(
        n10459) );
  INV_X1 U11778 ( .A(n11219), .ZN(n11209) );
  INV_X1 U11779 ( .A(n15648), .ZN(n13583) );
  AOI21_X1 U11780 ( .B1(n14043), .B2(n11924), .A(n11923), .ZN(n13572) );
  NOR2_X1 U11781 ( .A1(n10502), .A2(n10520), .ZN(n10500) );
  NAND2_X1 U11782 ( .A1(n10412), .A2(n16293), .ZN(n10242) );
  NOR2_X1 U11783 ( .A1(n16566), .A2(n17481), .ZN(n16565) );
  NAND2_X1 U11784 ( .A1(n18795), .A2(n17352), .ZN(n14315) );
  INV_X1 U11785 ( .A(n18163), .ZN(n18795) );
  AND2_X1 U11786 ( .A1(n11216), .A2(n13289), .ZN(n19854) );
  INV_X1 U11787 ( .A(n10996), .ZN(n19142) );
  INV_X1 U11788 ( .A(n16272), .ZN(n16285) );
  INV_X1 U11789 ( .A(n10596), .ZN(n10138) );
  INV_X1 U11791 ( .A(n13226), .ZN(n12474) );
  INV_X1 U11792 ( .A(n12394), .ZN(n12395) );
  MUX2_X1 U11793 ( .A(n13538), .B(n12397), .S(n12393), .Z(n12394) );
  OAI21_X1 U11794 ( .B1(n12401), .B2(n12387), .A(n13131), .ZN(n13541) );
  NAND2_X1 U11795 ( .A1(n20397), .A2(n20706), .ZN(n12555) );
  NAND2_X1 U11796 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n11546) );
  NAND2_X1 U11797 ( .A1(n18754), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11500) );
  NAND2_X1 U11798 ( .A1(n13567), .A2(n10160), .ZN(n13651) );
  NAND2_X1 U11799 ( .A1(n10159), .A2(n14615), .ZN(n10160) );
  NOR2_X1 U11800 ( .A1(n13570), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n10159) );
  NOR2_X1 U11801 ( .A1(n10118), .A2(n14745), .ZN(n10117) );
  INV_X1 U11802 ( .A(n10119), .ZN(n10118) );
  INV_X1 U11803 ( .A(n14266), .ZN(n12693) );
  INV_X1 U11804 ( .A(n13824), .ZN(n10114) );
  INV_X1 U11805 ( .A(n14011), .ZN(n10113) );
  NAND2_X1 U11806 ( .A1(n14909), .A2(n9849), .ZN(n10033) );
  INV_X1 U11807 ( .A(n10033), .ZN(n10032) );
  NOR2_X1 U11808 ( .A1(n10147), .A2(n14688), .ZN(n10146) );
  INV_X1 U11809 ( .A(n14762), .ZN(n10147) );
  NAND2_X1 U11810 ( .A1(n13225), .A2(n13232), .ZN(n14936) );
  AND2_X1 U11811 ( .A1(n10150), .A2(n14148), .ZN(n10149) );
  AND2_X1 U11812 ( .A1(n13997), .A2(n10151), .ZN(n10150) );
  INV_X1 U11813 ( .A(n14062), .ZN(n10151) );
  OR2_X1 U11814 ( .A1(n20146), .A2(n20124), .ZN(n14437) );
  NAND2_X1 U11815 ( .A1(n20150), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12542) );
  NAND2_X1 U11816 ( .A1(n12515), .A2(n12516), .ZN(n9985) );
  NAND2_X1 U11817 ( .A1(n10922), .A2(n10942), .ZN(n10919) );
  AND2_X1 U11818 ( .A1(n10865), .A2(n9913), .ZN(n10892) );
  INV_X1 U11819 ( .A(n12076), .ZN(n12049) );
  AND2_X1 U11820 ( .A1(n15267), .A2(n14503), .ZN(n10244) );
  NAND2_X1 U11821 ( .A1(n13580), .A2(n19169), .ZN(n12193) );
  NOR2_X1 U11822 ( .A1(n10207), .A2(n10206), .ZN(n10205) );
  INV_X1 U11823 ( .A(n15237), .ZN(n10206) );
  INV_X1 U11824 ( .A(n10208), .ZN(n10207) );
  NAND2_X1 U11825 ( .A1(n10236), .A2(n15325), .ZN(n10235) );
  INV_X1 U11826 ( .A(n15167), .ZN(n10236) );
  NOR2_X1 U11827 ( .A1(n16163), .A2(n10077), .ZN(n10076) );
  INV_X1 U11828 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11025) );
  OAI22_X1 U11829 ( .A1(n10487), .A2(n16293), .B1(n19853), .B2(n11933), .ZN(
        n11041) );
  INV_X1 U11830 ( .A(n13643), .ZN(n11049) );
  NAND2_X1 U11831 ( .A1(n10486), .A2(n10485), .ZN(n11040) );
  NAND2_X1 U11832 ( .A1(n10933), .A2(n10264), .ZN(n10263) );
  NOR2_X1 U11833 ( .A1(n10937), .A2(n10265), .ZN(n10264) );
  INV_X1 U11834 ( .A(n10932), .ZN(n10265) );
  INV_X1 U11835 ( .A(n15227), .ZN(n10214) );
  NAND2_X1 U11836 ( .A1(n10897), .A2(n16178), .ZN(n10048) );
  NAND2_X1 U11837 ( .A1(n10044), .A2(n14217), .ZN(n10043) );
  NOR2_X1 U11838 ( .A1(n16225), .A2(n10259), .ZN(n10258) );
  INV_X1 U11839 ( .A(n15631), .ZN(n10259) );
  INV_X1 U11840 ( .A(n13964), .ZN(n10241) );
  INV_X1 U11841 ( .A(n10275), .ZN(n10273) );
  INV_X1 U11842 ( .A(n11012), .ZN(n10828) );
  INV_X1 U11843 ( .A(n10829), .ZN(n9975) );
  AND2_X1 U11844 ( .A1(n11049), .A2(n10225), .ZN(n10224) );
  INV_X1 U11845 ( .A(n13637), .ZN(n10225) );
  INV_X1 U11846 ( .A(n13644), .ZN(n10226) );
  INV_X1 U11847 ( .A(n13851), .ZN(n10234) );
  OAI21_X1 U11848 ( .B1(n10600), .B2(n10599), .A(n10598), .ZN(n10646) );
  OAI21_X1 U11849 ( .B1(n10644), .B2(n10643), .A(n10642), .ZN(n10645) );
  NAND2_X1 U11850 ( .A1(n11189), .A2(n9894), .ZN(n9978) );
  NAND2_X1 U11851 ( .A1(n10454), .A2(n9890), .ZN(n9979) );
  AND3_X1 U11852 ( .A1(n10563), .A2(n10562), .A3(n10561), .ZN(n11227) );
  OR2_X1 U11853 ( .A1(n12193), .A2(n19173), .ZN(n11928) );
  OAI21_X1 U11854 ( .B1(n14598), .B2(n11938), .A(n11919), .ZN(n11932) );
  AND2_X1 U11855 ( .A1(n10439), .A2(n12237), .ZN(n10270) );
  NAND2_X1 U11856 ( .A1(n12225), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n9994) );
  NAND2_X1 U11857 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n9993) );
  NAND2_X1 U11858 ( .A1(n12225), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n9974) );
  AOI22_X1 U11859 ( .A1(n12094), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10553), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10366) );
  AOI21_X1 U11860 ( .B1(n12225), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10352) );
  NAND2_X1 U11861 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n10351) );
  NAND4_X1 U11862 ( .A1(n19199), .A2(n19180), .A3(n10441), .A4(n19174), .ZN(
        n10245) );
  INV_X1 U11863 ( .A(n11581), .ZN(n11715) );
  NAND2_X1 U11864 ( .A1(n17640), .A2(n9954), .ZN(n9957) );
  NOR2_X1 U11865 ( .A1(n17619), .A2(n9955), .ZN(n9954) );
  INV_X1 U11866 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n9955) );
  NOR2_X1 U11867 ( .A1(n17327), .A2(n11597), .ZN(n11601) );
  OR2_X1 U11868 ( .A1(n11615), .A2(n11614), .ZN(n11616) );
  NAND2_X1 U11869 ( .A1(n17528), .A2(n10092), .ZN(n10094) );
  AND2_X1 U11870 ( .A1(n11612), .A2(n10093), .ZN(n10092) );
  INV_X1 U11871 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10093) );
  AND2_X1 U11872 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n11595), .ZN(
        n11596) );
  XNOR2_X1 U11873 ( .A(n11765), .B(n11776), .ZN(n10086) );
  NOR2_X1 U11874 ( .A1(n17390), .A2(n15670), .ZN(n11737) );
  NAND2_X1 U11875 ( .A1(n14657), .A2(n10158), .ZN(n14641) );
  AND2_X1 U11876 ( .A1(n20012), .A2(n14601), .ZN(n13500) );
  AND2_X1 U11877 ( .A1(n20708), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13067) );
  AOI21_X1 U11878 ( .B1(n13920), .B2(n14859), .A(n13014), .ZN(n14450) );
  OAI21_X1 U11879 ( .B1(n13063), .B2(n14866), .A(n12996), .ZN(n14654) );
  AOI21_X1 U11880 ( .B1(n13920), .B2(n14874), .A(n12973), .ZN(n14668) );
  NAND2_X1 U11881 ( .A1(n12750), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12751) );
  NAND2_X1 U11882 ( .A1(n13225), .A2(n13240), .ZN(n15119) );
  NAND2_X1 U11883 ( .A1(n10158), .A2(n10154), .ZN(n10153) );
  INV_X1 U11884 ( .A(n14655), .ZN(n10154) );
  NAND2_X1 U11885 ( .A1(n14657), .A2(n10156), .ZN(n10155) );
  AND2_X1 U11886 ( .A1(n10158), .A2(n14616), .ZN(n10156) );
  INV_X1 U11887 ( .A(n10014), .ZN(n10010) );
  NAND2_X1 U11888 ( .A1(n14834), .A2(n9917), .ZN(n10008) );
  NAND2_X1 U11889 ( .A1(n10014), .A2(n14842), .ZN(n10009) );
  NAND2_X1 U11890 ( .A1(n14834), .A2(n14835), .ZN(n10006) );
  AND2_X1 U11891 ( .A1(n10017), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10012) );
  NAND2_X1 U11892 ( .A1(n10180), .A2(n13250), .ZN(n14844) );
  OR2_X1 U11893 ( .A1(n14834), .A2(n13225), .ZN(n10180) );
  INV_X1 U11894 ( .A(n15050), .ZN(n14886) );
  NAND2_X1 U11895 ( .A1(n14749), .A2(n14741), .ZN(n14742) );
  NOR2_X1 U11896 ( .A1(n10004), .A2(n10003), .ZN(n10002) );
  INV_X1 U11897 ( .A(n13231), .ZN(n10003) );
  NAND2_X1 U11898 ( .A1(n14282), .A2(n14283), .ZN(n14284) );
  NAND2_X1 U11899 ( .A1(n15943), .A2(n15942), .ZN(n15941) );
  NOR2_X1 U11900 ( .A1(n12487), .A2(n9983), .ZN(n9982) );
  INV_X1 U11901 ( .A(n12482), .ZN(n9983) );
  INV_X1 U11902 ( .A(n20503), .ZN(n20496) );
  INV_X1 U11903 ( .A(n20276), .ZN(n20528) );
  NOR2_X1 U11904 ( .A1(n20284), .A2(n20283), .ZN(n20599) );
  INV_X1 U11905 ( .A(n20172), .ZN(n20284) );
  NAND2_X1 U11906 ( .A1(n13122), .A2(n13121), .ZN(n14599) );
  NAND2_X1 U11907 ( .A1(n13138), .A2(n13078), .ZN(n13122) );
  AND2_X1 U11908 ( .A1(n10976), .A2(n10975), .ZN(n11146) );
  NAND2_X1 U11909 ( .A1(n14485), .A2(n10074), .ZN(n10073) );
  NOR2_X1 U11910 ( .A1(n14489), .A2(n18966), .ZN(n16127) );
  NAND2_X1 U11911 ( .A1(n10070), .A2(n15381), .ZN(n10071) );
  INV_X1 U11912 ( .A(n16127), .ZN(n10070) );
  NAND2_X1 U11913 ( .A1(n13323), .A2(n10079), .ZN(n10078) );
  INV_X1 U11914 ( .A(n10082), .ZN(n10079) );
  NAND2_X1 U11915 ( .A1(n10084), .A2(n16154), .ZN(n10085) );
  INV_X1 U11916 ( .A(n15169), .ZN(n10084) );
  AND2_X1 U11917 ( .A1(n9881), .A2(n10141), .ZN(n10140) );
  INV_X1 U11918 ( .A(n10842), .ZN(n10141) );
  OAI22_X1 U11919 ( .A1(n13282), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n19859), 
        .B2(n13281), .ZN(n13293) );
  NOR2_X1 U11920 ( .A1(n10201), .A2(n11441), .ZN(n10199) );
  AND2_X1 U11921 ( .A1(n10549), .A2(n10550), .ZN(n12065) );
  AND3_X1 U11922 ( .A1(n11421), .A2(n11420), .A3(n11419), .ZN(n15611) );
  AND3_X1 U11923 ( .A1(n11260), .A2(n11259), .A3(n11258), .ZN(n14025) );
  XNOR2_X1 U11924 ( .A(n11028), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13282) );
  NOR2_X1 U11925 ( .A1(n14473), .A2(n11869), .ZN(n11028) );
  AND2_X1 U11926 ( .A1(n9862), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10054) );
  OR2_X1 U11927 ( .A1(n10282), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10281) );
  NAND2_X1 U11928 ( .A1(n15360), .A2(n10280), .ZN(n10279) );
  AND2_X1 U11929 ( .A1(n10282), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10280) );
  OR2_X1 U11930 ( .A1(n10952), .A2(n10951), .ZN(n15366) );
  INV_X1 U11931 ( .A(n15410), .ZN(n10049) );
  INV_X1 U11932 ( .A(n9980), .ZN(n15416) );
  INV_X1 U11933 ( .A(n14133), .ZN(n10227) );
  AND2_X1 U11934 ( .A1(n13894), .A2(n9857), .ZN(n14156) );
  OR2_X1 U11935 ( .A1(n11801), .A2(n10048), .ZN(n10046) );
  NAND2_X1 U11936 ( .A1(n14218), .A2(n10845), .ZN(n10041) );
  NAND2_X1 U11937 ( .A1(n14113), .A2(n14112), .ZN(n10045) );
  XNOR2_X1 U11938 ( .A(n11003), .B(n14023), .ZN(n13886) );
  CLKBUF_X1 U11939 ( .A(n11215), .Z(n11216) );
  NAND2_X1 U11940 ( .A1(n13572), .A2(n13573), .ZN(n13575) );
  OR2_X1 U11941 ( .A1(n19296), .A2(n19826), .ZN(n19460) );
  AND2_X1 U11942 ( .A1(n19296), .A2(n19824), .ZN(n19589) );
  OR2_X1 U11943 ( .A1(n19449), .A2(n19837), .ZN(n19576) );
  NAND2_X1 U11944 ( .A1(n11162), .A2(n11152), .ZN(n16313) );
  NAND2_X1 U11945 ( .A1(n19065), .A2(n11151), .ZN(n11152) );
  INV_X1 U11946 ( .A(n17495), .ZN(n9969) );
  INV_X2 U11947 ( .A(n17004), .ZN(n17145) );
  NAND2_X1 U11948 ( .A1(n11671), .A2(n11670), .ZN(n17352) );
  NOR2_X2 U11949 ( .A1(n17588), .A2(n17589), .ZN(n17569) );
  NAND2_X1 U11950 ( .A1(n10089), .A2(n10087), .ZN(n10091) );
  AOI21_X1 U11951 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n10088), .A(
        n9864), .ZN(n10087) );
  OR2_X1 U11952 ( .A1(n18011), .A2(n17947), .ZN(n10089) );
  NOR2_X1 U11953 ( .A1(n10172), .A2(n10171), .ZN(n10170) );
  INV_X1 U11954 ( .A(n11697), .ZN(n10172) );
  NOR3_X1 U11955 ( .A1(n10169), .A2(n11689), .A3(n10167), .ZN(n10166) );
  INV_X1 U11956 ( .A(n18651), .ZN(n18643) );
  INV_X1 U11957 ( .A(n14774), .ZN(n14765) );
  NAND2_X1 U11958 ( .A1(n14774), .A2(n14452), .ZN(n14776) );
  OAI21_X1 U11959 ( .B1(n14902), .B2(n14903), .A(n10182), .ZN(n14904) );
  XNOR2_X1 U11960 ( .A(n14863), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15021) );
  NOR2_X1 U11961 ( .A1(n10182), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15747) );
  OR2_X1 U11962 ( .A1(n13258), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20102) );
  INV_X1 U11963 ( .A(n16014), .ZN(n20110) );
  AOI21_X1 U11964 ( .B1(n16062), .B2(n18984), .A(n16061), .ZN(n16063) );
  NOR2_X1 U11965 ( .A1(n16074), .A2(n18966), .ZN(n16057) );
  INV_X1 U11966 ( .A(n10039), .ZN(n10498) );
  NAND3_X1 U11967 ( .A1(n10216), .A2(n10215), .A3(n10217), .ZN(n16045) );
  NAND2_X1 U11968 ( .A1(n10221), .A2(n11132), .ZN(n10217) );
  OR2_X1 U11969 ( .A1(n11882), .A2(n10219), .ZN(n10216) );
  OR2_X1 U11970 ( .A1(n14475), .A2(n11884), .ZN(n16071) );
  NAND2_X1 U11971 ( .A1(n10315), .A2(n10202), .ZN(n10201) );
  INV_X1 U11972 ( .A(n13956), .ZN(n10202) );
  CLKBUF_X1 U11973 ( .A(n14077), .Z(n14078) );
  INV_X1 U11974 ( .A(n19837), .ZN(n19417) );
  OR2_X1 U11975 ( .A1(n19137), .A2(n13370), .ZN(n19150) );
  OR2_X1 U11976 ( .A1(n19827), .A2(n19585), .ZN(n19157) );
  NAND3_X1 U11977 ( .A1(n10132), .A2(n10131), .A3(n10964), .ZN(n10130) );
  NAND2_X1 U11978 ( .A1(n11889), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14516) );
  INV_X1 U11979 ( .A(n10949), .ZN(n11879) );
  AOI21_X1 U11980 ( .B1(n15580), .B2(n16285), .A(n10022), .ZN(n10021) );
  INV_X1 U11981 ( .A(n15578), .ZN(n10022) );
  OR2_X1 U11982 ( .A1(n15575), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10024) );
  INV_X1 U11983 ( .A(n16280), .ZN(n16271) );
  NAND2_X1 U11984 ( .A1(n11209), .A2(n11183), .ZN(n16278) );
  NAND2_X1 U11985 ( .A1(n11209), .A2(n11188), .ZN(n16272) );
  INV_X1 U11986 ( .A(n16278), .ZN(n16283) );
  INV_X1 U11987 ( .A(n19826), .ZN(n19824) );
  OR2_X1 U11988 ( .A1(n15646), .A2(n11938), .ZN(n11927) );
  XNOR2_X1 U11989 ( .A(n9952), .B(n9951), .ZN(n9950) );
  INV_X1 U11990 ( .A(n16534), .ZN(n9951) );
  NAND2_X1 U11991 ( .A1(n9953), .A2(n16837), .ZN(n9952) );
  INV_X1 U11992 ( .A(n16540), .ZN(n9947) );
  NOR2_X1 U11993 ( .A1(n17160), .A2(n17011), .ZN(n16997) );
  NAND2_X1 U11994 ( .A1(n17023), .A2(P3_EBX_REG_19__SCAN_IN), .ZN(n17011) );
  NOR2_X2 U11995 ( .A1(n16381), .A2(n17321), .ZN(n17724) );
  INV_X1 U11996 ( .A(n13079), .ZN(n13092) );
  INV_X1 U11997 ( .A(n19210), .ZN(n10794) );
  INV_X1 U11998 ( .A(n13509), .ZN(n13125) );
  NOR2_X1 U11999 ( .A1(n13092), .A2(n13134), .ZN(n13106) );
  INV_X1 U12000 ( .A(n19547), .ZN(n10788) );
  OR2_X1 U12001 ( .A1(n12553), .A2(n12552), .ZN(n13194) );
  AND3_X1 U12002 ( .A1(n12453), .A2(n12452), .A3(n12451), .ZN(n12475) );
  INV_X1 U12003 ( .A(n12558), .ZN(n12556) );
  NAND2_X1 U12004 ( .A1(n13537), .A2(n12509), .ZN(n13539) );
  INV_X1 U12005 ( .A(n20644), .ZN(n12534) );
  INV_X1 U12006 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13071) );
  NAND2_X1 U12007 ( .A1(n12409), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12479) );
  NOR2_X1 U12008 ( .A1(n14214), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10275) );
  NAND2_X1 U12009 ( .A1(n10778), .A2(n9998), .ZN(n10829) );
  OAI22_X1 U12010 ( .A1(n10617), .A2(n10754), .B1(n10752), .B2(n10616), .ZN(
        n10618) );
  OAI22_X1 U12011 ( .A1(n10609), .A2(n19580), .B1(n19630), .B2(n10608), .ZN(
        n10610) );
  NOR2_X1 U12012 ( .A1(n10480), .A2(n10319), .ZN(n10482) );
  NAND2_X1 U12013 ( .A1(n10521), .A2(n14043), .ZN(n10602) );
  OAI21_X1 U12014 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18762), .A(
        n11638), .ZN(n11639) );
  OR2_X1 U12015 ( .A1(n11642), .A2(n11643), .ZN(n11638) );
  OAI21_X1 U12016 ( .B1(n16490), .B2(n11731), .A(n18644), .ZN(n15670) );
  NAND2_X1 U12017 ( .A1(n12402), .A2(n20150), .ZN(n10109) );
  NOR2_X1 U12018 ( .A1(n14637), .A2(n10127), .ZN(n10126) );
  NOR2_X1 U12019 ( .A1(n14748), .A2(n10120), .ZN(n10119) );
  INV_X1 U12020 ( .A(n14752), .ZN(n10120) );
  OR2_X1 U12021 ( .A1(n13225), .A2(n13240), .ZN(n14937) );
  AND2_X1 U12022 ( .A1(n12631), .A2(n13984), .ZN(n10112) );
  INV_X1 U12023 ( .A(n12525), .ZN(n12909) );
  AND2_X1 U12024 ( .A1(n12607), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12623) );
  AND2_X1 U12025 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n12579), .ZN(
        n12607) );
  NOR2_X1 U12026 ( .A1(n12502), .A2(n12501), .ZN(n13179) );
  NOR2_X1 U12027 ( .A1(n14638), .A2(n10157), .ZN(n10158) );
  AND2_X1 U12028 ( .A1(n14423), .A2(n14422), .ZN(n14714) );
  INV_X1 U12029 ( .A(n13209), .ZN(n10189) );
  INV_X1 U12030 ( .A(n15942), .ZN(n10185) );
  NAND2_X1 U12031 ( .A1(n13209), .A2(n10188), .ZN(n10187) );
  INV_X1 U12032 ( .A(n13202), .ZN(n10188) );
  NOR2_X1 U12033 ( .A1(n12604), .A2(n12633), .ZN(n10192) );
  INV_X1 U12034 ( .A(n14437), .ZN(n14411) );
  AND2_X1 U12035 ( .A1(n10164), .A2(n13840), .ZN(n10163) );
  NAND2_X1 U12036 ( .A1(n14441), .A2(n14404), .ZN(n14431) );
  INV_X1 U12037 ( .A(n13658), .ZN(n10165) );
  OR2_X1 U12038 ( .A1(n13628), .A2(n13627), .ZN(n14957) );
  AND3_X1 U12039 ( .A1(n13535), .A2(n13130), .A3(n13129), .ZN(n13504) );
  OR2_X1 U12040 ( .A1(n13165), .A2(n20139), .ZN(n13199) );
  AOI22_X1 U12041 ( .A1(n12594), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12364), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12336) );
  NAND2_X1 U12042 ( .A1(n13221), .A2(n13108), .ZN(n13109) );
  AOI221_X1 U12043 ( .B1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n13081), 
        .C1(n13738), .C2(n13081), .A(n13077), .ZN(n13138) );
  INV_X1 U12044 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12532) );
  INV_X1 U12045 ( .A(n15712), .ZN(n13759) );
  OR2_X1 U12046 ( .A1(n10730), .A2(n10729), .ZN(n10732) );
  NAND2_X1 U12047 ( .A1(n10083), .A2(n16154), .ZN(n10082) );
  INV_X1 U12048 ( .A(n18858), .ZN(n10083) );
  NAND2_X1 U12049 ( .A1(n10082), .A2(n18858), .ZN(n10081) );
  AND2_X1 U12050 ( .A1(n10850), .A2(n13823), .ZN(n10854) );
  AND2_X1 U12051 ( .A1(n10784), .A2(n10142), .ZN(n10852) );
  NOR2_X1 U12052 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12095) );
  OR2_X1 U12053 ( .A1(n12193), .A2(n11939), .ZN(n11944) );
  BUF_X1 U12054 ( .A(n10347), .Z(n14538) );
  CLKBUF_X1 U12055 ( .A(n14532), .Z(n14543) );
  NOR2_X1 U12056 ( .A1(n12024), .A2(n10209), .ZN(n10208) );
  INV_X1 U12057 ( .A(n14209), .ZN(n10209) );
  NOR2_X1 U12058 ( .A1(n16085), .A2(n10067), .ZN(n10066) );
  NOR2_X1 U12059 ( .A1(n13327), .A2(n10056), .ZN(n10055) );
  INV_X1 U12060 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10056) );
  INV_X1 U12061 ( .A(n10060), .ZN(n10059) );
  NAND2_X1 U12062 ( .A1(n10134), .A2(n10133), .ZN(n10699) );
  NAND2_X1 U12063 ( .A1(n10689), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10133) );
  NAND2_X1 U12064 ( .A1(n10973), .A2(n9827), .ZN(n10134) );
  NOR2_X1 U12065 ( .A1(n10595), .A2(n10137), .ZN(n11245) );
  NOR2_X1 U12066 ( .A1(n11024), .A2(n10284), .ZN(n10282) );
  NOR2_X1 U12067 ( .A1(n10253), .A2(n11845), .ZN(n10251) );
  NOR2_X1 U12068 ( .A1(n15485), .A2(n15484), .ZN(n15283) );
  NAND2_X1 U12069 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n10278) );
  NOR2_X1 U12070 ( .A1(n13958), .A2(n10212), .ZN(n10210) );
  INV_X1 U12071 ( .A(n11018), .ZN(n11021) );
  AND2_X1 U12072 ( .A1(n9883), .A2(n13669), .ZN(n10240) );
  NOR2_X1 U12073 ( .A1(n10960), .A2(n10689), .ZN(n11269) );
  AND3_X1 U12074 ( .A1(n10825), .A2(n10312), .A3(n10824), .ZN(n11265) );
  AND3_X1 U12075 ( .A1(n11053), .A2(n11052), .A3(n11051), .ZN(n13637) );
  OR2_X1 U12076 ( .A1(n10689), .A2(n10781), .ZN(n11261) );
  NAND2_X1 U12077 ( .A1(n11005), .A2(n11004), .ZN(n11008) );
  NAND2_X1 U12078 ( .A1(n10688), .A2(n13856), .ZN(n10702) );
  AND2_X1 U12079 ( .A1(n10649), .A2(n10960), .ZN(n10286) );
  NAND2_X1 U12080 ( .A1(n10492), .A2(n10039), .ZN(n10477) );
  AND4_X1 U12081 ( .A1(n10445), .A2(n11194), .A3(n10425), .A4(n12239), .ZN(
        n10418) );
  NOR2_X1 U12082 ( .A1(n10326), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10540) );
  OR2_X1 U12083 ( .A1(n12193), .A2(n11920), .ZN(n11930) );
  NOR2_X1 U12084 ( .A1(n10502), .A2(n14043), .ZN(n10499) );
  NOR2_X1 U12085 ( .A1(n14598), .A2(n10531), .ZN(n10511) );
  INV_X1 U12086 ( .A(n10523), .ZN(n10527) );
  AOI21_X1 U12087 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n20915), .A(
        n11637), .ZN(n11643) );
  NOR2_X1 U12088 ( .A1(n11752), .A2(n11644), .ZN(n11637) );
  NAND2_X1 U12089 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18392), .ZN(
        n11644) );
  INV_X1 U12090 ( .A(n11543), .ZN(n11550) );
  AND3_X1 U12091 ( .A1(n9889), .A2(n11748), .A3(n18788), .ZN(n15676) );
  NOR2_X1 U12092 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n11618), .ZN(
        n11619) );
  NAND2_X1 U12093 ( .A1(n15682), .A2(n10102), .ZN(n10104) );
  NOR2_X1 U12094 ( .A1(n17465), .A2(n11759), .ZN(n10102) );
  NAND2_X1 U12095 ( .A1(n16388), .A2(n16380), .ZN(n11618) );
  NAND4_X1 U12096 ( .A1(n18754), .A2(n18769), .A3(n18762), .A4(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10288) );
  NAND2_X1 U12097 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14306) );
  NAND2_X1 U12098 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n10168) );
  INV_X1 U12099 ( .A(n11690), .ZN(n10169) );
  NOR2_X1 U12100 ( .A1(n12745), .A2(n14290), .ZN(n12750) );
  INV_X1 U12101 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19900) );
  INV_X1 U12102 ( .A(n15796), .ZN(n19932) );
  NOR2_X1 U12103 ( .A1(n13654), .A2(n13653), .ZN(n13659) );
  INV_X1 U12104 ( .A(n20117), .ZN(n20119) );
  NAND2_X1 U12105 ( .A1(n14391), .A2(n10126), .ZN(n10125) );
  NAND2_X1 U12106 ( .A1(n12974), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12997) );
  AND2_X1 U12107 ( .A1(n12954), .A2(n12953), .ZN(n14711) );
  OR2_X1 U12108 ( .A1(n15779), .A2(n13063), .ZN(n12953) );
  NOR2_X1 U12109 ( .A1(n12884), .A2(n12883), .ZN(n12885) );
  AND2_X1 U12110 ( .A1(n10117), .A2(n14737), .ZN(n10116) );
  NOR2_X1 U12111 ( .A1(n12846), .A2(n15824), .ZN(n12847) );
  NAND2_X1 U12112 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n12847), .ZN(
        n12884) );
  NAND2_X1 U12113 ( .A1(n12827), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12846) );
  OR2_X1 U12114 ( .A1(n12797), .A2(n14687), .ZN(n12798) );
  NOR2_X1 U12115 ( .A1(n20923), .A2(n12798), .ZN(n12827) );
  AND2_X1 U12116 ( .A1(n12767), .A2(n12766), .ZN(n14302) );
  CLKBUF_X1 U12117 ( .A(n14240), .Z(n14241) );
  NOR2_X1 U12118 ( .A1(n12734), .A2(n10123), .ZN(n10122) );
  NOR2_X1 U12119 ( .A1(n9859), .A2(n9919), .ZN(n10123) );
  AND2_X1 U12120 ( .A1(n14279), .A2(n14278), .ZN(n14281) );
  AND2_X1 U12121 ( .A1(n12687), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12688) );
  NOR2_X1 U12122 ( .A1(n12670), .A2(n19900), .ZN(n12687) );
  CLKBUF_X1 U12123 ( .A(n13986), .Z(n13987) );
  NAND2_X1 U12124 ( .A1(n12637), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12656) );
  AND2_X1 U12125 ( .A1(n12623), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12637) );
  NAND2_X1 U12126 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12560) );
  NAND2_X1 U12127 ( .A1(n14738), .A2(n14730), .ZN(n14731) );
  AND2_X1 U12128 ( .A1(n10029), .A2(n13225), .ZN(n10028) );
  OR2_X1 U12129 ( .A1(n13245), .A2(n10033), .ZN(n10029) );
  OAI21_X1 U12130 ( .B1(n13246), .B2(n9944), .A(n15895), .ZN(n14894) );
  AND2_X1 U12131 ( .A1(n21010), .A2(n13248), .ZN(n10005) );
  NOR2_X1 U12132 ( .A1(n14739), .A2(n14742), .ZN(n14738) );
  AND2_X1 U12133 ( .A1(n14769), .A2(n9925), .ZN(n14749) );
  INV_X1 U12134 ( .A(n14750), .ZN(n10145) );
  NAND2_X1 U12135 ( .A1(n14769), .A2(n9863), .ZN(n14754) );
  NAND2_X1 U12136 ( .A1(n14769), .A2(n14762), .ZN(n14763) );
  NAND2_X1 U12137 ( .A1(n14270), .A2(n14254), .ZN(n14770) );
  NAND2_X1 U12138 ( .A1(n15119), .A2(n14936), .ZN(n10001) );
  NOR2_X1 U12139 ( .A1(n14271), .A2(n14284), .ZN(n14270) );
  AND2_X1 U12140 ( .A1(n14013), .A2(n9902), .ZN(n14282) );
  INV_X1 U12141 ( .A(n14276), .ZN(n10148) );
  NAND2_X1 U12142 ( .A1(n14013), .A2(n10149), .ZN(n14275) );
  NAND2_X1 U12143 ( .A1(n14013), .A2(n13997), .ZN(n14061) );
  NAND2_X1 U12144 ( .A1(n13659), .A2(n10163), .ZN(n13841) );
  AND2_X1 U12145 ( .A1(n10161), .A2(n13659), .ZN(n13993) );
  AND2_X1 U12146 ( .A1(n10163), .A2(n10162), .ZN(n10161) );
  INV_X1 U12147 ( .A(n13834), .ZN(n10162) );
  AND2_X1 U12148 ( .A1(n13659), .A2(n10164), .ZN(n13839) );
  NAND2_X1 U12149 ( .A1(n13659), .A2(n13658), .ZN(n13724) );
  OR2_X1 U12150 ( .A1(n13628), .A2(n14606), .ZN(n20104) );
  AND2_X1 U12151 ( .A1(n14958), .A2(n14957), .ZN(n14972) );
  INV_X1 U12152 ( .A(n20104), .ZN(n20078) );
  INV_X1 U12153 ( .A(n14957), .ZN(n15103) );
  NAND2_X1 U12154 ( .A1(n12524), .A2(n20706), .ZN(n12470) );
  CLKBUF_X1 U12155 ( .A(n13739), .Z(n15161) );
  NAND2_X1 U12156 ( .A1(n12488), .A2(n12487), .ZN(n13513) );
  OR2_X1 U12157 ( .A1(n20197), .A2(n13164), .ZN(n20310) );
  INV_X1 U12158 ( .A(n20310), .ZN(n20562) );
  INV_X1 U12159 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20563) );
  INV_X1 U12160 ( .A(n20241), .ZN(n20640) );
  NAND2_X1 U12161 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20172), .ZN(n20158) );
  AND2_X1 U12162 ( .A1(n20197), .A2(n13164), .ZN(n20591) );
  NOR2_X1 U12163 ( .A1(n20121), .A2(n13772), .ZN(n20637) );
  INV_X1 U12164 ( .A(n20158), .ZN(n20163) );
  AND2_X1 U12165 ( .A1(n14599), .A2(n14602), .ZN(n15724) );
  NAND2_X1 U12166 ( .A1(n10136), .A2(n10135), .ZN(n10973) );
  NAND2_X1 U12167 ( .A1(n13299), .A2(n11142), .ZN(n10135) );
  NAND2_X1 U12168 ( .A1(n11245), .A2(n19845), .ZN(n10136) );
  AND2_X1 U12169 ( .A1(n10244), .A2(n12238), .ZN(n10243) );
  NAND2_X1 U12170 ( .A1(n10139), .A2(n9895), .ZN(n16077) );
  INV_X1 U12171 ( .A(n10957), .ZN(n10139) );
  OR2_X1 U12172 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n10943), .ZN(n16088) );
  NAND2_X1 U12173 ( .A1(n10942), .A2(n16088), .ZN(n10965) );
  OR2_X1 U12174 ( .A1(n10927), .A2(n10926), .ZN(n10938) );
  NAND2_X1 U12175 ( .A1(n10919), .A2(n10920), .ZN(n10927) );
  AND2_X1 U12176 ( .A1(n10885), .A2(n9930), .ZN(n10876) );
  AND2_X1 U12177 ( .A1(n10885), .A2(n10882), .ZN(n10896) );
  NAND2_X1 U12178 ( .A1(n10865), .A2(n9860), .ZN(n10880) );
  AND2_X1 U12179 ( .A1(n10865), .A2(n10867), .ZN(n10894) );
  AND3_X1 U12180 ( .A1(n11338), .A2(n11337), .A3(n11336), .ZN(n13676) );
  AND2_X1 U12181 ( .A1(n10220), .A2(n10219), .ZN(n10218) );
  AND2_X1 U12182 ( .A1(n12095), .A2(n10539), .ZN(n12066) );
  NAND2_X1 U12183 ( .A1(n13586), .A2(n13587), .ZN(n13689) );
  AND2_X1 U12184 ( .A1(n15275), .A2(n10244), .ZN(n14505) );
  AOI21_X1 U12185 ( .B1(n15215), .B2(n15218), .A(n12139), .ZN(n12158) );
  NOR2_X1 U12186 ( .A1(n15166), .A2(n9911), .ZN(n15298) );
  INV_X1 U12187 ( .A(n11830), .ZN(n10237) );
  AND2_X1 U12188 ( .A1(n15298), .A2(n15299), .ZN(n15301) );
  NOR2_X1 U12189 ( .A1(n10204), .A2(n15233), .ZN(n10203) );
  INV_X1 U12190 ( .A(n10205), .ZN(n10204) );
  NOR3_X1 U12191 ( .A1(n15166), .A2(n10235), .A3(n15317), .ZN(n15316) );
  AND2_X1 U12192 ( .A1(n11449), .A2(n11448), .ZN(n15167) );
  NOR2_X1 U12193 ( .A1(n15166), .A2(n15167), .ZN(n15324) );
  NAND2_X1 U12194 ( .A1(n13811), .A2(n13812), .ZN(n15610) );
  OAI211_X1 U12195 ( .C1(n11440), .C2(n11227), .A(n11243), .B(n11226), .ZN(
        n13475) );
  AND2_X1 U12196 ( .A1(n19860), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19065) );
  AOI21_X1 U12197 ( .B1(n19063), .B2(n19062), .A(n19061), .ZN(n19100) );
  AND2_X1 U12198 ( .A1(n13285), .A2(n13289), .ZN(n13358) );
  NAND2_X1 U12199 ( .A1(n14487), .A2(n10065), .ZN(n14473) );
  AND2_X1 U12200 ( .A1(n9861), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10065) );
  NAND2_X1 U12201 ( .A1(n14487), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14492) );
  AND3_X1 U12202 ( .A1(n11110), .A2(n11109), .A3(n11108), .ZN(n15206) );
  NAND2_X1 U12203 ( .A1(n14157), .A2(n13315), .ZN(n14232) );
  AND3_X1 U12204 ( .A1(n11088), .A2(n11087), .A3(n11086), .ZN(n14233) );
  AND2_X1 U12205 ( .A1(n15568), .A2(n15557), .ZN(n10285) );
  AND2_X1 U12206 ( .A1(n9854), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10075) );
  NAND2_X1 U12207 ( .A1(n13894), .A2(n10211), .ZN(n13957) );
  AND2_X1 U12208 ( .A1(n13894), .A2(n13893), .ZN(n13912) );
  NOR2_X1 U12209 ( .A1(n10060), .A2(n9920), .ZN(n10057) );
  AND2_X1 U12210 ( .A1(n13729), .A2(n13728), .ZN(n13818) );
  NAND2_X1 U12211 ( .A1(n13818), .A2(n13817), .ZN(n13819) );
  INV_X1 U12212 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n14220) );
  AND2_X1 U12213 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10062) );
  NOR2_X1 U12214 ( .A1(n18964), .A2(n10063), .ZN(n10061) );
  AND3_X1 U12215 ( .A1(n11048), .A2(n11047), .A3(n11046), .ZN(n13643) );
  NAND2_X1 U12216 ( .A1(n11044), .A2(n11043), .ZN(n13644) );
  NAND2_X1 U12217 ( .A1(n10226), .A2(n11049), .ZN(n13646) );
  NOR2_X1 U12218 ( .A1(n10963), .A2(n10962), .ZN(n10964) );
  NAND2_X1 U12219 ( .A1(n10248), .A2(n10247), .ZN(n11844) );
  INV_X1 U12220 ( .A(n10253), .ZN(n10247) );
  NAND2_X1 U12221 ( .A1(n10250), .A2(n10249), .ZN(n10248) );
  INV_X1 U12222 ( .A(n10955), .ZN(n10250) );
  INV_X1 U12223 ( .A(n10936), .ZN(n10262) );
  NAND2_X1 U12224 ( .A1(n15301), .A2(n13343), .ZN(n15485) );
  AND3_X1 U12225 ( .A1(n11107), .A2(n11106), .A3(n11105), .ZN(n15211) );
  NOR2_X1 U12226 ( .A1(n9941), .A2(n11831), .ZN(n9999) );
  AND2_X1 U12227 ( .A1(n9915), .A2(n13342), .ZN(n10213) );
  AND3_X1 U12228 ( .A1(n11099), .A2(n11098), .A3(n11097), .ZN(n15227) );
  NAND2_X1 U12229 ( .A1(n15241), .A2(n9906), .ZN(n15228) );
  AND2_X1 U12230 ( .A1(n15241), .A2(n9915), .ZN(n15229) );
  NAND2_X1 U12231 ( .A1(n10267), .A2(n10266), .ZN(n15398) );
  AND2_X1 U12232 ( .A1(n10904), .A2(n16178), .ZN(n10266) );
  CLKBUF_X1 U12233 ( .A(n15530), .Z(n15531) );
  AOI21_X1 U12234 ( .B1(n15583), .B2(n11806), .A(n11805), .ZN(n15429) );
  AND2_X1 U12235 ( .A1(n11444), .A2(n11443), .ZN(n14133) );
  AND2_X1 U12236 ( .A1(n14156), .A2(n14155), .ZN(n14157) );
  NAND2_X1 U12237 ( .A1(n9972), .A2(n10047), .ZN(n15583) );
  AOI21_X1 U12238 ( .B1(n9851), .B2(n10048), .A(n11804), .ZN(n10047) );
  NAND2_X1 U12239 ( .A1(n11801), .A2(n9851), .ZN(n9972) );
  INV_X1 U12240 ( .A(n15611), .ZN(n10228) );
  NAND2_X1 U12241 ( .A1(n13811), .A2(n9909), .ZN(n14132) );
  NAND2_X1 U12242 ( .A1(n15598), .A2(n15568), .ZN(n15423) );
  NAND2_X1 U12243 ( .A1(n11801), .A2(n10268), .ZN(n10267) );
  AND2_X1 U12244 ( .A1(n9858), .A2(n11802), .ZN(n10268) );
  AND2_X1 U12245 ( .A1(n16195), .A2(n15606), .ZN(n15621) );
  AND2_X1 U12246 ( .A1(n9923), .A2(n10043), .ZN(n10042) );
  NAND2_X1 U12247 ( .A1(n9976), .A2(n9892), .ZN(n9977) );
  AND2_X1 U12248 ( .A1(n10859), .A2(n11037), .ZN(n16191) );
  AND2_X1 U12249 ( .A1(n13674), .A2(n10238), .ZN(n13693) );
  AND2_X1 U12250 ( .A1(n10240), .A2(n10239), .ZN(n10238) );
  INV_X1 U12251 ( .A(n13676), .ZN(n10239) );
  NAND2_X1 U12252 ( .A1(n13693), .A2(n13694), .ZN(n13766) );
  AND2_X1 U12253 ( .A1(n16212), .A2(n16255), .ZN(n16195) );
  NOR2_X1 U12254 ( .A1(n13819), .A2(n13784), .ZN(n13869) );
  AND2_X1 U12255 ( .A1(n13870), .A2(n13869), .ZN(n13894) );
  NAND2_X1 U12256 ( .A1(n13674), .A2(n10240), .ZN(n13675) );
  AND3_X1 U12257 ( .A1(n11296), .A2(n11295), .A3(n11294), .ZN(n13964) );
  AND2_X1 U12258 ( .A1(n13674), .A2(n9883), .ZN(n13962) );
  NAND2_X1 U12259 ( .A1(n13674), .A2(n13673), .ZN(n13963) );
  AND2_X1 U12260 ( .A1(n13696), .A2(n13695), .ZN(n13729) );
  INV_X1 U12261 ( .A(n14022), .ZN(n14189) );
  AND3_X1 U12262 ( .A1(n11056), .A2(n11055), .A3(n11054), .ZN(n13683) );
  NAND2_X1 U12263 ( .A1(n10223), .A2(n10224), .ZN(n10222) );
  INV_X1 U12264 ( .A(n13683), .ZN(n10223) );
  NAND2_X1 U12265 ( .A1(n10226), .A2(n10224), .ZN(n13682) );
  INV_X1 U12266 ( .A(n11015), .ZN(n9997) );
  XNOR2_X1 U12267 ( .A(n10785), .B(n21044), .ZN(n14113) );
  AND2_X1 U12268 ( .A1(n10232), .A2(n14115), .ZN(n10231) );
  NOR2_X1 U12269 ( .A1(n14070), .A2(n10230), .ZN(n14116) );
  NAND2_X1 U12270 ( .A1(n10233), .A2(n10232), .ZN(n10230) );
  XNOR2_X1 U12271 ( .A(n11008), .B(n11007), .ZN(n14018) );
  NAND2_X1 U12272 ( .A1(n15572), .A2(n11211), .ZN(n15604) );
  NAND2_X1 U12273 ( .A1(n11189), .A2(n11194), .ZN(n10468) );
  NAND2_X1 U12274 ( .A1(n11917), .A2(n20990), .ZN(n11936) );
  CLKBUF_X1 U12275 ( .A(n10540), .Z(n14170) );
  INV_X1 U12276 ( .A(n10792), .ZN(n19329) );
  OR2_X1 U12277 ( .A1(n19296), .A2(n19824), .ZN(n19522) );
  INV_X1 U12278 ( .A(n19589), .ZN(n19575) );
  NAND2_X2 U12279 ( .A1(n10345), .A2(n10344), .ZN(n19174) );
  NAND2_X1 U12280 ( .A1(n10362), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10369) );
  NAND4_X1 U12281 ( .A1(n10298), .A2(n10350), .A3(n10349), .A4(n10348), .ZN(
        n10357) );
  NAND2_X1 U12282 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19672), .ZN(n19184) );
  INV_X1 U12283 ( .A(n19203), .ZN(n19195) );
  OR2_X1 U12285 ( .A1(n19449), .A2(n19417), .ZN(n19622) );
  INV_X1 U12286 ( .A(n19516), .ZN(n19675) );
  INV_X1 U12287 ( .A(n19585), .ZN(n19672) );
  OR2_X1 U12288 ( .A1(n19576), .A2(n19621), .ZN(n19159) );
  INV_X1 U12289 ( .A(n19184), .ZN(n19198) );
  AND2_X1 U12290 ( .A1(n11150), .A2(n10986), .ZN(n13353) );
  NOR2_X1 U12291 ( .A1(n18608), .A2(n16505), .ZN(n18630) );
  NOR2_X1 U12292 ( .A1(n16555), .A2(n16853), .ZN(n16545) );
  OR2_X1 U12293 ( .A1(n16618), .A2(n17547), .ZN(n9968) );
  OR2_X1 U12294 ( .A1(n16640), .A2(n16529), .ZN(n9963) );
  NOR2_X1 U12295 ( .A1(n16647), .A2(n17574), .ZN(n16640) );
  NOR2_X1 U12296 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16805), .ZN(n16787) );
  INV_X1 U12297 ( .A(n16842), .ZN(n16887) );
  NOR2_X1 U12298 ( .A1(n16614), .A2(n10174), .ZN(n10173) );
  INV_X1 U12299 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n10174) );
  NAND2_X1 U12300 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17106), .ZN(n15664) );
  NAND2_X1 U12301 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17174), .ZN(n17164) );
  NOR2_X1 U12302 ( .A1(n17391), .A2(n17351), .ZN(n17369) );
  AOI221_X1 U12303 ( .B1(n18796), .B2(n18644), .C1(n17392), .C2(n18644), .A(
        n17391), .ZN(n17393) );
  NOR2_X1 U12304 ( .A1(n16552), .A2(n16517), .ZN(n16360) );
  OR2_X1 U12305 ( .A1(n9961), .A2(n9960), .ZN(n17468) );
  NAND2_X1 U12306 ( .A1(n17532), .A2(n9958), .ZN(n9961) );
  NOR2_X1 U12307 ( .A1(n17506), .A2(n9959), .ZN(n9958) );
  NOR2_X1 U12308 ( .A1(n16375), .A2(n17878), .ZN(n17463) );
  AND3_X1 U12309 ( .A1(n17562), .A2(n10094), .A3(n9870), .ZN(n17510) );
  NAND2_X1 U12310 ( .A1(n17532), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17505) );
  OR2_X1 U12311 ( .A1(n9957), .A2(n9956), .ZN(n17588) );
  NAND2_X1 U12312 ( .A1(n17640), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17618) );
  NOR2_X1 U12313 ( .A1(n17660), .A2(n17662), .ZN(n17640) );
  INV_X1 U12314 ( .A(n17467), .ZN(n17661) );
  NAND2_X1 U12315 ( .A1(n10104), .A2(n10103), .ZN(n15754) );
  INV_X1 U12316 ( .A(n11619), .ZN(n10103) );
  NAND2_X1 U12317 ( .A1(n17747), .A2(n11601), .ZN(n16381) );
  INV_X1 U12318 ( .A(n10094), .ZN(n17517) );
  AND2_X1 U12319 ( .A1(n10308), .A2(n9938), .ZN(n10090) );
  NOR2_X1 U12320 ( .A1(n16383), .A2(n18785), .ZN(n17989) );
  NAND2_X1 U12321 ( .A1(n17678), .A2(n17679), .ZN(n17672) );
  NOR2_X1 U12322 ( .A1(n17736), .A2(n10098), .ZN(n17703) );
  NAND2_X1 U12323 ( .A1(n10101), .A2(n18057), .ZN(n10099) );
  NAND2_X1 U12324 ( .A1(n10107), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10106) );
  INV_X1 U12325 ( .A(n17753), .ZN(n10107) );
  NOR2_X1 U12326 ( .A1(n17760), .A2(n18088), .ZN(n17759) );
  NAND2_X1 U12327 ( .A1(n10097), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10096) );
  NAND2_X1 U12328 ( .A1(n11593), .A2(n10097), .ZN(n10095) );
  NOR2_X1 U12329 ( .A1(n18811), .A2(n14311), .ZN(n18606) );
  NOR2_X1 U12330 ( .A1(n17787), .A2(n17788), .ZN(n17786) );
  NOR2_X1 U12331 ( .A1(n18795), .A2(n18091), .ZN(n18111) );
  INV_X1 U12332 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20915) );
  NOR2_X1 U12333 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18157), .ZN(n18393) );
  INV_X1 U12334 ( .A(n11729), .ZN(n18171) );
  NOR2_X1 U12335 ( .A1(n11682), .A2(n11681), .ZN(n18175) );
  INV_X1 U12336 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15852) );
  INV_X1 U12337 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15860) );
  AND2_X1 U12338 ( .A1(n15796), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19964) );
  NOR2_X1 U12339 ( .A1(n19932), .A2(n19878), .ZN(n19948) );
  AND2_X1 U12340 ( .A1(n13933), .A2(n13926), .ZN(n19960) );
  OR2_X1 U12341 ( .A1(n19928), .A2(n13924), .ZN(n19952) );
  XNOR2_X1 U12342 ( .A(n14447), .B(n14616), .ZN(n14990) );
  INV_X1 U12343 ( .A(n14776), .ZN(n14767) );
  NAND2_X1 U12344 ( .A1(n13564), .A2(n13563), .ZN(n14774) );
  INV_X1 U12345 ( .A(n12509), .ZN(n14452) );
  CLKBUF_X1 U12346 ( .A(n13155), .Z(n14829) );
  INV_X1 U12347 ( .A(n14810), .ZN(n14828) );
  NAND2_X1 U12348 ( .A1(n13144), .A2(n13143), .ZN(n14808) );
  OR2_X1 U12349 ( .A1(n20013), .A2(n13500), .ZN(n13144) );
  OR2_X1 U12350 ( .A1(n20013), .A2(n13613), .ZN(n20064) );
  INV_X1 U12351 ( .A(n14391), .ZN(n14392) );
  OR2_X1 U12352 ( .A1(n14449), .A2(n14450), .ZN(n14451) );
  AND2_X1 U12353 ( .A1(n12976), .A2(n12957), .ZN(n14874) );
  NAND2_X1 U12354 ( .A1(n10111), .A2(n12631), .ZN(n14010) );
  INV_X1 U12355 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13792) );
  AND2_X1 U12356 ( .A1(n15724), .A2(n14611), .ZN(n20072) );
  NAND2_X1 U12357 ( .A1(n10155), .A2(n10152), .ZN(n14619) );
  OAI21_X1 U12358 ( .B1(n14669), .B2(n10153), .A(n14615), .ZN(n10152) );
  XNOR2_X1 U12359 ( .A(n9991), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14989) );
  NAND2_X1 U12360 ( .A1(n14833), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10027) );
  OAI211_X1 U12361 ( .C1(n14870), .C2(n10015), .A(n10013), .B(n10011), .ZN(
        n14998) );
  NAND2_X1 U12362 ( .A1(n10006), .A2(n10016), .ZN(n10015) );
  INV_X1 U12363 ( .A(n14948), .ZN(n10037) );
  OR2_X1 U12364 ( .A1(n13246), .A2(n14909), .ZN(n15087) );
  NAND2_X1 U12365 ( .A1(n9990), .A2(n13230), .ZN(n14204) );
  NAND2_X1 U12366 ( .A1(n15941), .A2(n13202), .ZN(n15938) );
  NOR2_X1 U12367 ( .A1(n15996), .A2(n20100), .ZN(n20089) );
  AND2_X1 U12368 ( .A1(n14972), .A2(n20104), .ZN(n15142) );
  INV_X1 U12369 ( .A(n20105), .ZN(n20087) );
  OR2_X1 U12370 ( .A1(n13628), .A2(n15158), .ZN(n14958) );
  OR2_X1 U12371 ( .A1(n20122), .A2(n13771), .ZN(n20503) );
  OAI21_X1 U12372 ( .B1(n13763), .B2(n16043), .A(n20284), .ZN(n20115) );
  NAND2_X1 U12373 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n14599), .ZN(n20794) );
  OAI221_X1 U12374 ( .B1(n10300), .B2(n20537), .C1(n10300), .C2(n20285), .A(
        n20599), .ZN(n20302) );
  INV_X1 U12375 ( .A(n20275), .ZN(n20301) );
  OAI211_X1 U12376 ( .C1(n10305), .C2(n20537), .A(n20456), .B(n20403), .ZN(
        n20420) );
  INV_X1 U12377 ( .A(n20384), .ZN(n20419) );
  OAI211_X1 U12378 ( .C1(n20628), .C2(n20600), .A(n20599), .B(n20598), .ZN(
        n20632) );
  INV_X1 U12379 ( .A(n20448), .ZN(n20650) );
  AND2_X1 U12380 ( .A1(n12396), .A2(n20163), .ZN(n20664) );
  AND2_X1 U12381 ( .A1(n20146), .A2(n20163), .ZN(n20670) );
  AND2_X1 U12382 ( .A1(n20154), .A2(n20163), .ZN(n20682) );
  INV_X1 U12383 ( .A(n20483), .ZN(n20688) );
  AND2_X1 U12384 ( .A1(n12509), .A2(n20163), .ZN(n20695) );
  INV_X1 U12385 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20706) );
  INV_X2 U12386 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20708) );
  INV_X1 U12387 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n18818) );
  OAI22_X1 U12388 ( .A1(n16127), .A2(n10068), .B1(n18954), .B2(n16112), .ZN(
        n16110) );
  NAND2_X1 U12389 ( .A1(n10069), .A2(n15381), .ZN(n10068) );
  INV_X1 U12390 ( .A(n16112), .ZN(n10069) );
  AND2_X1 U12391 ( .A1(n10071), .A2(n18954), .ZN(n16111) );
  INV_X1 U12392 ( .A(n10071), .ZN(n16126) );
  AND2_X1 U12393 ( .A1(n16048), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n18928) );
  AND2_X1 U12394 ( .A1(n10085), .A2(n18954), .ZN(n18857) );
  NOR2_X1 U12395 ( .A1(n18966), .A2(n13323), .ZN(n15169) );
  NAND2_X1 U12396 ( .A1(n10784), .A2(n9881), .ZN(n10843) );
  CLKBUF_X1 U12397 ( .A(n13293), .Z(n18954) );
  INV_X1 U12398 ( .A(n18990), .ZN(n18968) );
  INV_X1 U12399 ( .A(n18978), .ZN(n18950) );
  AND2_X1 U12400 ( .A1(n19854), .A2(n13300), .ZN(n18984) );
  OR2_X1 U12401 ( .A1(n18993), .A2(n20990), .ZN(n18990) );
  XNOR2_X1 U12402 ( .A(n14478), .B(n11850), .ZN(n14564) );
  AND3_X1 U12403 ( .A1(n11418), .A2(n11417), .A3(n11416), .ZN(n13956) );
  NAND2_X1 U12404 ( .A1(n10200), .A2(n10315), .ZN(n13915) );
  CLKBUF_X1 U12405 ( .A(n13865), .Z(n13866) );
  OR2_X1 U12406 ( .A1(n11311), .A2(n11310), .ZN(n13814) );
  NOR2_X1 U12407 ( .A1(n13670), .A2(n19156), .ZN(n18999) );
  AOI21_X1 U12408 ( .B1(n13383), .B2(n12236), .A(n16341), .ZN(n15340) );
  INV_X1 U12409 ( .A(n15340), .ZN(n19050) );
  AND2_X1 U12410 ( .A1(n19033), .A2(n12237), .ZN(n19051) );
  AND2_X1 U12411 ( .A1(n13359), .A2(n19169), .ZN(n19132) );
  INV_X1 U12412 ( .A(n19157), .ZN(n19146) );
  NAND2_X1 U12413 ( .A1(n14478), .A2(n14477), .ZN(n16059) );
  NAND2_X1 U12414 ( .A1(n10252), .A2(n10249), .ZN(n14471) );
  NAND2_X1 U12415 ( .A1(n10955), .A2(n10255), .ZN(n10252) );
  OR2_X1 U12416 ( .A1(n11882), .A2(n15191), .ZN(n16094) );
  NAND2_X1 U12417 ( .A1(n10263), .A2(n10936), .ZN(n15369) );
  NAND2_X1 U12418 ( .A1(n10050), .A2(n10051), .ZN(n15409) );
  NAND2_X1 U12419 ( .A1(n10046), .A2(n9851), .ZN(n15601) );
  NAND2_X1 U12420 ( .A1(n11801), .A2(n11802), .ZN(n16179) );
  AND2_X1 U12421 ( .A1(n10260), .A2(n10261), .ZN(n15630) );
  NOR2_X1 U12422 ( .A1(n14182), .A2(n14189), .ZN(n16288) );
  NOR2_X1 U12423 ( .A1(n14070), .A2(n11250), .ZN(n13852) );
  AND2_X1 U12424 ( .A1(n11006), .A2(n10649), .ZN(n13885) );
  INV_X1 U12425 ( .A(n15604), .ZN(n15575) );
  NAND2_X1 U12426 ( .A1(n10496), .A2(n10495), .ZN(n10497) );
  INV_X1 U12427 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19841) );
  NAND2_X1 U12428 ( .A1(n13583), .A2(n13582), .ZN(n19837) );
  INV_X1 U12429 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19831) );
  INV_X1 U12430 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19822) );
  INV_X1 U12431 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16325) );
  NAND2_X1 U12432 ( .A1(n13575), .A2(n13574), .ZN(n19826) );
  INV_X1 U12433 ( .A(n19293), .ZN(n19281) );
  AND2_X1 U12434 ( .A1(n19395), .A2(n19517), .ZN(n19319) );
  INV_X1 U12435 ( .A(n19343), .ZN(n19353) );
  OAI21_X1 U12436 ( .B1(n19379), .B2(n20990), .A(n19363), .ZN(n19382) );
  AND2_X1 U12437 ( .A1(n19395), .A2(n19589), .ZN(n19381) );
  NOR2_X1 U12438 ( .A1(n19621), .A2(n19356), .ZN(n19404) );
  INV_X1 U12439 ( .A(n19444), .ZN(n19440) );
  AND2_X1 U12440 ( .A1(n19395), .A2(n19811), .ZN(n19444) );
  OAI22_X1 U12441 ( .A1(n19488), .A2(n19487), .B1(n19486), .B2(n21095), .ZN(
        n19506) );
  OAI22_X1 U12442 ( .A1(n19197), .A2(n19202), .B1(n20974), .B2(n19195), .ZN(
        n19615) );
  INV_X1 U12443 ( .A(n19680), .ZN(n19625) );
  INV_X1 U12444 ( .A(n19662), .ZN(n19647) );
  OAI21_X1 U12445 ( .B1(n19635), .B2(n19634), .A(n19633), .ZN(n19658) );
  INV_X1 U12446 ( .A(n19638), .ZN(n19677) );
  AND2_X1 U12447 ( .A1(n19169), .A2(n19198), .ZN(n19681) );
  INV_X1 U12448 ( .A(n19600), .ZN(n19689) );
  AND2_X1 U12449 ( .A1(n19180), .A2(n19198), .ZN(n19693) );
  AND2_X1 U12450 ( .A1(n9827), .A2(n19198), .ZN(n19705) );
  INV_X1 U12451 ( .A(n19612), .ZN(n19713) );
  OR2_X1 U12452 ( .A1(n19622), .A2(n19621), .ZN(n19726) );
  INV_X1 U12453 ( .A(n19620), .ZN(n19721) );
  INV_X1 U12454 ( .A(n19159), .ZN(n19722) );
  NOR2_X1 U12455 ( .A1(n11153), .A2(n20990), .ZN(n16334) );
  INV_X1 U12456 ( .A(n16313), .ZN(n11153) );
  NAND2_X1 U12457 ( .A1(n18643), .A2(n18631), .ZN(n17391) );
  OR2_X1 U12458 ( .A1(n11739), .A2(n11740), .ZN(n18811) );
  INV_X1 U12459 ( .A(n9971), .ZN(n16556) );
  INV_X1 U12460 ( .A(n9970), .ZN(n16577) );
  NOR2_X1 U12461 ( .A1(n16585), .A2(n16586), .ZN(n16584) );
  NAND2_X1 U12462 ( .A1(n9967), .A2(n9965), .ZN(n16609) );
  NAND2_X1 U12463 ( .A1(n16853), .A2(n9966), .ZN(n9965) );
  OR2_X1 U12464 ( .A1(n16618), .A2(n9921), .ZN(n9967) );
  INV_X1 U12465 ( .A(n17533), .ZN(n9966) );
  AND2_X1 U12466 ( .A1(n9968), .A2(n16837), .ZN(n16610) );
  INV_X1 U12467 ( .A(n9963), .ZN(n16630) );
  INV_X1 U12468 ( .A(n16895), .ZN(n16886) );
  AND2_X1 U12469 ( .A1(n17545), .A2(n16686), .ZN(n9964) );
  NOR2_X1 U12470 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16830), .ZN(n16817) );
  INV_X1 U12471 ( .A(n16893), .ZN(n16864) );
  AOI211_X1 U12472 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18795), .A(n16509), .B(
        n16508), .ZN(n16896) );
  NAND3_X1 U12473 ( .A1(n16850), .A2(n16846), .A3(n18649), .ZN(n16897) );
  AND2_X1 U12474 ( .A1(n16960), .A2(n9873), .ZN(n16952) );
  NOR2_X1 U12475 ( .A1(n17050), .A2(n10176), .ZN(n17023) );
  AOI211_X1 U12476 ( .C1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .C2(n9834), .A(
        n11710), .B(n11709), .ZN(n11711) );
  NAND2_X1 U12477 ( .A1(n17065), .A2(P3_EBX_REG_15__SCAN_IN), .ZN(n17050) );
  NAND2_X1 U12478 ( .A1(n17136), .A2(P3_EBX_REG_10__SCAN_IN), .ZN(n17119) );
  NOR2_X1 U12479 ( .A1(n17157), .A2(n16775), .ZN(n17136) );
  NAND2_X1 U12480 ( .A1(n17163), .A2(P3_EBX_REG_8__SCAN_IN), .ZN(n17157) );
  NOR2_X1 U12481 ( .A1(n17164), .A2(n10175), .ZN(n17163) );
  NAND2_X1 U12482 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_7__SCAN_IN), 
        .ZN(n10175) );
  AND2_X1 U12483 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n17176), .ZN(n17171) );
  AND2_X1 U12484 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17171), .ZN(n17174) );
  AND2_X1 U12485 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n17181), .ZN(n17176) );
  INV_X2 U12486 ( .A(n17160), .ZN(n18188) );
  AND3_X1 U12487 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(n17190), .ZN(n17181) );
  NAND2_X1 U12488 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17226), .ZN(n17222) );
  INV_X1 U12489 ( .A(n17281), .ZN(n17268) );
  OR2_X1 U12490 ( .A1(n17397), .A2(n17269), .ZN(n17270) );
  NOR2_X1 U12491 ( .A1(n18188), .A2(n17344), .ZN(n17319) );
  NOR2_X1 U12492 ( .A1(n11518), .A2(n11517), .ZN(n17327) );
  INV_X1 U12493 ( .A(n17319), .ZN(n17339) );
  INV_X1 U12494 ( .A(n17345), .ZN(n17343) );
  NOR2_X1 U12495 ( .A1(n11540), .A2(n11539), .ZN(n11589) );
  NAND2_X1 U12496 ( .A1(n18616), .A2(n17195), .ZN(n17350) );
  NOR2_X1 U12497 ( .A1(n17339), .A2(n18616), .ZN(n17345) );
  CLKBUF_X1 U12498 ( .A(n17379), .Z(n17386) );
  NAND2_X1 U12500 ( .A1(n10100), .A2(n9935), .ZN(n17722) );
  INV_X1 U12501 ( .A(n17736), .ZN(n10100) );
  NAND2_X1 U12502 ( .A1(n9848), .A2(n16383), .ZN(n17726) );
  INV_X1 U12503 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17757) );
  NOR2_X1 U12504 ( .A1(n17775), .A2(n17777), .ZN(n17758) );
  INV_X1 U12505 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17777) );
  NAND2_X1 U12506 ( .A1(n18393), .A2(n18211), .ZN(n18499) );
  INV_X1 U12507 ( .A(n17822), .ZN(n17806) );
  NAND2_X1 U12508 ( .A1(n17817), .A2(n17715), .ZN(n17804) );
  NAND2_X1 U12509 ( .A1(n17562), .A2(n11613), .ZN(n17529) );
  NOR2_X1 U12510 ( .A1(n18606), .A2(n18615), .ZN(n18129) );
  INV_X1 U12511 ( .A(n17989), .ZN(n18010) );
  INV_X1 U12512 ( .A(n18121), .ZN(n18130) );
  INV_X1 U12513 ( .A(n18138), .ZN(n18140) );
  AOI21_X2 U12514 ( .B1(n11902), .B2(n11901), .A(n18651), .ZN(n18136) );
  INV_X1 U12515 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18392) );
  INV_X1 U12516 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18626) );
  INV_X1 U12517 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18154) );
  AOI211_X1 U12518 ( .C1(n18643), .C2(n18613), .A(n18159), .B(n15677), .ZN(
        n18775) );
  INV_X1 U12519 ( .A(n17193), .ZN(n18182) );
  AND2_X1 U12520 ( .A1(n13154), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20117)
         );
  INV_X1 U12521 ( .A(n19158), .ZN(n19156) );
  OAI21_X1 U12522 ( .B1(n15021), .B2(n20105), .A(n10193), .ZN(P1_U3004) );
  NOR2_X1 U12523 ( .A1(n15022), .A2(n10194), .ZN(n10193) );
  NOR2_X1 U12524 ( .A1(n15007), .A2(n14853), .ZN(n10194) );
  AOI21_X1 U12525 ( .B1(n16069), .B2(n16068), .A(n16067), .ZN(n16070) );
  NOR2_X1 U12526 ( .A1(n13865), .A2(n10201), .ZN(n14080) );
  NAND2_X1 U12527 ( .A1(n10197), .A2(n10196), .ZN(n13590) );
  NAND2_X1 U12528 ( .A1(n14598), .A2(n15201), .ZN(n10197) );
  OR2_X1 U12529 ( .A1(n15201), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10196) );
  INV_X1 U12530 ( .A(n11156), .ZN(n11157) );
  NAND2_X1 U12531 ( .A1(n11891), .A2(n16228), .ZN(n11892) );
  INV_X1 U12532 ( .A(n11860), .ZN(n11861) );
  AOI21_X1 U12533 ( .B1(n14517), .B2(n14516), .A(n14515), .ZN(n14518) );
  NAND2_X1 U12534 ( .A1(n14514), .A2(n14513), .ZN(n14515) );
  AND2_X1 U12535 ( .A1(n14502), .A2(n11843), .ZN(n14517) );
  AOI21_X1 U12536 ( .B1(n10023), .B2(n15577), .A(n10020), .ZN(n15581) );
  OAI21_X1 U12537 ( .B1(n15579), .B2(n16271), .A(n10021), .ZN(n10020) );
  NAND2_X1 U12538 ( .A1(n14588), .A2(n10198), .ZN(P2_U3044) );
  OR2_X1 U12539 ( .A1(n16272), .A2(n14598), .ZN(n10198) );
  NOR4_X1 U12540 ( .A1(n9948), .A2(n16538), .A3(n16537), .A4(n9947), .ZN(n9946) );
  NAND2_X1 U12541 ( .A1(n9950), .A2(n16874), .ZN(n9949) );
  NOR2_X1 U12542 ( .A1(n16542), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n9948) );
  NOR2_X1 U12543 ( .A1(n14306), .A2(n11499), .ZN(n11655) );
  INV_X1 U12544 ( .A(n13565), .ZN(n14615) );
  NAND2_X1 U12545 ( .A1(n14680), .A2(n14752), .ZN(n14747) );
  NAND2_X1 U12546 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13277) );
  NAND2_X1 U12547 ( .A1(n12686), .A2(n9859), .ZN(n14265) );
  AND2_X1 U12548 ( .A1(n15074), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9849) );
  NAND2_X1 U12549 ( .A1(n14128), .A2(n14209), .ZN(n14208) );
  INV_X1 U12550 ( .A(n11716), .ZN(n17004) );
  OR2_X1 U12551 ( .A1(n14306), .A2(n16880), .ZN(n9850) );
  OR2_X1 U12552 ( .A1(n10322), .A2(n15619), .ZN(n9851) );
  NAND2_X1 U12553 ( .A1(n11026), .A2(n10307), .ZN(n13272) );
  AND2_X1 U12554 ( .A1(n14680), .A2(n10117), .ZN(n14736) );
  NAND2_X1 U12555 ( .A1(n12686), .A2(n12685), .ZN(n14139) );
  NAND2_X1 U12556 ( .A1(n10000), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11817) );
  AND3_X1 U12557 ( .A1(n10064), .A2(n10061), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n9852) );
  AND2_X1 U12558 ( .A1(n16960), .A2(P3_EBX_REG_22__SCAN_IN), .ZN(n9853) );
  INV_X1 U12559 ( .A(n11544), .ZN(n17142) );
  NAND2_X1 U12560 ( .A1(n10041), .A2(n10044), .ZN(n10260) );
  AND2_X1 U12561 ( .A1(n10076), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9854) );
  OAI21_X1 U12562 ( .B1(n14218), .B2(n14216), .A(n10845), .ZN(n16223) );
  NOR2_X1 U12563 ( .A1(n16224), .A2(n14217), .ZN(n9855) );
  AND2_X1 U12564 ( .A1(n10233), .A2(n10231), .ZN(n9856) );
  INV_X1 U12565 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13276) );
  INV_X1 U12566 ( .A(n16974), .ZN(n11534) );
  AND2_X1 U12567 ( .A1(n10210), .A2(n13296), .ZN(n9857) );
  AOI21_X1 U12568 ( .B1(n10845), .B2(n14216), .A(n9855), .ZN(n10044) );
  INV_X1 U12569 ( .A(n17724), .ZN(n10101) );
  OR2_X1 U12570 ( .A1(n14051), .A2(n10869), .ZN(n9858) );
  NAND2_X1 U12571 ( .A1(n14128), .A2(n10205), .ZN(n15231) );
  NAND2_X1 U12572 ( .A1(n13270), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13268) );
  NAND2_X1 U12573 ( .A1(n13270), .A2(n9854), .ZN(n13309) );
  NAND2_X1 U12574 ( .A1(n13321), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11822) );
  AND2_X1 U12575 ( .A1(n12685), .A2(n12693), .ZN(n9859) );
  AND2_X1 U12576 ( .A1(n10847), .A2(n11063), .ZN(n16225) );
  AND2_X1 U12577 ( .A1(n9913), .A2(n10871), .ZN(n9860) );
  AND2_X1 U12578 ( .A1(n10066), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9861) );
  AND2_X1 U12579 ( .A1(n10055), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9862) );
  AND2_X1 U12580 ( .A1(n10146), .A2(n14753), .ZN(n9863) );
  AND2_X1 U12581 ( .A1(n17724), .A2(n17947), .ZN(n9864) );
  AND2_X1 U12582 ( .A1(n17678), .A2(n9938), .ZN(n9865) );
  AND2_X1 U12583 ( .A1(n13641), .A2(n11949), .ZN(n9866) );
  AND2_X1 U12584 ( .A1(n9860), .A2(n9933), .ZN(n9867) );
  NAND2_X1 U12585 ( .A1(n14487), .A2(n9861), .ZN(n11886) );
  NAND2_X1 U12586 ( .A1(n13321), .A2(n9862), .ZN(n13335) );
  AND2_X1 U12587 ( .A1(n12157), .A2(n15205), .ZN(n9868) );
  AND2_X1 U12588 ( .A1(n14476), .A2(n11883), .ZN(n9869) );
  AND2_X1 U12589 ( .A1(n11613), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9870) );
  AND2_X1 U12590 ( .A1(n10285), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9871) );
  AND2_X1 U12591 ( .A1(n10173), .A2(P3_EBX_REG_24__SCAN_IN), .ZN(n9872) );
  AND2_X1 U12592 ( .A1(n9872), .A2(P3_EBX_REG_25__SCAN_IN), .ZN(n9873) );
  INV_X2 U12593 ( .A(n19869), .ZN(n19792) );
  INV_X2 U12594 ( .A(n11075), .ZN(n11125) );
  INV_X1 U12595 ( .A(n11233), .ZN(n11355) );
  CLKBUF_X3 U12596 ( .A(n11124), .Z(n11131) );
  XNOR2_X1 U12597 ( .A(n11589), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11774) );
  NOR2_X1 U12598 ( .A1(n17737), .A2(n18071), .ZN(n17736) );
  OR2_X1 U12599 ( .A1(n14653), .A2(n10125), .ZN(n9874) );
  AND2_X1 U12600 ( .A1(n10260), .A2(n10258), .ZN(n15629) );
  OR2_X1 U12601 ( .A1(n11817), .A2(n10278), .ZN(n15376) );
  NAND2_X1 U12602 ( .A1(n15598), .A2(n10285), .ZN(n15424) );
  NAND2_X1 U12603 ( .A1(n10129), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10767) );
  NOR2_X1 U12604 ( .A1(n16609), .A2(n16853), .ZN(n9875) );
  NOR2_X1 U12605 ( .A1(n13277), .A2(n13276), .ZN(n13278) );
  AND2_X1 U12606 ( .A1(n16960), .A2(n9872), .ZN(n9876) );
  AND2_X1 U12607 ( .A1(n16960), .A2(n10173), .ZN(n9877) );
  INV_X1 U12608 ( .A(n13277), .ZN(n10064) );
  NOR2_X1 U12609 ( .A1(n13225), .A2(n16006), .ZN(n9879) );
  INV_X1 U12610 ( .A(n20150), .ZN(n12392) );
  NAND2_X1 U12611 ( .A1(n9976), .A2(n10837), .ZN(n14218) );
  NOR2_X1 U12612 ( .A1(n10262), .A2(n15368), .ZN(n9880) );
  AND2_X1 U12613 ( .A1(n10142), .A2(n10841), .ZN(n9881) );
  NAND2_X1 U12614 ( .A1(n14948), .A2(n13231), .ZN(n14912) );
  XNOR2_X1 U12615 ( .A(n12158), .B(n12157), .ZN(n15204) );
  AND2_X1 U12616 ( .A1(n11748), .A2(n11738), .ZN(n9882) );
  NAND2_X1 U12617 ( .A1(n10933), .A2(n10932), .ZN(n15378) );
  AND2_X1 U12618 ( .A1(n10267), .A2(n16178), .ZN(n15617) );
  AND2_X1 U12619 ( .A1(n10241), .A2(n13673), .ZN(n9883) );
  AND4_X1 U12620 ( .A1(n12330), .A2(n12329), .A3(n12328), .A4(n12327), .ZN(
        n9884) );
  AND4_X1 U12622 ( .A1(n11688), .A2(n11687), .A3(n11686), .A4(n11685), .ZN(
        n9885) );
  AND4_X1 U12623 ( .A1(n10751), .A2(n10750), .A3(n10749), .A4(n10748), .ZN(
        n9886) );
  NOR2_X1 U12624 ( .A1(n16082), .A2(n18966), .ZN(n9887) );
  NOR3_X1 U12625 ( .A1(n14313), .A2(n17160), .A3(n14312), .ZN(n14314) );
  AND2_X1 U12626 ( .A1(n15357), .A2(n9880), .ZN(n9888) );
  AND2_X1 U12627 ( .A1(n11738), .A2(n18587), .ZN(n9889) );
  AND2_X1 U12628 ( .A1(n13299), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9890) );
  NAND2_X1 U12629 ( .A1(n14680), .A2(n10119), .ZN(n10121) );
  AND2_X1 U12630 ( .A1(n15366), .A2(n10954), .ZN(n9891) );
  AND2_X1 U12631 ( .A1(n10837), .A2(n10044), .ZN(n9892) );
  NOR2_X1 U12632 ( .A1(n10086), .A2(n18122), .ZN(n9893) );
  AND2_X1 U12633 ( .A1(n11194), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9894) );
  INV_X2 U12634 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n16293) );
  NAND2_X1 U12635 ( .A1(n16089), .A2(n10948), .ZN(n9895) );
  AND4_X1 U12636 ( .A1(n11695), .A2(n11694), .A3(n11693), .A4(n11692), .ZN(
        n9896) );
  AND4_X1 U12637 ( .A1(n10591), .A2(n10589), .A3(n10590), .A4(n10138), .ZN(
        n9897) );
  NAND2_X1 U12638 ( .A1(n9977), .A2(n10042), .ZN(n16187) );
  INV_X1 U12639 ( .A(n10212), .ZN(n10211) );
  NAND2_X1 U12640 ( .A1(n13893), .A2(n13911), .ZN(n10212) );
  NAND2_X1 U12641 ( .A1(n12483), .A2(n9982), .ZN(n9898) );
  NAND2_X1 U12642 ( .A1(n10263), .A2(n9880), .ZN(n9899) );
  AND2_X1 U12643 ( .A1(n12557), .A2(n10191), .ZN(n9900) );
  NAND2_X1 U12644 ( .A1(n15891), .A2(n10002), .ZN(n10035) );
  INV_X1 U12645 ( .A(n10035), .ZN(n10031) );
  AND2_X1 U12646 ( .A1(n11013), .A2(n11012), .ZN(n9901) );
  AND2_X1 U12647 ( .A1(n10149), .A2(n10148), .ZN(n9902) );
  INV_X1 U12648 ( .A(n10254), .ZN(n10249) );
  NAND2_X1 U12649 ( .A1(n10246), .A2(n9891), .ZN(n10254) );
  NAND2_X1 U12650 ( .A1(n14018), .A2(n14119), .ZN(n14017) );
  AND2_X1 U12651 ( .A1(n11026), .A2(n10057), .ZN(n13269) );
  BUF_X1 U12652 ( .A(n12332), .Z(n13050) );
  NAND2_X1 U12653 ( .A1(n17528), .A2(n17561), .ZN(n17562) );
  AND2_X1 U12654 ( .A1(n14128), .A2(n10208), .ZN(n15236) );
  NOR2_X1 U12655 ( .A1(n13322), .A2(n18865), .ZN(n13321) );
  AND2_X1 U12656 ( .A1(n13269), .A2(n11027), .ZN(n13270) );
  AND2_X1 U12657 ( .A1(n13270), .A2(n10075), .ZN(n13310) );
  AND2_X1 U12658 ( .A1(n11026), .A2(n10059), .ZN(n13273) );
  AND2_X1 U12659 ( .A1(n13270), .A2(n10076), .ZN(n9903) );
  NAND2_X1 U12660 ( .A1(n10784), .A2(n10783), .ZN(n9904) );
  AND2_X1 U12661 ( .A1(n13894), .A2(n10210), .ZN(n9905) );
  AND2_X1 U12662 ( .A1(n15242), .A2(n11819), .ZN(n9906) );
  NAND2_X1 U12663 ( .A1(n15241), .A2(n15242), .ZN(n9907) );
  AND2_X1 U12664 ( .A1(n10228), .A2(n13812), .ZN(n9908) );
  AND2_X1 U12665 ( .A1(n9908), .A2(n13303), .ZN(n9909) );
  OR2_X1 U12666 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n10910), .ZN(
        n9910) );
  OR3_X1 U12667 ( .A1(n10235), .A2(n15317), .A3(n10237), .ZN(n9911) );
  AND2_X1 U12668 ( .A1(n14769), .A2(n10146), .ZN(n9912) );
  NAND2_X1 U12669 ( .A1(n14179), .A2(n11017), .ZN(n14212) );
  NAND2_X1 U12670 ( .A1(n14017), .A2(n11010), .ZN(n14107) );
  AND2_X1 U12671 ( .A1(n10893), .A2(n10867), .ZN(n9913) );
  NAND2_X1 U12672 ( .A1(n17608), .A2(n10101), .ZN(n17528) );
  OR2_X1 U12673 ( .A1(n15166), .A2(n10235), .ZN(n9914) );
  INV_X1 U12674 ( .A(n10832), .ZN(n10143) );
  AND2_X1 U12675 ( .A1(n9906), .A2(n10214), .ZN(n9915) );
  AND2_X1 U12676 ( .A1(n13811), .A2(n9908), .ZN(n9916) );
  INV_X1 U12677 ( .A(n12604), .ZN(n12602) );
  AND2_X1 U12678 ( .A1(n14835), .A2(n10016), .ZN(n9917) );
  AND2_X1 U12679 ( .A1(n13225), .A2(n9987), .ZN(n9918) );
  AND2_X1 U12680 ( .A1(n12685), .A2(n12705), .ZN(n9919) );
  OR2_X1 U12681 ( .A1(n16199), .A2(n10058), .ZN(n9920) );
  INV_X1 U12682 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16219) );
  OR2_X1 U12683 ( .A1(n17533), .A2(n17547), .ZN(n9921) );
  OR2_X1 U12684 ( .A1(n14842), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9922) );
  NAND2_X1 U12685 ( .A1(n15222), .A2(n10293), .ZN(n15215) );
  NAND2_X1 U12686 ( .A1(n12402), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12748) );
  AND2_X1 U12687 ( .A1(n10258), .A2(n16203), .ZN(n9923) );
  AND2_X1 U12688 ( .A1(n10051), .A2(n10049), .ZN(n9924) );
  AND2_X1 U12689 ( .A1(n9863), .A2(n10145), .ZN(n9925) );
  AND2_X1 U12690 ( .A1(n9909), .A2(n10227), .ZN(n9926) );
  INV_X1 U12691 ( .A(n13875), .ZN(n12631) );
  AOI21_X1 U12692 ( .B1(n13203), .B2(n12760), .A(n12630), .ZN(n13875) );
  INV_X1 U12693 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18964) );
  AND2_X1 U12694 ( .A1(n11947), .A2(n11948), .ZN(n9927) );
  INV_X1 U12695 ( .A(n17188), .ZN(n17184) );
  INV_X1 U12696 ( .A(n12508), .ZN(n13063) );
  NOR2_X1 U12697 ( .A1(n20128), .A2(n20397), .ZN(n9928) );
  NAND2_X1 U12698 ( .A1(n10229), .A2(n10233), .ZN(n13853) );
  AND2_X1 U12699 ( .A1(n13321), .A2(n10054), .ZN(n13334) );
  AND2_X1 U12700 ( .A1(n14013), .A2(n10150), .ZN(n9929) );
  AND2_X1 U12701 ( .A1(n10882), .A2(n10874), .ZN(n9930) );
  OR2_X1 U12702 ( .A1(n12157), .A2(n15205), .ZN(n9931) );
  NAND2_X1 U12703 ( .A1(n13375), .A2(n20139), .ZN(n13139) );
  INV_X1 U12704 ( .A(n14456), .ZN(n10157) );
  NOR2_X1 U12705 ( .A1(n14486), .A2(n14488), .ZN(n14487) );
  NAND2_X1 U12706 ( .A1(n10080), .A2(n10078), .ZN(n18856) );
  OR2_X1 U12707 ( .A1(n10528), .A2(n10527), .ZN(n19451) );
  OR2_X1 U12708 ( .A1(n9827), .A2(n10873), .ZN(n9933) );
  NOR2_X1 U12709 ( .A1(n17759), .A2(n11600), .ZN(n9934) );
  NOR2_X1 U12710 ( .A1(n11607), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9935) );
  OR2_X1 U12711 ( .A1(n11436), .A2(n11435), .ZN(n14079) );
  INV_X1 U12712 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10058) );
  INV_X1 U12713 ( .A(n10221), .ZN(n10220) );
  NAND2_X1 U12714 ( .A1(n9869), .A2(n11850), .ZN(n10221) );
  AND2_X1 U12715 ( .A1(n13321), .A2(n10055), .ZN(n9936) );
  AND2_X1 U12716 ( .A1(n10725), .A2(n10724), .ZN(n11257) );
  AND2_X1 U12717 ( .A1(n9930), .A2(n15238), .ZN(n9937) );
  INV_X1 U12718 ( .A(n16225), .ZN(n10261) );
  INV_X1 U12719 ( .A(n9850), .ZN(n17054) );
  INV_X1 U12720 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n9959) );
  INV_X1 U12721 ( .A(n17556), .ZN(n9962) );
  AND2_X1 U12722 ( .A1(n17679), .A2(n17991), .ZN(n9938) );
  NOR2_X1 U12723 ( .A1(n17786), .A2(n11593), .ZN(n9939) );
  INV_X1 U12724 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10077) );
  AND2_X1 U12725 ( .A1(n14487), .A2(n10066), .ZN(n9940) );
  INV_X1 U12726 ( .A(n20071), .ZN(n20120) );
  AND2_X1 U12727 ( .A1(n13261), .A2(n20570), .ZN(n20071) );
  INV_X1 U12728 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n10181) );
  INV_X1 U12729 ( .A(n17613), .ZN(n10088) );
  INV_X1 U12730 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10067) );
  OR2_X1 U12731 ( .A1(n10278), .A2(n15482), .ZN(n9941) );
  OR2_X1 U12732 ( .A1(n15009), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9942) );
  OR2_X1 U12733 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n9943) );
  INV_X1 U12734 ( .A(n10179), .ZN(n10178) );
  NAND2_X1 U12735 ( .A1(n14984), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10179) );
  NAND2_X1 U12736 ( .A1(n13247), .A2(n10005), .ZN(n9944) );
  OR2_X1 U12737 ( .A1(n9943), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9945) );
  INV_X1 U12738 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10016) );
  INV_X1 U12739 ( .A(n10284), .ZN(n10283) );
  NAND2_X1 U12740 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10284) );
  AOI22_X2 U12741 ( .A1(DATAI_16_), .A2(n20118), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n20162), .ZN(n20603) );
  AOI22_X2 U12742 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20162), .B1(DATAI_30_), 
        .B2(n20118), .ZN(n20693) );
  AOI22_X2 U12743 ( .A1(DATAI_19_), .A2(n20118), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n20162), .ZN(n20615) );
  NOR3_X4 U12744 ( .A1(n14827), .A2(n14452), .A3(n20154), .ZN(n14830) );
  INV_X1 U12745 ( .A(n14808), .ZN(n14827) );
  AOI22_X2 U12746 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20162), .B1(DATAI_26_), 
        .B2(n20118), .ZN(n20669) );
  NOR2_X2 U12747 ( .A1(n18757), .A2(n18660), .ZN(n16874) );
  NAND2_X1 U12748 ( .A1(n9949), .A2(n9946), .ZN(P3_U2641) );
  INV_X1 U12749 ( .A(n16544), .ZN(n9953) );
  INV_X1 U12750 ( .A(n9957), .ZN(n17602) );
  INV_X1 U12751 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n9956) );
  INV_X1 U12752 ( .A(n9961), .ZN(n17494) );
  INV_X1 U12753 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n9960) );
  INV_X1 U12754 ( .A(n9968), .ZN(n16617) );
  OR2_X2 U12755 ( .A1(n16584), .A2(n16853), .ZN(n9970) );
  OR2_X2 U12756 ( .A1(n16565), .A2(n16853), .ZN(n9971) );
  NAND2_X1 U12757 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n9973) );
  AND2_X4 U12758 ( .A1(n10539), .A2(n16296), .ZN(n10545) );
  AND2_X2 U12759 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10539) );
  AND2_X4 U12760 ( .A1(n10549), .A2(n10469), .ZN(n12225) );
  INV_X1 U12761 ( .A(n16187), .ZN(n10861) );
  INV_X1 U12762 ( .A(n10462), .ZN(n10478) );
  OR2_X2 U12763 ( .A1(n15417), .A2(n15418), .ZN(n9980) );
  NAND2_X1 U12764 ( .A1(n12483), .A2(n12482), .ZN(n12488) );
  XNOR2_X2 U12765 ( .A(n12410), .B(n12479), .ZN(n20238) );
  OAI21_X4 U12766 ( .B1(n13249), .B2(n13225), .A(n9986), .ZN(n14870) );
  NAND2_X2 U12767 ( .A1(n9990), .A2(n9988), .ZN(n14948) );
  NAND4_X1 U12768 ( .A1(n10443), .A2(n9992), .A3(n19860), .A4(n10444), .ZN(
        n10257) );
  NAND2_X1 U12769 ( .A1(n10436), .A2(n10437), .ZN(n9992) );
  NAND2_X1 U12770 ( .A1(n11189), .A2(n9992), .ZN(n16308) );
  AOI21_X1 U12771 ( .B1(n10297), .B2(n11014), .A(n9901), .ZN(n9995) );
  NAND2_X1 U12772 ( .A1(n14178), .A2(n10018), .ZN(n10019) );
  NAND3_X1 U12773 ( .A1(n14017), .A2(n10276), .A3(n9997), .ZN(n9996) );
  NAND2_X1 U12774 ( .A1(n15598), .A2(n9871), .ZN(n15530) );
  NAND2_X2 U12775 ( .A1(n11023), .A2(n11022), .ZN(n15598) );
  NOR2_X4 U12776 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13740) );
  NOR2_X1 U12777 ( .A1(n10001), .A2(n14939), .ZN(n14924) );
  NOR2_X1 U12778 ( .A1(n15895), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10004) );
  NAND2_X2 U12779 ( .A1(n14894), .A2(n14878), .ZN(n15050) );
  NAND3_X1 U12780 ( .A1(n10008), .A2(n10007), .A3(n10009), .ZN(n10013) );
  OR2_X1 U12781 ( .A1(n14834), .A2(n10010), .ZN(n10007) );
  NAND2_X1 U12782 ( .A1(n14870), .A2(n10178), .ZN(n13250) );
  NAND2_X1 U12783 ( .A1(n14870), .A2(n10012), .ZN(n10011) );
  NAND2_X1 U12784 ( .A1(n16221), .A2(n16222), .ZN(n11023) );
  NAND3_X1 U12785 ( .A1(n15694), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n10024), .ZN(n10023) );
  NAND2_X2 U12786 ( .A1(n13487), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13486) );
  NAND2_X1 U12787 ( .A1(n15932), .A2(n15930), .ZN(n10026) );
  NAND2_X1 U12788 ( .A1(n10030), .A2(n10028), .ZN(n14895) );
  NAND3_X1 U12789 ( .A1(n14948), .A2(n10032), .A3(n10031), .ZN(n10030) );
  NAND2_X1 U12790 ( .A1(n14948), .A2(n10031), .ZN(n10038) );
  NAND2_X1 U12791 ( .A1(n10035), .A2(n13245), .ZN(n10034) );
  NAND2_X1 U12792 ( .A1(n10037), .A2(n13245), .ZN(n10036) );
  NAND3_X1 U12793 ( .A1(n10036), .A2(n14909), .A3(n10034), .ZN(n14902) );
  NAND2_X4 U12794 ( .A1(n10242), .A2(n10040), .ZN(n19169) );
  NAND2_X1 U12795 ( .A1(n10417), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10040) );
  AND2_X2 U12796 ( .A1(n10468), .A2(n11207), .ZN(n14089) );
  NAND2_X1 U12797 ( .A1(n10045), .A2(n10786), .ZN(n14180) );
  NAND2_X1 U12798 ( .A1(n15416), .A2(n10053), .ZN(n10050) );
  NAND3_X1 U12799 ( .A1(n11026), .A2(n10059), .A3(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n13271) );
  INV_X1 U12800 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10063) );
  NAND4_X1 U12801 ( .A1(n10064), .A2(n10062), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A4(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n13274) );
  NAND3_X1 U12802 ( .A1(n10064), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13275) );
  OAI21_X1 U12803 ( .B1(n16083), .B2(n10073), .A(n10072), .ZN(n16074) );
  NAND2_X1 U12804 ( .A1(n18966), .A2(n14485), .ZN(n10072) );
  INV_X1 U12805 ( .A(n16084), .ZN(n10074) );
  NOR2_X1 U12806 ( .A1(n16083), .A2(n16084), .ZN(n16082) );
  NAND2_X1 U12807 ( .A1(n18966), .A2(n10081), .ZN(n10080) );
  INV_X1 U12808 ( .A(n10085), .ZN(n15168) );
  XNOR2_X1 U12809 ( .A(n10086), .B(n18122), .ZN(n17798) );
  NAND2_X1 U12810 ( .A1(n17678), .A2(n10090), .ZN(n17614) );
  NOR2_X1 U12811 ( .A1(n17510), .A2(n10101), .ZN(n11615) );
  NAND2_X1 U12812 ( .A1(n17528), .A2(n11612), .ZN(n17518) );
  INV_X1 U12813 ( .A(n17773), .ZN(n10097) );
  NOR2_X1 U12814 ( .A1(n17736), .A2(n11607), .ZN(n11608) );
  NAND2_X1 U12815 ( .A1(n15682), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15681) );
  INV_X1 U12816 ( .A(n10104), .ZN(n11621) );
  NAND2_X1 U12817 ( .A1(n11600), .A2(n10107), .ZN(n10105) );
  NOR2_X2 U12818 ( .A1(n17752), .A2(n11603), .ZN(n11606) );
  INV_X2 U12819 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18774) );
  NAND2_X2 U12820 ( .A1(n12402), .A2(n13080), .ZN(n12393) );
  NAND3_X1 U12821 ( .A1(n13621), .A2(n13080), .A3(n13141), .ZN(n10110) );
  NAND2_X2 U12822 ( .A1(n12322), .A2(n9878), .ZN(n13080) );
  OR2_X2 U12823 ( .A1(n12343), .A2(n12342), .ZN(n12396) );
  CLKBUF_X1 U12824 ( .A(n10114), .Z(n10111) );
  NAND3_X1 U12825 ( .A1(n10113), .A2(n10111), .A3(n12631), .ZN(n10115) );
  AND3_X2 U12826 ( .A1(n10113), .A2(n10114), .A3(n10112), .ZN(n13986) );
  INV_X1 U12827 ( .A(n10115), .ZN(n13985) );
  INV_X1 U12828 ( .A(n10121), .ZN(n14744) );
  NOR2_X1 U12829 ( .A1(n14653), .A2(n10124), .ZN(n14636) );
  NOR2_X1 U12830 ( .A1(n14653), .A2(n14654), .ZN(n14449) );
  NAND2_X1 U12831 ( .A1(n10129), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12104) );
  NAND2_X1 U12832 ( .A1(n10129), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12097) );
  NAND2_X1 U12833 ( .A1(n10129), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12126) );
  NAND2_X1 U12834 ( .A1(n10129), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n12146) );
  NAND2_X1 U12835 ( .A1(n10129), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n12140) );
  NAND2_X1 U12836 ( .A1(n10129), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12179) );
  NAND2_X1 U12837 ( .A1(n10129), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12185) );
  NAND2_X1 U12838 ( .A1(n10129), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n12202) );
  NAND2_X1 U12839 ( .A1(n10129), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n12209) );
  NAND2_X1 U12840 ( .A1(n10129), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12227) );
  NAND2_X1 U12841 ( .A1(n10129), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n14545) );
  AOI22_X1 U12842 ( .A1(n10557), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10129), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12122) );
  AOI22_X1 U12843 ( .A1(n10557), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10129), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12162) );
  AOI22_X1 U12844 ( .A1(n10557), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10129), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12168) );
  NAND2_X1 U12845 ( .A1(n11184), .A2(n16283), .ZN(n11494) );
  NAND2_X1 U12846 ( .A1(n10251), .A2(n10955), .ZN(n10131) );
  NAND2_X1 U12847 ( .A1(n10251), .A2(n10254), .ZN(n10132) );
  NAND3_X1 U12848 ( .A1(n9897), .A2(n10592), .A3(n10597), .ZN(n10137) );
  NAND2_X1 U12849 ( .A1(n10885), .A2(n9937), .ZN(n10922) );
  NAND2_X1 U12850 ( .A1(n10865), .A2(n9867), .ZN(n10889) );
  NOR2_X2 U12851 ( .A1(n14404), .A2(n13570), .ZN(n14435) );
  INV_X2 U12852 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18754) );
  NAND2_X2 U12853 ( .A1(n9885), .A2(n10166), .ZN(n17193) );
  NAND3_X1 U12854 ( .A1(n11700), .A2(n11699), .A3(n11698), .ZN(n10171) );
  NAND2_X1 U12855 ( .A1(n9889), .A2(n11748), .ZN(n14311) );
  NAND3_X1 U12856 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(P3_EBX_REG_17__SCAN_IN), 
        .A3(P3_EBX_REG_16__SCAN_IN), .ZN(n10176) );
  AND2_X2 U12857 ( .A1(n12266), .A2(n13743), .ZN(n12595) );
  AND2_X1 U12858 ( .A1(n13141), .A2(n12509), .ZN(n12507) );
  AND2_X1 U12859 ( .A1(n12392), .A2(n12509), .ZN(n12399) );
  NAND3_X1 U12860 ( .A1(n12558), .A2(n12760), .A3(n13774), .ZN(n10177) );
  NAND2_X1 U12861 ( .A1(n10177), .A2(n12513), .ZN(n12514) );
  NOR2_X2 U12862 ( .A1(n13249), .A2(n9942), .ZN(n14834) );
  NAND2_X1 U12863 ( .A1(n15943), .A2(n10184), .ZN(n10183) );
  NAND2_X1 U12864 ( .A1(n12556), .A2(n12557), .ZN(n12577) );
  INV_X1 U12865 ( .A(n12576), .ZN(n10191) );
  NAND2_X1 U12866 ( .A1(n12603), .A2(n12602), .ZN(n12632) );
  AND2_X2 U12867 ( .A1(n10466), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10461) );
  AOI21_X2 U12868 ( .B1(n12158), .B2(n9931), .A(n9868), .ZN(n12177) );
  XNOR2_X1 U12869 ( .A(n12177), .B(n10321), .ZN(n15196) );
  AND2_X2 U12870 ( .A1(n14128), .A2(n10203), .ZN(n15232) );
  NAND3_X1 U12871 ( .A1(n11947), .A2(n11948), .A3(n13641), .ZN(n13636) );
  NAND2_X1 U12872 ( .A1(n15241), .A2(n10213), .ZN(n15212) );
  NAND2_X1 U12873 ( .A1(n11882), .A2(n10218), .ZN(n10215) );
  NAND2_X1 U12874 ( .A1(n11882), .A2(n9869), .ZN(n14478) );
  AND2_X1 U12875 ( .A1(n11882), .A2(n11883), .ZN(n14475) );
  INV_X1 U12876 ( .A(n14070), .ZN(n10229) );
  NAND2_X1 U12877 ( .A1(n10229), .A2(n9856), .ZN(n14114) );
  NAND2_X1 U12878 ( .A1(n15275), .A2(n10243), .ZN(n11852) );
  AND2_X1 U12879 ( .A1(n15275), .A2(n15267), .ZN(n14504) );
  INV_X1 U12880 ( .A(n11852), .ZN(n11478) );
  NOR2_X1 U12881 ( .A1(n10245), .A2(n10439), .ZN(n10992) );
  NOR2_X2 U12882 ( .A1(n10245), .A2(n10440), .ZN(n10434) );
  NAND2_X1 U12883 ( .A1(n10257), .A2(n10448), .ZN(n10256) );
  NAND2_X1 U12884 ( .A1(n10269), .A2(n10490), .ZN(n10486) );
  XNOR2_X1 U12885 ( .A(n10491), .B(n10269), .ZN(n10504) );
  NAND2_X1 U12886 ( .A1(n10428), .A2(n10439), .ZN(n10449) );
  NAND2_X1 U12887 ( .A1(n10272), .A2(n10273), .ZN(n10271) );
  NAND2_X1 U12888 ( .A1(n11017), .A2(n10274), .ZN(n10272) );
  NAND2_X1 U12889 ( .A1(n9838), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14179) );
  NAND2_X1 U12890 ( .A1(n14214), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10274) );
  NOR2_X1 U12891 ( .A1(n11817), .A2(n15509), .ZN(n15386) );
  OAI211_X1 U12892 ( .C1(n15360), .C2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n10281), .B(n10279), .ZN(n11186) );
  NAND2_X1 U12893 ( .A1(n15360), .A2(n10283), .ZN(n11890) );
  AND2_X1 U12894 ( .A1(n15360), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15350) );
  NAND3_X1 U12895 ( .A1(n11006), .A2(n13886), .A3(n10649), .ZN(n11005) );
  NAND2_X1 U12896 ( .A1(n10286), .A2(n11006), .ZN(n10688) );
  INV_X1 U12897 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10287) );
  XNOR2_X1 U12898 ( .A(n11932), .B(n11930), .ZN(n13586) );
  NOR2_X1 U12899 ( .A1(n14862), .A2(n14861), .ZN(n14863) );
  OR2_X1 U12900 ( .A1(n14476), .A2(n14475), .ZN(n14477) );
  NAND2_X1 U12901 ( .A1(n15224), .A2(n15223), .ZN(n15222) );
  XNOR2_X1 U12902 ( .A(n11849), .B(n11848), .ZN(n11865) );
  OAI21_X1 U12903 ( .B1(n20121), .B2(n13199), .A(n13176), .ZN(n13701) );
  XNOR2_X1 U12904 ( .A(n12515), .B(n12516), .ZN(n13764) );
  NAND2_X4 U12905 ( .A1(n13224), .A2(n13223), .ZN(n13225) );
  NAND2_X1 U12906 ( .A1(n9898), .A2(n13513), .ZN(n13752) );
  INV_X1 U12907 ( .A(n18979), .ZN(n18958) );
  AND2_X1 U12908 ( .A1(n11818), .A2(n16228), .ZN(n10289) );
  INV_X1 U12909 ( .A(n16228), .ZN(n19140) );
  INV_X1 U12910 ( .A(n19169), .ZN(n10512) );
  OR2_X1 U12911 ( .A1(n11914), .A2(n17979), .ZN(n10290) );
  OR2_X1 U12912 ( .A1(n11914), .A2(n17725), .ZN(n10291) );
  INV_X1 U12913 ( .A(n19418), .ZN(n19474) );
  OR2_X1 U12914 ( .A1(n19356), .A2(n19575), .ZN(n19297) );
  OR2_X1 U12915 ( .A1(n16047), .A2(n19150), .ZN(n10292) );
  AND2_X1 U12916 ( .A1(n11915), .A2(n10290), .ZN(n10294) );
  NOR2_X1 U12917 ( .A1(n11910), .A2(n10317), .ZN(n10295) );
  OR2_X1 U12918 ( .A1(n10101), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10296) );
  AND2_X1 U12919 ( .A1(n11015), .A2(n14109), .ZN(n10297) );
  AND2_X1 U12920 ( .A1(n10346), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10298) );
  NOR2_X1 U12921 ( .A1(n20529), .A2(n20642), .ZN(n10299) );
  NOR2_X1 U12922 ( .A1(n20529), .A2(n20331), .ZN(n10300) );
  NAND2_X1 U12923 ( .A1(n10405), .A2(n10404), .ZN(n10407) );
  AND2_X1 U12924 ( .A1(n11870), .A2(n10292), .ZN(n10301) );
  INV_X1 U12925 ( .A(n11221), .ZN(n11313) );
  AND3_X1 U12926 ( .A1(n10353), .A2(n10352), .A3(n10351), .ZN(n10302) );
  AND2_X1 U12927 ( .A1(n10577), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n10304) );
  NOR2_X1 U12928 ( .A1(n20529), .A2(n20497), .ZN(n10305) );
  AND2_X1 U12929 ( .A1(n14419), .A2(n14418), .ZN(n10306) );
  NOR2_X1 U12930 ( .A1(n11025), .A2(n14220), .ZN(n10307) );
  AND3_X1 U12931 ( .A1(n21186), .A2(n17971), .A3(n17950), .ZN(n10308) );
  NAND2_X1 U12932 ( .A1(n13558), .A2(n13557), .ZN(n13649) );
  INV_X1 U12933 ( .A(n13649), .ZN(n12530) );
  AND2_X1 U12934 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10309) );
  AND4_X1 U12935 ( .A1(n10758), .A2(n10757), .A3(n10756), .A4(n10755), .ZN(
        n10311) );
  OR2_X1 U12936 ( .A1(n19100), .A2(n19856), .ZN(n19094) );
  AND4_X1 U12937 ( .A1(n10820), .A2(n10819), .A3(n10818), .A4(n10817), .ZN(
        n10312) );
  INV_X1 U12938 ( .A(n15637), .ZN(n11843) );
  NAND2_X1 U12939 ( .A1(n17652), .A2(n17817), .ZN(n17603) );
  AND2_X1 U12940 ( .A1(n12086), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10313) );
  AND2_X1 U12941 ( .A1(n10654), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10314) );
  AND2_X1 U12942 ( .A1(n11953), .A2(n11952), .ZN(n10315) );
  INV_X1 U12943 ( .A(n11225), .ZN(n11314) );
  AND2_X1 U12944 ( .A1(n19169), .A2(n20990), .ZN(n11225) );
  INV_X1 U12945 ( .A(n11314), .ZN(n11272) );
  INV_X1 U12946 ( .A(n14301), .ZN(n14760) );
  AND2_X1 U12947 ( .A1(n11762), .A2(n10291), .ZN(n10316) );
  OR2_X1 U12948 ( .A1(n11909), .A2(n11908), .ZN(n10317) );
  OR2_X1 U12949 ( .A1(n11911), .A2(n17822), .ZN(n10318) );
  NOR2_X1 U12950 ( .A1(n11124), .A2(n13589), .ZN(n10319) );
  AND2_X1 U12951 ( .A1(n11031), .A2(n14175), .ZN(n19138) );
  AND2_X1 U12952 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n10320) );
  CLKBUF_X3 U12953 ( .A(n13565), .Z(n14404) );
  INV_X1 U12954 ( .A(n13375), .ZN(n13376) );
  AND2_X1 U12955 ( .A1(n12174), .A2(n12194), .ZN(n10321) );
  AND3_X1 U12956 ( .A1(n11803), .A2(n11802), .A3(n9858), .ZN(n10322) );
  OR2_X1 U12957 ( .A1(n13106), .A2(n13105), .ZN(n13107) );
  OAI22_X1 U12958 ( .A1(n11968), .A2(n10754), .B1(n19154), .B2(n19173), .ZN(
        n10509) );
  OR2_X1 U12959 ( .A1(n12575), .A2(n12574), .ZN(n13195) );
  AND2_X1 U12960 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n19822), .ZN(
        n10675) );
  OR2_X1 U12961 ( .A1(n10509), .A2(n10508), .ZN(n10600) );
  AOI22_X1 U12962 ( .A1(n12094), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10548), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10390) );
  OR2_X1 U12963 ( .A1(n12601), .A2(n12600), .ZN(n13204) );
  INV_X1 U12964 ( .A(n13167), .ZN(n12450) );
  INV_X1 U12965 ( .A(n13136), .ZN(n13115) );
  OAI21_X1 U12966 ( .B1(n10682), .B2(n10675), .A(n10680), .ZN(n10730) );
  INV_X1 U12967 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11933) );
  OR2_X1 U12968 ( .A1(n11131), .A2(n13855), .ZN(n10489) );
  NAND2_X1 U12969 ( .A1(n9886), .A2(n10311), .ZN(n10777) );
  NAND2_X1 U12970 ( .A1(n10983), .A2(n10674), .ZN(n10682) );
  AND2_X1 U12971 ( .A1(n13102), .A2(n13101), .ZN(n13104) );
  INV_X1 U12972 ( .A(n14727), .ZN(n12912) );
  INV_X1 U12973 ( .A(n14141), .ZN(n12685) );
  OR2_X1 U12974 ( .A1(n12622), .A2(n12621), .ZN(n13213) );
  NOR2_X1 U12975 ( .A1(n12509), .A2(n20708), .ZN(n12525) );
  INV_X1 U12976 ( .A(n13199), .ZN(n13221) );
  OR2_X1 U12977 ( .A1(n12436), .A2(n12435), .ZN(n13167) );
  AND4_X1 U12978 ( .A1(n12317), .A2(n12316), .A3(n12315), .A4(n12314), .ZN(
        n12322) );
  OR2_X1 U12979 ( .A1(n11269), .A2(n10838), .ZN(n10841) );
  AOI21_X1 U12980 ( .B1(n11945), .B2(n11941), .A(n11940), .ZN(n11943) );
  OR2_X1 U12981 ( .A1(n12173), .A2(n12175), .ZN(n12194) );
  INV_X1 U12982 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10947) );
  INV_X1 U12983 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10326) );
  AOI22_X1 U12984 ( .A1(n12094), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10548), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10395) );
  AOI22_X1 U12985 ( .A1(n12094), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10553), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10361) );
  AOI21_X1 U12986 ( .B1(n20453), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n13104), .ZN(n13081) );
  NOR2_X1 U12987 ( .A1(n10306), .A2(n14728), .ZN(n14422) );
  NAND2_X1 U12988 ( .A1(n13045), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12376) );
  INV_X1 U12989 ( .A(n12976), .ZN(n12974) );
  INV_X1 U12990 ( .A(n14761), .ZN(n12783) );
  INV_X1 U12991 ( .A(n14274), .ZN(n12705) );
  OR2_X1 U12992 ( .A1(n13225), .A2(n13241), .ZN(n14934) );
  OR2_X1 U12993 ( .A1(n12449), .A2(n12448), .ZN(n13226) );
  INV_X1 U12994 ( .A(n12587), .ZN(n12588) );
  NOR2_X1 U12995 ( .A1(n15892), .A2(n13244), .ZN(n13245) );
  INV_X1 U12996 ( .A(n13108), .ZN(n13116) );
  AND2_X1 U12997 ( .A1(n10732), .A2(n10731), .ZN(n10978) );
  AND2_X1 U12998 ( .A1(n12112), .A2(n12117), .ZN(n12135) );
  INV_X1 U12999 ( .A(n12081), .ZN(n12051) );
  INV_X1 U13000 ( .A(n11050), .ZN(n11075) );
  INV_X1 U13001 ( .A(n14469), .ZN(n10962) );
  AND2_X1 U13002 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n11602), .ZN(
        n11603) );
  INV_X1 U13003 ( .A(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n21009) );
  INV_X1 U13004 ( .A(n12928), .ZN(n12929) );
  NAND2_X1 U13005 ( .A1(n15796), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13929) );
  INV_X1 U13006 ( .A(n12507), .ZN(n13599) );
  OR2_X1 U13007 ( .A1(n13016), .A2(n13015), .ZN(n13256) );
  INV_X1 U13008 ( .A(n12956), .ZN(n12955) );
  NAND2_X1 U13009 ( .A1(n12784), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12797) );
  NOR2_X1 U13010 ( .A1(n12560), .A2(n13792), .ZN(n12579) );
  INV_X1 U13011 ( .A(n12748), .ZN(n12760) );
  NAND2_X1 U13012 ( .A1(n14404), .A2(n14437), .ZN(n14617) );
  OAI211_X1 U13013 ( .C1(n15736), .C2(n20398), .A(n12486), .B(n12485), .ZN(
        n12487) );
  INV_X1 U13014 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20453) );
  AND3_X1 U13015 ( .A1(n11114), .A2(n11113), .A3(n11112), .ZN(n15198) );
  NOR2_X1 U13016 ( .A1(n13679), .A2(n19194), .ZN(n11949) );
  NAND2_X1 U13017 ( .A1(n11873), .A2(n9891), .ZN(n11876) );
  INV_X1 U13018 ( .A(n16191), .ZN(n10860) );
  NOR2_X1 U13019 ( .A1(n16287), .A2(n11482), .ZN(n16254) );
  XNOR2_X1 U13020 ( .A(n11249), .B(n11248), .ZN(n14069) );
  XNOR2_X1 U13021 ( .A(n15648), .B(n11928), .ZN(n13573) );
  OAI21_X1 U13022 ( .B1(n15680), .B2(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n11648), .ZN(n11753) );
  AOI21_X1 U13023 ( .B1(n11643), .B2(n11642), .A(n11641), .ZN(n11754) );
  OAI21_X1 U13024 ( .B1(n11911), .B2(n18144), .A(n10295), .ZN(n11912) );
  INV_X1 U13025 ( .A(n18167), .ZN(n11701) );
  NOR2_X1 U13026 ( .A1(n18178), .A2(n11701), .ZN(n11900) );
  AND2_X1 U13027 ( .A1(n13504), .A2(n13509), .ZN(n14602) );
  AND2_X1 U13028 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n12929), .ZN(
        n12949) );
  INV_X1 U13029 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14290) );
  OR3_X1 U13030 ( .A1(n20816), .A2(n13703), .A3(n13922), .ZN(n15796) );
  INV_X1 U13031 ( .A(n19960), .ZN(n15859) );
  AND2_X1 U13032 ( .A1(n13569), .A2(n13568), .ZN(n13610) );
  NAND2_X1 U13033 ( .A1(n13518), .A2(n13538), .ZN(n13123) );
  INV_X1 U13034 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n20923) );
  NOR2_X1 U13035 ( .A1(n15852), .A2(n12751), .ZN(n12784) );
  OR2_X1 U13036 ( .A1(n12729), .A2(n15860), .ZN(n12745) );
  OR2_X1 U13037 ( .A1(n12656), .A2(n12651), .ZN(n12670) );
  OR2_X1 U13038 ( .A1(n20072), .A2(n13252), .ZN(n14940) );
  NOR2_X1 U13039 ( .A1(n15116), .A2(n20078), .ZN(n15996) );
  XNOR2_X1 U13040 ( .A(n13486), .B(n13171), .ZN(n13632) );
  AND2_X1 U13041 ( .A1(n13512), .A2(n13559), .ZN(n15712) );
  NAND2_X1 U13042 ( .A1(n12558), .A2(n13772), .ZN(n13776) );
  INV_X1 U13043 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20638) );
  AND2_X1 U13044 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20644) );
  AND2_X1 U13045 ( .A1(n19861), .A2(n19858), .ZN(n13379) );
  INV_X1 U13046 ( .A(n13783), .ZN(n11951) );
  AND2_X1 U13047 ( .A1(n12154), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13641) );
  AND3_X1 U13048 ( .A1(n11379), .A2(n11378), .A3(n11377), .ZN(n13767) );
  NAND2_X1 U13049 ( .A1(n15452), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14513) );
  AND2_X1 U13050 ( .A1(n16189), .A2(n16188), .ZN(n11802) );
  AND2_X1 U13051 ( .A1(n11481), .A2(n15604), .ZN(n14022) );
  AND2_X1 U13052 ( .A1(n11206), .A2(n11205), .ZN(n15645) );
  NAND2_X1 U13053 ( .A1(n21095), .A2(n20990), .ZN(n19810) );
  OR2_X1 U13054 ( .A1(n19622), .A2(n19460), .ZN(n19418) );
  AND2_X1 U13055 ( .A1(n19580), .A2(n19579), .ZN(n19587) );
  AND2_X1 U13056 ( .A1(n19296), .A2(n19826), .ZN(n19811) );
  INV_X1 U13057 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n21095) );
  NOR2_X1 U13058 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16700), .ZN(n16684) );
  NOR2_X1 U13059 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16732), .ZN(n16709) );
  NAND2_X1 U13060 ( .A1(n18812), .A2(n17352), .ZN(n16508) );
  AOI21_X1 U13061 ( .B1(n11649), .B2(n11754), .A(n11753), .ZN(n18631) );
  NAND2_X1 U13062 ( .A1(n11792), .A2(n17717), .ZN(n17626) );
  INV_X1 U13063 ( .A(n17655), .ZN(n17667) );
  INV_X1 U13064 ( .A(n17626), .ZN(n18008) );
  AOI22_X1 U13065 ( .A1(n18786), .A2(n11913), .B1(n18788), .B2(n9828), .ZN(
        n11757) );
  OR2_X1 U13066 ( .A1(n17860), .A2(n11611), .ZN(n11612) );
  NOR2_X1 U13067 ( .A1(n11750), .A2(n18600), .ZN(n18593) );
  INV_X1 U13068 ( .A(n11913), .ZN(n18785) );
  NOR3_X1 U13069 ( .A1(n15676), .A2(n15675), .A3(n15674), .ZN(n18633) );
  INV_X1 U13070 ( .A(n19875), .ZN(n14611) );
  NAND2_X1 U13071 ( .A1(n12949), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12956) );
  NOR2_X1 U13072 ( .A1(n20744), .A2(n15862), .ZN(n14684) );
  AND2_X1 U13073 ( .A1(n15796), .A2(n13923), .ZN(n19928) );
  AND2_X1 U13074 ( .A1(n15796), .A2(n13935), .ZN(n19971) );
  OR2_X1 U13075 ( .A1(n13559), .A2(n19875), .ZN(n13564) );
  AND2_X1 U13076 ( .A1(n13520), .A2(n13592), .ZN(n19976) );
  AND2_X1 U13077 ( .A1(n13016), .A2(n12998), .ZN(n14859) );
  NAND2_X1 U13078 ( .A1(n12885), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12928) );
  NAND2_X1 U13079 ( .A1(n12688), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12729) );
  AND2_X1 U13080 ( .A1(n14940), .A2(n13255), .ZN(n15917) );
  INV_X1 U13081 ( .A(n14940), .ZN(n20065) );
  INV_X1 U13082 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13251) );
  INV_X1 U13083 ( .A(n14958), .ZN(n15971) );
  INV_X1 U13084 ( .A(n14972), .ZN(n20096) );
  NOR2_X1 U13085 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13553) );
  OR2_X1 U13086 ( .A1(n20197), .A2(n20123), .ZN(n20276) );
  OAI22_X1 U13087 ( .A1(n20205), .A2(n20204), .B1(n20459), .B2(n20337), .ZN(
        n20229) );
  NAND2_X1 U13088 ( .A1(n20122), .A2(n20121), .ZN(n20239) );
  INV_X1 U13089 ( .A(n20362), .ZN(n20342) );
  AND2_X1 U13090 ( .A1(n20644), .A2(n12533), .ZN(n20391) );
  NOR2_X1 U13091 ( .A1(n13776), .A2(n13775), .ZN(n20374) );
  INV_X1 U13092 ( .A(n20494), .ZN(n20450) );
  OAI22_X1 U13093 ( .A1(n20461), .A2(n20460), .B1(n20459), .B2(n20594), .ZN(
        n20490) );
  INV_X1 U13094 ( .A(n20527), .ZN(n20512) );
  AND2_X1 U13095 ( .A1(n20197), .A2(n20123), .ZN(n20495) );
  AND2_X1 U13096 ( .A1(n20637), .A2(n20528), .ZN(n20587) );
  INV_X1 U13097 ( .A(n20595), .ZN(n20631) );
  INV_X1 U13098 ( .A(n20475), .ZN(n20676) );
  AND2_X1 U13099 ( .A1(n20637), .A2(n20495), .ZN(n20699) );
  AND2_X1 U13100 ( .A1(n20705), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15736) );
  INV_X1 U13101 ( .A(n16046), .ZN(n16068) );
  INV_X1 U13102 ( .A(n18928), .ZN(n18982) );
  AND2_X1 U13103 ( .A1(n13358), .A2(n13288), .ZN(n18978) );
  AND2_X1 U13104 ( .A1(n19854), .A2(n16332), .ZN(n18979) );
  INV_X1 U13105 ( .A(n15261), .ZN(n15247) );
  NOR2_X1 U13106 ( .A1(n13670), .A2(n19158), .ZN(n18998) );
  INV_X1 U13107 ( .A(n16136), .ZN(n19052) );
  CLKBUF_X1 U13108 ( .A(n19087), .Z(n19856) );
  OAI21_X1 U13109 ( .B1(n15239), .B2(n19157), .A(n11824), .ZN(n11825) );
  INV_X1 U13110 ( .A(n19150), .ZN(n16234) );
  AND2_X1 U13111 ( .A1(n13356), .A2(n11029), .ZN(n19137) );
  INV_X1 U13112 ( .A(n19810), .ZN(n19813) );
  XNOR2_X1 U13113 ( .A(n13586), .B(n13588), .ZN(n19296) );
  OAI21_X1 U13114 ( .B1(n19166), .B2(n19165), .A(n19164), .ZN(n19204) );
  NOR2_X2 U13115 ( .A1(n19460), .A2(n19356), .ZN(n19232) );
  AND2_X1 U13116 ( .A1(n19449), .A2(n19417), .ZN(n19395) );
  NAND2_X1 U13117 ( .A1(n19449), .A2(n19837), .ZN(n19356) );
  INV_X1 U13118 ( .A(n19301), .ZN(n19320) );
  INV_X1 U13119 ( .A(n19297), .ZN(n19351) );
  OR2_X1 U13120 ( .A1(n19390), .A2(n19389), .ZN(n19413) );
  OAI21_X1 U13121 ( .B1(n19443), .B2(n19422), .A(n19672), .ZN(n19446) );
  INV_X1 U13122 ( .A(n19465), .ZN(n19479) );
  INV_X1 U13123 ( .A(n19510), .ZN(n19501) );
  AND2_X1 U13124 ( .A1(n19520), .A2(n19514), .ZN(n19538) );
  INV_X1 U13125 ( .A(n19726), .ZN(n19657) );
  INV_X1 U13126 ( .A(n19811), .ZN(n19621) );
  AND3_X1 U13127 ( .A1(n18818), .A2(n19794), .A3(n19748), .ZN(n19861) );
  NOR2_X1 U13128 ( .A1(n18795), .A2(n18160), .ZN(n11739) );
  INV_X1 U13129 ( .A(n16529), .ZN(n16837) );
  AND2_X1 U13130 ( .A1(n16842), .A2(n16514), .ZN(n16569) );
  NOR2_X1 U13131 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16654), .ZN(n16637) );
  NOR2_X1 U13132 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16674), .ZN(n16665) );
  NOR2_X1 U13133 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16756), .ZN(n16738) );
  NOR2_X1 U13134 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16773), .ZN(n16761) );
  NOR2_X1 U13135 ( .A1(n18645), .A2(n16508), .ZN(n16842) );
  INV_X1 U13136 ( .A(n16882), .ZN(n16872) );
  INV_X1 U13137 ( .A(n17214), .ZN(n17209) );
  NOR2_X1 U13138 ( .A1(n17399), .A2(n17270), .ZN(n17263) );
  INV_X1 U13139 ( .A(n17350), .ZN(n17317) );
  NAND2_X1 U13140 ( .A1(n17613), .A2(n17626), .ZN(n17878) );
  NOR2_X2 U13141 ( .A1(n18757), .A2(n17804), .ZN(n17655) );
  NOR2_X1 U13142 ( .A1(n18163), .A2(n16491), .ZN(n17809) );
  NOR2_X1 U13143 ( .A1(n17493), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17492) );
  NOR2_X1 U13144 ( .A1(n18128), .A2(n17887), .ZN(n17919) );
  INV_X1 U13145 ( .A(n18045), .ZN(n18024) );
  NOR2_X1 U13146 ( .A1(n11894), .A2(n18091), .ZN(n11913) );
  NOR2_X1 U13147 ( .A1(n18785), .A2(n18128), .ZN(n18135) );
  INV_X1 U13148 ( .A(n18393), .ZN(n18441) );
  NOR2_X1 U13149 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18748), .ZN(
        n18770) );
  INV_X1 U13150 ( .A(n18299), .ZN(n18290) );
  INV_X1 U13151 ( .A(n18497), .ZN(n18485) );
  OR2_X1 U13152 ( .A1(n20013), .A2(n13374), .ZN(n20011) );
  NAND2_X1 U13153 ( .A1(n20011), .A2(n13456), .ZN(n20816) );
  INV_X1 U13154 ( .A(n19964), .ZN(n19899) );
  OR2_X1 U13155 ( .A1(n14281), .A2(n14280), .ZN(n15914) );
  OR2_X1 U13156 ( .A1(n14827), .A2(n13664), .ZN(n14305) );
  NAND2_X1 U13157 ( .A1(n19976), .A2(n13620), .ZN(n13719) );
  INV_X1 U13158 ( .A(n19976), .ZN(n20007) );
  INV_X1 U13159 ( .A(n13260), .ZN(n13263) );
  OAI21_X1 U13160 ( .B1(n14281), .B2(n14269), .A(n14268), .ZN(n14945) );
  INV_X1 U13161 ( .A(n15917), .ZN(n20076) );
  INV_X1 U13162 ( .A(n20072), .ZN(n19882) );
  OR2_X1 U13163 ( .A1(n13628), .A2(n13616), .ZN(n16014) );
  OR2_X1 U13164 ( .A1(n13628), .A2(n13609), .ZN(n20105) );
  INV_X1 U13165 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20398) );
  INV_X1 U13166 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13738) );
  OR2_X1 U13167 ( .A1(n20239), .A2(n20276), .ZN(n20190) );
  OR2_X1 U13168 ( .A1(n20239), .A2(n20310), .ZN(n20233) );
  OR2_X1 U13169 ( .A1(n20239), .A2(n20198), .ZN(n20269) );
  OR2_X1 U13170 ( .A1(n20239), .A2(n20234), .ZN(n20275) );
  NAND2_X1 U13171 ( .A1(n20374), .A2(n20528), .ZN(n20330) );
  NAND2_X1 U13172 ( .A1(n20374), .A2(n20591), .ZN(n20396) );
  NAND2_X1 U13173 ( .A1(n20496), .A2(n20528), .ZN(n20447) );
  NAND2_X1 U13174 ( .A1(n20496), .A2(n20562), .ZN(n20494) );
  NAND2_X1 U13175 ( .A1(n20496), .A2(n20591), .ZN(n20527) );
  NAND2_X1 U13176 ( .A1(n20496), .A2(n20495), .ZN(n20561) );
  NAND2_X1 U13177 ( .A1(n20637), .A2(n20562), .ZN(n20595) );
  AND2_X1 U13178 ( .A1(n20641), .A2(n20640), .ZN(n20659) );
  NAND2_X1 U13179 ( .A1(n20637), .A2(n20591), .ZN(n20703) );
  INV_X1 U13180 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20705) );
  INV_X1 U13181 ( .A(n20769), .ZN(n20775) );
  OR2_X1 U13182 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n19872), .ZN(n20810) );
  OR2_X1 U13183 ( .A1(n11177), .A2(n10995), .ZN(n13356) );
  OR4_X1 U13184 ( .A1(n16261), .A2(n19854), .A3(n18961), .A4(n16328), .ZN(
        n18938) );
  INV_X1 U13185 ( .A(n18984), .ZN(n18973) );
  INV_X1 U13186 ( .A(n16151), .ZN(n15562) );
  XNOR2_X1 U13187 ( .A(n13687), .B(n13690), .ZN(n19449) );
  NOR2_X1 U13188 ( .A1(n12254), .A2(n12253), .ZN(n12255) );
  NAND2_X1 U13189 ( .A1(n11224), .A2(n19033), .ZN(n16136) );
  INV_X1 U13190 ( .A(n19050), .ZN(n19033) );
  AND2_X1 U13191 ( .A1(n19034), .A2(n16136), .ZN(n19021) );
  AND2_X1 U13192 ( .A1(n16134), .A2(n13670), .ZN(n19057) );
  INV_X1 U13193 ( .A(n19068), .ZN(n19098) );
  INV_X1 U13194 ( .A(n19100), .ZN(n19130) );
  OR2_X1 U13195 ( .A1(n13359), .A2(n13451), .ZN(n13415) );
  NOR2_X1 U13196 ( .A1(n10289), .A2(n11825), .ZN(n11826) );
  INV_X1 U13197 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16163) );
  INV_X1 U13198 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16199) );
  INV_X1 U13199 ( .A(n19137), .ZN(n16243) );
  INV_X1 U13200 ( .A(n11839), .ZN(n11840) );
  NAND2_X1 U13201 ( .A1(n11209), .A2(n11185), .ZN(n15637) );
  INV_X1 U13202 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16316) );
  AOI211_X2 U13203 ( .C1(n19162), .C2(n19165), .A(n19585), .B(n19155), .ZN(
        n19208) );
  NAND2_X1 U13204 ( .A1(n19209), .A2(n19395), .ZN(n19263) );
  OR2_X1 U13205 ( .A1(n19356), .A2(n19522), .ZN(n19293) );
  INV_X1 U13206 ( .A(n19319), .ZN(n19316) );
  AND2_X1 U13207 ( .A1(n19328), .A2(n19327), .ZN(n19343) );
  INV_X1 U13208 ( .A(n19381), .ZN(n19378) );
  INV_X1 U13209 ( .A(n19404), .ZN(n19416) );
  AND2_X1 U13210 ( .A1(n19455), .A2(n19454), .ZN(n19465) );
  OR2_X1 U13211 ( .A1(n19576), .A2(n19460), .ZN(n19510) );
  OR2_X1 U13212 ( .A1(n19622), .A2(n19522), .ZN(n19542) );
  AOI21_X1 U13213 ( .B1(n19549), .B2(n19550), .A(n19548), .ZN(n19574) );
  INV_X1 U13214 ( .A(n19701), .ZN(n19651) );
  OR2_X1 U13215 ( .A1(n19576), .A2(n19575), .ZN(n19662) );
  INV_X1 U13216 ( .A(n19643), .ZN(n19698) );
  INV_X1 U13217 ( .A(n19807), .ZN(n19804) );
  NOR2_X1 U13218 ( .A1(n18630), .A2(n17391), .ZN(n18812) );
  INV_X1 U13219 ( .A(n11794), .ZN(n16491) );
  NAND2_X1 U13220 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n16897), .ZN(n16882) );
  INV_X1 U13221 ( .A(n16896), .ZN(n16893) );
  AND2_X1 U13222 ( .A1(n17190), .A2(n17160), .ZN(n17188) );
  INV_X1 U13223 ( .A(n17188), .ZN(n17178) );
  NOR2_X1 U13224 ( .A1(n11529), .A2(n11528), .ZN(n17334) );
  NOR2_X1 U13225 ( .A1(n18804), .A2(n17369), .ZN(n17379) );
  INV_X1 U13226 ( .A(n17369), .ZN(n17389) );
  NAND2_X1 U13227 ( .A1(n17613), .A2(n17713), .ZN(n17625) );
  NAND2_X1 U13228 ( .A1(n17321), .A2(n9848), .ZN(n17725) );
  NOR2_X1 U13229 ( .A1(n17573), .A2(n17655), .ZN(n17800) );
  OAI21_X2 U13230 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18801), .A(n16491), 
        .ZN(n17817) );
  INV_X1 U13231 ( .A(n18136), .ZN(n18128) );
  NAND3_X1 U13232 ( .A1(n11913), .A2(n18136), .A3(n16383), .ZN(n18045) );
  NAND2_X1 U13233 ( .A1(n18138), .A2(n18128), .ZN(n18121) );
  INV_X1 U13234 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21022) );
  INV_X1 U13235 ( .A(n18534), .ZN(n18474) );
  INV_X1 U13236 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18757) );
  INV_X1 U13237 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18748) );
  INV_X1 U13238 ( .A(n18745), .ZN(n18742) );
  INV_X1 U13239 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18674) );
  NAND2_X1 U13240 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18674), .ZN(n18807) );
  INV_X1 U13241 ( .A(n16445), .ZN(n16442) );
  INV_X1 U13242 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11968) );
  AND2_X4 U13243 ( .A1(n10538), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14532) );
  AOI22_X1 U13244 ( .A1(n10347), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10325) );
  AOI22_X1 U13245 ( .A1(n12225), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10545), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10324) );
  AND2_X2 U13246 ( .A1(n10326), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14169) );
  AND2_X4 U13247 ( .A1(n14169), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10548) );
  AND2_X4 U13248 ( .A1(n10539), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10556) );
  AOI22_X1 U13249 ( .A1(n10548), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10556), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10323) );
  NAND3_X1 U13250 ( .A1(n10325), .A2(n10324), .A3(n10323), .ZN(n10329) );
  AND2_X4 U13251 ( .A1(n14088), .A2(n10469), .ZN(n10553) );
  AND2_X4 U13252 ( .A1(n10540), .A2(n16296), .ZN(n12094) );
  AOI22_X1 U13253 ( .A1(n10553), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n12094), .ZN(n10327) );
  INV_X1 U13254 ( .A(n10327), .ZN(n10328) );
  OAI21_X2 U13255 ( .B1(n10329), .B2(n10328), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10336) );
  AOI22_X1 U13256 ( .A1(n10347), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10333) );
  AOI22_X1 U13257 ( .A1(n12094), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10553), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10332) );
  AOI22_X1 U13258 ( .A1(n12225), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10545), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10331) );
  AOI22_X1 U13259 ( .A1(n10548), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10556), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10330) );
  NAND4_X1 U13260 ( .A1(n10333), .A2(n10332), .A3(n10331), .A4(n10330), .ZN(
        n10334) );
  NAND2_X4 U13261 ( .A1(n10336), .A2(n10335), .ZN(n19199) );
  AOI22_X1 U13262 ( .A1(n12094), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10553), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10339) );
  AOI22_X1 U13263 ( .A1(n10548), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10556), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10338) );
  AOI22_X1 U13264 ( .A1(n10347), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10337) );
  NAND4_X1 U13265 ( .A1(n10303), .A2(n10339), .A3(n10338), .A4(n10337), .ZN(
        n10345) );
  AOI22_X1 U13266 ( .A1(n12094), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10553), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10342) );
  AOI22_X1 U13267 ( .A1(n10548), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10556), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10341) );
  AOI22_X1 U13268 ( .A1(n10347), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10340) );
  NAND4_X1 U13269 ( .A1(n10343), .A2(n10342), .A3(n10341), .A4(n10340), .ZN(
        n10344) );
  AOI22_X1 U13270 ( .A1(n12225), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10545), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10346) );
  AOI22_X1 U13271 ( .A1(n12094), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10553), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10350) );
  AOI22_X1 U13272 ( .A1(n10548), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10556), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10349) );
  AOI22_X1 U13273 ( .A1(n10347), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10348) );
  AOI22_X1 U13274 ( .A1(n10548), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10556), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10353) );
  AOI22_X1 U13275 ( .A1(n12094), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10553), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10355) );
  AOI22_X1 U13276 ( .A1(n10347), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10354) );
  AOI22_X1 U13277 ( .A1(n10347), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10360) );
  AOI22_X1 U13278 ( .A1(n10548), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10556), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10359) );
  AOI22_X1 U13279 ( .A1(n12225), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10545), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10358) );
  NAND4_X1 U13280 ( .A1(n10361), .A2(n10360), .A3(n10359), .A4(n10358), .ZN(
        n10362) );
  AOI22_X1 U13281 ( .A1(n10347), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10365) );
  AOI22_X1 U13282 ( .A1(n10548), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10556), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10364) );
  AOI22_X1 U13283 ( .A1(n12225), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10545), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10363) );
  NAND4_X1 U13284 ( .A1(n10366), .A2(n10365), .A3(n10364), .A4(n10363), .ZN(
        n10367) );
  NAND2_X1 U13285 ( .A1(n10367), .A2(n16293), .ZN(n10368) );
  AOI22_X1 U13286 ( .A1(n10347), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10373) );
  AOI22_X1 U13287 ( .A1(n10548), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10553), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10372) );
  AOI22_X1 U13288 ( .A1(n12094), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10556), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10371) );
  AOI22_X1 U13289 ( .A1(n12225), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10545), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10370) );
  NAND4_X1 U13290 ( .A1(n10373), .A2(n10372), .A3(n10371), .A4(n10370), .ZN(
        n10374) );
  NAND2_X1 U13291 ( .A1(n10374), .A2(n16293), .ZN(n10381) );
  AOI22_X1 U13292 ( .A1(n10548), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10347), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10378) );
  AOI22_X1 U13293 ( .A1(n12094), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10377) );
  AOI22_X1 U13294 ( .A1(n12225), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10545), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10376) );
  AOI22_X1 U13295 ( .A1(n10553), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10556), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10375) );
  NAND4_X1 U13296 ( .A1(n10378), .A2(n10377), .A3(n10376), .A4(n10375), .ZN(
        n10379) );
  NAND2_X1 U13297 ( .A1(n10379), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10380) );
  NAND2_X2 U13298 ( .A1(n10381), .A2(n10380), .ZN(n10425) );
  AOI22_X1 U13299 ( .A1(n12094), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10548), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10385) );
  AOI22_X1 U13300 ( .A1(n10553), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10556), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10384) );
  AOI22_X1 U13301 ( .A1(n10347), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10383) );
  AOI22_X1 U13302 ( .A1(n12225), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10545), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10382) );
  NAND4_X1 U13303 ( .A1(n10385), .A2(n10384), .A3(n10383), .A4(n10382), .ZN(
        n10386) );
  NAND2_X1 U13304 ( .A1(n10386), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10393) );
  AOI22_X1 U13305 ( .A1(n10347), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10556), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10389) );
  AOI22_X1 U13306 ( .A1(n12225), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10545), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10388) );
  AOI22_X1 U13307 ( .A1(n10553), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10387) );
  NAND4_X1 U13308 ( .A1(n10390), .A2(n10389), .A3(n10388), .A4(n10387), .ZN(
        n10391) );
  NAND2_X1 U13309 ( .A1(n10391), .A2(n16293), .ZN(n10392) );
  NAND2_X2 U13310 ( .A1(n10393), .A2(n10392), .ZN(n10672) );
  OR2_X2 U13311 ( .A1(n10425), .A2(n10672), .ZN(n10440) );
  AOI22_X1 U13312 ( .A1(n12225), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10545), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10394) );
  AOI22_X1 U13313 ( .A1(n10347), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10556), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10397) );
  AOI22_X1 U13314 ( .A1(n12093), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10396) );
  NAND4_X1 U13315 ( .A1(n10398), .A2(n10397), .A3(n10396), .A4(n10395), .ZN(
        n10405) );
  AOI22_X1 U13316 ( .A1(n12094), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10347), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10403) );
  AOI22_X1 U13317 ( .A1(n12093), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10402) );
  AOI22_X1 U13318 ( .A1(n10548), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12225), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10401) );
  AOI22_X1 U13319 ( .A1(n10556), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10545), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10399) );
  AND2_X1 U13320 ( .A1(n10399), .A2(n16293), .ZN(n10400) );
  NAND4_X1 U13321 ( .A1(n10403), .A2(n10402), .A3(n10401), .A4(n10400), .ZN(
        n10404) );
  INV_X2 U13322 ( .A(n10407), .ZN(n10438) );
  NAND2_X1 U13323 ( .A1(n10434), .A2(n10438), .ZN(n13284) );
  NAND4_X1 U13324 ( .A1(n11161), .A2(n11197), .A3(n10441), .A4(n19199), .ZN(
        n10406) );
  NOR2_X1 U13325 ( .A1(n10406), .A2(n10439), .ZN(n10451) );
  NAND2_X1 U13326 ( .A1(n10451), .A2(n19160), .ZN(n11166) );
  NAND2_X1 U13327 ( .A1(n13284), .A2(n11166), .ZN(n11215) );
  AOI22_X1 U13328 ( .A1(n10347), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10411) );
  AOI22_X1 U13329 ( .A1(n10548), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10553), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10410) );
  AOI22_X1 U13330 ( .A1(n12094), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10556), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10409) );
  AOI22_X1 U13331 ( .A1(n12225), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10545), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10408) );
  NAND4_X1 U13332 ( .A1(n10411), .A2(n10410), .A3(n10409), .A4(n10408), .ZN(
        n10412) );
  AOI22_X1 U13333 ( .A1(n10347), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12225), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10416) );
  AOI22_X1 U13334 ( .A1(n12094), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10415) );
  AOI22_X1 U13335 ( .A1(n10548), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10553), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10414) );
  AOI22_X1 U13336 ( .A1(n10556), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10545), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10413) );
  NAND4_X1 U13337 ( .A1(n10416), .A2(n10415), .A3(n10414), .A4(n10413), .ZN(
        n10417) );
  INV_X1 U13338 ( .A(n10425), .ZN(n10419) );
  NAND2_X2 U13339 ( .A1(n10419), .A2(n11190), .ZN(n10446) );
  INV_X1 U13340 ( .A(n10446), .ZN(n11224) );
  NOR2_X1 U13341 ( .A1(n10440), .A2(n10438), .ZN(n10420) );
  INV_X1 U13342 ( .A(n10445), .ZN(n11143) );
  NOR2_X1 U13343 ( .A1(n12237), .A2(n10441), .ZN(n10421) );
  AND3_X2 U13344 ( .A1(n10422), .A2(n11199), .A3(n10421), .ZN(n11189) );
  NAND2_X1 U13345 ( .A1(n10462), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10433) );
  NOR2_X1 U13346 ( .A1(n13299), .A2(n19859), .ZN(n10423) );
  AOI22_X1 U13347 ( .A1(n11050), .A2(P2_REIP_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10432) );
  NAND2_X1 U13348 ( .A1(n10424), .A2(n19199), .ZN(n10427) );
  NAND2_X1 U13349 ( .A1(n10425), .A2(n10441), .ZN(n10426) );
  NAND2_X1 U13350 ( .A1(n10427), .A2(n10426), .ZN(n10428) );
  AND2_X2 U13351 ( .A1(n11192), .A2(n11194), .ZN(n12235) );
  NAND2_X2 U13352 ( .A1(n12235), .A2(n19845), .ZN(n11207) );
  NAND2_X2 U13353 ( .A1(n10429), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11124) );
  INV_X1 U13354 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n10430) );
  OR2_X2 U13355 ( .A1(n11124), .A2(n10430), .ZN(n10431) );
  AND3_X2 U13356 ( .A1(n10433), .A2(n10432), .A3(n10431), .ZN(n10473) );
  INV_X1 U13357 ( .A(n10434), .ZN(n10437) );
  NAND2_X1 U13358 ( .A1(n19174), .A2(n19169), .ZN(n10435) );
  INV_X1 U13359 ( .A(n11192), .ZN(n10447) );
  NAND2_X1 U13360 ( .A1(n10447), .A2(n11197), .ZN(n10444) );
  NAND2_X1 U13361 ( .A1(n10440), .A2(n10439), .ZN(n11169) );
  NAND2_X1 U13362 ( .A1(n10446), .A2(n10424), .ZN(n11167) );
  AND2_X1 U13363 ( .A1(n19199), .A2(n11167), .ZN(n10442) );
  NAND2_X1 U13364 ( .A1(n11165), .A2(n10442), .ZN(n11196) );
  NAND2_X1 U13365 ( .A1(n11196), .A2(n19180), .ZN(n10443) );
  NAND3_X1 U13366 ( .A1(n10447), .A2(n13389), .A3(n10446), .ZN(n10448) );
  NAND2_X1 U13367 ( .A1(n10446), .A2(n19180), .ZN(n10450) );
  NAND2_X1 U13368 ( .A1(n10450), .A2(n19174), .ZN(n10453) );
  NOR2_X1 U13369 ( .A1(n10451), .A2(n19860), .ZN(n10452) );
  NAND2_X1 U13370 ( .A1(n19859), .A2(n16335), .ZN(n19853) );
  INV_X1 U13371 ( .A(n19853), .ZN(n16331) );
  XNOR2_X2 U13372 ( .A(n10473), .B(n10474), .ZN(n10492) );
  NAND2_X1 U13373 ( .A1(n11066), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10460) );
  NAND2_X1 U13374 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10457) );
  NAND2_X1 U13375 ( .A1(n19853), .A2(n10457), .ZN(n10458) );
  NAND2_X1 U13376 ( .A1(n10462), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10463) );
  OAI21_X1 U13377 ( .B1(n10465), .B2(n13299), .A(n10468), .ZN(n10467) );
  OAI21_X1 U13378 ( .B1(n10467), .B2(n10466), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n10472) );
  OR2_X1 U13379 ( .A1(n19853), .A2(n19841), .ZN(n10470) );
  INV_X1 U13380 ( .A(n10473), .ZN(n10475) );
  INV_X1 U13381 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14579) );
  AOI22_X1 U13382 ( .A1(n11050), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10479) );
  OAI21_X1 U13383 ( .B1(n10478), .B2(n14579), .A(n10479), .ZN(n10480) );
  INV_X1 U13384 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13589) );
  AOI21_X1 U13385 ( .B1(n19859), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10481) );
  INV_X1 U13386 ( .A(n10482), .ZN(n10484) );
  INV_X1 U13387 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14023) );
  INV_X1 U13388 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13855) );
  AOI22_X1 U13389 ( .A1(n11050), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10488) );
  XNOR2_X2 U13390 ( .A(n11040), .B(n11038), .ZN(n10522) );
  INV_X1 U13391 ( .A(n10490), .ZN(n10491) );
  INV_X1 U13392 ( .A(n10504), .ZN(n10502) );
  INV_X1 U13393 ( .A(n10493), .ZN(n10496) );
  INV_X1 U13394 ( .A(n10494), .ZN(n10495) );
  INV_X1 U13395 ( .A(n15646), .ZN(n18985) );
  AND2_X1 U13396 ( .A1(n10492), .A2(n18985), .ZN(n10510) );
  INV_X1 U13397 ( .A(n10510), .ZN(n10531) );
  INV_X1 U13398 ( .A(n10492), .ZN(n10501) );
  XNOR2_X2 U13399 ( .A(n10501), .B(n10498), .ZN(n14043) );
  INV_X1 U13400 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11976) );
  AND2_X1 U13401 ( .A1(n10502), .A2(n10523), .ZN(n10503) );
  NAND2_X1 U13402 ( .A1(n19329), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10507) );
  AND2_X1 U13403 ( .A1(n14598), .A2(n10510), .ZN(n10505) );
  NAND2_X1 U13404 ( .A1(n19269), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10506) );
  OAI211_X1 U13405 ( .C1(n19240), .C2(n11976), .A(n10507), .B(n10506), .ZN(
        n10508) );
  NAND2_X1 U13406 ( .A1(n10520), .A2(n15646), .ZN(n10530) );
  INV_X1 U13407 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11299) );
  NOR2_X1 U13408 ( .A1(n10601), .A2(n11299), .ZN(n10518) );
  NOR2_X2 U13409 ( .A1(n10519), .A2(n14043), .ZN(n10603) );
  NAND2_X1 U13410 ( .A1(n10603), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10516) );
  AOI21_X1 U13411 ( .B1(n19388), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A(
        n10512), .ZN(n10515) );
  AND2_X1 U13412 ( .A1(n14598), .A2(n10523), .ZN(n10513) );
  NAND2_X1 U13413 ( .A1(n19210), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10514) );
  NAND3_X1 U13414 ( .A1(n10516), .A2(n10515), .A3(n10514), .ZN(n10517) );
  NOR2_X1 U13415 ( .A1(n10518), .A2(n10517), .ZN(n10537) );
  INV_X1 U13416 ( .A(n10519), .ZN(n10521) );
  INV_X1 U13417 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11977) );
  NOR2_X1 U13418 ( .A1(n10602), .A2(n11977), .ZN(n10525) );
  INV_X1 U13419 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11969) );
  NAND2_X1 U13420 ( .A1(n14043), .A2(n15646), .ZN(n10526) );
  INV_X1 U13421 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11970) );
  OAI22_X1 U13422 ( .A1(n11969), .A2(n19580), .B1(n10752), .B2(n11970), .ZN(
        n10524) );
  NOR2_X1 U13423 ( .A1(n10525), .A2(n10524), .ZN(n10536) );
  INV_X1 U13424 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10529) );
  INV_X1 U13425 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n20917) );
  OAI22_X1 U13426 ( .A1(n10529), .A2(n19630), .B1(n19451), .B2(n20917), .ZN(
        n10534) );
  INV_X1 U13427 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11967) );
  INV_X1 U13428 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10571) );
  OAI22_X1 U13429 ( .A1(n11967), .A2(n19547), .B1(n19664), .B2(n10571), .ZN(
        n10533) );
  NOR2_X1 U13430 ( .A1(n10534), .A2(n10533), .ZN(n10535) );
  NAND3_X1 U13431 ( .A1(n10537), .A2(n10536), .A3(n10535), .ZN(n10599) );
  AND2_X1 U13432 ( .A1(n12095), .A2(n10538), .ZN(n10588) );
  AOI22_X1 U13433 ( .A1(n10588), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12066), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10544) );
  AND2_X1 U13434 ( .A1(n14532), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10626) );
  NAND2_X1 U13435 ( .A1(n10626), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10543) );
  NAND2_X1 U13436 ( .A1(n12064), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n10542) );
  AND2_X1 U13437 ( .A1(n14170), .A2(n12095), .ZN(n10574) );
  NAND2_X1 U13438 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10541) );
  NAND4_X1 U13439 ( .A1(n10544), .A2(n10543), .A3(n10542), .A4(n10541), .ZN(
        n10547) );
  NAND2_X1 U13440 ( .A1(n14542), .A2(n16293), .ZN(n11975) );
  INV_X1 U13441 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n21089) );
  INV_X1 U13442 ( .A(n10545), .ZN(n14536) );
  INV_X1 U13443 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n19555) );
  OAI22_X1 U13444 ( .A1(n11975), .A2(n21089), .B1(n10767), .B2(n19555), .ZN(
        n10546) );
  NOR2_X1 U13445 ( .A1(n10547), .A2(n10546), .ZN(n10563) );
  AND2_X2 U13446 ( .A1(n14539), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10654) );
  AND2_X2 U13447 ( .A1(n14539), .A2(n16293), .ZN(n10577) );
  AND2_X1 U13448 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10550) );
  AOI22_X1 U13449 ( .A1(n12085), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12065), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10551) );
  INV_X1 U13450 ( .A(n10551), .ZN(n10552) );
  AND2_X2 U13451 ( .A1(n14538), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12086) );
  NOR4_X1 U13452 ( .A1(n10314), .A2(n10304), .A3(n10552), .A4(n10313), .ZN(
        n10562) );
  NAND2_X2 U13453 ( .A1(n14537), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12078) );
  INV_X1 U13454 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10555) );
  INV_X1 U13455 ( .A(n10553), .ZN(n10554) );
  OR2_X1 U13456 ( .A1(n10554), .A2(n16293), .ZN(n12076) );
  INV_X1 U13457 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n20926) );
  OAI22_X1 U13458 ( .A1(n12078), .A2(n10555), .B1(n12076), .B2(n20926), .ZN(
        n10560) );
  INV_X1 U13459 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10558) );
  INV_X1 U13460 ( .A(n10556), .ZN(n12099) );
  NAND2_X2 U13461 ( .A1(n10557), .A2(n16293), .ZN(n12080) );
  INV_X1 U13462 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11280) );
  OAI22_X1 U13463 ( .A1(n12081), .A2(n10558), .B1(n12080), .B2(n11280), .ZN(
        n10559) );
  NOR2_X1 U13464 ( .A1(n10560), .A2(n10559), .ZN(n10561) );
  NOR2_X1 U13465 ( .A1(n11227), .A2(n19169), .ZN(n13365) );
  NAND2_X1 U13466 ( .A1(n10626), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10567) );
  NAND2_X1 U13467 ( .A1(n12064), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10566) );
  INV_X1 U13468 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19173) );
  AOI22_X1 U13469 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12065), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10565) );
  NAND2_X1 U13470 ( .A1(n10588), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10564) );
  NAND4_X1 U13471 ( .A1(n10567), .A2(n10566), .A3(n10565), .A4(n10564), .ZN(
        n10570) );
  INV_X1 U13472 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10568) );
  OAI22_X1 U13473 ( .A1(n10568), .A2(n11975), .B1(n10767), .B2(n11967), .ZN(
        n10569) );
  NOR2_X1 U13474 ( .A1(n10570), .A2(n10569), .ZN(n10581) );
  OAI22_X1 U13475 ( .A1(n12078), .A2(n11968), .B1(n12076), .B2(n20917), .ZN(
        n10573) );
  OAI22_X1 U13476 ( .A1(n10571), .A2(n12081), .B1(n12080), .B2(n11299), .ZN(
        n10572) );
  NOR2_X1 U13477 ( .A1(n10573), .A2(n10572), .ZN(n10580) );
  AOI22_X1 U13478 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10574), .B1(
        n12085), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10576) );
  NAND2_X1 U13479 ( .A1(n12086), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10575) );
  AND2_X1 U13480 ( .A1(n10576), .A2(n10575), .ZN(n10579) );
  AOI22_X1 U13481 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10577), .B1(
        n10654), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10578) );
  NAND4_X1 U13482 ( .A1(n10581), .A2(n10580), .A3(n10579), .A4(n10578), .ZN(
        n11236) );
  NAND2_X1 U13483 ( .A1(n13365), .A2(n11236), .ZN(n11000) );
  NAND2_X1 U13484 ( .A1(n10626), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n10585) );
  NAND2_X1 U13485 ( .A1(n12064), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n10584) );
  AOI22_X1 U13486 ( .A1(n12085), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12065), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10583) );
  NAND2_X1 U13487 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n10582) );
  NAND4_X1 U13488 ( .A1(n10585), .A2(n10584), .A3(n10583), .A4(n10582), .ZN(
        n10587) );
  INV_X1 U13489 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12016) );
  INV_X1 U13490 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11323) );
  OAI22_X1 U13491 ( .A1(n12016), .A2(n11975), .B1(n12080), .B2(n11323), .ZN(
        n10586) );
  NOR2_X1 U13492 ( .A1(n10587), .A2(n10586), .ZN(n10597) );
  NAND2_X1 U13493 ( .A1(n10577), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n10592) );
  NAND2_X1 U13494 ( .A1(n10654), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n10591) );
  AOI22_X1 U13495 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12066), .B1(
        n10588), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10590) );
  NAND2_X1 U13496 ( .A1(n12086), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n10589) );
  INV_X1 U13497 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10593) );
  INV_X1 U13498 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12017) );
  OAI22_X1 U13499 ( .A1(n12078), .A2(n10593), .B1(n12076), .B2(n12017), .ZN(
        n10596) );
  INV_X1 U13500 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12011) );
  INV_X1 U13501 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10594) );
  OAI22_X1 U13502 ( .A1(n12011), .A2(n10767), .B1(n12081), .B2(n10594), .ZN(
        n10595) );
  NAND2_X1 U13503 ( .A1(n11000), .A2(n11245), .ZN(n10598) );
  INV_X1 U13504 ( .A(n19664), .ZN(n10787) );
  AOI22_X1 U13505 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n10788), .B1(
        n10787), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10607) );
  INV_X1 U13506 ( .A(n10601), .ZN(n19425) );
  AOI22_X1 U13507 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19456), .B1(
        n19425), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10606) );
  NAND2_X1 U13508 ( .A1(n19358), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n10605) );
  NAND2_X1 U13509 ( .A1(n10603), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n10604) );
  NAND4_X1 U13510 ( .A1(n10607), .A2(n10606), .A3(n10605), .A4(n10604), .ZN(
        n10644) );
  INV_X1 U13511 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10609) );
  INV_X1 U13512 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10608) );
  INV_X1 U13513 ( .A(n10610), .ZN(n10625) );
  INV_X1 U13514 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10612) );
  INV_X1 U13515 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10613) );
  INV_X1 U13516 ( .A(n19388), .ZN(n10742) );
  INV_X1 U13517 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12002) );
  OAI22_X1 U13518 ( .A1(n10613), .A2(n10791), .B1(n10742), .B2(n12002), .ZN(
        n10614) );
  NOR2_X1 U13519 ( .A1(n10615), .A2(n10614), .ZN(n10624) );
  INV_X1 U13520 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10617) );
  INV_X1 U13521 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10616) );
  INV_X1 U13522 ( .A(n10618), .ZN(n10623) );
  INV_X1 U13523 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10619) );
  INV_X1 U13524 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11939) );
  NOR2_X1 U13525 ( .A1(n19154), .A2(n11939), .ZN(n10620) );
  NOR2_X1 U13526 ( .A1(n10621), .A2(n10620), .ZN(n10622) );
  NAND4_X1 U13527 ( .A1(n10625), .A2(n10624), .A3(n10623), .A4(n10622), .ZN(
        n10643) );
  NAND2_X1 U13528 ( .A1(n10626), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n10630) );
  NAND2_X1 U13529 ( .A1(n12064), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n10629) );
  AOI22_X1 U13530 ( .A1(n12085), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12065), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10628) );
  NAND2_X1 U13531 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n10627) );
  NAND4_X1 U13532 ( .A1(n10630), .A2(n10629), .A3(n10628), .A4(n10627), .ZN(
        n10634) );
  INV_X1 U13533 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11998) );
  NAND2_X1 U13534 ( .A1(n10588), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n10632) );
  NAND2_X1 U13535 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n10631) );
  OAI211_X1 U13536 ( .C1(n10767), .C2(n11998), .A(n10632), .B(n10631), .ZN(
        n10633) );
  NOR2_X1 U13537 ( .A1(n10634), .A2(n10633), .ZN(n10641) );
  INV_X1 U13538 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11999) );
  INV_X1 U13539 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10635) );
  OAI22_X1 U13540 ( .A1(n11999), .A2(n12076), .B1(n12081), .B2(n10635), .ZN(
        n10637) );
  INV_X1 U13541 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11343) );
  OAI22_X1 U13542 ( .A1(n12002), .A2(n11975), .B1(n12080), .B2(n11343), .ZN(
        n10636) );
  NOR2_X1 U13543 ( .A1(n10637), .A2(n10636), .ZN(n10640) );
  AOI22_X1 U13544 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10577), .B1(
        n12086), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10639) );
  AOI22_X1 U13545 ( .A1(n12050), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10654), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10638) );
  NAND4_X1 U13546 ( .A1(n10641), .A2(n10640), .A3(n10639), .A4(n10638), .ZN(
        n10670) );
  INV_X1 U13547 ( .A(n10670), .ZN(n11255) );
  NAND2_X1 U13548 ( .A1(n11255), .A2(n10512), .ZN(n10642) );
  NAND2_X1 U13549 ( .A1(n10646), .A2(n10645), .ZN(n10649) );
  INV_X1 U13550 ( .A(n10645), .ZN(n10648) );
  AOI22_X1 U13551 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10574), .B1(
        n10588), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10653) );
  NAND2_X1 U13552 ( .A1(n10577), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10652) );
  NAND2_X1 U13553 ( .A1(n12049), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10651) );
  NAND2_X1 U13554 ( .A1(n12086), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10650) );
  NAND4_X1 U13555 ( .A1(n10653), .A2(n10652), .A3(n10651), .A4(n10650), .ZN(
        n10660) );
  INV_X1 U13556 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12075) );
  OR2_X1 U13557 ( .A1(n12078), .A2(n12075), .ZN(n10658) );
  NAND2_X1 U13558 ( .A1(n10654), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10657) );
  NAND2_X1 U13559 ( .A1(n11278), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10656) );
  NAND2_X1 U13560 ( .A1(n12051), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10655) );
  NAND4_X1 U13561 ( .A1(n10658), .A2(n10657), .A3(n10656), .A4(n10655), .ZN(
        n10659) );
  AOI22_X1 U13562 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n12085), .B1(
        n12066), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10664) );
  NAND2_X1 U13563 ( .A1(n10626), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10663) );
  NAND2_X1 U13564 ( .A1(n12064), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10662) );
  NAND2_X1 U13565 ( .A1(n12065), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10661) );
  NAND4_X1 U13566 ( .A1(n10664), .A2(n10663), .A3(n10662), .A4(n10661), .ZN(
        n10667) );
  INV_X1 U13567 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10665) );
  INV_X1 U13568 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11424) );
  OAI22_X1 U13569 ( .A1(n11975), .A2(n10665), .B1(n12080), .B2(n11424), .ZN(
        n10666) );
  NOR2_X1 U13570 ( .A1(n10667), .A2(n10666), .ZN(n10668) );
  NOR2_X1 U13571 ( .A1(n13299), .A2(n10670), .ZN(n10671) );
  MUX2_X1 U13572 ( .A(n10671), .B(P2_EBX_REG_3__SCAN_IN), .S(n10689), .Z(
        n10678) );
  NAND2_X1 U13573 ( .A1(n13299), .A2(n9827), .ZN(n10728) );
  MUX2_X1 U13574 ( .A(n19831), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n11138) );
  NAND2_X1 U13575 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19841), .ZN(
        n10971) );
  INV_X1 U13576 ( .A(n10971), .ZN(n10673) );
  NAND2_X1 U13577 ( .A1(n11138), .A2(n10673), .ZN(n10983) );
  NAND2_X1 U13578 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n19831), .ZN(
        n10674) );
  NAND2_X1 U13579 ( .A1(n16296), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10680) );
  MUX2_X1 U13580 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n11933), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10729) );
  INV_X1 U13581 ( .A(n10729), .ZN(n10676) );
  XNOR2_X1 U13582 ( .A(n10730), .B(n10676), .ZN(n10975) );
  NOR2_X1 U13583 ( .A1(n10728), .A2(n10975), .ZN(n10677) );
  NOR2_X1 U13584 ( .A1(n10678), .A2(n10677), .ZN(n10684) );
  INV_X1 U13585 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13584) );
  NOR2_X1 U13586 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n10679) );
  MUX2_X1 U13587 ( .A(n10679), .B(n11236), .S(n9827), .Z(n10695) );
  NAND2_X1 U13588 ( .A1(n10684), .A2(n10695), .ZN(n10683) );
  OAI21_X1 U13589 ( .B1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n16296), .A(
        n10680), .ZN(n10681) );
  XNOR2_X1 U13590 ( .A(n10682), .B(n10681), .ZN(n11133) );
  INV_X1 U13591 ( .A(n11133), .ZN(n11142) );
  INV_X1 U13592 ( .A(n10780), .ZN(n10687) );
  INV_X1 U13593 ( .A(n10695), .ZN(n10698) );
  INV_X1 U13594 ( .A(n10684), .ZN(n10685) );
  OAI21_X1 U13595 ( .B1(n10699), .B2(n10698), .A(n10685), .ZN(n10686) );
  NAND2_X1 U13596 ( .A1(n10687), .A2(n10686), .ZN(n13856) );
  NAND2_X1 U13597 ( .A1(n10702), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13881) );
  NOR2_X1 U13598 ( .A1(n11227), .A2(n13299), .ZN(n10690) );
  MUX2_X1 U13599 ( .A(n10690), .B(P2_EBX_REG_0__SCAN_IN), .S(n10689), .Z(
        n10692) );
  OAI21_X1 U13600 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19841), .A(
        n10971), .ZN(n11135) );
  NOR2_X1 U13601 ( .A1(n10728), .A2(n11135), .ZN(n10691) );
  NOR2_X1 U13602 ( .A1(n10692), .A2(n10691), .ZN(n18981) );
  INV_X1 U13603 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13462) );
  OR2_X1 U13604 ( .A1(n18981), .A2(n13462), .ZN(n13364) );
  NAND2_X1 U13605 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n10693) );
  NOR2_X1 U13606 ( .A1(n9827), .A2(n10693), .ZN(n10694) );
  NOR2_X1 U13607 ( .A1(n10695), .A2(n10694), .ZN(n10696) );
  INV_X1 U13608 ( .A(n10696), .ZN(n14041) );
  NOR2_X1 U13609 ( .A1(n13364), .A2(n14041), .ZN(n10697) );
  INV_X1 U13610 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14096) );
  XOR2_X1 U13611 ( .A(n10696), .B(n13364), .Z(n13408) );
  NOR2_X1 U13612 ( .A1(n14096), .A2(n13408), .ZN(n13407) );
  NOR2_X1 U13613 ( .A1(n10697), .A2(n13407), .ZN(n14578) );
  XNOR2_X1 U13614 ( .A(n10699), .B(n10698), .ZN(n14577) );
  OR2_X1 U13615 ( .A1(n14578), .A2(n14577), .ZN(n14575) );
  NAND2_X1 U13616 ( .A1(n14578), .A2(n14577), .ZN(n10700) );
  NAND2_X1 U13617 ( .A1(n10700), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10701) );
  AND2_X1 U13618 ( .A1(n14575), .A2(n10701), .ZN(n13883) );
  NAND2_X1 U13619 ( .A1(n13881), .A2(n13883), .ZN(n10704) );
  INV_X1 U13620 ( .A(n10702), .ZN(n10703) );
  NAND2_X1 U13621 ( .A1(n10703), .A2(n14023), .ZN(n13882) );
  NAND2_X1 U13622 ( .A1(n10704), .A2(n13882), .ZN(n14020) );
  INV_X1 U13623 ( .A(n14020), .ZN(n10738) );
  INV_X1 U13624 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10705) );
  OR2_X1 U13625 ( .A1(n12078), .A2(n10705), .ZN(n10709) );
  AOI22_X1 U13626 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10574), .B1(
        n10588), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10708) );
  NAND2_X1 U13627 ( .A1(n12086), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10707) );
  NAND2_X1 U13628 ( .A1(n10654), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10706) );
  NAND4_X1 U13629 ( .A1(n10709), .A2(n10708), .A3(n10707), .A4(n10706), .ZN(
        n10715) );
  NAND2_X1 U13630 ( .A1(n10577), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10713) );
  NAND2_X1 U13631 ( .A1(n12049), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10712) );
  INV_X1 U13632 ( .A(n12080), .ZN(n13807) );
  NAND2_X1 U13633 ( .A1(n13807), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10711) );
  NAND2_X1 U13634 ( .A1(n11278), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n10710) );
  NAND4_X1 U13635 ( .A1(n10713), .A2(n10712), .A3(n10711), .A4(n10710), .ZN(
        n10714) );
  NOR2_X1 U13636 ( .A1(n10715), .A2(n10714), .ZN(n10725) );
  AOI22_X1 U13637 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n12085), .B1(
        n12066), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10719) );
  NAND2_X1 U13638 ( .A1(n10626), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10718) );
  NAND2_X1 U13639 ( .A1(n12064), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10717) );
  NAND2_X1 U13640 ( .A1(n12065), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10716) );
  NAND4_X1 U13641 ( .A1(n10719), .A2(n10718), .A3(n10717), .A4(n10716), .ZN(
        n10723) );
  INV_X1 U13642 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10721) );
  INV_X1 U13643 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10720) );
  OAI22_X1 U13644 ( .A1(n10721), .A2(n11975), .B1(n12081), .B2(n10720), .ZN(
        n10722) );
  NOR2_X1 U13645 ( .A1(n10723), .A2(n10722), .ZN(n10724) );
  INV_X1 U13646 ( .A(n11257), .ZN(n10726) );
  NAND2_X1 U13647 ( .A1(n19845), .A2(n10726), .ZN(n10727) );
  MUX2_X1 U13648 ( .A(n10727), .B(P2_EBX_REG_4__SCAN_IN), .S(n10689), .Z(
        n10736) );
  INV_X1 U13649 ( .A(n10728), .ZN(n10734) );
  NAND2_X1 U13650 ( .A1(n11933), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10731) );
  NOR2_X1 U13651 ( .A1(n16325), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10733) );
  NAND2_X1 U13652 ( .A1(n10978), .A2(n10733), .ZN(n10976) );
  NAND2_X1 U13653 ( .A1(n10734), .A2(n10976), .ZN(n10735) );
  NAND2_X1 U13654 ( .A1(n10736), .A2(n10735), .ZN(n10779) );
  XNOR2_X1 U13655 ( .A(n10780), .B(n10779), .ZN(n18971) );
  INV_X1 U13656 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n14119) );
  XNOR2_X1 U13657 ( .A(n18971), .B(n14119), .ZN(n14021) );
  INV_X1 U13658 ( .A(n14021), .ZN(n10737) );
  NAND2_X1 U13659 ( .A1(n10738), .A2(n10737), .ZN(n10740) );
  OR2_X1 U13660 ( .A1(n18971), .A2(n14119), .ZN(n10739) );
  NAND2_X1 U13661 ( .A1(n10740), .A2(n10739), .ZN(n14112) );
  INV_X1 U13662 ( .A(n19580), .ZN(n10789) );
  AOI22_X1 U13663 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n10789), .B1(
        n10787), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10751) );
  INV_X1 U13664 ( .A(n19630), .ZN(n10741) );
  AOI22_X1 U13665 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n10741), .B1(
        n19425), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10750) );
  INV_X1 U13666 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10743) );
  INV_X1 U13667 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10768) );
  OAI22_X1 U13668 ( .A1(n10743), .A2(n10791), .B1(n10742), .B2(n10768), .ZN(
        n10746) );
  INV_X1 U13669 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10744) );
  INV_X1 U13670 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12031) );
  OAI22_X1 U13671 ( .A1(n10744), .A2(n10792), .B1(n10794), .B2(n12031), .ZN(
        n10745) );
  NOR2_X1 U13672 ( .A1(n10746), .A2(n10745), .ZN(n10749) );
  INV_X1 U13673 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12036) );
  INV_X1 U13674 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13679) );
  OAI22_X1 U13675 ( .A1(n12036), .A2(n19240), .B1(n19154), .B2(n13679), .ZN(
        n10747) );
  INV_X1 U13676 ( .A(n10747), .ZN(n10748) );
  INV_X1 U13677 ( .A(n10752), .ZN(n10753) );
  AOI22_X1 U13678 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19456), .B1(
        n10753), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10758) );
  INV_X1 U13679 ( .A(n10754), .ZN(n10804) );
  AOI22_X1 U13680 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n10788), .B1(
        n10804), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10757) );
  NAND2_X1 U13681 ( .A1(n19358), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10756) );
  NAND2_X1 U13682 ( .A1(n10603), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n10755) );
  AOI22_X1 U13683 ( .A1(n10577), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10654), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10766) );
  INV_X1 U13684 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12028) );
  AOI22_X1 U13685 ( .A1(n10588), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12066), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10759) );
  OAI21_X1 U13686 ( .B1(n12078), .B2(n12028), .A(n10759), .ZN(n10760) );
  INV_X1 U13687 ( .A(n10760), .ZN(n10765) );
  AOI22_X1 U13688 ( .A1(n12049), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12086), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10764) );
  INV_X1 U13689 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10761) );
  INV_X1 U13690 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11384) );
  OAI22_X1 U13691 ( .A1(n12081), .A2(n10761), .B1(n12080), .B2(n11384), .ZN(
        n10762) );
  INV_X1 U13692 ( .A(n10762), .ZN(n10763) );
  NAND4_X1 U13693 ( .A1(n10766), .A2(n10765), .A3(n10764), .A4(n10763), .ZN(
        n10775) );
  INV_X1 U13694 ( .A(n10767), .ZN(n11278) );
  INV_X1 U13695 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12027) );
  OAI22_X1 U13696 ( .A1(n11975), .A2(n10768), .B1(n10767), .B2(n12027), .ZN(
        n10769) );
  INV_X1 U13697 ( .A(n10769), .ZN(n10773) );
  AOI22_X1 U13698 ( .A1(n10626), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10574), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10772) );
  AOI22_X1 U13699 ( .A1(n12085), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12065), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10771) );
  NAND2_X1 U13700 ( .A1(n12064), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n10770) );
  NAND4_X1 U13701 ( .A1(n10773), .A2(n10772), .A3(n10771), .A4(n10770), .ZN(
        n10774) );
  NOR2_X1 U13702 ( .A1(n10775), .A2(n10774), .ZN(n10781) );
  NAND2_X1 U13703 ( .A1(n10781), .A2(n10512), .ZN(n10776) );
  INV_X1 U13704 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n18951) );
  NAND2_X1 U13705 ( .A1(n10689), .A2(n18951), .ZN(n10782) );
  NAND2_X1 U13706 ( .A1(n11261), .A2(n10782), .ZN(n10783) );
  OAI21_X1 U13707 ( .B1(n10784), .B2(n10783), .A(n9904), .ZN(n18949) );
  INV_X1 U13708 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21044) );
  NAND2_X1 U13709 ( .A1(n10785), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10786) );
  AOI22_X1 U13710 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n10788), .B1(
        n10787), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10803) );
  AOI22_X1 U13711 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n10789), .B1(
        n19425), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10802) );
  INV_X1 U13712 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10793) );
  INV_X1 U13713 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10790) );
  OAI22_X1 U13714 ( .A1(n10793), .A2(n10792), .B1(n10791), .B2(n10790), .ZN(
        n10797) );
  INV_X1 U13715 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10795) );
  INV_X1 U13716 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12056) );
  OAI22_X1 U13717 ( .A1(n10795), .A2(n10794), .B1(n10742), .B2(n12056), .ZN(
        n10796) );
  NOR2_X1 U13718 ( .A1(n10797), .A2(n10796), .ZN(n10801) );
  INV_X1 U13719 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10798) );
  INV_X1 U13720 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19194) );
  OAI22_X1 U13721 ( .A1(n10798), .A2(n19240), .B1(n19154), .B2(n19194), .ZN(
        n10799) );
  INV_X1 U13722 ( .A(n10799), .ZN(n10800) );
  NAND4_X1 U13723 ( .A1(n10803), .A2(n10802), .A3(n10801), .A4(n10800), .ZN(
        n10810) );
  AOI22_X1 U13724 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n10741), .B1(
        n19456), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10808) );
  AOI22_X1 U13725 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n10804), .B1(
        n10753), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10807) );
  NAND2_X1 U13726 ( .A1(n10603), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n10806) );
  NAND2_X1 U13727 ( .A1(n19358), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n10805) );
  NAND4_X1 U13728 ( .A1(n10808), .A2(n10807), .A3(n10806), .A4(n10805), .ZN(
        n10809) );
  NAND2_X1 U13729 ( .A1(n10626), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n10814) );
  NAND2_X1 U13730 ( .A1(n12064), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n10813) );
  AOI22_X1 U13731 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12065), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10812) );
  NAND2_X1 U13732 ( .A1(n10588), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n10811) );
  NAND4_X1 U13733 ( .A1(n10814), .A2(n10813), .A3(n10812), .A4(n10811), .ZN(
        n10816) );
  INV_X1 U13734 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12047) );
  OAI22_X1 U13735 ( .A1(n11975), .A2(n12056), .B1(n10767), .B2(n12047), .ZN(
        n10815) );
  NOR2_X1 U13736 ( .A1(n10816), .A2(n10815), .ZN(n10825) );
  AOI22_X1 U13737 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12085), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10820) );
  NAND2_X1 U13738 ( .A1(n10577), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n10819) );
  NAND2_X1 U13739 ( .A1(n10654), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n10818) );
  NAND2_X1 U13740 ( .A1(n12086), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n10817) );
  INV_X1 U13741 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10821) );
  INV_X1 U13742 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12059) );
  OAI22_X1 U13743 ( .A1(n12078), .A2(n10821), .B1(n12076), .B2(n12059), .ZN(
        n10823) );
  INV_X1 U13744 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12222) );
  INV_X1 U13745 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11406) );
  OAI22_X1 U13746 ( .A1(n12081), .A2(n12222), .B1(n12080), .B2(n11406), .ZN(
        n10822) );
  NOR2_X1 U13747 ( .A1(n10823), .A2(n10822), .ZN(n10824) );
  NAND2_X1 U13748 ( .A1(n11265), .A2(n10512), .ZN(n10826) );
  NAND2_X1 U13749 ( .A1(n10829), .A2(n11012), .ZN(n10830) );
  NAND2_X1 U13750 ( .A1(n11015), .A2(n10960), .ZN(n10835) );
  INV_X1 U13751 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n13686) );
  INV_X1 U13752 ( .A(n11265), .ZN(n10831) );
  MUX2_X1 U13753 ( .A(n13686), .B(n10831), .S(n9827), .Z(n10832) );
  INV_X1 U13754 ( .A(n10852), .ZN(n10834) );
  NAND2_X1 U13755 ( .A1(n9904), .A2(n10143), .ZN(n10833) );
  NAND2_X1 U13756 ( .A1(n10834), .A2(n10833), .ZN(n18937) );
  NAND2_X1 U13757 ( .A1(n10835), .A2(n18937), .ZN(n10836) );
  INV_X1 U13758 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14186) );
  XNOR2_X1 U13759 ( .A(n10836), .B(n14186), .ZN(n14181) );
  NAND2_X1 U13760 ( .A1(n10836), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10837) );
  NOR2_X1 U13761 ( .A1(n9827), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n10838) );
  INV_X1 U13762 ( .A(n10841), .ZN(n10839) );
  XNOR2_X1 U13763 ( .A(n10852), .B(n10839), .ZN(n18929) );
  AND2_X1 U13764 ( .A1(n18929), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14216) );
  INV_X1 U13765 ( .A(n18929), .ZN(n10840) );
  INV_X1 U13766 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n14213) );
  NAND2_X1 U13767 ( .A1(n10840), .A2(n14213), .ZN(n10845) );
  INV_X1 U13768 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n11060) );
  NOR2_X1 U13769 ( .A1(n9827), .A2(n11060), .ZN(n10842) );
  AND2_X1 U13770 ( .A1(n10843), .A2(n10842), .ZN(n10844) );
  OR2_X1 U13771 ( .A1(n10844), .A2(n10850), .ZN(n13969) );
  NOR2_X1 U13772 ( .A1(n13969), .A2(n10960), .ZN(n10846) );
  NAND2_X1 U13773 ( .A1(n10846), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16224) );
  INV_X1 U13774 ( .A(n10845), .ZN(n14217) );
  INV_X1 U13775 ( .A(n10846), .ZN(n10847) );
  INV_X1 U13776 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11063) );
  INV_X1 U13777 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n13823) );
  NOR2_X1 U13778 ( .A1(n9827), .A2(n13823), .ZN(n10848) );
  XNOR2_X1 U13779 ( .A(n10850), .B(n10848), .ZN(n18917) );
  NAND2_X1 U13780 ( .A1(n18917), .A2(n11020), .ZN(n10849) );
  INV_X1 U13781 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16257) );
  NAND2_X1 U13782 ( .A1(n10849), .A2(n16257), .ZN(n15631) );
  NAND2_X1 U13783 ( .A1(n10689), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10851) );
  MUX2_X1 U13784 ( .A(n10851), .B(P2_EBX_REG_10__SCAN_IN), .S(n10854), .Z(
        n10853) );
  AND2_X1 U13785 ( .A1(n10853), .A2(n10942), .ZN(n13949) );
  NAND2_X1 U13786 ( .A1(n13949), .A2(n11020), .ZN(n10864) );
  INV_X1 U13787 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16268) );
  NAND2_X1 U13788 ( .A1(n10864), .A2(n16268), .ZN(n16203) );
  INV_X1 U13789 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n13951) );
  INV_X1 U13790 ( .A(n10866), .ZN(n10855) );
  INV_X1 U13791 ( .A(n10865), .ZN(n10858) );
  NAND3_X1 U13792 ( .A1(n10689), .A2(P2_EBX_REG_11__SCAN_IN), .A3(n10856), 
        .ZN(n10857) );
  NAND2_X1 U13793 ( .A1(n10858), .A2(n10857), .ZN(n18902) );
  OR2_X1 U13794 ( .A1(n18902), .A2(n10960), .ZN(n10859) );
  INV_X1 U13795 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11037) );
  NAND2_X1 U13796 ( .A1(n10861), .A2(n10860), .ZN(n11801) );
  NAND2_X1 U13797 ( .A1(n11020), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10862) );
  OR2_X1 U13798 ( .A1(n18902), .A2(n10862), .ZN(n16189) );
  NOR2_X1 U13799 ( .A1(n10960), .A2(n16257), .ZN(n10863) );
  NAND2_X1 U13800 ( .A1(n18917), .A2(n10863), .ZN(n16200) );
  OR2_X1 U13801 ( .A1(n16268), .A2(n10864), .ZN(n16202) );
  AND2_X1 U13802 ( .A1(n16200), .A2(n16202), .ZN(n16188) );
  NAND2_X1 U13803 ( .A1(n10689), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10867) );
  NOR2_X1 U13804 ( .A1(n10867), .A2(n10866), .ZN(n10868) );
  OR2_X1 U13805 ( .A1(n10894), .A2(n10868), .ZN(n14051) );
  NAND2_X1 U13806 ( .A1(n11020), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10869) );
  INV_X1 U13807 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16176) );
  OAI21_X1 U13808 ( .B1(n14051), .B2(n10960), .A(n16176), .ZN(n16178) );
  NAND2_X1 U13809 ( .A1(n10689), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10893) );
  INV_X1 U13810 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n10870) );
  NAND2_X1 U13811 ( .A1(n10892), .A2(n10870), .ZN(n10901) );
  NAND3_X1 U13812 ( .A1(n10901), .A2(P2_EBX_REG_15__SCAN_IN), .A3(n10689), 
        .ZN(n10872) );
  OAI21_X1 U13813 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(P2_EBX_REG_14__SCAN_IN), 
        .A(n10689), .ZN(n10871) );
  NAND2_X1 U13814 ( .A1(n10872), .A2(n10880), .ZN(n13295) );
  NOR2_X1 U13815 ( .A1(n10960), .A2(n13295), .ZN(n10906) );
  NOR2_X1 U13816 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n10906), .ZN(
        n11805) );
  INV_X1 U13817 ( .A(n11805), .ZN(n15584) );
  NOR2_X1 U13818 ( .A1(P2_EBX_REG_16__SCAN_IN), .A2(P2_EBX_REG_17__SCAN_IN), 
        .ZN(n10873) );
  INV_X1 U13819 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n11085) );
  NOR2_X1 U13820 ( .A1(n9827), .A2(n11085), .ZN(n10884) );
  NAND2_X1 U13821 ( .A1(n10689), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n10882) );
  INV_X1 U13822 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n10874) );
  INV_X1 U13823 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n15238) );
  NAND2_X1 U13824 ( .A1(n10689), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10875) );
  NOR2_X1 U13825 ( .A1(n10876), .A2(n10875), .ZN(n10877) );
  NOR2_X1 U13826 ( .A1(n10919), .A2(n10877), .ZN(n13326) );
  AOI21_X1 U13827 ( .B1(n13326), .B2(n11020), .A(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11813) );
  OR2_X1 U13828 ( .A1(n10880), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10888) );
  INV_X1 U13829 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n11078) );
  NOR2_X1 U13830 ( .A1(n9827), .A2(n11078), .ZN(n10879) );
  INV_X1 U13831 ( .A(n10942), .ZN(n10878) );
  AOI21_X1 U13832 ( .B1(n10880), .B2(n10879), .A(n10878), .ZN(n10881) );
  AND2_X1 U13833 ( .A1(n10888), .A2(n10881), .ZN(n18869) );
  NAND2_X1 U13834 ( .A1(n18869), .A2(n11020), .ZN(n10912) );
  XNOR2_X1 U13835 ( .A(n10912), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15428) );
  NOR2_X1 U13836 ( .A1(n10885), .A2(n10882), .ZN(n10883) );
  OR2_X1 U13837 ( .A1(n10896), .A2(n10883), .ZN(n18854) );
  NOR2_X1 U13838 ( .A1(n18854), .A2(n10960), .ZN(n10908) );
  NOR2_X1 U13839 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n10908), .ZN(
        n15532) );
  AND2_X1 U13840 ( .A1(n10889), .A2(n10884), .ZN(n10886) );
  OR2_X1 U13841 ( .A1(n10886), .A2(n10885), .ZN(n15173) );
  NOR2_X1 U13842 ( .A1(n15173), .A2(n10960), .ZN(n10909) );
  NOR2_X1 U13843 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n10909), .ZN(
        n15549) );
  NOR2_X1 U13844 ( .A1(n15532), .A2(n15549), .ZN(n11809) );
  INV_X1 U13845 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n11081) );
  NOR2_X1 U13846 ( .A1(n9827), .A2(n11081), .ZN(n10887) );
  NAND2_X1 U13847 ( .A1(n10888), .A2(n10887), .ZN(n10890) );
  NAND2_X1 U13848 ( .A1(n10890), .A2(n10889), .ZN(n13314) );
  NOR2_X1 U13849 ( .A1(n13314), .A2(n10960), .ZN(n10910) );
  NAND3_X1 U13850 ( .A1(n15428), .A2(n11809), .A3(n9910), .ZN(n10891) );
  NOR2_X1 U13851 ( .A1(n11813), .A2(n10891), .ZN(n10898) );
  INV_X1 U13852 ( .A(n10892), .ZN(n10900) );
  OAI21_X1 U13853 ( .B1(n10894), .B2(n10893), .A(n10900), .ZN(n18889) );
  NOR2_X1 U13854 ( .A1(n10960), .A2(n18889), .ZN(n10907) );
  NOR2_X1 U13855 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n10907), .ZN(
        n15619) );
  INV_X1 U13856 ( .A(n15619), .ZN(n10897) );
  NOR2_X1 U13857 ( .A1(n9827), .A2(n10874), .ZN(n10895) );
  XNOR2_X1 U13858 ( .A(n10896), .B(n10895), .ZN(n18842) );
  NAND2_X1 U13859 ( .A1(n18842), .A2(n11020), .ZN(n10911) );
  INV_X1 U13860 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15523) );
  NAND2_X1 U13861 ( .A1(n10911), .A2(n15523), .ZN(n11799) );
  NAND4_X1 U13862 ( .A1(n15584), .A2(n10898), .A3(n10897), .A4(n11799), .ZN(
        n10903) );
  NAND2_X1 U13863 ( .A1(n10900), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10899) );
  MUX2_X1 U13864 ( .A(n10900), .B(n10899), .S(n10689), .Z(n10902) );
  NAND2_X1 U13865 ( .A1(n10902), .A2(n10901), .ZN(n18879) );
  NOR2_X1 U13866 ( .A1(n10960), .A2(n18879), .ZN(n10905) );
  NOR2_X1 U13867 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n10905), .ZN(
        n11804) );
  NOR2_X1 U13868 ( .A1(n10903), .A2(n11804), .ZN(n10904) );
  NAND2_X1 U13869 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n10905), .ZN(
        n15600) );
  NAND2_X1 U13870 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n10906), .ZN(
        n15585) );
  NAND2_X1 U13871 ( .A1(n15600), .A2(n15585), .ZN(n11800) );
  AND2_X1 U13872 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n10907), .ZN(
        n15618) );
  INV_X1 U13873 ( .A(n15618), .ZN(n11803) );
  NAND2_X1 U13874 ( .A1(n10908), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15533) );
  NAND2_X1 U13875 ( .A1(n10909), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15551) );
  NAND2_X1 U13876 ( .A1(n15533), .A2(n15551), .ZN(n11810) );
  NAND2_X1 U13877 ( .A1(n10910), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11808) );
  NOR2_X1 U13878 ( .A1(n15523), .A2(n10911), .ZN(n11811) );
  INV_X1 U13879 ( .A(n11811), .ZN(n11798) );
  INV_X1 U13880 ( .A(n10912), .ZN(n10913) );
  NAND2_X1 U13881 ( .A1(n10913), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11807) );
  NAND3_X1 U13882 ( .A1(n11808), .A2(n11798), .A3(n11807), .ZN(n10914) );
  NOR2_X1 U13883 ( .A1(n11810), .A2(n10914), .ZN(n10917) );
  INV_X1 U13884 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11831) );
  NOR2_X1 U13885 ( .A1(n10960), .A2(n11831), .ZN(n10915) );
  AND2_X1 U13886 ( .A1(n13326), .A2(n10915), .ZN(n11812) );
  INV_X1 U13887 ( .A(n11812), .ZN(n10916) );
  NAND3_X1 U13888 ( .A1(n11803), .A2(n10917), .A3(n10916), .ZN(n10918) );
  NOR2_X1 U13889 ( .A1(n11800), .A2(n10918), .ZN(n15397) );
  NAND2_X1 U13890 ( .A1(n10689), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10920) );
  INV_X1 U13891 ( .A(n10920), .ZN(n10921) );
  NAND2_X1 U13892 ( .A1(n10922), .A2(n10921), .ZN(n10923) );
  NAND2_X1 U13893 ( .A1(n10927), .A2(n10923), .ZN(n15704) );
  INV_X1 U13894 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15509) );
  OR3_X1 U13895 ( .A1(n15704), .A2(n10960), .A3(n15509), .ZN(n15395) );
  AND2_X1 U13896 ( .A1(n15397), .A2(n15395), .ZN(n10924) );
  NAND2_X1 U13897 ( .A1(n15398), .A2(n10924), .ZN(n15387) );
  OR2_X1 U13898 ( .A1(n15704), .A2(n10960), .ZN(n10925) );
  NAND2_X1 U13899 ( .A1(n10925), .A2(n15509), .ZN(n15396) );
  INV_X1 U13900 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n11100) );
  NOR2_X1 U13901 ( .A1(n9827), .A2(n11100), .ZN(n10926) );
  NAND2_X1 U13902 ( .A1(n10927), .A2(n10926), .ZN(n10928) );
  NAND2_X1 U13903 ( .A1(n10938), .A2(n10928), .ZN(n13340) );
  OR2_X1 U13904 ( .A1(n13340), .A2(n10960), .ZN(n10929) );
  XNOR2_X1 U13905 ( .A(n10929), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15389) );
  AND2_X1 U13906 ( .A1(n15396), .A2(n15389), .ZN(n10930) );
  NAND2_X1 U13907 ( .A1(n15387), .A2(n10930), .ZN(n10933) );
  INV_X1 U13908 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11103) );
  OR2_X1 U13909 ( .A1(n10960), .A2(n11103), .ZN(n10931) );
  OR2_X1 U13910 ( .A1(n13340), .A2(n10931), .ZN(n10932) );
  NAND2_X1 U13911 ( .A1(n10689), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10934) );
  MUX2_X1 U13912 ( .A(P2_EBX_REG_24__SCAN_IN), .B(n10934), .S(n10938), .Z(
        n10935) );
  AND2_X1 U13913 ( .A1(n10935), .A2(n10942), .ZN(n16123) );
  NAND2_X1 U13914 ( .A1(n16123), .A2(n11020), .ZN(n15379) );
  INV_X1 U13915 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15482) );
  NOR2_X1 U13916 ( .A1(n15379), .A2(n15482), .ZN(n10937) );
  NAND2_X1 U13917 ( .A1(n15379), .A2(n15482), .ZN(n10936) );
  NAND2_X1 U13918 ( .A1(n10689), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n10939) );
  MUX2_X1 U13919 ( .A(n10939), .B(P2_EBX_REG_25__SCAN_IN), .S(n10941), .Z(
        n10940) );
  AOI21_X1 U13920 ( .B1(n16117), .B2(n11020), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15368) );
  INV_X1 U13921 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n15209) );
  NAND2_X1 U13922 ( .A1(n10941), .A2(n15209), .ZN(n10943) );
  NAND2_X1 U13923 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n10943), .ZN(n10944) );
  NOR2_X1 U13924 ( .A1(n9827), .A2(n10944), .ZN(n10945) );
  NOR2_X1 U13925 ( .A1(n10965), .A2(n10945), .ZN(n16099) );
  NAND2_X1 U13926 ( .A1(n16099), .A2(n11020), .ZN(n10953) );
  XNOR2_X1 U13927 ( .A(n10953), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15357) );
  NAND2_X1 U13928 ( .A1(n10689), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n16091) );
  NAND2_X1 U13929 ( .A1(n16089), .A2(n11020), .ZN(n11875) );
  INV_X1 U13930 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11210) );
  NOR2_X2 U13931 ( .A1(n11873), .A2(n10946), .ZN(n10955) );
  NAND2_X1 U13932 ( .A1(n10947), .A2(n11210), .ZN(n10950) );
  INV_X1 U13933 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n11118) );
  NOR2_X1 U13934 ( .A1(n9827), .A2(n11118), .ZN(n10948) );
  NOR2_X2 U13935 ( .A1(n16089), .A2(n10948), .ZN(n10957) );
  INV_X1 U13936 ( .A(n16117), .ZN(n10952) );
  INV_X1 U13937 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15459) );
  OR2_X1 U13938 ( .A1(n10960), .A2(n15459), .ZN(n10951) );
  INV_X1 U13939 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15464) );
  OR2_X1 U13940 ( .A1(n10953), .A2(n15464), .ZN(n10954) );
  NAND2_X1 U13941 ( .A1(n10689), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n10956) );
  XNOR2_X1 U13942 ( .A(n10957), .B(n10956), .ZN(n16064) );
  INV_X1 U13943 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14482) );
  OAI21_X1 U13944 ( .B1(n16064), .B2(n10960), .A(n14482), .ZN(n14470) );
  NAND2_X1 U13945 ( .A1(n10957), .A2(n10956), .ZN(n10966) );
  INV_X1 U13946 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n11123) );
  NOR2_X1 U13947 ( .A1(n9827), .A2(n11123), .ZN(n10958) );
  XNOR2_X1 U13948 ( .A(n10966), .B(n10958), .ZN(n14495) );
  INV_X1 U13949 ( .A(n14495), .ZN(n10959) );
  AOI21_X1 U13950 ( .B1(n10959), .B2(n11020), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11845) );
  INV_X1 U13951 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11858) );
  OR3_X1 U13952 ( .A1(n14495), .A2(n10960), .A3(n11858), .ZN(n11846) );
  INV_X1 U13953 ( .A(n11846), .ZN(n10963) );
  INV_X1 U13954 ( .A(n16064), .ZN(n10961) );
  NAND3_X1 U13955 ( .A1(n10961), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n11020), .ZN(n14469) );
  INV_X1 U13956 ( .A(n10965), .ZN(n10968) );
  NOR2_X1 U13957 ( .A1(n10966), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10967) );
  MUX2_X1 U13958 ( .A(n10968), .B(n10967), .S(n10689), .Z(n16049) );
  NAND2_X1 U13959 ( .A1(n16049), .A2(n11020), .ZN(n10969) );
  XOR2_X1 U13960 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n10969), .Z(
        n10970) );
  INV_X1 U13961 ( .A(n11138), .ZN(n10972) );
  NAND2_X1 U13962 ( .A1(n10972), .A2(n10971), .ZN(n10984) );
  INV_X1 U13963 ( .A(n10984), .ZN(n10974) );
  OAI21_X1 U13964 ( .B1(n11135), .B2(n10974), .A(n10973), .ZN(n10977) );
  NAND2_X1 U13965 ( .A1(n10977), .A2(n11146), .ZN(n10982) );
  NAND2_X1 U13966 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16316), .ZN(
        n10980) );
  NAND2_X1 U13967 ( .A1(n10982), .A2(n11150), .ZN(n19846) );
  NAND2_X1 U13968 ( .A1(n10512), .A2(n19860), .ZN(n13302) );
  NAND2_X1 U13969 ( .A1(n11146), .A2(n11133), .ZN(n10987) );
  AND2_X1 U13970 ( .A1(n10984), .A2(n10983), .ZN(n11136) );
  INV_X1 U13971 ( .A(n10987), .ZN(n10985) );
  NAND2_X1 U13972 ( .A1(n11136), .A2(n10985), .ZN(n10986) );
  OAI21_X1 U13973 ( .B1(n11135), .B2(n10987), .A(n13353), .ZN(n10988) );
  INV_X1 U13974 ( .A(n10988), .ZN(n10991) );
  NAND2_X1 U13975 ( .A1(n10549), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10989) );
  NAND2_X1 U13976 ( .A1(n10989), .A2(n16316), .ZN(n13388) );
  INV_X1 U13977 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n10990) );
  OAI21_X1 U13978 ( .B1(n10654), .B2(n13388), .A(n10990), .ZN(n19833) );
  MUX2_X1 U13979 ( .A(n10991), .B(n19833), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n16330) );
  INV_X1 U13980 ( .A(n16330), .ZN(n19844) );
  OAI22_X1 U13981 ( .A1(n19846), .A2(n13302), .B1(n10512), .B2(n19844), .ZN(
        n10993) );
  NAND2_X1 U13982 ( .A1(n10993), .A2(n16321), .ZN(n11177) );
  NAND2_X1 U13983 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16335), .ZN(n19735) );
  INV_X1 U13984 ( .A(n19735), .ZN(n10994) );
  NAND2_X1 U13985 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n10994), .ZN(n16341) );
  INV_X1 U13986 ( .A(n16341), .ZN(n13387) );
  NAND2_X1 U13987 ( .A1(n19860), .A2(n13387), .ZN(n10995) );
  NAND2_X1 U13988 ( .A1(n11184), .A2(n10996), .ZN(n11160) );
  XNOR2_X1 U13989 ( .A(n11227), .B(n11236), .ZN(n10998) );
  OR2_X1 U13990 ( .A1(n13365), .A2(n13462), .ZN(n13367) );
  INV_X1 U13991 ( .A(n13367), .ZN(n10997) );
  NAND2_X1 U13992 ( .A1(n10998), .A2(n10997), .ZN(n10999) );
  XOR2_X1 U13993 ( .A(n10998), .B(n10997), .Z(n13410) );
  NAND2_X1 U13994 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13410), .ZN(
        n13409) );
  NAND2_X1 U13995 ( .A1(n10999), .A2(n13409), .ZN(n11001) );
  XNOR2_X1 U13996 ( .A(n14579), .B(n11001), .ZN(n14570) );
  XNOR2_X1 U13997 ( .A(n11245), .B(n11000), .ZN(n14569) );
  NAND2_X1 U13998 ( .A1(n14570), .A2(n14569), .ZN(n14568) );
  NAND2_X1 U13999 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11001), .ZN(
        n11002) );
  NAND2_X1 U14000 ( .A1(n14568), .A2(n11002), .ZN(n11003) );
  NAND2_X1 U14001 ( .A1(n11003), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11004) );
  INV_X1 U14002 ( .A(n11007), .ZN(n11009) );
  INV_X1 U14003 ( .A(n14109), .ZN(n11013) );
  NAND2_X1 U14004 ( .A1(n11014), .A2(n14109), .ZN(n11016) );
  NAND2_X1 U14005 ( .A1(n11016), .A2(n11015), .ZN(n11017) );
  NAND2_X1 U14006 ( .A1(n11021), .A2(n11020), .ZN(n11019) );
  NAND3_X1 U14007 ( .A1(n11021), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n11020), .ZN(n11022) );
  NOR2_X1 U14008 ( .A1(n16268), .A2(n11037), .ZN(n16255) );
  NAND2_X1 U14009 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16255), .ZN(
        n15605) );
  INV_X1 U14010 ( .A(n15605), .ZN(n15603) );
  NAND3_X1 U14011 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n15603), .ZN(n15555) );
  INV_X1 U14012 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15608) );
  NOR2_X1 U14013 ( .A1(n15555), .A2(n15608), .ZN(n15568) );
  AND3_X1 U14014 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15557) );
  INV_X1 U14015 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15556) );
  INV_X1 U14016 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15543) );
  NAND2_X1 U14017 ( .A1(n15406), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11816) );
  NOR2_X2 U14018 ( .A1(n15371), .A2(n15459), .ZN(n15360) );
  OR2_X1 U14019 ( .A1(n10947), .A2(n14482), .ZN(n11842) );
  OR2_X1 U14020 ( .A1(n11842), .A2(n11858), .ZN(n11024) );
  NOR2_X2 U14021 ( .A1(n13356), .A2(n19169), .ZN(n16228) );
  OR2_X1 U14022 ( .A1(n11186), .A2(n19140), .ZN(n11158) );
  INV_X1 U14023 ( .A(n13274), .ZN(n11026) );
  AND2_X1 U14024 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11027) );
  INV_X1 U14025 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15419) );
  NAND2_X1 U14026 ( .A1(n13310), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13322) );
  INV_X1 U14027 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18865) );
  INV_X1 U14028 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n13327) );
  INV_X1 U14029 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n13341) );
  NAND2_X1 U14030 ( .A1(n13334), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14486) );
  INV_X1 U14031 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14488) );
  INV_X1 U14032 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16085) );
  INV_X1 U14033 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n21072) );
  INV_X1 U14034 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n11869) );
  NOR2_X1 U14035 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n14175) );
  INV_X1 U14036 ( .A(n14175), .ZN(n19809) );
  NAND2_X1 U14037 ( .A1(n19810), .A2(n19809), .ZN(n19823) );
  NAND2_X1 U14038 ( .A1(n19823), .A2(n19859), .ZN(n11029) );
  NAND2_X1 U14039 ( .A1(n19859), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n11938) );
  NAND2_X1 U14040 ( .A1(n19626), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n11030) );
  AND2_X1 U14041 ( .A1(n11938), .A2(n11030), .ZN(n13370) );
  NAND2_X1 U14042 ( .A1(n21095), .A2(n19859), .ZN(n15763) );
  INV_X1 U14043 ( .A(n15763), .ZN(n11031) );
  INV_X2 U14044 ( .A(n19138), .ZN(n18878) );
  AND2_X1 U14045 ( .A1(P2_REIP_REG_31__SCAN_IN), .A2(n16261), .ZN(n11486) );
  AOI21_X1 U14046 ( .B1(n19137), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n11486), .ZN(n11155) );
  INV_X1 U14047 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11034) );
  INV_X1 U14048 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n14083) );
  OR2_X1 U14049 ( .A1(n11131), .A2(n14083), .ZN(n11033) );
  AOI22_X1 U14050 ( .A1(n11125), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n11032) );
  OAI211_X1 U14051 ( .C1(n11128), .C2(n11034), .A(n11033), .B(n11032), .ZN(
        n13296) );
  INV_X1 U14052 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13874) );
  OR2_X1 U14053 ( .A1(n11131), .A2(n13874), .ZN(n11036) );
  AOI22_X1 U14054 ( .A1(n11125), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11035) );
  OAI211_X1 U14055 ( .C1(n11117), .C2(n11037), .A(n11036), .B(n11035), .ZN(
        n13870) );
  INV_X1 U14056 ( .A(n11038), .ZN(n11039) );
  NAND2_X1 U14057 ( .A1(n11040), .A2(n11039), .ZN(n11044) );
  OR2_X1 U14058 ( .A1(n11042), .A2(n11041), .ZN(n11043) );
  INV_X1 U14059 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n11045) );
  OR2_X1 U14060 ( .A1(n11131), .A2(n11045), .ZN(n11048) );
  AOI22_X1 U14061 ( .A1(n11050), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11047) );
  OR2_X1 U14062 ( .A1(n11117), .A2(n14119), .ZN(n11046) );
  OR2_X1 U14063 ( .A1(n11131), .A2(n18951), .ZN(n11053) );
  AOI22_X1 U14064 ( .A1(n11050), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11052) );
  OR2_X1 U14065 ( .A1(n11117), .A2(n21044), .ZN(n11051) );
  OR2_X1 U14066 ( .A1(n11131), .A2(n13686), .ZN(n11056) );
  AOI22_X1 U14067 ( .A1(n11125), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11055) );
  OR2_X1 U14068 ( .A1(n11128), .A2(n14186), .ZN(n11054) );
  INV_X1 U14069 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n11057) );
  OR2_X1 U14070 ( .A1(n11131), .A2(n11057), .ZN(n11059) );
  AOI22_X1 U14071 ( .A1(n11125), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11058) );
  OAI211_X1 U14072 ( .C1(n11128), .C2(n14213), .A(n11059), .B(n11058), .ZN(
        n13695) );
  OR2_X1 U14073 ( .A1(n11131), .A2(n11060), .ZN(n11062) );
  AOI22_X1 U14074 ( .A1(n11125), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11061) );
  OAI211_X1 U14075 ( .C1(n11128), .C2(n11063), .A(n11062), .B(n11061), .ZN(
        n13728) );
  OR2_X1 U14076 ( .A1(n11131), .A2(n13823), .ZN(n11065) );
  AOI22_X1 U14077 ( .A1(n11125), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11064) );
  OAI211_X1 U14078 ( .C1(n11128), .C2(n16257), .A(n11065), .B(n11064), .ZN(
        n13817) );
  INV_X1 U14079 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n11318) );
  INV_X1 U14080 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n16335) );
  OAI22_X1 U14081 ( .A1(n11075), .A2(n11318), .B1(n16335), .B2(n10058), .ZN(
        n11068) );
  NOR2_X1 U14082 ( .A1(n11128), .A2(n16268), .ZN(n11067) );
  AOI211_X1 U14083 ( .C1(n11066), .C2(P2_EBX_REG_10__SCAN_IN), .A(n11068), .B(
        n11067), .ZN(n13784) );
  INV_X1 U14084 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n14049) );
  OR2_X1 U14085 ( .A1(n11131), .A2(n14049), .ZN(n11070) );
  AOI22_X1 U14086 ( .A1(n11125), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n11069) );
  OAI211_X1 U14087 ( .C1(n11128), .C2(n16176), .A(n11070), .B(n11069), .ZN(
        n13893) );
  INV_X1 U14088 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11074) );
  INV_X1 U14089 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n11071) );
  OR2_X1 U14090 ( .A1(n11131), .A2(n11071), .ZN(n11073) );
  AOI22_X1 U14091 ( .A1(n11125), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n11072) );
  OAI211_X1 U14092 ( .C1(n11117), .C2(n11074), .A(n11073), .B(n11072), .ZN(
        n13911) );
  INV_X1 U14093 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n11400) );
  OAI22_X1 U14094 ( .A1(n11075), .A2(n11400), .B1(n16335), .B2(n10077), .ZN(
        n11077) );
  NOR2_X1 U14095 ( .A1(n11128), .A2(n15608), .ZN(n11076) );
  AOI211_X1 U14096 ( .C1(n11066), .C2(P2_EBX_REG_14__SCAN_IN), .A(n11077), .B(
        n11076), .ZN(n13958) );
  INV_X1 U14097 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15695) );
  OR2_X1 U14098 ( .A1(n11131), .A2(n11078), .ZN(n11080) );
  AOI22_X1 U14099 ( .A1(n11125), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n11079) );
  OAI211_X1 U14100 ( .C1(n11128), .C2(n15695), .A(n11080), .B(n11079), .ZN(
        n14155) );
  INV_X1 U14101 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11084) );
  OR2_X1 U14102 ( .A1(n11131), .A2(n11081), .ZN(n11083) );
  AOI22_X1 U14103 ( .A1(n11125), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n11082) );
  OAI211_X1 U14104 ( .C1(n11128), .C2(n11084), .A(n11083), .B(n11082), .ZN(
        n13315) );
  OR2_X1 U14105 ( .A1(n11131), .A2(n11085), .ZN(n11088) );
  AOI22_X1 U14106 ( .A1(n11125), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11087) );
  OR2_X1 U14107 ( .A1(n11128), .A2(n15556), .ZN(n11086) );
  NOR2_X2 U14108 ( .A1(n14232), .A2(n14233), .ZN(n14234) );
  INV_X1 U14109 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n11089) );
  OR2_X1 U14110 ( .A1(n11131), .A2(n11089), .ZN(n11091) );
  AOI22_X1 U14111 ( .A1(n11125), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n11090) );
  OAI211_X1 U14112 ( .C1(n11117), .C2(n15543), .A(n11091), .B(n11090), .ZN(
        n15253) );
  AND2_X2 U14113 ( .A1(n14234), .A2(n15253), .ZN(n15241) );
  OR2_X1 U14114 ( .A1(n11131), .A2(n10874), .ZN(n11093) );
  AOI22_X1 U14115 ( .A1(n11125), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n11092) );
  OAI211_X1 U14116 ( .C1(n11128), .C2(n15523), .A(n11093), .B(n11092), .ZN(
        n15242) );
  OR2_X1 U14117 ( .A1(n11131), .A2(n15238), .ZN(n11095) );
  AOI22_X1 U14118 ( .A1(n11125), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n11094) );
  OAI211_X1 U14119 ( .C1(n11117), .C2(n11831), .A(n11095), .B(n11094), .ZN(
        n11819) );
  INV_X1 U14120 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n11096) );
  OR2_X1 U14121 ( .A1(n11124), .A2(n11096), .ZN(n11099) );
  AOI22_X1 U14122 ( .A1(n11125), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11098) );
  OR2_X1 U14123 ( .A1(n11128), .A2(n15509), .ZN(n11097) );
  OR2_X1 U14124 ( .A1(n11131), .A2(n11100), .ZN(n11102) );
  AOI22_X1 U14125 ( .A1(n11125), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n11101) );
  OAI211_X1 U14126 ( .C1(n11128), .C2(n11103), .A(n11102), .B(n11101), .ZN(
        n13342) );
  INV_X1 U14127 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n11104) );
  OR2_X1 U14128 ( .A1(n11131), .A2(n11104), .ZN(n11107) );
  AOI22_X1 U14129 ( .A1(n11125), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n11106) );
  OR2_X1 U14130 ( .A1(n11128), .A2(n15482), .ZN(n11105) );
  OR2_X1 U14131 ( .A1(n11131), .A2(n15209), .ZN(n11110) );
  AOI22_X1 U14132 ( .A1(n11125), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n11109) );
  OR2_X1 U14133 ( .A1(n11128), .A2(n15459), .ZN(n11108) );
  OR2_X2 U14134 ( .A1(n15214), .A2(n15206), .ZN(n15208) );
  INV_X1 U14135 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n11111) );
  OR2_X1 U14136 ( .A1(n11131), .A2(n11111), .ZN(n11114) );
  AOI22_X1 U14137 ( .A1(n11125), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n11113) );
  OR2_X1 U14138 ( .A1(n11128), .A2(n15464), .ZN(n11112) );
  INV_X1 U14139 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n16086) );
  OR2_X1 U14140 ( .A1(n11131), .A2(n16086), .ZN(n11116) );
  AOI22_X1 U14141 ( .A1(n11125), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n11115) );
  OAI211_X1 U14142 ( .C1(n11117), .C2(n11210), .A(n11116), .B(n11115), .ZN(
        n15190) );
  OR2_X1 U14143 ( .A1(n11131), .A2(n11118), .ZN(n11120) );
  AOI22_X1 U14144 ( .A1(n11125), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n11119) );
  OAI211_X1 U14145 ( .C1(n11128), .C2(n10947), .A(n11120), .B(n11119), .ZN(
        n11883) );
  INV_X1 U14146 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n21118) );
  OR2_X1 U14147 ( .A1(n11131), .A2(n21118), .ZN(n11122) );
  AOI22_X1 U14148 ( .A1(n11125), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n11121) );
  OAI211_X1 U14149 ( .C1(n11128), .C2(n14482), .A(n11122), .B(n11121), .ZN(
        n14476) );
  OR2_X1 U14150 ( .A1(n11124), .A2(n11123), .ZN(n11127) );
  AOI22_X1 U14151 ( .A1(n11125), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11126) );
  OAI211_X1 U14152 ( .C1(n11128), .C2(n11858), .A(n11127), .B(n11126), .ZN(
        n11850) );
  INV_X1 U14153 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n16050) );
  AOI22_X1 U14154 ( .A1(n11125), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n11130) );
  INV_X1 U14155 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13281) );
  OR2_X1 U14156 ( .A1(n11128), .A2(n13281), .ZN(n11129) );
  OAI211_X1 U14157 ( .C1(n11131), .C2(n16050), .A(n11130), .B(n11129), .ZN(
        n11132) );
  NAND2_X1 U14158 ( .A1(n19813), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19827) );
  NOR2_X1 U14159 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16333) );
  INV_X1 U14160 ( .A(n16333), .ZN(n19857) );
  NAND2_X1 U14161 ( .A1(n19160), .A2(n19169), .ZN(n11134) );
  MUX2_X1 U14162 ( .A(n11134), .B(n13299), .S(n11133), .Z(n11145) );
  INV_X1 U14163 ( .A(n11135), .ZN(n11137) );
  OAI211_X1 U14164 ( .C1(n19169), .C2(n11137), .A(n19160), .B(n11136), .ZN(
        n11141) );
  NAND2_X1 U14165 ( .A1(n11138), .A2(n11137), .ZN(n11139) );
  NAND2_X1 U14166 ( .A1(n19845), .A2(n11139), .ZN(n11140) );
  OAI211_X1 U14167 ( .C1(n11143), .C2(n11142), .A(n11141), .B(n11140), .ZN(
        n11144) );
  NAND2_X1 U14168 ( .A1(n11145), .A2(n11144), .ZN(n11147) );
  MUX2_X1 U14169 ( .A(n13299), .B(n11147), .S(n11146), .Z(n11148) );
  NAND2_X1 U14170 ( .A1(n11148), .A2(n11150), .ZN(n11149) );
  MUX2_X1 U14171 ( .A(n11149), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n19859), .Z(n11162) );
  INV_X1 U14172 ( .A(n11150), .ZN(n11151) );
  NAND2_X1 U14173 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19834) );
  OAI221_X4 U14174 ( .B1(n19857), .B2(n16334), .C1(n19834), .C2(n16334), .A(
        n19859), .ZN(n19585) );
  NAND2_X1 U14175 ( .A1(n16045), .A2(n19146), .ZN(n11154) );
  OAI211_X1 U14176 ( .C1(n13282), .C2(n19150), .A(n11155), .B(n11154), .ZN(
        n11156) );
  NAND2_X1 U14177 ( .A1(n11160), .A2(n11159), .ZN(P2_U2983) );
  NAND2_X1 U14178 ( .A1(n16313), .A2(n19169), .ZN(n19058) );
  NAND2_X1 U14179 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n18818), .ZN(n19869) );
  NAND2_X2 U14180 ( .A1(n19792), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n19794) );
  INV_X1 U14181 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19736) );
  INV_X1 U14182 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19752) );
  NAND2_X1 U14183 ( .A1(n19736), .A2(n19752), .ZN(n19748) );
  NAND2_X1 U14184 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19858) );
  NAND2_X1 U14185 ( .A1(n11161), .A2(n13379), .ZN(n11181) );
  AOI21_X1 U14186 ( .B1(n11162), .B2(n19160), .A(n10441), .ZN(n11179) );
  AOI21_X1 U14187 ( .B1(n10512), .B2(n10424), .A(n19860), .ZN(n11163) );
  OAI21_X1 U14188 ( .B1(n11163), .B2(n12237), .A(n19174), .ZN(n11164) );
  AND3_X1 U14189 ( .A1(n11165), .A2(n10465), .A3(n11164), .ZN(n11173) );
  NAND2_X1 U14190 ( .A1(n11167), .A2(n19174), .ZN(n11168) );
  NAND2_X1 U14191 ( .A1(n11166), .A2(n11168), .ZN(n11172) );
  NAND2_X1 U14192 ( .A1(n11169), .A2(n19199), .ZN(n11170) );
  INV_X1 U14193 ( .A(n13302), .ZN(n19865) );
  NAND2_X1 U14194 ( .A1(n11170), .A2(n19865), .ZN(n11198) );
  NAND3_X1 U14195 ( .A1(n10434), .A2(n13353), .A3(n13379), .ZN(n11171) );
  NAND4_X1 U14196 ( .A1(n11173), .A2(n11172), .A3(n11198), .A4(n11171), .ZN(
        n13381) );
  INV_X1 U14197 ( .A(n13381), .ZN(n11176) );
  MUX2_X1 U14198 ( .A(n10434), .B(n11161), .S(n10512), .Z(n11174) );
  NAND3_X1 U14199 ( .A1(n11174), .A2(n13353), .A3(n19858), .ZN(n11175) );
  NAND3_X1 U14200 ( .A1(n11177), .A2(n11176), .A3(n11175), .ZN(n11178) );
  AOI21_X1 U14201 ( .B1(n19058), .B2(n11179), .A(n11178), .ZN(n11180) );
  OAI21_X1 U14202 ( .B1(n19058), .B2(n11181), .A(n11180), .ZN(n11182) );
  NAND2_X1 U14203 ( .A1(n11182), .A2(n13387), .ZN(n11219) );
  INV_X1 U14204 ( .A(n16321), .ZN(n19849) );
  NOR2_X1 U14205 ( .A1(n19849), .A2(n13299), .ZN(n11183) );
  AND2_X1 U14206 ( .A1(n16321), .A2(n19865), .ZN(n11185) );
  OR2_X1 U14207 ( .A1(n11186), .A2(n15637), .ZN(n11492) );
  INV_X1 U14208 ( .A(n16045), .ZN(n11489) );
  NAND2_X1 U14209 ( .A1(n14166), .A2(n10512), .ZN(n11187) );
  NAND2_X1 U14210 ( .A1(n11187), .A2(n10468), .ZN(n11188) );
  AND3_X1 U14211 ( .A1(n10512), .A2(n19174), .A3(n9827), .ZN(n11191) );
  AND2_X1 U14212 ( .A1(n11189), .A2(n11191), .ZN(n13796) );
  NAND2_X1 U14213 ( .A1(n11209), .A2(n13796), .ZN(n15572) );
  NAND2_X1 U14214 ( .A1(n10446), .A2(n10512), .ZN(n11193) );
  MUX2_X1 U14215 ( .A(n11193), .B(n13389), .S(n11192), .Z(n11195) );
  NAND2_X1 U14216 ( .A1(n11195), .A2(n11194), .ZN(n11206) );
  NAND2_X1 U14217 ( .A1(n11196), .A2(n19169), .ZN(n14167) );
  AOI21_X1 U14218 ( .B1(n14167), .B2(n11198), .A(n11197), .ZN(n11204) );
  INV_X1 U14219 ( .A(n11199), .ZN(n13352) );
  NAND2_X1 U14220 ( .A1(n10465), .A2(n10441), .ZN(n11200) );
  AOI22_X1 U14221 ( .A1(n13352), .A2(n11200), .B1(n19860), .B2(n11161), .ZN(
        n11201) );
  NAND2_X1 U14222 ( .A1(n11202), .A2(n11201), .ZN(n11203) );
  NOR2_X1 U14223 ( .A1(n11204), .A2(n11203), .ZN(n11205) );
  NAND2_X1 U14224 ( .A1(n15645), .A2(n11207), .ZN(n11208) );
  NAND2_X1 U14225 ( .A1(n11209), .A2(n11208), .ZN(n11211) );
  NOR2_X1 U14226 ( .A1(n10947), .A2(n11210), .ZN(n15436) );
  NAND2_X1 U14227 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15436), .ZN(
        n15434) );
  NOR3_X1 U14228 ( .A1(n15464), .A2(n15482), .A3(n15459), .ZN(n11484) );
  NOR2_X1 U14229 ( .A1(n14096), .A2(n13462), .ZN(n13461) );
  NOR2_X1 U14230 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13461), .ZN(
        n13900) );
  NOR3_X1 U14231 ( .A1(n14119), .A2(n14023), .A3(n21044), .ZN(n14187) );
  NAND2_X1 U14232 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14187), .ZN(
        n14182) );
  NAND2_X1 U14233 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16287) );
  NOR3_X1 U14234 ( .A1(n13900), .A2(n14182), .A3(n16287), .ZN(n11212) );
  INV_X1 U14235 ( .A(n11211), .ZN(n15574) );
  NAND2_X1 U14236 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13461), .ZN(
        n14572) );
  NAND2_X1 U14237 ( .A1(n11219), .A2(n18878), .ZN(n13483) );
  INV_X1 U14238 ( .A(n13483), .ZN(n14582) );
  AOI21_X1 U14239 ( .B1(n15574), .B2(n14572), .A(n14582), .ZN(n13901) );
  OAI21_X1 U14240 ( .B1(n15575), .B2(n11212), .A(n13901), .ZN(n16258) );
  NAND3_X1 U14241 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15568), .A3(
        n15557), .ZN(n15518) );
  NAND2_X1 U14242 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15520) );
  NOR3_X1 U14243 ( .A1(n16258), .A2(n15518), .A3(n15520), .ZN(n15494) );
  NAND4_X1 U14244 ( .A1(n15494), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A4(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11213) );
  NOR2_X1 U14245 ( .A1(n15604), .A2(n14582), .ZN(n15493) );
  INV_X1 U14246 ( .A(n15493), .ZN(n16256) );
  NAND2_X1 U14247 ( .A1(n11213), .A2(n16256), .ZN(n15481) );
  OAI21_X1 U14248 ( .B1(n15575), .B2(n11484), .A(n15481), .ZN(n15452) );
  AOI21_X1 U14249 ( .B1(n15434), .B2(n15604), .A(n15452), .ZN(n11859) );
  OAI21_X1 U14250 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15575), .A(
        n11859), .ZN(n11214) );
  NAND2_X1 U14251 ( .A1(n11214), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11488) );
  NAND2_X1 U14252 ( .A1(n11216), .A2(n19169), .ZN(n11217) );
  AND2_X1 U14253 ( .A1(n16308), .A2(n11217), .ZN(n11218) );
  NOR2_X2 U14254 ( .A1(n11219), .A2(n11218), .ZN(n16280) );
  INV_X1 U14255 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19786) );
  OR2_X1 U14256 ( .A1(n11233), .A2(n19786), .ZN(n11223) );
  NOR2_X1 U14257 ( .A1(n19199), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11221) );
  AOI22_X1 U14258 ( .A1(n11273), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n11225), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11222) );
  NAND2_X1 U14259 ( .A1(n11223), .A2(n11222), .ZN(n15282) );
  NAND2_X1 U14260 ( .A1(n11224), .A2(n11225), .ZN(n11243) );
  MUX2_X1 U14261 ( .A(n19199), .B(n19841), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n11226) );
  INV_X1 U14262 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18836) );
  OR2_X1 U14263 ( .A1(n11233), .A2(n18836), .ZN(n11232) );
  INV_X1 U14264 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n11229) );
  NAND2_X1 U14265 ( .A1(n19169), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11228) );
  OAI211_X1 U14266 ( .C1(n19199), .C2(n11229), .A(n11228), .B(n20990), .ZN(
        n11230) );
  INV_X1 U14267 ( .A(n11230), .ZN(n11231) );
  NAND2_X1 U14268 ( .A1(n11232), .A2(n11231), .ZN(n13474) );
  INV_X1 U14269 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19754) );
  OR2_X1 U14270 ( .A1(n11233), .A2(n19754), .ZN(n11235) );
  AOI22_X1 U14271 ( .A1(n11221), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n11225), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11234) );
  NAND2_X1 U14272 ( .A1(n11235), .A2(n11234), .ZN(n11240) );
  XNOR2_X1 U14273 ( .A(n13477), .B(n11240), .ZN(n13464) );
  INV_X1 U14274 ( .A(n11236), .ZN(n11239) );
  NAND2_X1 U14275 ( .A1(n10446), .A2(n19199), .ZN(n11237) );
  MUX2_X1 U14276 ( .A(n11237), .B(n19831), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n11238) );
  OAI21_X1 U14277 ( .B1(n11239), .B2(n11440), .A(n11238), .ZN(n13463) );
  NOR2_X1 U14278 ( .A1(n13464), .A2(n13463), .ZN(n11242) );
  NOR2_X1 U14279 ( .A1(n13477), .A2(n11240), .ZN(n11241) );
  NAND2_X1 U14280 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11244) );
  OAI211_X1 U14281 ( .C1(n11440), .C2(n11245), .A(n11244), .B(n11243), .ZN(
        n11248) );
  INV_X1 U14282 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19756) );
  OR2_X1 U14283 ( .A1(n11233), .A2(n19756), .ZN(n11247) );
  INV_X2 U14284 ( .A(n11313), .ZN(n11273) );
  AOI22_X1 U14285 ( .A1(n11273), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n11272), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11246) );
  NAND2_X1 U14286 ( .A1(n11247), .A2(n11246), .ZN(n14068) );
  NOR2_X1 U14287 ( .A1(n14069), .A2(n14068), .ZN(n14070) );
  NOR2_X1 U14288 ( .A1(n11249), .A2(n11248), .ZN(n11250) );
  INV_X1 U14289 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n13887) );
  OR2_X1 U14290 ( .A1(n11233), .A2(n13887), .ZN(n11254) );
  AOI22_X1 U14291 ( .A1(n11272), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11252) );
  NAND2_X1 U14292 ( .A1(n11273), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11251) );
  AND2_X1 U14293 ( .A1(n11252), .A2(n11251), .ZN(n11253) );
  OAI211_X1 U14294 ( .C1(n11255), .C2(n11440), .A(n11254), .B(n11253), .ZN(
        n13851) );
  INV_X1 U14295 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n11256) );
  OR2_X1 U14296 ( .A1(n11233), .A2(n11256), .ZN(n11260) );
  AOI22_X1 U14297 ( .A1(n11273), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n11272), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11259) );
  OR2_X1 U14298 ( .A1(n11440), .A2(n11257), .ZN(n11258) );
  INV_X1 U14299 ( .A(n11261), .ZN(n11262) );
  AOI22_X1 U14300 ( .A1(n11262), .A2(n11220), .B1(n11272), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11264) );
  AOI22_X1 U14301 ( .A1(n11355), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n11273), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n11263) );
  NAND2_X1 U14302 ( .A1(n11264), .A2(n11263), .ZN(n14115) );
  OR2_X1 U14303 ( .A1(n11440), .A2(n11265), .ZN(n11266) );
  NAND2_X1 U14304 ( .A1(n14114), .A2(n11266), .ZN(n13672) );
  INV_X1 U14305 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19760) );
  OR2_X1 U14306 ( .A1(n11233), .A2(n19760), .ZN(n11268) );
  AOI22_X1 U14307 ( .A1(n11273), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n11272), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11267) );
  NAND2_X1 U14308 ( .A1(n11268), .A2(n11267), .ZN(n13671) );
  AOI22_X1 U14309 ( .A1(n13672), .A2(n13671), .B1(n11220), .B2(n11269), .ZN(
        n11270) );
  INV_X1 U14310 ( .A(n11270), .ZN(n13674) );
  INV_X1 U14311 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19117) );
  INV_X1 U14312 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19762) );
  OAI222_X1 U14313 ( .A1(n11314), .A2(n14213), .B1(n11313), .B2(n19117), .C1(
        n11233), .C2(n19762), .ZN(n13673) );
  INV_X1 U14314 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n11271) );
  OR2_X1 U14315 ( .A1(n11233), .A2(n11271), .ZN(n11296) );
  AOI22_X1 U14316 ( .A1(n11273), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n11272), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11295) );
  NAND2_X1 U14317 ( .A1(n10626), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11277) );
  NAND2_X1 U14318 ( .A1(n12064), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11276) );
  AOI22_X1 U14319 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12065), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11275) );
  NAND2_X1 U14320 ( .A1(n10588), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11274) );
  NAND4_X1 U14321 ( .A1(n11277), .A2(n11276), .A3(n11275), .A4(n11274), .ZN(
        n11282) );
  INV_X1 U14322 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11279) );
  OAI22_X1 U14323 ( .A1(n11975), .A2(n11280), .B1(n10767), .B2(n11279), .ZN(
        n11281) );
  NOR2_X1 U14324 ( .A1(n11282), .A2(n11281), .ZN(n11292) );
  INV_X1 U14325 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11283) );
  OAI22_X1 U14326 ( .A1(n12078), .A2(n19555), .B1(n12076), .B2(n11283), .ZN(
        n11286) );
  INV_X1 U14327 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11284) );
  OAI22_X1 U14328 ( .A1(n12081), .A2(n11284), .B1(n12080), .B2(n20926), .ZN(
        n11285) );
  NOR2_X1 U14329 ( .A1(n11286), .A2(n11285), .ZN(n11291) );
  AOI22_X1 U14330 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12085), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11288) );
  NAND2_X1 U14331 ( .A1(n12086), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11287) );
  AND2_X1 U14332 ( .A1(n11288), .A2(n11287), .ZN(n11290) );
  AOI22_X1 U14333 ( .A1(n10577), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10654), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11289) );
  NAND4_X1 U14334 ( .A1(n11292), .A2(n11291), .A3(n11290), .A4(n11289), .ZN(
        n13815) );
  INV_X1 U14335 ( .A(n13815), .ZN(n11293) );
  OR2_X1 U14336 ( .A1(n11440), .A2(n11293), .ZN(n11294) );
  AOI22_X1 U14337 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12066), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11297) );
  OAI21_X1 U14338 ( .B1(n11967), .B2(n12078), .A(n11297), .ZN(n11298) );
  INV_X1 U14339 ( .A(n11298), .ZN(n11304) );
  AOI22_X1 U14340 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10577), .B1(
        n12049), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11303) );
  AOI22_X1 U14341 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n10654), .B1(
        n12086), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11302) );
  OAI22_X1 U14342 ( .A1(n11299), .A2(n11975), .B1(n12081), .B2(n19173), .ZN(
        n11300) );
  INV_X1 U14343 ( .A(n11300), .ZN(n11301) );
  NAND4_X1 U14344 ( .A1(n11304), .A2(n11303), .A3(n11302), .A4(n11301), .ZN(
        n11311) );
  OAI22_X1 U14345 ( .A1(n11969), .A2(n10767), .B1(n12080), .B2(n20917), .ZN(
        n11305) );
  INV_X1 U14346 ( .A(n11305), .ZN(n11309) );
  AOI22_X1 U14347 ( .A1(n12064), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n12065), .ZN(n11308) );
  AOI22_X1 U14348 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12085), .B1(
        n10588), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11307) );
  NAND2_X1 U14349 ( .A1(n10626), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11306) );
  NAND4_X1 U14350 ( .A1(n11309), .A2(n11308), .A3(n11307), .A4(n11306), .ZN(
        n11310) );
  INV_X1 U14351 ( .A(n13814), .ZN(n11317) );
  INV_X1 U14352 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n11312) );
  OR2_X1 U14353 ( .A1(n11233), .A2(n11312), .ZN(n11316) );
  AOI22_X1 U14354 ( .A1(n11273), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n11272), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11315) );
  OAI211_X1 U14355 ( .C1(n11317), .C2(n11440), .A(n11316), .B(n11315), .ZN(
        n13669) );
  OR2_X1 U14356 ( .A1(n11233), .A2(n11318), .ZN(n11338) );
  AOI22_X1 U14357 ( .A1(n11273), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n11272), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11337) );
  NAND2_X1 U14358 ( .A1(n10626), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11322) );
  NAND2_X1 U14359 ( .A1(n12064), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n11321) );
  AOI22_X1 U14360 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12065), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11320) );
  NAND2_X1 U14361 ( .A1(n10588), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11319) );
  NAND4_X1 U14362 ( .A1(n11322), .A2(n11321), .A3(n11320), .A4(n11319), .ZN(
        n11326) );
  INV_X1 U14363 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11324) );
  OAI22_X1 U14364 ( .A1(n11324), .A2(n10767), .B1(n11975), .B2(n11323), .ZN(
        n11325) );
  NOR2_X1 U14365 ( .A1(n11326), .A2(n11325), .ZN(n11335) );
  INV_X1 U14366 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11327) );
  OAI22_X1 U14367 ( .A1(n12078), .A2(n12011), .B1(n12076), .B2(n11327), .ZN(
        n11329) );
  INV_X1 U14368 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11920) );
  OAI22_X1 U14369 ( .A1(n11920), .A2(n12081), .B1(n12080), .B2(n12017), .ZN(
        n11328) );
  NOR2_X1 U14370 ( .A1(n11329), .A2(n11328), .ZN(n11334) );
  AOI22_X1 U14371 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10574), .B1(
        n12085), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11331) );
  NAND2_X1 U14372 ( .A1(n12086), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n11330) );
  AND2_X1 U14373 ( .A1(n11331), .A2(n11330), .ZN(n11333) );
  AOI22_X1 U14374 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10577), .B1(
        n10654), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11332) );
  NAND4_X1 U14375 ( .A1(n11335), .A2(n11334), .A3(n11333), .A4(n11332), .ZN(
        n13783) );
  OR2_X1 U14376 ( .A1(n11440), .A2(n11951), .ZN(n11336) );
  NAND2_X1 U14377 ( .A1(n12064), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11342) );
  NAND2_X1 U14378 ( .A1(n10626), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11341) );
  AOI22_X1 U14379 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12065), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11340) );
  NAND2_X1 U14380 ( .A1(n10588), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11339) );
  NAND4_X1 U14381 ( .A1(n11342), .A2(n11341), .A3(n11340), .A4(n11339), .ZN(
        n11345) );
  OAI22_X1 U14382 ( .A1(n11939), .A2(n12081), .B1(n11975), .B2(n11343), .ZN(
        n11344) );
  NOR2_X1 U14383 ( .A1(n11345), .A2(n11344), .ZN(n11354) );
  AOI22_X1 U14384 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10574), .B1(
        n12085), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11349) );
  NAND2_X1 U14385 ( .A1(n10577), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n11348) );
  NAND2_X1 U14386 ( .A1(n12049), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11347) );
  NAND2_X1 U14387 ( .A1(n12086), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n11346) );
  AND4_X1 U14388 ( .A1(n11349), .A2(n11348), .A3(n11347), .A4(n11346), .ZN(
        n11353) );
  AOI22_X1 U14389 ( .A1(n12050), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10654), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11352) );
  OAI22_X1 U14390 ( .A1(n11999), .A2(n12080), .B1(n10767), .B2(n10609), .ZN(
        n11350) );
  INV_X1 U14391 ( .A(n11350), .ZN(n11351) );
  NAND4_X1 U14392 ( .A1(n11354), .A2(n11353), .A3(n11352), .A4(n11351), .ZN(
        n13867) );
  NAND2_X1 U14393 ( .A1(n11355), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n11357) );
  AOI22_X1 U14394 ( .A1(n11273), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n11272), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11356) );
  OAI211_X1 U14395 ( .C1(n9833), .C2(n11440), .A(n11357), .B(n11356), .ZN(
        n13694) );
  INV_X1 U14396 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n11358) );
  OR2_X1 U14397 ( .A1(n11233), .A2(n11358), .ZN(n11379) );
  AOI22_X1 U14398 ( .A1(n11273), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n11272), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11378) );
  NAND2_X1 U14399 ( .A1(n10626), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11362) );
  NAND2_X1 U14400 ( .A1(n12064), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11361) );
  AOI22_X1 U14401 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12065), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11360) );
  NAND2_X1 U14402 ( .A1(n10588), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11359) );
  NAND4_X1 U14403 ( .A1(n11362), .A2(n11361), .A3(n11360), .A4(n11359), .ZN(
        n11366) );
  INV_X1 U14404 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11364) );
  INV_X1 U14405 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11363) );
  OAI22_X1 U14406 ( .A1(n11364), .A2(n10767), .B1(n11975), .B2(n11363), .ZN(
        n11365) );
  NOR2_X1 U14407 ( .A1(n11366), .A2(n11365), .ZN(n11376) );
  INV_X1 U14408 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11985) );
  INV_X1 U14409 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11367) );
  OAI22_X1 U14410 ( .A1(n12078), .A2(n11985), .B1(n12076), .B2(n11367), .ZN(
        n11370) );
  INV_X1 U14411 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11368) );
  INV_X1 U14412 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11990) );
  OAI22_X1 U14413 ( .A1(n11368), .A2(n12081), .B1(n12080), .B2(n11990), .ZN(
        n11369) );
  NOR2_X1 U14414 ( .A1(n11370), .A2(n11369), .ZN(n11375) );
  AOI22_X1 U14415 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10574), .B1(
        n12085), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11372) );
  NAND2_X1 U14416 ( .A1(n12086), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11371) );
  AND2_X1 U14417 ( .A1(n11372), .A2(n11371), .ZN(n11374) );
  AOI22_X1 U14418 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n10654), .B1(
        n10577), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11373) );
  NAND4_X1 U14419 ( .A1(n11376), .A2(n11375), .A3(n11374), .A4(n11373), .ZN(
        n11953) );
  INV_X1 U14420 ( .A(n11953), .ZN(n13914) );
  OR2_X1 U14421 ( .A1(n11440), .A2(n13914), .ZN(n11377) );
  NAND2_X1 U14422 ( .A1(n12064), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11383) );
  NAND2_X1 U14423 ( .A1(n10626), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11382) );
  AOI22_X1 U14424 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12065), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11381) );
  NAND2_X1 U14425 ( .A1(n10588), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11380) );
  NAND4_X1 U14426 ( .A1(n11383), .A2(n11382), .A3(n11381), .A4(n11380), .ZN(
        n11386) );
  INV_X1 U14427 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12029) );
  OAI22_X1 U14428 ( .A1(n11975), .A2(n11384), .B1(n10767), .B2(n12029), .ZN(
        n11385) );
  NOR2_X1 U14429 ( .A1(n11386), .A2(n11385), .ZN(n11396) );
  AOI22_X1 U14430 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12085), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11390) );
  NAND2_X1 U14431 ( .A1(n10654), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11389) );
  NAND2_X1 U14432 ( .A1(n12049), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11388) );
  NAND2_X1 U14433 ( .A1(n12086), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11387) );
  AND4_X1 U14434 ( .A1(n11390), .A2(n11389), .A3(n11388), .A4(n11387), .ZN(
        n11395) );
  AOI22_X1 U14435 ( .A1(n12050), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10577), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11394) );
  INV_X1 U14436 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11391) );
  OAI22_X1 U14437 ( .A1(n12081), .A2(n13679), .B1(n12080), .B2(n11391), .ZN(
        n11392) );
  INV_X1 U14438 ( .A(n11392), .ZN(n11393) );
  NAND4_X1 U14439 ( .A1(n11396), .A2(n11395), .A3(n11394), .A4(n11393), .ZN(
        n11952) );
  INV_X1 U14440 ( .A(n11952), .ZN(n13913) );
  INV_X1 U14441 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n11397) );
  OR2_X1 U14442 ( .A1(n11233), .A2(n11397), .ZN(n11399) );
  AOI22_X1 U14443 ( .A1(n11273), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n11272), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11398) );
  OAI211_X1 U14444 ( .C1(n13913), .C2(n11440), .A(n11399), .B(n11398), .ZN(
        n13812) );
  OR2_X1 U14445 ( .A1(n11233), .A2(n11400), .ZN(n11421) );
  AOI22_X1 U14446 ( .A1(n11273), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n11272), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11420) );
  NAND2_X1 U14447 ( .A1(n10626), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11404) );
  NAND2_X1 U14448 ( .A1(n12064), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11403) );
  AOI22_X1 U14449 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12065), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11402) );
  NAND2_X1 U14450 ( .A1(n10588), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11401) );
  NAND4_X1 U14451 ( .A1(n11404), .A2(n11403), .A3(n11402), .A4(n11401), .ZN(
        n11408) );
  INV_X1 U14452 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11405) );
  OAI22_X1 U14453 ( .A1(n11975), .A2(n11406), .B1(n10767), .B2(n11405), .ZN(
        n11407) );
  NOR2_X1 U14454 ( .A1(n11408), .A2(n11407), .ZN(n11418) );
  AOI22_X1 U14455 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12085), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11412) );
  NAND2_X1 U14456 ( .A1(n10577), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n11411) );
  NAND2_X1 U14457 ( .A1(n10654), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11410) );
  NAND2_X1 U14458 ( .A1(n12086), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11409) );
  AND4_X1 U14459 ( .A1(n11412), .A2(n11411), .A3(n11410), .A4(n11409), .ZN(
        n11417) );
  INV_X1 U14460 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11413) );
  OAI22_X1 U14461 ( .A1(n12078), .A2(n12047), .B1(n12076), .B2(n11413), .ZN(
        n11415) );
  OAI22_X1 U14462 ( .A1(n12081), .A2(n19194), .B1(n12080), .B2(n12059), .ZN(
        n11414) );
  NOR2_X1 U14463 ( .A1(n11415), .A2(n11414), .ZN(n11416) );
  OR2_X1 U14464 ( .A1(n11440), .A2(n13956), .ZN(n11419) );
  AOI22_X1 U14465 ( .A1(n12050), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10577), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11429) );
  AOI22_X1 U14466 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n10654), .B1(
        n12049), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11428) );
  AOI22_X1 U14467 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10574), .B1(
        n10588), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11423) );
  NAND2_X1 U14468 ( .A1(n12086), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11422) );
  AND2_X1 U14469 ( .A1(n11423), .A2(n11422), .ZN(n11427) );
  INV_X1 U14470 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12077) );
  OAI22_X1 U14471 ( .A1(n11975), .A2(n11424), .B1(n10767), .B2(n12077), .ZN(
        n11425) );
  INV_X1 U14472 ( .A(n11425), .ZN(n11426) );
  NAND4_X1 U14473 ( .A1(n11429), .A2(n11428), .A3(n11427), .A4(n11426), .ZN(
        n11436) );
  INV_X1 U14474 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12072) );
  OAI22_X1 U14475 ( .A1(n12072), .A2(n12080), .B1(n12081), .B2(n19207), .ZN(
        n11430) );
  INV_X1 U14476 ( .A(n11430), .ZN(n11434) );
  AOI22_X1 U14477 ( .A1(n12064), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12065), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11433) );
  AOI22_X1 U14478 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n12085), .B1(
        n12066), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11432) );
  NAND2_X1 U14479 ( .A1(n10626), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11431) );
  NAND4_X1 U14480 ( .A1(n11434), .A2(n11433), .A3(n11432), .A4(n11431), .ZN(
        n11435) );
  INV_X1 U14481 ( .A(n14079), .ZN(n11441) );
  INV_X1 U14482 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n11437) );
  OR2_X1 U14483 ( .A1(n11233), .A2(n11437), .ZN(n11439) );
  AOI22_X1 U14484 ( .A1(n11273), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n11272), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11438) );
  OAI211_X1 U14485 ( .C1(n11441), .C2(n11440), .A(n11439), .B(n11438), .ZN(
        n13303) );
  INV_X1 U14486 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n11442) );
  OR2_X1 U14487 ( .A1(n11233), .A2(n11442), .ZN(n11444) );
  AOI22_X1 U14488 ( .A1(n11273), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n11272), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11443) );
  INV_X1 U14489 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19773) );
  OR2_X1 U14490 ( .A1(n11233), .A2(n19773), .ZN(n11446) );
  AOI22_X1 U14491 ( .A1(n11273), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n11225), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11445) );
  NAND2_X1 U14492 ( .A1(n11446), .A2(n11445), .ZN(n13316) );
  INV_X1 U14493 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n11447) );
  OR2_X1 U14494 ( .A1(n11233), .A2(n11447), .ZN(n11449) );
  AOI22_X1 U14495 ( .A1(n11273), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n11272), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11448) );
  INV_X1 U14496 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19776) );
  OR2_X1 U14497 ( .A1(n11233), .A2(n19776), .ZN(n11451) );
  AOI22_X1 U14498 ( .A1(n11273), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n11272), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11450) );
  NAND2_X1 U14499 ( .A1(n11451), .A2(n11450), .ZN(n15325) );
  INV_X1 U14500 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n11452) );
  OR2_X1 U14501 ( .A1(n11233), .A2(n11452), .ZN(n11454) );
  AOI22_X1 U14502 ( .A1(n11273), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n11272), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11453) );
  AND2_X1 U14503 ( .A1(n11454), .A2(n11453), .ZN(n15317) );
  INV_X1 U14504 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19779) );
  OR2_X1 U14505 ( .A1(n11233), .A2(n19779), .ZN(n11456) );
  AOI22_X1 U14506 ( .A1(n11273), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n11272), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11455) );
  NAND2_X1 U14507 ( .A1(n11456), .A2(n11455), .ZN(n11830) );
  OR2_X1 U14508 ( .A1(n11233), .A2(n19781), .ZN(n11458) );
  AOI22_X1 U14509 ( .A1(n11273), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n11225), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11457) );
  NAND2_X1 U14510 ( .A1(n11458), .A2(n11457), .ZN(n15299) );
  INV_X1 U14511 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19783) );
  OR2_X1 U14512 ( .A1(n11233), .A2(n19783), .ZN(n11460) );
  AOI22_X1 U14513 ( .A1(n11273), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n11225), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11459) );
  NAND2_X1 U14514 ( .A1(n11460), .A2(n11459), .ZN(n13343) );
  INV_X1 U14515 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n11461) );
  OR2_X1 U14516 ( .A1(n11233), .A2(n11461), .ZN(n11463) );
  AOI22_X1 U14517 ( .A1(n11273), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n11225), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11462) );
  AND2_X1 U14518 ( .A1(n11463), .A2(n11462), .ZN(n15484) );
  NAND2_X1 U14519 ( .A1(n15282), .A2(n15283), .ZN(n15285) );
  INV_X1 U14520 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n11464) );
  OR2_X1 U14521 ( .A1(n11233), .A2(n11464), .ZN(n11466) );
  AOI22_X1 U14522 ( .A1(n11273), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n11225), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11465) );
  AND2_X1 U14523 ( .A1(n11466), .A2(n11465), .ZN(n15276) );
  INV_X1 U14524 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19790) );
  OR2_X1 U14525 ( .A1(n11233), .A2(n19790), .ZN(n11468) );
  AOI22_X1 U14526 ( .A1(n11273), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n11225), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11467) );
  NAND2_X1 U14527 ( .A1(n11468), .A2(n11467), .ZN(n15267) );
  INV_X1 U14528 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n11469) );
  OR2_X1 U14529 ( .A1(n11233), .A2(n11469), .ZN(n11471) );
  AOI22_X1 U14530 ( .A1(n11273), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n11225), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11470) );
  NAND2_X1 U14531 ( .A1(n11471), .A2(n11470), .ZN(n14503) );
  INV_X1 U14532 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n21124) );
  OR2_X1 U14533 ( .A1(n11233), .A2(n21124), .ZN(n11473) );
  AOI22_X1 U14534 ( .A1(n11273), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n11225), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11472) );
  NAND2_X1 U14535 ( .A1(n11473), .A2(n11472), .ZN(n12238) );
  INV_X1 U14536 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n11474) );
  OR2_X1 U14537 ( .A1(n11233), .A2(n11474), .ZN(n11476) );
  AOI22_X1 U14538 ( .A1(n11273), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n11225), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11475) );
  AND2_X1 U14539 ( .A1(n11476), .A2(n11475), .ZN(n11851) );
  INV_X1 U14540 ( .A(n11851), .ZN(n11477) );
  NAND2_X1 U14541 ( .A1(n11478), .A2(n11477), .ZN(n11854) );
  INV_X1 U14542 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19796) );
  AOI22_X1 U14543 ( .A1(n11273), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n11225), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11479) );
  OAI21_X1 U14544 ( .B1(n11233), .B2(n19796), .A(n11479), .ZN(n11480) );
  INV_X1 U14545 ( .A(n15520), .ZN(n11483) );
  AOI21_X1 U14546 ( .B1(n15572), .B2(n14572), .A(n13900), .ZN(n11481) );
  INV_X1 U14547 ( .A(n16288), .ZN(n11482) );
  INV_X1 U14548 ( .A(n16254), .ZN(n15554) );
  NOR2_X1 U14549 ( .A1(n15518), .A2(n15554), .ZN(n15544) );
  NAND2_X1 U14550 ( .A1(n11483), .A2(n15544), .ZN(n11834) );
  NOR2_X1 U14551 ( .A1(n11831), .A2(n11834), .ZN(n15508) );
  NAND3_X1 U14552 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n15508), .ZN(n15483) );
  INV_X1 U14553 ( .A(n15483), .ZN(n15457) );
  NAND2_X1 U14554 ( .A1(n11484), .A2(n15457), .ZN(n15447) );
  NOR4_X1 U14555 ( .A1(n15447), .A2(n15434), .A3(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A4(n11858), .ZN(n11485) );
  OAI211_X1 U14556 ( .C1(n11489), .C2(n16272), .A(n11488), .B(n11487), .ZN(
        n11490) );
  INV_X1 U14557 ( .A(n11490), .ZN(n11491) );
  NAND2_X1 U14558 ( .A1(n11494), .A2(n11493), .ZN(P2_U3015) );
  NOR2_X4 U14559 ( .A1(n18754), .A2(n11495), .ZN(n15657) );
  AOI22_X1 U14560 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11508) );
  NOR4_X4 U14561 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(n18774), .A4(n18754), .ZN(
        n11716) );
  INV_X2 U14562 ( .A(n9850), .ZN(n17137) );
  AOI22_X1 U14563 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9834), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11497) );
  NOR3_X4 U14564 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n18601), .ZN(n17122) );
  AOI22_X1 U14565 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11496) );
  OAI211_X1 U14566 ( .C1(n10288), .C2(n21009), .A(n11497), .B(n11496), .ZN(
        n11506) );
  NOR2_X2 U14567 ( .A1(n16880), .A2(n11498), .ZN(n11519) );
  BUF_X4 U14568 ( .A(n11519), .Z(n17108) );
  AOI22_X1 U14569 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11504) );
  AOI22_X1 U14570 ( .A1(n9831), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17139), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11503) );
  AOI22_X1 U14571 ( .A1(n17128), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17107), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11502) );
  INV_X2 U14572 ( .A(n11702), .ZN(n17138) );
  INV_X2 U14573 ( .A(n16974), .ZN(n17144) );
  AOI22_X1 U14574 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11501) );
  NAND4_X1 U14575 ( .A1(n11504), .A2(n11503), .A3(n11502), .A4(n11501), .ZN(
        n11505) );
  AOI211_X1 U14576 ( .C1(n17145), .C2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A(
        n11506), .B(n11505), .ZN(n11507) );
  NAND2_X1 U14577 ( .A1(n11508), .A2(n11507), .ZN(n17747) );
  AOI22_X1 U14578 ( .A1(n17128), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17107), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11512) );
  AOI22_X1 U14579 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11511) );
  AOI22_X1 U14580 ( .A1(n17139), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9834), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11510) );
  AOI22_X1 U14581 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11509) );
  NAND4_X1 U14582 ( .A1(n11512), .A2(n11511), .A3(n11510), .A4(n11509), .ZN(
        n11518) );
  AOI22_X1 U14583 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11516) );
  AOI22_X1 U14584 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9831), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11515) );
  AOI22_X1 U14585 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9832), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11514) );
  AOI22_X1 U14586 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11513) );
  NAND4_X1 U14587 ( .A1(n11516), .A2(n11515), .A3(n11514), .A4(n11513), .ZN(
        n11517) );
  AOI22_X1 U14588 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9832), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11523) );
  AOI22_X1 U14589 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11522) );
  AOI22_X1 U14590 ( .A1(n17139), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11521) );
  BUF_X4 U14591 ( .A(n17122), .Z(n17094) );
  AOI22_X1 U14592 ( .A1(n17094), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17107), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11520) );
  NAND4_X1 U14593 ( .A1(n11523), .A2(n11522), .A3(n11521), .A4(n11520), .ZN(
        n11529) );
  AOI22_X1 U14594 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11527) );
  AOI22_X1 U14595 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17140), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11526) );
  AOI22_X1 U14596 ( .A1(n9831), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9834), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11525) );
  AOI22_X1 U14597 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11716), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11524) );
  NAND4_X1 U14598 ( .A1(n11527), .A2(n11526), .A3(n11525), .A4(n11524), .ZN(
        n11528) );
  INV_X1 U14599 ( .A(n11684), .ZN(n11696) );
  AOI22_X1 U14600 ( .A1(n9831), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9824), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11533) );
  AOI22_X1 U14601 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9834), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11532) );
  AOI22_X1 U14602 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11581), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11531) );
  INV_X2 U14603 ( .A(n17142), .ZN(n17123) );
  AOI22_X1 U14604 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11530) );
  NAND4_X1 U14605 ( .A1(n11533), .A2(n11532), .A3(n11531), .A4(n11530), .ZN(
        n11540) );
  AOI22_X1 U14606 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n15657), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11538) );
  AOI22_X1 U14607 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11537) );
  AOI22_X1 U14608 ( .A1(n11545), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11534), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11536) );
  AOI22_X1 U14609 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11716), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11535) );
  NAND4_X1 U14610 ( .A1(n11538), .A2(n11537), .A3(n11536), .A4(n11535), .ZN(
        n11539) );
  AOI22_X1 U14611 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9824), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11553) );
  INV_X1 U14612 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17183) );
  AOI22_X1 U14613 ( .A1(n11581), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9834), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11541) );
  OAI21_X1 U14614 ( .B1(n11702), .B2(n17183), .A(n11541), .ZN(n11542) );
  INV_X1 U14615 ( .A(n11542), .ZN(n11552) );
  AOI22_X1 U14616 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11716), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11543) );
  AOI22_X1 U14617 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n15657), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11548) );
  AOI22_X1 U14618 ( .A1(n11545), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11544), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11547) );
  NAND3_X1 U14619 ( .A1(n11548), .A2(n11547), .A3(n11546), .ZN(n11549) );
  NOR2_X1 U14620 ( .A1(n11550), .A2(n11549), .ZN(n11551) );
  AOI22_X1 U14621 ( .A1(n9831), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11555) );
  AOI22_X1 U14622 ( .A1(n17094), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11554) );
  AOI22_X1 U14623 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11566) );
  INV_X1 U14624 ( .A(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n20900) );
  AOI22_X1 U14625 ( .A1(n17094), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11558) );
  AOI22_X1 U14626 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9832), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11557) );
  OAI211_X1 U14627 ( .C1(n17004), .C2(n20900), .A(n11558), .B(n11557), .ZN(
        n11564) );
  AOI22_X1 U14628 ( .A1(n9834), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17107), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11562) );
  AOI22_X1 U14629 ( .A1(n9831), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11561) );
  AOI22_X1 U14630 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17140), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11560) );
  AOI22_X1 U14631 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17139), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11559) );
  NAND4_X1 U14632 ( .A1(n11562), .A2(n11561), .A3(n11560), .A4(n11559), .ZN(
        n11563) );
  AOI211_X1 U14633 ( .C1(n17146), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n11564), .B(n11563), .ZN(n11565) );
  NAND2_X1 U14634 ( .A1(n11566), .A2(n11565), .ZN(n11767) );
  NAND2_X1 U14635 ( .A1(n11594), .A2(n11767), .ZN(n11597) );
  AOI22_X1 U14636 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17140), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11570) );
  AOI22_X1 U14637 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17153), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11569) );
  AOI22_X1 U14638 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17139), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11568) );
  AOI22_X1 U14639 ( .A1(n9831), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9832), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11567) );
  NAND4_X1 U14640 ( .A1(n11570), .A2(n11569), .A3(n11568), .A4(n11567), .ZN(
        n11576) );
  AOI22_X1 U14641 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n9830), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11574) );
  AOI22_X1 U14642 ( .A1(n9834), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17094), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11573) );
  AOI22_X1 U14643 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11572) );
  AOI22_X1 U14644 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n17146), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11571) );
  NAND4_X1 U14645 ( .A1(n11574), .A2(n11573), .A3(n11572), .A4(n11571), .ZN(
        n11575) );
  INV_X1 U14646 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18071) );
  INV_X1 U14647 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21073) );
  NOR2_X1 U14648 ( .A1(n11776), .A2(n21073), .ZN(n11588) );
  AOI22_X1 U14649 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17094), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11580) );
  AOI22_X1 U14650 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17107), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11579) );
  AOI22_X1 U14651 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17139), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11578) );
  AOI22_X1 U14652 ( .A1(n9831), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11577) );
  NAND4_X1 U14653 ( .A1(n11580), .A2(n11579), .A3(n11578), .A4(n11577), .ZN(
        n11587) );
  AOI22_X1 U14654 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11585) );
  AOI22_X1 U14655 ( .A1(n9834), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11584) );
  AOI22_X1 U14656 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11581), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11583) );
  AOI22_X1 U14657 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11716), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11582) );
  NAND4_X1 U14658 ( .A1(n11585), .A2(n11584), .A3(n11583), .A4(n11582), .ZN(
        n11586) );
  NOR2_X1 U14659 ( .A1(n11587), .A2(n11586), .ZN(n11772) );
  NAND2_X1 U14660 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15768), .ZN(
        n17816) );
  NOR2_X1 U14661 ( .A1(n17816), .A2(n11774), .ZN(n17807) );
  NOR2_X1 U14662 ( .A1(n11588), .A2(n17807), .ZN(n17797) );
  INV_X1 U14663 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18122) );
  NOR2_X1 U14664 ( .A1(n17797), .A2(n17798), .ZN(n11590) );
  XNOR2_X1 U14665 ( .A(n11773), .B(n17334), .ZN(n11591) );
  INV_X1 U14666 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n17788) );
  NOR2_X1 U14667 ( .A1(n11592), .A2(n11591), .ZN(n11593) );
  INV_X1 U14668 ( .A(n11767), .ZN(n17331) );
  XNOR2_X1 U14669 ( .A(n11594), .B(n17331), .ZN(n11595) );
  XNOR2_X1 U14670 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n11595), .ZN(
        n17773) );
  NOR2_X2 U14671 ( .A1(n17772), .A2(n11596), .ZN(n11599) );
  XNOR2_X1 U14672 ( .A(n11597), .B(n17327), .ZN(n11598) );
  NOR2_X1 U14673 ( .A1(n11599), .A2(n11598), .ZN(n11600) );
  INV_X1 U14674 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18088) );
  XOR2_X1 U14675 ( .A(n11601), .B(n17747), .Z(n11602) );
  XNOR2_X1 U14676 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n11602), .ZN(
        n17753) );
  AOI21_X1 U14677 ( .B1(n16381), .B2(n17321), .A(n17724), .ZN(n11604) );
  INV_X1 U14678 ( .A(n11604), .ZN(n11605) );
  XNOR2_X1 U14679 ( .A(n11606), .B(n11605), .ZN(n17737) );
  NOR2_X1 U14680 ( .A1(n11606), .A2(n11605), .ZN(n11607) );
  INV_X1 U14681 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18057) );
  INV_X1 U14682 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18021) );
  NAND2_X1 U14683 ( .A1(n17703), .A2(n18021), .ZN(n17692) );
  INV_X1 U14684 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17679) );
  INV_X1 U14685 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21186) );
  INV_X1 U14686 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17971) );
  INV_X1 U14687 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17950) );
  NOR2_X2 U14688 ( .A1(n11608), .A2(n18057), .ZN(n18011) );
  NAND2_X1 U14689 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18014) );
  NOR2_X1 U14690 ( .A1(n18014), .A2(n17679), .ZN(n17658) );
  NAND2_X1 U14691 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17658), .ZN(
        n17965) );
  INV_X1 U14692 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17991) );
  NOR2_X1 U14693 ( .A1(n17965), .A2(n17991), .ZN(n17637) );
  NAND2_X1 U14694 ( .A1(n17637), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17951) );
  NOR2_X1 U14695 ( .A1(n17951), .A2(n17950), .ZN(n17613) );
  INV_X1 U14696 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17947) );
  INV_X1 U14697 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17931) );
  NAND2_X1 U14698 ( .A1(n17609), .A2(n17931), .ZN(n17608) );
  NOR2_X1 U14699 ( .A1(n17947), .A2(n17931), .ZN(n17923) );
  NAND2_X1 U14700 ( .A1(n17923), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17896) );
  INV_X1 U14701 ( .A(n17896), .ZN(n17585) );
  INV_X1 U14702 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17584) );
  INV_X1 U14703 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17568) );
  NOR2_X1 U14704 ( .A1(n17584), .A2(n17568), .ZN(n17898) );
  AND2_X1 U14705 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17898), .ZN(
        n17884) );
  NAND2_X1 U14706 ( .A1(n17585), .A2(n17884), .ZN(n17886) );
  INV_X1 U14707 ( .A(n17886), .ZN(n17544) );
  NAND2_X1 U14708 ( .A1(n17544), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17871) );
  INV_X1 U14709 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17863) );
  OR2_X1 U14710 ( .A1(n17871), .A2(n17863), .ZN(n17524) );
  NOR2_X1 U14711 ( .A1(n17724), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17598) );
  NAND2_X1 U14712 ( .A1(n17598), .A2(n17584), .ZN(n11610) );
  NOR2_X1 U14713 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n11610), .ZN(
        n17563) );
  INV_X1 U14714 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17555) );
  NAND2_X1 U14715 ( .A1(n17563), .A2(n17555), .ZN(n17542) );
  NOR3_X1 U14716 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n17542), .ZN(n11611) );
  INV_X1 U14717 ( .A(n11609), .ZN(n17953) );
  NAND2_X1 U14718 ( .A1(n17953), .A2(n17923), .ZN(n17561) );
  AND2_X1 U14719 ( .A1(n17884), .A2(n10309), .ZN(n11613) );
  INV_X1 U14720 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17850) );
  OR2_X1 U14721 ( .A1(n17724), .A2(n17517), .ZN(n17509) );
  OAI211_X1 U14722 ( .C1(n17510), .C2(n17850), .A(n17509), .B(n10296), .ZN(
        n17493) );
  INV_X1 U14723 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17831) );
  NOR2_X1 U14724 ( .A1(n17850), .A2(n17831), .ZN(n11760) );
  INV_X1 U14725 ( .A(n11760), .ZN(n17825) );
  AND2_X1 U14726 ( .A1(n17724), .A2(n17825), .ZN(n11614) );
  NOR2_X1 U14727 ( .A1(n17492), .A2(n11616), .ZN(n11617) );
  NOR2_X2 U14728 ( .A1(n11617), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16388) );
  NOR2_X1 U14729 ( .A1(n17724), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16380) );
  NOR2_X1 U14730 ( .A1(n17724), .A2(n11619), .ZN(n11625) );
  NAND2_X1 U14731 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n11617), .ZN(
        n17483) );
  NAND2_X1 U14732 ( .A1(n17724), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16378) );
  OAI21_X1 U14733 ( .B1(n17483), .B2(n16378), .A(n11618), .ZN(n15682) );
  INV_X1 U14734 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17465) );
  INV_X1 U14735 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18758) );
  AOI22_X1 U14736 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17724), .B1(
        n10101), .B2(n18758), .ZN(n11622) );
  NAND2_X1 U14737 ( .A1(n15753), .A2(n11622), .ZN(n11624) );
  INV_X1 U14738 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16348) );
  NAND2_X1 U14739 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16348), .ZN(
        n11907) );
  NOR2_X1 U14740 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16348), .ZN(
        n11620) );
  AOI211_X1 U14741 ( .C1(n11907), .C2(n11621), .A(n11625), .B(n11620), .ZN(
        n11623) );
  OAI22_X1 U14742 ( .A1(n11625), .A2(n11624), .B1(n11623), .B2(n11622), .ZN(
        n11916) );
  AOI22_X1 U14743 ( .A1(n9834), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11629) );
  AOI22_X1 U14744 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17139), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11628) );
  AOI22_X1 U14745 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9832), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11627) );
  AOI22_X1 U14746 ( .A1(n17094), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11626) );
  NAND4_X1 U14747 ( .A1(n11629), .A2(n11628), .A3(n11627), .A4(n11626), .ZN(
        n11636) );
  AOI22_X1 U14748 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n15657), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11634) );
  AOI22_X1 U14749 ( .A1(n9831), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11633) );
  INV_X2 U14750 ( .A(n11715), .ZN(n17128) );
  AOI22_X1 U14751 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17128), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11632) );
  AOI22_X1 U14752 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11631) );
  NAND4_X1 U14753 ( .A1(n11634), .A2(n11633), .A3(n11632), .A4(n11631), .ZN(
        n11635) );
  AOI22_X1 U14754 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(n18626), .B2(n18762), .ZN(
        n11642) );
  OAI22_X1 U14755 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18154), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n11639), .ZN(n11645) );
  NOR2_X1 U14756 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18154), .ZN(
        n11640) );
  NAND2_X1 U14757 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11639), .ZN(
        n11646) );
  AOI22_X1 U14758 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n11645), .B1(
        n11640), .B2(n11646), .ZN(n11756) );
  OAI21_X1 U14759 ( .B1(n11643), .B2(n11642), .A(n11756), .ZN(n11641) );
  OAI21_X1 U14760 ( .B1(n18392), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n11644), .ZN(n11751) );
  INV_X1 U14761 ( .A(n11751), .ZN(n11650) );
  XOR2_X1 U14762 ( .A(n11752), .B(n11644), .Z(n11649) );
  INV_X1 U14763 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15680) );
  AOI21_X1 U14764 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n11646), .A(
        n11645), .ZN(n11647) );
  INV_X1 U14765 ( .A(n11647), .ZN(n11648) );
  INV_X1 U14766 ( .A(n18631), .ZN(n16488) );
  AOI21_X1 U14767 ( .B1(n11754), .B2(n11650), .A(n16488), .ZN(n18786) );
  AOI22_X1 U14768 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11654) );
  AOI22_X1 U14769 ( .A1(n9824), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17107), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11653) );
  AOI22_X1 U14770 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9832), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11652) );
  AOI22_X1 U14771 ( .A1(n9831), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11651) );
  NAND4_X1 U14772 ( .A1(n11654), .A2(n11653), .A3(n11652), .A4(n11651), .ZN(
        n11661) );
  AOI22_X1 U14773 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n15657), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11659) );
  AOI22_X1 U14774 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17094), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11658) );
  AOI22_X1 U14775 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9834), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11657) );
  AOI22_X1 U14776 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11716), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11656) );
  NAND4_X1 U14777 ( .A1(n11659), .A2(n11658), .A3(n11657), .A4(n11656), .ZN(
        n11660) );
  XOR2_X1 U14778 ( .A(n18163), .B(n11701), .Z(n11894) );
  AOI22_X1 U14779 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11671) );
  INV_X1 U14780 ( .A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n21041) );
  AOI22_X1 U14781 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11663) );
  AOI22_X1 U14782 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11544), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11662) );
  OAI211_X1 U14783 ( .C1(n17004), .C2(n21041), .A(n11663), .B(n11662), .ZN(
        n11669) );
  AOI22_X1 U14784 ( .A1(n9831), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17139), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11667) );
  AOI22_X1 U14785 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9832), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11666) );
  AOI22_X1 U14786 ( .A1(n9834), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17094), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11665) );
  AOI22_X1 U14787 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17128), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11664) );
  NAND4_X1 U14788 ( .A1(n11667), .A2(n11666), .A3(n11665), .A4(n11664), .ZN(
        n11668) );
  AOI211_X1 U14789 ( .C1(n17146), .C2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n11669), .B(n11668), .ZN(n11670) );
  NAND2_X1 U14790 ( .A1(n18160), .A2(n18795), .ZN(n11731) );
  INV_X1 U14791 ( .A(n11731), .ZN(n11740) );
  AOI22_X1 U14792 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17139), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11676) );
  AOI22_X1 U14793 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11675) );
  AOI22_X1 U14794 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9831), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11674) );
  AOI22_X1 U14795 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11673) );
  NAND4_X1 U14796 ( .A1(n11676), .A2(n11675), .A3(n11674), .A4(n11673), .ZN(
        n11682) );
  AOI22_X1 U14797 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11680) );
  AOI22_X1 U14798 ( .A1(n9834), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11679) );
  AOI22_X1 U14799 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11678) );
  AOI22_X1 U14800 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11716), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11677) );
  NAND4_X1 U14801 ( .A1(n11680), .A2(n11679), .A3(n11678), .A4(n11677), .ZN(
        n11681) );
  AOI22_X1 U14802 ( .A1(n9834), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11544), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11691) );
  AOI22_X1 U14803 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17140), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11690) );
  AOI22_X1 U14804 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9831), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11683) );
  OAI21_X1 U14805 ( .B1(n11684), .B2(n21009), .A(n11683), .ZN(n11689) );
  AOI22_X1 U14806 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n15657), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11688) );
  AOI22_X1 U14807 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17094), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11687) );
  AOI22_X1 U14808 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11686) );
  AOI22_X1 U14809 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11716), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11685) );
  AOI22_X1 U14810 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9834), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11695) );
  AOI22_X1 U14811 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11694) );
  AOI22_X1 U14812 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17128), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11693) );
  AOI22_X1 U14813 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17107), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11692) );
  AOI22_X1 U14814 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n15657), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11700) );
  AOI22_X1 U14815 ( .A1(n9831), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17094), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11699) );
  AOI22_X1 U14816 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9824), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11698) );
  AOI22_X1 U14817 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11716), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11697) );
  AOI22_X1 U14818 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__7__SCAN_IN), .B2(n17108), .ZN(n11713) );
  AOI22_X1 U14819 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n17128), .ZN(n11712) );
  INV_X1 U14820 ( .A(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11704) );
  AOI22_X1 U14821 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17123), .B1(
        n17054), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11703) );
  OAI21_X1 U14822 ( .B1(n11704), .B2(n10310), .A(n11703), .ZN(n11710) );
  AOI22_X1 U14823 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11708) );
  AOI22_X1 U14824 ( .A1(n9831), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n9832), .ZN(n11707) );
  AOI22_X1 U14825 ( .A1(n9824), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n17094), .ZN(n11706) );
  AOI22_X1 U14826 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n17146), .B1(
        n11716), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11705) );
  NAND4_X1 U14827 ( .A1(n11708), .A2(n11707), .A3(n11706), .A4(n11705), .ZN(
        n11709) );
  NAND3_X2 U14828 ( .A1(n11713), .A2(n11712), .A3(n11711), .ZN(n17160) );
  AOI22_X1 U14829 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11725) );
  AOI22_X1 U14830 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17107), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11724) );
  INV_X1 U14831 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17179) );
  AOI22_X1 U14832 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11714) );
  OAI21_X1 U14833 ( .B1(n11715), .B2(n17179), .A(n11714), .ZN(n11722) );
  AOI22_X1 U14834 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15657), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11720) );
  AOI22_X1 U14835 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17139), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11719) );
  AOI22_X1 U14836 ( .A1(n9831), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9834), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11718) );
  AOI22_X1 U14837 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11716), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11717) );
  NAND4_X1 U14838 ( .A1(n11720), .A2(n11719), .A3(n11718), .A4(n11717), .ZN(
        n11721) );
  AOI211_X1 U14839 ( .C1(n17153), .C2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A(
        n11722), .B(n11721), .ZN(n11723) );
  NAND3_X1 U14840 ( .A1(n11725), .A2(n11724), .A3(n11723), .ZN(n11729) );
  NAND2_X1 U14841 ( .A1(n18167), .A2(n18171), .ZN(n18589) );
  NAND2_X1 U14842 ( .A1(n17193), .A2(n17201), .ZN(n11741) );
  AOI21_X1 U14843 ( .B1(n17160), .B2(n11741), .A(n18175), .ZN(n11727) );
  AOI21_X1 U14844 ( .B1(n11728), .B2(n18160), .A(n11727), .ZN(n11744) );
  INV_X1 U14845 ( .A(n18175), .ZN(n14313) );
  NAND2_X1 U14846 ( .A1(n17160), .A2(n18160), .ZN(n11747) );
  NOR4_X2 U14847 ( .A1(n14313), .A2(n11729), .A3(n11747), .A4(n11741), .ZN(
        n11750) );
  INV_X1 U14848 ( .A(n11750), .ZN(n15672) );
  AOI21_X2 U14849 ( .B1(n11730), .B2(n11744), .A(n11898), .ZN(n16490) );
  INV_X1 U14850 ( .A(n18589), .ZN(n11732) );
  NAND2_X1 U14851 ( .A1(n11733), .A2(n11732), .ZN(n14312) );
  INV_X1 U14852 ( .A(n14312), .ZN(n11735) );
  NAND2_X1 U14853 ( .A1(n18163), .A2(n18160), .ZN(n15766) );
  INV_X1 U14854 ( .A(n15766), .ZN(n11734) );
  NAND3_X1 U14855 ( .A1(n11735), .A2(n17160), .A3(n11734), .ZN(n11736) );
  INV_X1 U14856 ( .A(n11737), .ZN(n16505) );
  NOR3_X1 U14857 ( .A1(n11738), .A2(n18163), .A3(n16505), .ZN(n11749) );
  NOR2_X1 U14858 ( .A1(n18178), .A2(n17193), .ZN(n18616) );
  OAI21_X1 U14859 ( .B1(n18188), .B2(n18616), .A(n11739), .ZN(n11896) );
  AOI21_X1 U14860 ( .B1(n18175), .B2(n17201), .A(n11740), .ZN(n11743) );
  INV_X1 U14861 ( .A(n11741), .ZN(n11742) );
  AOI21_X1 U14862 ( .B1(n18167), .B2(n11743), .A(n11742), .ZN(n11746) );
  INV_X1 U14863 ( .A(n11744), .ZN(n11745) );
  AOI211_X1 U14864 ( .C1(n18171), .C2(n11747), .A(n11746), .B(n11745), .ZN(
        n11897) );
  OAI211_X1 U14865 ( .C1(n18171), .C2(n11748), .A(n11896), .B(n11897), .ZN(
        n15671) );
  NOR2_X1 U14866 ( .A1(n11752), .A2(n11751), .ZN(n11755) );
  NAND3_X1 U14867 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .A3(n18757), .ZN(n18651) );
  INV_X1 U14868 ( .A(n17321), .ZN(n16383) );
  NOR2_X1 U14869 ( .A1(n11916), .A2(n17726), .ZN(n11797) );
  INV_X1 U14870 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16552) );
  NAND2_X1 U14871 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17775) );
  NAND2_X1 U14872 ( .A1(n17758), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17742) );
  NAND2_X1 U14873 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17719) );
  NAND2_X1 U14874 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16749) );
  NOR2_X1 U14875 ( .A1(n17719), .A2(n16749), .ZN(n17681) );
  NAND3_X1 U14876 ( .A1(n17716), .A2(n17681), .A3(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17660) );
  NAND2_X1 U14877 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17662) );
  NAND2_X1 U14878 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17619) );
  NAND2_X1 U14879 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17589) );
  NAND2_X1 U14880 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17549) );
  NAND2_X1 U14881 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17506) );
  INV_X1 U14882 ( .A(n17468), .ZN(n17460) );
  NAND3_X1 U14883 ( .A1(n17460), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16359) );
  NOR2_X1 U14884 ( .A1(n16552), .A2(n16359), .ZN(n11758) );
  INV_X1 U14885 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17812) );
  INV_X1 U14886 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18809) );
  NOR2_X1 U14887 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18809), .ZN(n17652) );
  NAND2_X1 U14888 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18146) );
  NAND2_X1 U14889 ( .A1(n18748), .A2(n18146), .ZN(n18801) );
  NAND2_X1 U14890 ( .A1(n18757), .A2(n18809), .ZN(n18798) );
  AOI21_X1 U14891 ( .B1(n18798), .B2(n18146), .A(n18770), .ZN(n18157) );
  INV_X1 U14892 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n16507) );
  NOR3_X1 U14893 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n16507), .ZN(n18211) );
  OAI21_X1 U14894 ( .B1(n17812), .B2(n17603), .A(n18499), .ZN(n17467) );
  NAND2_X1 U14895 ( .A1(n11758), .A2(n17467), .ZN(n11763) );
  NOR2_X1 U14896 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n11763), .ZN(
        n16350) );
  NAND3_X1 U14897 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A3(n16520), .ZN(n16517) );
  NOR2_X1 U14898 ( .A1(n11758), .A2(n18499), .ZN(n16370) );
  INV_X1 U14899 ( .A(n17817), .ZN(n17774) );
  AOI211_X1 U14900 ( .C1(n17652), .C2(n16517), .A(n16370), .B(n17774), .ZN(
        n16363) );
  OAI21_X1 U14901 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n17603), .A(
        n16363), .ZN(n16351) );
  OAI21_X1 U14902 ( .B1(n16350), .B2(n16351), .A(
        P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11762) );
  NAND2_X1 U14903 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16364) );
  INV_X1 U14904 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11759) );
  NOR2_X1 U14905 ( .A1(n16364), .A2(n11759), .ZN(n15755) );
  NAND2_X1 U14906 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17824) );
  NOR2_X1 U14907 ( .A1(n17871), .A2(n17824), .ZN(n17512) );
  NAND2_X1 U14908 ( .A1(n17512), .A2(n11760), .ZN(n16375) );
  NOR2_X1 U14909 ( .A1(n11609), .A2(n16375), .ZN(n17464) );
  NAND3_X1 U14910 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15755), .A3(
        n17464), .ZN(n11761) );
  XOR2_X1 U14911 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n11761), .Z(
        n11914) );
  NAND2_X1 U14912 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n17715) );
  NAND2_X1 U14913 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16360), .ZN(
        n16349) );
  INV_X1 U14914 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18729) );
  NOR2_X1 U14915 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18810) );
  INV_X1 U14916 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18799) );
  NOR2_X1 U14917 ( .A1(n18729), .A2(n18138), .ZN(n11908) );
  INV_X1 U14918 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16536) );
  NOR3_X1 U14919 ( .A1(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n16536), .A3(
        n11763), .ZN(n11764) );
  AOI211_X1 U14920 ( .C1(n17655), .C2(n16837), .A(n11908), .B(n11764), .ZN(
        n11795) );
  NAND2_X1 U14921 ( .A1(n11776), .A2(n15768), .ZN(n11775) );
  INV_X1 U14922 ( .A(n11765), .ZN(n17340) );
  NAND2_X1 U14923 ( .A1(n11775), .A2(n17340), .ZN(n11771) );
  INV_X1 U14924 ( .A(n11771), .ZN(n11766) );
  NOR2_X1 U14925 ( .A1(n17334), .A2(n11766), .ZN(n11770) );
  NAND2_X1 U14926 ( .A1(n11770), .A2(n11767), .ZN(n11769) );
  NOR2_X1 U14927 ( .A1(n17327), .A2(n11769), .ZN(n17745) );
  NAND2_X1 U14928 ( .A1(n17745), .A2(n17747), .ZN(n11768) );
  NOR2_X1 U14929 ( .A1(n17321), .A2(n11768), .ZN(n11791) );
  XOR2_X1 U14930 ( .A(n17321), .B(n11768), .Z(n11787) );
  XOR2_X1 U14931 ( .A(n17327), .B(n11769), .Z(n11783) );
  AND2_X1 U14932 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n11783), .ZN(
        n11784) );
  XNOR2_X1 U14933 ( .A(n17331), .B(n11770), .ZN(n11781) );
  AND2_X1 U14934 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n11781), .ZN(
        n11782) );
  XNOR2_X1 U14935 ( .A(n17334), .B(n11771), .ZN(n11779) );
  AND2_X1 U14936 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n11779), .ZN(
        n11780) );
  OAI21_X1 U14937 ( .B1(n11773), .B2(n11772), .A(n11771), .ZN(n11777) );
  AND2_X1 U14938 ( .A1(n11777), .A2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11778) );
  NOR2_X1 U14939 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15768), .ZN(
        n17814) );
  NAND2_X1 U14940 ( .A1(n17814), .A2(n11774), .ZN(n17805) );
  OAI211_X1 U14941 ( .C1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n11776), .A(
        n11775), .B(n17805), .ZN(n17796) );
  XNOR2_X1 U14942 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n11777), .ZN(
        n17795) );
  NOR2_X1 U14943 ( .A1(n17796), .A2(n17795), .ZN(n17794) );
  NOR2_X1 U14944 ( .A1(n11778), .A2(n17794), .ZN(n17785) );
  XNOR2_X1 U14945 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n11779), .ZN(
        n17784) );
  NOR2_X1 U14946 ( .A1(n17785), .A2(n17784), .ZN(n17783) );
  NOR2_X1 U14947 ( .A1(n11780), .A2(n17783), .ZN(n17771) );
  XNOR2_X1 U14948 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n11781), .ZN(
        n17770) );
  NOR2_X1 U14949 ( .A1(n17771), .A2(n17770), .ZN(n17769) );
  NOR2_X1 U14950 ( .A1(n11782), .A2(n17769), .ZN(n17763) );
  XNOR2_X1 U14951 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n11783), .ZN(
        n17762) );
  NOR2_X1 U14952 ( .A1(n17763), .A2(n17762), .ZN(n17761) );
  NOR2_X1 U14953 ( .A1(n11784), .A2(n17761), .ZN(n17744) );
  INV_X1 U14954 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18064) );
  INV_X1 U14955 ( .A(n17747), .ZN(n17746) );
  XOR2_X1 U14956 ( .A(n17746), .B(n17745), .Z(n11785) );
  AOI222_X1 U14957 ( .A1(n17744), .A2(n18064), .B1(n17744), .B2(n11785), .C1(
        n18064), .C2(n11785), .ZN(n11788) );
  NOR2_X1 U14958 ( .A1(n11787), .A2(n11788), .ZN(n17731) );
  NOR2_X1 U14959 ( .A1(n17731), .A2(n18071), .ZN(n11786) );
  NAND2_X1 U14960 ( .A1(n11791), .A2(n11786), .ZN(n11792) );
  INV_X1 U14961 ( .A(n11786), .ZN(n11790) );
  AND2_X1 U14962 ( .A1(n11788), .A2(n11787), .ZN(n17732) );
  AOI21_X1 U14963 ( .B1(n11791), .B2(n11790), .A(n17732), .ZN(n11789) );
  OAI21_X1 U14964 ( .B1(n11791), .B2(n11790), .A(n11789), .ZN(n17718) );
  NAND2_X1 U14965 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17718), .ZN(
        n17717) );
  NAND3_X1 U14966 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n17463), .A3(
        n15755), .ZN(n11793) );
  XOR2_X1 U14967 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n11793), .Z(
        n11911) );
  NAND2_X1 U14968 ( .A1(n18163), .A2(n11794), .ZN(n17822) );
  NAND3_X1 U14969 ( .A1(n10316), .A2(n11795), .A3(n10318), .ZN(n11796) );
  OR2_X1 U14970 ( .A1(n11797), .A2(n11796), .ZN(P3_U2799) );
  NAND2_X1 U14971 ( .A1(n11799), .A2(n11798), .ZN(n15410) );
  INV_X1 U14972 ( .A(n11800), .ZN(n11806) );
  INV_X1 U14973 ( .A(n11804), .ZN(n15599) );
  NAND2_X1 U14974 ( .A1(n15427), .A2(n11807), .ZN(n15417) );
  NAND2_X1 U14975 ( .A1(n9910), .A2(n11808), .ZN(n15418) );
  NOR2_X1 U14976 ( .A1(n11813), .A2(n11812), .ZN(n11814) );
  NAND2_X1 U14977 ( .A1(n11828), .A2(n10996), .ZN(n11827) );
  OAI21_X1 U14978 ( .B1(n10000), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n11817), .ZN(n11838) );
  INV_X1 U14979 ( .A(n11838), .ZN(n11818) );
  INV_X1 U14980 ( .A(n11819), .ZN(n11820) );
  NAND2_X1 U14981 ( .A1(n9907), .A2(n11820), .ZN(n11821) );
  NAND2_X1 U14982 ( .A1(n15228), .A2(n11821), .ZN(n15239) );
  AOI21_X1 U14983 ( .B1(n13327), .B2(n11822), .A(n9936), .ZN(n13325) );
  OAI22_X1 U14984 ( .A1(n19779), .A2(n18878), .B1(n13327), .B2(n16243), .ZN(
        n11823) );
  AOI21_X1 U14985 ( .B1(n16234), .B2(n13325), .A(n11823), .ZN(n11824) );
  NAND2_X1 U14986 ( .A1(n11827), .A2(n11826), .ZN(P2_U2993) );
  NAND2_X1 U14987 ( .A1(n11828), .A2(n16283), .ZN(n11841) );
  INV_X1 U14988 ( .A(n15298), .ZN(n11829) );
  OAI21_X1 U14989 ( .B1(n11830), .B2(n15316), .A(n11829), .ZN(n13329) );
  INV_X1 U14990 ( .A(n13329), .ZN(n15312) );
  NOR3_X1 U14991 ( .A1(n15493), .A2(n15494), .A3(n11831), .ZN(n11832) );
  AOI21_X1 U14992 ( .B1(P2_REIP_REG_21__SCAN_IN), .B2(n19138), .A(n11832), 
        .ZN(n11833) );
  OAI21_X1 U14993 ( .B1(n15239), .B2(n16272), .A(n11833), .ZN(n11836) );
  NOR2_X1 U14994 ( .A1(n11834), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11835) );
  AOI211_X1 U14995 ( .C1(n16280), .C2(n15312), .A(n11836), .B(n11835), .ZN(
        n11837) );
  OAI21_X1 U14996 ( .B1(n11838), .B2(n15637), .A(n11837), .ZN(n11839) );
  NAND2_X1 U14997 ( .A1(n11841), .A2(n11840), .ZN(P2_U3025) );
  NOR2_X2 U14998 ( .A1(n11890), .A2(n11842), .ZN(n14481) );
  XNOR2_X1 U14999 ( .A(n14481), .B(n11858), .ZN(n11864) );
  NAND2_X1 U15000 ( .A1(n11864), .A2(n11843), .ZN(n11863) );
  NAND2_X1 U15001 ( .A1(n11844), .A2(n14469), .ZN(n11849) );
  INV_X1 U15002 ( .A(n11845), .ZN(n11847) );
  NAND2_X1 U15003 ( .A1(n11847), .A2(n11846), .ZN(n11848) );
  NAND2_X1 U15004 ( .A1(n11865), .A2(n16283), .ZN(n11862) );
  NAND2_X1 U15005 ( .A1(n11852), .A2(n11851), .ZN(n11853) );
  NAND2_X1 U15006 ( .A1(n11854), .A2(n11853), .ZN(n14555) );
  NAND2_X1 U15007 ( .A1(P2_REIP_REG_30__SCAN_IN), .A2(n16261), .ZN(n11866) );
  OR3_X1 U15008 ( .A1(n15447), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n15434), .ZN(n11855) );
  OAI211_X1 U15009 ( .C1(n16271), .C2(n14555), .A(n11866), .B(n11855), .ZN(
        n11856) );
  AOI21_X1 U15010 ( .B1(n14564), .B2(n16285), .A(n11856), .ZN(n11857) );
  OAI21_X1 U15011 ( .B1(n11859), .B2(n11858), .A(n11857), .ZN(n11860) );
  NAND3_X1 U15012 ( .A1(n11863), .A2(n11862), .A3(n11861), .ZN(P2_U3016) );
  NAND2_X1 U15013 ( .A1(n11864), .A2(n16228), .ZN(n11872) );
  NAND2_X1 U15014 ( .A1(n11865), .A2(n10996), .ZN(n11871) );
  NAND2_X1 U15015 ( .A1(n14564), .A2(n19146), .ZN(n11867) );
  OAI211_X1 U15016 ( .C1(n16243), .C2(n11869), .A(n11867), .B(n11866), .ZN(
        n11868) );
  INV_X1 U15017 ( .A(n11868), .ZN(n11870) );
  XNOR2_X1 U15018 ( .A(n14473), .B(n11869), .ZN(n16047) );
  NAND3_X1 U15019 ( .A1(n11872), .A2(n11871), .A3(n10301), .ZN(P2_U2984) );
  INV_X1 U15020 ( .A(n11875), .ZN(n11874) );
  NAND2_X1 U15021 ( .A1(n11876), .A2(n11874), .ZN(n11878) );
  NAND2_X1 U15022 ( .A1(n15351), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15352) );
  NAND2_X1 U15023 ( .A1(n15352), .A2(n11878), .ZN(n11881) );
  XNOR2_X1 U15024 ( .A(n11879), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11880) );
  XNOR2_X1 U15025 ( .A(n11881), .B(n11880), .ZN(n14519) );
  NOR2_X1 U15026 ( .A1(n11882), .A2(n11883), .ZN(n11884) );
  NAND2_X1 U15027 ( .A1(P2_REIP_REG_28__SCAN_IN), .A2(n16261), .ZN(n14508) );
  NAND2_X1 U15028 ( .A1(n19137), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11885) );
  OAI211_X1 U15029 ( .C1(n16071), .C2(n19157), .A(n14508), .B(n11885), .ZN(
        n11888) );
  OAI21_X1 U15030 ( .B1(n9940), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n11886), .ZN(n14485) );
  NOR2_X1 U15031 ( .A1(n14485), .A2(n19150), .ZN(n11887) );
  NOR2_X1 U15032 ( .A1(n11888), .A2(n11887), .ZN(n11893) );
  INV_X1 U15033 ( .A(n11890), .ZN(n11889) );
  NAND2_X1 U15034 ( .A1(n11890), .A2(n10947), .ZN(n14502) );
  AND2_X1 U15035 ( .A1(n14516), .A2(n14502), .ZN(n11891) );
  OAI211_X1 U15036 ( .C1(n14519), .C2(n19142), .A(n11893), .B(n11892), .ZN(
        P2_U2986) );
  INV_X2 U15037 ( .A(n18807), .ZN(n18739) );
  NAND2_X2 U15038 ( .A1(n18739), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18732) );
  INV_X1 U15039 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n16480) );
  INV_X1 U15040 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18677) );
  NAND2_X1 U15041 ( .A1(n16480), .A2(n18677), .ZN(n16487) );
  NAND3_X1 U15042 ( .A1(n18674), .A2(n18732), .A3(n16487), .ZN(n18668) );
  NAND2_X1 U15043 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18803) );
  INV_X1 U15044 ( .A(n18803), .ZN(n18796) );
  AOI21_X1 U15045 ( .B1(n18668), .B2(n11894), .A(n18796), .ZN(n16489) );
  INV_X1 U15046 ( .A(n16489), .ZN(n11895) );
  NOR3_X1 U15047 ( .A1(n11900), .A2(n16488), .A3(n11895), .ZN(n11899) );
  OAI211_X1 U15048 ( .C1(n11898), .C2(n9882), .A(n11897), .B(n11896), .ZN(
        n15675) );
  AOI211_X1 U15049 ( .C1(n18788), .C2(n11900), .A(n11899), .B(n15675), .ZN(
        n11902) );
  NAND4_X1 U15050 ( .A1(n18786), .A2(n18167), .A3(n18795), .A4(n17193), .ZN(
        n11901) );
  NAND2_X1 U15051 ( .A1(n9828), .A2(n18136), .ZN(n18144) );
  NAND3_X1 U15052 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15755), .A3(
        n18758), .ZN(n11903) );
  INV_X1 U15053 ( .A(n18606), .ZN(n18629) );
  AOI21_X1 U15054 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18053) );
  NAND3_X1 U15055 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18073) );
  NOR3_X1 U15056 ( .A1(n18064), .A2(n18071), .A3(n18073), .ZN(n18058) );
  NAND2_X1 U15057 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18058), .ZN(
        n17949) );
  NOR2_X1 U15058 ( .A1(n18053), .A2(n17949), .ZN(n17938) );
  NAND2_X1 U15059 ( .A1(n17613), .A2(n17938), .ZN(n17864) );
  INV_X1 U15060 ( .A(n18600), .ZN(n18603) );
  OAI21_X1 U15061 ( .B1(n15672), .B2(n15671), .A(n18603), .ZN(n18594) );
  INV_X1 U15062 ( .A(n18615), .ZN(n18033) );
  NAND2_X1 U15063 ( .A1(n18033), .A2(n18593), .ZN(n18113) );
  OAI21_X1 U15064 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18594), .A(
        n18113), .ZN(n18106) );
  NOR2_X1 U15065 ( .A1(n18122), .A2(n21073), .ZN(n18050) );
  NAND2_X1 U15066 ( .A1(n18058), .A2(n18050), .ZN(n18036) );
  NOR2_X1 U15067 ( .A1(n18057), .A2(n18036), .ZN(n17939) );
  NAND2_X1 U15068 ( .A1(n17613), .A2(n17939), .ZN(n17920) );
  OAI22_X1 U15069 ( .A1(n18629), .A2(n17864), .B1(n18106), .B2(n17920), .ZN(
        n15685) );
  NAND2_X1 U15070 ( .A1(n17512), .A2(n15685), .ZN(n17846) );
  NOR4_X1 U15071 ( .A1(n17825), .A2(n11903), .A3(n18128), .A4(n17846), .ZN(
        n11910) );
  INV_X1 U15072 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n20889) );
  NAND2_X1 U15073 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17939), .ZN(
        n17964) );
  INV_X1 U15074 ( .A(n17964), .ZN(n18032) );
  NAND2_X1 U15075 ( .A1(n17613), .A2(n18032), .ZN(n17940) );
  NOR3_X1 U15076 ( .A1(n16375), .A2(n20889), .A3(n17940), .ZN(n11905) );
  OAI21_X1 U15077 ( .B1(n16375), .B2(n17920), .A(n18594), .ZN(n11904) );
  INV_X1 U15078 ( .A(n17864), .ZN(n17879) );
  NAND2_X1 U15079 ( .A1(n17512), .A2(n17879), .ZN(n17845) );
  OAI21_X1 U15080 ( .B1(n17825), .B2(n17845), .A(n18606), .ZN(n17828) );
  OAI211_X1 U15081 ( .C1(n18033), .C2(n11905), .A(n11904), .B(n17828), .ZN(
        n15683) );
  NAND2_X1 U15082 ( .A1(n18136), .A2(n18091), .ZN(n18055) );
  OAI21_X1 U15083 ( .B1(n15755), .B2(n18055), .A(n18121), .ZN(n11906) );
  AOI21_X1 U15084 ( .B1(n18136), .B2(n15683), .A(n11906), .ZN(n15757) );
  OAI22_X1 U15085 ( .A1(n15757), .A2(n18758), .B1(n11907), .B2(n18055), .ZN(
        n11909) );
  INV_X1 U15086 ( .A(n11912), .ZN(n11915) );
  NAND2_X1 U15087 ( .A1(n17321), .A2(n18135), .ZN(n17979) );
  OAI21_X1 U15088 ( .B1(n11916), .B2(n18045), .A(n10294), .ZN(P3_U2831) );
  NAND2_X1 U15089 ( .A1(n10425), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11917) );
  NAND2_X1 U15090 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19387) );
  XNOR2_X1 U15091 ( .A(n19387), .B(n19822), .ZN(n19294) );
  NOR2_X1 U15092 ( .A1(n19294), .A2(n19810), .ZN(n11918) );
  AOI21_X1 U15093 ( .B1(n11936), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11918), .ZN(n11919) );
  NOR2_X1 U15094 ( .A1(n10425), .A2(n19859), .ZN(n13580) );
  INV_X1 U15095 ( .A(n11938), .ZN(n11924) );
  NAND2_X1 U15096 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19841), .ZN(
        n19623) );
  NAND2_X1 U15097 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19831), .ZN(
        n19577) );
  NAND2_X1 U15098 ( .A1(n19623), .A2(n19577), .ZN(n19628) );
  INV_X1 U15099 ( .A(n19628), .ZN(n11922) );
  NAND2_X1 U15100 ( .A1(n11936), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11921) );
  OAI21_X1 U15101 ( .B1(n11922), .B2(n19810), .A(n11921), .ZN(n11923) );
  NOR2_X1 U15102 ( .A1(n19810), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11925) );
  AOI21_X1 U15103 ( .B1(n11936), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n11925), .ZN(n11926) );
  NAND2_X1 U15104 ( .A1(n13583), .A2(n11928), .ZN(n11929) );
  INV_X1 U15105 ( .A(n11930), .ZN(n11931) );
  NAND2_X1 U15106 ( .A1(n11932), .A2(n11931), .ZN(n13688) );
  INV_X1 U15107 ( .A(n19387), .ZN(n19511) );
  AND2_X1 U15108 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19665) );
  NAND2_X1 U15109 ( .A1(n19511), .A2(n19665), .ZN(n19667) );
  OAI21_X1 U15110 ( .B1(n19387), .B2(n19822), .A(n11933), .ZN(n11934) );
  AND3_X1 U15111 ( .A1(n19813), .A2(n19667), .A3(n11934), .ZN(n11935) );
  AOI21_X1 U15112 ( .B1(n11936), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11935), .ZN(n11937) );
  INV_X1 U15113 ( .A(n11944), .ZN(n11941) );
  AND2_X1 U15114 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n10425), .ZN(
        n11940) );
  AND2_X1 U15115 ( .A1(n13688), .A2(n11943), .ZN(n11942) );
  INV_X1 U15116 ( .A(n11943), .ZN(n11946) );
  XNOR2_X1 U15117 ( .A(n11945), .B(n11944), .ZN(n13687) );
  INV_X1 U15118 ( .A(n12193), .ZN(n12154) );
  NOR2_X2 U15119 ( .A1(n13680), .A2(n19207), .ZN(n13727) );
  AND2_X1 U15120 ( .A1(n13814), .A2(n13815), .ZN(n11950) );
  NAND2_X1 U15121 ( .A1(n13727), .A2(n11950), .ZN(n13781) );
  NOR2_X1 U15122 ( .A1(n13781), .A2(n11951), .ZN(n13868) );
  INV_X1 U15123 ( .A(n12086), .ZN(n12048) );
  AOI22_X1 U15124 ( .A1(n10577), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10654), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11955) );
  AOI22_X1 U15125 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12085), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11954) );
  OAI211_X1 U15126 ( .C1(n12048), .C2(n19555), .A(n11955), .B(n11954), .ZN(
        n11964) );
  AOI22_X1 U15127 ( .A1(n12050), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12049), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11957) );
  AOI22_X1 U15128 ( .A1(n12051), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13807), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11956) );
  NAND2_X1 U15129 ( .A1(n11957), .A2(n11956), .ZN(n11963) );
  INV_X1 U15130 ( .A(n12064), .ZN(n12057) );
  AOI22_X1 U15131 ( .A1(n10626), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10588), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11959) );
  AOI22_X1 U15132 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12065), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11958) );
  OAI211_X1 U15133 ( .C1(n12057), .C2(n21089), .A(n11959), .B(n11958), .ZN(
        n11962) );
  INV_X1 U15134 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11960) );
  OAI22_X1 U15135 ( .A1(n11975), .A2(n20926), .B1(n10767), .B2(n11960), .ZN(
        n11961) );
  NOR4_X1 U15136 ( .A1(n11964), .A2(n11963), .A3(n11962), .A4(n11961), .ZN(
        n14129) );
  AOI22_X1 U15137 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n10577), .B1(
        n10654), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11966) );
  AOI22_X1 U15138 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10574), .B1(
        n12085), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11965) );
  OAI211_X1 U15139 ( .C1(n11967), .C2(n12048), .A(n11966), .B(n11965), .ZN(
        n11974) );
  OAI22_X1 U15140 ( .A1(n12078), .A2(n11969), .B1(n12076), .B2(n11968), .ZN(
        n11973) );
  INV_X1 U15141 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11971) );
  OAI22_X1 U15142 ( .A1(n11971), .A2(n12081), .B1(n12080), .B2(n11970), .ZN(
        n11972) );
  NOR3_X1 U15143 ( .A1(n11974), .A2(n11973), .A3(n11972), .ZN(n11982) );
  INV_X1 U15144 ( .A(n11975), .ZN(n12035) );
  AOI22_X1 U15145 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n11278), .B1(
        n12035), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11981) );
  AOI22_X1 U15146 ( .A1(n10626), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n10588), .ZN(n11980) );
  INV_X1 U15147 ( .A(n12066), .ZN(n12039) );
  INV_X1 U15148 ( .A(n12065), .ZN(n12037) );
  OAI22_X1 U15149 ( .A1(n12039), .A2(n11977), .B1(n12037), .B2(n11976), .ZN(
        n11978) );
  AOI21_X1 U15150 ( .B1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n12064), .A(
        n11978), .ZN(n11979) );
  NAND4_X1 U15151 ( .A1(n11982), .A2(n11981), .A3(n11980), .A4(n11979), .ZN(
        n14209) );
  AOI22_X1 U15152 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10654), .B1(
        n10577), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11984) );
  AOI22_X1 U15153 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10574), .B1(
        n12085), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11983) );
  OAI211_X1 U15154 ( .C1(n11985), .C2(n12048), .A(n11984), .B(n11983), .ZN(
        n11995) );
  AOI22_X1 U15155 ( .A1(n12050), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12049), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11987) );
  AOI22_X1 U15156 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n12051), .B1(
        n13807), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11986) );
  NAND2_X1 U15157 ( .A1(n11987), .A2(n11986), .ZN(n11994) );
  AOI22_X1 U15158 ( .A1(n10626), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__4__SCAN_IN), .B2(n10588), .ZN(n11989) );
  AOI22_X1 U15159 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12065), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11988) );
  OAI211_X1 U15160 ( .C1(n12057), .C2(n10721), .A(n11989), .B(n11988), .ZN(
        n11993) );
  INV_X1 U15161 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11991) );
  OAI22_X1 U15162 ( .A1(n11991), .A2(n10767), .B1(n11975), .B2(n11990), .ZN(
        n11992) );
  NOR4_X1 U15163 ( .A1(n11995), .A2(n11994), .A3(n11993), .A4(n11992), .ZN(
        n15246) );
  AOI22_X1 U15164 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10654), .B1(
        n10577), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11997) );
  AOI22_X1 U15165 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12085), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11996) );
  OAI211_X1 U15166 ( .C1(n11998), .C2(n12048), .A(n11997), .B(n11996), .ZN(
        n12008) );
  OAI22_X1 U15167 ( .A1(n11999), .A2(n11975), .B1(n10767), .B2(n10608), .ZN(
        n12007) );
  AOI22_X1 U15168 ( .A1(n10626), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__3__SCAN_IN), .B2(n10588), .ZN(n12001) );
  AOI22_X1 U15169 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12065), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12000) );
  OAI211_X1 U15170 ( .C1(n12057), .C2(n12002), .A(n12001), .B(n12000), .ZN(
        n12006) );
  AOI22_X1 U15171 ( .A1(n12050), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12049), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12004) );
  AOI22_X1 U15172 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n12051), .B1(
        n13807), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12003) );
  NAND2_X1 U15173 ( .A1(n12004), .A2(n12003), .ZN(n12005) );
  OR4_X1 U15174 ( .A1(n12008), .A2(n12007), .A3(n12006), .A4(n12005), .ZN(
        n15251) );
  INV_X1 U15175 ( .A(n15251), .ZN(n12023) );
  AOI22_X1 U15176 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10654), .B1(
        n10577), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12010) );
  AOI22_X1 U15177 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10574), .B1(
        n12085), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12009) );
  OAI211_X1 U15178 ( .C1(n12011), .C2(n12048), .A(n12010), .B(n12009), .ZN(
        n12022) );
  AOI22_X1 U15179 ( .A1(n12050), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12049), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12013) );
  AOI22_X1 U15180 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n12051), .B1(
        n13807), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12012) );
  NAND2_X1 U15181 ( .A1(n12013), .A2(n12012), .ZN(n12021) );
  AOI22_X1 U15182 ( .A1(n10626), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__2__SCAN_IN), .B2(n10588), .ZN(n12015) );
  AOI22_X1 U15183 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12065), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12014) );
  OAI211_X1 U15184 ( .C1(n12057), .C2(n12016), .A(n12015), .B(n12014), .ZN(
        n12020) );
  INV_X1 U15185 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12018) );
  OAI22_X1 U15186 ( .A1(n12018), .A2(n10767), .B1(n11975), .B2(n12017), .ZN(
        n12019) );
  NOR4_X1 U15187 ( .A1(n12022), .A2(n12021), .A3(n12020), .A4(n12019), .ZN(
        n14236) );
  OR2_X1 U15188 ( .A1(n12023), .A2(n14236), .ZN(n15245) );
  OR2_X1 U15189 ( .A1(n15246), .A2(n15245), .ZN(n12024) );
  AOI22_X1 U15190 ( .A1(n10577), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10654), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12026) );
  AOI22_X1 U15191 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12085), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12025) );
  OAI211_X1 U15192 ( .C1(n12048), .C2(n12027), .A(n12026), .B(n12025), .ZN(
        n12034) );
  OAI22_X1 U15193 ( .A1(n12078), .A2(n12029), .B1(n12076), .B2(n12028), .ZN(
        n12033) );
  INV_X1 U15194 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12030) );
  OAI22_X1 U15195 ( .A1(n12081), .A2(n12031), .B1(n12080), .B2(n12030), .ZN(
        n12032) );
  NOR3_X1 U15196 ( .A1(n12034), .A2(n12033), .A3(n12032), .ZN(n12044) );
  AOI22_X1 U15197 ( .A1(n12035), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11278), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12043) );
  AOI22_X1 U15198 ( .A1(n10626), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10588), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12042) );
  INV_X1 U15199 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12038) );
  OAI22_X1 U15200 ( .A1(n12039), .A2(n12038), .B1(n12037), .B2(n12036), .ZN(
        n12040) );
  AOI21_X1 U15201 ( .B1(n12064), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A(
        n12040), .ZN(n12041) );
  NAND4_X1 U15202 ( .A1(n12044), .A2(n12043), .A3(n12042), .A4(n12041), .ZN(
        n15237) );
  AOI22_X1 U15203 ( .A1(n10577), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10654), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12046) );
  AOI22_X1 U15204 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12085), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12045) );
  OAI211_X1 U15205 ( .C1(n12048), .C2(n12047), .A(n12046), .B(n12045), .ZN(
        n12063) );
  AOI22_X1 U15206 ( .A1(n12050), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12049), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12053) );
  AOI22_X1 U15207 ( .A1(n12051), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13807), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12052) );
  NAND2_X1 U15208 ( .A1(n12053), .A2(n12052), .ZN(n12062) );
  AOI22_X1 U15209 ( .A1(n10626), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10588), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12055) );
  AOI22_X1 U15210 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12065), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12054) );
  OAI211_X1 U15211 ( .C1(n12057), .C2(n12056), .A(n12055), .B(n12054), .ZN(
        n12061) );
  INV_X1 U15212 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12058) );
  OAI22_X1 U15213 ( .A1(n11975), .A2(n12059), .B1(n10767), .B2(n12058), .ZN(
        n12060) );
  NOR4_X1 U15214 ( .A1(n12063), .A2(n12062), .A3(n12061), .A4(n12060), .ZN(
        n15233) );
  NAND2_X1 U15215 ( .A1(n10626), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12070) );
  NAND2_X1 U15216 ( .A1(n12064), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12069) );
  AOI22_X1 U15217 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12065), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12068) );
  NAND2_X1 U15218 ( .A1(n10588), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n12067) );
  NAND4_X1 U15219 ( .A1(n12070), .A2(n12069), .A3(n12068), .A4(n12067), .ZN(
        n12074) );
  INV_X1 U15220 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12071) );
  OAI22_X1 U15221 ( .A1(n12072), .A2(n11975), .B1(n10767), .B2(n12071), .ZN(
        n12073) );
  NOR2_X1 U15222 ( .A1(n12074), .A2(n12073), .ZN(n12092) );
  OAI22_X1 U15223 ( .A1(n12078), .A2(n12077), .B1(n12076), .B2(n12075), .ZN(
        n12084) );
  INV_X1 U15224 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12082) );
  INV_X1 U15225 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12079) );
  OAI22_X1 U15226 ( .A1(n12082), .A2(n12081), .B1(n12080), .B2(n12079), .ZN(
        n12083) );
  NOR2_X1 U15227 ( .A1(n12084), .A2(n12083), .ZN(n12091) );
  AOI22_X1 U15228 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10574), .B1(
        n12085), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12088) );
  NAND2_X1 U15229 ( .A1(n12086), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n12087) );
  AND2_X1 U15230 ( .A1(n12088), .A2(n12087), .ZN(n12090) );
  INV_X1 U15231 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n19207) );
  AOI22_X1 U15232 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n10577), .B1(
        n10654), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12089) );
  NAND4_X1 U15233 ( .A1(n12092), .A2(n12091), .A3(n12090), .A4(n12089), .ZN(
        n12112) );
  AOI22_X1 U15234 ( .A1(n12093), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14539), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12103) );
  BUF_X1 U15235 ( .A(n12094), .Z(n14537) );
  AOI22_X1 U15236 ( .A1(n14537), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12102) );
  AND2_X1 U15237 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12096) );
  OR2_X1 U15238 ( .A1(n12096), .A2(n12095), .ZN(n14546) );
  INV_X1 U15239 ( .A(n14546), .ZN(n12204) );
  NAND2_X1 U15240 ( .A1(n14532), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12098) );
  AND3_X1 U15241 ( .A1(n12204), .A2(n12098), .A3(n12097), .ZN(n12101) );
  AOI22_X1 U15242 ( .A1(n10557), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14542), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12100) );
  NAND4_X1 U15243 ( .A1(n12103), .A2(n12102), .A3(n12101), .A4(n12100), .ZN(
        n12111) );
  AOI22_X1 U15244 ( .A1(n12093), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14539), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12109) );
  AOI22_X1 U15245 ( .A1(n14537), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12108) );
  AOI22_X1 U15246 ( .A1(n10557), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14542), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12107) );
  NAND2_X1 U15247 ( .A1(n14532), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12105) );
  AND3_X1 U15248 ( .A1(n12105), .A2(n14546), .A3(n12104), .ZN(n12106) );
  NAND4_X1 U15249 ( .A1(n12109), .A2(n12108), .A3(n12107), .A4(n12106), .ZN(
        n12110) );
  AND2_X1 U15250 ( .A1(n12111), .A2(n12110), .ZN(n12117) );
  NAND2_X1 U15251 ( .A1(n12135), .A2(n19169), .ZN(n12116) );
  INV_X1 U15252 ( .A(n12112), .ZN(n12114) );
  NAND2_X1 U15253 ( .A1(n19169), .A2(n12117), .ZN(n12113) );
  NAND2_X1 U15254 ( .A1(n12114), .A2(n12113), .ZN(n12115) );
  NAND2_X1 U15255 ( .A1(n12116), .A2(n12115), .ZN(n12138) );
  XNOR2_X1 U15256 ( .A(n15232), .B(n12138), .ZN(n15224) );
  INV_X1 U15257 ( .A(n12117), .ZN(n12118) );
  NOR2_X1 U15258 ( .A1(n19169), .A2(n12118), .ZN(n15223) );
  INV_X1 U15259 ( .A(n15232), .ZN(n12119) );
  AOI22_X1 U15260 ( .A1(n14537), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14539), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12125) );
  AOI22_X1 U15261 ( .A1(n12093), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12124) );
  NAND2_X1 U15262 ( .A1(n14543), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12121) );
  NAND2_X1 U15263 ( .A1(n14542), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12120) );
  AND3_X1 U15264 ( .A1(n12204), .A2(n12121), .A3(n12120), .ZN(n12123) );
  NAND4_X1 U15265 ( .A1(n12125), .A2(n12124), .A3(n12123), .A4(n12122), .ZN(
        n12133) );
  AOI22_X1 U15266 ( .A1(n12093), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n14539), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12131) );
  AOI22_X1 U15267 ( .A1(n14537), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12130) );
  AOI22_X1 U15268 ( .A1(n10557), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n14542), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12129) );
  NAND2_X1 U15269 ( .A1(n14543), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12127) );
  AND3_X1 U15270 ( .A1(n12127), .A2(n14546), .A3(n12126), .ZN(n12128) );
  NAND4_X1 U15271 ( .A1(n12131), .A2(n12130), .A3(n12129), .A4(n12128), .ZN(
        n12132) );
  AND2_X1 U15272 ( .A1(n12133), .A2(n12132), .ZN(n12134) );
  INV_X1 U15273 ( .A(n12134), .ZN(n15216) );
  INV_X1 U15274 ( .A(n12135), .ZN(n12136) );
  AND2_X1 U15275 ( .A1(n12135), .A2(n12134), .ZN(n12155) );
  AOI211_X1 U15276 ( .C1(n15216), .C2(n12136), .A(n12193), .B(n12155), .ZN(
        n15218) );
  INV_X1 U15277 ( .A(n15223), .ZN(n12137) );
  NOR3_X1 U15278 ( .A1(n12138), .A2(n15216), .A3(n12137), .ZN(n12139) );
  AOI22_X1 U15279 ( .A1(n12093), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14539), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12145) );
  AOI22_X1 U15280 ( .A1(n14537), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12144) );
  NAND2_X1 U15281 ( .A1(n14543), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n12141) );
  AND3_X1 U15282 ( .A1(n12204), .A2(n12141), .A3(n12140), .ZN(n12143) );
  AOI22_X1 U15283 ( .A1(n10557), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14542), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12142) );
  NAND4_X1 U15284 ( .A1(n12145), .A2(n12144), .A3(n12143), .A4(n12142), .ZN(
        n12153) );
  AOI22_X1 U15285 ( .A1(n12093), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14539), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12151) );
  AOI22_X1 U15286 ( .A1(n14537), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12150) );
  AOI22_X1 U15287 ( .A1(n10557), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n14542), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12149) );
  NAND2_X1 U15288 ( .A1(n14543), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12147) );
  AND3_X1 U15289 ( .A1(n12147), .A2(n14546), .A3(n12146), .ZN(n12148) );
  NAND4_X1 U15290 ( .A1(n12151), .A2(n12150), .A3(n12149), .A4(n12148), .ZN(
        n12152) );
  AND2_X1 U15291 ( .A1(n12153), .A2(n12152), .ZN(n12156) );
  NAND2_X1 U15292 ( .A1(n12155), .A2(n12156), .ZN(n12173) );
  OAI211_X1 U15293 ( .C1(n12155), .C2(n12156), .A(n12154), .B(n12173), .ZN(
        n12157) );
  NAND2_X1 U15294 ( .A1(n10512), .A2(n12156), .ZN(n15205) );
  AOI22_X1 U15295 ( .A1(n12093), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14537), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12164) );
  AOI22_X1 U15296 ( .A1(n14539), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12163) );
  NAND2_X1 U15297 ( .A1(n14543), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n12160) );
  NAND2_X1 U15298 ( .A1(n14542), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12159) );
  AND3_X1 U15299 ( .A1(n12204), .A2(n12160), .A3(n12159), .ZN(n12161) );
  NAND4_X1 U15300 ( .A1(n12164), .A2(n12163), .A3(n12162), .A4(n12161), .ZN(
        n12172) );
  AOI22_X1 U15301 ( .A1(n12093), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14539), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12170) );
  AOI22_X1 U15302 ( .A1(n14537), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12169) );
  NAND2_X1 U15303 ( .A1(n14543), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12166) );
  NAND2_X1 U15304 ( .A1(n14542), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n12165) );
  AND3_X1 U15305 ( .A1(n12166), .A2(n14546), .A3(n12165), .ZN(n12167) );
  NAND4_X1 U15306 ( .A1(n12170), .A2(n12169), .A3(n12168), .A4(n12167), .ZN(
        n12171) );
  NAND2_X1 U15307 ( .A1(n12172), .A2(n12171), .ZN(n12175) );
  AOI21_X1 U15308 ( .B1(n12173), .B2(n12175), .A(n12193), .ZN(n12174) );
  INV_X1 U15309 ( .A(n12175), .ZN(n12176) );
  NAND2_X1 U15310 ( .A1(n10512), .A2(n12176), .ZN(n15195) );
  NOR2_X2 U15311 ( .A1(n15194), .A2(n12178), .ZN(n12200) );
  AOI22_X1 U15312 ( .A1(n12093), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14539), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12184) );
  AOI22_X1 U15313 ( .A1(n14537), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12183) );
  NAND2_X1 U15314 ( .A1(n14543), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12180) );
  AND3_X1 U15315 ( .A1(n12204), .A2(n12180), .A3(n12179), .ZN(n12182) );
  AOI22_X1 U15316 ( .A1(n10557), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12225), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12181) );
  NAND4_X1 U15317 ( .A1(n12184), .A2(n12183), .A3(n12182), .A4(n12181), .ZN(
        n12192) );
  AOI22_X1 U15318 ( .A1(n12093), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n14539), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12190) );
  AOI22_X1 U15319 ( .A1(n14537), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12189) );
  AOI22_X1 U15320 ( .A1(n10557), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12225), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12188) );
  NAND2_X1 U15321 ( .A1(n14543), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12186) );
  AND3_X1 U15322 ( .A1(n12186), .A2(n12185), .A3(n14546), .ZN(n12187) );
  NAND4_X1 U15323 ( .A1(n12190), .A2(n12189), .A3(n12188), .A4(n12187), .ZN(
        n12191) );
  NAND2_X1 U15324 ( .A1(n12192), .A2(n12191), .ZN(n12195) );
  AOI21_X1 U15325 ( .B1(n12194), .B2(n12195), .A(n12193), .ZN(n12197) );
  INV_X1 U15326 ( .A(n12194), .ZN(n12196) );
  INV_X1 U15327 ( .A(n12195), .ZN(n12198) );
  NAND2_X1 U15328 ( .A1(n12196), .A2(n12198), .ZN(n15182) );
  NAND2_X1 U15329 ( .A1(n12197), .A2(n15182), .ZN(n12199) );
  XNOR2_X1 U15330 ( .A(n12200), .B(n12199), .ZN(n15188) );
  NAND2_X1 U15331 ( .A1(n10512), .A2(n12198), .ZN(n15189) );
  INV_X1 U15332 ( .A(n15181), .ZN(n12201) );
  AOI22_X1 U15333 ( .A1(n12093), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14537), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12208) );
  AOI22_X1 U15334 ( .A1(n14539), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10347), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12207) );
  AOI22_X1 U15335 ( .A1(n10557), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12225), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12206) );
  NAND2_X1 U15336 ( .A1(n14543), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n12203) );
  AND3_X1 U15337 ( .A1(n12204), .A2(n12203), .A3(n12202), .ZN(n12205) );
  NAND4_X1 U15338 ( .A1(n12208), .A2(n12207), .A3(n12206), .A4(n12205), .ZN(
        n12216) );
  AOI22_X1 U15339 ( .A1(n12093), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14539), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12214) );
  AOI22_X1 U15340 ( .A1(n14537), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12213) );
  AOI22_X1 U15341 ( .A1(n10557), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12225), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12212) );
  NAND2_X1 U15342 ( .A1(n14543), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12210) );
  AND3_X1 U15343 ( .A1(n12210), .A2(n14546), .A3(n12209), .ZN(n12211) );
  NAND4_X1 U15344 ( .A1(n12214), .A2(n12213), .A3(n12212), .A4(n12211), .ZN(
        n12215) );
  AND2_X1 U15345 ( .A1(n12216), .A2(n12215), .ZN(n12233) );
  NAND2_X1 U15346 ( .A1(n12217), .A2(n12233), .ZN(n14529) );
  AOI22_X1 U15347 ( .A1(n10553), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14539), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12219) );
  AOI22_X1 U15348 ( .A1(n14537), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10347), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12218) );
  NAND2_X1 U15349 ( .A1(n12219), .A2(n12218), .ZN(n12232) );
  AOI21_X1 U15350 ( .B1(n14532), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n14546), .ZN(n12221) );
  AOI22_X1 U15351 ( .A1(n10557), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12225), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12220) );
  OAI211_X1 U15352 ( .C1(n14536), .C2(n12222), .A(n12221), .B(n12220), .ZN(
        n12231) );
  AOI22_X1 U15353 ( .A1(n12093), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n14539), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12224) );
  AOI22_X1 U15354 ( .A1(n14537), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10347), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12223) );
  NAND2_X1 U15355 ( .A1(n12224), .A2(n12223), .ZN(n12230) );
  AOI22_X1 U15356 ( .A1(n10557), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12225), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12228) );
  NAND2_X1 U15357 ( .A1(n14543), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12226) );
  NAND4_X1 U15358 ( .A1(n12228), .A2(n14546), .A3(n12227), .A4(n12226), .ZN(
        n12229) );
  OAI22_X1 U15359 ( .A1(n12232), .A2(n12231), .B1(n12230), .B2(n12229), .ZN(
        n14526) );
  INV_X1 U15360 ( .A(n12233), .ZN(n15184) );
  NOR3_X1 U15361 ( .A1(n15182), .A2(n10512), .A3(n15184), .ZN(n14525) );
  XOR2_X1 U15362 ( .A(n14526), .B(n14525), .Z(n14528) );
  XNOR2_X1 U15363 ( .A(n14529), .B(n14528), .ZN(n15180) );
  AND2_X1 U15364 ( .A1(n11199), .A2(n19858), .ZN(n13354) );
  AND2_X1 U15365 ( .A1(n13354), .A2(n13353), .ZN(n12234) );
  AOI22_X1 U15366 ( .A1(n16313), .A2(n13796), .B1(n12234), .B2(n11216), .ZN(
        n13383) );
  NAND2_X1 U15367 ( .A1(n12235), .A2(n13389), .ZN(n12236) );
  XOR2_X1 U15368 ( .A(n12238), .B(n14505), .Z(n16058) );
  NAND2_X1 U15369 ( .A1(n19033), .A2(n12239), .ZN(n16134) );
  NOR4_X1 U15370 ( .A1(P2_ADDRESS_REG_16__SCAN_IN), .A2(
        P2_ADDRESS_REG_14__SCAN_IN), .A3(P2_ADDRESS_REG_13__SCAN_IN), .A4(
        P2_ADDRESS_REG_12__SCAN_IN), .ZN(n12243) );
  NOR4_X1 U15371 ( .A1(P2_ADDRESS_REG_20__SCAN_IN), .A2(
        P2_ADDRESS_REG_19__SCAN_IN), .A3(P2_ADDRESS_REG_18__SCAN_IN), .A4(
        P2_ADDRESS_REG_17__SCAN_IN), .ZN(n12242) );
  NOR4_X1 U15372 ( .A1(P2_ADDRESS_REG_7__SCAN_IN), .A2(
        P2_ADDRESS_REG_6__SCAN_IN), .A3(P2_ADDRESS_REG_5__SCAN_IN), .A4(
        P2_ADDRESS_REG_4__SCAN_IN), .ZN(n12241) );
  NOR4_X1 U15373 ( .A1(P2_ADDRESS_REG_11__SCAN_IN), .A2(
        P2_ADDRESS_REG_10__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n12240) );
  NAND4_X1 U15374 ( .A1(n12243), .A2(n12242), .A3(n12241), .A4(n12240), .ZN(
        n12248) );
  NOR4_X1 U15375 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_15__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n12246) );
  NOR4_X1 U15376 ( .A1(P2_ADDRESS_REG_24__SCAN_IN), .A2(
        P2_ADDRESS_REG_23__SCAN_IN), .A3(P2_ADDRESS_REG_22__SCAN_IN), .A4(
        P2_ADDRESS_REG_21__SCAN_IN), .ZN(n12245) );
  NOR4_X1 U15377 ( .A1(P2_ADDRESS_REG_3__SCAN_IN), .A2(
        P2_ADDRESS_REG_27__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_25__SCAN_IN), .ZN(n12244) );
  INV_X1 U15378 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19757) );
  NAND4_X1 U15379 ( .A1(n12246), .A2(n12245), .A3(n12244), .A4(n19757), .ZN(
        n12247) );
  AOI22_X1 U15380 ( .A1(n19156), .A2(BUF1_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n19158), .ZN(n13813) );
  INV_X1 U15381 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n19070) );
  OAI22_X1 U15382 ( .A1(n16134), .A2(n13813), .B1(n15340), .B2(n19070), .ZN(
        n12249) );
  AOI21_X1 U15383 ( .B1(n19051), .B2(n16058), .A(n12249), .ZN(n12250) );
  INV_X1 U15384 ( .A(n12250), .ZN(n12254) );
  AND2_X1 U15385 ( .A1(n19199), .A2(n10425), .ZN(n12251) );
  NAND2_X1 U15386 ( .A1(n19033), .A2(n12251), .ZN(n13670) );
  AOI22_X1 U15387 ( .A1(n18999), .A2(BUF2_REG_29__SCAN_IN), .B1(n18998), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n12252) );
  INV_X1 U15388 ( .A(n12252), .ZN(n12253) );
  OAI21_X1 U15389 ( .B1(n15180), .B2(n16136), .A(n12255), .ZN(P2_U2890) );
  NAND2_X1 U15390 ( .A1(n12594), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12259) );
  AND2_X2 U15391 ( .A1(n12272), .A2(n12266), .ZN(n12364) );
  NAND2_X1 U15392 ( .A1(n12364), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n12258) );
  NAND2_X1 U15393 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n12257) );
  NAND2_X1 U15394 ( .A1(n12984), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n12256) );
  AND2_X2 U15395 ( .A1(n12273), .A2(n12266), .ZN(n12438) );
  NAND2_X1 U15396 ( .A1(n12438), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n12264) );
  AND2_X4 U15397 ( .A1(n12271), .A2(n13743), .ZN(n12490) );
  NAND2_X1 U15398 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n12263) );
  AND2_X2 U15399 ( .A1(n12266), .A2(n13740), .ZN(n12425) );
  NAND2_X1 U15400 ( .A1(n12425), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12262) );
  AND2_X4 U15401 ( .A1(n13739), .A2(n13743), .ZN(n12430) );
  NAND2_X1 U15402 ( .A1(n12430), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n12261) );
  NAND2_X1 U15403 ( .A1(n12424), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n12270) );
  AND2_X2 U15404 ( .A1(n12271), .A2(n13740), .ZN(n12332) );
  NAND2_X1 U15405 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n12269) );
  NAND2_X1 U15407 ( .A1(n13045), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n12268) );
  NAND2_X1 U15408 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n12267) );
  AND2_X2 U15409 ( .A1(n12272), .A2(n12271), .ZN(n12337) );
  NAND2_X1 U15410 ( .A1(n12337), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n12279) );
  NAND2_X1 U15411 ( .A1(n12489), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12278) );
  NAND2_X1 U15412 ( .A1(n12491), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12277) );
  AND2_X2 U15413 ( .A1(n13745), .A2(n12275), .ZN(n12853) );
  NAND2_X1 U15414 ( .A1(n12853), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n12276) );
  AOI22_X1 U15415 ( .A1(n12337), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12287) );
  AOI22_X1 U15416 ( .A1(n12438), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12490), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12286) );
  AOI22_X1 U15417 ( .A1(n12491), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12853), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12285) );
  AOI22_X1 U15418 ( .A1(n12425), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12284) );
  NAND4_X1 U15419 ( .A1(n12287), .A2(n12286), .A3(n12285), .A4(n12284), .ZN(
        n12293) );
  AOI22_X1 U15420 ( .A1(n12594), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12364), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12291) );
  AOI22_X1 U15421 ( .A1(n12424), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13045), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12290) );
  AOI22_X1 U15422 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12595), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12289) );
  AOI22_X1 U15423 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12984), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12288) );
  NAND4_X1 U15424 ( .A1(n12291), .A2(n12290), .A3(n12289), .A4(n12288), .ZN(
        n12292) );
  NAND2_X1 U15425 ( .A1(n12594), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12297) );
  NAND2_X1 U15426 ( .A1(n12364), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12296) );
  NAND2_X1 U15427 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n12295) );
  NAND2_X1 U15428 ( .A1(n12984), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n12294) );
  NAND2_X1 U15429 ( .A1(n12337), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n12301) );
  NAND2_X1 U15430 ( .A1(n12489), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12300) );
  NAND2_X1 U15431 ( .A1(n12491), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12299) );
  NAND2_X1 U15432 ( .A1(n12853), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n12298) );
  NAND2_X1 U15433 ( .A1(n12424), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n12305) );
  NAND2_X1 U15434 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12304) );
  NAND2_X1 U15435 ( .A1(n13045), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12303) );
  NAND2_X1 U15436 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n12302) );
  NAND2_X1 U15437 ( .A1(n12438), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n12309) );
  NAND2_X1 U15438 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n12308) );
  NAND2_X1 U15439 ( .A1(n12425), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12307) );
  NAND2_X1 U15440 ( .A1(n12430), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12306) );
  AOI22_X1 U15441 ( .A1(n12594), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12364), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12317) );
  AOI22_X1 U15442 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12425), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12316) );
  AOI22_X1 U15443 ( .A1(n12424), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12595), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12315) );
  AOI22_X1 U15444 ( .A1(n12337), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12314) );
  AOI22_X1 U15445 ( .A1(n12489), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12490), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12321) );
  AOI22_X1 U15446 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13045), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12320) );
  AOI22_X1 U15447 ( .A1(n12438), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12984), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12319) );
  AOI22_X1 U15448 ( .A1(n12491), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12853), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12318) );
  AOI22_X1 U15449 ( .A1(n12594), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12364), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12326) );
  AOI22_X1 U15450 ( .A1(n12337), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12325) );
  AOI22_X1 U15451 ( .A1(n12424), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12425), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12324) );
  AOI22_X1 U15452 ( .A1(n12438), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12332), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12323) );
  AOI22_X1 U15453 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12984), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12330) );
  AOI22_X1 U15454 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13045), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12329) );
  AOI22_X1 U15455 ( .A1(n12491), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12853), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12328) );
  AOI22_X1 U15456 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12327) );
  NAND2_X2 U15457 ( .A1(n12331), .A2(n9884), .ZN(n20146) );
  AOI22_X1 U15458 ( .A1(n12424), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13045), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12335) );
  AOI22_X1 U15459 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12595), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12334) );
  AOI22_X1 U15460 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12984), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12333) );
  NAND4_X1 U15461 ( .A1(n12336), .A2(n12335), .A3(n12334), .A4(n12333), .ZN(
        n12343) );
  AOI22_X1 U15462 ( .A1(n12337), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12341) );
  AOI22_X1 U15463 ( .A1(n12438), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12490), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12340) );
  AOI22_X1 U15464 ( .A1(n12491), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12853), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12339) );
  AOI22_X1 U15465 ( .A1(n12425), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12338) );
  NAND4_X1 U15466 ( .A1(n12341), .A2(n12340), .A3(n12339), .A4(n12338), .ZN(
        n12342) );
  AND2_X1 U15467 ( .A1(n13125), .A2(n12396), .ZN(n12387) );
  NAND2_X1 U15468 ( .A1(n12594), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12347) );
  NAND2_X1 U15469 ( .A1(n12364), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12346) );
  NAND2_X1 U15470 ( .A1(n13045), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12345) );
  NAND2_X1 U15471 ( .A1(n12984), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12344) );
  NAND2_X1 U15472 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12351) );
  NAND2_X1 U15473 ( .A1(n12337), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12350) );
  NAND2_X1 U15474 ( .A1(n12489), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12349) );
  NAND2_X1 U15475 ( .A1(n12438), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12348) );
  NAND2_X1 U15476 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12355) );
  NAND2_X1 U15477 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12354) );
  NAND2_X1 U15478 ( .A1(n12425), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12353) );
  NAND2_X1 U15479 ( .A1(n12430), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12352) );
  NAND2_X1 U15480 ( .A1(n12424), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12359) );
  NAND2_X1 U15481 ( .A1(n12853), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12358) );
  NAND2_X1 U15482 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12357) );
  NAND2_X1 U15483 ( .A1(n12491), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12356) );
  NAND2_X1 U15484 ( .A1(n12364), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12366) );
  NAND2_X1 U15485 ( .A1(n12594), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12365) );
  NAND2_X1 U15486 ( .A1(n12366), .A2(n12365), .ZN(n12370) );
  NAND2_X1 U15487 ( .A1(n12984), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12368) );
  NAND2_X1 U15488 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12367) );
  NAND2_X1 U15489 ( .A1(n12368), .A2(n12367), .ZN(n12369) );
  NOR2_X1 U15490 ( .A1(n12370), .A2(n12369), .ZN(n12386) );
  NAND2_X1 U15491 ( .A1(n12337), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12374) );
  NAND2_X1 U15492 ( .A1(n12489), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12373) );
  NAND2_X1 U15493 ( .A1(n12491), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12372) );
  NAND2_X1 U15494 ( .A1(n12853), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12371) );
  NAND2_X1 U15495 ( .A1(n12424), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12378) );
  NAND2_X1 U15496 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12377) );
  NAND2_X1 U15497 ( .A1(n12595), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12375) );
  NAND2_X1 U15498 ( .A1(n12438), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12382) );
  NAND2_X1 U15499 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12381) );
  NAND2_X1 U15500 ( .A1(n12425), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12380) );
  NAND2_X1 U15501 ( .A1(n12430), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12379) );
  NAND2_X2 U15502 ( .A1(n20139), .A2(n20124), .ZN(n14609) );
  NAND2_X1 U15503 ( .A1(n13538), .A2(n20124), .ZN(n13928) );
  NAND2_X1 U15504 ( .A1(n13541), .A2(n13928), .ZN(n12390) );
  INV_X1 U15505 ( .A(n20146), .ZN(n12388) );
  NAND2_X1 U15506 ( .A1(n14615), .A2(n13509), .ZN(n13622) );
  NAND2_X1 U15507 ( .A1(n13620), .A2(n12396), .ZN(n12389) );
  NAND2_X1 U15508 ( .A1(n13622), .A2(n12389), .ZN(n13546) );
  NOR2_X2 U15509 ( .A1(n12390), .A2(n13546), .ZN(n12421) );
  NAND2_X1 U15510 ( .A1(n13165), .A2(n13141), .ZN(n12391) );
  NAND2_X1 U15511 ( .A1(n12391), .A2(n12509), .ZN(n13124) );
  NOR2_X1 U15512 ( .A1(n13124), .A2(n12392), .ZN(n12397) );
  NOR2_X2 U15513 ( .A1(n12396), .A2(n20146), .ZN(n12404) );
  INV_X1 U15514 ( .A(n12404), .ZN(n13753) );
  INV_X1 U15515 ( .A(n12397), .ZN(n12415) );
  INV_X1 U15516 ( .A(n12393), .ZN(n12398) );
  NAND2_X1 U15517 ( .A1(n12415), .A2(n15156), .ZN(n12418) );
  NAND4_X1 U15518 ( .A1(n12421), .A2(n13544), .A3(n13753), .A4(n12418), .ZN(
        n12406) );
  NAND2_X1 U15519 ( .A1(n13509), .A2(n20124), .ZN(n12400) );
  NAND4_X1 U15520 ( .A1(n12402), .A2(n13165), .A3(n20150), .A4(n12509), .ZN(
        n12403) );
  AND2_X2 U15521 ( .A1(n13501), .A2(n13620), .ZN(n13518) );
  INV_X1 U15522 ( .A(n13518), .ZN(n13374) );
  XNOR2_X1 U15523 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n13497) );
  OAI21_X1 U15524 ( .B1(n13374), .B2(n13497), .A(n13614), .ZN(n12405) );
  NAND2_X1 U15525 ( .A1(n13553), .A2(n20706), .ZN(n13258) );
  NAND2_X1 U15526 ( .A1(n20638), .A2(n20563), .ZN(n20529) );
  NAND2_X1 U15527 ( .A1(n20529), .A2(n12534), .ZN(n20454) );
  OR2_X1 U15528 ( .A1(n15736), .A2(n20638), .ZN(n12478) );
  OAI21_X1 U15529 ( .B1(n13258), .B2(n20454), .A(n12478), .ZN(n12407) );
  INV_X1 U15530 ( .A(n12407), .ZN(n12408) );
  MUX2_X1 U15531 ( .A(n13258), .B(n15736), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n12411) );
  OAI21_X2 U15532 ( .B1(n12484), .B2(n13554), .A(n12411), .ZN(n12454) );
  NAND2_X1 U15533 ( .A1(n14404), .A2(n14609), .ZN(n13458) );
  INV_X1 U15534 ( .A(n13553), .ZN(n20790) );
  NOR2_X1 U15535 ( .A1(n20790), .A2(n20706), .ZN(n12413) );
  NAND2_X1 U15536 ( .A1(n12404), .A2(n12402), .ZN(n13623) );
  OAI211_X1 U15537 ( .C1(n9840), .C2(n13458), .A(n12413), .B(n13623), .ZN(
        n12414) );
  INV_X1 U15538 ( .A(n12414), .ZN(n12417) );
  AND2_X1 U15539 ( .A1(n13620), .A2(n20139), .ZN(n20009) );
  NAND2_X1 U15540 ( .A1(n12415), .A2(n20009), .ZN(n12416) );
  OAI211_X1 U15541 ( .C1(n20139), .C2(n12418), .A(n12417), .B(n12416), .ZN(
        n12419) );
  INV_X1 U15542 ( .A(n12419), .ZN(n12420) );
  NAND2_X1 U15543 ( .A1(n12421), .A2(n12420), .ZN(n12455) );
  INV_X1 U15544 ( .A(n20238), .ZN(n12423) );
  AOI22_X1 U15545 ( .A1(n12982), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13039), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12429) );
  AOI22_X1 U15546 ( .A1(n13040), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12490), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12428) );
  AOI22_X1 U15547 ( .A1(n12443), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13049), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12427) );
  AOI22_X1 U15548 ( .A1(n13046), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12871), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12426) );
  NAND4_X1 U15549 ( .A1(n12429), .A2(n12428), .A3(n12427), .A4(n12426), .ZN(
        n12436) );
  AOI22_X1 U15550 ( .A1(n13047), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13022), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12434) );
  AOI22_X1 U15551 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13050), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12433) );
  INV_X1 U15552 ( .A(n12430), .ZN(n12543) );
  AOI22_X1 U15553 ( .A1(n13038), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12432) );
  AOI22_X1 U15554 ( .A1(n13045), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13048), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12431) );
  NAND4_X1 U15555 ( .A1(n12434), .A2(n12433), .A3(n12432), .A4(n12431), .ZN(
        n12435) );
  OR2_X1 U15556 ( .A1(n12450), .A2(n12542), .ZN(n12437) );
  AOI22_X1 U15557 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13047), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12442) );
  AOI22_X1 U15558 ( .A1(n13022), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13038), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12441) );
  AOI22_X1 U15559 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12440) );
  AOI22_X1 U15560 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13046), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12439) );
  NAND4_X1 U15561 ( .A1(n12442), .A2(n12441), .A3(n12440), .A4(n12439), .ZN(
        n12449) );
  AOI22_X1 U15562 ( .A1(n12337), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13039), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12447) );
  AOI22_X1 U15563 ( .A1(n13040), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12871), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12446) );
  AOI22_X1 U15564 ( .A1(n13045), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13048), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12445) );
  BUF_X1 U15565 ( .A(n12491), .Z(n12443) );
  AOI22_X1 U15566 ( .A1(n12443), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13049), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12444) );
  NAND4_X1 U15567 ( .A1(n12447), .A2(n12446), .A3(n12445), .A4(n12444), .ZN(
        n12448) );
  OR2_X1 U15568 ( .A1(n12542), .A2(n13226), .ZN(n12453) );
  NAND2_X1 U15569 ( .A1(n20124), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12541) );
  OR2_X1 U15570 ( .A1(n12450), .A2(n12541), .ZN(n12452) );
  NAND2_X1 U15571 ( .A1(n13108), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12451) );
  INV_X1 U15572 ( .A(n12455), .ZN(n12456) );
  XNOR2_X2 U15573 ( .A(n12454), .B(n12456), .ZN(n12524) );
  AOI22_X1 U15574 ( .A1(n13047), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13022), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12460) );
  AOI22_X1 U15575 ( .A1(n12982), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13050), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12459) );
  AOI22_X1 U15576 ( .A1(n13040), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12490), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12458) );
  AOI22_X1 U15577 ( .A1(n13046), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13048), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12457) );
  NAND4_X1 U15578 ( .A1(n12460), .A2(n12459), .A3(n12458), .A4(n12457), .ZN(
        n12466) );
  AOI22_X1 U15579 ( .A1(n13039), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13038), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12464) );
  AOI22_X1 U15580 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12983), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12463) );
  AOI22_X1 U15581 ( .A1(n12443), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13049), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12462) );
  AOI22_X1 U15582 ( .A1(n12871), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12461) );
  NAND4_X1 U15583 ( .A1(n12464), .A2(n12463), .A3(n12462), .A4(n12461), .ZN(
        n12465) );
  XNOR2_X1 U15584 ( .A(n12474), .B(n13166), .ZN(n12468) );
  INV_X1 U15585 ( .A(n12542), .ZN(n12467) );
  NAND2_X1 U15586 ( .A1(n12468), .A2(n12467), .ZN(n12469) );
  INV_X1 U15587 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12473) );
  AOI21_X1 U15588 ( .B1(n20124), .B2(n13166), .A(n20706), .ZN(n12472) );
  NAND2_X1 U15589 ( .A1(n20150), .A2(n13226), .ZN(n12471) );
  OAI211_X1 U15590 ( .C1(n13116), .C2(n12473), .A(n12472), .B(n12471), .ZN(
        n12521) );
  NOR2_X1 U15591 ( .A1(n12542), .A2(n12474), .ZN(n13222) );
  INV_X1 U15592 ( .A(n13170), .ZN(n12476) );
  NAND2_X1 U15593 ( .A1(n12476), .A2(n12475), .ZN(n12477) );
  INV_X1 U15594 ( .A(n12478), .ZN(n12481) );
  INV_X1 U15595 ( .A(n12479), .ZN(n12480) );
  OAI21_X1 U15596 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n12481), .A(
        n12480), .ZN(n12482) );
  OR2_X1 U15597 ( .A1(n12484), .A2(n10190), .ZN(n12486) );
  INV_X1 U15598 ( .A(n13258), .ZN(n12538) );
  XNOR2_X1 U15599 ( .A(n12534), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20133) );
  NAND2_X1 U15600 ( .A1(n12538), .A2(n20133), .ZN(n12485) );
  AOI22_X1 U15601 ( .A1(n12982), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13039), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12495) );
  AOI22_X1 U15602 ( .A1(n13038), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12490), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12494) );
  AOI22_X1 U15603 ( .A1(n12443), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13049), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12493) );
  AOI22_X1 U15604 ( .A1(n13046), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12492) );
  NAND4_X1 U15605 ( .A1(n12495), .A2(n12494), .A3(n12493), .A4(n12492), .ZN(
        n12502) );
  AOI22_X1 U15606 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13047), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12500) );
  AOI22_X1 U15607 ( .A1(n13040), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12983), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12499) );
  AOI22_X1 U15608 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12871), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12498) );
  AOI22_X1 U15609 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13048), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12497) );
  NAND4_X1 U15610 ( .A1(n12500), .A2(n12499), .A3(n12498), .A4(n12497), .ZN(
        n12501) );
  INV_X1 U15611 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12503) );
  OAI22_X1 U15612 ( .A1(n12541), .A2(n13179), .B1(n13116), .B2(n12503), .ZN(
        n12504) );
  NAND2_X1 U15613 ( .A1(n12506), .A2(n12505), .ZN(n13774) );
  NAND2_X1 U15614 ( .A1(n12507), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12585) );
  NOR2_X1 U15615 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12508) );
  INV_X1 U15616 ( .A(n13063), .ZN(n13920) );
  XNOR2_X1 U15617 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13936) );
  AOI21_X1 U15618 ( .B1(n13920), .B2(n13936), .A(n13067), .ZN(n12511) );
  NAND2_X1 U15619 ( .A1(n13068), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n12510) );
  OAI211_X1 U15620 ( .C1(n12585), .C2(n10190), .A(n12511), .B(n12510), .ZN(
        n12512) );
  INV_X1 U15621 ( .A(n12512), .ZN(n12513) );
  NAND2_X1 U15622 ( .A1(n13067), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12531) );
  NAND2_X1 U15623 ( .A1(n13764), .A2(n12760), .ZN(n12520) );
  AOI22_X1 U15624 ( .A1(n13068), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20708), .ZN(n12518) );
  INV_X1 U15625 ( .A(n12585), .ZN(n12559) );
  NAND2_X1 U15626 ( .A1(n12559), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12517) );
  AND2_X1 U15627 ( .A1(n12518), .A2(n12517), .ZN(n12519) );
  NAND2_X1 U15628 ( .A1(n12520), .A2(n12519), .ZN(n13558) );
  NAND2_X1 U15629 ( .A1(n13164), .A2(n12402), .ZN(n12523) );
  NAND2_X1 U15630 ( .A1(n12523), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13490) );
  NAND2_X1 U15631 ( .A1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20708), .ZN(
        n12527) );
  NAND2_X1 U15632 ( .A1(n12525), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n12526) );
  OAI211_X1 U15633 ( .C1(n12585), .C2(n13554), .A(n12527), .B(n12526), .ZN(
        n12528) );
  AOI21_X1 U15634 ( .B1(n12524), .B2(n12760), .A(n12528), .ZN(n13491) );
  OR2_X1 U15635 ( .A1(n13490), .A2(n13491), .ZN(n13488) );
  NAND2_X1 U15636 ( .A1(n13491), .A2(n12508), .ZN(n12529) );
  NAND2_X1 U15637 ( .A1(n13488), .A2(n12529), .ZN(n13557) );
  NAND2_X1 U15638 ( .A1(n9932), .A2(n12530), .ZN(n13650) );
  OR2_X1 U15639 ( .A1(n12484), .A2(n12532), .ZN(n12540) );
  NAND2_X1 U15640 ( .A1(n20453), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20331) );
  INV_X1 U15641 ( .A(n20331), .ZN(n12533) );
  INV_X1 U15642 ( .A(n20391), .ZN(n12536) );
  OAI21_X1 U15643 ( .B1(n12534), .B2(n20398), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12535) );
  NAND2_X1 U15644 ( .A1(n12536), .A2(n12535), .ZN(n20399) );
  NOR2_X1 U15645 ( .A1(n15736), .A2(n20453), .ZN(n12537) );
  AOI21_X1 U15646 ( .B1(n20399), .B2(n12538), .A(n12537), .ZN(n12539) );
  AOI22_X1 U15647 ( .A1(n12982), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13039), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12547) );
  AOI22_X1 U15648 ( .A1(n13038), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12490), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12546) );
  AOI22_X1 U15649 ( .A1(n12443), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13049), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12545) );
  AOI22_X1 U15650 ( .A1(n13046), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12544) );
  NAND4_X1 U15651 ( .A1(n12547), .A2(n12546), .A3(n12545), .A4(n12544), .ZN(
        n12553) );
  AOI22_X1 U15652 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13047), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12551) );
  AOI22_X1 U15653 ( .A1(n13040), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12983), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12550) );
  AOI22_X1 U15654 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12871), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12549) );
  AOI22_X1 U15655 ( .A1(n13022), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13048), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12548) );
  NAND4_X1 U15656 ( .A1(n12551), .A2(n12550), .A3(n12549), .A4(n12548), .ZN(
        n12552) );
  AOI22_X1 U15657 ( .A1(n13079), .A2(n13194), .B1(n13108), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12554) );
  INV_X1 U15658 ( .A(n12557), .ZN(n13772) );
  NAND2_X1 U15659 ( .A1(n12559), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12564) );
  NAND2_X1 U15660 ( .A1(n13792), .A2(n12560), .ZN(n12561) );
  INV_X1 U15661 ( .A(n12579), .ZN(n12580) );
  AND2_X1 U15662 ( .A1(n12561), .A2(n12580), .ZN(n19972) );
  INV_X1 U15663 ( .A(n13067), .ZN(n12690) );
  OAI22_X1 U15664 ( .A1(n19972), .A2(n13063), .B1(n12690), .B2(n13792), .ZN(
        n12562) );
  AOI21_X1 U15665 ( .B1(n13068), .B2(P1_EAX_REG_3__SCAN_IN), .A(n12562), .ZN(
        n12563) );
  AND2_X1 U15666 ( .A1(n12564), .A2(n12563), .ZN(n12565) );
  AOI22_X1 U15667 ( .A1(n12982), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12490), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12569) );
  AOI22_X1 U15668 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n13040), .B1(
        n13038), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12568) );
  AOI22_X1 U15669 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12496), .B1(
        n13050), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12567) );
  AOI22_X1 U15670 ( .A1(n12443), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13049), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12566) );
  NAND4_X1 U15671 ( .A1(n12569), .A2(n12568), .A3(n12567), .A4(n12566), .ZN(
        n12575) );
  AOI22_X1 U15672 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n13047), .B1(
        n9829), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12573) );
  AOI22_X1 U15673 ( .A1(n13039), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12871), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12572) );
  AOI22_X1 U15674 ( .A1(n13046), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13048), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12571) );
  AOI22_X1 U15675 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12570) );
  NAND4_X1 U15676 ( .A1(n12573), .A2(n12572), .A3(n12571), .A4(n12570), .ZN(
        n12574) );
  AOI22_X1 U15677 ( .A1(n13079), .A2(n13195), .B1(
        P1_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n13108), .ZN(n12576) );
  NAND2_X1 U15678 ( .A1(n12577), .A2(n12576), .ZN(n12578) );
  NAND2_X1 U15679 ( .A1(n12605), .A2(n12578), .ZN(n13187) );
  INV_X1 U15680 ( .A(n13187), .ZN(n12589) );
  INV_X1 U15681 ( .A(n12607), .ZN(n12609) );
  INV_X1 U15682 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n12581) );
  NAND2_X1 U15683 ( .A1(n12581), .A2(n12580), .ZN(n12582) );
  NAND2_X1 U15684 ( .A1(n12609), .A2(n12582), .ZN(n20075) );
  INV_X1 U15685 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20200) );
  OAI21_X1 U15686 ( .B1(n20200), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20708), .ZN(n12584) );
  NAND2_X1 U15687 ( .A1(n13068), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n12583) );
  OAI211_X1 U15688 ( .C1(n12585), .C2(n13738), .A(n12584), .B(n12583), .ZN(
        n12586) );
  OAI21_X1 U15689 ( .B1(n13063), .B2(n20075), .A(n12586), .ZN(n12587) );
  AOI21_X1 U15690 ( .B1(n12589), .B2(n12760), .A(n12588), .ZN(n13843) );
  NOR2_X2 U15691 ( .A1(n13720), .A2(n13843), .ZN(n13826) );
  INV_X1 U15692 ( .A(n12605), .ZN(n12603) );
  INV_X1 U15693 ( .A(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n21081) );
  AOI22_X1 U15694 ( .A1(n12982), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13039), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12593) );
  AOI22_X1 U15695 ( .A1(n13038), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12490), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12592) );
  AOI22_X1 U15696 ( .A1(n12443), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13049), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12591) );
  AOI22_X1 U15697 ( .A1(n13046), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12590) );
  NAND4_X1 U15698 ( .A1(n12593), .A2(n12592), .A3(n12591), .A4(n12590), .ZN(
        n12601) );
  AOI22_X1 U15699 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13047), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12599) );
  AOI22_X1 U15700 ( .A1(n13040), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12983), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12598) );
  AOI22_X1 U15701 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12871), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12597) );
  AOI22_X1 U15702 ( .A1(n13022), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13048), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12596) );
  NAND4_X1 U15703 ( .A1(n12599), .A2(n12598), .A3(n12597), .A4(n12596), .ZN(
        n12600) );
  AOI22_X1 U15704 ( .A1(n13079), .A2(n13204), .B1(n13108), .B2(
        P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12604) );
  NAND2_X1 U15705 ( .A1(n12605), .A2(n12604), .ZN(n12606) );
  NAND2_X1 U15706 ( .A1(n12632), .A2(n12606), .ZN(n13200) );
  INV_X1 U15707 ( .A(n12623), .ZN(n12625) );
  INV_X1 U15708 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12608) );
  NAND2_X1 U15709 ( .A1(n12609), .A2(n12608), .ZN(n12610) );
  NAND2_X1 U15710 ( .A1(n12625), .A2(n12610), .ZN(n19937) );
  AOI22_X1 U15711 ( .A1(n19937), .A2(n12508), .B1(n13067), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12612) );
  NAND2_X1 U15712 ( .A1(n13068), .A2(P1_EAX_REG_5__SCAN_IN), .ZN(n12611) );
  OAI211_X1 U15713 ( .C1(n13200), .C2(n12748), .A(n12612), .B(n12611), .ZN(
        n13825) );
  NAND2_X1 U15714 ( .A1(n13826), .A2(n13825), .ZN(n13824) );
  AOI22_X1 U15715 ( .A1(n12982), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13047), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12616) );
  AOI22_X1 U15716 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13038), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12615) );
  AOI22_X1 U15717 ( .A1(n13039), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12490), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12614) );
  AOI22_X1 U15718 ( .A1(n13040), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12983), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12613) );
  NAND4_X1 U15719 ( .A1(n12616), .A2(n12615), .A3(n12614), .A4(n12613), .ZN(
        n12622) );
  AOI22_X1 U15720 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13048), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12620) );
  AOI22_X1 U15721 ( .A1(n13022), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12871), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12619) );
  AOI22_X1 U15722 ( .A1(n12443), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13049), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12618) );
  AOI22_X1 U15723 ( .A1(n13046), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12617) );
  NAND4_X1 U15724 ( .A1(n12620), .A2(n12619), .A3(n12618), .A4(n12617), .ZN(
        n12621) );
  AOI22_X1 U15725 ( .A1(n13079), .A2(n13213), .B1(n13108), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12633) );
  NAND2_X1 U15726 ( .A1(n12632), .A2(n12633), .ZN(n13203) );
  INV_X1 U15727 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n12629) );
  INV_X1 U15728 ( .A(n12637), .ZN(n12627) );
  INV_X1 U15729 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12624) );
  NAND2_X1 U15730 ( .A1(n12625), .A2(n12624), .ZN(n12626) );
  NAND2_X1 U15731 ( .A1(n12627), .A2(n12626), .ZN(n19931) );
  AOI22_X1 U15732 ( .A1(n19931), .A2(n12508), .B1(n13067), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12628) );
  OAI21_X1 U15733 ( .B1(n12909), .B2(n12629), .A(n12628), .ZN(n12630) );
  INV_X1 U15734 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12635) );
  NAND2_X1 U15735 ( .A1(n13079), .A2(n13226), .ZN(n12634) );
  OAI21_X1 U15736 ( .B1(n12635), .B2(n13116), .A(n12634), .ZN(n12636) );
  INV_X1 U15737 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n12639) );
  OAI21_X1 U15738 ( .B1(n12637), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n12656), .ZN(n19912) );
  AOI22_X1 U15739 ( .A1(n19912), .A2(n12508), .B1(n13067), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12638) );
  OAI21_X1 U15740 ( .B1(n12909), .B2(n12639), .A(n12638), .ZN(n12640) );
  AOI21_X1 U15741 ( .B1(n13212), .B2(n12760), .A(n12640), .ZN(n14011) );
  AOI22_X1 U15742 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13040), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12644) );
  AOI22_X1 U15743 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13046), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12643) );
  AOI22_X1 U15744 ( .A1(n12443), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13049), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12642) );
  AOI22_X1 U15745 ( .A1(n12337), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12641) );
  NAND4_X1 U15746 ( .A1(n12644), .A2(n12643), .A3(n12642), .A4(n12641), .ZN(
        n12650) );
  AOI22_X1 U15747 ( .A1(n13022), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13039), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12648) );
  AOI22_X1 U15748 ( .A1(n13038), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12490), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12647) );
  AOI22_X1 U15749 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12871), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12646) );
  AOI22_X1 U15750 ( .A1(n13047), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13048), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12645) );
  NAND4_X1 U15751 ( .A1(n12648), .A2(n12647), .A3(n12646), .A4(n12645), .ZN(
        n12649) );
  OAI21_X1 U15752 ( .B1(n12650), .B2(n12649), .A(n12760), .ZN(n12655) );
  NAND2_X1 U15753 ( .A1(n13068), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n12654) );
  INV_X1 U15754 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12651) );
  XNOR2_X1 U15755 ( .A(n12656), .B(n12651), .ZN(n14103) );
  NAND2_X1 U15756 ( .A1(n14103), .A2(n12508), .ZN(n12653) );
  NAND2_X1 U15757 ( .A1(n13067), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12652) );
  NAND4_X1 U15758 ( .A1(n12655), .A2(n12654), .A3(n12653), .A4(n12652), .ZN(
        n13984) );
  XNOR2_X1 U15759 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n12670), .ZN(
        n19905) );
  AOI22_X1 U15760 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13022), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12660) );
  AOI22_X1 U15761 ( .A1(n13047), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13038), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12659) );
  AOI22_X1 U15762 ( .A1(n13045), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13048), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12658) );
  AOI22_X1 U15763 ( .A1(n13039), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12657) );
  NAND4_X1 U15764 ( .A1(n12660), .A2(n12659), .A3(n12658), .A4(n12657), .ZN(
        n12666) );
  AOI22_X1 U15765 ( .A1(n12337), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12490), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12664) );
  AOI22_X1 U15766 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13046), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12663) );
  AOI22_X1 U15767 ( .A1(n13040), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12871), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12662) );
  AOI22_X1 U15768 ( .A1(n12443), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13049), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12661) );
  NAND4_X1 U15769 ( .A1(n12664), .A2(n12663), .A3(n12662), .A4(n12661), .ZN(
        n12665) );
  OR2_X1 U15770 ( .A1(n12666), .A2(n12665), .ZN(n12667) );
  AOI22_X1 U15771 ( .A1(n12760), .A2(n12667), .B1(n13067), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12669) );
  NAND2_X1 U15772 ( .A1(n12525), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12668) );
  OAI211_X1 U15773 ( .C1(n19905), .C2(n13063), .A(n12669), .B(n12668), .ZN(
        n14057) );
  NAND2_X1 U15774 ( .A1(n13986), .A2(n14057), .ZN(n14056) );
  INV_X2 U15775 ( .A(n14056), .ZN(n12686) );
  XNOR2_X1 U15776 ( .A(n12687), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14951) );
  AOI22_X1 U15777 ( .A1(n13040), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12983), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12674) );
  AOI22_X1 U15778 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13046), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12673) );
  AOI22_X1 U15779 ( .A1(n12443), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13049), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12672) );
  AOI22_X1 U15780 ( .A1(n13038), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12671) );
  NAND4_X1 U15781 ( .A1(n12674), .A2(n12673), .A3(n12672), .A4(n12671), .ZN(
        n12680) );
  AOI22_X1 U15782 ( .A1(n13047), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13022), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12678) );
  AOI22_X1 U15783 ( .A1(n13039), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13050), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12677) );
  BUF_X1 U15784 ( .A(n12337), .Z(n12982) );
  AOI22_X1 U15785 ( .A1(n12982), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13048), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12676) );
  AOI22_X1 U15786 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12871), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12675) );
  NAND4_X1 U15787 ( .A1(n12678), .A2(n12677), .A3(n12676), .A4(n12675), .ZN(
        n12679) );
  OAI21_X1 U15788 ( .B1(n12680), .B2(n12679), .A(n12760), .ZN(n12683) );
  NAND2_X1 U15789 ( .A1(n12525), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n12682) );
  NAND2_X1 U15790 ( .A1(n13067), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12681) );
  NAND3_X1 U15791 ( .A1(n12683), .A2(n12682), .A3(n12681), .ZN(n12684) );
  AOI21_X1 U15792 ( .B1(n14951), .B2(n12508), .A(n12684), .ZN(n14141) );
  INV_X1 U15793 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12691) );
  OAI21_X1 U15794 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n12688), .A(
        n12729), .ZN(n15928) );
  NAND2_X1 U15795 ( .A1(n15928), .A2(n12508), .ZN(n12689) );
  OAI21_X1 U15796 ( .B1(n12691), .B2(n12690), .A(n12689), .ZN(n12692) );
  AOI21_X1 U15797 ( .B1(n12525), .B2(P1_EAX_REG_11__SCAN_IN), .A(n12692), .ZN(
        n14266) );
  AOI22_X1 U15798 ( .A1(n12982), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13039), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12697) );
  AOI22_X1 U15799 ( .A1(n13038), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12490), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12696) );
  AOI22_X1 U15800 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13050), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12695) );
  AOI22_X1 U15801 ( .A1(n12443), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13049), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12694) );
  NAND4_X1 U15802 ( .A1(n12697), .A2(n12696), .A3(n12695), .A4(n12694), .ZN(
        n12703) );
  AOI22_X1 U15803 ( .A1(n13022), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12983), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12701) );
  AOI22_X1 U15804 ( .A1(n13046), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13048), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12700) );
  AOI22_X1 U15805 ( .A1(n13047), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12871), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12699) );
  AOI22_X1 U15806 ( .A1(n13040), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12698) );
  NAND4_X1 U15807 ( .A1(n12701), .A2(n12700), .A3(n12699), .A4(n12698), .ZN(
        n12702) );
  NOR2_X1 U15808 ( .A1(n12703), .A2(n12702), .ZN(n12704) );
  OR2_X1 U15809 ( .A1(n12748), .A2(n12704), .ZN(n14274) );
  XNOR2_X1 U15810 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n12745), .ZN(
        n14942) );
  AOI22_X1 U15811 ( .A1(n12982), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13039), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12709) );
  AOI22_X1 U15812 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13040), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12708) );
  AOI22_X1 U15813 ( .A1(n13038), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13046), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12707) );
  AOI22_X1 U15814 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13048), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12706) );
  NAND4_X1 U15815 ( .A1(n12709), .A2(n12708), .A3(n12707), .A4(n12706), .ZN(
        n12715) );
  AOI22_X1 U15816 ( .A1(n13047), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12490), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12713) );
  AOI22_X1 U15817 ( .A1(n13022), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12871), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12712) );
  AOI22_X1 U15818 ( .A1(n12443), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13049), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12711) );
  AOI22_X1 U15819 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12710) );
  NAND4_X1 U15820 ( .A1(n12713), .A2(n12712), .A3(n12711), .A4(n12710), .ZN(
        n12714) );
  OR2_X1 U15821 ( .A1(n12715), .A2(n12714), .ZN(n12716) );
  AOI22_X1 U15822 ( .A1(n12760), .A2(n12716), .B1(n13067), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12718) );
  NAND2_X1 U15823 ( .A1(n12525), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n12717) );
  OAI211_X1 U15824 ( .C1(n14942), .C2(n13063), .A(n12718), .B(n12717), .ZN(
        n14269) );
  AOI22_X1 U15825 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12496), .B1(
        n13047), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12722) );
  AOI22_X1 U15826 ( .A1(n12982), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13039), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12721) );
  AOI22_X1 U15827 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n13038), .B1(
        n13050), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12720) );
  AOI22_X1 U15828 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12983), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12719) );
  NAND4_X1 U15829 ( .A1(n12722), .A2(n12721), .A3(n12720), .A4(n12719), .ZN(
        n12728) );
  AOI22_X1 U15830 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n13040), .B1(
        n12871), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12726) );
  AOI22_X1 U15831 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n9829), .B1(
        n13048), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12725) );
  AOI22_X1 U15832 ( .A1(n12443), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13049), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12724) );
  AOI22_X1 U15833 ( .A1(n13046), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12723) );
  NAND4_X1 U15834 ( .A1(n12726), .A2(n12725), .A3(n12724), .A4(n12723), .ZN(
        n12727) );
  NOR2_X1 U15835 ( .A1(n12728), .A2(n12727), .ZN(n12733) );
  XNOR2_X1 U15836 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n12729), .ZN(
        n15916) );
  INV_X1 U15837 ( .A(n15916), .ZN(n12730) );
  AOI22_X1 U15838 ( .A1(n13067), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n13920), .B2(n12730), .ZN(n12732) );
  NAND2_X1 U15839 ( .A1(n13068), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n12731) );
  OAI211_X1 U15840 ( .C1(n12748), .C2(n12733), .A(n12732), .B(n12731), .ZN(
        n14278) );
  NAND2_X1 U15841 ( .A1(n14269), .A2(n14278), .ZN(n12734) );
  AOI22_X1 U15842 ( .A1(n12982), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13022), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12738) );
  AOI22_X1 U15843 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13050), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12737) );
  AOI22_X1 U15844 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13046), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12736) );
  AOI22_X1 U15845 ( .A1(n13045), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13048), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12735) );
  NAND4_X1 U15846 ( .A1(n12738), .A2(n12737), .A3(n12736), .A4(n12735), .ZN(
        n12744) );
  AOI22_X1 U15847 ( .A1(n13039), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13038), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12742) );
  AOI22_X1 U15848 ( .A1(n12443), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13049), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12741) );
  AOI22_X1 U15849 ( .A1(n13047), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12871), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12740) );
  AOI22_X1 U15850 ( .A1(n13040), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12739) );
  NAND4_X1 U15851 ( .A1(n12742), .A2(n12741), .A3(n12740), .A4(n12739), .ZN(
        n12743) );
  NOR2_X1 U15852 ( .A1(n12744), .A2(n12743), .ZN(n12749) );
  XNOR2_X1 U15853 ( .A(n12750), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14928) );
  NAND2_X1 U15854 ( .A1(n14928), .A2(n13920), .ZN(n12747) );
  AOI22_X1 U15855 ( .A1(n13068), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n13067), 
        .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12746) );
  OAI211_X1 U15856 ( .C1(n12749), .C2(n12748), .A(n12747), .B(n12746), .ZN(
        n14242) );
  NAND2_X1 U15857 ( .A1(n14239), .A2(n14242), .ZN(n14240) );
  AOI21_X1 U15858 ( .B1(n15852), .B2(n12751), .A(n12784), .ZN(n15910) );
  OR2_X1 U15859 ( .A1(n15910), .A2(n13063), .ZN(n12767) );
  AOI22_X1 U15860 ( .A1(n13022), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13040), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12755) );
  AOI22_X1 U15861 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13046), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12754) );
  AOI22_X1 U15862 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12871), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12753) );
  AOI22_X1 U15863 ( .A1(n12443), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12853), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12752) );
  NAND4_X1 U15864 ( .A1(n12755), .A2(n12754), .A3(n12753), .A4(n12752), .ZN(
        n12762) );
  AOI22_X1 U15865 ( .A1(n12982), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12594), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12759) );
  AOI22_X1 U15866 ( .A1(n13047), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12983), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12758) );
  AOI22_X1 U15867 ( .A1(n13038), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13048), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12757) );
  AOI22_X1 U15868 ( .A1(n13039), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12756) );
  NAND4_X1 U15869 ( .A1(n12759), .A2(n12758), .A3(n12757), .A4(n12756), .ZN(
        n12761) );
  OAI21_X1 U15870 ( .B1(n12762), .B2(n12761), .A(n12760), .ZN(n12765) );
  NAND2_X1 U15871 ( .A1(n13068), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12764) );
  NAND2_X1 U15872 ( .A1(n13067), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12763) );
  AND3_X1 U15873 ( .A1(n12765), .A2(n12764), .A3(n12763), .ZN(n12766) );
  NOR2_X2 U15874 ( .A1(n14240), .A2(n14302), .ZN(n14301) );
  INV_X1 U15875 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15841) );
  XNOR2_X1 U15876 ( .A(n12784), .B(n15841), .ZN(n15846) );
  NAND2_X1 U15877 ( .A1(n15846), .A2(n13920), .ZN(n12782) );
  AOI22_X1 U15878 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13047), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12771) );
  AOI22_X1 U15879 ( .A1(n12982), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13050), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12770) );
  AOI22_X1 U15880 ( .A1(n12443), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12853), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12769) );
  AOI22_X1 U15881 ( .A1(n13038), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13048), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12768) );
  NAND4_X1 U15882 ( .A1(n12771), .A2(n12770), .A3(n12769), .A4(n12768), .ZN(
        n12777) );
  AOI22_X1 U15883 ( .A1(n13022), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12983), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12775) );
  AOI22_X1 U15884 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13046), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12774) );
  AOI22_X1 U15885 ( .A1(n13040), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12871), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12773) );
  AOI22_X1 U15886 ( .A1(n13039), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12772) );
  NAND4_X1 U15887 ( .A1(n12775), .A2(n12774), .A3(n12773), .A4(n12772), .ZN(
        n12776) );
  NOR2_X1 U15888 ( .A1(n12777), .A2(n12776), .ZN(n12780) );
  AOI21_X1 U15889 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15841), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12778) );
  AOI21_X1 U15890 ( .B1(n12525), .B2(P1_EAX_REG_16__SCAN_IN), .A(n12778), .ZN(
        n12779) );
  OAI21_X1 U15891 ( .B1(n13033), .B2(n12780), .A(n12779), .ZN(n12781) );
  NAND2_X1 U15892 ( .A1(n12782), .A2(n12781), .ZN(n14761) );
  XNOR2_X1 U15893 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n12797), .ZN(
        n14686) );
  AOI22_X1 U15894 ( .A1(n13068), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n13067), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12796) );
  AOI22_X1 U15895 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13022), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12788) );
  AOI22_X1 U15896 ( .A1(n12982), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12871), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12787) );
  AOI22_X1 U15897 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13048), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12786) );
  AOI22_X1 U15898 ( .A1(n12491), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12853), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12785) );
  NAND4_X1 U15899 ( .A1(n12788), .A2(n12787), .A3(n12786), .A4(n12785), .ZN(
        n12794) );
  AOI22_X1 U15900 ( .A1(n13047), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13038), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12792) );
  AOI22_X1 U15901 ( .A1(n13039), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12490), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12791) );
  AOI22_X1 U15902 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13046), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12790) );
  AOI22_X1 U15903 ( .A1(n13040), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12789) );
  NAND4_X1 U15904 ( .A1(n12792), .A2(n12791), .A3(n12790), .A4(n12789), .ZN(
        n12793) );
  INV_X1 U15905 ( .A(n13033), .ZN(n13059) );
  OAI21_X1 U15906 ( .B1(n12794), .B2(n12793), .A(n13059), .ZN(n12795) );
  OAI211_X1 U15907 ( .C1(n14686), .C2(n13063), .A(n12796), .B(n12795), .ZN(
        n14682) );
  INV_X1 U15908 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14687) );
  AOI21_X1 U15909 ( .B1(n12798), .B2(n20923), .A(n12827), .ZN(n15837) );
  AOI22_X1 U15910 ( .A1(n13068), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n20708), .ZN(n12812) );
  AOI22_X1 U15911 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13050), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12802) );
  AOI22_X1 U15912 ( .A1(n12982), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13046), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12801) );
  AOI22_X1 U15913 ( .A1(n13022), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12871), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12800) );
  AOI22_X1 U15914 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12853), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12799) );
  NAND4_X1 U15915 ( .A1(n12802), .A2(n12801), .A3(n12800), .A4(n12799), .ZN(
        n12810) );
  AOI22_X1 U15916 ( .A1(n13040), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12983), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12808) );
  AOI21_X1 U15917 ( .B1(n12443), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n12508), .ZN(n12804) );
  NAND2_X1 U15918 ( .A1(n13047), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n12803) );
  AND2_X1 U15919 ( .A1(n12804), .A2(n12803), .ZN(n12807) );
  AOI22_X1 U15920 ( .A1(n13039), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12984), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12806) );
  AOI22_X1 U15921 ( .A1(n13038), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12805) );
  NAND4_X1 U15922 ( .A1(n12808), .A2(n12807), .A3(n12806), .A4(n12805), .ZN(
        n12809) );
  NAND2_X1 U15923 ( .A1(n13033), .A2(n13063), .ZN(n12876) );
  OAI21_X1 U15924 ( .B1(n12810), .B2(n12809), .A(n12876), .ZN(n12811) );
  AOI22_X1 U15925 ( .A1(n15837), .A2(n12508), .B1(n12812), .B2(n12811), .ZN(
        n14752) );
  AOI22_X1 U15926 ( .A1(n12982), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13047), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12816) );
  AOI22_X1 U15927 ( .A1(n13039), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13038), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12815) );
  AOI22_X1 U15928 ( .A1(n13040), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13050), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12814) );
  AOI22_X1 U15929 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12984), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12813) );
  NAND4_X1 U15930 ( .A1(n12816), .A2(n12815), .A3(n12814), .A4(n12813), .ZN(
        n12822) );
  AOI22_X1 U15931 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12983), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12820) );
  AOI22_X1 U15932 ( .A1(n13046), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12871), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12819) );
  AOI22_X1 U15933 ( .A1(n12443), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12853), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12818) );
  AOI22_X1 U15934 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12817) );
  NAND4_X1 U15935 ( .A1(n12820), .A2(n12819), .A3(n12818), .A4(n12817), .ZN(
        n12821) );
  NOR2_X1 U15936 ( .A1(n12822), .A2(n12821), .ZN(n12826) );
  OAI21_X1 U15937 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n20200), .A(
        n20708), .ZN(n12823) );
  INV_X1 U15938 ( .A(n12823), .ZN(n12824) );
  AOI21_X1 U15939 ( .B1(n12525), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12824), .ZN(
        n12825) );
  OAI21_X1 U15940 ( .B1(n13033), .B2(n12826), .A(n12825), .ZN(n12829) );
  OAI21_X1 U15941 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n12827), .A(
        n12846), .ZN(n15890) );
  OR2_X1 U15942 ( .A1(n13063), .A2(n15890), .ZN(n12828) );
  NAND2_X1 U15943 ( .A1(n12829), .A2(n12828), .ZN(n14748) );
  AOI22_X1 U15944 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n12496), .B1(
        n13047), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12833) );
  AOI22_X1 U15945 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n9829), .B1(
        n13046), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12832) );
  AOI22_X1 U15946 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n13045), .B1(
        n12984), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12831) );
  AOI22_X1 U15947 ( .A1(n12982), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12853), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12830) );
  NAND4_X1 U15948 ( .A1(n12833), .A2(n12832), .A3(n12831), .A4(n12830), .ZN(
        n12841) );
  AOI22_X1 U15949 ( .A1(n13039), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13038), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12839) );
  AOI22_X1 U15950 ( .A1(n13040), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13050), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12838) );
  AOI22_X1 U15951 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12837) );
  NAND2_X1 U15952 ( .A1(n12871), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12835) );
  NAND2_X1 U15953 ( .A1(n12443), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12834) );
  AND3_X1 U15954 ( .A1(n12835), .A2(n12834), .A3(n13063), .ZN(n12836) );
  NAND4_X1 U15955 ( .A1(n12839), .A2(n12838), .A3(n12837), .A4(n12836), .ZN(
        n12840) );
  OAI21_X1 U15956 ( .B1(n12841), .B2(n12840), .A(n12876), .ZN(n12843) );
  AOI22_X1 U15957 ( .A1(n13068), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20708), .ZN(n12842) );
  NAND2_X1 U15958 ( .A1(n12843), .A2(n12842), .ZN(n12845) );
  XNOR2_X1 U15959 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n12846), .ZN(
        n15814) );
  NAND2_X1 U15960 ( .A1(n15814), .A2(n13920), .ZN(n12844) );
  NAND2_X1 U15961 ( .A1(n12845), .A2(n12844), .ZN(n14745) );
  INV_X1 U15962 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15824) );
  OR2_X1 U15963 ( .A1(n12847), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12848) );
  NAND2_X1 U15964 ( .A1(n12848), .A2(n12884), .ZN(n15883) );
  INV_X1 U15965 ( .A(n15883), .ZN(n12864) );
  AOI22_X1 U15966 ( .A1(n12982), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13038), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12852) );
  AOI22_X1 U15967 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13040), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12851) );
  AOI22_X1 U15968 ( .A1(n13046), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12850) );
  AOI22_X1 U15969 ( .A1(n13047), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12984), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12849) );
  NAND4_X1 U15970 ( .A1(n12852), .A2(n12851), .A3(n12850), .A4(n12849), .ZN(
        n12859) );
  AOI22_X1 U15971 ( .A1(n13039), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13050), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12857) );
  AOI22_X1 U15972 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12983), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12856) );
  AOI22_X1 U15973 ( .A1(n12496), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12871), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12855) );
  AOI22_X1 U15974 ( .A1(n12443), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12853), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12854) );
  NAND4_X1 U15975 ( .A1(n12857), .A2(n12856), .A3(n12855), .A4(n12854), .ZN(
        n12858) );
  OR2_X1 U15976 ( .A1(n12859), .A2(n12858), .ZN(n12862) );
  INV_X1 U15977 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n14809) );
  NAND2_X1 U15978 ( .A1(n20708), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12860) );
  OAI211_X1 U15979 ( .C1(n12909), .C2(n14809), .A(n13063), .B(n12860), .ZN(
        n12861) );
  AOI21_X1 U15980 ( .B1(n13059), .B2(n12862), .A(n12861), .ZN(n12863) );
  AOI21_X1 U15981 ( .B1(n12864), .B2(n13920), .A(n12863), .ZN(n14737) );
  AOI22_X1 U15982 ( .A1(n13047), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13038), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12868) );
  AOI22_X1 U15983 ( .A1(n13040), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12490), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12867) );
  AOI22_X1 U15984 ( .A1(n12337), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13049), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12866) );
  AOI22_X1 U15985 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13048), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12865) );
  NAND4_X1 U15986 ( .A1(n12868), .A2(n12867), .A3(n12866), .A4(n12865), .ZN(
        n12878) );
  AOI22_X1 U15987 ( .A1(n13039), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13050), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12875) );
  AOI21_X1 U15988 ( .B1(n12491), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n12508), .ZN(n12870) );
  NAND2_X1 U15989 ( .A1(n13022), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12869) );
  AND2_X1 U15990 ( .A1(n12870), .A2(n12869), .ZN(n12874) );
  AOI22_X1 U15991 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13046), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12873) );
  AOI22_X1 U15992 ( .A1(n12871), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12872) );
  NAND4_X1 U15993 ( .A1(n12875), .A2(n12874), .A3(n12873), .A4(n12872), .ZN(
        n12877) );
  OAI21_X1 U15994 ( .B1(n12878), .B2(n12877), .A(n12876), .ZN(n12880) );
  AOI22_X1 U15995 ( .A1(n13068), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20708), .ZN(n12879) );
  NAND2_X1 U15996 ( .A1(n12880), .A2(n12879), .ZN(n12882) );
  XNOR2_X1 U15997 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B(n12884), .ZN(
        n15798) );
  NAND2_X1 U15998 ( .A1(n15798), .A2(n13920), .ZN(n12881) );
  NAND2_X1 U15999 ( .A1(n12882), .A2(n12881), .ZN(n14734) );
  INV_X1 U16000 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12883) );
  OR2_X1 U16001 ( .A1(n12885), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12886) );
  NAND2_X1 U16002 ( .A1(n12886), .A2(n12928), .ZN(n15878) );
  AOI22_X1 U16003 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13050), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12890) );
  AOI22_X1 U16004 ( .A1(n13040), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12983), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12889) );
  AOI22_X1 U16005 ( .A1(n13047), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13048), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12888) );
  AOI22_X1 U16006 ( .A1(n12982), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12887) );
  NAND4_X1 U16007 ( .A1(n12890), .A2(n12889), .A3(n12888), .A4(n12887), .ZN(
        n12896) );
  AOI22_X1 U16008 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13038), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12894) );
  AOI22_X1 U16009 ( .A1(n13039), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13046), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12893) );
  AOI22_X1 U16010 ( .A1(n13022), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12871), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12892) );
  AOI22_X1 U16011 ( .A1(n12443), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13049), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12891) );
  NAND4_X1 U16012 ( .A1(n12894), .A2(n12893), .A3(n12892), .A4(n12891), .ZN(
        n12895) );
  NOR2_X1 U16013 ( .A1(n12896), .A2(n12895), .ZN(n12913) );
  AOI22_X1 U16014 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13047), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12900) );
  AOI22_X1 U16015 ( .A1(n13039), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13038), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12899) );
  AOI22_X1 U16016 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12898) );
  AOI22_X1 U16017 ( .A1(n13040), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12871), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12897) );
  NAND4_X1 U16018 ( .A1(n12900), .A2(n12899), .A3(n12898), .A4(n12897), .ZN(
        n12906) );
  AOI22_X1 U16019 ( .A1(n13022), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12983), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12904) );
  AOI22_X1 U16020 ( .A1(n12982), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13046), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12903) );
  AOI22_X1 U16021 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13048), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12902) );
  AOI22_X1 U16022 ( .A1(n12443), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13049), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12901) );
  NAND4_X1 U16023 ( .A1(n12904), .A2(n12903), .A3(n12902), .A4(n12901), .ZN(
        n12905) );
  NOR2_X1 U16024 ( .A1(n12906), .A2(n12905), .ZN(n12914) );
  XNOR2_X1 U16025 ( .A(n12913), .B(n12914), .ZN(n12907) );
  NOR2_X1 U16026 ( .A1(n12907), .A2(n13033), .ZN(n12911) );
  INV_X1 U16027 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14798) );
  NAND2_X1 U16028 ( .A1(n20708), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12908) );
  OAI211_X1 U16029 ( .C1(n12909), .C2(n14798), .A(n13063), .B(n12908), .ZN(
        n12910) );
  OAI22_X1 U16030 ( .A1(n15878), .A2(n13063), .B1(n12911), .B2(n12910), .ZN(
        n14727) );
  NAND2_X1 U16031 ( .A1(n14725), .A2(n12912), .ZN(n14719) );
  NOR2_X1 U16032 ( .A1(n12914), .A2(n12913), .ZN(n12944) );
  AOI22_X1 U16033 ( .A1(n12982), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13039), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12918) );
  AOI22_X1 U16034 ( .A1(n13038), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12490), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12917) );
  AOI22_X1 U16035 ( .A1(n12443), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13049), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12916) );
  AOI22_X1 U16036 ( .A1(n13046), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12915) );
  NAND4_X1 U16037 ( .A1(n12918), .A2(n12917), .A3(n12916), .A4(n12915), .ZN(
        n12924) );
  AOI22_X1 U16038 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13047), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12922) );
  AOI22_X1 U16039 ( .A1(n13040), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13045), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12921) );
  AOI22_X1 U16040 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12871), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12920) );
  AOI22_X1 U16041 ( .A1(n13022), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13048), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12919) );
  NAND4_X1 U16042 ( .A1(n12922), .A2(n12921), .A3(n12920), .A4(n12919), .ZN(
        n12923) );
  OR2_X1 U16043 ( .A1(n12924), .A2(n12923), .ZN(n12943) );
  XNOR2_X1 U16044 ( .A(n12944), .B(n12943), .ZN(n12927) );
  INV_X1 U16045 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n20903) );
  AOI21_X1 U16046 ( .B1(n20903), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12925) );
  AOI21_X1 U16047 ( .B1(n12525), .B2(P1_EAX_REG_24__SCAN_IN), .A(n12925), .ZN(
        n12926) );
  OAI21_X1 U16048 ( .B1(n12927), .B2(n13033), .A(n12926), .ZN(n12932) );
  NOR2_X1 U16049 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n12929), .ZN(
        n12930) );
  NOR2_X1 U16050 ( .A1(n12949), .A2(n12930), .ZN(n15786) );
  NAND2_X1 U16051 ( .A1(n15786), .A2(n13920), .ZN(n12931) );
  NAND2_X1 U16052 ( .A1(n12932), .A2(n12931), .ZN(n14720) );
  AOI22_X1 U16053 ( .A1(n13047), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13022), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12936) );
  AOI22_X1 U16054 ( .A1(n13039), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13038), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12935) );
  AOI22_X1 U16055 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13045), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12934) );
  AOI22_X1 U16056 ( .A1(n13040), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12933) );
  NAND4_X1 U16057 ( .A1(n12936), .A2(n12935), .A3(n12934), .A4(n12933), .ZN(
        n12942) );
  AOI22_X1 U16058 ( .A1(n12982), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13050), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12940) );
  AOI22_X1 U16059 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12871), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12939) );
  AOI22_X1 U16060 ( .A1(n13046), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13048), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12938) );
  AOI22_X1 U16061 ( .A1(n12491), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13049), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12937) );
  NAND4_X1 U16062 ( .A1(n12940), .A2(n12939), .A3(n12938), .A4(n12937), .ZN(
        n12941) );
  NOR2_X1 U16063 ( .A1(n12942), .A2(n12941), .ZN(n12959) );
  NAND2_X1 U16064 ( .A1(n12944), .A2(n12943), .ZN(n12958) );
  XNOR2_X1 U16065 ( .A(n12959), .B(n12958), .ZN(n12948) );
  NAND2_X1 U16066 ( .A1(n20708), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12945) );
  NAND2_X1 U16067 ( .A1(n13063), .A2(n12945), .ZN(n12946) );
  AOI21_X1 U16068 ( .B1(n12525), .B2(P1_EAX_REG_25__SCAN_IN), .A(n12946), .ZN(
        n12947) );
  OAI21_X1 U16069 ( .B1(n12948), .B2(n13033), .A(n12947), .ZN(n12954) );
  INV_X1 U16070 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12951) );
  INV_X1 U16071 ( .A(n12949), .ZN(n12950) );
  NAND2_X1 U16072 ( .A1(n12951), .A2(n12950), .ZN(n12952) );
  NAND2_X1 U16073 ( .A1(n12956), .A2(n12952), .ZN(n15779) );
  INV_X1 U16074 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n20887) );
  NAND2_X1 U16075 ( .A1(n12956), .A2(n20887), .ZN(n12957) );
  OAI21_X1 U16076 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20887), .A(n13063), 
        .ZN(n12972) );
  NOR2_X1 U16077 ( .A1(n12959), .A2(n12958), .ZN(n12992) );
  AOI22_X1 U16078 ( .A1(n12337), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13039), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12963) );
  AOI22_X1 U16079 ( .A1(n13038), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12490), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12962) );
  AOI22_X1 U16080 ( .A1(n12491), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13049), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12961) );
  AOI22_X1 U16081 ( .A1(n13046), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12960) );
  NAND4_X1 U16082 ( .A1(n12963), .A2(n12962), .A3(n12961), .A4(n12960), .ZN(
        n12969) );
  AOI22_X1 U16083 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13047), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12967) );
  AOI22_X1 U16084 ( .A1(n13040), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13045), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12966) );
  AOI22_X1 U16085 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12871), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12965) );
  AOI22_X1 U16086 ( .A1(n13022), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13048), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12964) );
  NAND4_X1 U16087 ( .A1(n12967), .A2(n12966), .A3(n12965), .A4(n12964), .ZN(
        n12968) );
  OR2_X1 U16088 ( .A1(n12969), .A2(n12968), .ZN(n12991) );
  XNOR2_X1 U16089 ( .A(n12992), .B(n12991), .ZN(n12970) );
  NOR2_X1 U16090 ( .A1(n12970), .A2(n13033), .ZN(n12971) );
  AOI211_X1 U16091 ( .C1(n12525), .C2(P1_EAX_REG_26__SCAN_IN), .A(n12972), .B(
        n12971), .ZN(n12973) );
  INV_X1 U16092 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12975) );
  NAND2_X1 U16093 ( .A1(n12976), .A2(n12975), .ZN(n12977) );
  NAND2_X1 U16094 ( .A1(n12997), .A2(n12977), .ZN(n14866) );
  AOI22_X1 U16095 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n12496), .B1(
        n13047), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12981) );
  AOI22_X1 U16096 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13050), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12980) );
  AOI22_X1 U16097 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n9829), .B1(
        n13046), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12979) );
  AOI22_X1 U16098 ( .A1(n13039), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12978) );
  NAND4_X1 U16099 ( .A1(n12981), .A2(n12980), .A3(n12979), .A4(n12978), .ZN(
        n12990) );
  AOI22_X1 U16100 ( .A1(n12982), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13040), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12988) );
  AOI22_X1 U16101 ( .A1(n13038), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12983), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12987) );
  AOI22_X1 U16102 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n12984), .B1(
        n12871), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12986) );
  AOI22_X1 U16103 ( .A1(n12491), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13049), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12985) );
  NAND4_X1 U16104 ( .A1(n12988), .A2(n12987), .A3(n12986), .A4(n12985), .ZN(
        n12989) );
  NOR2_X1 U16105 ( .A1(n12990), .A2(n12989), .ZN(n13000) );
  NAND2_X1 U16106 ( .A1(n12992), .A2(n12991), .ZN(n12999) );
  XNOR2_X1 U16107 ( .A(n13000), .B(n12999), .ZN(n12995) );
  AOI21_X1 U16108 ( .B1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n20708), .A(
        n13920), .ZN(n12994) );
  NAND2_X1 U16109 ( .A1(n13068), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n12993) );
  OAI211_X1 U16110 ( .C1(n12995), .C2(n13033), .A(n12994), .B(n12993), .ZN(
        n12996) );
  INV_X1 U16111 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n20977) );
  NAND2_X1 U16112 ( .A1(n12997), .A2(n20977), .ZN(n12998) );
  AOI21_X1 U16113 ( .B1(n20977), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13013) );
  NOR2_X1 U16114 ( .A1(n13000), .A2(n12999), .ZN(n13030) );
  AOI22_X1 U16115 ( .A1(n12337), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13039), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13004) );
  AOI22_X1 U16116 ( .A1(n13038), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12490), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13003) );
  AOI22_X1 U16117 ( .A1(n12491), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13049), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13002) );
  AOI22_X1 U16118 ( .A1(n13046), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13001) );
  NAND4_X1 U16119 ( .A1(n13004), .A2(n13003), .A3(n13002), .A4(n13001), .ZN(
        n13010) );
  AOI22_X1 U16120 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13047), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13008) );
  AOI22_X1 U16121 ( .A1(n13040), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13045), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13007) );
  AOI22_X1 U16122 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12871), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13006) );
  AOI22_X1 U16123 ( .A1(n13022), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13048), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13005) );
  NAND4_X1 U16124 ( .A1(n13008), .A2(n13007), .A3(n13006), .A4(n13005), .ZN(
        n13009) );
  OR2_X1 U16125 ( .A1(n13010), .A2(n13009), .ZN(n13029) );
  XNOR2_X1 U16126 ( .A(n13030), .B(n13029), .ZN(n13011) );
  NOR2_X1 U16127 ( .A1(n13011), .A2(n13033), .ZN(n13012) );
  AOI211_X1 U16128 ( .C1(n13068), .C2(P1_EAX_REG_28__SCAN_IN), .A(n13013), .B(
        n13012), .ZN(n13014) );
  INV_X1 U16129 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n13015) );
  NAND2_X1 U16130 ( .A1(n13016), .A2(n13015), .ZN(n13017) );
  NAND2_X1 U16131 ( .A1(n13256), .A2(n13017), .ZN(n14846) );
  AOI22_X1 U16132 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13046), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13021) );
  AOI22_X1 U16133 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13048), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13020) );
  AOI22_X1 U16134 ( .A1(n12337), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13019) );
  AOI22_X1 U16135 ( .A1(n13038), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13018) );
  NAND4_X1 U16136 ( .A1(n13021), .A2(n13020), .A3(n13019), .A4(n13018), .ZN(
        n13028) );
  AOI22_X1 U16137 ( .A1(n13047), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13040), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13026) );
  AOI22_X1 U16138 ( .A1(n13022), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13045), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13025) );
  AOI22_X1 U16139 ( .A1(n13039), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12871), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13024) );
  AOI22_X1 U16140 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13049), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13023) );
  NAND4_X1 U16141 ( .A1(n13026), .A2(n13025), .A3(n13024), .A4(n13023), .ZN(
        n13027) );
  NOR2_X1 U16142 ( .A1(n13028), .A2(n13027), .ZN(n13037) );
  NAND2_X1 U16143 ( .A1(n13030), .A2(n13029), .ZN(n13036) );
  XNOR2_X1 U16144 ( .A(n13037), .B(n13036), .ZN(n13034) );
  AOI21_X1 U16145 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20708), .A(
        n13920), .ZN(n13032) );
  NAND2_X1 U16146 ( .A1(n13068), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n13031) );
  OAI211_X1 U16147 ( .C1(n13034), .C2(n13033), .A(n13032), .B(n13031), .ZN(
        n13035) );
  OAI21_X1 U16148 ( .B1(n13063), .B2(n14846), .A(n13035), .ZN(n14637) );
  NOR2_X1 U16149 ( .A1(n13037), .A2(n13036), .ZN(n13058) );
  AOI22_X1 U16150 ( .A1(n13039), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13038), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13044) );
  AOI22_X1 U16151 ( .A1(n12337), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12491), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13043) );
  AOI22_X1 U16152 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12871), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13042) );
  AOI22_X1 U16153 ( .A1(n13040), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13041) );
  NAND4_X1 U16154 ( .A1(n13044), .A2(n13043), .A3(n13042), .A4(n13041), .ZN(
        n13056) );
  AOI22_X1 U16155 ( .A1(n12490), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13045), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13054) );
  AOI22_X1 U16156 ( .A1(n13047), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13046), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13053) );
  AOI22_X1 U16157 ( .A1(n13022), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13048), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13052) );
  AOI22_X1 U16158 ( .A1(n13050), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13049), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13051) );
  NAND4_X1 U16159 ( .A1(n13054), .A2(n13053), .A3(n13052), .A4(n13051), .ZN(
        n13055) );
  NOR2_X1 U16160 ( .A1(n13056), .A2(n13055), .ZN(n13057) );
  XNOR2_X1 U16161 ( .A(n13058), .B(n13057), .ZN(n13060) );
  NAND2_X1 U16162 ( .A1(n13060), .A2(n13059), .ZN(n13066) );
  NAND2_X1 U16163 ( .A1(n20708), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13061) );
  NAND2_X1 U16164 ( .A1(n13063), .A2(n13061), .ZN(n13062) );
  AOI21_X1 U16165 ( .B1(n13068), .B2(P1_EAX_REG_30__SCAN_IN), .A(n13062), .ZN(
        n13065) );
  INV_X1 U16166 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14627) );
  XNOR2_X1 U16167 ( .A(n13256), .B(n14627), .ZN(n14837) );
  NOR2_X1 U16168 ( .A1(n14837), .A2(n13063), .ZN(n13064) );
  AOI21_X1 U16169 ( .B1(n13066), .B2(n13065), .A(n13064), .ZN(n14391) );
  AOI22_X1 U16170 ( .A1(n13068), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n13067), .ZN(n13069) );
  INV_X1 U16171 ( .A(n13069), .ZN(n13070) );
  XNOR2_X1 U16172 ( .A(n13071), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n13085) );
  INV_X1 U16173 ( .A(n13085), .ZN(n13073) );
  NAND2_X1 U16174 ( .A1(n20563), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13084) );
  INV_X1 U16175 ( .A(n13084), .ZN(n13072) );
  NAND2_X1 U16176 ( .A1(n13073), .A2(n13072), .ZN(n13086) );
  NAND2_X1 U16177 ( .A1(n20638), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13074) );
  NAND2_X1 U16178 ( .A1(n13086), .A2(n13074), .ZN(n13083) );
  XNOR2_X1 U16179 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n13082) );
  NAND2_X1 U16180 ( .A1(n13083), .A2(n13082), .ZN(n13076) );
  NAND2_X1 U16181 ( .A1(n20398), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13075) );
  NAND2_X1 U16182 ( .A1(n13076), .A2(n13075), .ZN(n13102) );
  XNOR2_X1 U16183 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n13101) );
  INV_X1 U16184 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20116) );
  NOR2_X1 U16185 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20116), .ZN(
        n13077) );
  INV_X1 U16186 ( .A(n13109), .ZN(n13078) );
  NAND2_X1 U16187 ( .A1(n13138), .A2(n13079), .ZN(n13120) );
  OAI22_X1 U16188 ( .A1(n13092), .A2(n20139), .B1(n20706), .B2(n20154), .ZN(
        n13095) );
  NOR2_X1 U16189 ( .A1(n20139), .A2(n13095), .ZN(n13112) );
  NAND3_X1 U16190 ( .A1(n13738), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(
        n13081), .ZN(n13136) );
  XNOR2_X1 U16191 ( .A(n13083), .B(n13082), .ZN(n13134) );
  AOI21_X1 U16192 ( .B1(n20139), .B2(n20154), .A(n13131), .ZN(n13089) );
  INV_X1 U16193 ( .A(n13089), .ZN(n13105) );
  NAND2_X1 U16194 ( .A1(n13085), .A2(n13084), .ZN(n13087) );
  NAND2_X1 U16195 ( .A1(n13087), .A2(n13086), .ZN(n13135) );
  INV_X1 U16196 ( .A(n13135), .ZN(n13088) );
  NOR2_X1 U16197 ( .A1(n13088), .A2(n13112), .ZN(n13098) );
  XNOR2_X1 U16198 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n13090) );
  OAI211_X1 U16199 ( .C1(n20124), .C2(n13125), .A(n13089), .B(n13090), .ZN(
        n13094) );
  INV_X1 U16200 ( .A(n13090), .ZN(n13091) );
  OAI21_X1 U16201 ( .B1(n13092), .B2(n13091), .A(n13109), .ZN(n13093) );
  NAND2_X1 U16202 ( .A1(n13094), .A2(n13093), .ZN(n13097) );
  NOR2_X1 U16203 ( .A1(n13098), .A2(n13097), .ZN(n13100) );
  AOI21_X1 U16204 ( .B1(n13108), .B2(n13135), .A(n13095), .ZN(n13096) );
  AOI21_X1 U16205 ( .B1(n13098), .B2(n13097), .A(n13096), .ZN(n13099) );
  AOI211_X1 U16206 ( .C1(n13106), .C2(n13105), .A(n13100), .B(n13099), .ZN(
        n13111) );
  NOR2_X1 U16207 ( .A1(n13102), .A2(n13101), .ZN(n13103) );
  NOR2_X1 U16208 ( .A1(n13104), .A2(n13103), .ZN(n13132) );
  AOI22_X1 U16209 ( .A1(n13108), .A2(n13134), .B1(n13132), .B2(n13107), .ZN(
        n13110) );
  OAI22_X1 U16210 ( .A1(n13111), .A2(n13110), .B1(n13132), .B2(n13109), .ZN(
        n13113) );
  AOI21_X1 U16211 ( .B1(n13112), .B2(n13115), .A(n13113), .ZN(n13117) );
  INV_X1 U16212 ( .A(n13113), .ZN(n13114) );
  OAI22_X1 U16213 ( .A1(n13117), .A2(n13116), .B1(n13115), .B2(n13114), .ZN(
        n13118) );
  AOI21_X1 U16214 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20706), .A(
        n13118), .ZN(n13119) );
  NAND2_X1 U16215 ( .A1(n13120), .A2(n13119), .ZN(n13121) );
  NAND2_X1 U16216 ( .A1(n15736), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n19875) );
  NAND2_X1 U16217 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20818) );
  INV_X1 U16218 ( .A(n20818), .ZN(n15760) );
  OR2_X1 U16219 ( .A1(n13123), .A2(n15760), .ZN(n20012) );
  INV_X1 U16220 ( .A(n13124), .ZN(n13127) );
  OR2_X1 U16221 ( .A1(n13125), .A2(n13141), .ZN(n13126) );
  AND2_X1 U16222 ( .A1(n13127), .A2(n13126), .ZN(n13535) );
  INV_X1 U16223 ( .A(n13128), .ZN(n13130) );
  NAND2_X1 U16224 ( .A1(n15156), .A2(n20124), .ZN(n13129) );
  NAND2_X1 U16225 ( .A1(n13504), .A2(n13131), .ZN(n14601) );
  INV_X1 U16226 ( .A(n13132), .ZN(n13133) );
  NOR3_X1 U16227 ( .A1(n13135), .A2(n13134), .A3(n13133), .ZN(n13137) );
  OAI21_X1 U16228 ( .B1(n13138), .B2(n13137), .A(n13136), .ZN(n14607) );
  NOR2_X1 U16229 ( .A1(n13139), .A2(n15760), .ZN(n13140) );
  NAND2_X1 U16230 ( .A1(n14607), .A2(n13140), .ZN(n13506) );
  NAND4_X1 U16231 ( .A1(n14452), .A2(n20150), .A3(n13141), .A4(n14611), .ZN(
        n13560) );
  OAI22_X1 U16232 ( .A1(n13506), .A2(n19875), .B1(n13547), .B2(n13560), .ZN(
        n13142) );
  INV_X1 U16233 ( .A(n13142), .ZN(n13143) );
  NAND3_X1 U16234 ( .A1(n14625), .A2(n14452), .A3(n14808), .ZN(n13161) );
  NOR4_X1 U16235 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(
        P1_ADDRESS_REG_15__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_13__SCAN_IN), .ZN(n13148) );
  NOR4_X1 U16236 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(
        P1_ADDRESS_REG_19__SCAN_IN), .A3(P1_ADDRESS_REG_18__SCAN_IN), .A4(
        P1_ADDRESS_REG_17__SCAN_IN), .ZN(n13147) );
  NOR4_X1 U16237 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(
        P1_ADDRESS_REG_6__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13146) );
  NOR4_X1 U16238 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(
        P1_ADDRESS_REG_10__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n13145) );
  AND4_X1 U16239 ( .A1(n13148), .A2(n13147), .A3(n13146), .A4(n13145), .ZN(
        n13153) );
  NOR4_X1 U16240 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_5__SCAN_IN), .A4(
        P1_ADDRESS_REG_12__SCAN_IN), .ZN(n13151) );
  NOR4_X1 U16241 ( .A1(P1_ADDRESS_REG_25__SCAN_IN), .A2(
        P1_ADDRESS_REG_24__SCAN_IN), .A3(P1_ADDRESS_REG_23__SCAN_IN), .A4(
        P1_ADDRESS_REG_21__SCAN_IN), .ZN(n13150) );
  NOR4_X1 U16242 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_28__SCAN_IN), .A3(P1_ADDRESS_REG_27__SCAN_IN), .A4(
        P1_ADDRESS_REG_26__SCAN_IN), .ZN(n13149) );
  INV_X1 U16243 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20728) );
  AND4_X1 U16244 ( .A1(n13151), .A2(n13150), .A3(n13149), .A4(n20728), .ZN(
        n13152) );
  NAND2_X1 U16245 ( .A1(n13153), .A2(n13152), .ZN(n13154) );
  NOR3_X1 U16246 ( .A1(n14827), .A2(n20117), .A3(n13599), .ZN(n13155) );
  AOI22_X1 U16247 ( .A1(n14829), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14827), .ZN(n13156) );
  INV_X1 U16248 ( .A(n13156), .ZN(n13159) );
  NOR2_X1 U16249 ( .A1(n13599), .A2(n20119), .ZN(n13157) );
  NAND2_X1 U16250 ( .A1(n14808), .A2(n13157), .ZN(n14810) );
  INV_X1 U16251 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n19197) );
  NOR2_X1 U16252 ( .A1(n14810), .A2(n19197), .ZN(n13158) );
  NOR2_X1 U16253 ( .A1(n13159), .A2(n13158), .ZN(n13160) );
  NAND2_X1 U16254 ( .A1(n13161), .A2(n13160), .ZN(P1_U2873) );
  INV_X1 U16255 ( .A(n13166), .ZN(n13162) );
  AND2_X1 U16256 ( .A1(n20124), .A2(n20146), .ZN(n13174) );
  AOI21_X1 U16257 ( .B1(n20009), .B2(n13162), .A(n13174), .ZN(n13163) );
  NOR2_X1 U16258 ( .A1(n13128), .A2(n13165), .ZN(n13169) );
  NAND2_X1 U16259 ( .A1(n13166), .A2(n13167), .ZN(n13180) );
  OAI211_X1 U16260 ( .C1(n13167), .C2(n13166), .A(n20009), .B(n13180), .ZN(
        n13168) );
  OAI211_X1 U16261 ( .C1(n13170), .C2(n20139), .A(n13169), .B(n13168), .ZN(
        n13171) );
  NAND2_X1 U16262 ( .A1(n13632), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13633) );
  INV_X1 U16263 ( .A(n13486), .ZN(n13172) );
  NAND2_X1 U16264 ( .A1(n13172), .A2(n13171), .ZN(n13173) );
  INV_X1 U16265 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20113) );
  XNOR2_X1 U16266 ( .A(n13180), .B(n13179), .ZN(n13175) );
  AOI21_X1 U16267 ( .B1(n20009), .B2(n13175), .A(n13174), .ZN(n13176) );
  NAND2_X1 U16268 ( .A1(n13702), .A2(n13701), .ZN(n13700) );
  NAND2_X1 U16269 ( .A1(n13177), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13178) );
  INV_X1 U16270 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20092) );
  OR2_X1 U16271 ( .A1(n20122), .A2(n13199), .ZN(n13184) );
  NAND2_X1 U16272 ( .A1(n13180), .A2(n13179), .ZN(n13197) );
  INV_X1 U16273 ( .A(n13194), .ZN(n13181) );
  XNOR2_X1 U16274 ( .A(n13197), .B(n13181), .ZN(n13182) );
  NAND2_X1 U16275 ( .A1(n13182), .A2(n20009), .ZN(n13183) );
  NAND2_X1 U16276 ( .A1(n13184), .A2(n13183), .ZN(n13788) );
  NAND2_X1 U16277 ( .A1(n13789), .A2(n13788), .ZN(n13787) );
  NAND2_X1 U16278 ( .A1(n13185), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13186) );
  NAND2_X1 U16279 ( .A1(n13787), .A2(n13186), .ZN(n20068) );
  OR2_X1 U16280 ( .A1(n13187), .A2(n13199), .ZN(n13191) );
  NAND2_X1 U16281 ( .A1(n13197), .A2(n13194), .ZN(n13188) );
  XNOR2_X1 U16282 ( .A(n13188), .B(n13195), .ZN(n13189) );
  NAND2_X1 U16283 ( .A1(n13189), .A2(n20009), .ZN(n13190) );
  NAND2_X1 U16284 ( .A1(n13191), .A2(n13190), .ZN(n13192) );
  INV_X1 U16285 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20084) );
  XNOR2_X1 U16286 ( .A(n13192), .B(n20084), .ZN(n20067) );
  NAND2_X1 U16287 ( .A1(n20068), .A2(n20067), .ZN(n20066) );
  NAND2_X1 U16288 ( .A1(n13192), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13193) );
  NAND2_X1 U16289 ( .A1(n20066), .A2(n13193), .ZN(n15943) );
  AND2_X1 U16290 ( .A1(n13195), .A2(n13194), .ZN(n13196) );
  AND2_X1 U16291 ( .A1(n13197), .A2(n13196), .ZN(n13205) );
  XNOR2_X1 U16292 ( .A(n13205), .B(n13204), .ZN(n13198) );
  INV_X1 U16293 ( .A(n20009), .ZN(n20812) );
  OAI22_X1 U16294 ( .A1(n13200), .A2(n13199), .B1(n13198), .B2(n20812), .ZN(
        n13201) );
  INV_X1 U16295 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16035) );
  XNOR2_X1 U16296 ( .A(n13201), .B(n16035), .ZN(n15942) );
  NAND2_X1 U16297 ( .A1(n13201), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13202) );
  NAND3_X1 U16298 ( .A1(n13224), .A2(n13221), .A3(n13203), .ZN(n13208) );
  NAND2_X1 U16299 ( .A1(n13205), .A2(n13204), .ZN(n13214) );
  XNOR2_X1 U16300 ( .A(n13213), .B(n13214), .ZN(n13206) );
  NAND2_X1 U16301 ( .A1(n20009), .A2(n13206), .ZN(n13207) );
  INV_X1 U16302 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15935) );
  NAND2_X1 U16303 ( .A1(n15936), .A2(n15935), .ZN(n13209) );
  INV_X1 U16304 ( .A(n15936), .ZN(n13210) );
  NAND2_X1 U16305 ( .A1(n13210), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13211) );
  NAND2_X1 U16306 ( .A1(n13212), .A2(n13221), .ZN(n13219) );
  INV_X1 U16307 ( .A(n13213), .ZN(n13215) );
  NOR2_X1 U16308 ( .A1(n13215), .A2(n13214), .ZN(n13227) );
  INV_X1 U16309 ( .A(n13227), .ZN(n13216) );
  XNOR2_X1 U16310 ( .A(n13226), .B(n13216), .ZN(n13217) );
  NAND2_X1 U16311 ( .A1(n20009), .A2(n13217), .ZN(n13218) );
  NAND2_X1 U16312 ( .A1(n13219), .A2(n13218), .ZN(n13220) );
  OR2_X1 U16313 ( .A1(n13220), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15930) );
  NAND2_X1 U16314 ( .A1(n13220), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15929) );
  AND2_X1 U16315 ( .A1(n13222), .A2(n13221), .ZN(n13223) );
  NAND3_X1 U16316 ( .A1(n20009), .A2(n13227), .A3(n13226), .ZN(n13228) );
  NAND2_X1 U16317 ( .A1(n13225), .A2(n13228), .ZN(n14099) );
  OR2_X1 U16318 ( .A1(n14099), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13229) );
  NAND2_X1 U16319 ( .A1(n14099), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13230) );
  INV_X1 U16320 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16006) );
  NAND2_X1 U16321 ( .A1(n13225), .A2(n16006), .ZN(n13231) );
  INV_X1 U16322 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15970) );
  INV_X1 U16323 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n13240) );
  NAND2_X1 U16324 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n13232) );
  INV_X1 U16325 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14244) );
  NAND2_X1 U16326 ( .A1(n13225), .A2(n14244), .ZN(n13233) );
  NAND2_X1 U16327 ( .A1(n14924), .A2(n13233), .ZN(n14913) );
  OR2_X1 U16328 ( .A1(n13225), .A2(n14244), .ZN(n13235) );
  NAND2_X1 U16329 ( .A1(n13234), .A2(n13235), .ZN(n15904) );
  INV_X1 U16330 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n13237) );
  NOR2_X1 U16331 ( .A1(n13225), .A2(n13237), .ZN(n13236) );
  NOR2_X1 U16332 ( .A1(n15904), .A2(n13236), .ZN(n13239) );
  XNOR2_X1 U16333 ( .A(n13225), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14917) );
  NAND2_X1 U16334 ( .A1(n13225), .A2(n13237), .ZN(n15907) );
  NAND2_X1 U16335 ( .A1(n14917), .A2(n15907), .ZN(n13238) );
  INV_X1 U16336 ( .A(n13239), .ZN(n15892) );
  NOR2_X1 U16337 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n13241) );
  NAND2_X1 U16338 ( .A1(n14937), .A2(n14934), .ZN(n14914) );
  NOR2_X1 U16339 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n13242) );
  NOR2_X1 U16340 ( .A1(n13225), .A2(n13242), .ZN(n13243) );
  XNOR2_X1 U16341 ( .A(n13225), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14909) );
  INV_X1 U16342 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n21010) );
  AND2_X1 U16343 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15074) );
  INV_X1 U16344 ( .A(n15074), .ZN(n15745) );
  NAND2_X1 U16345 ( .A1(n14895), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14878) );
  INV_X1 U16346 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n13248) );
  INV_X1 U16347 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15094) );
  INV_X1 U16348 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15885) );
  NAND2_X1 U16349 ( .A1(n15094), .A2(n15885), .ZN(n14901) );
  INV_X1 U16350 ( .A(n14901), .ZN(n13247) );
  AND2_X1 U16351 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14962) );
  NAND2_X1 U16352 ( .A1(n14962), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14977) );
  AND2_X1 U16353 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14984) );
  NAND2_X1 U16354 ( .A1(n13225), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14841) );
  INV_X1 U16355 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14436) );
  INV_X1 U16356 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14853) );
  NAND2_X1 U16357 ( .A1(n14436), .A2(n14853), .ZN(n15009) );
  INV_X1 U16358 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14964) );
  NAND2_X1 U16359 ( .A1(n15895), .A2(n14964), .ZN(n14842) );
  INV_X1 U16360 ( .A(n20570), .ZN(n20648) );
  NAND2_X1 U16361 ( .A1(n20648), .A2(n13258), .ZN(n20817) );
  AND2_X1 U16362 ( .A1(n20817), .A2(n20706), .ZN(n13252) );
  NAND2_X1 U16363 ( .A1(n20706), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13254) );
  NAND2_X1 U16364 ( .A1(n20200), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13253) );
  AND2_X1 U16365 ( .A1(n13254), .A2(n13253), .ZN(n13492) );
  INV_X1 U16366 ( .A(n13492), .ZN(n13255) );
  NOR2_X1 U16367 ( .A1(n13256), .A2(n14627), .ZN(n13257) );
  XNOR2_X1 U16368 ( .A(n13257), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13934) );
  INV_X1 U16369 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20772) );
  NOR2_X1 U16370 ( .A1(n20102), .A2(n20772), .ZN(n14966) );
  AOI21_X1 U16371 ( .B1(n20065), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14966), .ZN(n13259) );
  OAI21_X1 U16372 ( .B1(n20076), .B2(n13934), .A(n13259), .ZN(n13260) );
  NAND3_X1 U16373 ( .A1(n20706), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16038) );
  INV_X1 U16374 ( .A(n16038), .ZN(n13261) );
  NAND2_X1 U16375 ( .A1(n14625), .A2(n20071), .ZN(n13262) );
  OAI211_X1 U16376 ( .C1(n14989), .C2(n19882), .A(n13263), .B(n13262), .ZN(
        P1_U2968) );
  INV_X1 U16377 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20811) );
  NOR3_X1 U16378 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20811), .ZN(n13265) );
  NOR4_X1 U16379 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13264) );
  NAND4_X1 U16380 ( .A1(n20117), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13265), .A4(
        n13264), .ZN(U214) );
  NOR4_X1 U16381 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13266) );
  NAND3_X1 U16382 ( .A1(P2_W_R_N_REG_SCAN_IN), .A2(P2_M_IO_N_REG_SCAN_IN), 
        .A3(n13266), .ZN(n13267) );
  NOR3_X1 U16383 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .A3(n13267), .ZN(n16395) );
  NAND3_X1 U16384 ( .A1(n16395), .A2(n19156), .A3(U214), .ZN(U212) );
  AOI21_X1 U16385 ( .B1(n16163), .B2(n13268), .A(n9903), .ZN(n16155) );
  INV_X1 U16386 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18890) );
  NAND2_X1 U16387 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n13269), .ZN(
        n13280) );
  AOI21_X1 U16388 ( .B1(n18890), .B2(n13280), .A(n13270), .ZN(n18894) );
  AOI21_X1 U16389 ( .B1(n16199), .B2(n13271), .A(n13269), .ZN(n18907) );
  AOI21_X1 U16390 ( .B1(n16219), .B2(n13272), .A(n13273), .ZN(n18915) );
  NOR2_X1 U16391 ( .A1(n14220), .A2(n13274), .ZN(n13279) );
  AOI21_X1 U16392 ( .B1(n14220), .B2(n13274), .A(n13279), .ZN(n18926) );
  AOI21_X1 U16393 ( .B1(n18964), .B2(n13275), .A(n9852), .ZN(n18956) );
  AOI21_X1 U16394 ( .B1(n13276), .B2(n13277), .A(n13278), .ZN(n13889) );
  INV_X1 U16395 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n18988) );
  AOI22_X1 U16396 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13462), .B1(n18988), 
        .B2(n19859), .ZN(n14034) );
  AOI22_X1 U16397 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14096), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19859), .ZN(n14035) );
  NOR2_X1 U16398 ( .A1(n14034), .A2(n14035), .ZN(n14036) );
  OAI21_X1 U16399 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n13277), .ZN(n14065) );
  NAND2_X1 U16400 ( .A1(n14036), .A2(n14065), .ZN(n13849) );
  NOR2_X1 U16401 ( .A1(n13889), .A2(n13849), .ZN(n18965) );
  OAI21_X1 U16402 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n13278), .A(
        n13275), .ZN(n19149) );
  NAND2_X1 U16403 ( .A1(n18965), .A2(n19149), .ZN(n18953) );
  NOR2_X1 U16404 ( .A1(n18956), .A2(n18953), .ZN(n18941) );
  OAI21_X1 U16405 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n9852), .A(
        n13274), .ZN(n18942) );
  NAND2_X1 U16406 ( .A1(n18941), .A2(n18942), .ZN(n18925) );
  NOR2_X1 U16407 ( .A1(n18926), .A2(n18925), .ZN(n13965) );
  OAI21_X1 U16408 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n13279), .A(
        n13272), .ZN(n16233) );
  NAND2_X1 U16409 ( .A1(n13965), .A2(n16233), .ZN(n18914) );
  NOR2_X1 U16410 ( .A1(n18915), .A2(n18914), .ZN(n13945) );
  OAI21_X1 U16411 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n13273), .A(
        n13271), .ZN(n16211) );
  NAND2_X1 U16412 ( .A1(n13945), .A2(n16211), .ZN(n18908) );
  NOR2_X1 U16413 ( .A1(n18907), .A2(n18908), .ZN(n14046) );
  OAI21_X1 U16414 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n13269), .A(
        n13280), .ZN(n16186) );
  NAND2_X1 U16415 ( .A1(n14046), .A2(n16186), .ZN(n18892) );
  NOR2_X1 U16416 ( .A1(n18894), .A2(n18892), .ZN(n18882) );
  OAI21_X1 U16417 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n13270), .A(
        n13268), .ZN(n18883) );
  NAND2_X1 U16418 ( .A1(n18882), .A2(n18883), .ZN(n13283) );
  NOR2_X1 U16419 ( .A1(n16155), .A2(n13283), .ZN(n18866) );
  NOR3_X4 U16420 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n16335), .A3(n15763), 
        .ZN(n18961) );
  NAND2_X1 U16421 ( .A1(n18961), .A2(n18954), .ZN(n18995) );
  AOI211_X1 U16422 ( .C1(n16155), .C2(n13283), .A(n18866), .B(n18995), .ZN(
        n13308) );
  INV_X1 U16423 ( .A(n13284), .ZN(n13285) );
  AND2_X1 U16424 ( .A1(n13353), .A2(n13387), .ZN(n13289) );
  INV_X1 U16425 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19626) );
  NAND2_X1 U16426 ( .A1(n19626), .A2(n19858), .ZN(n13298) );
  NAND2_X1 U16427 ( .A1(n16050), .A2(n13298), .ZN(n13287) );
  NAND2_X1 U16428 ( .A1(n13379), .A2(n19626), .ZN(n13301) );
  INV_X1 U16429 ( .A(n13301), .ZN(n13286) );
  AOI21_X1 U16430 ( .B1(n19169), .B2(n13287), .A(n13286), .ZN(n13288) );
  NAND2_X1 U16431 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n21095), .ZN(n19728) );
  NOR2_X1 U16432 ( .A1(n19735), .A2(n19728), .ZN(n16328) );
  INV_X2 U16433 ( .A(n18938), .ZN(n18993) );
  AOI22_X1 U16434 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18968), .B1(
        P2_REIP_REG_15__SCAN_IN), .B2(n18993), .ZN(n13290) );
  OAI211_X1 U16435 ( .C1(n14083), .C2(n18950), .A(n13290), .B(n18878), .ZN(
        n13307) );
  INV_X1 U16436 ( .A(n13298), .ZN(n13291) );
  NOR2_X1 U16437 ( .A1(n13299), .A2(n13291), .ZN(n13292) );
  AND2_X1 U16438 ( .A1(n19854), .A2(n13292), .ZN(n16048) );
  INV_X1 U16439 ( .A(n16155), .ZN(n13294) );
  NAND2_X1 U16440 ( .A1(n18961), .A2(n18966), .ZN(n18989) );
  OAI22_X1 U16441 ( .A1(n13295), .A2(n18982), .B1(n13294), .B2(n18989), .ZN(
        n13306) );
  NOR2_X1 U16442 ( .A1(n13296), .A2(n9905), .ZN(n13297) );
  NOR2_X1 U16443 ( .A1(n13297), .A2(n14156), .ZN(n16156) );
  INV_X1 U16444 ( .A(n16156), .ZN(n13304) );
  NOR2_X1 U16445 ( .A1(n13299), .A2(n13298), .ZN(n13300) );
  NOR2_X1 U16446 ( .A1(n13302), .A2(n13301), .ZN(n16332) );
  OAI21_X1 U16447 ( .B1(n13303), .B2(n9916), .A(n14132), .ZN(n15595) );
  OAI22_X1 U16448 ( .A1(n13304), .A2(n18973), .B1(n18958), .B2(n15595), .ZN(
        n13305) );
  OR4_X1 U16449 ( .A1(n13308), .A2(n13307), .A3(n13306), .A4(n13305), .ZN(
        P2_U2840) );
  AOI21_X1 U16450 ( .B1(n15419), .B2(n13309), .A(n13310), .ZN(n15422) );
  OAI21_X1 U16451 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n9903), .A(
        n13309), .ZN(n18867) );
  NAND2_X1 U16452 ( .A1(n18866), .A2(n18867), .ZN(n13311) );
  NOR2_X1 U16453 ( .A1(n15422), .A2(n13311), .ZN(n13323) );
  AOI211_X1 U16454 ( .C1(n15422), .C2(n13311), .A(n13323), .B(n18995), .ZN(
        n13320) );
  AOI22_X1 U16455 ( .A1(P2_REIP_REG_17__SCAN_IN), .A2(n18993), .B1(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n18968), .ZN(n13312) );
  OAI211_X1 U16456 ( .C1(n11081), .C2(n18950), .A(n13312), .B(n18878), .ZN(
        n13319) );
  INV_X1 U16457 ( .A(n15422), .ZN(n13313) );
  OAI22_X1 U16458 ( .A1(n13314), .A2(n18982), .B1(n13313), .B2(n18989), .ZN(
        n13318) );
  OAI21_X1 U16459 ( .B1(n14157), .B2(n13315), .A(n14232), .ZN(n15567) );
  OAI21_X1 U16460 ( .B1(n13316), .B2(n14131), .A(n15166), .ZN(n15579) );
  OAI22_X1 U16461 ( .A1(n15567), .A2(n18973), .B1(n18958), .B2(n15579), .ZN(
        n13317) );
  OR4_X1 U16462 ( .A1(n13320), .A2(n13319), .A3(n13318), .A4(n13317), .ZN(
        P2_U2838) );
  OAI21_X1 U16463 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n13321), .A(
        n11822), .ZN(n15411) );
  INV_X1 U16464 ( .A(n15411), .ZN(n18848) );
  AOI21_X1 U16465 ( .B1(n18865), .B2(n13322), .A(n13321), .ZN(n18858) );
  OAI21_X1 U16466 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n13310), .A(
        n13322), .ZN(n16154) );
  INV_X1 U16467 ( .A(n16154), .ZN(n15170) );
  NOR2_X1 U16468 ( .A1(n18966), .A2(n18856), .ZN(n18846) );
  NOR2_X1 U16469 ( .A1(n18848), .A2(n18846), .ZN(n18847) );
  NOR2_X1 U16470 ( .A1(n18966), .A2(n18847), .ZN(n13324) );
  NOR2_X1 U16471 ( .A1(n13324), .A2(n13325), .ZN(n13337) );
  INV_X1 U16472 ( .A(n18961), .ZN(n19732) );
  AOI211_X1 U16473 ( .C1(n13325), .C2(n13324), .A(n13337), .B(n19732), .ZN(
        n13333) );
  OAI22_X1 U16474 ( .A1(n19779), .A2(n18938), .B1(n15238), .B2(n18950), .ZN(
        n13332) );
  INV_X1 U16475 ( .A(n13326), .ZN(n13328) );
  OAI22_X1 U16476 ( .A1(n13328), .A2(n18982), .B1(n13327), .B2(n18990), .ZN(
        n13331) );
  OAI22_X1 U16477 ( .A1(n15239), .A2(n18973), .B1(n13329), .B2(n18958), .ZN(
        n13330) );
  OR4_X1 U16478 ( .A1(n13333), .A2(n13332), .A3(n13331), .A4(n13330), .ZN(
        P2_U2834) );
  AND2_X1 U16479 ( .A1(n13335), .A2(n13341), .ZN(n13336) );
  OR2_X1 U16480 ( .A1(n13334), .A2(n13336), .ZN(n15390) );
  INV_X1 U16481 ( .A(n15390), .ZN(n13339) );
  OAI21_X1 U16482 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n9936), .A(
        n13335), .ZN(n15401) );
  INV_X1 U16483 ( .A(n15401), .ZN(n15702) );
  NOR2_X1 U16484 ( .A1(n13337), .A2(n18966), .ZN(n15700) );
  NOR2_X1 U16485 ( .A1(n15702), .A2(n15700), .ZN(n15701) );
  NOR2_X1 U16486 ( .A1(n18966), .A2(n15701), .ZN(n13338) );
  NOR2_X1 U16487 ( .A1(n13339), .A2(n13338), .ZN(n14489) );
  AOI211_X1 U16488 ( .C1(n13339), .C2(n13338), .A(n14489), .B(n19732), .ZN(
        n13347) );
  OAI22_X1 U16489 ( .A1(n19783), .A2(n18938), .B1(n11100), .B2(n18950), .ZN(
        n13346) );
  OAI22_X1 U16490 ( .A1(n13341), .A2(n18990), .B1(n13340), .B2(n18982), .ZN(
        n13345) );
  OAI21_X1 U16491 ( .B1(n15229), .B2(n13342), .A(n15212), .ZN(n15495) );
  OAI21_X1 U16492 ( .B1(n15301), .B2(n13343), .A(n15485), .ZN(n15499) );
  OAI22_X1 U16493 ( .A1(n15495), .A2(n18973), .B1(n18958), .B2(n15499), .ZN(
        n13344) );
  OR4_X1 U16494 ( .A1(n13347), .A2(n13346), .A3(n13345), .A4(n13344), .ZN(
        P2_U2832) );
  INV_X1 U16495 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19795) );
  AND2_X2 U16496 ( .A1(n16395), .A2(n19795), .ZN(n21215) );
  INV_X2 U16497 ( .A(n21215), .ZN(U215) );
  NOR2_X1 U16498 ( .A1(n11166), .A2(n16341), .ZN(n19059) );
  NAND2_X1 U16499 ( .A1(n19059), .A2(n13353), .ZN(n18987) );
  INV_X1 U16500 ( .A(n18987), .ZN(n13348) );
  INV_X1 U16501 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n19871) );
  INV_X1 U16502 ( .A(n13358), .ZN(n13357) );
  NAND2_X1 U16503 ( .A1(n19813), .A2(n16335), .ZN(n18819) );
  OAI211_X1 U16504 ( .C1(n13348), .C2(n19871), .A(n13357), .B(n18819), .ZN(
        P2_U2814) );
  INV_X1 U16505 ( .A(n19854), .ZN(n13351) );
  INV_X1 U16506 ( .A(n18819), .ZN(n13349) );
  OAI21_X1 U16507 ( .B1(n13349), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n13351), 
        .ZN(n13350) );
  OAI21_X1 U16508 ( .B1(n13352), .B2(n13351), .A(n13350), .ZN(P2_U3612) );
  INV_X1 U16509 ( .A(n11216), .ZN(n13355) );
  INV_X1 U16510 ( .A(n13353), .ZN(n16309) );
  NOR4_X1 U16511 ( .A1(n13355), .A2(n13354), .A3(n13379), .A4(n16309), .ZN(
        n16314) );
  NOR2_X1 U16512 ( .A1(n16314), .A2(n16341), .ZN(n19851) );
  OAI21_X1 U16513 ( .B1(n19851), .B2(n10990), .A(n13356), .ZN(P2_U2819) );
  INV_X1 U16514 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13362) );
  INV_X1 U16515 ( .A(n19858), .ZN(n19731) );
  NOR2_X1 U16516 ( .A1(n13357), .A2(n19731), .ZN(n13359) );
  NAND2_X1 U16517 ( .A1(n13358), .A2(n10512), .ZN(n19062) );
  INV_X1 U16518 ( .A(n19132), .ZN(n13361) );
  AOI22_X1 U16519 ( .A1(n19156), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19158), .ZN(n13899) );
  INV_X1 U16520 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13360) );
  OAI222_X1 U16521 ( .A1(n13362), .A2(n13415), .B1(n13361), .B2(n13899), .C1(
        n13360), .C2(n19062), .ZN(P2_U2982) );
  NAND2_X1 U16522 ( .A1(n18981), .A2(n13462), .ZN(n13363) );
  AND2_X1 U16523 ( .A1(n13364), .A2(n13363), .ZN(n13482) );
  NAND2_X1 U16524 ( .A1(n13365), .A2(n13462), .ZN(n13366) );
  NAND2_X1 U16525 ( .A1(n13367), .A2(n13366), .ZN(n13478) );
  INV_X1 U16526 ( .A(n13478), .ZN(n13368) );
  NAND2_X1 U16527 ( .A1(n16228), .A2(n13368), .ZN(n13369) );
  NAND2_X1 U16528 ( .A1(n16261), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n13473) );
  NAND2_X1 U16529 ( .A1(n13369), .A2(n13473), .ZN(n13372) );
  AOI21_X1 U16530 ( .B1(n16243), .B2(n13370), .A(n18988), .ZN(n13371) );
  AOI211_X1 U16531 ( .C1(n13482), .C2(n10996), .A(n13372), .B(n13371), .ZN(
        n13373) );
  OAI21_X1 U16532 ( .B1(n15646), .B2(n19157), .A(n13373), .ZN(P2_U3014) );
  NOR2_X1 U16533 ( .A1(n13376), .A2(n19875), .ZN(n13377) );
  NAND2_X1 U16534 ( .A1(n14607), .A2(n13377), .ZN(n13456) );
  NAND2_X1 U16535 ( .A1(n20570), .A2(n20705), .ZN(n19878) );
  INV_X1 U16536 ( .A(n19878), .ZN(n13457) );
  AOI21_X1 U16537 ( .B1(n13456), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n13457), 
        .ZN(n13378) );
  NAND2_X1 U16538 ( .A1(n20011), .A2(n13378), .ZN(P1_U2801) );
  INV_X1 U16539 ( .A(n13379), .ZN(n13380) );
  OR2_X1 U16540 ( .A1(n11166), .A2(n13380), .ZN(n13384) );
  NOR2_X1 U16541 ( .A1(n16313), .A2(n16308), .ZN(n13576) );
  NOR2_X1 U16542 ( .A1(n13576), .A2(n13381), .ZN(n13382) );
  OAI211_X1 U16543 ( .C1(n13384), .C2(n19058), .A(n13383), .B(n13382), .ZN(
        n16315) );
  NOR2_X1 U16544 ( .A1(n19859), .A2(n19834), .ZN(n16329) );
  NAND2_X1 U16545 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(n16329), .ZN(n13385) );
  OAI21_X1 U16546 ( .B1(n20990), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n13385), 
        .ZN(n13386) );
  AOI21_X1 U16547 ( .B1(n16315), .B2(n13387), .A(n13386), .ZN(n15651) );
  INV_X1 U16548 ( .A(n15651), .ZN(n13391) );
  AND3_X1 U16549 ( .A1(n10451), .A2(n13389), .A3(n13388), .ZN(n16319) );
  NAND3_X1 U16550 ( .A1(n13391), .A2(n14175), .A3(n16319), .ZN(n13390) );
  OAI21_X1 U16551 ( .B1(n13391), .B2(n16316), .A(n13390), .ZN(P2_U3595) );
  INV_X1 U16552 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n19080) );
  INV_X2 U16553 ( .A(n13415), .ZN(n19134) );
  NAND2_X1 U16554 ( .A1(n19134), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13392) );
  INV_X1 U16555 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16430) );
  INV_X1 U16556 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n16454) );
  AOI22_X1 U16557 ( .A1(n19156), .A2(n16430), .B1(n16454), .B2(n19158), .ZN(
        n19006) );
  NAND2_X1 U16558 ( .A1(n19132), .A2(n19006), .ZN(n13393) );
  OAI211_X1 U16559 ( .C1(n19080), .C2(n19062), .A(n13392), .B(n13393), .ZN(
        P2_U2960) );
  INV_X1 U16560 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19115) );
  NAND2_X1 U16561 ( .A1(n19134), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13394) );
  OAI211_X1 U16562 ( .C1(n19115), .C2(n19062), .A(n13394), .B(n13393), .ZN(
        P2_U2975) );
  AOI22_X1 U16563 ( .A1(n19134), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(
        P2_EAX_REG_10__SCAN_IN), .B2(n13451), .ZN(n13396) );
  AOI22_X1 U16564 ( .A1(n19156), .A2(BUF1_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n19158), .ZN(n15277) );
  INV_X1 U16565 ( .A(n15277), .ZN(n13395) );
  NAND2_X1 U16566 ( .A1(n19132), .A2(n13395), .ZN(n13439) );
  NAND2_X1 U16567 ( .A1(n13396), .A2(n13439), .ZN(P2_U2977) );
  AOI22_X1 U16568 ( .A1(n19134), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_16__SCAN_IN), .B2(n13451), .ZN(n13398) );
  AOI22_X1 U16569 ( .A1(n19156), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n19158), .ZN(n19161) );
  INV_X1 U16570 ( .A(n19161), .ZN(n13397) );
  NAND2_X1 U16571 ( .A1(n19132), .A2(n13397), .ZN(n13424) );
  NAND2_X1 U16572 ( .A1(n13398), .A2(n13424), .ZN(P2_U2952) );
  AOI22_X1 U16573 ( .A1(n19134), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n13451), .ZN(n13400) );
  AOI22_X1 U16574 ( .A1(n19156), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n19158), .ZN(n19175) );
  INV_X1 U16575 ( .A(n19175), .ZN(n13399) );
  NAND2_X1 U16576 ( .A1(n19132), .A2(n13399), .ZN(n13426) );
  NAND2_X1 U16577 ( .A1(n13400), .A2(n13426), .ZN(P2_U2954) );
  AOI22_X1 U16578 ( .A1(n19134), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n13451), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n13402) );
  AOI22_X1 U16579 ( .A1(n19156), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19158), .ZN(n19170) );
  INV_X1 U16580 ( .A(n19170), .ZN(n13401) );
  NAND2_X1 U16581 ( .A1(n19132), .A2(n13401), .ZN(n13454) );
  NAND2_X1 U16582 ( .A1(n13402), .A2(n13454), .ZN(P2_U2953) );
  AOI22_X1 U16583 ( .A1(n19134), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_3__SCAN_IN), .B2(n13451), .ZN(n13404) );
  AOI22_X1 U16584 ( .A1(n19156), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n19158), .ZN(n19181) );
  INV_X1 U16585 ( .A(n19181), .ZN(n13403) );
  NAND2_X1 U16586 ( .A1(n19132), .A2(n13403), .ZN(n13420) );
  NAND2_X1 U16587 ( .A1(n13404), .A2(n13420), .ZN(P2_U2970) );
  AOI22_X1 U16588 ( .A1(n19134), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n13451), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n13406) );
  AOI22_X1 U16589 ( .A1(n19156), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n19158), .ZN(n19191) );
  INV_X1 U16590 ( .A(n19191), .ZN(n13405) );
  NAND2_X1 U16591 ( .A1(n19132), .A2(n13405), .ZN(n13443) );
  NAND2_X1 U16592 ( .A1(n13406), .A2(n13443), .ZN(P2_U2973) );
  AOI21_X1 U16593 ( .B1(n14096), .B2(n13408), .A(n13407), .ZN(n13470) );
  OAI21_X1 U16594 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13410), .A(
        n13409), .ZN(n13465) );
  MUX2_X1 U16595 ( .A(n19150), .B(n16243), .S(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n13412) );
  NOR2_X1 U16596 ( .A1(n18878), .A2(n19754), .ZN(n13469) );
  INV_X1 U16597 ( .A(n13469), .ZN(n13411) );
  OAI211_X1 U16598 ( .C1(n13465), .C2(n19140), .A(n13412), .B(n13411), .ZN(
        n13413) );
  AOI21_X1 U16599 ( .B1(n13470), .B2(n10996), .A(n13413), .ZN(n13414) );
  OAI21_X1 U16600 ( .B1(n10520), .B2(n19157), .A(n13414), .ZN(P2_U3013) );
  AOI22_X1 U16601 ( .A1(n19134), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_11__SCAN_IN), .B2(n13451), .ZN(n13417) );
  AOI22_X1 U16602 ( .A1(n19156), .A2(BUF1_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n19158), .ZN(n15270) );
  INV_X1 U16603 ( .A(n15270), .ZN(n13416) );
  NAND2_X1 U16604 ( .A1(n19132), .A2(n13416), .ZN(n13437) );
  NAND2_X1 U16605 ( .A1(n13417), .A2(n13437), .ZN(P2_U2978) );
  AOI22_X1 U16606 ( .A1(n19134), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n13451), 
        .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n13419) );
  AOI22_X1 U16607 ( .A1(n19156), .A2(BUF1_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n19158), .ZN(n15287) );
  INV_X1 U16608 ( .A(n15287), .ZN(n13418) );
  NAND2_X1 U16609 ( .A1(n19132), .A2(n13418), .ZN(n13445) );
  NAND2_X1 U16610 ( .A1(n13419), .A2(n13445), .ZN(P2_U2961) );
  AOI22_X1 U16611 ( .A1(n19134), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n13451), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n13421) );
  NAND2_X1 U16612 ( .A1(n13421), .A2(n13420), .ZN(P2_U2955) );
  AOI22_X1 U16613 ( .A1(n19134), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_4__SCAN_IN), .B2(n13451), .ZN(n13423) );
  AOI22_X1 U16614 ( .A1(n19156), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n19158), .ZN(n19185) );
  INV_X1 U16615 ( .A(n19185), .ZN(n13422) );
  NAND2_X1 U16616 ( .A1(n19132), .A2(n13422), .ZN(n13447) );
  NAND2_X1 U16617 ( .A1(n13423), .A2(n13447), .ZN(P2_U2971) );
  AOI22_X1 U16618 ( .A1(n19134), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_0__SCAN_IN), .B2(n13451), .ZN(n13425) );
  NAND2_X1 U16619 ( .A1(n13425), .A2(n13424), .ZN(P2_U2967) );
  AOI22_X1 U16620 ( .A1(n19134), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_2__SCAN_IN), .B2(n13451), .ZN(n13427) );
  NAND2_X1 U16621 ( .A1(n13427), .A2(n13426), .ZN(P2_U2969) );
  AOI22_X1 U16622 ( .A1(n19134), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n13451), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n13428) );
  AOI22_X1 U16623 ( .A1(n19156), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n19158), .ZN(n19188) );
  INV_X1 U16624 ( .A(n19188), .ZN(n19009) );
  NAND2_X1 U16625 ( .A1(n19132), .A2(n19009), .ZN(n13452) );
  NAND2_X1 U16626 ( .A1(n13428), .A2(n13452), .ZN(P2_U2957) );
  AOI22_X1 U16627 ( .A1(n19134), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_13__SCAN_IN), .B2(n13451), .ZN(n13430) );
  INV_X1 U16628 ( .A(n13813), .ZN(n13429) );
  NAND2_X1 U16629 ( .A1(n19132), .A2(n13429), .ZN(n13433) );
  NAND2_X1 U16630 ( .A1(n13430), .A2(n13433), .ZN(P2_U2980) );
  AOI22_X1 U16631 ( .A1(n19134), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_12__SCAN_IN), .B2(n13451), .ZN(n13432) );
  AOI22_X1 U16632 ( .A1(n19156), .A2(BUF1_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n19158), .ZN(n15262) );
  INV_X1 U16633 ( .A(n15262), .ZN(n13431) );
  NAND2_X1 U16634 ( .A1(n19132), .A2(n13431), .ZN(n13435) );
  NAND2_X1 U16635 ( .A1(n13432), .A2(n13435), .ZN(P2_U2979) );
  AOI22_X1 U16636 ( .A1(n19134), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n13451), .ZN(n13434) );
  NAND2_X1 U16637 ( .A1(n13434), .A2(n13433), .ZN(P2_U2965) );
  AOI22_X1 U16638 ( .A1(n19134), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_28__SCAN_IN), .B2(n13451), .ZN(n13436) );
  NAND2_X1 U16639 ( .A1(n13436), .A2(n13435), .ZN(P2_U2964) );
  AOI22_X1 U16640 ( .A1(n19134), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n13451), .ZN(n13438) );
  NAND2_X1 U16641 ( .A1(n13438), .A2(n13437), .ZN(P2_U2963) );
  AOI22_X1 U16642 ( .A1(n19134), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(
        P2_EAX_REG_26__SCAN_IN), .B2(n13451), .ZN(n13440) );
  NAND2_X1 U16643 ( .A1(n13440), .A2(n13439), .ZN(P2_U2962) );
  AOI22_X1 U16644 ( .A1(n19134), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n13451), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n13442) );
  AOI22_X1 U16645 ( .A1(n19156), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n19158), .ZN(n19201) );
  INV_X1 U16646 ( .A(n19201), .ZN(n13441) );
  NAND2_X1 U16647 ( .A1(n19132), .A2(n13441), .ZN(n13449) );
  NAND2_X1 U16648 ( .A1(n13442), .A2(n13449), .ZN(P2_U2959) );
  AOI22_X1 U16649 ( .A1(n19134), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n13451), .ZN(n13444) );
  NAND2_X1 U16650 ( .A1(n13444), .A2(n13443), .ZN(P2_U2958) );
  AOI22_X1 U16651 ( .A1(n19134), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_9__SCAN_IN), .B2(n13451), .ZN(n13446) );
  NAND2_X1 U16652 ( .A1(n13446), .A2(n13445), .ZN(P2_U2976) );
  AOI22_X1 U16653 ( .A1(n19134), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n13451), .ZN(n13448) );
  NAND2_X1 U16654 ( .A1(n13448), .A2(n13447), .ZN(P2_U2956) );
  AOI22_X1 U16655 ( .A1(n19134), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n13451), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n13450) );
  NAND2_X1 U16656 ( .A1(n13450), .A2(n13449), .ZN(P2_U2974) );
  AOI22_X1 U16657 ( .A1(n19134), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_5__SCAN_IN), .B2(n13451), .ZN(n13453) );
  NAND2_X1 U16658 ( .A1(n13453), .A2(n13452), .ZN(P2_U2972) );
  AOI22_X1 U16659 ( .A1(n19134), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_1__SCAN_IN), .B2(n13451), .ZN(n13455) );
  NAND2_X1 U16660 ( .A1(n13455), .A2(n13454), .ZN(P2_U2968) );
  NOR2_X1 U16661 ( .A1(n13457), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n13460)
         );
  NAND2_X1 U16662 ( .A1(n20816), .A2(n13458), .ZN(n13459) );
  OAI21_X1 U16663 ( .B1(n20816), .B2(n13460), .A(n13459), .ZN(P1_U3487) );
  AOI211_X1 U16664 ( .C1(n14096), .C2(n13462), .A(n13461), .B(n15575), .ZN(
        n13467) );
  XNOR2_X1 U16665 ( .A(n13464), .B(n13463), .ZN(n19829) );
  INV_X1 U16666 ( .A(n19829), .ZN(n19012) );
  OAI22_X1 U16667 ( .A1(n16271), .A2(n19012), .B1(n13465), .B2(n15637), .ZN(
        n13466) );
  NOR2_X1 U16668 ( .A1(n13467), .A2(n13466), .ZN(n13472) );
  NOR2_X1 U16669 ( .A1(n13483), .A2(n14096), .ZN(n13468) );
  AOI211_X1 U16670 ( .C1(n13470), .C2(n16283), .A(n13469), .B(n13468), .ZN(
        n13471) );
  OAI211_X1 U16671 ( .C1(n10520), .C2(n16272), .A(n13472), .B(n13471), .ZN(
        P2_U3045) );
  OAI21_X1 U16672 ( .B1(n16272), .B2(n15646), .A(n13473), .ZN(n13481) );
  NOR2_X1 U16673 ( .A1(n13475), .A2(n13474), .ZN(n13476) );
  NOR2_X1 U16674 ( .A1(n13477), .A2(n13476), .ZN(n19054) );
  INV_X1 U16675 ( .A(n19054), .ZN(n13479) );
  OAI22_X1 U16676 ( .A1(n16271), .A2(n13479), .B1(n15637), .B2(n13478), .ZN(
        n13480) );
  AOI211_X1 U16677 ( .C1(n16283), .C2(n13482), .A(n13481), .B(n13480), .ZN(
        n13485) );
  MUX2_X1 U16678 ( .A(n15575), .B(n13483), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n13484) );
  NAND2_X1 U16679 ( .A1(n13485), .A2(n13484), .ZN(P2_U3046) );
  OAI21_X1 U16680 ( .B1(n13487), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13486), .ZN(n13630) );
  INV_X1 U16681 ( .A(n13488), .ZN(n13489) );
  AOI21_X1 U16682 ( .B1(n13491), .B2(n13490), .A(n13489), .ZN(n14702) );
  NAND2_X1 U16683 ( .A1(n14702), .A2(n20071), .ZN(n13496) );
  NAND2_X1 U16684 ( .A1(n13492), .A2(n14940), .ZN(n13494) );
  INV_X1 U16685 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13493) );
  NOR2_X1 U16686 ( .A1(n20102), .A2(n13493), .ZN(n13618) );
  AOI21_X1 U16687 ( .B1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n13494), .A(
        n13618), .ZN(n13495) );
  OAI211_X1 U16688 ( .C1(n19882), .C2(n13630), .A(n13496), .B(n13495), .ZN(
        P1_U2999) );
  INV_X1 U16689 ( .A(n13497), .ZN(n13499) );
  INV_X1 U16690 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n13498) );
  NAND2_X1 U16691 ( .A1(n13499), .A2(n13498), .ZN(n15761) );
  OAI21_X1 U16692 ( .B1(n15760), .B2(n15761), .A(n13500), .ZN(n13503) );
  INV_X1 U16693 ( .A(n13501), .ZN(n15732) );
  NAND2_X1 U16694 ( .A1(n13375), .A2(n13538), .ZN(n15158) );
  NAND3_X1 U16695 ( .A1(n14601), .A2(n15732), .A3(n15158), .ZN(n13502) );
  AND2_X1 U16696 ( .A1(n13503), .A2(n13502), .ZN(n13508) );
  NAND2_X1 U16697 ( .A1(n13544), .A2(n13504), .ZN(n13505) );
  NAND2_X1 U16698 ( .A1(n13505), .A2(n13376), .ZN(n13596) );
  OAI211_X1 U16699 ( .C1(n13928), .C2(n12396), .A(n13506), .B(n13596), .ZN(
        n13507) );
  AOI21_X1 U16700 ( .B1(n14599), .B2(n13508), .A(n13507), .ZN(n13512) );
  OR2_X1 U16701 ( .A1(n13509), .A2(n13928), .ZN(n13511) );
  NAND2_X1 U16702 ( .A1(n14617), .A2(n13128), .ZN(n13510) );
  AND2_X1 U16703 ( .A1(n13511), .A2(n13510), .ZN(n13542) );
  NOR2_X1 U16704 ( .A1(n15156), .A2(n20139), .ZN(n13591) );
  NAND2_X1 U16705 ( .A1(n13542), .A2(n13591), .ZN(n14606) );
  OR2_X1 U16706 ( .A1(n14599), .A2(n14606), .ZN(n13559) );
  INV_X1 U16707 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19883) );
  NOR2_X1 U16708 ( .A1(n20708), .A2(n20705), .ZN(n15149) );
  NAND2_X1 U16709 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15149), .ZN(n16043) );
  OAI22_X1 U16710 ( .A1(n15712), .A2(n19875), .B1(n19883), .B2(n16043), .ZN(
        n13515) );
  AOI21_X1 U16711 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20706), .A(n13515), 
        .ZN(n20799) );
  INV_X1 U16712 ( .A(n20799), .ZN(n20797) );
  INV_X1 U16713 ( .A(n20277), .ZN(n20533) );
  NOR2_X1 U16714 ( .A1(n13513), .A2(n20533), .ZN(n13514) );
  XOR2_X1 U16715 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n13514), .Z(
        n19947) );
  INV_X1 U16716 ( .A(n13139), .ZN(n13734) );
  NAND2_X1 U16717 ( .A1(n13553), .A2(n13515), .ZN(n20801) );
  INV_X1 U16718 ( .A(n20801), .ZN(n13516) );
  NAND3_X1 U16719 ( .A1(n19947), .A2(n13734), .A3(n13516), .ZN(n13517) );
  OAI21_X1 U16720 ( .B1(n20797), .B2(n13738), .A(n13517), .ZN(P1_U3468) );
  INV_X1 U16721 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13522) );
  NAND2_X1 U16722 ( .A1(n13518), .A2(n20139), .ZN(n13613) );
  OR2_X1 U16723 ( .A1(n20013), .A2(n15158), .ZN(n13519) );
  NAND2_X1 U16724 ( .A1(n20064), .A2(n13519), .ZN(n13520) );
  INV_X1 U16725 ( .A(n15761), .ZN(n13592) );
  INV_X1 U16726 ( .A(n15149), .ZN(n16039) );
  NOR2_X1 U16727 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16039), .ZN(n20005) );
  NOR2_X4 U16728 ( .A1(n19976), .A2(n20819), .ZN(n20004) );
  AOI22_X1 U16729 ( .A1(n20819), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13521) );
  OAI21_X1 U16730 ( .B1(n13522), .B2(n13719), .A(n13521), .ZN(P1_U2912) );
  INV_X1 U16731 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13524) );
  AOI22_X1 U16732 ( .A1(n20819), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13523) );
  OAI21_X1 U16733 ( .B1(n13524), .B2(n13719), .A(n13523), .ZN(P1_U2906) );
  INV_X1 U16734 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13526) );
  AOI22_X1 U16735 ( .A1(n20819), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13525) );
  OAI21_X1 U16736 ( .B1(n13526), .B2(n13719), .A(n13525), .ZN(P1_U2907) );
  INV_X1 U16737 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13528) );
  AOI22_X1 U16738 ( .A1(n20819), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13527) );
  OAI21_X1 U16739 ( .B1(n13528), .B2(n13719), .A(n13527), .ZN(P1_U2908) );
  INV_X1 U16740 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13530) );
  AOI22_X1 U16741 ( .A1(n20819), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13529) );
  OAI21_X1 U16742 ( .B1(n13530), .B2(n13719), .A(n13529), .ZN(P1_U2909) );
  INV_X1 U16743 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13532) );
  AOI22_X1 U16744 ( .A1(n20819), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13531) );
  OAI21_X1 U16745 ( .B1(n13532), .B2(n13719), .A(n13531), .ZN(P1_U2910) );
  INV_X1 U16746 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13534) );
  AOI22_X1 U16747 ( .A1(n20819), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13533) );
  OAI21_X1 U16748 ( .B1(n13534), .B2(n13719), .A(n13533), .ZN(P1_U2911) );
  INV_X1 U16749 ( .A(n12524), .ZN(n13551) );
  INV_X1 U16750 ( .A(n13535), .ZN(n13536) );
  NAND2_X1 U16751 ( .A1(n13536), .A2(n14615), .ZN(n13543) );
  NAND2_X1 U16752 ( .A1(n12402), .A2(n12396), .ZN(n13537) );
  OAI21_X1 U16753 ( .B1(n12404), .B2(n13539), .A(n13538), .ZN(n13540) );
  AND4_X1 U16754 ( .A1(n13543), .A2(n13542), .A3(n13541), .A4(n13540), .ZN(
        n13545) );
  NAND2_X1 U16755 ( .A1(n13545), .A2(n13544), .ZN(n13626) );
  INV_X1 U16756 ( .A(n13546), .ZN(n13548) );
  NAND4_X1 U16757 ( .A1(n13139), .A2(n13548), .A3(n15732), .A4(n13547), .ZN(
        n13549) );
  OR2_X1 U16758 ( .A1(n13626), .A2(n13549), .ZN(n15160) );
  INV_X1 U16759 ( .A(n15160), .ZN(n13550) );
  OAI22_X1 U16760 ( .A1(n13551), .A2(n13550), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15156), .ZN(n15709) );
  OAI22_X1 U16761 ( .A1(n20705), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20794), .ZN(n13552) );
  AOI21_X1 U16762 ( .B1(n15709), .B2(n13553), .A(n13552), .ZN(n13556) );
  INV_X1 U16763 ( .A(n15158), .ZN(n15710) );
  AOI21_X1 U16764 ( .B1(n15710), .B2(n13553), .A(n20799), .ZN(n13555) );
  OAI22_X1 U16765 ( .A1(n13556), .A2(n20799), .B1(n13555), .B2(n13554), .ZN(
        P1_U3474) );
  OAI21_X1 U16766 ( .B1(n13558), .B2(n13557), .A(n13649), .ZN(n13983) );
  NOR2_X1 U16767 ( .A1(n13560), .A2(n13570), .ZN(n13561) );
  NAND2_X1 U16768 ( .A1(n13562), .A2(n13561), .ZN(n13563) );
  INV_X1 U16769 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13973) );
  INV_X1 U16770 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20098) );
  NAND2_X1 U16771 ( .A1(n14437), .A2(n20098), .ZN(n13566) );
  OAI211_X1 U16772 ( .C1(n13570), .C2(P1_EBX_REG_1__SCAN_IN), .A(n13566), .B(
        n14404), .ZN(n13567) );
  INV_X1 U16773 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n14698) );
  NAND2_X1 U16774 ( .A1(n14404), .A2(n14698), .ZN(n13569) );
  NAND2_X1 U16775 ( .A1(n14437), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n13568) );
  XNOR2_X1 U16776 ( .A(n13652), .B(n14441), .ZN(n13974) );
  INV_X1 U16777 ( .A(n13974), .ZN(n15140) );
  AOI22_X1 U16778 ( .A1(n14767), .A2(n15140), .B1(n14765), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13571) );
  OAI21_X1 U16779 ( .B1(n13983), .B2(n14773), .A(n13571), .ZN(P1_U2871) );
  OR2_X1 U16780 ( .A1(n13573), .A2(n13572), .ZN(n13574) );
  INV_X1 U16781 ( .A(n13576), .ZN(n13577) );
  AOI21_X4 U16782 ( .B1(n13577), .B2(n11207), .A(n16341), .ZN(n15201) );
  NAND2_X1 U16783 ( .A1(n15201), .A2(n19199), .ZN(n15261) );
  NOR2_X1 U16784 ( .A1(n10520), .A2(n15259), .ZN(n13578) );
  AOI21_X1 U16785 ( .B1(P2_EBX_REG_1__SCAN_IN), .B2(n15259), .A(n13578), .ZN(
        n13579) );
  OAI21_X1 U16786 ( .B1(n19824), .B2(n15261), .A(n13579), .ZN(P2_U2886) );
  NOR2_X1 U16787 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13581) );
  OAI21_X1 U16788 ( .B1(n11220), .B2(n13581), .A(n13580), .ZN(n13582) );
  MUX2_X1 U16789 ( .A(n13584), .B(n15646), .S(n15201), .Z(n13585) );
  OAI21_X1 U16790 ( .B1(n19837), .B2(n15261), .A(n13585), .ZN(P2_U2887) );
  INV_X1 U16791 ( .A(n13587), .ZN(n13588) );
  INV_X1 U16792 ( .A(n19296), .ZN(n19817) );
  OAI21_X1 U16793 ( .B1(n19817), .B2(n15261), .A(n13590), .ZN(P2_U2885) );
  INV_X1 U16794 ( .A(n13591), .ZN(n13597) );
  OAI211_X1 U16795 ( .C1(n20139), .C2(n13592), .A(n20818), .B(n12396), .ZN(
        n13593) );
  INV_X1 U16796 ( .A(n13593), .ZN(n13594) );
  NAND2_X1 U16797 ( .A1(n14607), .A2(n13594), .ZN(n13595) );
  OAI211_X1 U16798 ( .C1(n14599), .C2(n13597), .A(n13596), .B(n13595), .ZN(
        n13598) );
  NAND2_X1 U16799 ( .A1(n13598), .A2(n14611), .ZN(n13603) );
  AOI21_X1 U16800 ( .B1(n20139), .B2(n15761), .A(n15760), .ZN(n13925) );
  NAND2_X1 U16801 ( .A1(n13599), .A2(n13620), .ZN(n13600) );
  AOI21_X1 U16802 ( .B1(n13501), .B2(n13925), .A(n13600), .ZN(n13601) );
  INV_X1 U16803 ( .A(n14602), .ZN(n13608) );
  INV_X1 U16804 ( .A(n13604), .ZN(n13607) );
  INV_X1 U16805 ( .A(n13614), .ZN(n13605) );
  NAND2_X1 U16806 ( .A1(n13605), .A2(n12392), .ZN(n13606) );
  AND4_X1 U16807 ( .A1(n13608), .A2(n13607), .A3(n14601), .A4(n13606), .ZN(
        n13609) );
  INV_X1 U16808 ( .A(n13610), .ZN(n13612) );
  INV_X1 U16809 ( .A(n14617), .ZN(n14432) );
  INV_X1 U16810 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20099) );
  NAND2_X1 U16811 ( .A1(n14432), .A2(n20099), .ZN(n13611) );
  NAND2_X1 U16812 ( .A1(n13612), .A2(n13611), .ZN(n14696) );
  INV_X1 U16813 ( .A(n14696), .ZN(n13619) );
  OAI21_X1 U16814 ( .B1(n13614), .B2(n12392), .A(n13613), .ZN(n13615) );
  INV_X1 U16815 ( .A(n13615), .ZN(n13616) );
  NAND2_X1 U16816 ( .A1(n13628), .A2(n20102), .ZN(n15136) );
  AOI21_X1 U16817 ( .B1(n14958), .B2(n15136), .A(n20099), .ZN(n13617) );
  AOI211_X1 U16818 ( .C1(n13619), .C2(n20110), .A(n13618), .B(n13617), .ZN(
        n13629) );
  MUX2_X1 U16819 ( .A(n13622), .B(n13621), .S(n13620), .Z(n13624) );
  NAND2_X1 U16820 ( .A1(n13624), .A2(n13623), .ZN(n13625) );
  NOR2_X1 U16821 ( .A1(n13626), .A2(n13625), .ZN(n13627) );
  OAI21_X1 U16822 ( .B1(n20078), .B2(n15103), .A(n20099), .ZN(n15137) );
  OAI211_X1 U16823 ( .C1(n13630), .C2(n20105), .A(n13629), .B(n15137), .ZN(
        P1_U3031) );
  INV_X1 U16824 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n13981) );
  NOR2_X1 U16825 ( .A1(n20102), .A2(n13981), .ZN(n15139) );
  NOR2_X1 U16826 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13631) );
  AOI211_X1 U16827 ( .C1(n20065), .C2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n15139), .B(n13631), .ZN(n13635) );
  OR2_X1 U16828 ( .A1(n13632), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15135) );
  NAND3_X1 U16829 ( .A1(n15135), .A2(n20072), .A3(n13633), .ZN(n13634) );
  OAI211_X1 U16830 ( .C1(n13983), .C2(n20120), .A(n13635), .B(n13634), .ZN(
        P1_U2998) );
  XOR2_X1 U16831 ( .A(n13636), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n13640)
         );
  NAND2_X1 U16832 ( .A1(n13646), .A2(n13637), .ZN(n13638) );
  AND2_X1 U16833 ( .A1(n13682), .A2(n13638), .ZN(n16235) );
  INV_X1 U16834 ( .A(n16235), .ZN(n18957) );
  MUX2_X1 U16835 ( .A(n18957), .B(n18951), .S(n15259), .Z(n13639) );
  OAI21_X1 U16836 ( .B1(n13640), .B2(n15261), .A(n13639), .ZN(P2_U2882) );
  OR2_X1 U16837 ( .A1(n9927), .A2(n13641), .ZN(n13642) );
  NAND2_X1 U16838 ( .A1(n13636), .A2(n13642), .ZN(n19023) );
  NAND2_X1 U16839 ( .A1(n13644), .A2(n13643), .ZN(n13645) );
  AND2_X1 U16840 ( .A1(n13646), .A2(n13645), .ZN(n19145) );
  INV_X1 U16841 ( .A(n19145), .ZN(n18972) );
  NOR2_X1 U16842 ( .A1(n18972), .A2(n15259), .ZN(n13647) );
  AOI21_X1 U16843 ( .B1(P2_EBX_REG_4__SCAN_IN), .B2(n15259), .A(n13647), .ZN(
        n13648) );
  OAI21_X1 U16844 ( .B1(n19023), .B2(n15261), .A(n13648), .ZN(P2_U2883) );
  OAI21_X1 U16845 ( .B1(n9932), .B2(n12530), .A(n13650), .ZN(n13944) );
  INV_X1 U16846 ( .A(n13651), .ZN(n13654) );
  NOR2_X1 U16847 ( .A1(n13652), .A2(n13570), .ZN(n13653) );
  INV_X1 U16848 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13661) );
  NAND2_X1 U16849 ( .A1(n14435), .A2(n13661), .ZN(n13657) );
  NAND2_X1 U16850 ( .A1(n14437), .A2(n20113), .ZN(n13655) );
  OAI211_X1 U16851 ( .C1(n13570), .C2(P1_EBX_REG_2__SCAN_IN), .A(n13655), .B(
        n14404), .ZN(n13656) );
  NAND2_X1 U16852 ( .A1(n13657), .A2(n13656), .ZN(n13658) );
  OR2_X1 U16853 ( .A1(n13659), .A2(n13658), .ZN(n13660) );
  NAND2_X1 U16854 ( .A1(n13660), .A2(n13724), .ZN(n20097) );
  OAI22_X1 U16855 ( .A1(n20097), .A2(n14776), .B1(n13661), .B2(n14774), .ZN(
        n13662) );
  INV_X1 U16856 ( .A(n13662), .ZN(n13663) );
  OAI21_X1 U16857 ( .B1(n13944), .B2(n14773), .A(n13663), .ZN(P1_U2870) );
  INV_X1 U16858 ( .A(n14702), .ZN(n13733) );
  NAND2_X1 U16859 ( .A1(n12393), .A2(n12509), .ZN(n13664) );
  NAND2_X2 U16860 ( .A1(n14808), .A2(n13664), .ZN(n14818) );
  INV_X1 U16861 ( .A(DATAI_0_), .ZN(n13666) );
  NAND2_X1 U16862 ( .A1(n20117), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13665) );
  OAI21_X1 U16863 ( .B1(n20117), .B2(n13666), .A(n13665), .ZN(n20014) );
  INV_X1 U16864 ( .A(n20014), .ZN(n20131) );
  INV_X1 U16865 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20008) );
  OAI222_X1 U16866 ( .A1(n13733), .A2(n14818), .B1(n14305), .B2(n20131), .C1(
        n14808), .C2(n20008), .ZN(P1_U2904) );
  INV_X1 U16867 ( .A(DATAI_1_), .ZN(n13668) );
  NAND2_X1 U16868 ( .A1(n20117), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13667) );
  OAI21_X1 U16869 ( .B1(n20117), .B2(n13668), .A(n13667), .ZN(n20017) );
  INV_X1 U16870 ( .A(n20017), .ZN(n20140) );
  INV_X1 U16871 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20003) );
  OAI222_X1 U16872 ( .A1(n13983), .A2(n14818), .B1(n14305), .B2(n20140), .C1(
        n14808), .C2(n20003), .ZN(P1_U2903) );
  OAI21_X1 U16873 ( .B1(n13669), .B2(n13962), .A(n13675), .ZN(n18919) );
  INV_X1 U16874 ( .A(n19051), .ZN(n19034) );
  INV_X1 U16875 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19113) );
  OAI222_X1 U16876 ( .A1(n18919), .A2(n19021), .B1(n15287), .B2(n19057), .C1(
        n19113), .C2(n19033), .ZN(P2_U2910) );
  XNOR2_X1 U16877 ( .A(n13672), .B(n13671), .ZN(n18948) );
  INV_X1 U16878 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19119) );
  OAI222_X1 U16879 ( .A1(n18948), .A2(n19021), .B1(n19033), .B2(n19119), .C1(
        n19057), .C2(n19191), .ZN(P2_U2913) );
  OAI21_X1 U16880 ( .B1(n13674), .B2(n13673), .A(n13963), .ZN(n18932) );
  OAI222_X1 U16881 ( .A1(n18932), .A2(n19021), .B1(n19201), .B2(n19057), .C1(
        n19117), .C2(n19033), .ZN(P2_U2912) );
  AOI21_X1 U16882 ( .B1(n13676), .B2(n13675), .A(n13693), .ZN(n13948) );
  INV_X1 U16883 ( .A(n13948), .ZN(n16270) );
  INV_X1 U16884 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19111) );
  OAI222_X1 U16885 ( .A1(n16270), .A2(n19021), .B1(n15277), .B2(n19057), .C1(
        n19111), .C2(n19033), .ZN(P2_U2909) );
  INV_X1 U16886 ( .A(DATAI_2_), .ZN(n13678) );
  NAND2_X1 U16887 ( .A1(n20117), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13677) );
  OAI21_X1 U16888 ( .B1(n20117), .B2(n13678), .A(n13677), .ZN(n20020) );
  INV_X1 U16889 ( .A(n20020), .ZN(n20143) );
  INV_X1 U16890 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20001) );
  OAI222_X1 U16891 ( .A1(n13944), .A2(n14818), .B1(n14305), .B2(n20143), .C1(
        n14808), .C2(n20001), .ZN(P1_U2902) );
  NOR2_X1 U16892 ( .A1(n13636), .A2(n13679), .ZN(n13681) );
  OAI211_X1 U16893 ( .C1(n13681), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n15247), .B(n13680), .ZN(n13685) );
  AOI21_X1 U16894 ( .B1(n13683), .B2(n13682), .A(n13696), .ZN(n18944) );
  NAND2_X1 U16895 ( .A1(n18944), .A2(n15201), .ZN(n13684) );
  OAI211_X1 U16896 ( .C1(n15201), .C2(n13686), .A(n13685), .B(n13684), .ZN(
        P2_U2881) );
  NAND2_X1 U16897 ( .A1(n13689), .A2(n13688), .ZN(n13690) );
  MUX2_X1 U16898 ( .A(n13855), .B(n13691), .S(n15201), .Z(n13692) );
  OAI21_X1 U16899 ( .B1(n19449), .B2(n15261), .A(n13692), .ZN(P2_U2884) );
  OAI21_X1 U16900 ( .B1(n13694), .B2(n13693), .A(n13766), .ZN(n18901) );
  INV_X1 U16901 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19109) );
  OAI222_X1 U16902 ( .A1(n18901), .A2(n19021), .B1(n15270), .B2(n19057), .C1(
        n19109), .C2(n19033), .ZN(P2_U2908) );
  XOR2_X1 U16903 ( .A(n13680), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n13699)
         );
  NOR2_X1 U16904 ( .A1(n13696), .A2(n13695), .ZN(n13697) );
  OR2_X1 U16905 ( .A1(n13729), .A2(n13697), .ZN(n18931) );
  MUX2_X1 U16906 ( .A(n18931), .B(n11057), .S(n15259), .Z(n13698) );
  OAI21_X1 U16907 ( .B1(n13699), .B2(n15261), .A(n13698), .ZN(P2_U2880) );
  OAI21_X1 U16908 ( .B1(n13702), .B2(n13701), .A(n13700), .ZN(n20106) );
  INV_X1 U16909 ( .A(n13944), .ZN(n13706) );
  AOI22_X1 U16910 ( .A1(n20065), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n13703), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13704) );
  OAI21_X1 U16911 ( .B1(n20076), .B2(n13936), .A(n13704), .ZN(n13705) );
  AOI21_X1 U16912 ( .B1(n13706), .B2(n20071), .A(n13705), .ZN(n13707) );
  OAI21_X1 U16913 ( .B1(n19882), .B2(n20106), .A(n13707), .ZN(P1_U2997) );
  INV_X1 U16914 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n20016) );
  AOI22_X1 U16915 ( .A1(n20005), .A2(P1_UWORD_REG_0__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13708) );
  OAI21_X1 U16916 ( .B1(n20016), .B2(n13719), .A(n13708), .ZN(P1_U2920) );
  INV_X1 U16917 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n20019) );
  AOI22_X1 U16918 ( .A1(n20005), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13709) );
  OAI21_X1 U16919 ( .B1(n20019), .B2(n13719), .A(n13709), .ZN(P1_U2919) );
  AOI22_X1 U16920 ( .A1(n20819), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13710) );
  OAI21_X1 U16921 ( .B1(n14798), .B2(n13719), .A(n13710), .ZN(P1_U2913) );
  INV_X1 U16922 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13712) );
  AOI22_X1 U16923 ( .A1(n20819), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13711) );
  OAI21_X1 U16924 ( .B1(n13712), .B2(n13719), .A(n13711), .ZN(P1_U2914) );
  AOI22_X1 U16925 ( .A1(n20819), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13713) );
  OAI21_X1 U16926 ( .B1(n14809), .B2(n13719), .A(n13713), .ZN(P1_U2915) );
  INV_X1 U16927 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13715) );
  AOI22_X1 U16928 ( .A1(n20819), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13714) );
  OAI21_X1 U16929 ( .B1(n13715), .B2(n13719), .A(n13714), .ZN(P1_U2917) );
  INV_X1 U16930 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13717) );
  AOI22_X1 U16931 ( .A1(n20819), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13716) );
  OAI21_X1 U16932 ( .B1(n13717), .B2(n13719), .A(n13716), .ZN(P1_U2916) );
  INV_X1 U16933 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n20023) );
  AOI22_X1 U16934 ( .A1(n20819), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13718) );
  OAI21_X1 U16935 ( .B1(n20023), .B2(n13719), .A(n13718), .ZN(P1_U2918) );
  OAI21_X1 U16936 ( .B1(n13721), .B2(n13722), .A(n13720), .ZN(n19968) );
  MUX2_X1 U16937 ( .A(n14431), .B(n14404), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n13723) );
  OAI21_X1 U16938 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14617), .A(
        n13723), .ZN(n13725) );
  AOI21_X1 U16939 ( .B1(n13725), .B2(n13724), .A(n13839), .ZN(n20086) );
  AOI22_X1 U16940 ( .A1(n14767), .A2(n20086), .B1(n14765), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n13726) );
  OAI21_X1 U16941 ( .B1(n19968), .B2(n14773), .A(n13726), .ZN(P1_U2869) );
  XNOR2_X1 U16942 ( .A(n13727), .B(n13815), .ZN(n13732) );
  NOR2_X1 U16943 ( .A1(n13729), .A2(n13728), .ZN(n13730) );
  OR2_X1 U16944 ( .A1(n13818), .A2(n13730), .ZN(n16220) );
  MUX2_X1 U16945 ( .A(n16220), .B(n11060), .S(n15259), .Z(n13731) );
  OAI21_X1 U16946 ( .B1(n13732), .B2(n15261), .A(n13731), .ZN(P2_U2879) );
  OAI222_X1 U16947 ( .A1(n14696), .A2(n14776), .B1(n14774), .B2(n14698), .C1(
        n14773), .C2(n13733), .ZN(P1_U2872) );
  NAND2_X1 U16948 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n19883), .ZN(n13760) );
  AOI21_X1 U16949 ( .B1(n19947), .B2(n13734), .A(n15712), .ZN(n13735) );
  NOR2_X1 U16950 ( .A1(n13735), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13736) );
  OAI21_X1 U16951 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n13759), .A(
        n13736), .ZN(n13737) );
  OAI21_X1 U16952 ( .B1(n13760), .B2(n13738), .A(n13737), .ZN(n13761) );
  INV_X1 U16953 ( .A(n13761), .ZN(n15150) );
  NOR2_X1 U16954 ( .A1(n15161), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13741) );
  NOR2_X1 U16955 ( .A1(n13741), .A2(n13740), .ZN(n13742) );
  AND2_X1 U16956 ( .A1(n13742), .A2(n12543), .ZN(n20788) );
  NAND2_X1 U16957 ( .A1(n12404), .A2(n20788), .ZN(n13750) );
  AND2_X1 U16958 ( .A1(n14601), .A2(n14606), .ZN(n13756) );
  INV_X1 U16959 ( .A(n13756), .ZN(n13748) );
  MUX2_X1 U16960 ( .A(n13740), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15161), .Z(n13744) );
  NOR2_X1 U16961 ( .A1(n13744), .A2(n13743), .ZN(n13747) );
  XNOR2_X1 U16962 ( .A(n13745), .B(n12532), .ZN(n13746) );
  AOI22_X1 U16963 ( .A1(n13748), .A2(n13747), .B1(n15710), .B2(n13746), .ZN(
        n13749) );
  OAI21_X1 U16964 ( .B1(n15160), .B2(n13750), .A(n13749), .ZN(n13751) );
  AOI21_X1 U16965 ( .B1(n20397), .B2(n15160), .A(n13751), .ZN(n20791) );
  MUX2_X1 U16966 ( .A(n12532), .B(n20791), .S(n13759), .Z(n15722) );
  OAI22_X1 U16967 ( .A1(n15722), .A2(P1_STATE2_REG_1__SCAN_IN), .B1(n13760), 
        .B2(n12532), .ZN(n15146) );
  INV_X1 U16968 ( .A(n20534), .ZN(n20128) );
  XNOR2_X1 U16969 ( .A(n15161), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n20793) );
  NOR3_X1 U16970 ( .A1(n15160), .A2(n13753), .A3(n20793), .ZN(n13758) );
  INV_X1 U16971 ( .A(n20793), .ZN(n13755) );
  XNOR2_X1 U16972 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13754) );
  OAI22_X1 U16973 ( .A1(n13756), .A2(n13755), .B1(n15158), .B2(n13754), .ZN(
        n13757) );
  AOI211_X1 U16974 ( .C1(n20128), .C2(n15160), .A(n13758), .B(n13757), .ZN(
        n20802) );
  MUX2_X1 U16975 ( .A(n10190), .B(n20802), .S(n13759), .Z(n15718) );
  OAI22_X1 U16976 ( .A1(n15718), .A2(P1_STATE2_REG_1__SCAN_IN), .B1(n13760), 
        .B2(n10190), .ZN(n15147) );
  AOI21_X1 U16977 ( .B1(n15146), .B2(n15147), .A(n13761), .ZN(n15728) );
  AOI21_X1 U16978 ( .B1(n12266), .B2(n15150), .A(n15728), .ZN(n13762) );
  NOR2_X1 U16979 ( .A1(n13762), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(n13763) );
  OAI21_X1 U16980 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(
        P1_STATE2_REG_1__SCAN_IN), .A(n20706), .ZN(n20813) );
  INV_X1 U16981 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20537) );
  NAND2_X1 U16982 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20537), .ZN(n15151) );
  NAND2_X1 U16983 ( .A1(n20115), .A2(n15151), .ZN(n14524) );
  NAND2_X1 U16984 ( .A1(n20115), .A2(n20570), .ZN(n13770) );
  NAND2_X1 U16985 ( .A1(n20197), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20502) );
  XNOR2_X1 U16986 ( .A(n20121), .B(n20502), .ZN(n13765) );
  OAI222_X1 U16987 ( .A1(n14524), .A2(n20534), .B1(n20115), .B2(n20398), .C1(
        n13770), .C2(n13765), .ZN(P1_U3476) );
  AOI21_X1 U16988 ( .B1(n13767), .B2(n13766), .A(n13811), .ZN(n14048) );
  INV_X1 U16989 ( .A(n14048), .ZN(n16247) );
  INV_X1 U16990 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19107) );
  OAI222_X1 U16991 ( .A1(n16247), .A2(n19021), .B1(n15262), .B2(n19057), .C1(
        n19107), .C2(n19033), .ZN(P2_U2907) );
  NAND2_X1 U16992 ( .A1(n20119), .A2(DATAI_3_), .ZN(n13769) );
  NAND2_X1 U16993 ( .A1(n20117), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13768) );
  AND2_X1 U16994 ( .A1(n13769), .A2(n13768), .ZN(n20147) );
  INV_X1 U16995 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n19999) );
  OAI222_X1 U16996 ( .A1(n19968), .A2(n14818), .B1(n14305), .B2(n20147), .C1(
        n14808), .C2(n19999), .ZN(P1_U2901) );
  INV_X1 U16997 ( .A(n20397), .ZN(n13780) );
  INV_X1 U16998 ( .A(n13770), .ZN(n14520) );
  INV_X1 U16999 ( .A(n20121), .ZN(n13771) );
  OR2_X1 U17000 ( .A1(n20197), .A2(n20200), .ZN(n20425) );
  INV_X1 U17001 ( .A(n20425), .ZN(n13773) );
  NAND2_X1 U17002 ( .A1(n20637), .A2(n13773), .ZN(n20567) );
  INV_X1 U17003 ( .A(n13774), .ZN(n13775) );
  INV_X1 U17004 ( .A(n20502), .ZN(n20636) );
  NAND2_X1 U17005 ( .A1(n20374), .A2(n20636), .ZN(n20371) );
  OR2_X1 U17006 ( .A1(n20122), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13777) );
  NAND4_X1 U17007 ( .A1(n20503), .A2(n20567), .A3(n20371), .A4(n13777), .ZN(
        n13778) );
  INV_X1 U17008 ( .A(n20115), .ZN(n14521) );
  AOI22_X1 U17009 ( .A1(n14520), .A2(n13778), .B1(n14521), .B2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n13779) );
  OAI21_X1 U17010 ( .B1(n13780), .B2(n14524), .A(n13779), .ZN(P1_U3475) );
  INV_X1 U17011 ( .A(n13781), .ZN(n13782) );
  XNOR2_X1 U17012 ( .A(n13782), .B(n13783), .ZN(n13786) );
  AOI21_X1 U17013 ( .B1(n13784), .B2(n13819), .A(n13869), .ZN(n16208) );
  INV_X1 U17014 ( .A(n16208), .ZN(n16273) );
  MUX2_X1 U17015 ( .A(n13951), .B(n16273), .S(n15201), .Z(n13785) );
  OAI21_X1 U17016 ( .B1(n13786), .B2(n15261), .A(n13785), .ZN(P2_U2877) );
  OAI21_X1 U17017 ( .B1(n13789), .B2(n13788), .A(n13787), .ZN(n13790) );
  INV_X1 U17018 ( .A(n13790), .ZN(n20088) );
  NAND2_X1 U17019 ( .A1(n20088), .A2(n20072), .ZN(n13795) );
  INV_X1 U17020 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n13791) );
  NOR2_X1 U17021 ( .A1(n20102), .A2(n13791), .ZN(n20085) );
  NOR2_X1 U17022 ( .A1(n14940), .A2(n13792), .ZN(n13793) );
  AOI211_X1 U17023 ( .C1(n15917), .C2(n19972), .A(n20085), .B(n13793), .ZN(
        n13794) );
  OAI211_X1 U17024 ( .C1(n20120), .C2(n19968), .A(n13795), .B(n13794), .ZN(
        P1_U2996) );
  INV_X1 U17025 ( .A(n19449), .ZN(n19815) );
  INV_X1 U17026 ( .A(n14089), .ZN(n13806) );
  INV_X1 U17027 ( .A(n13796), .ZN(n16312) );
  NAND2_X1 U17028 ( .A1(n16312), .A2(n16308), .ZN(n14092) );
  INV_X1 U17029 ( .A(n10539), .ZN(n13797) );
  NAND2_X1 U17030 ( .A1(n13797), .A2(n16296), .ZN(n14087) );
  INV_X1 U17031 ( .A(n14087), .ZN(n13801) );
  NAND2_X1 U17032 ( .A1(n14092), .A2(n13801), .ZN(n13799) );
  INV_X1 U17033 ( .A(n10549), .ZN(n13800) );
  NAND2_X1 U17034 ( .A1(n14166), .A2(n13800), .ZN(n13798) );
  OAI211_X1 U17035 ( .C1(n14089), .C2(n10557), .A(n13799), .B(n13798), .ZN(
        n13804) );
  INV_X1 U17036 ( .A(n14092), .ZN(n13802) );
  INV_X1 U17037 ( .A(n14166), .ZN(n15642) );
  OAI22_X1 U17038 ( .A1(n13802), .A2(n13801), .B1(n15642), .B2(n13800), .ZN(
        n13803) );
  MUX2_X1 U17039 ( .A(n13804), .B(n13803), .S(n16293), .Z(n13805) );
  AOI21_X1 U17040 ( .B1(n13807), .B2(n13806), .A(n13805), .ZN(n13808) );
  OAI21_X1 U17041 ( .B1(n13691), .B2(n15645), .A(n13808), .ZN(n16295) );
  AOI22_X1 U17042 ( .A1(n19815), .A2(n16334), .B1(n14175), .B2(n16295), .ZN(
        n13810) );
  NAND2_X1 U17043 ( .A1(n15651), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13809) );
  OAI21_X1 U17044 ( .B1(n13810), .B2(n15651), .A(n13809), .ZN(P2_U3596) );
  OAI21_X1 U17045 ( .B1(n13812), .B2(n13811), .A(n15610), .ZN(n18895) );
  INV_X1 U17046 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19105) );
  OAI222_X1 U17047 ( .A1(n18895), .A2(n19021), .B1(n13813), .B2(n19057), .C1(
        n19105), .C2(n19033), .ZN(P2_U2906) );
  AOI21_X1 U17048 ( .B1(n13727), .B2(n13815), .A(n13814), .ZN(n13816) );
  OR3_X1 U17049 ( .A1(n13782), .A2(n13816), .A3(n15261), .ZN(n13822) );
  OR2_X1 U17050 ( .A1(n13818), .A2(n13817), .ZN(n13820) );
  NAND2_X1 U17051 ( .A1(n13820), .A2(n13819), .ZN(n18920) );
  INV_X1 U17052 ( .A(n18920), .ZN(n15634) );
  NAND2_X1 U17053 ( .A1(n15634), .A2(n15201), .ZN(n13821) );
  OAI211_X1 U17054 ( .C1(n15201), .C2(n13823), .A(n13822), .B(n13821), .ZN(
        P2_U2878) );
  OR2_X1 U17055 ( .A1(n13826), .A2(n13825), .ZN(n13827) );
  AND2_X1 U17056 ( .A1(n13824), .A2(n13827), .ZN(n19939) );
  INV_X1 U17057 ( .A(n19939), .ZN(n13838) );
  INV_X1 U17058 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n13828) );
  NAND2_X1 U17059 ( .A1(n14441), .A2(n13828), .ZN(n13829) );
  OAI211_X1 U17060 ( .C1(n14615), .C2(n16035), .A(n13829), .B(n14437), .ZN(
        n13830) );
  OAI21_X1 U17061 ( .B1(n14431), .B2(P1_EBX_REG_5__SCAN_IN), .A(n13830), .ZN(
        n13834) );
  INV_X1 U17062 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13845) );
  NAND2_X1 U17063 ( .A1(n14435), .A2(n13845), .ZN(n13833) );
  NAND2_X1 U17064 ( .A1(n14411), .A2(n13570), .ZN(n14414) );
  NAND2_X1 U17065 ( .A1(n14411), .A2(P1_EBX_REG_4__SCAN_IN), .ZN(n13832) );
  NAND2_X1 U17066 ( .A1(n13570), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13831) );
  NAND4_X1 U17067 ( .A1(n13833), .A2(n14414), .A3(n13832), .A4(n13831), .ZN(
        n13840) );
  AOI21_X1 U17068 ( .B1(n13834), .B2(n13841), .A(n13993), .ZN(n19936) );
  AOI22_X1 U17069 ( .A1(n14767), .A2(n19936), .B1(n14765), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n13835) );
  OAI21_X1 U17070 ( .B1(n13838), .B2(n14773), .A(n13835), .ZN(P1_U2867) );
  NAND2_X1 U17071 ( .A1(n20119), .A2(DATAI_5_), .ZN(n13837) );
  NAND2_X1 U17072 ( .A1(n20117), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13836) );
  AND2_X1 U17073 ( .A1(n13837), .A2(n13836), .ZN(n20155) );
  INV_X1 U17074 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n19995) );
  OAI222_X1 U17075 ( .A1(n13838), .A2(n14818), .B1(n14305), .B2(n20155), .C1(
        n14808), .C2(n19995), .ZN(P1_U2899) );
  OR2_X1 U17076 ( .A1(n13840), .A2(n13839), .ZN(n13842) );
  NAND2_X1 U17077 ( .A1(n13842), .A2(n13841), .ZN(n19946) );
  INV_X1 U17078 ( .A(n13843), .ZN(n13844) );
  XNOR2_X1 U17079 ( .A(n13720), .B(n13844), .ZN(n20070) );
  INV_X1 U17080 ( .A(n20070), .ZN(n13848) );
  OAI222_X1 U17081 ( .A1(n19946), .A2(n14776), .B1(n14773), .B2(n13848), .C1(
        n14774), .C2(n13845), .ZN(P1_U2868) );
  INV_X1 U17082 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n19997) );
  NAND2_X1 U17083 ( .A1(n20119), .A2(DATAI_4_), .ZN(n13847) );
  NAND2_X1 U17084 ( .A1(n20117), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13846) );
  AND2_X1 U17085 ( .A1(n13847), .A2(n13846), .ZN(n20151) );
  OAI222_X1 U17086 ( .A1(n14808), .A2(n19997), .B1(n14305), .B2(n20151), .C1(
        n14818), .C2(n13848), .ZN(P1_U2900) );
  NAND2_X1 U17087 ( .A1(n18954), .A2(n13849), .ZN(n13850) );
  XNOR2_X1 U17088 ( .A(n13889), .B(n13850), .ZN(n13863) );
  OR2_X1 U17089 ( .A1(n13852), .A2(n13851), .ZN(n13854) );
  NAND2_X1 U17090 ( .A1(n13854), .A2(n13853), .ZN(n19035) );
  INV_X1 U17091 ( .A(n19035), .ZN(n19814) );
  OAI22_X1 U17092 ( .A1(n13887), .A2(n18938), .B1(n13855), .B2(n18950), .ZN(
        n13858) );
  OAI22_X1 U17093 ( .A1(n13276), .A2(n18990), .B1(n13856), .B2(n18982), .ZN(
        n13857) );
  AOI211_X1 U17094 ( .C1(n18979), .C2(n19814), .A(n13858), .B(n13857), .ZN(
        n13861) );
  INV_X1 U17095 ( .A(n13691), .ZN(n13859) );
  NAND2_X1 U17096 ( .A1(n13859), .A2(n18984), .ZN(n13860) );
  OAI211_X1 U17097 ( .C1(n18987), .C2(n19449), .A(n13861), .B(n13860), .ZN(
        n13862) );
  AOI21_X1 U17098 ( .B1(n13863), .B2(n18961), .A(n13862), .ZN(n13864) );
  INV_X1 U17099 ( .A(n13864), .ZN(P2_U2852) );
  OAI211_X1 U17100 ( .C1(n13868), .C2(n13867), .A(n13866), .B(n15247), .ZN(
        n13873) );
  NOR2_X1 U17101 ( .A1(n13870), .A2(n13869), .ZN(n13871) );
  NOR2_X1 U17102 ( .A1(n13871), .A2(n13894), .ZN(n18905) );
  NAND2_X1 U17103 ( .A1(n18905), .A2(n15201), .ZN(n13872) );
  OAI211_X1 U17104 ( .C1(n15201), .C2(n13874), .A(n13873), .B(n13872), .ZN(
        P2_U2876) );
  XOR2_X1 U17105 ( .A(n13824), .B(n13875), .Z(n19927) );
  INV_X1 U17106 ( .A(n19927), .ZN(n13910) );
  INV_X1 U17107 ( .A(n14435), .ZN(n13879) );
  INV_X1 U17108 ( .A(n14414), .ZN(n13876) );
  AOI21_X1 U17109 ( .B1(n14411), .B2(P1_EBX_REG_6__SCAN_IN), .A(n13876), .ZN(
        n13878) );
  NAND2_X1 U17110 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13570), .ZN(
        n13877) );
  OAI211_X1 U17111 ( .C1(P1_EBX_REG_6__SCAN_IN), .C2(n13879), .A(n13878), .B(
        n13877), .ZN(n13992) );
  XOR2_X1 U17112 ( .A(n13993), .B(n13992), .Z(n19922) );
  AOI22_X1 U17113 ( .A1(n14767), .A2(n19922), .B1(n14765), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n13880) );
  OAI21_X1 U17114 ( .B1(n13910), .B2(n14773), .A(n13880), .ZN(P1_U2866) );
  NAND2_X1 U17115 ( .A1(n13882), .A2(n13881), .ZN(n13884) );
  XNOR2_X1 U17116 ( .A(n13884), .B(n13883), .ZN(n13907) );
  XOR2_X1 U17117 ( .A(n13885), .B(n13886), .Z(n13904) );
  OAI22_X1 U17118 ( .A1(n16243), .A2(n13276), .B1(n13887), .B2(n18878), .ZN(
        n13888) );
  AOI21_X1 U17119 ( .B1(n16234), .B2(n13889), .A(n13888), .ZN(n13890) );
  OAI21_X1 U17120 ( .B1(n13691), .B2(n19157), .A(n13890), .ZN(n13891) );
  AOI21_X1 U17121 ( .B1(n13904), .B2(n16228), .A(n13891), .ZN(n13892) );
  OAI21_X1 U17122 ( .B1(n13907), .B2(n19142), .A(n13892), .ZN(P2_U3011) );
  XNOR2_X1 U17123 ( .A(n13866), .B(n13914), .ZN(n13898) );
  INV_X1 U17124 ( .A(n13893), .ZN(n13896) );
  INV_X1 U17125 ( .A(n13894), .ZN(n13895) );
  AOI21_X1 U17126 ( .B1(n13896), .B2(n13895), .A(n13912), .ZN(n16183) );
  INV_X1 U17127 ( .A(n16183), .ZN(n16248) );
  MUX2_X1 U17128 ( .A(n14049), .B(n16248), .S(n15201), .Z(n13897) );
  OAI21_X1 U17129 ( .B1(n13898), .B2(n15261), .A(n13897), .ZN(P2_U2875) );
  OAI222_X1 U17130 ( .A1(n15595), .A2(n19021), .B1(n19033), .B2(n13360), .C1(
        n13899), .C2(n19057), .ZN(P2_U2904) );
  INV_X1 U17131 ( .A(n13900), .ZN(n14571) );
  OAI21_X1 U17132 ( .B1(n14571), .B2(n15572), .A(n13901), .ZN(n14183) );
  MUX2_X1 U17133 ( .A(n14022), .B(n14183), .S(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(n13903) );
  OAI22_X1 U17134 ( .A1(n19035), .A2(n16271), .B1(n13887), .B2(n18878), .ZN(
        n13902) );
  AOI211_X1 U17135 ( .C1(n16285), .C2(n13859), .A(n13903), .B(n13902), .ZN(
        n13906) );
  NAND2_X1 U17136 ( .A1(n13904), .A2(n11843), .ZN(n13905) );
  OAI211_X1 U17137 ( .C1(n13907), .C2(n16278), .A(n13906), .B(n13905), .ZN(
        P2_U3043) );
  NAND2_X1 U17138 ( .A1(n20119), .A2(DATAI_6_), .ZN(n13909) );
  NAND2_X1 U17139 ( .A1(n20117), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13908) );
  AND2_X1 U17140 ( .A1(n13909), .A2(n13908), .ZN(n20159) );
  OAI222_X1 U17141 ( .A1(n14818), .A2(n13910), .B1(n14305), .B2(n20159), .C1(
        n14808), .C2(n12629), .ZN(P1_U2898) );
  OAI21_X1 U17142 ( .B1(n13912), .B2(n13911), .A(n13957), .ZN(n18896) );
  OAI21_X1 U17143 ( .B1(n13866), .B2(n13914), .A(n13913), .ZN(n13916) );
  NAND3_X1 U17144 ( .A1(n13916), .A2(n15247), .A3(n13915), .ZN(n13918) );
  NAND2_X1 U17145 ( .A1(n15259), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n13917) );
  OAI211_X1 U17146 ( .C1(n18896), .C2(n15259), .A(n13918), .B(n13917), .ZN(
        P2_U2874) );
  NAND3_X1 U17147 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20708), .A3(n20705), 
        .ZN(n15739) );
  AND2_X1 U17148 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20706), .ZN(n13919) );
  NAND2_X1 U17149 ( .A1(n13920), .A2(n13919), .ZN(n13921) );
  OAI21_X1 U17150 ( .B1(n15739), .B2(n20706), .A(n13921), .ZN(n13922) );
  NOR2_X1 U17151 ( .A1(n13934), .A2(n20705), .ZN(n13923) );
  NOR2_X1 U17152 ( .A1(n13929), .A2(n14609), .ZN(n13924) );
  INV_X1 U17153 ( .A(n19952), .ZN(n19969) );
  NOR2_X1 U17154 ( .A1(n13929), .A2(n20124), .ZN(n13933) );
  AND2_X1 U17155 ( .A1(n13925), .A2(n20200), .ZN(n13931) );
  AOI21_X1 U17156 ( .B1(n19945), .B2(n13981), .A(n19932), .ZN(n19975) );
  INV_X1 U17157 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20727) );
  INV_X1 U17158 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14704) );
  NOR2_X1 U17159 ( .A1(n20139), .A2(n14704), .ZN(n13930) );
  NAND2_X1 U17160 ( .A1(n20818), .A2(n20200), .ZN(n15731) );
  AND2_X1 U17161 ( .A1(n13930), .A2(n15731), .ZN(n13926) );
  OAI22_X1 U17162 ( .A1(n19975), .A2(n20727), .B1(n15859), .B2(n20097), .ZN(
        n13927) );
  INV_X1 U17163 ( .A(n13927), .ZN(n13943) );
  NOR2_X1 U17164 ( .A1(n19934), .A2(n13981), .ZN(n19963) );
  NOR2_X1 U17165 ( .A1(n13929), .A2(n13928), .ZN(n19965) );
  INV_X1 U17166 ( .A(n19965), .ZN(n13940) );
  NOR2_X1 U17167 ( .A1(n13931), .A2(n13930), .ZN(n13932) );
  AND2_X2 U17168 ( .A1(n13933), .A2(n13932), .ZN(n19961) );
  NAND2_X1 U17169 ( .A1(n19961), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n13939) );
  AND2_X1 U17170 ( .A1(n13934), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13935) );
  INV_X1 U17171 ( .A(n13936), .ZN(n13937) );
  AOI22_X1 U17172 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n19964), .B1(
        n19971), .B2(n13937), .ZN(n13938) );
  OAI211_X1 U17173 ( .C1(n13940), .C2(n20534), .A(n13939), .B(n13938), .ZN(
        n13941) );
  AOI21_X1 U17174 ( .B1(n19963), .B2(n20727), .A(n13941), .ZN(n13942) );
  OAI211_X1 U17175 ( .C1(n19969), .C2(n13944), .A(n13943), .B(n13942), .ZN(
        P1_U2838) );
  NOR2_X1 U17176 ( .A1(n18966), .A2(n13945), .ZN(n13946) );
  XNOR2_X1 U17177 ( .A(n13946), .B(n16211), .ZN(n13947) );
  AOI22_X1 U17178 ( .A1(n18979), .A2(n13948), .B1(n18961), .B2(n13947), .ZN(
        n13955) );
  OAI21_X1 U17179 ( .B1(n16273), .B2(n18973), .A(n18878), .ZN(n13953) );
  AOI22_X1 U17180 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n18968), .B1(
        n13949), .B2(n18928), .ZN(n13950) );
  OAI21_X1 U17181 ( .B1(n13951), .B2(n18950), .A(n13950), .ZN(n13952) );
  AOI211_X1 U17182 ( .C1(n18993), .C2(P2_REIP_REG_10__SCAN_IN), .A(n13953), 
        .B(n13952), .ZN(n13954) );
  NAND2_X1 U17183 ( .A1(n13955), .A2(n13954), .ZN(P2_U2845) );
  XNOR2_X1 U17184 ( .A(n13915), .B(n13956), .ZN(n13961) );
  AOI21_X1 U17185 ( .B1(n13958), .B2(n13957), .A(n9905), .ZN(n18885) );
  NOR2_X1 U17186 ( .A1(n15201), .A2(n10870), .ZN(n13959) );
  AOI21_X1 U17187 ( .B1(n18885), .B2(n15201), .A(n13959), .ZN(n13960) );
  OAI21_X1 U17188 ( .B1(n13961), .B2(n15261), .A(n13960), .ZN(P2_U2873) );
  AOI21_X1 U17189 ( .B1(n13964), .B2(n13963), .A(n13962), .ZN(n19005) );
  NOR2_X1 U17190 ( .A1(n18966), .A2(n13965), .ZN(n13966) );
  XNOR2_X1 U17191 ( .A(n13966), .B(n16233), .ZN(n13967) );
  AOI22_X1 U17192 ( .A1(n18979), .A2(n19005), .B1(n18961), .B2(n13967), .ZN(
        n13972) );
  AOI22_X1 U17193 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18968), .B1(
        P2_EBX_REG_8__SCAN_IN), .B2(n18978), .ZN(n13968) );
  OAI21_X1 U17194 ( .B1(n13969), .B2(n18982), .A(n13968), .ZN(n13970) );
  AOI211_X1 U17195 ( .C1(P2_REIP_REG_8__SCAN_IN), .C2(n18993), .A(n16261), .B(
        n13970), .ZN(n13971) );
  OAI211_X1 U17196 ( .C1(n18973), .C2(n16220), .A(n13972), .B(n13971), .ZN(
        P2_U2847) );
  INV_X1 U17197 ( .A(n19961), .ZN(n14697) );
  OAI22_X1 U17198 ( .A1(n13974), .A2(n15859), .B1(n13973), .B2(n14697), .ZN(
        n13976) );
  NOR2_X1 U17199 ( .A1(n15796), .A2(n13981), .ZN(n13975) );
  AOI211_X1 U17200 ( .C1(n19964), .C2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13976), .B(n13975), .ZN(n13979) );
  INV_X1 U17201 ( .A(n20535), .ZN(n20592) );
  NAND2_X1 U17202 ( .A1(n19965), .A2(n20592), .ZN(n13978) );
  OAI211_X1 U17203 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n19959), .A(
        n13979), .B(n13978), .ZN(n13980) );
  AOI21_X1 U17204 ( .B1(n19945), .B2(n13981), .A(n13980), .ZN(n13982) );
  OAI21_X1 U17205 ( .B1(n13983), .B2(n19969), .A(n13982), .ZN(P1_U2839) );
  INV_X1 U17206 ( .A(n13984), .ZN(n13988) );
  AOI21_X1 U17207 ( .B1(n13988), .B2(n10115), .A(n13987), .ZN(n14105) );
  INV_X1 U17208 ( .A(n14105), .ZN(n14084) );
  INV_X1 U17209 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20735) );
  INV_X1 U17210 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20732) );
  NAND4_X1 U17211 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n19933)
         );
  NOR2_X1 U17212 ( .A1(n20732), .A2(n19933), .ZN(n19921) );
  NAND2_X1 U17213 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n19921), .ZN(n19919) );
  NOR2_X1 U17214 ( .A1(n20735), .A2(n19919), .ZN(n14005) );
  NAND2_X1 U17215 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n14005), .ZN(n14258) );
  AND2_X1 U17216 ( .A1(n14258), .A2(n19945), .ZN(n14006) );
  INV_X1 U17217 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n14002) );
  INV_X1 U17218 ( .A(n14103), .ZN(n14000) );
  NAND2_X1 U17219 ( .A1(n14435), .A2(n14002), .ZN(n13991) );
  NAND2_X1 U17220 ( .A1(n14411), .A2(P1_EBX_REG_8__SCAN_IN), .ZN(n13990) );
  NAND2_X1 U17221 ( .A1(n13570), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13989) );
  NAND4_X1 U17222 ( .A1(n13991), .A2(n14414), .A3(n13990), .A4(n13989), .ZN(
        n13997) );
  NAND2_X1 U17223 ( .A1(n13993), .A2(n13992), .ZN(n14014) );
  INV_X1 U17224 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16024) );
  INV_X1 U17225 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n13994) );
  NAND2_X1 U17226 ( .A1(n14441), .A2(n13994), .ZN(n13995) );
  OAI211_X1 U17227 ( .C1(n14615), .C2(n16024), .A(n13995), .B(n14437), .ZN(
        n13996) );
  OAI21_X1 U17228 ( .B1(n14431), .B2(P1_EBX_REG_7__SCAN_IN), .A(n13996), .ZN(
        n14015) );
  NOR2_X2 U17229 ( .A1(n14014), .A2(n14015), .ZN(n14013) );
  OR2_X1 U17230 ( .A1(n13997), .A2(n14013), .ZN(n13998) );
  NAND2_X1 U17231 ( .A1(n13998), .A2(n14061), .ZN(n16015) );
  INV_X1 U17232 ( .A(n19948), .ZN(n19923) );
  OAI21_X1 U17233 ( .B1(n15859), .B2(n16015), .A(n19923), .ZN(n13999) );
  AOI21_X1 U17234 ( .B1(n19971), .B2(n14000), .A(n13999), .ZN(n14001) );
  OAI21_X1 U17235 ( .B1(n14697), .B2(n14002), .A(n14001), .ZN(n14004) );
  AOI21_X1 U17236 ( .B1(n19945), .B2(n14258), .A(n19932), .ZN(n19901) );
  INV_X1 U17237 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20737) );
  OAI22_X1 U17238 ( .A1(n19901), .A2(n20737), .B1(n12651), .B2(n19899), .ZN(
        n14003) );
  AOI211_X1 U17239 ( .C1(n14006), .C2(n14005), .A(n14004), .B(n14003), .ZN(
        n14007) );
  OAI21_X1 U17240 ( .B1(n14084), .B2(n15867), .A(n14007), .ZN(P1_U2832) );
  NAND2_X1 U17241 ( .A1(n20119), .A2(DATAI_8_), .ZN(n14009) );
  NAND2_X1 U17242 ( .A1(n20117), .A2(BUF1_REG_8__SCAN_IN), .ZN(n14008) );
  AND2_X1 U17243 ( .A1(n14009), .A2(n14008), .ZN(n20045) );
  INV_X1 U17244 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n19991) );
  OAI222_X1 U17245 ( .A1(n14084), .A2(n14818), .B1(n14305), .B2(n20045), .C1(
        n14808), .C2(n19991), .ZN(P1_U2896) );
  AND2_X1 U17246 ( .A1(n14011), .A2(n14010), .ZN(n14012) );
  NOR2_X1 U17247 ( .A1(n13985), .A2(n14012), .ZN(n19917) );
  INV_X1 U17248 ( .A(n19917), .ZN(n14033) );
  AOI21_X1 U17249 ( .B1(n14015), .B2(n14014), .A(n14013), .ZN(n19910) );
  AOI22_X1 U17250 ( .A1(n14767), .A2(n19910), .B1(n14765), .B2(
        P1_EBX_REG_7__SCAN_IN), .ZN(n14016) );
  OAI21_X1 U17251 ( .B1(n14033), .B2(n14773), .A(n14016), .ZN(P1_U2865) );
  OAI21_X1 U17252 ( .B1(n14018), .B2(n14119), .A(n14017), .ZN(n14019) );
  INV_X1 U17253 ( .A(n14019), .ZN(n19141) );
  XOR2_X1 U17254 ( .A(n14020), .B(n14021), .Z(n19139) );
  NAND2_X1 U17255 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n14022), .ZN(
        n14118) );
  AOI21_X1 U17256 ( .B1(n14023), .B2(n15604), .A(n14183), .ZN(n14117) );
  NAND2_X1 U17257 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n16261), .ZN(n14024) );
  OAI221_X1 U17258 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n14118), .C1(
        n14119), .C2(n14117), .A(n14024), .ZN(n14029) );
  NAND2_X1 U17259 ( .A1(n14025), .A2(n13853), .ZN(n14027) );
  INV_X1 U17260 ( .A(n14116), .ZN(n14026) );
  AND2_X1 U17261 ( .A1(n14027), .A2(n14026), .ZN(n19022) );
  INV_X1 U17262 ( .A(n19022), .ZN(n19015) );
  OAI22_X1 U17263 ( .A1(n18972), .A2(n16272), .B1(n16271), .B2(n19015), .ZN(
        n14028) );
  AOI211_X1 U17264 ( .C1(n19139), .C2(n16283), .A(n14029), .B(n14028), .ZN(
        n14030) );
  OAI21_X1 U17265 ( .B1(n19141), .B2(n15637), .A(n14030), .ZN(P2_U3042) );
  NAND2_X1 U17266 ( .A1(n20119), .A2(DATAI_7_), .ZN(n14032) );
  NAND2_X1 U17267 ( .A1(n20117), .A2(BUF1_REG_7__SCAN_IN), .ZN(n14031) );
  AND2_X1 U17268 ( .A1(n14032), .A2(n14031), .ZN(n20165) );
  OAI222_X1 U17269 ( .A1(n14033), .A2(n14818), .B1(n14305), .B2(n20165), .C1(
        n14808), .C2(n12639), .ZN(P1_U2897) );
  INV_X1 U17270 ( .A(n14034), .ZN(n18996) );
  INV_X1 U17271 ( .A(n14035), .ZN(n14037) );
  NOR2_X1 U17272 ( .A1(n18966), .A2(n14036), .ZN(n14066) );
  OAI21_X1 U17273 ( .B1(n18996), .B2(n14037), .A(n14066), .ZN(n14095) );
  OAI22_X1 U17274 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18989), .B1(
        n14095), .B2(n19732), .ZN(n14038) );
  INV_X1 U17275 ( .A(n14038), .ZN(n14045) );
  AOI22_X1 U17276 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18968), .B1(
        n18979), .B2(n19829), .ZN(n14040) );
  AOI22_X1 U17277 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18993), .B1(
        P2_EBX_REG_1__SCAN_IN), .B2(n18978), .ZN(n14039) );
  OAI211_X1 U17278 ( .C1(n18982), .C2(n14041), .A(n14040), .B(n14039), .ZN(
        n14042) );
  AOI21_X1 U17279 ( .B1(n14043), .B2(n18984), .A(n14042), .ZN(n14044) );
  OAI211_X1 U17280 ( .C1(n19824), .C2(n18987), .A(n14045), .B(n14044), .ZN(
        P2_U2854) );
  OR2_X1 U17281 ( .A1(n18966), .A2(n14046), .ZN(n18906) );
  XOR2_X1 U17282 ( .A(n18906), .B(n16186), .Z(n14047) );
  AOI22_X1 U17283 ( .A1(n14048), .A2(n18979), .B1(n18961), .B2(n14047), .ZN(
        n14055) );
  OAI21_X1 U17284 ( .B1(n18950), .B2(n14049), .A(n18878), .ZN(n14053) );
  AOI22_X1 U17285 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n18993), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18968), .ZN(n14050) );
  OAI21_X1 U17286 ( .B1(n14051), .B2(n18982), .A(n14050), .ZN(n14052) );
  AOI211_X1 U17287 ( .C1(n16183), .C2(n18984), .A(n14053), .B(n14052), .ZN(
        n14054) );
  NAND2_X1 U17288 ( .A1(n14055), .A2(n14054), .ZN(P2_U2843) );
  OAI21_X1 U17289 ( .B1(n13987), .B2(n14057), .A(n14056), .ZN(n19904) );
  INV_X1 U17290 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n14058) );
  NAND2_X1 U17291 ( .A1(n14441), .A2(n14058), .ZN(n14059) );
  OAI211_X1 U17292 ( .C1(n14615), .C2(n16006), .A(n14059), .B(n14437), .ZN(
        n14060) );
  OAI21_X1 U17293 ( .B1(n14431), .B2(P1_EBX_REG_9__SCAN_IN), .A(n14060), .ZN(
        n14062) );
  AOI21_X1 U17294 ( .B1(n14062), .B2(n14061), .A(n9929), .ZN(n19903) );
  AOI22_X1 U17295 ( .A1(n14767), .A2(n19903), .B1(n14765), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n14063) );
  OAI21_X1 U17296 ( .B1(n19904), .B2(n14773), .A(n14063), .ZN(P1_U2863) );
  INV_X1 U17297 ( .A(n14065), .ZN(n14591) );
  INV_X1 U17298 ( .A(n14066), .ZN(n14064) );
  AOI221_X1 U17299 ( .B1(n14591), .B2(n14066), .C1(n14065), .C2(n14064), .A(
        n19732), .ZN(n14067) );
  INV_X1 U17300 ( .A(n14067), .ZN(n14076) );
  NAND2_X1 U17301 ( .A1(n14069), .A2(n14068), .ZN(n14071) );
  NAND2_X1 U17302 ( .A1(n14071), .A2(n10229), .ZN(n19820) );
  AOI22_X1 U17303 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n18968), .B1(
        n18979), .B2(n19820), .ZN(n14073) );
  AOI22_X1 U17304 ( .A1(P2_REIP_REG_2__SCAN_IN), .A2(n18993), .B1(
        P2_EBX_REG_2__SCAN_IN), .B2(n18978), .ZN(n14072) );
  OAI211_X1 U17305 ( .C1(n18982), .C2(n14577), .A(n14073), .B(n14072), .ZN(
        n14074) );
  AOI21_X1 U17306 ( .B1(n10502), .B2(n18984), .A(n14074), .ZN(n14075) );
  OAI211_X1 U17307 ( .C1(n19817), .C2(n18987), .A(n14076), .B(n14075), .ZN(
        P2_U2853) );
  OAI211_X1 U17308 ( .C1(n14080), .C2(n14079), .A(n14078), .B(n15247), .ZN(
        n14082) );
  NAND2_X1 U17309 ( .A1(n16156), .A2(n15201), .ZN(n14081) );
  OAI211_X1 U17310 ( .C1(n15201), .C2(n14083), .A(n14082), .B(n14081), .ZN(
        P2_U2872) );
  OAI222_X1 U17311 ( .A1(n16015), .A2(n14776), .B1(n14774), .B2(n14002), .C1(
        n14773), .C2(n14084), .ZN(P1_U2864) );
  NAND2_X1 U17312 ( .A1(n20119), .A2(DATAI_9_), .ZN(n14086) );
  NAND2_X1 U17313 ( .A1(n20117), .A2(BUF1_REG_9__SCAN_IN), .ZN(n14085) );
  AND2_X1 U17314 ( .A1(n14086), .A2(n14085), .ZN(n20047) );
  INV_X1 U17315 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n19989) );
  OAI222_X1 U17316 ( .A1(n19904), .A2(n14818), .B1(n14305), .B2(n20047), .C1(
        n14808), .C2(n19989), .ZN(P1_U2895) );
  NAND2_X1 U17317 ( .A1(n12099), .A2(n14087), .ZN(n14093) );
  NOR3_X1 U17318 ( .A1(n15642), .A2(n14088), .A3(n10549), .ZN(n14091) );
  NOR2_X1 U17319 ( .A1(n14089), .A2(n14093), .ZN(n14090) );
  AOI211_X1 U17320 ( .C1(n14093), .C2(n14092), .A(n14091), .B(n14090), .ZN(
        n14094) );
  OAI21_X1 U17321 ( .B1(n14598), .B2(n15645), .A(n14094), .ZN(n16304) );
  AOI221_X1 U17322 ( .B1(n18996), .B2(n18954), .C1(n13462), .C2(n18966), .A(
        n16335), .ZN(n15650) );
  OAI21_X1 U17323 ( .B1(n18954), .B2(n14096), .A(n14095), .ZN(n14173) );
  AOI222_X1 U17324 ( .A1(n16304), .A2(n14175), .B1(n15650), .B2(n14173), .C1(
        n19296), .C2(n16334), .ZN(n14098) );
  NAND2_X1 U17325 ( .A1(n15651), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14097) );
  OAI21_X1 U17326 ( .B1(n14098), .B2(n15651), .A(n14097), .ZN(P2_U3599) );
  XOR2_X1 U17327 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n14099), .Z(
        n14100) );
  XNOR2_X1 U17328 ( .A(n14101), .B(n14100), .ZN(n16013) );
  AOI22_X1 U17329 ( .A1(n20065), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n13703), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n14102) );
  OAI21_X1 U17330 ( .B1(n20076), .B2(n14103), .A(n14102), .ZN(n14104) );
  AOI21_X1 U17331 ( .B1(n14105), .B2(n20071), .A(n14104), .ZN(n14106) );
  OAI21_X1 U17332 ( .B1(n16013), .B2(n19882), .A(n14106), .ZN(P1_U2991) );
  INV_X1 U17333 ( .A(n14108), .ZN(n14110) );
  NAND2_X1 U17334 ( .A1(n14110), .A2(n14109), .ZN(n14111) );
  XNOR2_X1 U17335 ( .A(n14107), .B(n14111), .ZN(n16236) );
  XNOR2_X1 U17336 ( .A(n14113), .B(n14112), .ZN(n16239) );
  INV_X1 U17337 ( .A(n16239), .ZN(n14126) );
  OAI21_X1 U17338 ( .B1(n14116), .B2(n14115), .A(n14114), .ZN(n19020) );
  INV_X1 U17339 ( .A(n14117), .ZN(n14122) );
  AOI221_X1 U17340 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C1(n14119), .C2(n21044), .A(
        n14118), .ZN(n14121) );
  INV_X1 U17341 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n19758) );
  NOR2_X1 U17342 ( .A1(n19758), .A2(n18878), .ZN(n14120) );
  AOI211_X1 U17343 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n14122), .A(
        n14121), .B(n14120), .ZN(n14124) );
  NAND2_X1 U17344 ( .A1(n16235), .A2(n16285), .ZN(n14123) );
  OAI211_X1 U17345 ( .C1(n19020), .C2(n16271), .A(n14124), .B(n14123), .ZN(
        n14125) );
  AOI21_X1 U17346 ( .B1(n14126), .B2(n16283), .A(n14125), .ZN(n14127) );
  OAI21_X1 U17347 ( .B1(n15637), .B2(n16236), .A(n14127), .ZN(P2_U3041) );
  AOI21_X1 U17348 ( .B1(n14129), .B2(n14078), .A(n14128), .ZN(n14130) );
  INV_X1 U17349 ( .A(n14130), .ZN(n14162) );
  AOI21_X1 U17350 ( .B1(n14133), .B2(n14132), .A(n14131), .ZN(n18873) );
  INV_X1 U17351 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n19099) );
  OAI22_X1 U17352 ( .A1(n16134), .A2(n19161), .B1(n19033), .B2(n19099), .ZN(
        n14137) );
  INV_X1 U17353 ( .A(n18999), .ZN(n15344) );
  INV_X1 U17354 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n14135) );
  INV_X1 U17355 ( .A(n18998), .ZN(n15342) );
  INV_X1 U17356 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n14134) );
  OAI22_X1 U17357 ( .A1(n15344), .A2(n14135), .B1(n15342), .B2(n14134), .ZN(
        n14136) );
  AOI211_X1 U17358 ( .C1(n19051), .C2(n18873), .A(n14137), .B(n14136), .ZN(
        n14138) );
  OAI21_X1 U17359 ( .B1(n14162), .B2(n16136), .A(n14138), .ZN(P2_U2903) );
  INV_X1 U17360 ( .A(n14139), .ZN(n14140) );
  AOI21_X1 U17361 ( .B1(n14141), .B2(n14056), .A(n14140), .ZN(n14953) );
  INV_X1 U17362 ( .A(n14953), .ZN(n14165) );
  INV_X1 U17363 ( .A(n14951), .ZN(n14153) );
  INV_X1 U17364 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20740) );
  NOR2_X1 U17365 ( .A1(n19934), .A2(n14258), .ZN(n19898) );
  NAND2_X1 U17366 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n19898), .ZN(n14143) );
  INV_X1 U17367 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20739) );
  NOR3_X1 U17368 ( .A1(n20740), .A2(n20739), .A3(n14258), .ZN(n14259) );
  INV_X1 U17369 ( .A(n14259), .ZN(n14142) );
  AOI21_X1 U17370 ( .B1(n19945), .B2(n14142), .A(n19932), .ZN(n15869) );
  AOI21_X1 U17371 ( .B1(n20740), .B2(n14143), .A(n15869), .ZN(n14152) );
  INV_X1 U17372 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14144) );
  NAND2_X1 U17373 ( .A1(n14435), .A2(n14144), .ZN(n14147) );
  NAND2_X1 U17374 ( .A1(n14411), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n14146) );
  NAND2_X1 U17375 ( .A1(n13570), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14145) );
  NAND4_X1 U17376 ( .A1(n14147), .A2(n14414), .A3(n14146), .A4(n14145), .ZN(
        n14148) );
  OR2_X1 U17377 ( .A1(n14148), .A2(n9929), .ZN(n14149) );
  NAND2_X1 U17378 ( .A1(n14149), .A2(n14275), .ZN(n15992) );
  AOI22_X1 U17379 ( .A1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n19964), .B1(
        P1_EBX_REG_10__SCAN_IN), .B2(n19961), .ZN(n14150) );
  OAI211_X1 U17380 ( .C1(n15992), .C2(n15859), .A(n14150), .B(n19923), .ZN(
        n14151) );
  AOI211_X1 U17381 ( .C1(n19971), .C2(n14153), .A(n14152), .B(n14151), .ZN(
        n14154) );
  OAI21_X1 U17382 ( .B1(n14165), .B2(n15867), .A(n14154), .ZN(P1_U2830) );
  NAND2_X1 U17383 ( .A1(n15259), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n14161) );
  INV_X1 U17384 ( .A(n14155), .ZN(n14159) );
  INV_X1 U17385 ( .A(n14156), .ZN(n14158) );
  AOI21_X1 U17386 ( .B1(n14159), .B2(n14158), .A(n14157), .ZN(n18874) );
  NAND2_X1 U17387 ( .A1(n18874), .A2(n15201), .ZN(n14160) );
  OAI211_X1 U17388 ( .C1(n14162), .C2(n15261), .A(n14161), .B(n14160), .ZN(
        P2_U2871) );
  NAND2_X1 U17389 ( .A1(n20119), .A2(DATAI_10_), .ZN(n14164) );
  NAND2_X1 U17390 ( .A1(n20117), .A2(BUF1_REG_10__SCAN_IN), .ZN(n14163) );
  AND2_X1 U17391 ( .A1(n14164), .A2(n14163), .ZN(n20049) );
  INV_X1 U17392 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n19987) );
  OAI222_X1 U17393 ( .A1(n14165), .A2(n14818), .B1(n14305), .B2(n20049), .C1(
        n14808), .C2(n19987), .ZN(P1_U2894) );
  OAI222_X1 U17394 ( .A1(n15992), .A2(n14776), .B1(n14774), .B2(n14144), .C1(
        n14773), .C2(n14165), .ZN(P1_U2862) );
  NAND2_X1 U17395 ( .A1(n14166), .A2(n10287), .ZN(n14172) );
  INV_X1 U17396 ( .A(n11189), .ZN(n14168) );
  NAND2_X1 U17397 ( .A1(n14168), .A2(n14167), .ZN(n15641) );
  OAI21_X1 U17398 ( .B1(n14170), .B2(n14169), .A(n15641), .ZN(n14171) );
  OAI211_X1 U17399 ( .C1(n10520), .C2(n15645), .A(n14172), .B(n14171), .ZN(
        n16300) );
  INV_X1 U17400 ( .A(n14173), .ZN(n14174) );
  AOI222_X1 U17401 ( .A1(n16300), .A2(n14175), .B1(n19826), .B2(n16334), .C1(
        n14174), .C2(n15650), .ZN(n14177) );
  NAND2_X1 U17402 ( .A1(n15651), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14176) );
  OAI21_X1 U17403 ( .B1(n14177), .B2(n15651), .A(n14176), .ZN(P2_U3600) );
  OAI21_X1 U17404 ( .B1(n9838), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n14179), .ZN(n14202) );
  XOR2_X1 U17405 ( .A(n14180), .B(n14181), .Z(n14200) );
  INV_X1 U17406 ( .A(n14182), .ZN(n14185) );
  INV_X1 U17407 ( .A(n14183), .ZN(n14184) );
  OAI21_X1 U17408 ( .B1(n15575), .B2(n14185), .A(n14184), .ZN(n16281) );
  NOR2_X1 U17409 ( .A1(n19760), .A2(n18878), .ZN(n14191) );
  NAND2_X1 U17410 ( .A1(n14187), .A2(n14186), .ZN(n14188) );
  NOR2_X1 U17411 ( .A1(n14189), .A2(n14188), .ZN(n14190) );
  AOI211_X1 U17412 ( .C1(n16281), .C2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n14191), .B(n14190), .ZN(n14193) );
  NAND2_X1 U17413 ( .A1(n18944), .A2(n16285), .ZN(n14192) );
  OAI211_X1 U17414 ( .C1(n18948), .C2(n16271), .A(n14193), .B(n14192), .ZN(
        n14194) );
  AOI21_X1 U17415 ( .B1(n14200), .B2(n16283), .A(n14194), .ZN(n14195) );
  OAI21_X1 U17416 ( .B1(n15637), .B2(n14202), .A(n14195), .ZN(P2_U3040) );
  INV_X1 U17417 ( .A(n18944), .ZN(n14198) );
  OAI22_X1 U17418 ( .A1(n19760), .A2(n18878), .B1(n19150), .B2(n18942), .ZN(
        n14196) );
  AOI21_X1 U17419 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n19137), .A(
        n14196), .ZN(n14197) );
  OAI21_X1 U17420 ( .B1(n14198), .B2(n19157), .A(n14197), .ZN(n14199) );
  AOI21_X1 U17421 ( .B1(n14200), .B2(n10996), .A(n14199), .ZN(n14201) );
  OAI21_X1 U17422 ( .B1(n19140), .B2(n14202), .A(n14201), .ZN(P2_U3008) );
  XNOR2_X1 U17423 ( .A(n13225), .B(n16006), .ZN(n14203) );
  XNOR2_X1 U17424 ( .A(n14204), .B(n14203), .ZN(n16002) );
  NAND2_X1 U17425 ( .A1(n16002), .A2(n20072), .ZN(n14207) );
  NOR2_X1 U17426 ( .A1(n20102), .A2(n20739), .ZN(n16000) );
  AND2_X1 U17427 ( .A1(n20065), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14205) );
  AOI211_X1 U17428 ( .C1(n19905), .C2(n15917), .A(n16000), .B(n14205), .ZN(
        n14206) );
  OAI211_X1 U17429 ( .C1(n20120), .C2(n19904), .A(n14207), .B(n14206), .ZN(
        P1_U2990) );
  OAI21_X1 U17430 ( .B1(n14128), .B2(n14209), .A(n14208), .ZN(n15349) );
  NOR2_X1 U17431 ( .A1(n15567), .A2(n15259), .ZN(n14210) );
  AOI21_X1 U17432 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n15259), .A(n14210), .ZN(
        n14211) );
  OAI21_X1 U17433 ( .B1(n15349), .B2(n15261), .A(n14211), .ZN(P2_U2870) );
  XNOR2_X1 U17434 ( .A(n14214), .B(n14213), .ZN(n14215) );
  XNOR2_X1 U17435 ( .A(n14212), .B(n14215), .ZN(n14231) );
  NOR2_X1 U17436 ( .A1(n14217), .A2(n14216), .ZN(n14219) );
  XOR2_X1 U17437 ( .A(n14219), .B(n14218), .Z(n14229) );
  OAI22_X1 U17438 ( .A1(n19762), .A2(n18878), .B1(n14220), .B2(n16243), .ZN(
        n14221) );
  AOI21_X1 U17439 ( .B1(n16234), .B2(n18926), .A(n14221), .ZN(n14222) );
  OAI21_X1 U17440 ( .B1(n18931), .B2(n19157), .A(n14222), .ZN(n14223) );
  AOI21_X1 U17441 ( .B1(n14229), .B2(n10996), .A(n14223), .ZN(n14224) );
  OAI21_X1 U17442 ( .B1(n14231), .B2(n19140), .A(n14224), .ZN(P2_U3007) );
  NOR2_X1 U17443 ( .A1(n19762), .A2(n18878), .ZN(n14225) );
  AOI221_X1 U17444 ( .B1(n16288), .B2(n14213), .C1(n16281), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n14225), .ZN(n14226) );
  INV_X1 U17445 ( .A(n14226), .ZN(n14228) );
  OAI22_X1 U17446 ( .A1(n18932), .A2(n16271), .B1(n16272), .B2(n18931), .ZN(
        n14227) );
  AOI211_X1 U17447 ( .C1(n14229), .C2(n16283), .A(n14228), .B(n14227), .ZN(
        n14230) );
  OAI21_X1 U17448 ( .B1(n15637), .B2(n14231), .A(n14230), .ZN(P2_U3039) );
  NAND2_X1 U17449 ( .A1(n14233), .A2(n14232), .ZN(n14235) );
  INV_X1 U17450 ( .A(n14234), .ZN(n15254) );
  AND2_X1 U17451 ( .A1(n14235), .A2(n15254), .ZN(n16151) );
  NOR2_X1 U17452 ( .A1(n14208), .A2(n14236), .ZN(n15252) );
  AOI21_X1 U17453 ( .B1(n14236), .B2(n14208), .A(n15252), .ZN(n15333) );
  NAND2_X1 U17454 ( .A1(n15333), .A2(n15247), .ZN(n14238) );
  NAND2_X1 U17455 ( .A1(n15259), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n14237) );
  OAI211_X1 U17456 ( .C1(n15562), .C2(n15259), .A(n14238), .B(n14237), .ZN(
        P2_U2869) );
  OAI21_X1 U17457 ( .B1(n14239), .B2(n14242), .A(n14241), .ZN(n14933) );
  INV_X1 U17458 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14243) );
  NAND2_X1 U17459 ( .A1(n14435), .A2(n14243), .ZN(n14247) );
  NAND2_X1 U17460 ( .A1(n14437), .A2(n14244), .ZN(n14245) );
  OAI211_X1 U17461 ( .C1(n13570), .C2(P1_EBX_REG_14__SCAN_IN), .A(n14245), .B(
        n14404), .ZN(n14246) );
  NAND2_X1 U17462 ( .A1(n14247), .A2(n14246), .ZN(n14254) );
  MUX2_X1 U17463 ( .A(n14431), .B(n14404), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n14248) );
  OAI21_X1 U17464 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n14617), .A(
        n14248), .ZN(n14271) );
  MUX2_X1 U17465 ( .A(n14431), .B(n14404), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n14249) );
  OAI21_X1 U17466 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n14617), .A(
        n14249), .ZN(n14276) );
  INV_X1 U17467 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n14250) );
  NAND2_X1 U17468 ( .A1(n14435), .A2(n14250), .ZN(n14253) );
  NAND2_X1 U17469 ( .A1(n14411), .A2(P1_EBX_REG_12__SCAN_IN), .ZN(n14252) );
  NAND2_X1 U17470 ( .A1(n13570), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14251) );
  NAND4_X1 U17471 ( .A1(n14253), .A2(n14414), .A3(n14252), .A4(n14251), .ZN(
        n14283) );
  OR2_X1 U17472 ( .A1(n14254), .A2(n14270), .ZN(n14255) );
  NAND2_X1 U17473 ( .A1(n14255), .A2(n14770), .ZN(n15111) );
  INV_X1 U17474 ( .A(n15111), .ZN(n14256) );
  AOI22_X1 U17475 ( .A1(n14767), .A2(n14256), .B1(n14765), .B2(
        P1_EBX_REG_14__SCAN_IN), .ZN(n14257) );
  OAI21_X1 U17476 ( .B1(n14933), .B2(n14773), .A(n14257), .ZN(P1_U2858) );
  INV_X1 U17477 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n20744) );
  NOR4_X1 U17478 ( .A1(n19934), .A2(n20740), .A3(n20739), .A4(n14258), .ZN(
        n15871) );
  NAND2_X1 U17479 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n15871), .ZN(n15862) );
  NOR2_X1 U17480 ( .A1(n19932), .A2(n19945), .ZN(n14699) );
  INV_X1 U17481 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20743) );
  NOR2_X1 U17482 ( .A1(n20744), .A2(n20743), .ZN(n14288) );
  NAND4_X1 U17483 ( .A1(n14259), .A2(n14288), .A3(P1_REIP_REG_14__SCAN_IN), 
        .A4(P1_REIP_REG_13__SCAN_IN), .ZN(n14459) );
  NOR2_X1 U17484 ( .A1(n19932), .A2(n14459), .ZN(n14685) );
  NOR2_X1 U17485 ( .A1(n14699), .A2(n14685), .ZN(n15855) );
  OAI221_X1 U17486 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(P1_REIP_REG_13__SCAN_IN), .C1(P1_REIP_REG_14__SCAN_IN), .C2(n14684), .A(n15855), .ZN(n14264) );
  INV_X1 U17487 ( .A(n14928), .ZN(n14262) );
  AOI22_X1 U17488 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19964), .B1(
        P1_EBX_REG_14__SCAN_IN), .B2(n19961), .ZN(n14260) );
  OAI211_X1 U17489 ( .C1(n15111), .C2(n15859), .A(n14260), .B(n19923), .ZN(
        n14261) );
  AOI21_X1 U17490 ( .B1(n19971), .B2(n14262), .A(n14261), .ZN(n14263) );
  OAI211_X1 U17491 ( .C1(n14933), .C2(n15867), .A(n14264), .B(n14263), .ZN(
        P1_U2826) );
  NAND2_X1 U17492 ( .A1(n14139), .A2(n14266), .ZN(n14267) );
  NAND2_X1 U17493 ( .A1(n14265), .A2(n14267), .ZN(n14273) );
  OAI21_X1 U17494 ( .B1(n14273), .B2(n14274), .A(n14265), .ZN(n14279) );
  INV_X1 U17495 ( .A(n14239), .ZN(n14268) );
  AOI21_X1 U17496 ( .B1(n14271), .B2(n14284), .A(n14270), .ZN(n15976) );
  AOI22_X1 U17497 ( .A1(n14767), .A2(n15976), .B1(n14765), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14272) );
  OAI21_X1 U17498 ( .B1(n14945), .B2(n14773), .A(n14272), .ZN(P1_U2859) );
  XOR2_X1 U17499 ( .A(n14274), .B(n14273), .Z(n15925) );
  INV_X1 U17500 ( .A(n15925), .ZN(n14296) );
  AOI21_X1 U17501 ( .B1(n14276), .B2(n14275), .A(n14282), .ZN(n15982) );
  AOI22_X1 U17502 ( .A1(n14767), .A2(n15982), .B1(n14765), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n14277) );
  OAI21_X1 U17503 ( .B1(n14296), .B2(n14773), .A(n14277), .ZN(P1_U2861) );
  NOR2_X1 U17504 ( .A1(n14279), .A2(n14278), .ZN(n14280) );
  OR2_X1 U17505 ( .A1(n14283), .A2(n14282), .ZN(n14285) );
  NAND2_X1 U17506 ( .A1(n14285), .A2(n14284), .ZN(n15858) );
  OAI222_X1 U17507 ( .A1(n15914), .A2(n14773), .B1(n14774), .B2(n14250), .C1(
        n15858), .C2(n14776), .ZN(P1_U2860) );
  NAND2_X1 U17508 ( .A1(n20119), .A2(DATAI_12_), .ZN(n14287) );
  NAND2_X1 U17509 ( .A1(n20117), .A2(BUF1_REG_12__SCAN_IN), .ZN(n14286) );
  AND2_X1 U17510 ( .A1(n14287), .A2(n14286), .ZN(n20053) );
  INV_X1 U17511 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n19983) );
  OAI222_X1 U17512 ( .A1(n15914), .A2(n14818), .B1(n14305), .B2(n20053), .C1(
        n14808), .C2(n19983), .ZN(P1_U2892) );
  INV_X1 U17513 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20746) );
  OAI21_X1 U17514 ( .B1(n14699), .B2(n14288), .A(n15869), .ZN(n15864) );
  AOI22_X1 U17515 ( .A1(P1_EBX_REG_13__SCAN_IN), .A2(n19961), .B1(n19960), 
        .B2(n15976), .ZN(n14289) );
  OAI211_X1 U17516 ( .C1(n19899), .C2(n14290), .A(n14289), .B(n19923), .ZN(
        n14291) );
  AOI221_X1 U17517 ( .B1(n14684), .B2(n20746), .C1(n15864), .C2(
        P1_REIP_REG_13__SCAN_IN), .A(n14291), .ZN(n14293) );
  NAND2_X1 U17518 ( .A1(n19971), .A2(n14942), .ZN(n14292) );
  OAI211_X1 U17519 ( .C1(n14945), .C2(n15867), .A(n14293), .B(n14292), .ZN(
        P1_U2827) );
  NAND2_X1 U17520 ( .A1(n20119), .A2(DATAI_11_), .ZN(n14295) );
  NAND2_X1 U17521 ( .A1(n20117), .A2(BUF1_REG_11__SCAN_IN), .ZN(n14294) );
  AND2_X1 U17522 ( .A1(n14295), .A2(n14294), .ZN(n20051) );
  INV_X1 U17523 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n19985) );
  OAI222_X1 U17524 ( .A1(n14296), .A2(n14818), .B1(n14305), .B2(n20051), .C1(
        n14808), .C2(n19985), .ZN(P1_U2893) );
  NAND2_X1 U17525 ( .A1(n20119), .A2(DATAI_14_), .ZN(n14298) );
  NAND2_X1 U17526 ( .A1(n20117), .A2(BUF1_REG_14__SCAN_IN), .ZN(n14297) );
  AND2_X1 U17527 ( .A1(n14298), .A2(n14297), .ZN(n20058) );
  INV_X1 U17528 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n19979) );
  OAI222_X1 U17529 ( .A1(n14933), .A2(n14818), .B1(n14305), .B2(n20058), .C1(
        n14808), .C2(n19979), .ZN(P1_U2890) );
  NAND2_X1 U17530 ( .A1(n20119), .A2(DATAI_13_), .ZN(n14300) );
  NAND2_X1 U17531 ( .A1(n20117), .A2(BUF1_REG_13__SCAN_IN), .ZN(n14299) );
  AND2_X1 U17532 ( .A1(n14300), .A2(n14299), .ZN(n20055) );
  INV_X1 U17533 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n19981) );
  OAI222_X1 U17534 ( .A1(n14945), .A2(n14818), .B1(n14305), .B2(n20055), .C1(
        n14808), .C2(n19981), .ZN(P1_U2891) );
  AOI21_X1 U17535 ( .B1(n14302), .B2(n14241), .A(n14301), .ZN(n15911) );
  INV_X1 U17536 ( .A(n15911), .ZN(n14772) );
  NAND2_X1 U17537 ( .A1(n20119), .A2(DATAI_15_), .ZN(n14304) );
  NAND2_X1 U17538 ( .A1(n20117), .A2(BUF1_REG_15__SCAN_IN), .ZN(n14303) );
  AND2_X1 U17539 ( .A1(n14304), .A2(n14303), .ZN(n20061) );
  INV_X1 U17540 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n20063) );
  OAI222_X1 U17541 ( .A1(n14772), .A2(n14818), .B1(n14305), .B2(n20061), .C1(
        n14808), .C2(n20063), .ZN(P1_U2889) );
  OAI21_X1 U17542 ( .B1(n14306), .B2(n18769), .A(n15680), .ZN(n15678) );
  OR2_X1 U17543 ( .A1(n15678), .A2(n17143), .ZN(n18147) );
  NOR2_X1 U17544 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18147), .ZN(n14307) );
  NAND3_X1 U17545 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18746)
         );
  OAI21_X1 U17546 ( .B1(n14307), .B2(n18746), .A(n18441), .ZN(n18153) );
  INV_X1 U17547 ( .A(n18153), .ZN(n14308) );
  INV_X1 U17548 ( .A(n17715), .ZN(n17776) );
  NOR2_X1 U17549 ( .A1(n17776), .A2(n18801), .ZN(n15667) );
  AOI21_X1 U17550 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n15667), .ZN(n15668) );
  NOR2_X1 U17551 ( .A1(n14308), .A2(n15668), .ZN(n14310) );
  NOR2_X1 U17552 ( .A1(n18748), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18192) );
  OR2_X1 U17553 ( .A1(n18192), .A2(n14308), .ZN(n15666) );
  OR2_X1 U17554 ( .A1(n18211), .A2(n15666), .ZN(n14309) );
  MUX2_X1 U17555 ( .A(n14310), .B(n14309), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  AND2_X1 U17556 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n16931) );
  NAND2_X1 U17557 ( .A1(n18188), .A2(n17190), .ZN(n17192) );
  INV_X1 U17558 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16592) );
  INV_X1 U17559 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16614) );
  INV_X1 U17560 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16985) );
  INV_X1 U17561 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17024) );
  INV_X1 U17562 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16675) );
  INV_X1 U17563 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17053) );
  INV_X1 U17564 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n16714) );
  INV_X1 U17565 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16733) );
  INV_X1 U17566 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16759) );
  INV_X1 U17567 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16775) );
  INV_X1 U17568 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n16806) );
  INV_X1 U17569 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17167) );
  NAND2_X1 U17570 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16997), .ZN(n16986) );
  NAND2_X1 U17571 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16952), .ZN(n16944) );
  NAND2_X1 U17572 ( .A1(n17184), .A2(n16944), .ZN(n16942) );
  OAI21_X1 U17573 ( .B1(n16931), .B2(n17192), .A(n16942), .ZN(n16936) );
  AOI22_X1 U17574 ( .A1(n9834), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17107), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14319) );
  AOI22_X1 U17575 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9831), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14318) );
  AOI22_X1 U17576 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9832), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14317) );
  AOI22_X1 U17577 ( .A1(n17094), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14316) );
  NAND4_X1 U17578 ( .A1(n14319), .A2(n14318), .A3(n14317), .A4(n14316), .ZN(
        n14325) );
  AOI22_X1 U17579 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15657), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14323) );
  AOI22_X1 U17580 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14322) );
  AOI22_X1 U17581 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11696), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14321) );
  AOI22_X1 U17582 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14320) );
  NAND4_X1 U17583 ( .A1(n14323), .A2(n14322), .A3(n14321), .A4(n14320), .ZN(
        n14324) );
  NOR2_X1 U17584 ( .A1(n14325), .A2(n14324), .ZN(n16940) );
  AOI22_X1 U17585 ( .A1(n17094), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14329) );
  AOI22_X1 U17586 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14328) );
  AOI22_X1 U17587 ( .A1(n9834), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17107), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14327) );
  AOI22_X1 U17588 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9832), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14326) );
  NAND4_X1 U17589 ( .A1(n14329), .A2(n14328), .A3(n14327), .A4(n14326), .ZN(
        n14335) );
  AOI22_X1 U17590 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n15657), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14333) );
  AOI22_X1 U17591 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9831), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14332) );
  AOI22_X1 U17592 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11696), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14331) );
  AOI22_X1 U17593 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14330) );
  NAND4_X1 U17594 ( .A1(n14333), .A2(n14332), .A3(n14331), .A4(n14330), .ZN(
        n14334) );
  NOR2_X1 U17595 ( .A1(n14335), .A2(n14334), .ZN(n16950) );
  AOI22_X1 U17596 ( .A1(n17139), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14339) );
  AOI22_X1 U17597 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17137), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14338) );
  AOI22_X1 U17598 ( .A1(n9831), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14337) );
  AOI22_X1 U17599 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9834), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14336) );
  NAND4_X1 U17600 ( .A1(n14339), .A2(n14338), .A3(n14337), .A4(n14336), .ZN(
        n14345) );
  AOI22_X1 U17601 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n15657), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14343) );
  AOI22_X1 U17602 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17107), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14342) );
  AOI22_X1 U17603 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14341) );
  AOI22_X1 U17604 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14340) );
  NAND4_X1 U17605 ( .A1(n14343), .A2(n14342), .A3(n14341), .A4(n14340), .ZN(
        n14344) );
  NOR2_X1 U17606 ( .A1(n14345), .A2(n14344), .ZN(n16958) );
  AOI22_X1 U17607 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17144), .B1(
        n17128), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14349) );
  AOI22_X1 U17608 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n9832), .B1(
        n17153), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14348) );
  AOI22_X1 U17609 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n17094), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n17123), .ZN(n14347) );
  AOI22_X1 U17610 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__7__SCAN_IN), .B2(n9831), .ZN(n14346) );
  NAND4_X1 U17611 ( .A1(n14349), .A2(n14348), .A3(n14347), .A4(n14346), .ZN(
        n14355) );
  AOI22_X1 U17612 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n15657), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14353) );
  AOI22_X1 U17613 ( .A1(n17054), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n17108), .ZN(n14352) );
  AOI22_X1 U17614 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n9834), .B1(
        P3_INSTQUEUE_REG_5__7__SCAN_IN), .B2(n9824), .ZN(n14351) );
  AOI22_X1 U17615 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n17145), .B1(
        n17146), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14350) );
  NAND4_X1 U17616 ( .A1(n14353), .A2(n14352), .A3(n14351), .A4(n14350), .ZN(
        n14354) );
  NOR2_X1 U17617 ( .A1(n14355), .A2(n14354), .ZN(n16957) );
  NOR2_X1 U17618 ( .A1(n16958), .A2(n16957), .ZN(n16955) );
  AOI22_X1 U17619 ( .A1(n9824), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14367) );
  AOI22_X1 U17620 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17107), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14366) );
  AOI22_X1 U17621 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14356) );
  INV_X1 U17622 ( .A(n14356), .ZN(n14357) );
  AOI21_X1 U17623 ( .B1(n17094), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A(
        n14357), .ZN(n14358) );
  INV_X1 U17624 ( .A(n14358), .ZN(n14364) );
  AOI22_X1 U17625 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n15657), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14362) );
  AOI22_X1 U17626 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9831), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14361) );
  AOI22_X1 U17627 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9834), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14360) );
  AOI22_X1 U17628 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14359) );
  NAND4_X1 U17629 ( .A1(n14362), .A2(n14361), .A3(n14360), .A4(n14359), .ZN(
        n14363) );
  AOI211_X1 U17630 ( .C1(n17138), .C2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A(
        n14364), .B(n14363), .ZN(n14365) );
  NAND3_X1 U17631 ( .A1(n14367), .A2(n14366), .A3(n14365), .ZN(n16954) );
  NAND2_X1 U17632 ( .A1(n16955), .A2(n16954), .ZN(n16953) );
  NOR2_X1 U17633 ( .A1(n16950), .A2(n16953), .ZN(n16947) );
  AOI22_X1 U17634 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11696), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14377) );
  AOI22_X1 U17635 ( .A1(n9831), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14376) );
  AOI22_X1 U17636 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17107), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14368) );
  OAI21_X1 U17637 ( .B1(n9850), .B2(n17179), .A(n14368), .ZN(n14374) );
  AOI22_X1 U17638 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n15657), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14372) );
  AOI22_X1 U17639 ( .A1(n17128), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9834), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14371) );
  AOI22_X1 U17640 ( .A1(n17094), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14370) );
  AOI22_X1 U17641 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14369) );
  NAND4_X1 U17642 ( .A1(n14372), .A2(n14371), .A3(n14370), .A4(n14369), .ZN(
        n14373) );
  AOI211_X1 U17643 ( .C1(n17138), .C2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n14374), .B(n14373), .ZN(n14375) );
  NAND3_X1 U17644 ( .A1(n14377), .A2(n14376), .A3(n14375), .ZN(n16946) );
  NAND2_X1 U17645 ( .A1(n16947), .A2(n16946), .ZN(n16945) );
  NOR2_X1 U17646 ( .A1(n16940), .A2(n16945), .ZN(n16939) );
  AOI22_X1 U17647 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17153), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14381) );
  AOI22_X1 U17648 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17107), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14380) );
  AOI22_X1 U17649 ( .A1(n17094), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14379) );
  AOI22_X1 U17650 ( .A1(n9831), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11696), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14378) );
  NAND4_X1 U17651 ( .A1(n14381), .A2(n14380), .A3(n14379), .A4(n14378), .ZN(
        n14387) );
  AOI22_X1 U17652 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n15657), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14385) );
  AOI22_X1 U17653 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17140), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14384) );
  AOI22_X1 U17654 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9834), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14383) );
  AOI22_X1 U17655 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14382) );
  NAND4_X1 U17656 ( .A1(n14385), .A2(n14384), .A3(n14383), .A4(n14382), .ZN(
        n14386) );
  NOR2_X1 U17657 ( .A1(n14387), .A2(n14386), .ZN(n16932) );
  XNOR2_X1 U17658 ( .A(n16939), .B(n16932), .ZN(n17213) );
  AOI22_X1 U17659 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16936), .B1(n17188), 
        .B2(n17213), .ZN(n14390) );
  INV_X1 U17660 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n14388) );
  INV_X1 U17661 ( .A(n16944), .ZN(n16949) );
  NAND3_X1 U17662 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n14388), .A3(n16949), 
        .ZN(n14389) );
  NAND2_X1 U17663 ( .A1(n14390), .A2(n14389), .ZN(P3_U2675) );
  XNOR2_X1 U17664 ( .A(n14636), .B(n14392), .ZN(n14839) );
  INV_X1 U17665 ( .A(n14839), .ZN(n14780) );
  INV_X1 U17666 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14448) );
  MUX2_X1 U17667 ( .A(n14431), .B(n14404), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n14393) );
  OAI21_X1 U17668 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n14617), .A(
        n14393), .ZN(n14739) );
  MUX2_X1 U17669 ( .A(n14431), .B(n14404), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n14394) );
  OAI21_X1 U17670 ( .B1(n14617), .B2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n14394), .ZN(n14688) );
  MUX2_X1 U17671 ( .A(n14431), .B(n14404), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n14395) );
  OAI21_X1 U17672 ( .B1(n14617), .B2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n14395), .ZN(n14771) );
  INV_X1 U17673 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14396) );
  NAND2_X1 U17674 ( .A1(n14435), .A2(n14396), .ZN(n14399) );
  INV_X1 U17675 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15894) );
  NAND2_X1 U17676 ( .A1(n14437), .A2(n15894), .ZN(n14397) );
  OAI211_X1 U17677 ( .C1(n13570), .C2(P1_EBX_REG_16__SCAN_IN), .A(n14397), .B(
        n14404), .ZN(n14398) );
  NAND2_X1 U17678 ( .A1(n14399), .A2(n14398), .ZN(n14762) );
  INV_X1 U17679 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14400) );
  NAND2_X1 U17680 ( .A1(n14435), .A2(n14400), .ZN(n14403) );
  NAND2_X1 U17681 ( .A1(n14437), .A2(n15094), .ZN(n14401) );
  OAI211_X1 U17682 ( .C1(n13570), .C2(P1_EBX_REG_18__SCAN_IN), .A(n14401), .B(
        n14404), .ZN(n14402) );
  NAND2_X1 U17683 ( .A1(n14403), .A2(n14402), .ZN(n14753) );
  MUX2_X1 U17684 ( .A(n14431), .B(n14404), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n14405) );
  OAI21_X1 U17685 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n14617), .A(
        n14405), .ZN(n14750) );
  INV_X1 U17686 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14406) );
  NAND2_X1 U17687 ( .A1(n14435), .A2(n14406), .ZN(n14409) );
  NAND2_X1 U17688 ( .A1(n14411), .A2(P1_EBX_REG_20__SCAN_IN), .ZN(n14408) );
  NAND2_X1 U17689 ( .A1(n13570), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14407) );
  NAND4_X1 U17690 ( .A1(n14409), .A2(n14414), .A3(n14408), .A4(n14407), .ZN(
        n14741) );
  INV_X1 U17691 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14410) );
  NAND2_X1 U17692 ( .A1(n14435), .A2(n14410), .ZN(n14415) );
  NAND2_X1 U17693 ( .A1(n14411), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n14413) );
  NAND2_X1 U17694 ( .A1(n13570), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14412) );
  NAND4_X1 U17695 ( .A1(n14415), .A2(n14414), .A3(n14413), .A4(n14412), .ZN(
        n14730) );
  INV_X1 U17696 ( .A(n14731), .ZN(n14423) );
  INV_X1 U17697 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14416) );
  NAND2_X1 U17698 ( .A1(n14435), .A2(n14416), .ZN(n14419) );
  INV_X1 U17699 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15040) );
  NAND2_X1 U17700 ( .A1(n14437), .A2(n15040), .ZN(n14417) );
  OAI211_X1 U17701 ( .C1(n13570), .C2(P1_EBX_REG_24__SCAN_IN), .A(n14417), .B(
        n14404), .ZN(n14418) );
  MUX2_X1 U17702 ( .A(n14431), .B(n14404), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n14421) );
  NAND2_X1 U17703 ( .A1(n14432), .A2(n10181), .ZN(n14420) );
  NAND2_X1 U17704 ( .A1(n14421), .A2(n14420), .ZN(n14728) );
  MUX2_X1 U17705 ( .A(n14431), .B(n14404), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n14425) );
  INV_X1 U17706 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14882) );
  NAND2_X1 U17707 ( .A1(n14432), .A2(n14882), .ZN(n14424) );
  NAND2_X1 U17708 ( .A1(n14425), .A2(n14424), .ZN(n14715) );
  INV_X1 U17709 ( .A(n14715), .ZN(n14426) );
  INV_X1 U17710 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14427) );
  NAND2_X1 U17711 ( .A1(n14435), .A2(n14427), .ZN(n14430) );
  INV_X1 U17712 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14850) );
  NAND2_X1 U17713 ( .A1(n14437), .A2(n14850), .ZN(n14428) );
  OAI211_X1 U17714 ( .C1(n13570), .C2(P1_EBX_REG_26__SCAN_IN), .A(n14428), .B(
        n14404), .ZN(n14429) );
  NAND2_X1 U17715 ( .A1(n14430), .A2(n14429), .ZN(n14670) );
  MUX2_X1 U17716 ( .A(n14431), .B(n14404), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n14434) );
  NAND2_X1 U17717 ( .A1(n14432), .A2(n14853), .ZN(n14433) );
  NAND2_X1 U17718 ( .A1(n14434), .A2(n14433), .ZN(n14655) );
  INV_X1 U17719 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14458) );
  NAND2_X1 U17720 ( .A1(n14435), .A2(n14458), .ZN(n14440) );
  NAND2_X1 U17721 ( .A1(n14437), .A2(n14436), .ZN(n14438) );
  OAI211_X1 U17722 ( .C1(n13570), .C2(P1_EBX_REG_28__SCAN_IN), .A(n14438), .B(
        n14404), .ZN(n14439) );
  NAND2_X1 U17723 ( .A1(n14440), .A2(n14439), .ZN(n14456) );
  INV_X1 U17724 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14706) );
  NAND2_X1 U17725 ( .A1(n14441), .A2(n14706), .ZN(n14442) );
  OAI21_X1 U17726 ( .B1(n14617), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n14442), .ZN(n14443) );
  MUX2_X1 U17727 ( .A(n14443), .B(n14442), .S(n14615), .Z(n14638) );
  INV_X1 U17728 ( .A(n14641), .ZN(n14444) );
  OAI22_X1 U17729 ( .A1(n14444), .A2(n14404), .B1(n14443), .B2(n14639), .ZN(
        n14447) );
  NAND2_X1 U17730 ( .A1(n14617), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n14446) );
  NAND2_X1 U17731 ( .A1(n13570), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14445) );
  NAND2_X1 U17732 ( .A1(n14446), .A2(n14445), .ZN(n14616) );
  OAI222_X1 U17733 ( .A1(n14773), .A2(n14780), .B1(n14774), .B2(n14448), .C1(
        n14990), .C2(n14776), .ZN(P1_U2842) );
  NAND2_X2 U17734 ( .A1(n14635), .A2(n14451), .ZN(n14856) );
  AOI22_X1 U17735 ( .A1(n14828), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n14827), .ZN(n14455) );
  INV_X1 U17736 ( .A(n20053), .ZN(n14453) );
  AOI22_X1 U17737 ( .A1(n14830), .A2(n14453), .B1(n14829), .B2(DATAI_28_), 
        .ZN(n14454) );
  OAI211_X1 U17738 ( .C1(n14856), .C2(n14818), .A(n14455), .B(n14454), .ZN(
        P1_U2876) );
  OR2_X1 U17739 ( .A1(n14657), .A2(n14456), .ZN(n14457) );
  NAND2_X1 U17740 ( .A1(n14639), .A2(n14457), .ZN(n15013) );
  OAI222_X1 U17741 ( .A1(n14458), .A2(n14774), .B1(n14776), .B2(n15013), .C1(
        n14856), .C2(n14773), .ZN(P1_U2844) );
  INV_X1 U17742 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n14462) );
  INV_X1 U17743 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20763) );
  INV_X1 U17744 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20762) );
  INV_X1 U17745 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20752) );
  NAND2_X1 U17746 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n15847) );
  NOR2_X1 U17747 ( .A1(n20752), .A2(n15847), .ZN(n15816) );
  NAND4_X1 U17748 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n15816), .A3(
        P1_REIP_REG_19__SCAN_IN), .A4(P1_REIP_REG_18__SCAN_IN), .ZN(n15789) );
  NOR2_X1 U17749 ( .A1(n14459), .A2(n15789), .ZN(n15797) );
  NAND4_X1 U17750 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n15797), .A3(
        P1_REIP_REG_22__SCAN_IN), .A4(P1_REIP_REG_21__SCAN_IN), .ZN(n15781) );
  NOR2_X1 U17751 ( .A1(n20762), .A2(n15781), .ZN(n15770) );
  NAND2_X1 U17752 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n15770), .ZN(n14672) );
  NOR2_X1 U17753 ( .A1(n20763), .A2(n14672), .ZN(n14671) );
  NAND2_X1 U17754 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n14671), .ZN(n14463) );
  NOR2_X1 U17755 ( .A1(n14462), .A2(n14463), .ZN(n14646) );
  INV_X1 U17756 ( .A(n14646), .ZN(n14460) );
  NAND2_X1 U17757 ( .A1(n19945), .A2(n14460), .ZN(n14461) );
  NAND2_X1 U17758 ( .A1(n14461), .A2(n15796), .ZN(n14643) );
  OAI21_X1 U17759 ( .B1(n19934), .B2(n14463), .A(n14462), .ZN(n14467) );
  AOI22_X1 U17760 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19964), .B1(
        n19971), .B2(n14859), .ZN(n14465) );
  NAND2_X1 U17761 ( .A1(n19961), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n14464) );
  OAI211_X1 U17762 ( .C1(n15859), .C2(n15013), .A(n14465), .B(n14464), .ZN(
        n14466) );
  AOI21_X1 U17763 ( .B1(n14643), .B2(n14467), .A(n14466), .ZN(n14468) );
  OAI21_X1 U17764 ( .B1(n14856), .B2(n15867), .A(n14468), .ZN(P1_U2812) );
  NAND2_X1 U17765 ( .A1(n14470), .A2(n14469), .ZN(n14472) );
  XOR2_X1 U17766 ( .A(n14472), .B(n14471), .Z(n15445) );
  INV_X1 U17767 ( .A(n14473), .ZN(n14474) );
  AOI21_X1 U17768 ( .B1(n21072), .B2(n11886), .A(n14474), .ZN(n16056) );
  NAND2_X1 U17769 ( .A1(P2_REIP_REG_29__SCAN_IN), .A2(n19138), .ZN(n15437) );
  NAND2_X1 U17770 ( .A1(n19137), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14479) );
  OAI211_X1 U17771 ( .C1(n16059), .C2(n19157), .A(n15437), .B(n14479), .ZN(
        n14480) );
  AOI21_X1 U17772 ( .B1(n16056), .B2(n16234), .A(n14480), .ZN(n14484) );
  AOI21_X2 U17773 ( .B1(n14482), .B2(n14516), .A(n14481), .ZN(n15442) );
  NAND2_X1 U17774 ( .A1(n15442), .A2(n16228), .ZN(n14483) );
  OAI211_X1 U17775 ( .C1(n15445), .C2(n19142), .A(n14484), .B(n14483), .ZN(
        P2_U2985) );
  INV_X1 U17776 ( .A(n14485), .ZN(n16075) );
  INV_X1 U17777 ( .A(n14487), .ZN(n14490) );
  AOI21_X1 U17778 ( .B1(n14488), .B2(n14486), .A(n14487), .ZN(n16112) );
  OAI21_X1 U17779 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n13334), .A(
        n14486), .ZN(n15381) );
  INV_X1 U17780 ( .A(n15381), .ZN(n16128) );
  NOR2_X1 U17781 ( .A1(n18966), .A2(n16110), .ZN(n16103) );
  NAND2_X1 U17782 ( .A1(n14490), .A2(n10067), .ZN(n14491) );
  NAND2_X1 U17783 ( .A1(n14492), .A2(n14491), .ZN(n15363) );
  INV_X1 U17784 ( .A(n15363), .ZN(n16104) );
  NOR2_X1 U17785 ( .A1(n16103), .A2(n16104), .ZN(n16102) );
  NOR2_X1 U17786 ( .A1(n16102), .A2(n18966), .ZN(n16083) );
  AOI21_X1 U17787 ( .B1(n16085), .B2(n14492), .A(n9940), .ZN(n16084) );
  NOR2_X1 U17788 ( .A1(n16057), .A2(n16056), .ZN(n16046) );
  NOR2_X1 U17789 ( .A1(n16046), .A2(n18966), .ZN(n14493) );
  XNOR2_X1 U17790 ( .A(n14493), .B(n16047), .ZN(n14500) );
  AOI22_X1 U17791 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n18978), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n18993), .ZN(n14494) );
  OAI21_X1 U17792 ( .B1(n14495), .B2(n18982), .A(n14494), .ZN(n14496) );
  AOI21_X1 U17793 ( .B1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n18968), .A(
        n14496), .ZN(n14498) );
  NAND2_X1 U17794 ( .A1(n14564), .A2(n18984), .ZN(n14497) );
  OAI211_X1 U17795 ( .C1(n14555), .C2(n18958), .A(n14498), .B(n14497), .ZN(
        n14499) );
  AOI21_X1 U17796 ( .B1(n14500), .B2(n18961), .A(n14499), .ZN(n14501) );
  INV_X1 U17797 ( .A(n14501), .ZN(P2_U2825) );
  INV_X1 U17798 ( .A(n14503), .ZN(n14507) );
  INV_X1 U17799 ( .A(n14504), .ZN(n14506) );
  AOI21_X1 U17800 ( .B1(n14507), .B2(n14506), .A(n14505), .ZN(n16072) );
  XNOR2_X1 U17801 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14509) );
  OAI21_X1 U17802 ( .B1(n15447), .B2(n14509), .A(n14508), .ZN(n14510) );
  AOI21_X1 U17803 ( .B1(n16280), .B2(n16072), .A(n14510), .ZN(n14511) );
  OAI21_X1 U17804 ( .B1(n16071), .B2(n16272), .A(n14511), .ZN(n14512) );
  INV_X1 U17805 ( .A(n14512), .ZN(n14514) );
  OAI21_X1 U17806 ( .B1(n14519), .B2(n16278), .A(n14518), .ZN(P2_U3018) );
  OAI211_X1 U17807 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20197), .A(n14520), 
        .B(n20502), .ZN(n14523) );
  NAND2_X1 U17808 ( .A1(n14521), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n14522) );
  OAI211_X1 U17809 ( .C1(n14524), .C2(n20535), .A(n14523), .B(n14522), .ZN(
        P1_U3477) );
  INV_X1 U17810 ( .A(n14525), .ZN(n14527) );
  OAI22_X1 U17811 ( .A1(n14529), .A2(n14528), .B1(n14527), .B2(n14526), .ZN(
        n14554) );
  AOI22_X1 U17812 ( .A1(n10553), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14539), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14531) );
  AOI22_X1 U17813 ( .A1(n14537), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14530) );
  NAND2_X1 U17814 ( .A1(n14531), .A2(n14530), .ZN(n14551) );
  INV_X1 U17815 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14535) );
  AOI21_X1 U17816 ( .B1(n14532), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n14546), .ZN(n14534) );
  AOI22_X1 U17817 ( .A1(n10557), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14542), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14533) );
  OAI211_X1 U17818 ( .C1(n14536), .C2(n14535), .A(n14534), .B(n14533), .ZN(
        n14550) );
  AOI22_X1 U17819 ( .A1(n10553), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14537), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14541) );
  AOI22_X1 U17820 ( .A1(n14539), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14540) );
  NAND2_X1 U17821 ( .A1(n14541), .A2(n14540), .ZN(n14549) );
  AOI22_X1 U17822 ( .A1(n10557), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n14542), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14547) );
  NAND2_X1 U17823 ( .A1(n14543), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n14544) );
  NAND4_X1 U17824 ( .A1(n14547), .A2(n14546), .A3(n14545), .A4(n14544), .ZN(
        n14548) );
  OAI22_X1 U17825 ( .A1(n14551), .A2(n14550), .B1(n14549), .B2(n14548), .ZN(
        n14552) );
  INV_X1 U17826 ( .A(n14552), .ZN(n14553) );
  XNOR2_X1 U17827 ( .A(n14554), .B(n14553), .ZN(n14567) );
  INV_X1 U17828 ( .A(n14555), .ZN(n14561) );
  INV_X1 U17829 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n14556) );
  OR2_X1 U17830 ( .A1(n19158), .A2(n14556), .ZN(n14558) );
  NAND2_X1 U17831 ( .A1(n19158), .A2(BUF2_REG_14__SCAN_IN), .ZN(n14557) );
  AND2_X1 U17832 ( .A1(n14558), .A2(n14557), .ZN(n19002) );
  INV_X1 U17833 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n14559) );
  OAI22_X1 U17834 ( .A1(n16134), .A2(n19002), .B1(n15340), .B2(n14559), .ZN(
        n14560) );
  AOI21_X1 U17835 ( .B1(n14561), .B2(n19051), .A(n14560), .ZN(n14563) );
  AOI22_X1 U17836 ( .A1(n18999), .A2(BUF2_REG_30__SCAN_IN), .B1(n18998), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n14562) );
  OAI211_X1 U17837 ( .C1(n14567), .C2(n16136), .A(n14563), .B(n14562), .ZN(
        P2_U2889) );
  NAND2_X1 U17838 ( .A1(n14564), .A2(n15201), .ZN(n14566) );
  NAND2_X1 U17839 ( .A1(n15259), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14565) );
  OAI211_X1 U17840 ( .C1(n14567), .C2(n15261), .A(n14566), .B(n14565), .ZN(
        P2_U2857) );
  OAI21_X1 U17841 ( .B1(n14570), .B2(n14569), .A(n14568), .ZN(n14594) );
  INV_X1 U17842 ( .A(n15572), .ZN(n14573) );
  NAND2_X1 U17843 ( .A1(n14572), .A2(n14571), .ZN(n14581) );
  NAND2_X1 U17844 ( .A1(n14573), .A2(n14581), .ZN(n14574) );
  NAND2_X1 U17845 ( .A1(n19138), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n14589) );
  OAI211_X1 U17846 ( .C1(n14594), .C2(n15637), .A(n14574), .B(n14589), .ZN(
        n14587) );
  INV_X1 U17847 ( .A(n14575), .ZN(n14576) );
  AOI21_X1 U17848 ( .B1(n14578), .B2(n14577), .A(n14576), .ZN(n14580) );
  XNOR2_X1 U17849 ( .A(n14580), .B(n14579), .ZN(n14596) );
  INV_X1 U17850 ( .A(n14596), .ZN(n14585) );
  INV_X1 U17851 ( .A(n14581), .ZN(n14583) );
  AOI22_X1 U17852 ( .A1(n15574), .A2(n14583), .B1(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n14582), .ZN(n14584) );
  OAI21_X1 U17853 ( .B1(n14585), .B2(n16278), .A(n14584), .ZN(n14586) );
  AOI211_X1 U17854 ( .C1(n16280), .C2(n19820), .A(n14587), .B(n14586), .ZN(
        n14588) );
  INV_X1 U17855 ( .A(n14589), .ZN(n14590) );
  AOI21_X1 U17856 ( .B1(n19137), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n14590), .ZN(n14593) );
  NAND2_X1 U17857 ( .A1(n16234), .A2(n14591), .ZN(n14592) );
  OAI211_X1 U17858 ( .C1(n14594), .C2(n19140), .A(n14593), .B(n14592), .ZN(
        n14595) );
  AOI21_X1 U17859 ( .B1(n14596), .B2(n10996), .A(n14595), .ZN(n14597) );
  OAI21_X1 U17860 ( .B1(n14598), .B2(n19157), .A(n14597), .ZN(P2_U3012) );
  INV_X1 U17861 ( .A(n14599), .ZN(n15740) );
  INV_X1 U17862 ( .A(n14607), .ZN(n14600) );
  AOI22_X1 U17863 ( .A1(n15740), .A2(n13518), .B1(n13375), .B2(n14600), .ZN(
        n14605) );
  INV_X1 U17864 ( .A(n14601), .ZN(n14603) );
  OAI21_X1 U17865 ( .B1(n14603), .B2(n14602), .A(n15740), .ZN(n14604) );
  OAI211_X1 U17866 ( .C1(n15740), .C2(n14606), .A(n14605), .B(n14604), .ZN(
        n15723) );
  AOI21_X1 U17867 ( .B1(n14607), .B2(n13375), .A(n13518), .ZN(n14608) );
  AOI21_X1 U17868 ( .B1(n15740), .B2(n14609), .A(n14608), .ZN(n19874) );
  NAND3_X1 U17869 ( .A1(n13570), .A2(n14609), .A3(n15761), .ZN(n14610) );
  NAND2_X1 U17870 ( .A1(n14610), .A2(n20818), .ZN(n20815) );
  NAND2_X1 U17871 ( .A1(n19874), .A2(n20815), .ZN(n15729) );
  AND2_X1 U17872 ( .A1(n15729), .A2(n14611), .ZN(n19884) );
  MUX2_X1 U17873 ( .A(P1_MORE_REG_SCAN_IN), .B(n15723), .S(n19884), .Z(
        P1_U3484) );
  NAND2_X1 U17874 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(n14646), .ZN(n14630) );
  INV_X1 U17875 ( .A(n14630), .ZN(n14614) );
  NAND2_X1 U17876 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n14614), .ZN(n14612) );
  NAND2_X1 U17877 ( .A1(n19945), .A2(n14612), .ZN(n14613) );
  NAND2_X1 U17878 ( .A1(n14613), .A2(n15796), .ZN(n14631) );
  NAND2_X1 U17879 ( .A1(n14631), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n14623) );
  AOI22_X1 U17880 ( .A1(n19961), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19964), .ZN(n14622) );
  NAND4_X1 U17881 ( .A1(n19945), .A2(P1_REIP_REG_30__SCAN_IN), .A3(n20772), 
        .A4(n14614), .ZN(n14621) );
  AOI22_X1 U17882 ( .A1(n14617), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n13570), .ZN(n14618) );
  XNOR2_X1 U17883 ( .A(n14619), .B(n14618), .ZN(n14967) );
  NAND2_X1 U17884 ( .A1(n19960), .A2(n14967), .ZN(n14620) );
  NAND4_X1 U17885 ( .A1(n14623), .A2(n14622), .A3(n14621), .A4(n14620), .ZN(
        n14624) );
  AOI21_X1 U17886 ( .B1(n14625), .B2(n19928), .A(n14624), .ZN(n14626) );
  INV_X1 U17887 ( .A(n14626), .ZN(P1_U2809) );
  OAI22_X1 U17888 ( .A1(n14627), .A2(n19899), .B1(n19959), .B2(n14837), .ZN(
        n14629) );
  NOR2_X1 U17889 ( .A1(n15859), .A2(n14990), .ZN(n14628) );
  NOR2_X1 U17890 ( .A1(n19934), .A2(n14630), .ZN(n14632) );
  OAI21_X1 U17891 ( .B1(n14632), .B2(P1_REIP_REG_30__SCAN_IN), .A(n14631), 
        .ZN(n14633) );
  OAI211_X1 U17892 ( .C1(n14780), .C2(n15867), .A(n14634), .B(n14633), .ZN(
        P1_U2810) );
  NAND2_X1 U17893 ( .A1(n14639), .A2(n14638), .ZN(n14640) );
  NAND2_X1 U17894 ( .A1(n14641), .A2(n14640), .ZN(n15001) );
  INV_X1 U17895 ( .A(n15001), .ZN(n14642) );
  AOI22_X1 U17896 ( .A1(n14642), .A2(n19960), .B1(n19961), .B2(
        P1_EBX_REG_29__SCAN_IN), .ZN(n14650) );
  NAND2_X1 U17897 ( .A1(n14643), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14649) );
  INV_X1 U17898 ( .A(n14846), .ZN(n14644) );
  AOI22_X1 U17899 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19964), .B1(
        n19971), .B2(n14644), .ZN(n14648) );
  INV_X1 U17900 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n14645) );
  NAND3_X1 U17901 ( .A1(n19945), .A2(n14646), .A3(n14645), .ZN(n14647) );
  NAND4_X1 U17902 ( .A1(n14650), .A2(n14649), .A3(n14648), .A4(n14647), .ZN(
        n14651) );
  AOI21_X1 U17903 ( .B1(n14848), .B2(n19928), .A(n14651), .ZN(n14652) );
  INV_X1 U17904 ( .A(n14652), .ZN(P1_U2811) );
  AOI21_X1 U17905 ( .B1(n14654), .B2(n14653), .A(n14449), .ZN(n14868) );
  AND2_X1 U17906 ( .A1(n14669), .A2(n14655), .ZN(n14656) );
  NOR2_X1 U17907 ( .A1(n14657), .A2(n14656), .ZN(n15018) );
  AOI22_X1 U17908 ( .A1(n15018), .A2(n19960), .B1(n19961), .B2(
        P1_EBX_REG_27__SCAN_IN), .ZN(n14664) );
  INV_X1 U17909 ( .A(n14671), .ZN(n14658) );
  NAND2_X1 U17910 ( .A1(n19945), .A2(n14658), .ZN(n14659) );
  NAND2_X1 U17911 ( .A1(n14659), .A2(n15796), .ZN(n14674) );
  NAND2_X1 U17912 ( .A1(n14674), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14663) );
  INV_X1 U17913 ( .A(n14866), .ZN(n14660) );
  AOI22_X1 U17914 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n19964), .B1(
        n19971), .B2(n14660), .ZN(n14662) );
  INV_X1 U17915 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n14864) );
  NAND3_X1 U17916 ( .A1(n19945), .A2(n14671), .A3(n14864), .ZN(n14661) );
  NAND4_X1 U17917 ( .A1(n14664), .A2(n14663), .A3(n14662), .A4(n14661), .ZN(
        n14665) );
  AOI21_X1 U17918 ( .B1(n14868), .B2(n19928), .A(n14665), .ZN(n14666) );
  INV_X1 U17919 ( .A(n14666), .ZN(P1_U2813) );
  OAI21_X1 U17920 ( .B1(n14667), .B2(n14668), .A(n14653), .ZN(n14871) );
  OAI21_X1 U17921 ( .B1(n14713), .B2(n14670), .A(n14669), .ZN(n15025) );
  INV_X1 U17922 ( .A(n15025), .ZN(n14708) );
  NOR2_X1 U17923 ( .A1(n14672), .A2(n14671), .ZN(n14673) );
  AOI22_X1 U17924 ( .A1(n14708), .A2(n19960), .B1(n19945), .B2(n14673), .ZN(
        n14678) );
  NAND2_X1 U17925 ( .A1(n14674), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14677) );
  AOI22_X1 U17926 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19964), .B1(
        n19971), .B2(n14874), .ZN(n14676) );
  NAND2_X1 U17927 ( .A1(n19961), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n14675) );
  AND4_X1 U17928 ( .A1(n14678), .A2(n14677), .A3(n14676), .A4(n14675), .ZN(
        n14679) );
  OAI21_X1 U17929 ( .B1(n14871), .B2(n15867), .A(n14679), .ZN(P1_U2814) );
  NOR2_X1 U17930 ( .A1(n14681), .A2(n14682), .ZN(n14683) );
  OR2_X1 U17931 ( .A1(n14680), .A2(n14683), .ZN(n15900) );
  NAND3_X1 U17932 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(n14684), .ZN(n15815) );
  OAI21_X1 U17933 ( .B1(n15847), .B2(n15815), .A(n20752), .ZN(n14692) );
  AOI21_X1 U17934 ( .B1(n15816), .B2(n14685), .A(n14699), .ZN(n15831) );
  INV_X1 U17935 ( .A(n14686), .ZN(n15899) );
  OAI22_X1 U17936 ( .A1(n14687), .A2(n19899), .B1(n15899), .B2(n19959), .ZN(
        n14691) );
  AOI21_X1 U17937 ( .B1(n14688), .B2(n14763), .A(n9912), .ZN(n15956) );
  INV_X1 U17938 ( .A(n15956), .ZN(n14759) );
  AOI21_X1 U17939 ( .B1(n19961), .B2(P1_EBX_REG_17__SCAN_IN), .A(n19948), .ZN(
        n14689) );
  OAI21_X1 U17940 ( .B1(n15859), .B2(n14759), .A(n14689), .ZN(n14690) );
  AOI211_X1 U17941 ( .C1(n14692), .C2(n15831), .A(n14691), .B(n14690), .ZN(
        n14693) );
  OAI21_X1 U17942 ( .B1(n15900), .B2(n15867), .A(n14693), .ZN(P1_U2823) );
  NAND2_X1 U17943 ( .A1(n19899), .A2(n19959), .ZN(n14694) );
  AOI22_X1 U17944 ( .A1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n14694), .B1(
        n19965), .B2(n12524), .ZN(n14695) );
  OAI21_X1 U17945 ( .B1(n15859), .B2(n14696), .A(n14695), .ZN(n14701) );
  OAI22_X1 U17946 ( .A1(n14699), .A2(n13493), .B1(n14698), .B2(n14697), .ZN(
        n14700) );
  AOI211_X1 U17947 ( .C1(n14702), .C2(n19952), .A(n14701), .B(n14700), .ZN(
        n14703) );
  INV_X1 U17948 ( .A(n14703), .ZN(P1_U2840) );
  INV_X1 U17949 ( .A(n14967), .ZN(n14705) );
  OAI22_X1 U17950 ( .A1(n14705), .A2(n14776), .B1(n14704), .B2(n14774), .ZN(
        P1_U2841) );
  INV_X1 U17951 ( .A(n14848), .ZN(n14784) );
  OAI222_X1 U17952 ( .A1(n14706), .A2(n14774), .B1(n14776), .B2(n15001), .C1(
        n14784), .C2(n14773), .ZN(P1_U2843) );
  INV_X1 U17953 ( .A(n14868), .ZN(n14788) );
  AOI22_X1 U17954 ( .A1(n14767), .A2(n15018), .B1(n14765), .B2(
        P1_EBX_REG_27__SCAN_IN), .ZN(n14707) );
  OAI21_X1 U17955 ( .B1(n14788), .B2(n14773), .A(n14707), .ZN(P1_U2845) );
  AOI22_X1 U17956 ( .A1(n14767), .A2(n14708), .B1(n14765), .B2(
        P1_EBX_REG_26__SCAN_IN), .ZN(n14709) );
  OAI21_X1 U17957 ( .B1(n14871), .B2(n14773), .A(n14709), .ZN(P1_U2846) );
  NOR2_X1 U17958 ( .A1(n14710), .A2(n14711), .ZN(n14712) );
  OR2_X1 U17959 ( .A1(n14667), .A2(n14712), .ZN(n15775) );
  INV_X1 U17960 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14718) );
  INV_X1 U17961 ( .A(n14713), .ZN(n14717) );
  INV_X1 U17962 ( .A(n14714), .ZN(n14722) );
  NAND2_X1 U17963 ( .A1(n14722), .A2(n14715), .ZN(n14716) );
  NAND2_X1 U17964 ( .A1(n14717), .A2(n14716), .ZN(n15774) );
  OAI222_X1 U17965 ( .A1(n14773), .A2(n15775), .B1(n14774), .B2(n14718), .C1(
        n15774), .C2(n14776), .ZN(P1_U2847) );
  AOI21_X1 U17966 ( .B1(n14720), .B2(n14719), .A(n14710), .ZN(n14892) );
  INV_X1 U17967 ( .A(n14892), .ZN(n15784) );
  OAI21_X1 U17968 ( .B1(n14728), .B2(n14731), .A(n10306), .ZN(n14721) );
  NAND2_X1 U17969 ( .A1(n14722), .A2(n14721), .ZN(n15783) );
  INV_X1 U17970 ( .A(n15783), .ZN(n14723) );
  AOI22_X1 U17971 ( .A1(n14767), .A2(n14723), .B1(n14765), .B2(
        P1_EBX_REG_24__SCAN_IN), .ZN(n14724) );
  OAI21_X1 U17972 ( .B1(n15784), .B2(n14773), .A(n14724), .ZN(P1_U2848) );
  INV_X1 U17973 ( .A(n14719), .ZN(n14726) );
  AOI21_X1 U17974 ( .B1(n14727), .B2(n9847), .A(n14726), .ZN(n15875) );
  INV_X1 U17975 ( .A(n15875), .ZN(n14803) );
  XNOR2_X1 U17976 ( .A(n14728), .B(n14731), .ZN(n15790) );
  INV_X1 U17977 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14729) );
  OAI222_X1 U17978 ( .A1(n14773), .A2(n14803), .B1(n14776), .B2(n15790), .C1(
        n14729), .C2(n14774), .ZN(P1_U2849) );
  OR2_X1 U17979 ( .A1(n14730), .A2(n14738), .ZN(n14732) );
  NAND2_X1 U17980 ( .A1(n14732), .A2(n14731), .ZN(n15058) );
  NAND2_X1 U17981 ( .A1(n14733), .A2(n14734), .ZN(n14735) );
  AND2_X1 U17982 ( .A1(n9847), .A2(n14735), .ZN(n15800) );
  INV_X1 U17983 ( .A(n15800), .ZN(n14807) );
  OAI222_X1 U17984 ( .A1(n15058), .A2(n14776), .B1(n14774), .B2(n14410), .C1(
        n14773), .C2(n14807), .ZN(P1_U2850) );
  OAI21_X1 U17985 ( .B1(n14736), .B2(n14737), .A(n14733), .ZN(n15810) );
  AOI21_X1 U17986 ( .B1(n14739), .B2(n14742), .A(n14738), .ZN(n15811) );
  AOI22_X1 U17987 ( .A1(n14767), .A2(n15811), .B1(n14765), .B2(
        P1_EBX_REG_21__SCAN_IN), .ZN(n14740) );
  OAI21_X1 U17988 ( .B1(n15810), .B2(n14773), .A(n14740), .ZN(P1_U2851) );
  OR2_X1 U17989 ( .A1(n14741), .A2(n14749), .ZN(n14743) );
  NAND2_X1 U17990 ( .A1(n14743), .A2(n14742), .ZN(n15817) );
  AOI21_X1 U17991 ( .B1(n14745), .B2(n10121), .A(n14736), .ZN(n14746) );
  INV_X1 U17992 ( .A(n14746), .ZN(n15818) );
  OAI222_X1 U17993 ( .A1(n15817), .A2(n14776), .B1(n14774), .B2(n14406), .C1(
        n14773), .C2(n15818), .ZN(P1_U2852) );
  AOI21_X1 U17994 ( .B1(n14748), .B2(n14747), .A(n14744), .ZN(n15887) );
  INV_X1 U17995 ( .A(n15887), .ZN(n14822) );
  AOI21_X1 U17996 ( .B1(n14750), .B2(n14754), .A(n14749), .ZN(n15948) );
  AOI22_X1 U17997 ( .A1(n14767), .A2(n15948), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n14765), .ZN(n14751) );
  OAI21_X1 U17998 ( .B1(n14822), .B2(n14773), .A(n14751), .ZN(P1_U2853) );
  OAI21_X1 U17999 ( .B1(n14680), .B2(n14752), .A(n14747), .ZN(n15834) );
  OR2_X1 U18000 ( .A1(n14753), .A2(n9912), .ZN(n14755) );
  NAND2_X1 U18001 ( .A1(n14755), .A2(n14754), .ZN(n15833) );
  INV_X1 U18002 ( .A(n15833), .ZN(n14756) );
  AOI22_X1 U18003 ( .A1(n14767), .A2(n14756), .B1(n14765), .B2(
        P1_EBX_REG_18__SCAN_IN), .ZN(n14757) );
  OAI21_X1 U18004 ( .B1(n15834), .B2(n14773), .A(n14757), .ZN(P1_U2854) );
  INV_X1 U18005 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14758) );
  OAI222_X1 U18006 ( .A1(n14759), .A2(n14776), .B1(n14758), .B2(n14774), .C1(
        n15900), .C2(n14773), .ZN(P1_U2855) );
  AOI21_X1 U18007 ( .B1(n14761), .B2(n14760), .A(n14681), .ZN(n14920) );
  INV_X1 U18008 ( .A(n14920), .ZN(n15843) );
  OR2_X1 U18009 ( .A1(n14762), .A2(n14769), .ZN(n14764) );
  NAND2_X1 U18010 ( .A1(n14764), .A2(n14763), .ZN(n15842) );
  INV_X1 U18011 ( .A(n15842), .ZN(n14766) );
  AOI22_X1 U18012 ( .A1(n14767), .A2(n14766), .B1(n14765), .B2(
        P1_EBX_REG_16__SCAN_IN), .ZN(n14768) );
  OAI21_X1 U18013 ( .B1(n15843), .B2(n14773), .A(n14768), .ZN(P1_U2856) );
  AOI21_X1 U18014 ( .B1(n14771), .B2(n14770), .A(n14769), .ZN(n15850) );
  INV_X1 U18015 ( .A(n15850), .ZN(n15963) );
  INV_X1 U18016 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14775) );
  OAI222_X1 U18017 ( .A1(n15963), .A2(n14776), .B1(n14775), .B2(n14774), .C1(
        n14773), .C2(n14772), .ZN(P1_U2857) );
  AOI22_X1 U18018 ( .A1(n14828), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n14827), .ZN(n14779) );
  INV_X1 U18019 ( .A(n20058), .ZN(n14777) );
  AOI22_X1 U18020 ( .A1(n14830), .A2(n14777), .B1(n14829), .B2(DATAI_30_), 
        .ZN(n14778) );
  OAI211_X1 U18021 ( .C1(n14780), .C2(n14818), .A(n14779), .B(n14778), .ZN(
        P1_U2874) );
  AOI22_X1 U18022 ( .A1(n14828), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n14827), .ZN(n14783) );
  INV_X1 U18023 ( .A(n20055), .ZN(n14781) );
  AOI22_X1 U18024 ( .A1(n14830), .A2(n14781), .B1(n14829), .B2(DATAI_29_), 
        .ZN(n14782) );
  OAI211_X1 U18025 ( .C1(n14784), .C2(n14818), .A(n14783), .B(n14782), .ZN(
        P1_U2875) );
  AOI22_X1 U18026 ( .A1(n14828), .A2(BUF1_REG_27__SCAN_IN), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(n14827), .ZN(n14787) );
  INV_X1 U18027 ( .A(n20051), .ZN(n14785) );
  AOI22_X1 U18028 ( .A1(n14830), .A2(n14785), .B1(n14829), .B2(DATAI_27_), 
        .ZN(n14786) );
  OAI211_X1 U18029 ( .C1(n14788), .C2(n14818), .A(n14787), .B(n14786), .ZN(
        P1_U2877) );
  AOI22_X1 U18030 ( .A1(n14828), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n14827), .ZN(n14791) );
  INV_X1 U18031 ( .A(n20049), .ZN(n14789) );
  AOI22_X1 U18032 ( .A1(n14830), .A2(n14789), .B1(n14829), .B2(DATAI_26_), 
        .ZN(n14790) );
  OAI211_X1 U18033 ( .C1(n14871), .C2(n14818), .A(n14791), .B(n14790), .ZN(
        P1_U2878) );
  AOI22_X1 U18034 ( .A1(n14828), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n14827), .ZN(n14794) );
  INV_X1 U18035 ( .A(n20047), .ZN(n14792) );
  AOI22_X1 U18036 ( .A1(n14830), .A2(n14792), .B1(n14829), .B2(DATAI_25_), 
        .ZN(n14793) );
  OAI211_X1 U18037 ( .C1(n15775), .C2(n14818), .A(n14794), .B(n14793), .ZN(
        P1_U2879) );
  AOI22_X1 U18038 ( .A1(n14828), .A2(BUF1_REG_24__SCAN_IN), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(n14827), .ZN(n14797) );
  INV_X1 U18039 ( .A(n20045), .ZN(n14795) );
  AOI22_X1 U18040 ( .A1(n14830), .A2(n14795), .B1(n14829), .B2(DATAI_24_), 
        .ZN(n14796) );
  OAI211_X1 U18041 ( .C1(n15784), .C2(n14818), .A(n14797), .B(n14796), .ZN(
        P1_U2880) );
  INV_X1 U18042 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n14799) );
  OAI22_X1 U18043 ( .A1(n14810), .A2(n14799), .B1(n14798), .B2(n14808), .ZN(
        n14801) );
  INV_X1 U18044 ( .A(n14830), .ZN(n14811) );
  NOR2_X1 U18045 ( .A1(n14811), .A2(n20165), .ZN(n14800) );
  AOI211_X1 U18046 ( .C1(n14829), .C2(DATAI_23_), .A(n14801), .B(n14800), .ZN(
        n14802) );
  OAI21_X1 U18047 ( .B1(n14803), .B2(n14818), .A(n14802), .ZN(P1_U2881) );
  AOI22_X1 U18048 ( .A1(n14828), .A2(BUF1_REG_22__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n14827), .ZN(n14806) );
  INV_X1 U18049 ( .A(n20159), .ZN(n14804) );
  AOI22_X1 U18050 ( .A1(n14830), .A2(n14804), .B1(n14829), .B2(DATAI_22_), 
        .ZN(n14805) );
  OAI211_X1 U18051 ( .C1(n14807), .C2(n14818), .A(n14806), .B(n14805), .ZN(
        P1_U2882) );
  INV_X1 U18052 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n15308) );
  OAI22_X1 U18053 ( .A1(n14810), .A2(n15308), .B1(n14809), .B2(n14808), .ZN(
        n14813) );
  NOR2_X1 U18054 ( .A1(n14811), .A2(n20155), .ZN(n14812) );
  AOI211_X1 U18055 ( .C1(n14829), .C2(DATAI_21_), .A(n14813), .B(n14812), .ZN(
        n14814) );
  OAI21_X1 U18056 ( .B1(n15810), .B2(n14818), .A(n14814), .ZN(P1_U2883) );
  AOI22_X1 U18057 ( .A1(n14828), .A2(BUF1_REG_20__SCAN_IN), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(n14827), .ZN(n14817) );
  INV_X1 U18058 ( .A(n20151), .ZN(n14815) );
  AOI22_X1 U18059 ( .A1(n14830), .A2(n14815), .B1(n14829), .B2(DATAI_20_), 
        .ZN(n14816) );
  OAI211_X1 U18060 ( .C1(n15818), .C2(n14818), .A(n14817), .B(n14816), .ZN(
        P1_U2884) );
  AOI22_X1 U18061 ( .A1(n14828), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n14827), .ZN(n14821) );
  INV_X1 U18062 ( .A(n20147), .ZN(n14819) );
  AOI22_X1 U18063 ( .A1(n14830), .A2(n14819), .B1(n14829), .B2(DATAI_19_), 
        .ZN(n14820) );
  OAI211_X1 U18064 ( .C1(n14822), .C2(n14818), .A(n14821), .B(n14820), .ZN(
        P1_U2885) );
  AOI22_X1 U18065 ( .A1(n14828), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n14827), .ZN(n14824) );
  AOI22_X1 U18066 ( .A1(n14830), .A2(n20020), .B1(n14829), .B2(DATAI_18_), 
        .ZN(n14823) );
  OAI211_X1 U18067 ( .C1(n15834), .C2(n14818), .A(n14824), .B(n14823), .ZN(
        P1_U2886) );
  AOI22_X1 U18068 ( .A1(n14828), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n14827), .ZN(n14826) );
  AOI22_X1 U18069 ( .A1(n14830), .A2(n20017), .B1(n14829), .B2(DATAI_17_), 
        .ZN(n14825) );
  OAI211_X1 U18070 ( .C1(n15900), .C2(n14818), .A(n14826), .B(n14825), .ZN(
        P1_U2887) );
  AOI22_X1 U18071 ( .A1(n14828), .A2(BUF1_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n14827), .ZN(n14832) );
  AOI22_X1 U18072 ( .A1(n14830), .A2(n20014), .B1(n14829), .B2(DATAI_16_), 
        .ZN(n14831) );
  OAI211_X1 U18073 ( .C1(n15843), .C2(n14818), .A(n14832), .B(n14831), .ZN(
        P1_U2888) );
  INV_X1 U18074 ( .A(n14842), .ZN(n14835) );
  INV_X1 U18075 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n20774) );
  NOR2_X1 U18076 ( .A1(n20102), .A2(n20774), .ZN(n14991) );
  AOI21_X1 U18077 ( .B1(n20065), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n14991), .ZN(n14836) );
  OAI21_X1 U18078 ( .B1(n20076), .B2(n14837), .A(n14836), .ZN(n14838) );
  AOI21_X1 U18079 ( .B1(n14839), .B2(n20071), .A(n14838), .ZN(n14840) );
  OAI21_X1 U18080 ( .B1(n14998), .B2(n19882), .A(n14840), .ZN(P1_U2969) );
  NAND2_X1 U18081 ( .A1(n14842), .A2(n14841), .ZN(n14843) );
  XNOR2_X1 U18082 ( .A(n14844), .B(n14843), .ZN(n15006) );
  NAND2_X1 U18083 ( .A1(n13703), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n15000) );
  NAND2_X1 U18084 ( .A1(n20065), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14845) );
  OAI211_X1 U18085 ( .C1(n20076), .C2(n14846), .A(n15000), .B(n14845), .ZN(
        n14847) );
  AOI21_X1 U18086 ( .B1(n14848), .B2(n20071), .A(n14847), .ZN(n14849) );
  OAI21_X1 U18087 ( .B1(n19882), .B2(n15006), .A(n14849), .ZN(P1_U2970) );
  AOI21_X2 U18088 ( .B1(n13225), .B2(n14977), .A(n14886), .ZN(n14854) );
  NOR2_X1 U18089 ( .A1(n13225), .A2(n14853), .ZN(n14852) );
  NAND2_X1 U18090 ( .A1(n14882), .A2(n14850), .ZN(n15027) );
  NOR3_X1 U18091 ( .A1(n15027), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14851) );
  OAI22_X1 U18092 ( .A1(n14854), .A2(n14851), .B1(n15895), .B2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14861) );
  XNOR2_X1 U18093 ( .A(n14855), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15016) );
  NAND2_X1 U18094 ( .A1(n13703), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n15011) );
  OAI21_X1 U18095 ( .B1(n14940), .B2(n20977), .A(n15011), .ZN(n14858) );
  NOR2_X1 U18096 ( .A1(n14856), .A2(n20120), .ZN(n14857) );
  AOI211_X2 U18097 ( .C1(n15917), .C2(n14859), .A(n14858), .B(n14857), .ZN(
        n14860) );
  OAI21_X1 U18098 ( .B1(n19882), .B2(n15016), .A(n14860), .ZN(P1_U2971) );
  INV_X1 U18099 ( .A(n14870), .ZN(n14862) );
  NOR2_X1 U18100 ( .A1(n20102), .A2(n14864), .ZN(n15017) );
  AOI21_X1 U18101 ( .B1(n20065), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15017), .ZN(n14865) );
  OAI21_X1 U18102 ( .B1(n20076), .B2(n14866), .A(n14865), .ZN(n14867) );
  AOI21_X1 U18103 ( .B1(n14868), .B2(n20071), .A(n14867), .ZN(n14869) );
  OAI21_X1 U18104 ( .B1(n19882), .B2(n15021), .A(n14869), .ZN(P1_U2972) );
  XNOR2_X1 U18105 ( .A(n14870), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15031) );
  NAND2_X1 U18106 ( .A1(n13703), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n15024) );
  OAI21_X1 U18107 ( .B1(n14940), .B2(n20887), .A(n15024), .ZN(n14873) );
  NOR2_X1 U18108 ( .A1(n14871), .A2(n20120), .ZN(n14872) );
  OAI21_X1 U18109 ( .B1(n19882), .B2(n15031), .A(n14875), .ZN(P1_U2973) );
  INV_X1 U18110 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n14876) );
  NOR2_X1 U18111 ( .A1(n20102), .A2(n14876), .ZN(n15035) );
  NOR2_X1 U18112 ( .A1(n20076), .A2(n15779), .ZN(n14877) );
  AOI211_X1 U18113 ( .C1(n20065), .C2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n15035), .B(n14877), .ZN(n14885) );
  INV_X1 U18114 ( .A(n14878), .ZN(n14879) );
  OAI21_X1 U18115 ( .B1(n14879), .B2(n15895), .A(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14888) );
  MUX2_X1 U18116 ( .A(n15040), .B(n14880), .S(n15895), .Z(n14881) );
  XNOR2_X1 U18117 ( .A(n14883), .B(n14882), .ZN(n15033) );
  NAND2_X1 U18118 ( .A1(n15033), .A2(n20072), .ZN(n14884) );
  OAI211_X1 U18119 ( .C1(n15775), .C2(n20120), .A(n14885), .B(n14884), .ZN(
        P1_U2974) );
  NAND2_X1 U18120 ( .A1(n14888), .A2(n14886), .ZN(n14887) );
  MUX2_X1 U18121 ( .A(n14888), .B(n14887), .S(n15895), .Z(n14889) );
  XNOR2_X1 U18122 ( .A(n14889), .B(n15040), .ZN(n15048) );
  NAND2_X1 U18123 ( .A1(n15917), .A2(n15786), .ZN(n14890) );
  NAND2_X1 U18124 ( .A1(n13703), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n15043) );
  OAI211_X1 U18125 ( .C1(n14940), .C2(n20903), .A(n14890), .B(n15043), .ZN(
        n14891) );
  AOI21_X1 U18126 ( .B1(n14892), .B2(n20071), .A(n14891), .ZN(n14893) );
  OAI21_X1 U18127 ( .B1(n19882), .B2(n15048), .A(n14893), .ZN(P1_U2975) );
  NAND2_X1 U18128 ( .A1(n14895), .A2(n14894), .ZN(n14896) );
  XOR2_X1 U18129 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n14896), .Z(
        n15071) );
  INV_X1 U18130 ( .A(n15798), .ZN(n14898) );
  NAND2_X1 U18131 ( .A1(n20065), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14897) );
  NAND2_X1 U18132 ( .A1(n13703), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n15059) );
  OAI211_X1 U18133 ( .C1(n20076), .C2(n14898), .A(n14897), .B(n15059), .ZN(
        n14899) );
  AOI21_X1 U18134 ( .B1(n15800), .B2(n20071), .A(n14899), .ZN(n14900) );
  OAI21_X1 U18135 ( .B1(n19882), .B2(n15071), .A(n14900), .ZN(P1_U2977) );
  NAND2_X1 U18136 ( .A1(n13703), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15076) );
  OR2_X1 U18137 ( .A1(n13225), .A2(n14901), .ZN(n15746) );
  NAND2_X1 U18138 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n13225), .ZN(
        n14903) );
  XNOR2_X1 U18139 ( .A(n14904), .B(n13248), .ZN(n15075) );
  NAND2_X1 U18140 ( .A1(n20072), .A2(n15075), .ZN(n14905) );
  OAI211_X1 U18141 ( .C1(n14940), .C2(n15824), .A(n15076), .B(n14905), .ZN(
        n14906) );
  AOI21_X1 U18142 ( .B1(n15917), .B2(n15814), .A(n14906), .ZN(n14907) );
  OAI21_X1 U18143 ( .B1(n15818), .B2(n20120), .A(n14907), .ZN(P1_U2979) );
  NAND2_X1 U18144 ( .A1(n13703), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n15089) );
  OAI21_X1 U18145 ( .B1(n14940), .B2(n20923), .A(n15089), .ZN(n14908) );
  AOI21_X1 U18146 ( .B1(n15837), .B2(n15917), .A(n14908), .ZN(n14911) );
  NAND3_X1 U18147 ( .A1(n15087), .A2(n14902), .A3(n20072), .ZN(n14910) );
  OAI211_X1 U18148 ( .C1(n15834), .C2(n20120), .A(n14911), .B(n14910), .ZN(
        P1_U2981) );
  OR2_X1 U18149 ( .A1(n14912), .A2(n14913), .ZN(n14915) );
  INV_X1 U18150 ( .A(n14914), .ZN(n14922) );
  NAND2_X1 U18151 ( .A1(n14915), .A2(n14922), .ZN(n15905) );
  OAI21_X1 U18152 ( .B1(n15905), .B2(n15892), .A(n15907), .ZN(n14916) );
  XOR2_X1 U18153 ( .A(n14917), .B(n14916), .Z(n15101) );
  NAND2_X1 U18154 ( .A1(n15917), .A2(n15846), .ZN(n14918) );
  NAND2_X1 U18155 ( .A1(n13703), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n15096) );
  OAI211_X1 U18156 ( .C1(n14940), .C2(n15841), .A(n14918), .B(n15096), .ZN(
        n14919) );
  AOI21_X1 U18157 ( .B1(n14920), .B2(n20071), .A(n14919), .ZN(n14921) );
  OAI21_X1 U18158 ( .B1(n15101), .B2(n19882), .A(n14921), .ZN(P1_U2983) );
  NAND2_X1 U18159 ( .A1(n14912), .A2(n14922), .ZN(n15893) );
  INV_X1 U18160 ( .A(n13234), .ZN(n14923) );
  AOI21_X1 U18161 ( .B1(n15893), .B2(n14924), .A(n14923), .ZN(n14926) );
  XNOR2_X1 U18162 ( .A(n13225), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14925) );
  XNOR2_X1 U18163 ( .A(n14926), .B(n14925), .ZN(n15114) );
  NAND2_X1 U18164 ( .A1(n15114), .A2(n20072), .ZN(n14932) );
  INV_X1 U18165 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n14927) );
  OR2_X1 U18166 ( .A1(n20102), .A2(n14927), .ZN(n15110) );
  INV_X1 U18167 ( .A(n15110), .ZN(n14930) );
  NOR2_X1 U18168 ( .A1(n20076), .A2(n14928), .ZN(n14929) );
  AOI211_X1 U18169 ( .C1(n20065), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n14930), .B(n14929), .ZN(n14931) );
  OAI211_X1 U18170 ( .C1(n20120), .C2(n14933), .A(n14932), .B(n14931), .ZN(
        P1_U2985) );
  INV_X1 U18171 ( .A(n14912), .ZN(n15921) );
  INV_X1 U18172 ( .A(n14934), .ZN(n14935) );
  AOI21_X1 U18173 ( .B1(n15921), .B2(n14936), .A(n14935), .ZN(n15118) );
  NAND3_X1 U18174 ( .A1(n15118), .A2(n15119), .A3(n14937), .ZN(n15120) );
  NAND2_X1 U18175 ( .A1(n15120), .A2(n15119), .ZN(n14938) );
  XOR2_X1 U18176 ( .A(n14939), .B(n14938), .Z(n15975) );
  NAND2_X1 U18177 ( .A1(n15975), .A2(n20072), .ZN(n14944) );
  OAI22_X1 U18178 ( .A1(n14940), .A2(n14290), .B1(n20102), .B2(n20746), .ZN(
        n14941) );
  AOI21_X1 U18179 ( .B1(n15917), .B2(n14942), .A(n14941), .ZN(n14943) );
  OAI211_X1 U18180 ( .C1(n20120), .C2(n14945), .A(n14944), .B(n14943), .ZN(
        P1_U2986) );
  NAND2_X1 U18181 ( .A1(n14948), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14947) );
  XNOR2_X1 U18182 ( .A(n15921), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14946) );
  MUX2_X1 U18183 ( .A(n14947), .B(n14946), .S(n13225), .Z(n14949) );
  OR3_X1 U18184 ( .A1(n14948), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n13225), .ZN(n15922) );
  NAND2_X1 U18185 ( .A1(n14949), .A2(n15922), .ZN(n15994) );
  INV_X1 U18186 ( .A(n15994), .ZN(n14955) );
  AOI22_X1 U18187 ( .A1(n20065), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n13703), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14950) );
  OAI21_X1 U18188 ( .B1(n20076), .B2(n14951), .A(n14950), .ZN(n14952) );
  AOI21_X1 U18189 ( .B1(n14953), .B2(n20071), .A(n14952), .ZN(n14954) );
  OAI21_X1 U18190 ( .B1(n14955), .B2(n19882), .A(n14954), .ZN(P1_U2989) );
  INV_X1 U18191 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14956) );
  INV_X1 U18192 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16019) );
  NOR3_X1 U18193 ( .A1(n16019), .A2(n16024), .A3(n15935), .ZN(n15989) );
  NAND3_X1 U18194 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n15989), .ZN(n15125) );
  NOR2_X1 U18195 ( .A1(n14956), .A2(n15125), .ZN(n15131) );
  NAND2_X1 U18196 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15131), .ZN(
        n14968) );
  NAND2_X1 U18197 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20081) );
  NOR2_X1 U18198 ( .A1(n16035), .A2(n20081), .ZN(n15117) );
  INV_X1 U18199 ( .A(n15117), .ZN(n14959) );
  AOI21_X1 U18200 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20100) );
  NOR2_X1 U18201 ( .A1(n14959), .A2(n20100), .ZN(n15988) );
  INV_X1 U18202 ( .A(n15988), .ZN(n15124) );
  NOR2_X1 U18203 ( .A1(n14968), .A2(n15124), .ZN(n15106) );
  NAND2_X1 U18204 ( .A1(n20078), .A2(n15106), .ZN(n15060) );
  NOR2_X1 U18205 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15971), .ZN(
        n15141) );
  NOR3_X1 U18206 ( .A1(n14972), .A2(n15141), .A3(n20098), .ZN(n20094) );
  NAND2_X1 U18207 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n20094), .ZN(
        n16011) );
  NOR2_X1 U18208 ( .A1(n14959), .A2(n16011), .ZN(n15128) );
  NOR2_X1 U18209 ( .A1(n15970), .A2(n14968), .ZN(n14960) );
  NAND2_X1 U18210 ( .A1(n15128), .A2(n14960), .ZN(n15042) );
  OAI21_X1 U18211 ( .B1(n15970), .B2(n15060), .A(n15042), .ZN(n15109) );
  NAND4_X1 U18212 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15088) );
  NOR2_X1 U18213 ( .A1(n15094), .A2(n15088), .ZN(n14971) );
  AND4_X1 U18214 ( .A1(n14971), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A4(n15074), .ZN(n14961) );
  NAND2_X1 U18215 ( .A1(n15109), .A2(n14961), .ZN(n15057) );
  INV_X1 U18216 ( .A(n14962), .ZN(n14963) );
  NOR2_X1 U18217 ( .A1(n15057), .A2(n14963), .ZN(n15032) );
  AND2_X1 U18218 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14982) );
  NAND2_X1 U18219 ( .A1(n15032), .A2(n14982), .ZN(n15020) );
  INV_X1 U18220 ( .A(n14984), .ZN(n15008) );
  OR3_X1 U18221 ( .A1(n15020), .A2(n15008), .A3(n14964), .ZN(n14993) );
  NOR3_X1 U18222 ( .A1(n14993), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n10016), .ZN(n14965) );
  AOI211_X1 U18223 ( .C1(n20110), .C2(n14967), .A(n14966), .B(n14965), .ZN(
        n14988) );
  NAND3_X1 U18224 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n15117), .ZN(n15126) );
  NOR2_X1 U18225 ( .A1(n15126), .A2(n14968), .ZN(n15972) );
  NAND2_X1 U18226 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15972), .ZN(
        n15104) );
  NAND2_X1 U18227 ( .A1(n15103), .A2(n20099), .ZN(n14969) );
  NAND2_X1 U18228 ( .A1(n15136), .A2(n14969), .ZN(n20095) );
  AOI21_X1 U18229 ( .B1(n20096), .B2(n15104), .A(n20095), .ZN(n15083) );
  INV_X1 U18230 ( .A(n15106), .ZN(n15085) );
  NAND2_X1 U18231 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14971), .ZN(
        n15062) );
  OAI21_X1 U18232 ( .B1(n15085), .B2(n15062), .A(n20078), .ZN(n14970) );
  OAI211_X1 U18233 ( .C1(n14972), .C2(n14971), .A(n15083), .B(n14970), .ZN(
        n15947) );
  INV_X1 U18234 ( .A(n20095), .ZN(n15990) );
  NAND2_X1 U18235 ( .A1(n15142), .A2(n15990), .ZN(n15991) );
  OAI21_X1 U18236 ( .B1(n15745), .B2(n15947), .A(n15991), .ZN(n15752) );
  INV_X1 U18237 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14973) );
  NOR2_X1 U18238 ( .A1(n21010), .A2(n14973), .ZN(n15064) );
  OR2_X1 U18239 ( .A1(n15142), .A2(n15064), .ZN(n14974) );
  AND2_X1 U18240 ( .A1(n15752), .A2(n14974), .ZN(n15051) );
  NAND2_X1 U18241 ( .A1(n20078), .A2(n10181), .ZN(n14975) );
  AND2_X1 U18242 ( .A1(n15051), .A2(n14975), .ZN(n15041) );
  NAND2_X1 U18243 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14976) );
  NAND2_X1 U18244 ( .A1(n15103), .A2(n14976), .ZN(n14979) );
  NAND2_X1 U18245 ( .A1(n15971), .A2(n14977), .ZN(n14978) );
  OAI211_X1 U18246 ( .C1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n20104), .A(
        n14979), .B(n14978), .ZN(n14980) );
  INV_X1 U18247 ( .A(n14980), .ZN(n14981) );
  NAND2_X1 U18248 ( .A1(n15041), .A2(n14981), .ZN(n15036) );
  INV_X1 U18249 ( .A(n15142), .ZN(n16012) );
  OR2_X1 U18250 ( .A1(n15036), .A2(n16012), .ZN(n14986) );
  INV_X1 U18251 ( .A(n14982), .ZN(n15028) );
  OR2_X1 U18252 ( .A1(n15036), .A2(n15028), .ZN(n14983) );
  NAND2_X1 U18253 ( .A1(n14986), .A2(n14983), .ZN(n15007) );
  OR2_X1 U18254 ( .A1(n15142), .A2(n14984), .ZN(n14985) );
  AND2_X1 U18255 ( .A1(n15007), .A2(n14985), .ZN(n14999) );
  OAI211_X1 U18256 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15142), .A(
        n14999), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14994) );
  NAND3_X1 U18257 ( .A1(n14994), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14986), .ZN(n14987) );
  OAI211_X1 U18258 ( .C1(n14989), .C2(n20105), .A(n14988), .B(n14987), .ZN(
        P1_U3000) );
  INV_X1 U18259 ( .A(n14990), .ZN(n14992) );
  AOI21_X1 U18260 ( .B1(n14992), .B2(n20110), .A(n14991), .ZN(n14997) );
  INV_X1 U18261 ( .A(n14993), .ZN(n14995) );
  OAI21_X1 U18262 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n14995), .A(
        n14994), .ZN(n14996) );
  OAI211_X1 U18263 ( .C1(n14998), .C2(n20105), .A(n14997), .B(n14996), .ZN(
        P1_U3001) );
  INV_X1 U18264 ( .A(n14999), .ZN(n15004) );
  OAI21_X1 U18265 ( .B1(n16014), .B2(n15001), .A(n15000), .ZN(n15003) );
  NOR3_X1 U18266 ( .A1(n15020), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n15008), .ZN(n15002) );
  AOI211_X1 U18267 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15004), .A(
        n15003), .B(n15002), .ZN(n15005) );
  OAI21_X1 U18268 ( .B1(n15006), .B2(n20105), .A(n15005), .ZN(P1_U3002) );
  INV_X1 U18269 ( .A(n15007), .ZN(n15023) );
  INV_X1 U18270 ( .A(n15020), .ZN(n15010) );
  NAND3_X1 U18271 ( .A1(n15010), .A2(n15009), .A3(n15008), .ZN(n15012) );
  OAI211_X1 U18272 ( .C1(n16014), .C2(n15013), .A(n15012), .B(n15011), .ZN(
        n15014) );
  AOI21_X1 U18273 ( .B1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n15023), .A(
        n15014), .ZN(n15015) );
  OAI21_X1 U18274 ( .B1(n15016), .B2(n20105), .A(n15015), .ZN(P1_U3003) );
  AOI21_X1 U18275 ( .B1(n20110), .B2(n15018), .A(n15017), .ZN(n15019) );
  OAI21_X1 U18276 ( .B1(n15020), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15019), .ZN(n15022) );
  OAI21_X1 U18277 ( .B1(n16014), .B2(n15025), .A(n15024), .ZN(n15026) );
  AOI21_X1 U18278 ( .B1(n15036), .B2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15026), .ZN(n15030) );
  NAND3_X1 U18279 ( .A1(n15032), .A2(n15028), .A3(n15027), .ZN(n15029) );
  OAI211_X1 U18280 ( .C1(n15031), .C2(n20105), .A(n15030), .B(n15029), .ZN(
        P1_U3005) );
  INV_X1 U18281 ( .A(n15032), .ZN(n15039) );
  NAND2_X1 U18282 ( .A1(n15033), .A2(n20087), .ZN(n15038) );
  NOR2_X1 U18283 ( .A1(n16014), .A2(n15774), .ZN(n15034) );
  AOI211_X1 U18284 ( .C1(n15036), .C2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15035), .B(n15034), .ZN(n15037) );
  OAI211_X1 U18285 ( .C1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n15039), .A(
        n15038), .B(n15037), .ZN(P1_U3006) );
  OAI21_X1 U18286 ( .B1(n15057), .B2(n10181), .A(n15040), .ZN(n15046) );
  OAI211_X1 U18287 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n15042), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n15041), .ZN(n15045) );
  OAI21_X1 U18288 ( .B1(n16014), .B2(n15783), .A(n15043), .ZN(n15044) );
  AOI21_X1 U18289 ( .B1(n15046), .B2(n15045), .A(n15044), .ZN(n15047) );
  OAI21_X1 U18290 ( .B1(n15048), .B2(n20105), .A(n15047), .ZN(P1_U3007) );
  XNOR2_X1 U18291 ( .A(n13225), .B(n10181), .ZN(n15049) );
  XNOR2_X1 U18292 ( .A(n15050), .B(n15049), .ZN(n15874) );
  NAND2_X1 U18293 ( .A1(n15874), .A2(n20087), .ZN(n15056) );
  INV_X1 U18294 ( .A(n15051), .ZN(n15054) );
  INV_X1 U18295 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n15052) );
  OAI22_X1 U18296 ( .A1(n16014), .A2(n15790), .B1(n20102), .B2(n15052), .ZN(
        n15053) );
  AOI21_X1 U18297 ( .B1(n15054), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15053), .ZN(n15055) );
  OAI211_X1 U18298 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n15057), .A(
        n15056), .B(n15055), .ZN(P1_U3008) );
  INV_X1 U18299 ( .A(n15058), .ZN(n15799) );
  INV_X1 U18300 ( .A(n15059), .ZN(n15069) );
  NAND3_X1 U18301 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15972), .A3(
        n15103), .ZN(n15061) );
  NAND2_X1 U18302 ( .A1(n15061), .A2(n15060), .ZN(n15973) );
  INV_X1 U18303 ( .A(n15062), .ZN(n15063) );
  OAI221_X1 U18304 ( .B1(n15973), .B2(n15972), .C1(n15973), .C2(n15971), .A(
        n15063), .ZN(n15952) );
  NOR2_X1 U18305 ( .A1(n15952), .A2(n15745), .ZN(n15744) );
  INV_X1 U18306 ( .A(n15064), .ZN(n15065) );
  NAND2_X1 U18307 ( .A1(n15744), .A2(n15065), .ZN(n15067) );
  AOI21_X1 U18308 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n15744), .A(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15066) );
  AOI21_X1 U18309 ( .B1(n15752), .B2(n15067), .A(n15066), .ZN(n15068) );
  AOI211_X1 U18310 ( .C1(n20110), .C2(n15799), .A(n15069), .B(n15068), .ZN(
        n15070) );
  OAI21_X1 U18311 ( .B1(n15071), .B2(n20105), .A(n15070), .ZN(P1_U3009) );
  NOR2_X1 U18312 ( .A1(n15973), .A2(n15971), .ZN(n15073) );
  INV_X1 U18313 ( .A(n15947), .ZN(n15072) );
  OAI21_X1 U18314 ( .B1(n15074), .B2(n15073), .A(n15072), .ZN(n15080) );
  OAI21_X1 U18315 ( .B1(n15952), .B2(n15885), .A(n13248), .ZN(n15079) );
  NAND2_X1 U18316 ( .A1(n20087), .A2(n15075), .ZN(n15077) );
  OAI211_X1 U18317 ( .C1(n15817), .C2(n16014), .A(n15077), .B(n15076), .ZN(
        n15078) );
  AOI21_X1 U18318 ( .B1(n15080), .B2(n15079), .A(n15078), .ZN(n15081) );
  INV_X1 U18319 ( .A(n15081), .ZN(P1_U3011) );
  INV_X1 U18320 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15953) );
  NOR3_X1 U18321 ( .A1(n13237), .A2(n15953), .A3(n15894), .ZN(n15086) );
  INV_X1 U18322 ( .A(n15991), .ZN(n15082) );
  AOI21_X1 U18323 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n15083), .A(
        n15082), .ZN(n15084) );
  AOI221_X1 U18324 ( .B1(n15970), .B2(n20078), .C1(n15085), .C2(n20078), .A(
        n15084), .ZN(n15962) );
  OAI21_X1 U18325 ( .B1(n15142), .B2(n15086), .A(n15962), .ZN(n15958) );
  INV_X1 U18326 ( .A(n15958), .ZN(n15095) );
  NAND3_X1 U18327 ( .A1(n15087), .A2(n14902), .A3(n20087), .ZN(n15093) );
  NOR2_X1 U18328 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15088), .ZN(
        n15091) );
  OAI21_X1 U18329 ( .B1(n16014), .B2(n15833), .A(n15089), .ZN(n15090) );
  AOI21_X1 U18330 ( .B1(n15109), .B2(n15091), .A(n15090), .ZN(n15092) );
  OAI211_X1 U18331 ( .C1(n15095), .C2(n15094), .A(n15093), .B(n15092), .ZN(
        P1_U3013) );
  NAND2_X1 U18332 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15109), .ZN(
        n15954) );
  OR2_X1 U18333 ( .A1(n15954), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15968) );
  AOI21_X1 U18334 ( .B1(n15962), .B2(n15968), .A(n15894), .ZN(n15099) );
  NOR3_X1 U18335 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n13237), .A3(
        n15954), .ZN(n15098) );
  OAI21_X1 U18336 ( .B1(n16014), .B2(n15842), .A(n15096), .ZN(n15097) );
  NOR3_X1 U18337 ( .A1(n15099), .A2(n15098), .A3(n15097), .ZN(n15100) );
  OAI21_X1 U18338 ( .B1(n15101), .B2(n20105), .A(n15100), .ZN(P1_U3015) );
  INV_X1 U18339 ( .A(n15972), .ZN(n15102) );
  AOI22_X1 U18340 ( .A1(n15971), .A2(n15104), .B1(n15103), .B2(n15102), .ZN(
        n15105) );
  OAI211_X1 U18341 ( .C1(n15106), .C2(n20104), .A(n15990), .B(n15105), .ZN(
        n15974) );
  AOI21_X1 U18342 ( .B1(n15970), .B2(n15973), .A(n15974), .ZN(n15107) );
  INV_X1 U18343 ( .A(n15107), .ZN(n15108) );
  MUX2_X1 U18344 ( .A(n15109), .B(n15108), .S(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(n15113) );
  OAI21_X1 U18345 ( .B1(n16014), .B2(n15111), .A(n15110), .ZN(n15112) );
  AOI211_X1 U18346 ( .C1(n15114), .C2(n20087), .A(n15113), .B(n15112), .ZN(
        n15115) );
  INV_X1 U18347 ( .A(n15115), .ZN(P1_U3017) );
  INV_X1 U18348 ( .A(n16011), .ZN(n15116) );
  NAND2_X1 U18349 ( .A1(n15117), .A2(n20089), .ZN(n16030) );
  NOR2_X1 U18350 ( .A1(n16030), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15132) );
  INV_X1 U18351 ( .A(n15118), .ZN(n15123) );
  OAI21_X1 U18352 ( .B1(n13240), .B2(n13225), .A(n15119), .ZN(n15122) );
  INV_X1 U18353 ( .A(n15120), .ZN(n15121) );
  AOI21_X1 U18354 ( .B1(n15123), .B2(n15122), .A(n15121), .ZN(n15920) );
  NOR2_X1 U18355 ( .A1(n15125), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15981) );
  AOI21_X1 U18356 ( .B1(n20078), .B2(n15124), .A(n20095), .ZN(n16008) );
  OAI21_X1 U18357 ( .B1(n15126), .B2(n15125), .A(n20096), .ZN(n15127) );
  OAI211_X1 U18358 ( .C1(n15131), .C2(n20104), .A(n16008), .B(n15127), .ZN(
        n15984) );
  AOI21_X1 U18359 ( .B1(n15128), .B2(n15981), .A(n15984), .ZN(n15129) );
  OAI22_X1 U18360 ( .A1(n15920), .A2(n20105), .B1(n15129), .B2(n13240), .ZN(
        n15130) );
  AOI21_X1 U18361 ( .B1(n15132), .B2(n15131), .A(n15130), .ZN(n15134) );
  NAND2_X1 U18362 ( .A1(n13703), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n15133) );
  OAI211_X1 U18363 ( .C1(n16014), .C2(n15858), .A(n15134), .B(n15133), .ZN(
        P1_U3019) );
  NAND3_X1 U18364 ( .A1(n15135), .A2(n20087), .A3(n13633), .ZN(n15145) );
  AOI21_X1 U18365 ( .B1(n15137), .B2(n15136), .A(n20098), .ZN(n15138) );
  AOI211_X1 U18366 ( .C1(n20110), .C2(n15140), .A(n15139), .B(n15138), .ZN(
        n15144) );
  OR3_X1 U18367 ( .A1(n15142), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n15141), .ZN(n15143) );
  NAND3_X1 U18368 ( .A1(n15145), .A2(n15144), .A3(n15143), .ZN(P1_U3030) );
  INV_X1 U18369 ( .A(n12266), .ZN(n15155) );
  NAND3_X1 U18370 ( .A1(n15147), .A2(n15155), .A3(n15146), .ZN(n15148) );
  NAND3_X1 U18371 ( .A1(n15150), .A2(n15149), .A3(n15148), .ZN(n15742) );
  NAND2_X1 U18372 ( .A1(n12524), .A2(n15151), .ZN(n15152) );
  OAI211_X1 U18373 ( .C1(n20648), .C2(n13164), .A(n15742), .B(n15152), .ZN(
        n15153) );
  MUX2_X1 U18374 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n15153), .S(
        n20115), .Z(P1_U3478) );
  INV_X1 U18375 ( .A(n15161), .ZN(n15154) );
  NAND2_X1 U18376 ( .A1(n15155), .A2(n15154), .ZN(n15157) );
  OAI22_X1 U18377 ( .A1(n15158), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n15157), .B2(n15156), .ZN(n15159) );
  AOI21_X1 U18378 ( .B1(n20592), .B2(n15160), .A(n15159), .ZN(n15711) );
  AOI22_X1 U18379 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n20098), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13251), .ZN(n20796) );
  NAND2_X1 U18380 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20795) );
  INV_X1 U18381 ( .A(n20795), .ZN(n15163) );
  NOR3_X1 U18382 ( .A1(n12266), .A2(n15161), .A3(n20794), .ZN(n15162) );
  AOI21_X1 U18383 ( .B1(n20796), .B2(n15163), .A(n15162), .ZN(n15164) );
  OAI21_X1 U18384 ( .B1(n15711), .B2(n20790), .A(n15164), .ZN(n15165) );
  MUX2_X1 U18385 ( .A(n15165), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n20799), .Z(P1_U3473) );
  AOI21_X1 U18386 ( .B1(n15167), .B2(n15166), .A(n15324), .ZN(n15559) );
  AOI211_X1 U18387 ( .C1(n15170), .C2(n15169), .A(n15168), .B(n19732), .ZN(
        n15175) );
  AOI21_X1 U18388 ( .B1(P2_REIP_REG_18__SCAN_IN), .B2(n18993), .A(n16261), 
        .ZN(n15172) );
  AOI22_X1 U18389 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18968), .B1(
        P2_EBX_REG_18__SCAN_IN), .B2(n18978), .ZN(n15171) );
  OAI211_X1 U18390 ( .C1(n15173), .C2(n18982), .A(n15172), .B(n15171), .ZN(
        n15174) );
  AOI211_X1 U18391 ( .C1(n18979), .C2(n15559), .A(n15175), .B(n15174), .ZN(
        n15176) );
  OAI21_X1 U18392 ( .B1(n18973), .B2(n15562), .A(n15176), .ZN(P2_U2837) );
  NAND2_X1 U18393 ( .A1(n16045), .A2(n15201), .ZN(n15177) );
  OAI21_X1 U18394 ( .B1(n15201), .B2(n16050), .A(n15177), .ZN(P2_U2856) );
  NOR2_X1 U18395 ( .A1(n16059), .A2(n15259), .ZN(n15178) );
  AOI21_X1 U18396 ( .B1(P2_EBX_REG_29__SCAN_IN), .B2(n15259), .A(n15178), .ZN(
        n15179) );
  OAI21_X1 U18397 ( .B1(n15180), .B2(n15261), .A(n15179), .ZN(P2_U2858) );
  INV_X1 U18398 ( .A(n15182), .ZN(n15183) );
  NOR2_X1 U18399 ( .A1(n15181), .A2(n15183), .ZN(n15185) );
  XNOR2_X1 U18400 ( .A(n15185), .B(n15184), .ZN(n15266) );
  NOR2_X1 U18401 ( .A1(n16071), .A2(n15259), .ZN(n15186) );
  AOI21_X1 U18402 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n15259), .A(n15186), .ZN(
        n15187) );
  OAI21_X1 U18403 ( .B1(n15266), .B2(n15261), .A(n15187), .ZN(P2_U2859) );
  XNOR2_X1 U18404 ( .A(n15188), .B(n15189), .ZN(n15274) );
  NOR2_X1 U18405 ( .A1(n15200), .A2(n15190), .ZN(n15191) );
  NOR2_X1 U18406 ( .A1(n16094), .A2(n15259), .ZN(n15192) );
  AOI21_X1 U18407 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n15259), .A(n15192), .ZN(
        n15193) );
  OAI21_X1 U18408 ( .B1(n15274), .B2(n15261), .A(n15193), .ZN(P2_U2860) );
  AOI21_X1 U18409 ( .B1(n15196), .B2(n15195), .A(n15194), .ZN(n15197) );
  INV_X1 U18410 ( .A(n15197), .ZN(n15281) );
  NAND2_X1 U18411 ( .A1(n15259), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n15203) );
  AND2_X1 U18412 ( .A1(n15208), .A2(n15198), .ZN(n15199) );
  NOR2_X1 U18413 ( .A1(n15200), .A2(n15199), .ZN(n16101) );
  NAND2_X1 U18414 ( .A1(n16101), .A2(n15201), .ZN(n15202) );
  OAI211_X1 U18415 ( .C1(n15281), .C2(n15261), .A(n15203), .B(n15202), .ZN(
        P2_U2861) );
  XNOR2_X1 U18416 ( .A(n15204), .B(n15205), .ZN(n15291) );
  NAND2_X1 U18417 ( .A1(n15214), .A2(n15206), .ZN(n15207) );
  NAND2_X1 U18418 ( .A1(n15208), .A2(n15207), .ZN(n16115) );
  MUX2_X1 U18419 ( .A(n16115), .B(n15209), .S(n15259), .Z(n15210) );
  OAI21_X1 U18420 ( .B1(n15291), .B2(n15261), .A(n15210), .ZN(P2_U2862) );
  NAND2_X1 U18421 ( .A1(n15212), .A2(n15211), .ZN(n15213) );
  NAND2_X1 U18422 ( .A1(n15214), .A2(n15213), .ZN(n16124) );
  NOR2_X1 U18423 ( .A1(n15216), .A2(n19169), .ZN(n15217) );
  XNOR2_X1 U18424 ( .A(n15218), .B(n15217), .ZN(n15219) );
  XNOR2_X1 U18425 ( .A(n15215), .B(n15219), .ZN(n16139) );
  NAND2_X1 U18426 ( .A1(n16139), .A2(n15247), .ZN(n15221) );
  NAND2_X1 U18427 ( .A1(n15259), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n15220) );
  OAI211_X1 U18428 ( .C1(n16124), .C2(n15259), .A(n15221), .B(n15220), .ZN(
        P2_U2863) );
  OAI21_X1 U18429 ( .B1(n15224), .B2(n15223), .A(n15222), .ZN(n15296) );
  NOR2_X1 U18430 ( .A1(n15495), .A2(n15259), .ZN(n15225) );
  AOI21_X1 U18431 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n15259), .A(n15225), .ZN(
        n15226) );
  OAI21_X1 U18432 ( .B1(n15296), .B2(n15261), .A(n15226), .ZN(P2_U2864) );
  AND2_X1 U18433 ( .A1(n15228), .A2(n15227), .ZN(n15230) );
  OR2_X1 U18434 ( .A1(n15230), .A2(n15229), .ZN(n15697) );
  AOI21_X1 U18435 ( .B1(n15233), .B2(n15231), .A(n15232), .ZN(n15297) );
  NAND2_X1 U18436 ( .A1(n15297), .A2(n15247), .ZN(n15235) );
  NAND2_X1 U18437 ( .A1(n15259), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n15234) );
  OAI211_X1 U18438 ( .C1(n15697), .C2(n15259), .A(n15235), .B(n15234), .ZN(
        P2_U2865) );
  OAI21_X1 U18439 ( .B1(n15236), .B2(n15237), .A(n15231), .ZN(n15314) );
  MUX2_X1 U18440 ( .A(n15239), .B(n15238), .S(n15259), .Z(n15240) );
  OAI21_X1 U18441 ( .B1(n15314), .B2(n15261), .A(n15240), .ZN(P2_U2866) );
  INV_X1 U18442 ( .A(n15241), .ZN(n15257) );
  INV_X1 U18443 ( .A(n15242), .ZN(n15243) );
  NAND2_X1 U18444 ( .A1(n15257), .A2(n15243), .ZN(n15244) );
  NAND2_X1 U18445 ( .A1(n9907), .A2(n15244), .ZN(n18843) );
  OR2_X1 U18446 ( .A1(n14208), .A2(n15245), .ZN(n15250) );
  AOI21_X1 U18447 ( .B1(n15246), .B2(n15250), .A(n15236), .ZN(n15315) );
  NAND2_X1 U18448 ( .A1(n15315), .A2(n15247), .ZN(n15249) );
  NAND2_X1 U18449 ( .A1(n15259), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n15248) );
  OAI211_X1 U18450 ( .C1(n18843), .C2(n15259), .A(n15249), .B(n15248), .ZN(
        P2_U2867) );
  OAI21_X1 U18451 ( .B1(n15252), .B2(n15251), .A(n15250), .ZN(n15332) );
  INV_X1 U18452 ( .A(n15253), .ZN(n15255) );
  NAND2_X1 U18453 ( .A1(n15255), .A2(n15254), .ZN(n15256) );
  NAND2_X1 U18454 ( .A1(n15257), .A2(n15256), .ZN(n18860) );
  NOR2_X1 U18455 ( .A1(n15259), .A2(n18860), .ZN(n15258) );
  AOI21_X1 U18456 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n15259), .A(n15258), .ZN(
        n15260) );
  OAI21_X1 U18457 ( .B1(n15332), .B2(n15261), .A(n15260), .ZN(P2_U2868) );
  INV_X1 U18458 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n19072) );
  OAI22_X1 U18459 ( .A1(n16134), .A2(n15262), .B1(n15340), .B2(n19072), .ZN(
        n15263) );
  AOI21_X1 U18460 ( .B1(n19051), .B2(n16072), .A(n15263), .ZN(n15265) );
  AOI22_X1 U18461 ( .A1(n18999), .A2(BUF2_REG_28__SCAN_IN), .B1(n18998), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n15264) );
  OAI211_X1 U18462 ( .C1(n15266), .C2(n16136), .A(n15265), .B(n15264), .ZN(
        P2_U2891) );
  INV_X1 U18463 ( .A(n15267), .ZN(n15269) );
  INV_X1 U18464 ( .A(n15275), .ZN(n15268) );
  AOI21_X1 U18465 ( .B1(n15269), .B2(n15268), .A(n14504), .ZN(n16097) );
  INV_X1 U18466 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n19074) );
  OAI22_X1 U18467 ( .A1(n16134), .A2(n15270), .B1(n15340), .B2(n19074), .ZN(
        n15271) );
  AOI21_X1 U18468 ( .B1(n19051), .B2(n16097), .A(n15271), .ZN(n15273) );
  AOI22_X1 U18469 ( .A1(n18999), .A2(BUF2_REG_27__SCAN_IN), .B1(n18998), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n15272) );
  OAI211_X1 U18470 ( .C1(n15274), .C2(n16136), .A(n15273), .B(n15272), .ZN(
        P2_U2892) );
  AOI21_X1 U18471 ( .B1(n15276), .B2(n15285), .A(n15275), .ZN(n16100) );
  INV_X1 U18472 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n19076) );
  OAI22_X1 U18473 ( .A1(n16134), .A2(n15277), .B1(n15340), .B2(n19076), .ZN(
        n15278) );
  AOI21_X1 U18474 ( .B1(n19051), .B2(n16100), .A(n15278), .ZN(n15280) );
  AOI22_X1 U18475 ( .A1(n18999), .A2(BUF2_REG_26__SCAN_IN), .B1(n18998), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n15279) );
  OAI211_X1 U18476 ( .C1(n15281), .C2(n16136), .A(n15280), .B(n15279), .ZN(
        P2_U2893) );
  INV_X1 U18477 ( .A(n15282), .ZN(n15284) );
  INV_X1 U18478 ( .A(n15283), .ZN(n15486) );
  NAND2_X1 U18479 ( .A1(n15284), .A2(n15486), .ZN(n15286) );
  AND2_X1 U18480 ( .A1(n15286), .A2(n15285), .ZN(n16121) );
  INV_X1 U18481 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n19078) );
  OAI22_X1 U18482 ( .A1(n16134), .A2(n15287), .B1(n15340), .B2(n19078), .ZN(
        n15288) );
  AOI21_X1 U18483 ( .B1(n19051), .B2(n16121), .A(n15288), .ZN(n15290) );
  AOI22_X1 U18484 ( .A1(n18999), .A2(BUF2_REG_25__SCAN_IN), .B1(n18998), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n15289) );
  OAI211_X1 U18485 ( .C1(n15291), .C2(n16136), .A(n15290), .B(n15289), .ZN(
        P2_U2894) );
  INV_X1 U18486 ( .A(n15499), .ZN(n15293) );
  INV_X1 U18487 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n19082) );
  OAI22_X1 U18488 ( .A1(n16134), .A2(n19201), .B1(n15340), .B2(n19082), .ZN(
        n15292) );
  AOI21_X1 U18489 ( .B1(n19051), .B2(n15293), .A(n15292), .ZN(n15295) );
  AOI22_X1 U18490 ( .A1(n18999), .A2(BUF2_REG_23__SCAN_IN), .B1(n18998), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n15294) );
  OAI211_X1 U18491 ( .C1(n15296), .C2(n16136), .A(n15295), .B(n15294), .ZN(
        P2_U2896) );
  INV_X1 U18492 ( .A(n15297), .ZN(n15307) );
  NOR2_X1 U18493 ( .A1(n15299), .A2(n15298), .ZN(n15300) );
  NOR2_X1 U18494 ( .A1(n15301), .A2(n15300), .ZN(n15698) );
  INV_X1 U18495 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n19084) );
  OAI22_X1 U18496 ( .A1(n16134), .A2(n19191), .B1(n19033), .B2(n19084), .ZN(
        n15305) );
  INV_X1 U18497 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n15303) );
  INV_X1 U18498 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n15302) );
  OAI22_X1 U18499 ( .A1(n15344), .A2(n15303), .B1(n15342), .B2(n15302), .ZN(
        n15304) );
  AOI211_X1 U18500 ( .C1(n19051), .C2(n15698), .A(n15305), .B(n15304), .ZN(
        n15306) );
  OAI21_X1 U18501 ( .B1(n15307), .B2(n16136), .A(n15306), .ZN(P2_U2897) );
  INV_X1 U18502 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n19086) );
  OAI22_X1 U18503 ( .A1(n16134), .A2(n19188), .B1(n19033), .B2(n19086), .ZN(
        n15311) );
  INV_X1 U18504 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n15309) );
  OAI22_X1 U18505 ( .A1(n15344), .A2(n15309), .B1(n15342), .B2(n15308), .ZN(
        n15310) );
  AOI211_X1 U18506 ( .C1(n19051), .C2(n15312), .A(n15311), .B(n15310), .ZN(
        n15313) );
  OAI21_X1 U18507 ( .B1(n15314), .B2(n16136), .A(n15313), .ZN(P2_U2898) );
  INV_X1 U18508 ( .A(n15315), .ZN(n15323) );
  AOI21_X1 U18509 ( .B1(n15317), .B2(n9914), .A(n15316), .ZN(n18844) );
  INV_X1 U18510 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n19089) );
  OAI22_X1 U18511 ( .A1(n16134), .A2(n19185), .B1(n19033), .B2(n19089), .ZN(
        n15321) );
  INV_X1 U18512 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n15319) );
  INV_X1 U18513 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n15318) );
  OAI22_X1 U18514 ( .A1(n15344), .A2(n15319), .B1(n15342), .B2(n15318), .ZN(
        n15320) );
  AOI211_X1 U18515 ( .C1(n19051), .C2(n18844), .A(n15321), .B(n15320), .ZN(
        n15322) );
  OAI21_X1 U18516 ( .B1(n15323), .B2(n16136), .A(n15322), .ZN(P2_U2899) );
  OAI21_X1 U18517 ( .B1(n15325), .B2(n15324), .A(n9914), .ZN(n18859) );
  INV_X1 U18518 ( .A(n18859), .ZN(n15330) );
  INV_X1 U18519 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n19091) );
  OAI22_X1 U18520 ( .A1(n16134), .A2(n19181), .B1(n15340), .B2(n19091), .ZN(
        n15329) );
  INV_X1 U18521 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n15327) );
  INV_X1 U18522 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n15326) );
  OAI22_X1 U18523 ( .A1(n15344), .A2(n15327), .B1(n15342), .B2(n15326), .ZN(
        n15328) );
  AOI211_X1 U18524 ( .C1(n19051), .C2(n15330), .A(n15329), .B(n15328), .ZN(
        n15331) );
  OAI21_X1 U18525 ( .B1(n15332), .B2(n16136), .A(n15331), .ZN(P2_U2900) );
  INV_X1 U18526 ( .A(n15333), .ZN(n15339) );
  INV_X1 U18527 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n19093) );
  OAI22_X1 U18528 ( .A1(n16134), .A2(n19175), .B1(n15340), .B2(n19093), .ZN(
        n15337) );
  INV_X1 U18529 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n15335) );
  INV_X1 U18530 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n15334) );
  OAI22_X1 U18531 ( .A1(n15344), .A2(n15335), .B1(n15342), .B2(n15334), .ZN(
        n15336) );
  AOI211_X1 U18532 ( .C1(n19051), .C2(n15559), .A(n15337), .B(n15336), .ZN(
        n15338) );
  OAI21_X1 U18533 ( .B1(n15339), .B2(n16136), .A(n15338), .ZN(P2_U2901) );
  INV_X1 U18534 ( .A(n15579), .ZN(n15347) );
  INV_X1 U18535 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n19096) );
  OAI22_X1 U18536 ( .A1(n16134), .A2(n19170), .B1(n15340), .B2(n19096), .ZN(
        n15346) );
  INV_X1 U18537 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n15343) );
  INV_X1 U18538 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n15341) );
  OAI22_X1 U18539 ( .A1(n15344), .A2(n15343), .B1(n15342), .B2(n15341), .ZN(
        n15345) );
  AOI211_X1 U18540 ( .C1(n19051), .C2(n15347), .A(n15346), .B(n15345), .ZN(
        n15348) );
  OAI21_X1 U18541 ( .B1(n15349), .B2(n16136), .A(n15348), .ZN(P2_U2902) );
  OAI21_X1 U18542 ( .B1(n15350), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n11890), .ZN(n15455) );
  NAND3_X1 U18543 ( .A1(n15446), .A2(n10996), .A3(n15352), .ZN(n15356) );
  NOR2_X1 U18544 ( .A1(n19790), .A2(n18878), .ZN(n15449) );
  AOI21_X1 U18545 ( .B1(n19137), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15449), .ZN(n15353) );
  OAI21_X1 U18546 ( .B1(n16094), .B2(n19157), .A(n15353), .ZN(n15354) );
  AOI21_X1 U18547 ( .B1(n16084), .B2(n16234), .A(n15354), .ZN(n15355) );
  OAI211_X1 U18548 ( .C1(n19140), .C2(n15455), .A(n15356), .B(n15355), .ZN(
        P2_U2987) );
  NAND2_X1 U18549 ( .A1(n9899), .A2(n15366), .ZN(n15358) );
  MUX2_X1 U18550 ( .A(n15358), .B(n15366), .S(n15357), .Z(n15359) );
  NAND2_X1 U18551 ( .A1(n15359), .A2(n11873), .ZN(n15468) );
  INV_X1 U18552 ( .A(n15360), .ZN(n15470) );
  AOI21_X1 U18553 ( .B1(n15464), .B2(n15470), .A(n15350), .ZN(n15466) );
  AND2_X1 U18554 ( .A1(P2_REIP_REG_26__SCAN_IN), .A2(n16261), .ZN(n15461) );
  AOI21_X1 U18555 ( .B1(n19137), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15461), .ZN(n15362) );
  NAND2_X1 U18556 ( .A1(n16101), .A2(n19146), .ZN(n15361) );
  OAI211_X1 U18557 ( .C1(n15363), .C2(n19150), .A(n15362), .B(n15361), .ZN(
        n15364) );
  AOI21_X1 U18558 ( .B1(n15466), .B2(n16228), .A(n15364), .ZN(n15365) );
  OAI21_X1 U18559 ( .B1(n19142), .B2(n15468), .A(n15365), .ZN(P2_U2988) );
  INV_X1 U18560 ( .A(n15366), .ZN(n15367) );
  NOR2_X1 U18561 ( .A1(n15368), .A2(n15367), .ZN(n15370) );
  XOR2_X1 U18562 ( .A(n15370), .B(n15369), .Z(n15479) );
  NAND2_X1 U18563 ( .A1(n15371), .A2(n15459), .ZN(n15469) );
  NAND3_X1 U18564 ( .A1(n15470), .A2(n16228), .A3(n15469), .ZN(n15375) );
  NOR2_X1 U18565 ( .A1(n19786), .A2(n18878), .ZN(n15473) );
  AOI21_X1 U18566 ( .B1(n19137), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n15473), .ZN(n15372) );
  OAI21_X1 U18567 ( .B1(n16115), .B2(n19157), .A(n15372), .ZN(n15373) );
  AOI21_X1 U18568 ( .B1(n16112), .B2(n16234), .A(n15373), .ZN(n15374) );
  OAI211_X1 U18569 ( .C1(n19142), .C2(n15479), .A(n15375), .B(n15374), .ZN(
        P2_U2989) );
  INV_X1 U18570 ( .A(n15376), .ZN(n15377) );
  OAI21_X1 U18571 ( .B1(n15377), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15371), .ZN(n15492) );
  XNOR2_X1 U18572 ( .A(n15379), .B(n15482), .ZN(n15380) );
  XNOR2_X1 U18573 ( .A(n15378), .B(n15380), .ZN(n15490) );
  OAI22_X1 U18574 ( .A1(n11461), .A2(n18878), .B1(n19150), .B2(n15381), .ZN(
        n15384) );
  INV_X1 U18575 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15382) );
  OAI22_X1 U18576 ( .A1(n16124), .A2(n19157), .B1(n15382), .B2(n16243), .ZN(
        n15383) );
  AOI211_X1 U18577 ( .C1(n15490), .C2(n10996), .A(n15384), .B(n15383), .ZN(
        n15385) );
  OAI21_X1 U18578 ( .B1(n15492), .B2(n19140), .A(n15385), .ZN(P2_U2990) );
  OAI21_X1 U18579 ( .B1(n15386), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15376), .ZN(n15505) );
  AND2_X1 U18580 ( .A1(n15387), .A2(n15396), .ZN(n15388) );
  XOR2_X1 U18581 ( .A(n15389), .B(n15388), .Z(n15502) );
  NOR2_X1 U18582 ( .A1(n15390), .A2(n19150), .ZN(n15393) );
  NAND2_X1 U18583 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n16261), .ZN(n15498) );
  NAND2_X1 U18584 ( .A1(n19137), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15391) );
  OAI211_X1 U18585 ( .C1(n15495), .C2(n19157), .A(n15498), .B(n15391), .ZN(
        n15392) );
  AOI211_X1 U18586 ( .C1(n15502), .C2(n10996), .A(n15393), .B(n15392), .ZN(
        n15394) );
  OAI21_X1 U18587 ( .B1(n19140), .B2(n15505), .A(n15394), .ZN(P2_U2991) );
  NAND2_X1 U18588 ( .A1(n15396), .A2(n15395), .ZN(n15400) );
  NAND2_X1 U18589 ( .A1(n15398), .A2(n15397), .ZN(n15399) );
  XOR2_X1 U18590 ( .A(n15400), .B(n15399), .Z(n15516) );
  INV_X1 U18591 ( .A(n15386), .ZN(n15507) );
  NAND2_X1 U18592 ( .A1(n11817), .A2(n15509), .ZN(n15506) );
  NAND3_X1 U18593 ( .A1(n15507), .A2(n16228), .A3(n15506), .ZN(n15405) );
  NOR2_X1 U18594 ( .A1(n15697), .A2(n19157), .ZN(n15403) );
  INV_X1 U18595 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n19781) );
  OAI22_X1 U18596 ( .A1(n19781), .A2(n18878), .B1(n19150), .B2(n15401), .ZN(
        n15402) );
  AOI211_X1 U18597 ( .C1(n19137), .C2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15403), .B(n15402), .ZN(n15404) );
  OAI211_X1 U18598 ( .C1(n15516), .C2(n19142), .A(n15405), .B(n15404), .ZN(
        P2_U2992) );
  OR2_X1 U18599 ( .A1(n15406), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15407) );
  NAND2_X1 U18600 ( .A1(n11816), .A2(n15407), .ZN(n15529) );
  AOI21_X1 U18601 ( .B1(n15410), .B2(n15409), .A(n15408), .ZN(n15517) );
  NAND2_X1 U18602 ( .A1(n15517), .A2(n10996), .ZN(n15415) );
  NOR2_X1 U18603 ( .A1(n18843), .A2(n19157), .ZN(n15413) );
  NAND2_X1 U18604 ( .A1(P2_REIP_REG_20__SCAN_IN), .A2(n19138), .ZN(n15522) );
  OAI21_X1 U18605 ( .B1(n19150), .B2(n15411), .A(n15522), .ZN(n15412) );
  AOI211_X1 U18606 ( .C1(n19137), .C2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15413), .B(n15412), .ZN(n15414) );
  OAI211_X1 U18607 ( .C1(n19140), .C2(n15529), .A(n15415), .B(n15414), .ZN(
        P2_U2994) );
  AOI21_X1 U18608 ( .B1(n15418), .B2(n15417), .A(n15416), .ZN(n15582) );
  NOR2_X1 U18609 ( .A1(n15567), .A2(n19157), .ZN(n15421) );
  NAND2_X1 U18610 ( .A1(P2_REIP_REG_17__SCAN_IN), .A2(n19138), .ZN(n15578) );
  OAI21_X1 U18611 ( .B1(n16243), .B2(n15419), .A(n15578), .ZN(n15420) );
  AOI211_X1 U18612 ( .C1(n16234), .C2(n15422), .A(n15421), .B(n15420), .ZN(
        n15426) );
  OAI211_X1 U18613 ( .C1(n15571), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n16228), .B(n15424), .ZN(n15425) );
  OAI211_X1 U18614 ( .C1(n15582), .C2(n19142), .A(n15426), .B(n15425), .ZN(
        P2_U2997) );
  OAI21_X1 U18615 ( .B1(n15429), .B2(n15428), .A(n15427), .ZN(n15691) );
  NAND2_X1 U18616 ( .A1(P2_REIP_REG_16__SCAN_IN), .A2(n16261), .ZN(n15689) );
  NAND2_X1 U18617 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n19137), .ZN(
        n15430) );
  OAI211_X1 U18618 ( .C1(n19150), .C2(n18867), .A(n15689), .B(n15430), .ZN(
        n15432) );
  AOI211_X1 U18619 ( .C1(n15695), .C2(n15589), .A(n19140), .B(n15571), .ZN(
        n15431) );
  AOI211_X1 U18620 ( .C1(n19146), .C2(n18874), .A(n15432), .B(n15431), .ZN(
        n15433) );
  OAI21_X1 U18621 ( .B1(n15691), .B2(n19142), .A(n15433), .ZN(P2_U2998) );
  NOR2_X1 U18622 ( .A1(n16059), .A2(n16272), .ZN(n15441) );
  INV_X1 U18623 ( .A(n16058), .ZN(n15439) );
  INV_X1 U18624 ( .A(n15447), .ZN(n15435) );
  OAI211_X1 U18625 ( .C1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15436), .A(
        n15435), .B(n15434), .ZN(n15438) );
  OAI211_X1 U18626 ( .C1(n16271), .C2(n15439), .A(n15438), .B(n15437), .ZN(
        n15440) );
  AOI211_X1 U18627 ( .C1(n15452), .C2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15441), .B(n15440), .ZN(n15444) );
  NAND2_X1 U18628 ( .A1(n15442), .A2(n11843), .ZN(n15443) );
  OAI211_X1 U18629 ( .C1(n15445), .C2(n16278), .A(n15444), .B(n15443), .ZN(
        P2_U3017) );
  NAND3_X1 U18630 ( .A1(n15446), .A2(n15352), .A3(n16283), .ZN(n15454) );
  NOR2_X1 U18631 ( .A1(n15447), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15448) );
  AOI211_X1 U18632 ( .C1(n16280), .C2(n16097), .A(n15449), .B(n15448), .ZN(
        n15450) );
  OAI21_X1 U18633 ( .B1(n16094), .B2(n16272), .A(n15450), .ZN(n15451) );
  AOI21_X1 U18634 ( .B1(n15452), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15451), .ZN(n15453) );
  OAI211_X1 U18635 ( .C1(n15455), .C2(n15637), .A(n15454), .B(n15453), .ZN(
        P2_U3019) );
  INV_X1 U18636 ( .A(n15481), .ZN(n15456) );
  AOI21_X1 U18637 ( .B1(n15457), .B2(n15482), .A(n15456), .ZN(n15471) );
  AOI21_X1 U18638 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15464), .A(
        n15459), .ZN(n15458) );
  AOI211_X1 U18639 ( .C1(n15464), .C2(n15459), .A(n15483), .B(n15458), .ZN(
        n15460) );
  AOI211_X1 U18640 ( .C1(n16280), .C2(n16100), .A(n15461), .B(n15460), .ZN(
        n15463) );
  NAND2_X1 U18641 ( .A1(n16101), .A2(n16285), .ZN(n15462) );
  OAI211_X1 U18642 ( .C1(n15471), .C2(n15464), .A(n15463), .B(n15462), .ZN(
        n15465) );
  AOI21_X1 U18643 ( .B1(n15466), .B2(n11843), .A(n15465), .ZN(n15467) );
  OAI21_X1 U18644 ( .B1(n16278), .B2(n15468), .A(n15467), .ZN(P2_U3020) );
  NAND3_X1 U18645 ( .A1(n15470), .A2(n11843), .A3(n15469), .ZN(n15478) );
  INV_X1 U18646 ( .A(n15471), .ZN(n15476) );
  NOR3_X1 U18647 ( .A1(n15483), .A2(n15482), .A3(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15472) );
  AOI211_X1 U18648 ( .C1(n16280), .C2(n16121), .A(n15473), .B(n15472), .ZN(
        n15474) );
  OAI21_X1 U18649 ( .B1(n16115), .B2(n16272), .A(n15474), .ZN(n15475) );
  AOI21_X1 U18650 ( .B1(n15476), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15475), .ZN(n15477) );
  OAI211_X1 U18651 ( .C1(n15479), .C2(n16278), .A(n15478), .B(n15477), .ZN(
        P2_U3021) );
  NAND2_X1 U18652 ( .A1(P2_REIP_REG_24__SCAN_IN), .A2(n16261), .ZN(n15480) );
  OAI221_X1 U18653 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15483), 
        .C1(n15482), .C2(n15481), .A(n15480), .ZN(n15489) );
  NAND2_X1 U18654 ( .A1(n15485), .A2(n15484), .ZN(n15487) );
  NAND2_X1 U18655 ( .A1(n15487), .A2(n15486), .ZN(n16137) );
  OAI22_X1 U18656 ( .A1(n16124), .A2(n16272), .B1(n16271), .B2(n16137), .ZN(
        n15488) );
  AOI211_X1 U18657 ( .C1(n15490), .C2(n16283), .A(n15489), .B(n15488), .ZN(
        n15491) );
  OAI21_X1 U18658 ( .B1(n15492), .B2(n15637), .A(n15491), .ZN(P2_U3022) );
  AOI21_X1 U18659 ( .B1(n15494), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15493), .ZN(n15513) );
  NOR2_X1 U18660 ( .A1(n15495), .A2(n16272), .ZN(n15501) );
  XNOR2_X1 U18661 ( .A(n15509), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15496) );
  NAND2_X1 U18662 ( .A1(n15496), .A2(n15508), .ZN(n15497) );
  OAI211_X1 U18663 ( .C1(n16271), .C2(n15499), .A(n15498), .B(n15497), .ZN(
        n15500) );
  AOI211_X1 U18664 ( .C1(n15513), .C2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15501), .B(n15500), .ZN(n15504) );
  NAND2_X1 U18665 ( .A1(n15502), .A2(n16283), .ZN(n15503) );
  OAI211_X1 U18666 ( .C1(n15505), .C2(n15637), .A(n15504), .B(n15503), .ZN(
        P2_U3023) );
  NAND3_X1 U18667 ( .A1(n15507), .A2(n11843), .A3(n15506), .ZN(n15515) );
  AOI22_X1 U18668 ( .A1(n15509), .A2(n15508), .B1(n19138), .B2(
        P2_REIP_REG_22__SCAN_IN), .ZN(n15511) );
  NAND2_X1 U18669 ( .A1(n16280), .A2(n15698), .ZN(n15510) );
  OAI211_X1 U18670 ( .C1(n15697), .C2(n16272), .A(n15511), .B(n15510), .ZN(
        n15512) );
  AOI21_X1 U18671 ( .B1(n15513), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15512), .ZN(n15514) );
  OAI211_X1 U18672 ( .C1(n15516), .C2(n16278), .A(n15515), .B(n15514), .ZN(
        P2_U3024) );
  NAND2_X1 U18673 ( .A1(n15517), .A2(n16283), .ZN(n15528) );
  AND2_X1 U18674 ( .A1(n15604), .A2(n15518), .ZN(n15519) );
  OR2_X1 U18675 ( .A1(n16258), .A2(n15519), .ZN(n15558) );
  INV_X1 U18676 ( .A(n15558), .ZN(n15541) );
  OAI211_X1 U18677 ( .C1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(n15544), .B(n15520), .ZN(
        n15521) );
  OAI211_X1 U18678 ( .C1(n15541), .C2(n15523), .A(n15522), .B(n15521), .ZN(
        n15526) );
  NAND2_X1 U18679 ( .A1(n16280), .A2(n18844), .ZN(n15524) );
  OAI21_X1 U18680 ( .B1(n18843), .B2(n16272), .A(n15524), .ZN(n15525) );
  NOR2_X1 U18681 ( .A1(n15526), .A2(n15525), .ZN(n15527) );
  OAI211_X1 U18682 ( .C1(n15529), .C2(n15637), .A(n15528), .B(n15527), .ZN(
        P2_U3026) );
  AOI21_X1 U18683 ( .B1(n15543), .B2(n15531), .A(n15406), .ZN(n16144) );
  INV_X1 U18684 ( .A(n16144), .ZN(n15547) );
  INV_X1 U18685 ( .A(n15532), .ZN(n15534) );
  NAND2_X1 U18686 ( .A1(n15534), .A2(n15533), .ZN(n15536) );
  XNOR2_X1 U18687 ( .A(n15536), .B(n15535), .ZN(n16145) );
  NAND2_X1 U18688 ( .A1(n16145), .A2(n16283), .ZN(n15546) );
  INV_X1 U18689 ( .A(n18860), .ZN(n15539) );
  NOR2_X1 U18690 ( .A1(n19776), .A2(n18878), .ZN(n15538) );
  NOR2_X1 U18691 ( .A1(n16271), .A2(n18859), .ZN(n15537) );
  AOI211_X1 U18692 ( .C1(n16285), .C2(n15539), .A(n15538), .B(n15537), .ZN(
        n15540) );
  OAI21_X1 U18693 ( .B1(n15541), .B2(n15543), .A(n15540), .ZN(n15542) );
  AOI21_X1 U18694 ( .B1(n15544), .B2(n15543), .A(n15542), .ZN(n15545) );
  OAI211_X1 U18695 ( .C1(n15547), .C2(n15637), .A(n15546), .B(n15545), .ZN(
        P2_U3027) );
  NAND2_X1 U18696 ( .A1(n15424), .A2(n15556), .ZN(n15548) );
  NAND2_X1 U18697 ( .A1(n15531), .A2(n15548), .ZN(n16148) );
  INV_X1 U18698 ( .A(n15549), .ZN(n15550) );
  NAND2_X1 U18699 ( .A1(n15551), .A2(n15550), .ZN(n15552) );
  XNOR2_X1 U18700 ( .A(n15553), .B(n15552), .ZN(n16149) );
  OR2_X1 U18701 ( .A1(n16149), .A2(n16278), .ZN(n15566) );
  NOR2_X1 U18702 ( .A1(n15555), .A2(n15554), .ZN(n15609) );
  AND2_X1 U18703 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15609), .ZN(
        n15591) );
  AND2_X1 U18704 ( .A1(n15557), .A2(n15556), .ZN(n15564) );
  NAND2_X1 U18705 ( .A1(n15558), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15561) );
  AOI22_X1 U18706 ( .A1(n16280), .A2(n15559), .B1(n16261), .B2(
        P2_REIP_REG_18__SCAN_IN), .ZN(n15560) );
  OAI211_X1 U18707 ( .C1(n16272), .C2(n15562), .A(n15561), .B(n15560), .ZN(
        n15563) );
  AOI21_X1 U18708 ( .B1(n15591), .B2(n15564), .A(n15563), .ZN(n15565) );
  OAI211_X1 U18709 ( .C1(n16148), .C2(n15637), .A(n15566), .B(n15565), .ZN(
        P2_U3028) );
  INV_X1 U18710 ( .A(n15567), .ZN(n15580) );
  INV_X1 U18711 ( .A(n15568), .ZN(n15569) );
  OR2_X1 U18712 ( .A1(n16258), .A2(n15569), .ZN(n15570) );
  AND2_X1 U18713 ( .A1(n15570), .A2(n16256), .ZN(n15592) );
  AOI21_X1 U18714 ( .B1(n15637), .B2(n15572), .A(n15571), .ZN(n15573) );
  AOI211_X1 U18715 ( .C1(n11034), .C2(n15574), .A(n15592), .B(n15573), .ZN(
        n15694) );
  INV_X1 U18716 ( .A(n15589), .ZN(n15576) );
  AOI22_X1 U18717 ( .A1(n15576), .A2(n11843), .B1(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15591), .ZN(n15696) );
  OAI21_X1 U18718 ( .B1(n15696), .B2(n15695), .A(n11084), .ZN(n15577) );
  OAI21_X1 U18719 ( .B1(n15582), .B2(n16278), .A(n15581), .ZN(P2_U3029) );
  NAND2_X1 U18720 ( .A1(n15583), .A2(n15600), .ZN(n15587) );
  NAND2_X1 U18721 ( .A1(n15585), .A2(n15584), .ZN(n15586) );
  XOR2_X1 U18722 ( .A(n15587), .B(n15586), .Z(n16159) );
  NAND2_X1 U18723 ( .A1(n15423), .A2(n11034), .ZN(n15588) );
  AND2_X1 U18724 ( .A1(n15589), .A2(n15588), .ZN(n16157) );
  NOR2_X1 U18725 ( .A1(n11437), .A2(n18878), .ZN(n15590) );
  AOI221_X1 U18726 ( .B1(n15592), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), 
        .C1(n15591), .C2(n11034), .A(n15590), .ZN(n15594) );
  NAND2_X1 U18727 ( .A1(n16285), .A2(n16156), .ZN(n15593) );
  OAI211_X1 U18728 ( .C1(n16271), .C2(n15595), .A(n15594), .B(n15593), .ZN(
        n15596) );
  AOI21_X1 U18729 ( .B1(n16157), .B2(n11843), .A(n15596), .ZN(n15597) );
  OAI21_X1 U18730 ( .B1(n16159), .B2(n16278), .A(n15597), .ZN(P2_U3031) );
  NOR2_X1 U18731 ( .A1(n16176), .A2(n11074), .ZN(n15606) );
  OAI21_X1 U18732 ( .B1(n15621), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n15423), .ZN(n16164) );
  NAND2_X1 U18733 ( .A1(n15600), .A2(n15599), .ZN(n15602) );
  XOR2_X1 U18734 ( .A(n15602), .B(n15601), .Z(n16165) );
  NAND2_X1 U18735 ( .A1(n15603), .A2(n16254), .ZN(n16246) );
  AOI21_X1 U18736 ( .B1(n15605), .B2(n15604), .A(n16258), .ZN(n16245) );
  OAI21_X1 U18737 ( .B1(n15606), .B2(n16246), .A(n16245), .ZN(n15626) );
  NOR2_X1 U18738 ( .A1(n11400), .A2(n18878), .ZN(n15607) );
  AOI221_X1 U18739 ( .B1(n15609), .B2(n15608), .C1(n15626), .C2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(n15607), .ZN(n15614) );
  XNOR2_X1 U18740 ( .A(n15611), .B(n15610), .ZN(n19004) );
  INV_X1 U18741 ( .A(n19004), .ZN(n15612) );
  AOI22_X1 U18742 ( .A1(n18885), .A2(n16285), .B1(n16280), .B2(n15612), .ZN(
        n15613) );
  OAI211_X1 U18743 ( .C1(n16165), .C2(n16278), .A(n15614), .B(n15613), .ZN(
        n15615) );
  INV_X1 U18744 ( .A(n15615), .ZN(n15616) );
  OAI21_X1 U18745 ( .B1(n15637), .B2(n16164), .A(n15616), .ZN(P2_U3032) );
  NOR2_X1 U18746 ( .A1(n15619), .A2(n15618), .ZN(n15620) );
  XNOR2_X1 U18747 ( .A(n15617), .B(n15620), .ZN(n16169) );
  NAND2_X1 U18748 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n16195), .ZN(
        n16174) );
  AOI21_X1 U18749 ( .B1(n11074), .B2(n16174), .A(n15621), .ZN(n16171) );
  NAND2_X1 U18750 ( .A1(n16171), .A2(n11843), .ZN(n15628) );
  OAI21_X1 U18751 ( .B1(n16176), .B2(n16246), .A(n11074), .ZN(n15625) );
  INV_X1 U18752 ( .A(n18895), .ZN(n15622) );
  AOI22_X1 U18753 ( .A1(n16280), .A2(n15622), .B1(n16261), .B2(
        P2_REIP_REG_13__SCAN_IN), .ZN(n15623) );
  OAI21_X1 U18754 ( .B1(n18896), .B2(n16272), .A(n15623), .ZN(n15624) );
  AOI21_X1 U18755 ( .B1(n15626), .B2(n15625), .A(n15624), .ZN(n15627) );
  OAI211_X1 U18756 ( .C1(n16169), .C2(n16278), .A(n15628), .B(n15627), .ZN(
        P2_U3033) );
  AOI21_X1 U18757 ( .B1(n15631), .B2(n16200), .A(n15630), .ZN(n15632) );
  AOI21_X1 U18758 ( .B1(n15629), .B2(n16200), .A(n15632), .ZN(n16216) );
  NOR2_X1 U18759 ( .A1(n11312), .A2(n18878), .ZN(n15633) );
  AOI221_X1 U18760 ( .B1(n16254), .B2(n16257), .C1(n16258), .C2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n15633), .ZN(n15636) );
  NAND2_X1 U18761 ( .A1(n15634), .A2(n16285), .ZN(n15635) );
  OAI211_X1 U18762 ( .C1(n16271), .C2(n18919), .A(n15636), .B(n15635), .ZN(
        n15639) );
  NOR2_X1 U18763 ( .A1(n15598), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16213) );
  NOR3_X1 U18764 ( .A1(n16213), .A2(n16212), .A3(n15637), .ZN(n15638) );
  AOI211_X1 U18765 ( .C1(n16216), .C2(n16283), .A(n15639), .B(n15638), .ZN(
        n15640) );
  INV_X1 U18766 ( .A(n15640), .ZN(P2_U3037) );
  INV_X1 U18767 ( .A(n15641), .ZN(n15643) );
  MUX2_X1 U18768 ( .A(n15643), .B(n15642), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n15644) );
  OAI21_X1 U18769 ( .B1(n15646), .B2(n15645), .A(n15644), .ZN(n16299) );
  AOI21_X1 U18770 ( .B1(n16299), .B2(n20990), .A(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n15649) );
  INV_X1 U18771 ( .A(n16334), .ZN(n15647) );
  OAI22_X1 U18772 ( .A1(n15650), .A2(n15649), .B1(n15648), .B2(n15647), .ZN(
        n15652) );
  MUX2_X1 U18773 ( .A(n15652), .B(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .S(
        n15651), .Z(P2_U3601) );
  AOI22_X1 U18774 ( .A1(n11696), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9834), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15656) );
  AOI22_X1 U18775 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15655) );
  AOI22_X1 U18776 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17107), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15654) );
  AOI22_X1 U18777 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17140), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15653) );
  NAND4_X1 U18778 ( .A1(n15656), .A2(n15655), .A3(n15654), .A4(n15653), .ZN(
        n15663) );
  AOI22_X1 U18779 ( .A1(n11630), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n15657), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15661) );
  AOI22_X1 U18780 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9831), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15660) );
  AOI22_X1 U18781 ( .A1(n11534), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15659) );
  AOI22_X1 U18782 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15658) );
  NAND4_X1 U18783 ( .A1(n15661), .A2(n15660), .A3(n15659), .A4(n15658), .ZN(
        n15662) );
  NOR2_X1 U18784 ( .A1(n15663), .A2(n15662), .ZN(n17293) );
  AND2_X1 U18785 ( .A1(n17184), .A2(n15664), .ZN(n17091) );
  NOR2_X1 U18786 ( .A1(n17160), .A2(n15664), .ZN(n17068) );
  AOI22_X1 U18787 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17091), .B1(n17068), 
        .B2(n16733), .ZN(n15665) );
  OAI21_X1 U18788 ( .B1(n17293), .B2(n17178), .A(n15665), .ZN(P3_U2690) );
  NAND2_X1 U18789 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18300) );
  AOI221_X1 U18790 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18300), .C1(n15667), 
        .C2(n18300), .A(n15666), .ZN(n18152) );
  NOR2_X1 U18791 ( .A1(n15668), .A2(n20915), .ZN(n15669) );
  OAI21_X1 U18792 ( .B1(n15669), .B2(n18211), .A(n18153), .ZN(n18150) );
  AOI22_X1 U18793 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18152), .B1(
        n18150), .B2(n18626), .ZN(P3_U2865) );
  NAND2_X1 U18794 ( .A1(n18631), .A2(n18803), .ZN(n15673) );
  INV_X1 U18795 ( .A(n18668), .ZN(n18794) );
  NAND2_X1 U18796 ( .A1(n18794), .A2(n15670), .ZN(n17351) );
  OAI211_X1 U18797 ( .C1(n17390), .C2(n18608), .A(n18631), .B(n18803), .ZN(
        n15767) );
  OAI21_X1 U18798 ( .B1(n15673), .B2(n17351), .A(n15767), .ZN(n15674) );
  INV_X1 U18799 ( .A(n18633), .ZN(n18613) );
  NOR2_X1 U18800 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18748), .ZN(n18159) );
  INV_X1 U18801 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18148) );
  NOR2_X1 U18802 ( .A1(n18148), .A2(n18746), .ZN(n15677) );
  INV_X1 U18803 ( .A(n18775), .ZN(n18772) );
  AND2_X1 U18804 ( .A1(n15678), .A2(n18608), .ZN(n18632) );
  NAND3_X1 U18805 ( .A1(n18772), .A2(n18810), .A3(n18632), .ZN(n15679) );
  OAI21_X1 U18806 ( .B1(n18772), .B2(n15680), .A(n15679), .ZN(P3_U3284) );
  OAI21_X1 U18807 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15682), .A(
        n15681), .ZN(n16365) );
  INV_X1 U18808 ( .A(n18594), .ZN(n18617) );
  NAND2_X1 U18809 ( .A1(n18617), .A2(n18629), .ZN(n17990) );
  AOI21_X1 U18810 ( .B1(n20889), .B2(n17990), .A(n15683), .ZN(n16376) );
  INV_X1 U18811 ( .A(n18144), .ZN(n18125) );
  NAND2_X1 U18812 ( .A1(n15755), .A2(n17463), .ZN(n16347) );
  INV_X1 U18813 ( .A(n17979), .ZN(n18049) );
  NAND2_X1 U18814 ( .A1(n17464), .A2(n15755), .ZN(n16346) );
  AOI22_X1 U18815 ( .A1(n18125), .A2(n16347), .B1(n18049), .B2(n16346), .ZN(
        n15756) );
  INV_X1 U18816 ( .A(n18055), .ZN(n18127) );
  AOI21_X1 U18817 ( .B1(n18127), .B2(n17465), .A(n18130), .ZN(n15684) );
  OAI211_X1 U18818 ( .C1(n16376), .C2(n18128), .A(n15756), .B(n15684), .ZN(
        n15687) );
  INV_X1 U18819 ( .A(n9828), .ZN(n18787) );
  INV_X1 U18820 ( .A(n18011), .ZN(n17723) );
  OAI22_X1 U18821 ( .A1(n18787), .A2(n18008), .B1(n17723), .B2(n18010), .ZN(
        n17982) );
  AOI21_X1 U18822 ( .B1(n17982), .B2(n17613), .A(n15685), .ZN(n17887) );
  INV_X1 U18823 ( .A(n17919), .ZN(n17911) );
  NOR2_X1 U18824 ( .A1(n16375), .A2(n17911), .ZN(n17832) );
  NOR2_X1 U18825 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16364), .ZN(
        n15686) );
  AOI22_X1 U18826 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15687), .B1(
        n17832), .B2(n15686), .ZN(n15688) );
  INV_X2 U18827 ( .A(n18138), .ZN(n18126) );
  NAND2_X1 U18828 ( .A1(n18126), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16362) );
  OAI211_X1 U18829 ( .C1(n18045), .C2(n16365), .A(n15688), .B(n16362), .ZN(
        P3_U2833) );
  AOI22_X1 U18830 ( .A1(n18874), .A2(n16285), .B1(n16280), .B2(n18873), .ZN(
        n15690) );
  OAI211_X1 U18831 ( .C1(n15691), .C2(n16278), .A(n15690), .B(n15689), .ZN(
        n15692) );
  INV_X1 U18832 ( .A(n15692), .ZN(n15693) );
  OAI221_X1 U18833 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15696), 
        .C1(n15695), .C2(n15694), .A(n15693), .ZN(P2_U3030) );
  INV_X1 U18834 ( .A(n15697), .ZN(n15699) );
  AOI22_X1 U18835 ( .A1(n15699), .A2(n18984), .B1(n18979), .B2(n15698), .ZN(
        n15708) );
  AOI211_X1 U18836 ( .C1(n15702), .C2(n15700), .A(n15701), .B(n19732), .ZN(
        n15706) );
  AOI22_X1 U18837 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n18968), .B1(
        P2_EBX_REG_22__SCAN_IN), .B2(n18978), .ZN(n15703) );
  OAI21_X1 U18838 ( .B1(n15704), .B2(n18982), .A(n15703), .ZN(n15705) );
  AOI211_X1 U18839 ( .C1(n18993), .C2(P2_REIP_REG_22__SCAN_IN), .A(n15706), 
        .B(n15705), .ZN(n15707) );
  NAND2_X1 U18840 ( .A1(n15708), .A2(n15707), .ZN(P2_U2833) );
  NOR2_X1 U18841 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(P1_MORE_REG_SCAN_IN), .ZN(
        n15730) );
  INV_X1 U18842 ( .A(n15718), .ZN(n15720) );
  AOI21_X1 U18843 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15710), .A(
        n15709), .ZN(n15713) );
  INV_X1 U18844 ( .A(n15713), .ZN(n15716) );
  INV_X1 U18845 ( .A(n20529), .ZN(n15715) );
  AOI211_X1 U18846 ( .C1(n20644), .C2(n15713), .A(n15712), .B(n15711), .ZN(
        n15714) );
  AOI211_X1 U18847 ( .C1(n20638), .C2(n15716), .A(n15715), .B(n15714), .ZN(
        n15717) );
  OAI21_X1 U18848 ( .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15718), .A(
        n15717), .ZN(n15719) );
  OAI21_X1 U18849 ( .B1(n15720), .B2(n20398), .A(n15719), .ZN(n15721) );
  OAI21_X1 U18850 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15722), .A(
        n15721), .ZN(n15726) );
  AOI21_X1 U18851 ( .B1(n15722), .B2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15725) );
  AOI211_X1 U18852 ( .C1(n15726), .C2(n15725), .A(n15724), .B(n15723), .ZN(
        n15727) );
  OAI211_X1 U18853 ( .C1(n15730), .C2(n15729), .A(n15728), .B(n15727), .ZN(
        n15735) );
  NOR2_X1 U18854 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20708), .ZN(n15734) );
  OR4_X1 U18855 ( .A1(n15732), .A2(n20812), .A3(n15761), .A4(n15731), .ZN(
        n15733) );
  OAI221_X1 U18856 ( .B1(n15736), .B2(n15734), .C1(n15736), .C2(n15760), .A(
        n15733), .ZN(n16041) );
  AOI221_X1 U18857 ( .B1(n20706), .B2(n20705), .C1(n15735), .C2(n20705), .A(
        n16041), .ZN(n15737) );
  NOR2_X1 U18858 ( .A1(n15737), .A2(n20706), .ZN(n16044) );
  OAI211_X1 U18859 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20818), .A(n16044), 
        .B(n15739), .ZN(n16042) );
  AOI21_X1 U18860 ( .B1(n15736), .B2(n15735), .A(n16042), .ZN(n15743) );
  INV_X1 U18861 ( .A(n15737), .ZN(n15738) );
  OAI21_X1 U18862 ( .B1(n15740), .B2(n15739), .A(n15738), .ZN(n15741) );
  AOI22_X1 U18863 ( .A1(n15743), .A2(n15742), .B1(n20706), .B2(n15741), .ZN(
        P1_U3161) );
  AOI22_X1 U18864 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n13703), .B1(n15744), 
        .B2(n21010), .ZN(n15751) );
  NOR3_X1 U18865 ( .A1(n14902), .A2(n15895), .A3(n15745), .ZN(n15748) );
  NOR2_X1 U18866 ( .A1(n15748), .A2(n15747), .ZN(n15749) );
  XNOR2_X1 U18867 ( .A(n15749), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15879) );
  AOI22_X1 U18868 ( .A1(n15879), .A2(n20087), .B1(n20110), .B2(n15811), .ZN(
        n15750) );
  OAI211_X1 U18869 ( .C1(n21010), .C2(n15752), .A(n15751), .B(n15750), .ZN(
        P1_U3010) );
  OAI21_X1 U18870 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15754), .A(
        n15753), .ZN(n16358) );
  AND2_X1 U18871 ( .A1(n16348), .A2(n15755), .ZN(n16356) );
  AOI21_X1 U18872 ( .B1(n15757), .B2(n15756), .A(n16348), .ZN(n15758) );
  AOI21_X1 U18873 ( .B1(n17832), .B2(n16356), .A(n15758), .ZN(n15759) );
  NAND2_X1 U18874 ( .A1(n18126), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16352) );
  OAI211_X1 U18875 ( .C1(n18045), .C2(n16358), .A(n15759), .B(n16352), .ZN(
        P3_U2832) );
  INV_X1 U18876 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20724) );
  INV_X1 U18877 ( .A(HOLD), .ZN(n20723) );
  NOR2_X1 U18878 ( .A1(n20724), .A2(n20723), .ZN(n20711) );
  AOI22_X1 U18879 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n15762) );
  NAND2_X1 U18880 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n15760), .ZN(n20717) );
  OAI211_X1 U18881 ( .C1(n20711), .C2(n15762), .A(n15761), .B(n20717), .ZN(
        P1_U3195) );
  AND2_X1 U18882 ( .A1(n20004), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR3_X1 U18883 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19859), .A3(n19858), 
        .ZN(n16327) );
  INV_X1 U18884 ( .A(n16329), .ZN(n16344) );
  OAI211_X1 U18885 ( .C1(P2_STATEBS16_REG_SCAN_IN), .C2(n15763), .A(n16344), 
        .B(n19857), .ZN(n15764) );
  NOR2_X1 U18886 ( .A1(n16327), .A2(n15764), .ZN(P2_U3178) );
  OAI221_X1 U18887 ( .B1(n10990), .B2(n16344), .C1(n16330), .C2(n16344), .A(
        n19585), .ZN(n19842) );
  NOR2_X1 U18888 ( .A1(n16325), .A2(n19842), .ZN(P2_U3047) );
  OAI22_X2 U18889 ( .A1(n18651), .A2(n15767), .B1(n15766), .B2(n15765), .ZN(
        n17195) );
  NAND2_X1 U18890 ( .A1(n18188), .A2(n17195), .ZN(n17337) );
  INV_X1 U18891 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17424) );
  INV_X1 U18892 ( .A(n17195), .ZN(n17344) );
  AOI22_X1 U18893 ( .A1(n17345), .A2(BUF2_REG_0__SCAN_IN), .B1(n17317), .B2(
        n15768), .ZN(n15769) );
  OAI221_X1 U18894 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17337), .C1(n17424), 
        .C2(n17195), .A(n15769), .ZN(P3_U2735) );
  AOI21_X1 U18895 ( .B1(n19945), .B2(n15781), .A(n19932), .ZN(n15791) );
  NAND2_X1 U18896 ( .A1(n19945), .A2(n20762), .ZN(n15780) );
  AOI21_X1 U18897 ( .B1(n15791), .B2(n15780), .A(n14876), .ZN(n15773) );
  NAND2_X1 U18898 ( .A1(n19945), .A2(n15770), .ZN(n15771) );
  OAI22_X1 U18899 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n15771), .B1(n12951), 
        .B2(n19899), .ZN(n15772) );
  AOI211_X1 U18900 ( .C1(n19961), .C2(P1_EBX_REG_25__SCAN_IN), .A(n15773), .B(
        n15772), .ZN(n15778) );
  OAI22_X1 U18901 ( .A1(n15775), .A2(n15867), .B1(n15774), .B2(n15859), .ZN(
        n15776) );
  INV_X1 U18902 ( .A(n15776), .ZN(n15777) );
  OAI211_X1 U18903 ( .C1(n15779), .C2(n19959), .A(n15778), .B(n15777), .ZN(
        P1_U2815) );
  OAI22_X1 U18904 ( .A1(n15791), .A2(n20762), .B1(n15781), .B2(n15780), .ZN(
        n15782) );
  AOI21_X1 U18905 ( .B1(P1_EBX_REG_24__SCAN_IN), .B2(n19961), .A(n15782), .ZN(
        n15788) );
  OAI22_X1 U18906 ( .A1(n15784), .A2(n15867), .B1(n15783), .B2(n15859), .ZN(
        n15785) );
  AOI21_X1 U18907 ( .B1(n15786), .B2(n19971), .A(n15785), .ZN(n15787) );
  OAI211_X1 U18908 ( .C1(n20903), .C2(n19899), .A(n15788), .B(n15787), .ZN(
        P1_U2816) );
  AOI22_X1 U18909 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n19964), .B1(
        P1_EBX_REG_23__SCAN_IN), .B2(n19961), .ZN(n15795) );
  INV_X1 U18910 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21030) );
  INV_X1 U18911 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20759) );
  NOR2_X1 U18912 ( .A1(n21030), .A2(n20759), .ZN(n15801) );
  NOR2_X1 U18913 ( .A1(n15789), .A2(n15815), .ZN(n15809) );
  AOI21_X1 U18914 ( .B1(n15801), .B2(n15809), .A(P1_REIP_REG_23__SCAN_IN), 
        .ZN(n15792) );
  OAI22_X1 U18915 ( .A1(n15792), .A2(n15791), .B1(n15790), .B2(n15859), .ZN(
        n15793) );
  AOI21_X1 U18916 ( .B1(n15875), .B2(n19928), .A(n15793), .ZN(n15794) );
  OAI211_X1 U18917 ( .C1(n15878), .C2(n19959), .A(n15795), .B(n15794), .ZN(
        P1_U2817) );
  AOI22_X1 U18918 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19964), .B1(
        P1_EBX_REG_22__SCAN_IN), .B2(n19961), .ZN(n15806) );
  OAI21_X1 U18919 ( .B1(n15797), .B2(n19934), .A(n15796), .ZN(n15821) );
  AOI22_X1 U18920 ( .A1(n15798), .A2(n19971), .B1(P1_REIP_REG_22__SCAN_IN), 
        .B2(n15821), .ZN(n15805) );
  AOI22_X1 U18921 ( .A1(n15800), .A2(n19928), .B1(n19960), .B2(n15799), .ZN(
        n15804) );
  INV_X1 U18922 ( .A(n15801), .ZN(n15802) );
  OAI211_X1 U18923 ( .C1(P1_REIP_REG_22__SCAN_IN), .C2(P1_REIP_REG_21__SCAN_IN), .A(n15809), .B(n15802), .ZN(n15803) );
  NAND4_X1 U18924 ( .A1(n15806), .A2(n15805), .A3(n15804), .A4(n15803), .ZN(
        P1_U2818) );
  AOI22_X1 U18925 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n19964), .B1(
        P1_EBX_REG_21__SCAN_IN), .B2(n19961), .ZN(n15807) );
  OAI21_X1 U18926 ( .B1(n15883), .B2(n19959), .A(n15807), .ZN(n15808) );
  AOI221_X1 U18927 ( .B1(n15821), .B2(P1_REIP_REG_21__SCAN_IN), .C1(n15809), 
        .C2(n20759), .A(n15808), .ZN(n15813) );
  INV_X1 U18928 ( .A(n15810), .ZN(n15880) );
  AOI22_X1 U18929 ( .A1(n15880), .A2(n19928), .B1(n19960), .B2(n15811), .ZN(
        n15812) );
  NAND2_X1 U18930 ( .A1(n15813), .A2(n15812), .ZN(P1_U2819) );
  AOI22_X1 U18931 ( .A1(n15814), .A2(n19971), .B1(P1_EBX_REG_20__SCAN_IN), 
        .B2(n19961), .ZN(n15823) );
  NAND2_X1 U18932 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n15825) );
  INV_X1 U18933 ( .A(n15815), .ZN(n15854) );
  NAND2_X1 U18934 ( .A1(n15816), .A2(n15854), .ZN(n15839) );
  INV_X1 U18935 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20756) );
  OAI21_X1 U18936 ( .B1(n15825), .B2(n15839), .A(n20756), .ZN(n15820) );
  OAI22_X1 U18937 ( .A1(n15818), .A2(n15867), .B1(n15859), .B2(n15817), .ZN(
        n15819) );
  AOI21_X1 U18938 ( .B1(n15821), .B2(n15820), .A(n15819), .ZN(n15822) );
  OAI211_X1 U18939 ( .C1(n15824), .C2(n19899), .A(n15823), .B(n15822), .ZN(
        P1_U2820) );
  OAI21_X1 U18940 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(P1_REIP_REG_18__SCAN_IN), 
        .A(n15825), .ZN(n15830) );
  AOI22_X1 U18941 ( .A1(P1_EBX_REG_19__SCAN_IN), .A2(n19961), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n15831), .ZN(n15826) );
  OAI21_X1 U18942 ( .B1(n15890), .B2(n19959), .A(n15826), .ZN(n15827) );
  AOI211_X1 U18943 ( .C1(n19964), .C2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n19948), .B(n15827), .ZN(n15829) );
  AOI22_X1 U18944 ( .A1(n15887), .A2(n19928), .B1(n19960), .B2(n15948), .ZN(
        n15828) );
  OAI211_X1 U18945 ( .C1(n15839), .C2(n15830), .A(n15829), .B(n15828), .ZN(
        P1_U2821) );
  AOI22_X1 U18946 ( .A1(P1_EBX_REG_18__SCAN_IN), .A2(n19961), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n15831), .ZN(n15832) );
  OAI211_X1 U18947 ( .C1(n19899), .C2(n20923), .A(n15832), .B(n19923), .ZN(
        n15836) );
  OAI22_X1 U18948 ( .A1(n15834), .A2(n15867), .B1(n15859), .B2(n15833), .ZN(
        n15835) );
  AOI211_X1 U18949 ( .C1(n15837), .C2(n19971), .A(n15836), .B(n15835), .ZN(
        n15838) );
  OAI21_X1 U18950 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(n15839), .A(n15838), 
        .ZN(P1_U2822) );
  AOI22_X1 U18951 ( .A1(P1_EBX_REG_16__SCAN_IN), .A2(n19961), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n15855), .ZN(n15840) );
  OAI211_X1 U18952 ( .C1(n19899), .C2(n15841), .A(n15840), .B(n19923), .ZN(
        n15845) );
  OAI22_X1 U18953 ( .A1(n15843), .A2(n15867), .B1(n15859), .B2(n15842), .ZN(
        n15844) );
  AOI211_X1 U18954 ( .C1(n15846), .C2(n19971), .A(n15845), .B(n15844), .ZN(
        n15849) );
  OAI211_X1 U18955 ( .C1(P1_REIP_REG_16__SCAN_IN), .C2(P1_REIP_REG_15__SCAN_IN), .A(n15854), .B(n15847), .ZN(n15848) );
  NAND2_X1 U18956 ( .A1(n15849), .A2(n15848), .ZN(P1_U2824) );
  INV_X1 U18957 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20749) );
  AOI22_X1 U18958 ( .A1(P1_EBX_REG_15__SCAN_IN), .A2(n19961), .B1(n19960), 
        .B2(n15850), .ZN(n15851) );
  OAI211_X1 U18959 ( .C1(n19899), .C2(n15852), .A(n15851), .B(n19923), .ZN(
        n15853) );
  AOI221_X1 U18960 ( .B1(n15855), .B2(P1_REIP_REG_15__SCAN_IN), .C1(n15854), 
        .C2(n20749), .A(n15853), .ZN(n15857) );
  AOI22_X1 U18961 ( .A1(n15911), .A2(n19928), .B1(n19971), .B2(n15910), .ZN(
        n15856) );
  NAND2_X1 U18962 ( .A1(n15857), .A2(n15856), .ZN(P1_U2825) );
  OAI22_X1 U18963 ( .A1(n15860), .A2(n19899), .B1(n15859), .B2(n15858), .ZN(
        n15861) );
  AOI211_X1 U18964 ( .C1(n19961), .C2(P1_EBX_REG_12__SCAN_IN), .A(n19948), .B(
        n15861), .ZN(n15866) );
  NAND2_X1 U18965 ( .A1(n20744), .A2(n15862), .ZN(n15863) );
  AOI22_X1 U18966 ( .A1(n15916), .A2(n19971), .B1(n15864), .B2(n15863), .ZN(
        n15865) );
  OAI211_X1 U18967 ( .C1(n15867), .C2(n15914), .A(n15866), .B(n15865), .ZN(
        P1_U2828) );
  AOI22_X1 U18968 ( .A1(P1_EBX_REG_11__SCAN_IN), .A2(n19961), .B1(n19960), 
        .B2(n15982), .ZN(n15868) );
  OAI21_X1 U18969 ( .B1(n20743), .B2(n15869), .A(n15868), .ZN(n15870) );
  AOI211_X1 U18970 ( .C1(n19964), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n19948), .B(n15870), .ZN(n15873) );
  AOI22_X1 U18971 ( .A1(n15925), .A2(n19928), .B1(n15871), .B2(n20743), .ZN(
        n15872) );
  OAI211_X1 U18972 ( .C1(n15928), .C2(n19959), .A(n15873), .B(n15872), .ZN(
        P1_U2829) );
  AOI22_X1 U18973 ( .A1(n20065), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B1(
        n13703), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n15877) );
  AOI22_X1 U18974 ( .A1(n15875), .A2(n20071), .B1(n20072), .B2(n15874), .ZN(
        n15876) );
  OAI211_X1 U18975 ( .C1(n20076), .C2(n15878), .A(n15877), .B(n15876), .ZN(
        P1_U2976) );
  AOI22_X1 U18976 ( .A1(n20065), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n13703), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n15882) );
  AOI22_X1 U18977 ( .A1(n15880), .A2(n20071), .B1(n20072), .B2(n15879), .ZN(
        n15881) );
  OAI211_X1 U18978 ( .C1(n20076), .C2(n15883), .A(n15882), .B(n15881), .ZN(
        P1_U2978) );
  AOI22_X1 U18979 ( .A1(n20065), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n13703), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15889) );
  NOR2_X1 U18980 ( .A1(n13225), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15884) );
  MUX2_X1 U18981 ( .A(n13225), .B(n15884), .S(n14902), .Z(n15886) );
  XNOR2_X1 U18982 ( .A(n15886), .B(n15885), .ZN(n15949) );
  AOI22_X1 U18983 ( .A1(n15887), .A2(n20071), .B1(n20072), .B2(n15949), .ZN(
        n15888) );
  OAI211_X1 U18984 ( .C1(n20076), .C2(n15890), .A(n15889), .B(n15888), .ZN(
        P1_U2980) );
  OAI21_X1 U18985 ( .B1(n15893), .B2(n15892), .A(n15891), .ZN(n15897) );
  NAND2_X1 U18986 ( .A1(n15897), .A2(n15894), .ZN(n15896) );
  MUX2_X1 U18987 ( .A(n15897), .B(n15896), .S(n15895), .Z(n15898) );
  XOR2_X1 U18988 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B(n15898), .Z(
        n15961) );
  AOI22_X1 U18989 ( .A1(n20065), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n13703), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n15903) );
  OAI22_X1 U18990 ( .A1(n15900), .A2(n20120), .B1(n15899), .B2(n20076), .ZN(
        n15901) );
  INV_X1 U18991 ( .A(n15901), .ZN(n15902) );
  OAI211_X1 U18992 ( .C1(n15961), .C2(n19882), .A(n15903), .B(n15902), .ZN(
        P1_U2982) );
  OR2_X1 U18993 ( .A1(n15905), .A2(n15904), .ZN(n15909) );
  OR2_X1 U18994 ( .A1(n13225), .A2(n13237), .ZN(n15906) );
  AND2_X1 U18995 ( .A1(n15907), .A2(n15906), .ZN(n15908) );
  XNOR2_X1 U18996 ( .A(n15909), .B(n15908), .ZN(n15964) );
  AOI22_X1 U18997 ( .A1(n20065), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n13703), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n15913) );
  AOI22_X1 U18998 ( .A1(n15911), .A2(n20071), .B1(n15917), .B2(n15910), .ZN(
        n15912) );
  OAI211_X1 U18999 ( .C1(n15964), .C2(n19882), .A(n15913), .B(n15912), .ZN(
        P1_U2984) );
  AOI22_X1 U19000 ( .A1(n20065), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n13703), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15919) );
  INV_X1 U19001 ( .A(n15914), .ZN(n15915) );
  AOI22_X1 U19002 ( .A1(n15917), .A2(n15916), .B1(n20071), .B2(n15915), .ZN(
        n15918) );
  OAI211_X1 U19003 ( .C1(n15920), .C2(n19882), .A(n15919), .B(n15918), .ZN(
        P1_U2987) );
  AOI22_X1 U19004 ( .A1(n20065), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n13703), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15927) );
  NAND3_X1 U19005 ( .A1(n15921), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n13225), .ZN(n15923) );
  NAND2_X1 U19006 ( .A1(n15923), .A2(n15922), .ZN(n15924) );
  XOR2_X1 U19007 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n15924), .Z(
        n15983) );
  AOI22_X1 U19008 ( .A1(n20072), .A2(n15983), .B1(n20071), .B2(n15925), .ZN(
        n15926) );
  OAI211_X1 U19009 ( .C1(n20076), .C2(n15928), .A(n15927), .B(n15926), .ZN(
        P1_U2988) );
  AOI22_X1 U19010 ( .A1(n20065), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n13703), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15934) );
  NAND2_X1 U19011 ( .A1(n15930), .A2(n15929), .ZN(n15931) );
  XNOR2_X1 U19012 ( .A(n15932), .B(n15931), .ZN(n16021) );
  AOI22_X1 U19013 ( .A1(n16021), .A2(n20072), .B1(n20071), .B2(n19917), .ZN(
        n15933) );
  OAI211_X1 U19014 ( .C1(n20076), .C2(n19912), .A(n15934), .B(n15933), .ZN(
        P1_U2992) );
  AOI22_X1 U19015 ( .A1(n20065), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n13703), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n15940) );
  XNOR2_X1 U19016 ( .A(n15936), .B(n15935), .ZN(n15937) );
  XNOR2_X1 U19017 ( .A(n15938), .B(n15937), .ZN(n16027) );
  AOI22_X1 U19018 ( .A1(n16027), .A2(n20072), .B1(n20071), .B2(n19927), .ZN(
        n15939) );
  OAI211_X1 U19019 ( .C1(n20076), .C2(n19931), .A(n15940), .B(n15939), .ZN(
        P1_U2993) );
  AOI22_X1 U19020 ( .A1(n20065), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n13703), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n15946) );
  OAI21_X1 U19021 ( .B1(n15943), .B2(n15942), .A(n15941), .ZN(n15944) );
  INV_X1 U19022 ( .A(n15944), .ZN(n16031) );
  AOI22_X1 U19023 ( .A1(n16031), .A2(n20072), .B1(n20071), .B2(n19939), .ZN(
        n15945) );
  OAI211_X1 U19024 ( .C1(n20076), .C2(n19937), .A(n15946), .B(n15945), .ZN(
        P1_U2994) );
  AOI22_X1 U19025 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n15947), .B1(
        n13703), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15951) );
  AOI22_X1 U19026 ( .A1(n15949), .A2(n20087), .B1(n20110), .B2(n15948), .ZN(
        n15950) );
  OAI211_X1 U19027 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15952), .A(
        n15951), .B(n15950), .ZN(P1_U3012) );
  NAND2_X1 U19028 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15955) );
  OAI21_X1 U19029 ( .B1(n15955), .B2(n15954), .A(n15953), .ZN(n15957) );
  AOI22_X1 U19030 ( .A1(n15958), .A2(n15957), .B1(n20110), .B2(n15956), .ZN(
        n15960) );
  NAND2_X1 U19031 ( .A1(n13703), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n15959) );
  OAI211_X1 U19032 ( .C1(n15961), .C2(n20105), .A(n15960), .B(n15959), .ZN(
        P1_U3014) );
  INV_X1 U19033 ( .A(n15962), .ZN(n15967) );
  OAI22_X1 U19034 ( .A1(n16014), .A2(n15963), .B1(n20749), .B2(n20102), .ZN(
        n15966) );
  NOR2_X1 U19035 ( .A1(n15964), .A2(n20105), .ZN(n15965) );
  AOI211_X1 U19036 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15967), .A(
        n15966), .B(n15965), .ZN(n15969) );
  NAND2_X1 U19037 ( .A1(n15969), .A2(n15968), .ZN(P1_U3016) );
  OAI221_X1 U19038 ( .B1(n15973), .B2(n15972), .C1(n15973), .C2(n15971), .A(
        n15970), .ZN(n15980) );
  AOI22_X1 U19039 ( .A1(n15975), .A2(n20087), .B1(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n15974), .ZN(n15979) );
  NAND2_X1 U19040 ( .A1(n13703), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n15978) );
  NAND2_X1 U19041 ( .A1(n20110), .A2(n15976), .ZN(n15977) );
  NAND4_X1 U19042 ( .A1(n15980), .A2(n15979), .A3(n15978), .A4(n15977), .ZN(
        P1_U3018) );
  INV_X1 U19043 ( .A(n15981), .ZN(n15987) );
  AOI22_X1 U19044 ( .A1(n20110), .A2(n15982), .B1(n13703), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n15986) );
  AOI22_X1 U19045 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n15984), .B1(
        n20087), .B2(n15983), .ZN(n15985) );
  OAI211_X1 U19046 ( .C1(n16030), .C2(n15987), .A(n15986), .B(n15985), .ZN(
        P1_U3020) );
  INV_X1 U19047 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15999) );
  NAND2_X1 U19048 ( .A1(n15989), .A2(n15988), .ZN(n15995) );
  OAI21_X1 U19049 ( .B1(n20098), .B2(n20113), .A(n20096), .ZN(n16007) );
  NAND2_X1 U19050 ( .A1(n15990), .A2(n16007), .ZN(n20077) );
  OAI21_X1 U19051 ( .B1(n15995), .B2(n20077), .A(n15991), .ZN(n16005) );
  OAI22_X1 U19052 ( .A1(n16014), .A2(n15992), .B1(n20740), .B2(n20102), .ZN(
        n15993) );
  AOI21_X1 U19053 ( .B1(n20087), .B2(n15994), .A(n15993), .ZN(n15998) );
  NOR2_X1 U19054 ( .A1(n15996), .A2(n15995), .ZN(n16001) );
  OAI221_X1 U19055 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n15999), .C2(n16006), .A(
        n16001), .ZN(n15997) );
  OAI211_X1 U19056 ( .C1(n15999), .C2(n16005), .A(n15998), .B(n15997), .ZN(
        P1_U3021) );
  AOI21_X1 U19057 ( .B1(n20110), .B2(n19903), .A(n16000), .ZN(n16004) );
  AOI22_X1 U19058 ( .A1(n16002), .A2(n20087), .B1(n16001), .B2(n16006), .ZN(
        n16003) );
  OAI211_X1 U19059 ( .C1(n16006), .C2(n16005), .A(n16004), .B(n16003), .ZN(
        P1_U3022) );
  NOR2_X1 U19060 ( .A1(n20081), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16032) );
  INV_X1 U19061 ( .A(n16032), .ZN(n16010) );
  NAND2_X1 U19062 ( .A1(n16008), .A2(n16007), .ZN(n16009) );
  AOI21_X1 U19063 ( .B1(n20096), .B2(n20081), .A(n16009), .ZN(n16036) );
  OAI21_X1 U19064 ( .B1(n16011), .B2(n16010), .A(n16036), .ZN(n16026) );
  AOI21_X1 U19065 ( .B1(n15935), .B2(n16012), .A(n16026), .ZN(n16025) );
  OAI222_X1 U19066 ( .A1(n16015), .A2(n16014), .B1(n20102), .B2(n20737), .C1(
        n20105), .C2(n16013), .ZN(n16016) );
  INV_X1 U19067 ( .A(n16016), .ZN(n16018) );
  NOR2_X1 U19068 ( .A1(n15935), .A2(n16030), .ZN(n16020) );
  OAI221_X1 U19069 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16019), .C2(n16024), .A(
        n16020), .ZN(n16017) );
  OAI211_X1 U19070 ( .C1(n16025), .C2(n16019), .A(n16018), .B(n16017), .ZN(
        P1_U3023) );
  AOI22_X1 U19071 ( .A1(n20110), .A2(n19910), .B1(n13703), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n16023) );
  AOI22_X1 U19072 ( .A1(n16021), .A2(n20087), .B1(n16020), .B2(n16024), .ZN(
        n16022) );
  OAI211_X1 U19073 ( .C1(n16025), .C2(n16024), .A(n16023), .B(n16022), .ZN(
        P1_U3024) );
  AOI22_X1 U19074 ( .A1(n20110), .A2(n19922), .B1(n13703), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n16029) );
  AOI22_X1 U19075 ( .A1(n16027), .A2(n20087), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16026), .ZN(n16028) );
  OAI211_X1 U19076 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n16030), .A(
        n16029), .B(n16028), .ZN(P1_U3025) );
  AOI22_X1 U19077 ( .A1(n20110), .A2(n19936), .B1(n13703), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n16034) );
  AOI22_X1 U19078 ( .A1(n20089), .A2(n16032), .B1(n20087), .B2(n16031), .ZN(
        n16033) );
  OAI211_X1 U19079 ( .C1(n16036), .C2(n16035), .A(n16034), .B(n16033), .ZN(
        P1_U3026) );
  NAND4_X1 U19080 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n20708), .A4(n20818), .ZN(n16037) );
  AND2_X1 U19081 ( .A1(n16038), .A2(n16037), .ZN(n20707) );
  NAND2_X1 U19082 ( .A1(n20707), .A2(n16039), .ZN(n16040) );
  AOI22_X1 U19083 ( .A1(n20705), .A2(n16042), .B1(n16041), .B2(n16040), .ZN(
        P1_U3162) );
  OAI21_X1 U19084 ( .B1(n16044), .B2(n20537), .A(n16043), .ZN(P1_U3466) );
  AOI22_X1 U19085 ( .A1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n18968), .B1(
        P2_REIP_REG_31__SCAN_IN), .B2(n18993), .ZN(n16055) );
  AOI22_X1 U19086 ( .A1(n16045), .A2(n18984), .B1(n18979), .B2(n18997), .ZN(
        n16054) );
  NAND4_X1 U19087 ( .A1(n18961), .A2(n16046), .A3(n16047), .A4(n18954), .ZN(
        n16053) );
  AOI21_X1 U19088 ( .B1(n16049), .B2(n16048), .A(n18978), .ZN(n16051) );
  OR2_X1 U19089 ( .A1(n16051), .A2(n16050), .ZN(n16052) );
  NAND4_X1 U19090 ( .A1(n16055), .A2(n16054), .A3(n16053), .A4(n16052), .ZN(
        P2_U2824) );
  AOI21_X1 U19091 ( .B1(n16057), .B2(n16056), .A(n19732), .ZN(n16069) );
  INV_X1 U19092 ( .A(n16059), .ZN(n16062) );
  AOI22_X1 U19093 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18968), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n18993), .ZN(n16060) );
  OAI21_X1 U19094 ( .B1(n18950), .B2(n21118), .A(n16060), .ZN(n16061) );
  OAI21_X1 U19095 ( .B1(n16064), .B2(n18982), .A(n16063), .ZN(n16065) );
  INV_X1 U19096 ( .A(n16065), .ZN(n16066) );
  OAI21_X1 U19097 ( .B1(n15439), .B2(n18958), .A(n16066), .ZN(n16067) );
  INV_X1 U19098 ( .A(n16070), .ZN(P2_U2826) );
  INV_X1 U19099 ( .A(n16071), .ZN(n16073) );
  AOI22_X1 U19100 ( .A1(n16073), .A2(n18984), .B1(n16072), .B2(n18979), .ZN(
        n16081) );
  AOI211_X1 U19101 ( .C1(n16075), .C2(n9887), .A(n16074), .B(n19732), .ZN(
        n16079) );
  AOI22_X1 U19102 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18968), .B1(
        P2_EBX_REG_28__SCAN_IN), .B2(n18978), .ZN(n16076) );
  OAI21_X1 U19103 ( .B1(n16077), .B2(n18982), .A(n16076), .ZN(n16078) );
  AOI211_X1 U19104 ( .C1(n18993), .C2(P2_REIP_REG_28__SCAN_IN), .A(n16079), 
        .B(n16078), .ZN(n16080) );
  NAND2_X1 U19105 ( .A1(n16081), .A2(n16080), .ZN(P2_U2827) );
  AOI211_X1 U19106 ( .C1(n16084), .C2(n16083), .A(n16082), .B(n19732), .ZN(
        n16096) );
  OAI22_X1 U19107 ( .A1(n18950), .A2(n16086), .B1(n16085), .B2(n18990), .ZN(
        n16087) );
  AOI21_X1 U19108 ( .B1(n18993), .B2(P2_REIP_REG_27__SCAN_IN), .A(n16087), 
        .ZN(n16093) );
  INV_X1 U19109 ( .A(n16088), .ZN(n16090) );
  OAI211_X1 U19110 ( .C1(n16091), .C2(n16090), .A(n16089), .B(n18928), .ZN(
        n16092) );
  OAI211_X1 U19111 ( .C1(n16094), .C2(n18973), .A(n16093), .B(n16092), .ZN(
        n16095) );
  AOI211_X1 U19112 ( .C1(n18979), .C2(n16097), .A(n16096), .B(n16095), .ZN(
        n16098) );
  INV_X1 U19113 ( .A(n16098), .ZN(P2_U2828) );
  AOI22_X1 U19114 ( .A1(P2_REIP_REG_26__SCAN_IN), .A2(n18993), .B1(n16099), 
        .B2(n18928), .ZN(n16109) );
  AOI22_X1 U19115 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n18968), .B1(
        P2_EBX_REG_26__SCAN_IN), .B2(n18978), .ZN(n16108) );
  AOI22_X1 U19116 ( .A1(n16101), .A2(n18984), .B1(n18979), .B2(n16100), .ZN(
        n16107) );
  AOI21_X1 U19117 ( .B1(n16104), .B2(n16103), .A(n16102), .ZN(n16105) );
  NAND2_X1 U19118 ( .A1(n18961), .A2(n16105), .ZN(n16106) );
  NAND4_X1 U19119 ( .A1(n16109), .A2(n16108), .A3(n16107), .A4(n16106), .ZN(
        P2_U2829) );
  AOI211_X1 U19120 ( .C1(n16112), .C2(n16111), .A(n16110), .B(n19732), .ZN(
        n16120) );
  NAND2_X1 U19121 ( .A1(n18993), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n16114) );
  AOI22_X1 U19122 ( .A1(n18978), .A2(P2_EBX_REG_25__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n18968), .ZN(n16113) );
  OAI211_X1 U19123 ( .C1(n16115), .C2(n18973), .A(n16114), .B(n16113), .ZN(
        n16116) );
  AOI21_X1 U19124 ( .B1(n16117), .B2(n18928), .A(n16116), .ZN(n16118) );
  INV_X1 U19125 ( .A(n16118), .ZN(n16119) );
  AOI211_X1 U19126 ( .C1(n18979), .C2(n16121), .A(n16120), .B(n16119), .ZN(
        n16122) );
  INV_X1 U19127 ( .A(n16122), .ZN(P2_U2830) );
  AOI22_X1 U19128 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(n18978), .B1(n16123), 
        .B2(n18928), .ZN(n16133) );
  AOI22_X1 U19129 ( .A1(P2_REIP_REG_24__SCAN_IN), .A2(n18993), .B1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n18968), .ZN(n16132) );
  OAI22_X1 U19130 ( .A1(n16124), .A2(n18973), .B1(n18958), .B2(n16137), .ZN(
        n16125) );
  INV_X1 U19131 ( .A(n16125), .ZN(n16131) );
  AOI21_X1 U19132 ( .B1(n16128), .B2(n16127), .A(n16126), .ZN(n16129) );
  NAND2_X1 U19133 ( .A1(n18961), .A2(n16129), .ZN(n16130) );
  NAND4_X1 U19134 ( .A1(n16133), .A2(n16132), .A3(n16131), .A4(n16130), .ZN(
        P2_U2831) );
  INV_X1 U19135 ( .A(n16134), .ZN(n16135) );
  AOI22_X1 U19136 ( .A1(n16135), .A2(n19006), .B1(P2_EAX_REG_24__SCAN_IN), 
        .B2(n19050), .ZN(n16142) );
  AOI22_X1 U19137 ( .A1(n18998), .A2(BUF1_REG_24__SCAN_IN), .B1(n18999), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n16141) );
  INV_X1 U19138 ( .A(n16137), .ZN(n16138) );
  AOI22_X1 U19139 ( .A1(n16139), .A2(n19052), .B1(n19051), .B2(n16138), .ZN(
        n16140) );
  NAND3_X1 U19140 ( .A1(n16142), .A2(n16141), .A3(n16140), .ZN(P2_U2895) );
  OAI22_X1 U19141 ( .A1(n18865), .A2(n16243), .B1(n19776), .B2(n18878), .ZN(
        n16143) );
  AOI21_X1 U19142 ( .B1(n16234), .B2(n18858), .A(n16143), .ZN(n16147) );
  AOI22_X1 U19143 ( .A1(n16145), .A2(n10996), .B1(n16228), .B2(n16144), .ZN(
        n16146) );
  OAI211_X1 U19144 ( .C1(n19157), .C2(n18860), .A(n16147), .B(n16146), .ZN(
        P2_U2995) );
  AOI22_X1 U19145 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n19137), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n19138), .ZN(n16153) );
  OAI22_X1 U19146 ( .A1(n16149), .A2(n19142), .B1(n19140), .B2(n16148), .ZN(
        n16150) );
  AOI21_X1 U19147 ( .B1(n19146), .B2(n16151), .A(n16150), .ZN(n16152) );
  OAI211_X1 U19148 ( .C1(n19150), .C2(n16154), .A(n16153), .B(n16152), .ZN(
        P2_U2996) );
  AOI22_X1 U19149 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19138), .B1(n16234), 
        .B2(n16155), .ZN(n16162) );
  AOI22_X1 U19150 ( .A1(n16157), .A2(n16228), .B1(n19146), .B2(n16156), .ZN(
        n16158) );
  OAI21_X1 U19151 ( .B1(n16159), .B2(n19142), .A(n16158), .ZN(n16160) );
  INV_X1 U19152 ( .A(n16160), .ZN(n16161) );
  OAI211_X1 U19153 ( .C1(n16163), .C2(n16243), .A(n16162), .B(n16161), .ZN(
        P2_U2999) );
  AOI22_X1 U19154 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19137), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19138), .ZN(n16168) );
  OAI22_X1 U19155 ( .A1(n16165), .A2(n19142), .B1(n19140), .B2(n16164), .ZN(
        n16166) );
  AOI21_X1 U19156 ( .B1(n19146), .B2(n18885), .A(n16166), .ZN(n16167) );
  OAI211_X1 U19157 ( .C1(n19150), .C2(n18883), .A(n16168), .B(n16167), .ZN(
        P2_U3000) );
  AOI22_X1 U19158 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19138), .B1(n16234), 
        .B2(n18894), .ZN(n16173) );
  OAI22_X1 U19159 ( .A1(n16169), .A2(n19142), .B1(n19157), .B2(n18896), .ZN(
        n16170) );
  AOI21_X1 U19160 ( .B1(n16171), .B2(n16228), .A(n16170), .ZN(n16172) );
  OAI211_X1 U19161 ( .C1(n18890), .C2(n16243), .A(n16173), .B(n16172), .ZN(
        P2_U3001) );
  AOI22_X1 U19162 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n16261), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19137), .ZN(n16185) );
  INV_X1 U19163 ( .A(n16195), .ZN(n16177) );
  INV_X1 U19164 ( .A(n16174), .ZN(n16175) );
  AOI21_X1 U19165 ( .B1(n16177), .B2(n16176), .A(n16175), .ZN(n16251) );
  INV_X1 U19166 ( .A(n16251), .ZN(n16181) );
  NAND2_X1 U19167 ( .A1(n9858), .A2(n16178), .ZN(n16180) );
  XOR2_X1 U19168 ( .A(n16180), .B(n16179), .Z(n16253) );
  OAI22_X1 U19169 ( .A1(n16181), .A2(n19140), .B1(n16253), .B2(n19142), .ZN(
        n16182) );
  AOI21_X1 U19170 ( .B1(n19146), .B2(n16183), .A(n16182), .ZN(n16184) );
  OAI211_X1 U19171 ( .C1(n19150), .C2(n16186), .A(n16185), .B(n16184), .ZN(
        P2_U3002) );
  AOI22_X1 U19172 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19138), .B1(n16234), 
        .B2(n18907), .ZN(n16198) );
  NAND2_X1 U19173 ( .A1(n16187), .A2(n16188), .ZN(n16193) );
  INV_X1 U19174 ( .A(n16189), .ZN(n16190) );
  NOR2_X1 U19175 ( .A1(n16191), .A2(n16190), .ZN(n16192) );
  XNOR2_X1 U19176 ( .A(n16193), .B(n16192), .ZN(n16265) );
  INV_X1 U19177 ( .A(n16265), .ZN(n16196) );
  AOI21_X1 U19178 ( .B1(n16212), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16194) );
  NOR2_X1 U19179 ( .A1(n16195), .A2(n16194), .ZN(n16262) );
  AOI222_X1 U19180 ( .A1(n16196), .A2(n10996), .B1(n19146), .B2(n18905), .C1(
        n16228), .C2(n16262), .ZN(n16197) );
  OAI211_X1 U19181 ( .C1(n16199), .C2(n16243), .A(n16198), .B(n16197), .ZN(
        P2_U3003) );
  AOI22_X1 U19182 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n19137), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n16261), .ZN(n16210) );
  XNOR2_X1 U19183 ( .A(n16212), .B(n16268), .ZN(n16276) );
  INV_X1 U19184 ( .A(n16276), .ZN(n16206) );
  INV_X1 U19185 ( .A(n16200), .ZN(n16201) );
  NOR2_X1 U19186 ( .A1(n15629), .A2(n16201), .ZN(n16205) );
  NAND2_X1 U19187 ( .A1(n16203), .A2(n16202), .ZN(n16204) );
  XNOR2_X1 U19188 ( .A(n16205), .B(n16204), .ZN(n16279) );
  OAI22_X1 U19189 ( .A1(n16206), .A2(n19140), .B1(n16279), .B2(n19142), .ZN(
        n16207) );
  AOI21_X1 U19190 ( .B1(n19146), .B2(n16208), .A(n16207), .ZN(n16209) );
  OAI211_X1 U19191 ( .C1(n19150), .C2(n16211), .A(n16210), .B(n16209), .ZN(
        P2_U3004) );
  AOI22_X1 U19192 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19138), .B1(n16234), 
        .B2(n18915), .ZN(n16218) );
  NOR2_X1 U19193 ( .A1(n18920), .A2(n19157), .ZN(n16215) );
  NOR3_X1 U19194 ( .A1(n16213), .A2(n16212), .A3(n19140), .ZN(n16214) );
  AOI211_X1 U19195 ( .C1(n10996), .C2(n16216), .A(n16215), .B(n16214), .ZN(
        n16217) );
  OAI211_X1 U19196 ( .C1(n16219), .C2(n16243), .A(n16218), .B(n16217), .ZN(
        P2_U3005) );
  AOI22_X1 U19197 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n16261), .B1(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19137), .ZN(n16232) );
  INV_X1 U19198 ( .A(n16220), .ZN(n16284) );
  XOR2_X1 U19199 ( .A(n9837), .B(n16222), .Z(n16286) );
  INV_X1 U19200 ( .A(n16224), .ZN(n16226) );
  NOR2_X1 U19201 ( .A1(n16226), .A2(n16225), .ZN(n16227) );
  XNOR2_X1 U19202 ( .A(n16223), .B(n16227), .ZN(n16282) );
  AOI22_X1 U19203 ( .A1(n16286), .A2(n16228), .B1(n10996), .B2(n16282), .ZN(
        n16229) );
  INV_X1 U19204 ( .A(n16229), .ZN(n16230) );
  AOI21_X1 U19205 ( .B1(n19146), .B2(n16284), .A(n16230), .ZN(n16231) );
  OAI211_X1 U19206 ( .C1(n19150), .C2(n16233), .A(n16232), .B(n16231), .ZN(
        P2_U3006) );
  AOI22_X1 U19207 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19138), .B1(n16234), 
        .B2(n18956), .ZN(n16242) );
  NAND2_X1 U19208 ( .A1(n16235), .A2(n19146), .ZN(n16238) );
  OR2_X1 U19209 ( .A1(n16236), .A2(n19140), .ZN(n16237) );
  OAI211_X1 U19210 ( .C1(n16239), .C2(n19142), .A(n16238), .B(n16237), .ZN(
        n16240) );
  INV_X1 U19211 ( .A(n16240), .ZN(n16241) );
  OAI211_X1 U19212 ( .C1(n18964), .C2(n16243), .A(n16242), .B(n16241), .ZN(
        P2_U3009) );
  NAND2_X1 U19213 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n16261), .ZN(n16244) );
  OAI221_X1 U19214 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16246), 
        .C1(n16176), .C2(n16245), .A(n16244), .ZN(n16250) );
  OAI22_X1 U19215 ( .A1(n16248), .A2(n16272), .B1(n16271), .B2(n16247), .ZN(
        n16249) );
  AOI211_X1 U19216 ( .C1(n16251), .C2(n11843), .A(n16250), .B(n16249), .ZN(
        n16252) );
  OAI21_X1 U19217 ( .B1(n16253), .B2(n16278), .A(n16252), .ZN(P2_U3034) );
  NAND2_X1 U19218 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16254), .ZN(
        n16269) );
  AOI211_X1 U19219 ( .C1(n16268), .C2(n11037), .A(n16255), .B(n16269), .ZN(
        n16260) );
  OAI21_X1 U19220 ( .B1(n16258), .B2(n16257), .A(n16256), .ZN(n16267) );
  OAI22_X1 U19221 ( .A1(n16267), .A2(n11037), .B1(n16271), .B2(n18901), .ZN(
        n16259) );
  AOI211_X1 U19222 ( .C1(n16261), .C2(P2_REIP_REG_11__SCAN_IN), .A(n16260), 
        .B(n16259), .ZN(n16264) );
  AOI22_X1 U19223 ( .A1(n16262), .A2(n11843), .B1(n16285), .B2(n18905), .ZN(
        n16263) );
  OAI211_X1 U19224 ( .C1(n16265), .C2(n16278), .A(n16264), .B(n16263), .ZN(
        P2_U3035) );
  NAND2_X1 U19225 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n19138), .ZN(n16266) );
  OAI221_X1 U19226 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16269), 
        .C1(n16268), .C2(n16267), .A(n16266), .ZN(n16275) );
  OAI22_X1 U19227 ( .A1(n16273), .A2(n16272), .B1(n16271), .B2(n16270), .ZN(
        n16274) );
  AOI211_X1 U19228 ( .C1(n16276), .C2(n11843), .A(n16275), .B(n16274), .ZN(
        n16277) );
  OAI21_X1 U19229 ( .B1(n16279), .B2(n16278), .A(n16277), .ZN(P2_U3036) );
  AOI22_X1 U19230 ( .A1(n16281), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n16280), .B2(n19005), .ZN(n16292) );
  AOI222_X1 U19231 ( .A1(n16286), .A2(n11843), .B1(n16285), .B2(n16284), .C1(
        n16283), .C2(n16282), .ZN(n16291) );
  NAND2_X1 U19232 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19138), .ZN(n16290) );
  OAI211_X1 U19233 ( .C1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n16288), .B(n16287), .ZN(n16289) );
  NAND4_X1 U19234 ( .A1(n16292), .A2(n16291), .A3(n16290), .A4(n16289), .ZN(
        P2_U3038) );
  INV_X1 U19235 ( .A(n16315), .ZN(n16298) );
  NAND2_X1 U19236 ( .A1(n16298), .A2(n16293), .ZN(n16294) );
  OAI21_X1 U19237 ( .B1(n16295), .B2(n16298), .A(n16294), .ZN(n16318) );
  NAND2_X1 U19238 ( .A1(n16298), .A2(n16296), .ZN(n16297) );
  OAI21_X1 U19239 ( .B1(n16304), .B2(n16298), .A(n16297), .ZN(n16317) );
  OR2_X1 U19240 ( .A1(n16317), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n16305) );
  INV_X1 U19241 ( .A(n16300), .ZN(n16302) );
  OAI22_X1 U19242 ( .A1(n16300), .A2(n19831), .B1(n19841), .B2(n16299), .ZN(
        n16301) );
  OAI21_X1 U19243 ( .B1(n16302), .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n16301), .ZN(n16303) );
  OAI211_X1 U19244 ( .C1(n19822), .C2(n16304), .A(n16303), .B(n16315), .ZN(
        n16306) );
  AND3_X1 U19245 ( .A1(n16318), .A2(n16305), .A3(n16306), .ZN(n16307) );
  OAI22_X1 U19246 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n16307), .B1(
        n16318), .B2(n16306), .ZN(n16326) );
  INV_X1 U19247 ( .A(n16308), .ZN(n16310) );
  AOI22_X1 U19248 ( .A1(n16313), .A2(n16310), .B1(n11216), .B2(n16309), .ZN(
        n16311) );
  OAI21_X1 U19249 ( .B1(n16313), .B2(n16312), .A(n16311), .ZN(n19847) );
  OAI21_X1 U19250 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n16314), .ZN(n16323) );
  OAI22_X1 U19251 ( .A1(n16318), .A2(n16317), .B1(n16316), .B2(n16315), .ZN(
        n16320) );
  AOI211_X1 U19252 ( .C1(n16321), .C2(n19860), .A(n16320), .B(n16319), .ZN(
        n16322) );
  NAND2_X1 U19253 ( .A1(n16323), .A2(n16322), .ZN(n16324) );
  AOI211_X1 U19254 ( .C1(n16326), .C2(n16325), .A(n19847), .B(n16324), .ZN(
        n16342) );
  AOI211_X1 U19255 ( .C1(n16330), .C2(n16329), .A(n16328), .B(n16327), .ZN(
        n16340) );
  AOI22_X1 U19256 ( .A1(n16334), .A2(n16333), .B1(n19731), .B2(n16336), .ZN(
        n16338) );
  AND2_X1 U19257 ( .A1(n16342), .A2(n16335), .ZN(n16337) );
  OAI21_X1 U19258 ( .B1(n16337), .B2(n19859), .A(n16336), .ZN(n19729) );
  NAND2_X1 U19259 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19729), .ZN(n16343) );
  OAI21_X1 U19260 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n16338), .A(n16343), 
        .ZN(n16339) );
  OAI211_X1 U19261 ( .C1(n16342), .C2(n16341), .A(n16340), .B(n16339), .ZN(
        P2_U3176) );
  INV_X1 U19262 ( .A(n16343), .ZN(n16345) );
  INV_X1 U19263 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20990) );
  OAI21_X1 U19264 ( .B1(n16345), .B2(n20990), .A(n16344), .ZN(P2_U3593) );
  OAI22_X2 U19265 ( .A1(n18008), .A2(n17822), .B1(n17725), .B2(n17723), .ZN(
        n17713) );
  NOR2_X1 U19266 ( .A1(n16375), .A2(n17625), .ZN(n17488) );
  INV_X1 U19267 ( .A(n17725), .ZN(n17685) );
  NAND2_X1 U19268 ( .A1(n17685), .A2(n16346), .ZN(n16374) );
  NAND2_X1 U19269 ( .A1(n17806), .A2(n16347), .ZN(n16366) );
  AOI21_X1 U19270 ( .B1(n16374), .B2(n16366), .A(n16348), .ZN(n16355) );
  OAI21_X1 U19271 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16360), .A(
        n16349), .ZN(n16534) );
  AOI21_X1 U19272 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16351), .A(
        n16350), .ZN(n16353) );
  OAI211_X1 U19273 ( .C1(n17667), .C2(n16534), .A(n16353), .B(n16352), .ZN(
        n16354) );
  AOI211_X1 U19274 ( .C1(n16356), .C2(n17488), .A(n16355), .B(n16354), .ZN(
        n16357) );
  OAI21_X1 U19275 ( .B1(n17726), .B2(n16358), .A(n16357), .ZN(P3_U2800) );
  INV_X1 U19276 ( .A(n17464), .ZN(n17826) );
  NOR2_X1 U19277 ( .A1(n17826), .A2(n16364), .ZN(n16384) );
  NOR2_X1 U19278 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16384), .ZN(
        n16373) );
  INV_X1 U19279 ( .A(n16359), .ZN(n16371) );
  AOI21_X1 U19280 ( .B1(n16552), .B2(n16517), .A(n16360), .ZN(n16546) );
  OAI21_X1 U19281 ( .B1(n17573), .B2(n17655), .A(n16546), .ZN(n16361) );
  OAI211_X1 U19282 ( .C1(n16363), .C2(n16552), .A(n16362), .B(n16361), .ZN(
        n16369) );
  INV_X1 U19283 ( .A(n17463), .ZN(n17827) );
  NOR2_X1 U19284 ( .A1(n16364), .A2(n17827), .ZN(n16377) );
  NOR2_X1 U19285 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16377), .ZN(
        n16367) );
  OAI22_X1 U19286 ( .A1(n16367), .A2(n16366), .B1(n17726), .B2(n16365), .ZN(
        n16368) );
  AOI211_X1 U19287 ( .C1(n16371), .C2(n16370), .A(n16369), .B(n16368), .ZN(
        n16372) );
  OAI21_X1 U19288 ( .B1(n16374), .B2(n16373), .A(n16372), .ZN(P3_U2801) );
  NOR3_X1 U19289 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n20889), .A3(
        n16375), .ZN(n17459) );
  AOI22_X1 U19290 ( .A1(n18126), .A2(P3_REIP_REG_28__SCAN_IN), .B1(n17919), 
        .B2(n17459), .ZN(n16392) );
  OAI211_X1 U19291 ( .C1(n16377), .C2(n18787), .A(n16376), .B(n18121), .ZN(
        n16386) );
  INV_X1 U19292 ( .A(n16378), .ZN(n16379) );
  NOR2_X1 U19293 ( .A1(n16380), .A2(n16379), .ZN(n17477) );
  AOI21_X1 U19294 ( .B1(n17483), .B2(n17724), .A(n16388), .ZN(n16387) );
  INV_X1 U19295 ( .A(n16387), .ZN(n17476) );
  NAND2_X1 U19296 ( .A1(n17477), .A2(n17476), .ZN(n17475) );
  OAI21_X1 U19297 ( .B1(n17483), .B2(n16381), .A(n17475), .ZN(n16382) );
  AOI221_X1 U19298 ( .B1(n17321), .B2(n16384), .C1(n16383), .C2(n16382), .A(
        n18785), .ZN(n16385) );
  OAI211_X1 U19299 ( .C1(n16386), .C2(n16385), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18138), .ZN(n16391) );
  NAND4_X1 U19300 ( .A1(n17724), .A2(n18135), .A3(n16387), .A4(n17465), .ZN(
        n16390) );
  INV_X1 U19301 ( .A(n16388), .ZN(n17484) );
  OR3_X1 U19302 ( .A1(n18045), .A2(n17484), .A3(n17477), .ZN(n16389) );
  NAND4_X1 U19303 ( .A1(n16392), .A2(n16391), .A3(n16390), .A4(n16389), .ZN(
        P3_U2834) );
  NOR3_X1 U19304 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16394) );
  NOR4_X1 U19305 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16393) );
  NAND4_X1 U19306 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16394), .A3(n16393), .A4(
        U215), .ZN(U213) );
  INV_X1 U19307 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19064) );
  NAND2_X1 U19308 ( .A1(n19156), .A2(n16395), .ZN(n16396) );
  NAND2_X1 U19309 ( .A1(U214), .A2(n16396), .ZN(n16434) );
  INV_X1 U19310 ( .A(n16434), .ZN(n16445) );
  INV_X1 U19311 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16476) );
  OAI222_X1 U19312 ( .A1(U212), .A2(n19064), .B1(n16442), .B2(n19197), .C1(
        U214), .C2(n16476), .ZN(U216) );
  INV_X2 U19313 ( .A(U214), .ZN(n16444) );
  AOI222_X1 U19314 ( .A1(n16436), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n16445), 
        .B2(BUF1_REG_30__SCAN_IN), .C1(n16444), .C2(P1_DATAO_REG_30__SCAN_IN), 
        .ZN(n16397) );
  INV_X1 U19315 ( .A(n16397), .ZN(U217) );
  INV_X1 U19316 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16399) );
  AOI22_X1 U19317 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16444), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16436), .ZN(n16398) );
  OAI21_X1 U19318 ( .B1(n16399), .B2(n16442), .A(n16398), .ZN(U218) );
  INV_X1 U19319 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n16473) );
  INV_X1 U19320 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16400) );
  INV_X1 U19321 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n21093) );
  OAI222_X1 U19322 ( .A1(U212), .A2(n16473), .B1(n16442), .B2(n16400), .C1(
        U214), .C2(n21093), .ZN(U219) );
  INV_X1 U19323 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n19179) );
  AOI22_X1 U19324 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16444), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16436), .ZN(n16401) );
  OAI21_X1 U19325 ( .B1(n19179), .B2(n16442), .A(n16401), .ZN(U220) );
  INV_X1 U19326 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16403) );
  AOI22_X1 U19327 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16444), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16436), .ZN(n16402) );
  OAI21_X1 U19328 ( .B1(n16403), .B2(n16442), .A(n16402), .ZN(U221) );
  INV_X1 U19329 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16405) );
  AOI22_X1 U19330 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16444), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16436), .ZN(n16404) );
  OAI21_X1 U19331 ( .B1(n16405), .B2(n16442), .A(n16404), .ZN(U222) );
  INV_X1 U19332 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16407) );
  AOI22_X1 U19333 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16444), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16436), .ZN(n16406) );
  OAI21_X1 U19334 ( .B1(n16407), .B2(n16442), .A(n16406), .ZN(U223) );
  AOI22_X1 U19335 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16444), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16436), .ZN(n16408) );
  OAI21_X1 U19336 ( .B1(n14799), .B2(n16442), .A(n16408), .ZN(U224) );
  AOI22_X1 U19337 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16444), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16436), .ZN(n16409) );
  OAI21_X1 U19338 ( .B1(n15302), .B2(n16442), .A(n16409), .ZN(U225) );
  AOI22_X1 U19339 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16444), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16436), .ZN(n16410) );
  OAI21_X1 U19340 ( .B1(n15308), .B2(n16442), .A(n16410), .ZN(U226) );
  AOI22_X1 U19341 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16444), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16436), .ZN(n16411) );
  OAI21_X1 U19342 ( .B1(n15318), .B2(n16442), .A(n16411), .ZN(U227) );
  AOI22_X1 U19343 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16444), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16436), .ZN(n16412) );
  OAI21_X1 U19344 ( .B1(n15326), .B2(n16442), .A(n16412), .ZN(U228) );
  AOI22_X1 U19345 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16444), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16436), .ZN(n16413) );
  OAI21_X1 U19346 ( .B1(n15334), .B2(n16442), .A(n16413), .ZN(U229) );
  AOI22_X1 U19347 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16444), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16436), .ZN(n16414) );
  OAI21_X1 U19348 ( .B1(n15341), .B2(n16434), .A(n16414), .ZN(U230) );
  AOI222_X1 U19349 ( .A1(n16436), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n16445), 
        .B2(BUF1_REG_16__SCAN_IN), .C1(n16444), .C2(P1_DATAO_REG_16__SCAN_IN), 
        .ZN(n16415) );
  INV_X1 U19350 ( .A(n16415), .ZN(U231) );
  INV_X1 U19351 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n16417) );
  AOI22_X1 U19352 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16444), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16436), .ZN(n16416) );
  OAI21_X1 U19353 ( .B1(n16417), .B2(n16434), .A(n16416), .ZN(U232) );
  AOI22_X1 U19354 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16444), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16436), .ZN(n16418) );
  OAI21_X1 U19355 ( .B1(n14556), .B2(n16434), .A(n16418), .ZN(U233) );
  INV_X1 U19356 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16420) );
  AOI22_X1 U19357 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16444), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16436), .ZN(n16419) );
  OAI21_X1 U19358 ( .B1(n16420), .B2(n16434), .A(n16419), .ZN(U234) );
  INV_X1 U19359 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16422) );
  AOI22_X1 U19360 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16444), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16436), .ZN(n16421) );
  OAI21_X1 U19361 ( .B1(n16422), .B2(n16434), .A(n16421), .ZN(U235) );
  INV_X1 U19362 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n16424) );
  AOI22_X1 U19363 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16444), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16436), .ZN(n16423) );
  OAI21_X1 U19364 ( .B1(n16424), .B2(n16434), .A(n16423), .ZN(U236) );
  INV_X1 U19365 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16426) );
  AOI22_X1 U19366 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16444), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16436), .ZN(n16425) );
  OAI21_X1 U19367 ( .B1(n16426), .B2(n16434), .A(n16425), .ZN(U237) );
  INV_X1 U19368 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16428) );
  AOI22_X1 U19369 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16444), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16436), .ZN(n16427) );
  OAI21_X1 U19370 ( .B1(n16428), .B2(n16434), .A(n16427), .ZN(U238) );
  AOI22_X1 U19371 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16444), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16436), .ZN(n16429) );
  OAI21_X1 U19372 ( .B1(n16430), .B2(n16434), .A(n16429), .ZN(U239) );
  INV_X1 U19373 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16432) );
  AOI22_X1 U19374 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16444), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16436), .ZN(n16431) );
  OAI21_X1 U19375 ( .B1(n16432), .B2(n16434), .A(n16431), .ZN(U240) );
  INV_X1 U19376 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16435) );
  AOI22_X1 U19377 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16444), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16436), .ZN(n16433) );
  OAI21_X1 U19378 ( .B1(n16435), .B2(n16434), .A(n16433), .ZN(U241) );
  INV_X1 U19379 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n20913) );
  AOI22_X1 U19380 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16445), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16436), .ZN(n16437) );
  OAI21_X1 U19381 ( .B1(n20913), .B2(U214), .A(n16437), .ZN(U242) );
  INV_X1 U19382 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16450) );
  AOI22_X1 U19383 ( .A1(BUF1_REG_4__SCAN_IN), .A2(n16445), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n16444), .ZN(n16438) );
  OAI21_X1 U19384 ( .B1(n16450), .B2(U212), .A(n16438), .ZN(U243) );
  INV_X1 U19385 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n21040) );
  INV_X1 U19386 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16439) );
  INV_X1 U19387 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n21122) );
  OAI222_X1 U19388 ( .A1(U212), .A2(n21040), .B1(n16442), .B2(n16439), .C1(
        U214), .C2(n21122), .ZN(U244) );
  INV_X1 U19389 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16449) );
  AOI22_X1 U19390 ( .A1(BUF1_REG_2__SCAN_IN), .A2(n16445), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n16444), .ZN(n16440) );
  OAI21_X1 U19391 ( .B1(n16449), .B2(U212), .A(n16440), .ZN(U245) );
  INV_X1 U19392 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16443) );
  AOI22_X1 U19393 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16444), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16436), .ZN(n16441) );
  OAI21_X1 U19394 ( .B1(n16443), .B2(n16442), .A(n16441), .ZN(U246) );
  INV_X1 U19395 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n16447) );
  AOI22_X1 U19396 ( .A1(BUF1_REG_0__SCAN_IN), .A2(n16445), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n16444), .ZN(n16446) );
  OAI21_X1 U19397 ( .B1(n16447), .B2(U212), .A(n16446), .ZN(U247) );
  INV_X1 U19398 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18155) );
  AOI22_X1 U19399 ( .A1(n21215), .A2(n16447), .B1(n18155), .B2(U215), .ZN(U251) );
  OAI22_X1 U19400 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n21215), .ZN(n16448) );
  INV_X1 U19401 ( .A(n16448), .ZN(U252) );
  INV_X1 U19402 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18166) );
  AOI22_X1 U19403 ( .A1(n21215), .A2(n16449), .B1(n18166), .B2(U215), .ZN(U253) );
  INV_X1 U19404 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18170) );
  AOI22_X1 U19405 ( .A1(n21215), .A2(n21040), .B1(n18170), .B2(U215), .ZN(U254) );
  INV_X1 U19406 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18174) );
  AOI22_X1 U19407 ( .A1(n21215), .A2(n16450), .B1(n18174), .B2(U215), .ZN(U255) );
  INV_X1 U19408 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16451) );
  INV_X1 U19409 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n21103) );
  AOI22_X1 U19410 ( .A1(n21215), .A2(n16451), .B1(n21103), .B2(U215), .ZN(U256) );
  INV_X1 U19411 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16452) );
  INV_X1 U19412 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18181) );
  AOI22_X1 U19413 ( .A1(n21215), .A2(n16452), .B1(n18181), .B2(U215), .ZN(U257) );
  INV_X1 U19414 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16453) );
  INV_X1 U19415 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18185) );
  AOI22_X1 U19416 ( .A1(n21215), .A2(n16453), .B1(n18185), .B2(U215), .ZN(U258) );
  INV_X1 U19417 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16455) );
  AOI22_X1 U19418 ( .A1(n21215), .A2(n16455), .B1(n16454), .B2(U215), .ZN(U259) );
  INV_X1 U19419 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16456) );
  INV_X1 U19420 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17314) );
  AOI22_X1 U19421 ( .A1(n21215), .A2(n16456), .B1(n17314), .B2(U215), .ZN(U260) );
  INV_X1 U19422 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16457) );
  INV_X1 U19423 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17305) );
  AOI22_X1 U19424 ( .A1(n21215), .A2(n16457), .B1(n17305), .B2(U215), .ZN(U262) );
  INV_X1 U19425 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16458) );
  INV_X1 U19426 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17300) );
  AOI22_X1 U19427 ( .A1(n21215), .A2(n16458), .B1(n17300), .B2(U215), .ZN(U263) );
  INV_X1 U19428 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16459) );
  INV_X1 U19429 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17296) );
  AOI22_X1 U19430 ( .A1(n21215), .A2(n16459), .B1(n17296), .B2(U215), .ZN(U264) );
  OAI22_X1 U19431 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n21215), .ZN(n16460) );
  INV_X1 U19432 ( .A(n16460), .ZN(U265) );
  OAI22_X1 U19433 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n21215), .ZN(n16461) );
  INV_X1 U19434 ( .A(n16461), .ZN(U266) );
  INV_X1 U19435 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n21188) );
  AOI22_X1 U19436 ( .A1(n21215), .A2(n21188), .B1(n14135), .B2(U215), .ZN(U267) );
  INV_X1 U19437 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n16462) );
  AOI22_X1 U19438 ( .A1(n21215), .A2(n16462), .B1(n15343), .B2(U215), .ZN(U268) );
  OAI22_X1 U19439 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n21215), .ZN(n16463) );
  INV_X1 U19440 ( .A(n16463), .ZN(U269) );
  OAI22_X1 U19441 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n21215), .ZN(n16464) );
  INV_X1 U19442 ( .A(n16464), .ZN(U270) );
  INV_X1 U19443 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n16465) );
  AOI22_X1 U19444 ( .A1(n21215), .A2(n16465), .B1(n15319), .B2(U215), .ZN(U271) );
  INV_X1 U19445 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n16466) );
  AOI22_X1 U19446 ( .A1(n21215), .A2(n16466), .B1(n15309), .B2(U215), .ZN(U272) );
  INV_X1 U19447 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n16467) );
  AOI22_X1 U19448 ( .A1(n21215), .A2(n16467), .B1(n15303), .B2(U215), .ZN(U273) );
  OAI22_X1 U19449 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n21215), .ZN(n16468) );
  INV_X1 U19450 ( .A(n16468), .ZN(U274) );
  OAI22_X1 U19451 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n21215), .ZN(n16469) );
  INV_X1 U19452 ( .A(n16469), .ZN(U275) );
  OAI22_X1 U19453 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n21215), .ZN(n16470) );
  INV_X1 U19454 ( .A(n16470), .ZN(U276) );
  OAI22_X1 U19455 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n21215), .ZN(n16471) );
  INV_X1 U19456 ( .A(n16471), .ZN(U277) );
  INV_X1 U19457 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n16472) );
  INV_X1 U19458 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n19178) );
  AOI22_X1 U19459 ( .A1(n21215), .A2(n16472), .B1(n19178), .B2(U215), .ZN(U278) );
  INV_X1 U19460 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n21025) );
  AOI22_X1 U19461 ( .A1(n21215), .A2(n16473), .B1(n21025), .B2(U215), .ZN(U279) );
  INV_X1 U19462 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n16474) );
  INV_X1 U19463 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n17212) );
  AOI22_X1 U19464 ( .A1(n21215), .A2(n16474), .B1(n17212), .B2(U215), .ZN(U280) );
  INV_X1 U19465 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n19067) );
  INV_X1 U19466 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n17202) );
  AOI22_X1 U19467 ( .A1(n21215), .A2(n19067), .B1(n17202), .B2(U215), .ZN(U281) );
  INV_X1 U19468 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n20974) );
  AOI22_X1 U19469 ( .A1(n21215), .A2(n19064), .B1(n20974), .B2(U215), .ZN(U282) );
  INV_X1 U19470 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16475) );
  AOI222_X1 U19471 ( .A1(n16476), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16475), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .C1(n19064), .C2(
        P2_DATAO_REG_30__SCAN_IN), .ZN(n16477) );
  INV_X2 U19472 ( .A(n16479), .ZN(n16478) );
  INV_X1 U19473 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18692) );
  INV_X1 U19474 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19766) );
  AOI22_X1 U19475 ( .A1(n16478), .A2(n18692), .B1(n19766), .B2(n16479), .ZN(
        U347) );
  INV_X1 U19476 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18690) );
  INV_X1 U19477 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19765) );
  AOI22_X1 U19478 ( .A1(n16478), .A2(n18690), .B1(n19765), .B2(n16479), .ZN(
        U348) );
  INV_X1 U19479 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18688) );
  INV_X1 U19480 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19764) );
  AOI22_X1 U19481 ( .A1(n16478), .A2(n18688), .B1(n19764), .B2(n16479), .ZN(
        U349) );
  INV_X1 U19482 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18687) );
  INV_X1 U19483 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19763) );
  AOI22_X1 U19484 ( .A1(n16478), .A2(n18687), .B1(n19763), .B2(n16479), .ZN(
        U350) );
  INV_X1 U19485 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18685) );
  INV_X1 U19486 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19761) );
  AOI22_X1 U19487 ( .A1(n16478), .A2(n18685), .B1(n19761), .B2(n16479), .ZN(
        U351) );
  INV_X1 U19488 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18684) );
  INV_X1 U19489 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19759) );
  AOI22_X1 U19490 ( .A1(n16478), .A2(n18684), .B1(n19759), .B2(n16479), .ZN(
        U352) );
  INV_X1 U19491 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18682) );
  INV_X1 U19492 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n21027) );
  AOI22_X1 U19493 ( .A1(n16478), .A2(n18682), .B1(n21027), .B2(n16479), .ZN(
        U353) );
  INV_X1 U19494 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n21038) );
  AOI22_X1 U19495 ( .A1(n16478), .A2(n21038), .B1(n19757), .B2(n16479), .ZN(
        U354) );
  INV_X1 U19496 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18730) );
  AOI22_X1 U19497 ( .A1(n16478), .A2(n18730), .B1(n19795), .B2(n16479), .ZN(
        U355) );
  INV_X1 U19498 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18728) );
  INV_X1 U19499 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20955) );
  AOI22_X1 U19500 ( .A1(n16478), .A2(n18728), .B1(n20955), .B2(n16479), .ZN(
        U356) );
  INV_X1 U19501 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18725) );
  INV_X1 U19502 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19791) );
  AOI22_X1 U19503 ( .A1(n16478), .A2(n18725), .B1(n19791), .B2(n16479), .ZN(
        U357) );
  INV_X1 U19504 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18724) );
  INV_X1 U19505 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19789) );
  AOI22_X1 U19506 ( .A1(n16478), .A2(n18724), .B1(n19789), .B2(n16479), .ZN(
        U358) );
  INV_X1 U19507 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18722) );
  INV_X1 U19508 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19788) );
  AOI22_X1 U19509 ( .A1(n16478), .A2(n18722), .B1(n19788), .B2(n16479), .ZN(
        U359) );
  INV_X1 U19510 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18719) );
  INV_X1 U19511 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19787) );
  AOI22_X1 U19512 ( .A1(n16478), .A2(n18719), .B1(n19787), .B2(n16479), .ZN(
        U360) );
  INV_X1 U19513 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18717) );
  INV_X1 U19514 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19785) );
  AOI22_X1 U19515 ( .A1(n16478), .A2(n18717), .B1(n19785), .B2(n16479), .ZN(
        U361) );
  INV_X1 U19516 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18714) );
  INV_X1 U19517 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19784) );
  AOI22_X1 U19518 ( .A1(n16478), .A2(n18714), .B1(n19784), .B2(n16479), .ZN(
        U362) );
  INV_X1 U19519 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18713) );
  INV_X1 U19520 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19782) );
  AOI22_X1 U19521 ( .A1(n16478), .A2(n18713), .B1(n19782), .B2(n16479), .ZN(
        U363) );
  INV_X1 U19522 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18710) );
  INV_X1 U19523 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19780) );
  AOI22_X1 U19524 ( .A1(n16478), .A2(n18710), .B1(n19780), .B2(n16479), .ZN(
        U364) );
  INV_X1 U19525 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18679) );
  INV_X1 U19526 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19755) );
  AOI22_X1 U19527 ( .A1(n16478), .A2(n18679), .B1(n19755), .B2(n16479), .ZN(
        U365) );
  INV_X1 U19528 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18709) );
  INV_X1 U19529 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19778) );
  AOI22_X1 U19530 ( .A1(n16478), .A2(n18709), .B1(n19778), .B2(n16479), .ZN(
        U366) );
  INV_X1 U19531 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18706) );
  INV_X1 U19532 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19777) );
  AOI22_X1 U19533 ( .A1(n16478), .A2(n18706), .B1(n19777), .B2(n16479), .ZN(
        U367) );
  INV_X1 U19534 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18705) );
  INV_X1 U19535 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19775) );
  AOI22_X1 U19536 ( .A1(n16478), .A2(n18705), .B1(n19775), .B2(n16479), .ZN(
        U368) );
  INV_X1 U19537 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18703) );
  INV_X1 U19538 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19774) );
  AOI22_X1 U19539 ( .A1(n16478), .A2(n18703), .B1(n19774), .B2(n16479), .ZN(
        U369) );
  INV_X1 U19540 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18701) );
  INV_X1 U19541 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20935) );
  AOI22_X1 U19542 ( .A1(n16478), .A2(n18701), .B1(n20935), .B2(n16479), .ZN(
        U370) );
  INV_X1 U19543 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18700) );
  INV_X1 U19544 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19772) );
  AOI22_X1 U19545 ( .A1(n16478), .A2(n18700), .B1(n19772), .B2(n16479), .ZN(
        U371) );
  INV_X1 U19546 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18697) );
  INV_X1 U19547 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19771) );
  AOI22_X1 U19548 ( .A1(n16478), .A2(n18697), .B1(n19771), .B2(n16479), .ZN(
        U372) );
  INV_X1 U19549 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18695) );
  INV_X1 U19550 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19770) );
  AOI22_X1 U19551 ( .A1(n16478), .A2(n18695), .B1(n19770), .B2(n16479), .ZN(
        U373) );
  INV_X1 U19552 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18694) );
  INV_X1 U19553 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19769) );
  AOI22_X1 U19554 ( .A1(n16478), .A2(n18694), .B1(n19769), .B2(n16479), .ZN(
        U374) );
  INV_X1 U19555 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n20957) );
  INV_X1 U19556 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19768) );
  AOI22_X1 U19557 ( .A1(n16478), .A2(n20957), .B1(n19768), .B2(n16479), .ZN(
        U375) );
  INV_X1 U19558 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18678) );
  INV_X1 U19559 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19753) );
  AOI22_X1 U19560 ( .A1(n16478), .A2(n18678), .B1(n19753), .B2(n16479), .ZN(
        U376) );
  INV_X1 U19561 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16482) );
  NAND2_X1 U19562 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18677), .ZN(n16481) );
  NAND2_X1 U19563 ( .A1(n18674), .A2(n16480), .ZN(n18662) );
  OAI21_X1 U19564 ( .B1(n16481), .B2(n16480), .A(n18662), .ZN(n18745) );
  OAI21_X1 U19565 ( .B1(n18674), .B2(n16482), .A(n18742), .ZN(P3_U2633) );
  NOR2_X1 U19566 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18799), .ZN(n18656) );
  INV_X1 U19567 ( .A(n18656), .ZN(n16485) );
  NAND2_X1 U19568 ( .A1(n18809), .A2(n18748), .ZN(n16484) );
  OAI21_X1 U19569 ( .B1(n16490), .B2(n17391), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16483) );
  OAI21_X1 U19570 ( .B1(n16485), .B2(n16484), .A(n16483), .ZN(P3_U2634) );
  AOI21_X1 U19571 ( .B1(n18674), .B2(n18677), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16486) );
  AOI22_X1 U19572 ( .A1(n18739), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16486), 
        .B2(n18807), .ZN(P3_U2635) );
  INV_X1 U19573 ( .A(BS16), .ZN(n18822) );
  AOI21_X1 U19574 ( .B1(n16487), .B2(n18822), .A(n18742), .ZN(n18740) );
  INV_X1 U19575 ( .A(n18740), .ZN(n18743) );
  OAI21_X1 U19576 ( .B1(n18745), .B2(n16507), .A(n18743), .ZN(P3_U2636) );
  NOR3_X1 U19577 ( .A1(n16490), .A2(n16489), .A3(n16488), .ZN(n18634) );
  NOR2_X1 U19578 ( .A1(n18634), .A2(n18651), .ZN(n18793) );
  OAI21_X1 U19579 ( .B1(n18793), .B2(n18148), .A(n16491), .ZN(P3_U2637) );
  NOR4_X1 U19580 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_15__SCAN_IN), .A3(P3_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_20__SCAN_IN), .ZN(n16495) );
  NOR4_X1 U19581 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_11__SCAN_IN), .A3(P3_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_13__SCAN_IN), .ZN(n16494) );
  NOR4_X1 U19582 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_27__SCAN_IN), .A3(P3_DATAWIDTH_REG_28__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16493) );
  NOR4_X1 U19583 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_22__SCAN_IN), .A3(P3_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_24__SCAN_IN), .ZN(n16492) );
  NAND4_X1 U19584 ( .A1(n16495), .A2(n16494), .A3(n16493), .A4(n16492), .ZN(
        n16501) );
  NOR4_X1 U19585 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_19__SCAN_IN), .A3(P3_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_8__SCAN_IN), .ZN(n16499) );
  AOI211_X1 U19586 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_26__SCAN_IN), .B(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n16498) );
  NOR4_X1 U19587 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_6__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(n16497) );
  NOR4_X1 U19588 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_2__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_4__SCAN_IN), .ZN(n16496) );
  NAND4_X1 U19589 ( .A1(n16499), .A2(n16498), .A3(n16497), .A4(n16496), .ZN(
        n16500) );
  NOR2_X1 U19590 ( .A1(n16501), .A2(n16500), .ZN(n18783) );
  INV_X1 U19591 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18737) );
  NOR3_X1 U19592 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16503) );
  OAI21_X1 U19593 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16503), .A(n18783), .ZN(
        n16502) );
  OAI21_X1 U19594 ( .B1(n18783), .B2(n18737), .A(n16502), .ZN(P3_U2638) );
  INV_X1 U19595 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18776) );
  INV_X1 U19596 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18744) );
  AOI21_X1 U19597 ( .B1(n18776), .B2(n18744), .A(n16503), .ZN(n16504) );
  INV_X1 U19598 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18734) );
  INV_X1 U19599 ( .A(n18783), .ZN(n18778) );
  AOI22_X1 U19600 ( .A1(n18783), .A2(n16504), .B1(n18734), .B2(n18778), .ZN(
        P3_U2639) );
  NAND2_X1 U19601 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18795), .ZN(n16506) );
  AOI211_X4 U19602 ( .C1(n16507), .C2(n18803), .A(n16508), .B(n16506), .ZN(
        n16895) );
  NOR3_X1 U19603 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16869) );
  INV_X1 U19604 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17175) );
  NAND2_X1 U19605 ( .A1(n16869), .A2(n17175), .ZN(n16858) );
  NOR2_X1 U19606 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16858), .ZN(n16840) );
  INV_X1 U19607 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16831) );
  NAND2_X1 U19608 ( .A1(n16840), .A2(n16831), .ZN(n16830) );
  NAND2_X1 U19609 ( .A1(n16817), .A2(n16806), .ZN(n16805) );
  NAND2_X1 U19610 ( .A1(n16787), .A2(n16775), .ZN(n16773) );
  NAND2_X1 U19611 ( .A1(n16761), .A2(n16759), .ZN(n16756) );
  NAND2_X1 U19612 ( .A1(n16738), .A2(n16733), .ZN(n16732) );
  INV_X1 U19613 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16703) );
  NAND2_X1 U19614 ( .A1(n16709), .A2(n16703), .ZN(n16700) );
  NAND2_X1 U19615 ( .A1(n16684), .A2(n16675), .ZN(n16674) );
  INV_X1 U19616 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16655) );
  NAND2_X1 U19617 ( .A1(n16665), .A2(n16655), .ZN(n16654) );
  NAND2_X1 U19618 ( .A1(n16637), .A2(n16985), .ZN(n16633) );
  NOR2_X1 U19619 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16633), .ZN(n16619) );
  NAND2_X1 U19620 ( .A1(n16619), .A2(n16614), .ZN(n16613) );
  NOR2_X1 U19621 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16613), .ZN(n16599) );
  NAND2_X1 U19622 ( .A1(n16599), .A2(n16592), .ZN(n16591) );
  NOR2_X1 U19623 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16591), .ZN(n16575) );
  INV_X1 U19624 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16943) );
  NAND2_X1 U19625 ( .A1(n16575), .A2(n16943), .ZN(n16570) );
  NOR2_X1 U19626 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16570), .ZN(n16554) );
  INV_X1 U19627 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16930) );
  NAND2_X1 U19628 ( .A1(n16554), .A2(n16930), .ZN(n16533) );
  NOR2_X1 U19629 ( .A1(n16886), .A2(n16533), .ZN(n16539) );
  INV_X1 U19630 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16513) );
  INV_X1 U19631 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18731) );
  OAI211_X1 U19632 ( .C1(n18795), .C2(n18794), .A(n18803), .B(n16507), .ZN(
        n18645) );
  INV_X1 U19633 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18716) );
  INV_X1 U19634 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18712) );
  INV_X1 U19635 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18696) );
  INV_X1 U19636 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18698) );
  INV_X1 U19637 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n20924) );
  INV_X1 U19638 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18686) );
  INV_X1 U19639 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18683) );
  INV_X1 U19640 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n21028) );
  NOR2_X1 U19641 ( .A1(n21028), .A2(n18776), .ZN(n16868) );
  AND2_X1 U19642 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(n16868), .ZN(n16855) );
  NAND2_X1 U19643 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16855), .ZN(n16825) );
  NOR2_X1 U19644 ( .A1(n18683), .A2(n16825), .ZN(n16804) );
  NAND2_X1 U19645 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n16804), .ZN(n16801) );
  NOR2_X1 U19646 ( .A1(n18686), .A2(n16801), .ZN(n16796) );
  NAND2_X1 U19647 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16796), .ZN(n16795) );
  NAND2_X1 U19648 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n16760) );
  NOR3_X1 U19649 ( .A1(n20924), .A2(n16795), .A3(n16760), .ZN(n16745) );
  NAND2_X1 U19650 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16745), .ZN(n16717) );
  NOR3_X1 U19651 ( .A1(n18696), .A2(n18698), .A3(n16717), .ZN(n16683) );
  INV_X1 U19652 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18708) );
  INV_X1 U19653 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18702) );
  NAND2_X1 U19654 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16693) );
  NOR2_X1 U19655 ( .A1(n18702), .A2(n16693), .ZN(n16650) );
  NAND3_X1 U19656 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .A3(n16650), .ZN(n16636) );
  NOR2_X1 U19657 ( .A1(n18708), .A2(n16636), .ZN(n16626) );
  NAND3_X1 U19658 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n16683), .A3(n16626), 
        .ZN(n16620) );
  NOR2_X1 U19659 ( .A1(n18712), .A2(n16620), .ZN(n16606) );
  NAND2_X1 U19660 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16606), .ZN(n16596) );
  NOR2_X1 U19661 ( .A1(n18716), .A2(n16596), .ZN(n16573) );
  AND3_X1 U19662 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .A3(n16573), .ZN(n16514) );
  NAND4_X1 U19663 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16569), .ZN(n16516) );
  NOR3_X1 U19664 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18731), .A3(n16516), 
        .ZN(n16512) );
  NAND3_X1 U19665 ( .A1(n18799), .A2(n18809), .A3(n16507), .ZN(n18660) );
  NOR2_X1 U19666 ( .A1(n18140), .A2(n16874), .ZN(n16850) );
  INV_X1 U19667 ( .A(n18812), .ZN(n16846) );
  NOR2_X1 U19668 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18748), .ZN(n18654) );
  NAND2_X1 U19669 ( .A1(n18654), .A2(n18656), .ZN(n18649) );
  INV_X1 U19670 ( .A(n18645), .ZN(n16509) );
  AOI22_X1 U19671 ( .A1(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n16872), .B1(
        P3_EBX_REG_31__SCAN_IN), .B2(n16864), .ZN(n16510) );
  INV_X1 U19672 ( .A(n16510), .ZN(n16511) );
  AOI211_X1 U19673 ( .C1(n16539), .C2(n16513), .A(n16512), .B(n16511), .ZN(
        n16532) );
  NAND2_X1 U19674 ( .A1(n16514), .A2(n16897), .ZN(n16553) );
  NAND3_X1 U19675 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16515) );
  NAND2_X1 U19676 ( .A1(n16897), .A2(n16887), .ZN(n16894) );
  OAI21_X1 U19677 ( .B1(n16553), .B2(n16515), .A(n16894), .ZN(n16535) );
  INV_X1 U19678 ( .A(n16535), .ZN(n16549) );
  NOR2_X1 U19679 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16516), .ZN(n16538) );
  OAI21_X1 U19680 ( .B1(n16549), .B2(n16538), .A(P3_REIP_REG_31__SCAN_IN), 
        .ZN(n16531) );
  INV_X1 U19681 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17486) );
  INV_X1 U19682 ( .A(n16520), .ZN(n16519) );
  NOR2_X1 U19683 ( .A1(n17486), .A2(n16519), .ZN(n16518) );
  OAI21_X1 U19684 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16518), .A(
        n16517), .ZN(n17472) );
  INV_X1 U19685 ( .A(n17472), .ZN(n16557) );
  AOI21_X1 U19686 ( .B1(n17486), .B2(n16519), .A(n16518), .ZN(n17481) );
  NOR2_X1 U19687 ( .A1(n17812), .A2(n17505), .ZN(n16523) );
  INV_X1 U19688 ( .A(n16523), .ZN(n16522) );
  OR2_X1 U19689 ( .A1(n17506), .A2(n16522), .ZN(n17462) );
  AOI21_X1 U19690 ( .B1(n9960), .B2(n17462), .A(n16520), .ZN(n17495) );
  INV_X1 U19691 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17522) );
  NOR2_X1 U19692 ( .A1(n17522), .A2(n16522), .ZN(n16521) );
  OAI21_X1 U19693 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16521), .A(
        n17462), .ZN(n17508) );
  INV_X1 U19694 ( .A(n17508), .ZN(n16586) );
  AOI22_X1 U19695 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16522), .B1(
        n16523), .B2(n17522), .ZN(n17519) );
  INV_X1 U19696 ( .A(n17519), .ZN(n16598) );
  NAND2_X1 U19697 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17532), .ZN(
        n16524) );
  AOI21_X1 U19698 ( .B1(n9959), .B2(n16524), .A(n16523), .ZN(n17533) );
  INV_X1 U19699 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17559) );
  OR2_X1 U19700 ( .A1(n17812), .A2(n17548), .ZN(n16527) );
  NOR2_X1 U19701 ( .A1(n17559), .A2(n16527), .ZN(n16525) );
  OAI21_X1 U19702 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n16525), .A(
        n16524), .ZN(n16526) );
  INV_X1 U19703 ( .A(n16526), .ZN(n17547) );
  XNOR2_X1 U19704 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n16527), .ZN(
        n17556) );
  NOR2_X1 U19705 ( .A1(n17812), .A2(n17588), .ZN(n17579) );
  INV_X1 U19706 ( .A(n17579), .ZN(n16670) );
  NOR2_X1 U19707 ( .A1(n17589), .A2(n16670), .ZN(n17545) );
  OAI21_X1 U19708 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17545), .A(
        n16527), .ZN(n16528) );
  INV_X1 U19709 ( .A(n16528), .ZN(n17574) );
  NOR2_X1 U19710 ( .A1(n17812), .A2(n17618), .ZN(n17616) );
  NAND2_X1 U19711 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17616), .ZN(
        n16697) );
  NOR2_X1 U19712 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16697), .ZN(
        n16686) );
  NOR2_X1 U19713 ( .A1(n16598), .A2(n9875), .ZN(n16597) );
  NOR2_X1 U19714 ( .A1(n16576), .A2(n16853), .ZN(n16566) );
  NOR2_X1 U19715 ( .A1(n16546), .A2(n16545), .ZN(n16544) );
  NAND4_X1 U19716 ( .A1(n16837), .A2(n16874), .A3(n16544), .A4(n16534), .ZN(
        n16530) );
  NAND3_X1 U19717 ( .A1(n16532), .A2(n16531), .A3(n16530), .ZN(P3_U2640) );
  NAND2_X1 U19718 ( .A1(n16895), .A2(n16533), .ZN(n16542) );
  OAI22_X1 U19719 ( .A1(n16536), .A2(n16882), .B1(n18731), .B2(n16535), .ZN(
        n16537) );
  OAI21_X1 U19720 ( .B1(n16896), .B2(n16539), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16540) );
  NAND2_X1 U19721 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16561) );
  NOR2_X1 U19722 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16561), .ZN(n16541) );
  AOI22_X1 U19723 ( .A1(n16864), .A2(P3_EBX_REG_29__SCAN_IN), .B1(n16569), 
        .B2(n16541), .ZN(n16551) );
  INV_X1 U19724 ( .A(n16554), .ZN(n16543) );
  AOI21_X1 U19725 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n16543), .A(n16542), .ZN(
        n16548) );
  INV_X1 U19726 ( .A(n16874), .ZN(n18657) );
  AOI211_X1 U19727 ( .C1(n16546), .C2(n16545), .A(n16544), .B(n18657), .ZN(
        n16547) );
  AOI211_X1 U19728 ( .C1(n16549), .C2(P3_REIP_REG_29__SCAN_IN), .A(n16548), 
        .B(n16547), .ZN(n16550) );
  OAI211_X1 U19729 ( .C1(n16552), .C2(n16882), .A(n16551), .B(n16550), .ZN(
        P3_U2642) );
  AOI22_X1 U19730 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16872), .B1(
        n16864), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16564) );
  NAND2_X1 U19731 ( .A1(n16894), .A2(n16553), .ZN(n16582) );
  INV_X1 U19732 ( .A(n16582), .ZN(n16560) );
  AOI211_X1 U19733 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16570), .A(n16554), .B(
        n16886), .ZN(n16559) );
  AOI211_X1 U19734 ( .C1(n16557), .C2(n16556), .A(n16555), .B(n18657), .ZN(
        n16558) );
  AOI211_X1 U19735 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16560), .A(n16559), 
        .B(n16558), .ZN(n16563) );
  OAI211_X1 U19736 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16569), .B(n16561), .ZN(n16562) );
  NAND3_X1 U19737 ( .A1(n16564), .A2(n16563), .A3(n16562), .ZN(P3_U2643) );
  INV_X1 U19738 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18723) );
  AOI211_X1 U19739 ( .C1(n17481), .C2(n16566), .A(n16565), .B(n18657), .ZN(
        n16568) );
  OAI22_X1 U19740 ( .A1(n17486), .A2(n16882), .B1(n16893), .B2(n16943), .ZN(
        n16567) );
  AOI211_X1 U19741 ( .C1(n16569), .C2(n18723), .A(n16568), .B(n16567), .ZN(
        n16572) );
  OAI211_X1 U19742 ( .C1(n16575), .C2(n16943), .A(n16895), .B(n16570), .ZN(
        n16571) );
  OAI211_X1 U19743 ( .C1(n16582), .C2(n18723), .A(n16572), .B(n16571), .ZN(
        P3_U2644) );
  NAND2_X1 U19744 ( .A1(n16842), .A2(n16573), .ZN(n16595) );
  INV_X1 U19745 ( .A(n16595), .ZN(n16574) );
  AOI21_X1 U19746 ( .B1(P3_REIP_REG_25__SCAN_IN), .B2(n16574), .A(
        P3_REIP_REG_26__SCAN_IN), .ZN(n16583) );
  AOI22_X1 U19747 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n16872), .B1(
        n16864), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16581) );
  AOI211_X1 U19748 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16591), .A(n16575), .B(
        n16886), .ZN(n16579) );
  AOI211_X1 U19749 ( .C1(n17495), .C2(n16577), .A(n16576), .B(n18657), .ZN(
        n16578) );
  NOR2_X1 U19750 ( .A1(n16579), .A2(n16578), .ZN(n16580) );
  OAI211_X1 U19751 ( .C1(n16583), .C2(n16582), .A(n16581), .B(n16580), .ZN(
        P3_U2645) );
  INV_X1 U19752 ( .A(n16897), .ZN(n16881) );
  OAI21_X1 U19753 ( .B1(n16881), .B2(n16596), .A(n16894), .ZN(n16607) );
  OAI21_X1 U19754 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n16887), .A(n16607), 
        .ZN(n16590) );
  AOI211_X1 U19755 ( .C1(n16586), .C2(n16585), .A(n16584), .B(n18657), .ZN(
        n16589) );
  AOI22_X1 U19756 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n16872), .B1(
        n16864), .B2(P3_EBX_REG_25__SCAN_IN), .ZN(n16587) );
  INV_X1 U19757 ( .A(n16587), .ZN(n16588) );
  AOI211_X1 U19758 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n16590), .A(n16589), 
        .B(n16588), .ZN(n16594) );
  OAI211_X1 U19759 ( .C1(n16599), .C2(n16592), .A(n16895), .B(n16591), .ZN(
        n16593) );
  OAI211_X1 U19760 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n16595), .A(n16594), 
        .B(n16593), .ZN(P3_U2646) );
  AOI22_X1 U19761 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16872), .B1(
        n16864), .B2(P3_EBX_REG_24__SCAN_IN), .ZN(n16605) );
  NOR2_X1 U19762 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16887), .ZN(n16603) );
  INV_X1 U19763 ( .A(n16596), .ZN(n16602) );
  AOI211_X1 U19764 ( .C1(n16598), .C2(n9875), .A(n16597), .B(n18657), .ZN(
        n16601) );
  AOI211_X1 U19765 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16613), .A(n16599), .B(
        n16886), .ZN(n16600) );
  AOI211_X1 U19766 ( .C1(n16603), .C2(n16602), .A(n16601), .B(n16600), .ZN(
        n16604) );
  OAI211_X1 U19767 ( .C1(n18716), .C2(n16607), .A(n16605), .B(n16604), .ZN(
        P3_U2647) );
  AOI21_X1 U19768 ( .B1(n16606), .B2(n16842), .A(P3_REIP_REG_23__SCAN_IN), 
        .ZN(n16608) );
  NOR2_X1 U19769 ( .A1(n16608), .A2(n16607), .ZN(n16612) );
  AOI211_X1 U19770 ( .C1(n17533), .C2(n16610), .A(n16609), .B(n18657), .ZN(
        n16611) );
  AOI211_X1 U19771 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n16864), .A(n16612), .B(
        n16611), .ZN(n16616) );
  OAI211_X1 U19772 ( .C1(n16619), .C2(n16614), .A(n16895), .B(n16613), .ZN(
        n16615) );
  OAI211_X1 U19773 ( .C1(n16882), .C2(n9959), .A(n16616), .B(n16615), .ZN(
        P3_U2648) );
  AOI21_X1 U19774 ( .B1(n16842), .B2(n16620), .A(n16881), .ZN(n16627) );
  AOI22_X1 U19775 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n16872), .B1(
        n16864), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n16625) );
  AOI211_X1 U19776 ( .C1(n17547), .C2(n16618), .A(n16617), .B(n18657), .ZN(
        n16623) );
  AOI211_X1 U19777 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16633), .A(n16619), .B(
        n16886), .ZN(n16622) );
  NOR3_X1 U19778 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16887), .A3(n16620), 
        .ZN(n16621) );
  NOR3_X1 U19779 ( .A1(n16623), .A2(n16622), .A3(n16621), .ZN(n16624) );
  OAI211_X1 U19780 ( .C1(n18712), .C2(n16627), .A(n16625), .B(n16624), .ZN(
        P3_U2649) );
  INV_X1 U19781 ( .A(n16626), .ZN(n16628) );
  INV_X1 U19782 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18711) );
  NAND2_X1 U19783 ( .A1(n16842), .A2(n16683), .ZN(n16708) );
  AOI221_X1 U19784 ( .B1(n16628), .B2(n18711), .C1(n16708), .C2(n18711), .A(
        n16627), .ZN(n16632) );
  AOI211_X1 U19785 ( .C1(n17556), .C2(n16630), .A(n16629), .B(n18657), .ZN(
        n16631) );
  AOI211_X1 U19786 ( .C1(n16872), .C2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n16632), .B(n16631), .ZN(n16635) );
  OAI211_X1 U19787 ( .C1(n16637), .C2(n16985), .A(n16895), .B(n16633), .ZN(
        n16634) );
  OAI211_X1 U19788 ( .C1(n16985), .C2(n16893), .A(n16635), .B(n16634), .ZN(
        P3_U2650) );
  NOR3_X1 U19789 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16636), .A3(n16708), 
        .ZN(n16639) );
  AOI211_X1 U19790 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16654), .A(n16637), .B(
        n16886), .ZN(n16638) );
  AOI211_X1 U19791 ( .C1(n16872), .C2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16639), .B(n16638), .ZN(n16644) );
  INV_X1 U19792 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18704) );
  NAND3_X1 U19793 ( .A1(n16683), .A2(n16650), .A3(n16897), .ZN(n16679) );
  NOR2_X1 U19794 ( .A1(n18704), .A2(n16679), .ZN(n16648) );
  INV_X1 U19795 ( .A(n16894), .ZN(n16649) );
  AOI211_X1 U19796 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(n16648), .A(n16649), 
        .B(n18708), .ZN(n16642) );
  AOI211_X1 U19797 ( .C1(n17574), .C2(n16647), .A(n16640), .B(n18657), .ZN(
        n16641) );
  AOI211_X1 U19798 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16864), .A(n16642), .B(
        n16641), .ZN(n16643) );
  NAND2_X1 U19799 ( .A1(n16644), .A2(n16643), .ZN(P3_U2651) );
  INV_X1 U19800 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16651) );
  NAND2_X1 U19801 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17579), .ZN(
        n16660) );
  AOI21_X1 U19802 ( .B1(n16651), .B2(n16660), .A(n17545), .ZN(n17580) );
  INV_X1 U19803 ( .A(n17580), .ZN(n16646) );
  INV_X1 U19804 ( .A(n16686), .ZN(n16659) );
  OAI21_X1 U19805 ( .B1(n16660), .B2(n16659), .A(n16837), .ZN(n16645) );
  AOI221_X1 U19806 ( .B1(n16647), .B2(n16646), .C1(n16645), .C2(n17580), .A(
        n18126), .ZN(n16658) );
  NOR2_X1 U19807 ( .A1(n16649), .A2(n16648), .ZN(n16662) );
  INV_X1 U19808 ( .A(n16708), .ZN(n16694) );
  NAND2_X1 U19809 ( .A1(n16650), .A2(n16694), .ZN(n16664) );
  NOR3_X1 U19810 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n18704), .A3(n16664), 
        .ZN(n16653) );
  OAI22_X1 U19811 ( .A1(n16651), .A2(n16882), .B1(n16893), .B2(n16655), .ZN(
        n16652) );
  AOI211_X1 U19812 ( .C1(n16662), .C2(P3_REIP_REG_19__SCAN_IN), .A(n16653), 
        .B(n16652), .ZN(n16657) );
  OAI211_X1 U19813 ( .C1(n16665), .C2(n16655), .A(n16895), .B(n16654), .ZN(
        n16656) );
  OAI211_X1 U19814 ( .C1(n16850), .C2(n16658), .A(n16657), .B(n16656), .ZN(
        P3_U2652) );
  INV_X1 U19815 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17596) );
  OAI21_X1 U19816 ( .B1(n16670), .B2(n16659), .A(n16837), .ZN(n16672) );
  OAI21_X1 U19817 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17579), .A(
        n16660), .ZN(n17593) );
  XOR2_X1 U19818 ( .A(n16672), .B(n17593), .Z(n16661) );
  AOI21_X1 U19819 ( .B1(n16661), .B2(n16874), .A(n18140), .ZN(n16669) );
  INV_X1 U19820 ( .A(n16662), .ZN(n16663) );
  AOI21_X1 U19821 ( .B1(n18704), .B2(n16664), .A(n16663), .ZN(n16667) );
  AOI211_X1 U19822 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16674), .A(n16665), .B(
        n16886), .ZN(n16666) );
  AOI211_X1 U19823 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16864), .A(n16667), .B(
        n16666), .ZN(n16668) );
  OAI211_X1 U19824 ( .C1(n17596), .C2(n16882), .A(n16669), .B(n16668), .ZN(
        P3_U2653) );
  AND2_X1 U19825 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17602), .ZN(
        n16685) );
  OAI21_X1 U19826 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16685), .A(
        n16670), .ZN(n17604) );
  AOI211_X1 U19827 ( .C1(n16685), .C2(n16686), .A(n16853), .B(n17604), .ZN(
        n16671) );
  AOI211_X1 U19828 ( .C1(n16672), .C2(n17604), .A(n16671), .B(n18657), .ZN(
        n16673) );
  AOI211_X1 U19829 ( .C1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .C2(n16872), .A(
        n18126), .B(n16673), .ZN(n16682) );
  NOR3_X1 U19830 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n16693), .A3(n16708), 
        .ZN(n16678) );
  OAI211_X1 U19831 ( .C1(n16675), .C2(n16684), .A(n16674), .B(n16895), .ZN(
        n16676) );
  INV_X1 U19832 ( .A(n16676), .ZN(n16677) );
  AOI211_X1 U19833 ( .C1(P3_EBX_REG_17__SCAN_IN), .C2(n16864), .A(n16678), .B(
        n16677), .ZN(n16681) );
  NAND3_X1 U19834 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n16894), .A3(n16679), 
        .ZN(n16680) );
  NAND3_X1 U19835 ( .A1(n16682), .A2(n16681), .A3(n16680), .ZN(P3_U2654) );
  NAND2_X1 U19836 ( .A1(n16683), .A2(n16897), .ZN(n16718) );
  NAND2_X1 U19837 ( .A1(n16894), .A2(n16718), .ZN(n16721) );
  INV_X1 U19838 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n20890) );
  AOI211_X1 U19839 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16700), .A(n16684), .B(
        n16886), .ZN(n16692) );
  INV_X1 U19840 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16690) );
  AOI21_X1 U19841 ( .B1(n16690), .B2(n16697), .A(n16685), .ZN(n17617) );
  NOR2_X1 U19842 ( .A1(n16686), .A2(n16853), .ZN(n16688) );
  INV_X1 U19843 ( .A(n17617), .ZN(n16687) );
  INV_X1 U19844 ( .A(n16688), .ZN(n16699) );
  OAI221_X1 U19845 ( .B1(n17617), .B2(n16688), .C1(n16687), .C2(n16699), .A(
        n16874), .ZN(n16689) );
  OAI211_X1 U19846 ( .C1(n16690), .C2(n16882), .A(n18138), .B(n16689), .ZN(
        n16691) );
  AOI211_X1 U19847 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16864), .A(n16692), .B(
        n16691), .ZN(n16696) );
  OAI211_X1 U19848 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(P3_REIP_REG_15__SCAN_IN), .A(n16694), .B(n16693), .ZN(n16695) );
  OAI211_X1 U19849 ( .C1(n16721), .C2(n20890), .A(n16696), .B(n16695), .ZN(
        P3_U2655) );
  INV_X1 U19850 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18699) );
  INV_X1 U19851 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17627) );
  INV_X1 U19852 ( .A(n17616), .ZN(n16710) );
  INV_X1 U19853 ( .A(n16697), .ZN(n16698) );
  AOI21_X1 U19854 ( .B1(n17627), .B2(n16710), .A(n16698), .ZN(n17630) );
  NOR3_X1 U19855 ( .A1(n17630), .A2(n18657), .A3(n16699), .ZN(n16706) );
  OAI211_X1 U19856 ( .C1(n16709), .C2(n16703), .A(n16895), .B(n16700), .ZN(
        n16701) );
  OAI21_X1 U19857 ( .B1(n16882), .B2(n17627), .A(n16701), .ZN(n16705) );
  NOR2_X1 U19858 ( .A1(n16837), .A2(n18657), .ZN(n16866) );
  AOI21_X1 U19859 ( .B1(n16837), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n18657), .ZN(n16889) );
  OAI211_X1 U19860 ( .C1(n17616), .C2(n16866), .A(n17630), .B(n16889), .ZN(
        n16702) );
  OAI211_X1 U19861 ( .C1(n16893), .C2(n16703), .A(n18138), .B(n16702), .ZN(
        n16704) );
  NOR3_X1 U19862 ( .A1(n16706), .A2(n16705), .A3(n16704), .ZN(n16707) );
  OAI221_X1 U19863 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n16708), .C1(n18699), 
        .C2(n16721), .A(n16707), .ZN(P3_U2656) );
  AOI211_X1 U19864 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16732), .A(n16709), .B(
        n16886), .ZN(n16716) );
  NOR2_X1 U19865 ( .A1(n17812), .A2(n17660), .ZN(n16741) );
  INV_X1 U19866 ( .A(n16741), .ZN(n17651) );
  NOR2_X1 U19867 ( .A1(n17662), .A2(n17651), .ZN(n16722) );
  OAI21_X1 U19868 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16722), .A(
        n16710), .ZN(n17641) );
  NOR2_X1 U19869 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17812), .ZN(
        n16875) );
  NAND2_X1 U19870 ( .A1(n17640), .A2(n16875), .ZN(n16727) );
  NAND2_X1 U19871 ( .A1(n16837), .A2(n16727), .ZN(n16712) );
  AOI21_X1 U19872 ( .B1(n17641), .B2(n16712), .A(n18657), .ZN(n16711) );
  OAI21_X1 U19873 ( .B1(n17641), .B2(n16712), .A(n16711), .ZN(n16713) );
  OAI211_X1 U19874 ( .C1(n16893), .C2(n16714), .A(n18138), .B(n16713), .ZN(
        n16715) );
  AOI211_X1 U19875 ( .C1(n16872), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16716), .B(n16715), .ZN(n16720) );
  NOR2_X1 U19876 ( .A1(n16887), .A2(n16717), .ZN(n16729) );
  NAND3_X1 U19877 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16729), .A3(n16718), 
        .ZN(n16719) );
  OAI211_X1 U19878 ( .C1(n16721), .C2(n18698), .A(n16720), .B(n16719), .ZN(
        P3_U2657) );
  AOI22_X1 U19879 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n16872), .B1(
        n16864), .B2(P3_EBX_REG_13__SCAN_IN), .ZN(n16737) );
  INV_X1 U19880 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16723) );
  NAND2_X1 U19881 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16741), .ZN(
        n16740) );
  AOI21_X1 U19882 ( .B1(n16723), .B2(n16740), .A(n16722), .ZN(n17654) );
  NAND2_X1 U19883 ( .A1(n16837), .A2(n16874), .ZN(n16883) );
  NOR2_X1 U19884 ( .A1(n17654), .A2(n16883), .ZN(n16728) );
  INV_X1 U19885 ( .A(n16740), .ZN(n16724) );
  OAI211_X1 U19886 ( .C1(n16853), .C2(n16724), .A(n16889), .B(n17654), .ZN(
        n16725) );
  INV_X1 U19887 ( .A(n16725), .ZN(n16726) );
  AOI211_X1 U19888 ( .C1(n16728), .C2(n16727), .A(n18126), .B(n16726), .ZN(
        n16736) );
  INV_X1 U19889 ( .A(n16729), .ZN(n16731) );
  OAI21_X1 U19890 ( .B1(n16745), .B2(n16887), .A(n16897), .ZN(n16755) );
  NOR2_X1 U19891 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16887), .ZN(n16744) );
  NOR2_X1 U19892 ( .A1(n16755), .A2(n16744), .ZN(n16730) );
  MUX2_X1 U19893 ( .A(n16731), .B(n16730), .S(P3_REIP_REG_13__SCAN_IN), .Z(
        n16735) );
  OAI211_X1 U19894 ( .C1(n16738), .C2(n16733), .A(n16895), .B(n16732), .ZN(
        n16734) );
  NAND4_X1 U19895 ( .A1(n16737), .A2(n16736), .A3(n16735), .A4(n16734), .ZN(
        P3_U2658) );
  AOI211_X1 U19896 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16756), .A(n16738), .B(
        n16886), .ZN(n16739) );
  AOI21_X1 U19897 ( .B1(n16872), .B2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16739), .ZN(n16748) );
  OAI21_X1 U19898 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n16741), .A(
        n16740), .ZN(n17666) );
  OAI21_X1 U19899 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17651), .A(
        n16837), .ZN(n16742) );
  XOR2_X1 U19900 ( .A(n17666), .B(n16742), .Z(n16743) );
  AOI22_X1 U19901 ( .A1(n16864), .A2(P3_EBX_REG_12__SCAN_IN), .B1(n16874), 
        .B2(n16743), .ZN(n16747) );
  AOI22_X1 U19902 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16755), .B1(n16745), 
        .B2(n16744), .ZN(n16746) );
  NAND4_X1 U19903 ( .A1(n16748), .A2(n16747), .A3(n16746), .A4(n18138), .ZN(
        P3_U2659) );
  OR2_X1 U19904 ( .A1(n16887), .A2(n16795), .ZN(n16786) );
  OAI21_X1 U19905 ( .B1(n16760), .B2(n16786), .A(n20924), .ZN(n16754) );
  AND2_X1 U19906 ( .A1(n17716), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17720) );
  NAND2_X1 U19907 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17720), .ZN(
        n16800) );
  INV_X1 U19908 ( .A(n16800), .ZN(n16789) );
  NAND2_X1 U19909 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16789), .ZN(
        n16788) );
  NOR2_X1 U19910 ( .A1(n16749), .A2(n16788), .ZN(n16762) );
  OAI21_X1 U19911 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16762), .A(
        n17651), .ZN(n17682) );
  INV_X1 U19912 ( .A(n16788), .ZN(n16778) );
  NAND2_X1 U19913 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16778), .ZN(
        n16777) );
  OAI21_X1 U19914 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16777), .A(
        n16837), .ZN(n16776) );
  OAI21_X1 U19915 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16853), .A(
        n16776), .ZN(n16765) );
  OAI21_X1 U19916 ( .B1(n17682), .B2(n16765), .A(n18138), .ZN(n16750) );
  AOI21_X1 U19917 ( .B1(n17682), .B2(n16765), .A(n16750), .ZN(n16752) );
  INV_X1 U19918 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16751) );
  OAI22_X1 U19919 ( .A1(n16850), .A2(n16752), .B1(n16751), .B2(n16882), .ZN(
        n16753) );
  AOI21_X1 U19920 ( .B1(n16755), .B2(n16754), .A(n16753), .ZN(n16758) );
  OAI211_X1 U19921 ( .C1(n16761), .C2(n16759), .A(n16895), .B(n16756), .ZN(
        n16757) );
  OAI211_X1 U19922 ( .C1(n16759), .C2(n16893), .A(n16758), .B(n16757), .ZN(
        P3_U2660) );
  OAI21_X1 U19923 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(P3_REIP_REG_9__SCAN_IN), 
        .A(n16760), .ZN(n16772) );
  AOI22_X1 U19924 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n16872), .B1(
        n16864), .B2(P3_EBX_REG_10__SCAN_IN), .ZN(n16771) );
  AOI21_X1 U19925 ( .B1(n16795), .B2(n16842), .A(n16881), .ZN(n16799) );
  INV_X1 U19926 ( .A(n16799), .ZN(n16769) );
  AOI211_X1 U19927 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16773), .A(n16761), .B(
        n16886), .ZN(n16768) );
  INV_X1 U19928 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16763) );
  AOI21_X1 U19929 ( .B1(n16763), .B2(n16777), .A(n16762), .ZN(n17696) );
  INV_X1 U19930 ( .A(n17696), .ZN(n16764) );
  OAI221_X1 U19931 ( .B1(n17696), .B2(n16765), .C1(n16764), .C2(n16776), .A(
        n16874), .ZN(n16766) );
  NAND2_X1 U19932 ( .A1(n18138), .A2(n16766), .ZN(n16767) );
  AOI211_X1 U19933 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(n16769), .A(n16768), 
        .B(n16767), .ZN(n16770) );
  OAI211_X1 U19934 ( .C1(n16786), .C2(n16772), .A(n16771), .B(n16770), .ZN(
        P3_U2661) );
  INV_X1 U19935 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18689) );
  OAI211_X1 U19936 ( .C1(n16787), .C2(n16775), .A(n16895), .B(n16773), .ZN(
        n16774) );
  OAI21_X1 U19937 ( .B1(n16775), .B2(n16893), .A(n16774), .ZN(n16784) );
  INV_X1 U19938 ( .A(n16776), .ZN(n16780) );
  OAI21_X1 U19939 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16778), .A(
        n16777), .ZN(n17706) );
  NOR3_X1 U19940 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A3(n16788), .ZN(n16779) );
  AOI211_X1 U19941 ( .C1(n16780), .C2(n17706), .A(n18126), .B(n16779), .ZN(
        n16782) );
  INV_X1 U19942 ( .A(n16866), .ZN(n16781) );
  OAI22_X1 U19943 ( .A1(n16850), .A2(n16782), .B1(n16781), .B2(n17706), .ZN(
        n16783) );
  AOI211_X1 U19944 ( .C1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n16872), .A(
        n16784), .B(n16783), .ZN(n16785) );
  OAI221_X1 U19945 ( .B1(P3_REIP_REG_9__SCAN_IN), .B2(n16786), .C1(n18689), 
        .C2(n16799), .A(n16785), .ZN(P3_U2662) );
  INV_X1 U19946 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n21043) );
  AOI211_X1 U19947 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16805), .A(n16787), .B(
        n16886), .ZN(n16794) );
  AOI21_X1 U19948 ( .B1(n17720), .B2(n16875), .A(n16853), .ZN(n16791) );
  OAI21_X1 U19949 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16789), .A(
        n16788), .ZN(n17730) );
  OAI21_X1 U19950 ( .B1(n16791), .B2(n17730), .A(n18138), .ZN(n16790) );
  AOI21_X1 U19951 ( .B1(n16791), .B2(n17730), .A(n16790), .ZN(n16792) );
  INV_X1 U19952 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n20937) );
  OAI22_X1 U19953 ( .A1(n16850), .A2(n16792), .B1(n20937), .B2(n16882), .ZN(
        n16793) );
  AOI211_X1 U19954 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16864), .A(n16794), .B(
        n16793), .ZN(n16798) );
  NAND3_X1 U19955 ( .A1(n16796), .A2(n16842), .A3(n16795), .ZN(n16797) );
  OAI211_X1 U19956 ( .C1(n16799), .C2(n21043), .A(n16798), .B(n16797), .ZN(
        P3_U2663) );
  AOI22_X1 U19957 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n16872), .B1(
        n16864), .B2(P3_EBX_REG_7__SCAN_IN), .ZN(n16810) );
  NOR2_X1 U19958 ( .A1(n17812), .A2(n17742), .ZN(n16822) );
  INV_X1 U19959 ( .A(n16822), .ZN(n16812) );
  NOR2_X1 U19960 ( .A1(n17757), .A2(n16812), .ZN(n16811) );
  INV_X1 U19961 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16884) );
  AOI21_X1 U19962 ( .B1(n16811), .B2(n16884), .A(n16853), .ZN(n16813) );
  OAI21_X1 U19963 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16811), .A(
        n16800), .ZN(n17741) );
  XNOR2_X1 U19964 ( .A(n16813), .B(n17741), .ZN(n16803) );
  NOR3_X1 U19965 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n16887), .A3(n16801), .ZN(
        n16802) );
  AOI211_X1 U19966 ( .C1(n16874), .C2(n16803), .A(n18126), .B(n16802), .ZN(
        n16809) );
  OAI21_X1 U19967 ( .B1(n16804), .B2(n16887), .A(n16897), .ZN(n16829) );
  INV_X1 U19968 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n20952) );
  AND3_X1 U19969 ( .A1(n20952), .A2(n16842), .A3(n16804), .ZN(n16819) );
  OAI21_X1 U19970 ( .B1(n16829), .B2(n16819), .A(P3_REIP_REG_7__SCAN_IN), .ZN(
        n16808) );
  OAI211_X1 U19971 ( .C1(n16817), .C2(n16806), .A(n16895), .B(n16805), .ZN(
        n16807) );
  NAND4_X1 U19972 ( .A1(n16810), .A2(n16809), .A3(n16808), .A4(n16807), .ZN(
        P3_U2664) );
  AOI21_X1 U19973 ( .B1(n17757), .B2(n16812), .A(n16811), .ZN(n17754) );
  NAND2_X1 U19974 ( .A1(n16874), .A2(n16813), .ZN(n16815) );
  OAI211_X1 U19975 ( .C1(n16822), .C2(n16853), .A(n17754), .B(n16889), .ZN(
        n16814) );
  OAI21_X1 U19976 ( .B1(n17754), .B2(n16815), .A(n16814), .ZN(n16816) );
  AOI211_X1 U19977 ( .C1(n16864), .C2(P3_EBX_REG_6__SCAN_IN), .A(n18126), .B(
        n16816), .ZN(n16821) );
  AOI211_X1 U19978 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16830), .A(n16817), .B(
        n16886), .ZN(n16818) );
  AOI211_X1 U19979 ( .C1(n16829), .C2(P3_REIP_REG_6__SCAN_IN), .A(n16819), .B(
        n16818), .ZN(n16820) );
  OAI211_X1 U19980 ( .C1(n17757), .C2(n16882), .A(n16821), .B(n16820), .ZN(
        P3_U2665) );
  INV_X1 U19981 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16826) );
  NAND2_X1 U19982 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17758), .ZN(
        n16835) );
  AOI21_X1 U19983 ( .B1(n16826), .B2(n16835), .A(n16822), .ZN(n17764) );
  AOI21_X1 U19984 ( .B1(n17758), .B2(n16875), .A(n16853), .ZN(n16839) );
  INV_X1 U19985 ( .A(n16839), .ZN(n16824) );
  INV_X1 U19986 ( .A(n17764), .ZN(n16823) );
  AOI221_X1 U19987 ( .B1(n17764), .B2(n16824), .C1(n16823), .C2(n16839), .A(
        n18126), .ZN(n16834) );
  OAI21_X1 U19988 ( .B1(n16887), .B2(n16825), .A(n18683), .ZN(n16828) );
  OAI22_X1 U19989 ( .A1(n16826), .A2(n16882), .B1(n16893), .B2(n16831), .ZN(
        n16827) );
  AOI21_X1 U19990 ( .B1(n16829), .B2(n16828), .A(n16827), .ZN(n16833) );
  OAI211_X1 U19991 ( .C1(n16840), .C2(n16831), .A(n16895), .B(n16830), .ZN(
        n16832) );
  OAI211_X1 U19992 ( .C1(n16850), .C2(n16834), .A(n16833), .B(n16832), .ZN(
        P3_U2666) );
  NOR2_X1 U19993 ( .A1(n17812), .A2(n17775), .ZN(n16851) );
  OAI21_X1 U19994 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16851), .A(
        n16835), .ZN(n17778) );
  INV_X1 U19995 ( .A(n16875), .ZN(n16836) );
  OR2_X1 U19996 ( .A1(n17775), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17782) );
  OAI22_X1 U19997 ( .A1(n16837), .A2(n17778), .B1(n16836), .B2(n17782), .ZN(
        n16838) );
  AOI211_X1 U19998 ( .C1(n16839), .C2(n17778), .A(n18126), .B(n16838), .ZN(
        n16849) );
  OAI21_X1 U19999 ( .B1(n16855), .B2(n16887), .A(n16897), .ZN(n16857) );
  AOI211_X1 U20000 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16858), .A(n16840), .B(
        n16886), .ZN(n16841) );
  AOI21_X1 U20001 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n16864), .A(n16841), .ZN(
        n16844) );
  INV_X1 U20002 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18681) );
  NAND3_X1 U20003 ( .A1(n16842), .A2(n16855), .A3(n18681), .ZN(n16843) );
  OAI211_X1 U20004 ( .C1(n16882), .C2(n17777), .A(n16844), .B(n16843), .ZN(
        n16845) );
  AOI21_X1 U20005 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n16857), .A(n16845), .ZN(
        n16848) );
  NOR2_X1 U20006 ( .A1(n17352), .A2(n16846), .ZN(n18814) );
  OAI21_X1 U20007 ( .B1(n17138), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n18814), .ZN(n16847) );
  OAI211_X1 U20008 ( .C1(n16850), .C2(n16849), .A(n16848), .B(n16847), .ZN(
        P3_U2667) );
  AOI22_X1 U20009 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n16872), .B1(
        n16864), .B2(P3_EBX_REG_3__SCAN_IN), .ZN(n16862) );
  INV_X1 U20010 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16852) );
  NAND2_X1 U20011 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16865) );
  AOI21_X1 U20012 ( .B1(n16852), .B2(n16865), .A(n16851), .ZN(n17789) );
  AOI21_X1 U20013 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n16875), .A(
        n16853), .ZN(n16873) );
  XOR2_X1 U20014 ( .A(n17789), .B(n16873), .Z(n16854) );
  NOR2_X1 U20015 ( .A1(n18762), .A2(n18769), .ZN(n18595) );
  NAND2_X1 U20016 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18595), .ZN(
        n18591) );
  INV_X1 U20017 ( .A(n18591), .ZN(n16863) );
  OAI21_X1 U20018 ( .B1(n16863), .B2(n18754), .A(n17142), .ZN(n18752) );
  AOI22_X1 U20019 ( .A1(n16874), .A2(n16854), .B1(n18814), .B2(n18752), .ZN(
        n16861) );
  NOR2_X1 U20020 ( .A1(n16855), .A2(n16887), .ZN(n16856) );
  AOI22_X1 U20021 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(n16857), .B1(n16868), 
        .B2(n16856), .ZN(n16860) );
  OAI211_X1 U20022 ( .C1(n16869), .C2(n17175), .A(n16895), .B(n16858), .ZN(
        n16859) );
  NAND4_X1 U20023 ( .A1(n16862), .A2(n16861), .A3(n16860), .A4(n16859), .ZN(
        P3_U2668) );
  AND2_X1 U20024 ( .A1(n18762), .A2(n18601), .ZN(n18596) );
  NOR2_X1 U20025 ( .A1(n16863), .A2(n18596), .ZN(n18759) );
  AOI22_X1 U20026 ( .A1(n16864), .A2(P3_EBX_REG_2__SCAN_IN), .B1(n18759), .B2(
        n18814), .ZN(n16879) );
  OAI21_X1 U20027 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16865), .ZN(n17799) );
  INV_X1 U20028 ( .A(n17799), .ZN(n16867) );
  AOI22_X1 U20029 ( .A1(n16881), .A2(P3_REIP_REG_2__SCAN_IN), .B1(n16867), 
        .B2(n16866), .ZN(n16878) );
  AOI211_X1 U20030 ( .C1(n21028), .C2(n18776), .A(n16868), .B(n16887), .ZN(
        n16871) );
  INV_X1 U20031 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17191) );
  INV_X1 U20032 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17186) );
  NAND2_X1 U20033 ( .A1(n17191), .A2(n17186), .ZN(n16885) );
  AOI211_X1 U20034 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16885), .A(n16869), .B(
        n16886), .ZN(n16870) );
  AOI211_X1 U20035 ( .C1(n16872), .C2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n16871), .B(n16870), .ZN(n16877) );
  OAI211_X1 U20036 ( .C1(n16875), .C2(n17799), .A(n16874), .B(n16873), .ZN(
        n16876) );
  NAND4_X1 U20037 ( .A1(n16879), .A2(n16878), .A3(n16877), .A4(n16876), .ZN(
        P3_U2669) );
  NAND2_X1 U20038 ( .A1(n18601), .A2(n16880), .ZN(n18619) );
  INV_X1 U20039 ( .A(n18619), .ZN(n18766) );
  AOI22_X1 U20040 ( .A1(n16881), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n18766), 
        .B2(n18814), .ZN(n16892) );
  OAI211_X1 U20041 ( .C1(n16884), .C2(n16883), .A(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B(n16882), .ZN(n16890) );
  OAI21_X1 U20042 ( .B1(n17186), .B2(n17191), .A(n16885), .ZN(n17187) );
  OAI22_X1 U20043 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16887), .B1(n16886), 
        .B2(n17187), .ZN(n16888) );
  AOI221_X1 U20044 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16890), .C1(
        n16889), .C2(n16890), .A(n16888), .ZN(n16891) );
  OAI211_X1 U20045 ( .C1(n16893), .C2(n17186), .A(n16892), .B(n16891), .ZN(
        P3_U2670) );
  AOI22_X1 U20046 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n16894), .B1(n18814), 
        .B2(n18774), .ZN(n16900) );
  OAI21_X1 U20047 ( .B1(n16896), .B2(n16895), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n16899) );
  INV_X1 U20048 ( .A(n18810), .ZN(n18749) );
  NAND3_X1 U20049 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18749), .A3(
        n16897), .ZN(n16898) );
  NAND3_X1 U20050 ( .A1(n16900), .A2(n16899), .A3(n16898), .ZN(P3_U2671) );
  INV_X1 U20051 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n16972) );
  NAND4_X1 U20052 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .A4(P3_EBX_REG_21__SCAN_IN), .ZN(n16902)
         );
  NAND4_X1 U20053 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_26__SCAN_IN), 
        .A3(P3_EBX_REG_25__SCAN_IN), .A4(n16931), .ZN(n16901) );
  NOR4_X1 U20054 ( .A1(n16972), .A2(n17011), .A3(n16902), .A4(n16901), .ZN(
        n16928) );
  NAND2_X1 U20055 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16928), .ZN(n16927) );
  NAND2_X1 U20056 ( .A1(n16927), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16904) );
  OR2_X1 U20057 ( .A1(n17160), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16903) );
  OAI22_X1 U20058 ( .A1(n17188), .A2(n16904), .B1(n16927), .B2(n16903), .ZN(
        P3_U2672) );
  AOI22_X1 U20059 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n9834), .ZN(n16908) );
  AOI22_X1 U20060 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n17123), .B1(
        n9832), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16907) );
  AOI22_X1 U20061 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n9831), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16906) );
  AOI22_X1 U20062 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17128), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16905) );
  NAND4_X1 U20063 ( .A1(n16908), .A2(n16907), .A3(n16906), .A4(n16905), .ZN(
        n16914) );
  AOI22_X1 U20064 ( .A1(n11630), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16912) );
  AOI22_X1 U20065 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n11696), .B1(
        P3_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n17108), .ZN(n16911) );
  AOI22_X1 U20066 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n17054), .B1(
        P3_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n17094), .ZN(n16910) );
  AOI22_X1 U20067 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n17145), .B1(
        P3_INSTQUEUE_REG_5__7__SCAN_IN), .B2(n17146), .ZN(n16909) );
  NAND4_X1 U20068 ( .A1(n16912), .A2(n16911), .A3(n16910), .A4(n16909), .ZN(
        n16913) );
  NOR2_X1 U20069 ( .A1(n16914), .A2(n16913), .ZN(n16926) );
  AOI22_X1 U20070 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16918) );
  AOI22_X1 U20071 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9831), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16917) );
  AOI22_X1 U20072 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17128), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16916) );
  AOI22_X1 U20073 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17107), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16915) );
  NAND4_X1 U20074 ( .A1(n16918), .A2(n16917), .A3(n16916), .A4(n16915), .ZN(
        n16924) );
  AOI22_X1 U20075 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16922) );
  AOI22_X1 U20076 ( .A1(n11696), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11519), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16921) );
  AOI22_X1 U20077 ( .A1(n9834), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16920) );
  AOI22_X1 U20078 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16919) );
  NAND4_X1 U20079 ( .A1(n16922), .A2(n16921), .A3(n16920), .A4(n16919), .ZN(
        n16923) );
  NOR2_X1 U20080 ( .A1(n16924), .A2(n16923), .ZN(n16934) );
  INV_X1 U20081 ( .A(n16939), .ZN(n16933) );
  NOR3_X1 U20082 ( .A1(n16934), .A2(n16933), .A3(n16932), .ZN(n16925) );
  XOR2_X1 U20083 ( .A(n16926), .B(n16925), .Z(n17203) );
  OAI211_X1 U20084 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16928), .A(n16927), .B(
        n17178), .ZN(n16929) );
  OAI21_X1 U20085 ( .B1(n17203), .B2(n17178), .A(n16929), .ZN(P3_U2673) );
  NAND2_X1 U20086 ( .A1(n16931), .A2(n16930), .ZN(n16938) );
  NOR2_X1 U20087 ( .A1(n16933), .A2(n16932), .ZN(n16935) );
  XNOR2_X1 U20088 ( .A(n16935), .B(n16934), .ZN(n17207) );
  AOI22_X1 U20089 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16936), .B1(n17188), 
        .B2(n17207), .ZN(n16937) );
  OAI21_X1 U20090 ( .B1(n16944), .B2(n16938), .A(n16937), .ZN(P3_U2674) );
  AOI21_X1 U20091 ( .B1(n16940), .B2(n16945), .A(n16939), .ZN(n17217) );
  NAND2_X1 U20092 ( .A1(n17188), .A2(n17217), .ZN(n16941) );
  OAI221_X1 U20093 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n16944), .C1(n16943), 
        .C2(n16942), .A(n16941), .ZN(P3_U2676) );
  AOI21_X1 U20094 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17184), .A(n16952), .ZN(
        n16948) );
  OAI21_X1 U20095 ( .B1(n16947), .B2(n16946), .A(n16945), .ZN(n17225) );
  OAI22_X1 U20096 ( .A1(n16949), .A2(n16948), .B1(n17184), .B2(n17225), .ZN(
        P3_U2677) );
  AOI21_X1 U20097 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17184), .A(n9876), .ZN(
        n16951) );
  XNOR2_X1 U20098 ( .A(n16950), .B(n16953), .ZN(n17230) );
  OAI22_X1 U20099 ( .A1(n16952), .A2(n16951), .B1(n17184), .B2(n17230), .ZN(
        P3_U2678) );
  AOI21_X1 U20100 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17184), .A(n9877), .ZN(
        n16956) );
  OAI21_X1 U20101 ( .B1(n16955), .B2(n16954), .A(n16953), .ZN(n17236) );
  OAI22_X1 U20102 ( .A1(n9876), .A2(n16956), .B1(n17184), .B2(n17236), .ZN(
        P3_U2679) );
  AOI21_X1 U20103 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17184), .A(n9853), .ZN(
        n16959) );
  XNOR2_X1 U20104 ( .A(n16958), .B(n16957), .ZN(n17239) );
  OAI22_X1 U20105 ( .A1(n9877), .A2(n16959), .B1(n17184), .B2(n17239), .ZN(
        P3_U2680) );
  AOI21_X1 U20106 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17184), .A(n16960), .ZN(
        n16971) );
  AOI22_X1 U20107 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17107), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16964) );
  AOI22_X1 U20108 ( .A1(n11696), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16963) );
  AOI22_X1 U20109 ( .A1(n17128), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9831), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16962) );
  AOI22_X1 U20110 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9832), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16961) );
  NAND4_X1 U20111 ( .A1(n16964), .A2(n16963), .A3(n16962), .A4(n16961), .ZN(
        n16970) );
  AOI22_X1 U20112 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16968) );
  AOI22_X1 U20113 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9834), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16967) );
  AOI22_X1 U20114 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11519), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16966) );
  AOI22_X1 U20115 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16965) );
  NAND4_X1 U20116 ( .A1(n16968), .A2(n16967), .A3(n16966), .A4(n16965), .ZN(
        n16969) );
  NOR2_X1 U20117 ( .A1(n16970), .A2(n16969), .ZN(n17243) );
  OAI22_X1 U20118 ( .A1(n9853), .A2(n16971), .B1(n17243), .B2(n17178), .ZN(
        P3_U2681) );
  OAI21_X1 U20119 ( .B1(n16972), .B2(n17011), .A(n17178), .ZN(n16998) );
  AOI22_X1 U20120 ( .A1(n9831), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9832), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16983) );
  AOI22_X1 U20121 ( .A1(n17128), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17094), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16982) );
  INV_X1 U20122 ( .A(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n21185) );
  AOI22_X1 U20123 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17107), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n16973) );
  OAI21_X1 U20124 ( .B1(n16974), .B2(n21185), .A(n16973), .ZN(n16980) );
  AOI22_X1 U20125 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16978) );
  AOI22_X1 U20126 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9834), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16977) );
  AOI22_X1 U20127 ( .A1(n11696), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11519), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16976) );
  AOI22_X1 U20128 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16975) );
  NAND4_X1 U20129 ( .A1(n16978), .A2(n16977), .A3(n16976), .A4(n16975), .ZN(
        n16979) );
  AOI211_X1 U20130 ( .C1(n17153), .C2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A(
        n16980), .B(n16979), .ZN(n16981) );
  NAND3_X1 U20131 ( .A1(n16983), .A2(n16982), .A3(n16981), .ZN(n17248) );
  NAND2_X1 U20132 ( .A1(n17188), .A2(n17248), .ZN(n16984) );
  OAI221_X1 U20133 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n16986), .C1(n16985), 
        .C2(n16998), .A(n16984), .ZN(P3_U2682) );
  AOI22_X1 U20134 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16990) );
  AOI22_X1 U20135 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11519), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16989) );
  AOI22_X1 U20136 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17107), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16988) );
  AOI22_X1 U20137 ( .A1(n11534), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11696), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n16987) );
  NAND4_X1 U20138 ( .A1(n16990), .A2(n16989), .A3(n16988), .A4(n16987), .ZN(
        n16996) );
  AOI22_X1 U20139 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16994) );
  AOI22_X1 U20140 ( .A1(n17128), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9831), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16993) );
  AOI22_X1 U20141 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9834), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16992) );
  AOI22_X1 U20142 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16991) );
  NAND4_X1 U20143 ( .A1(n16994), .A2(n16993), .A3(n16992), .A4(n16991), .ZN(
        n16995) );
  NOR2_X1 U20144 ( .A1(n16996), .A2(n16995), .ZN(n17257) );
  NOR2_X1 U20145 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16997), .ZN(n16999) );
  OAI22_X1 U20146 ( .A1(n17257), .A2(n17178), .B1(n16999), .B2(n16998), .ZN(
        P3_U2683) );
  AOI22_X1 U20147 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9832), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17003) );
  AOI22_X1 U20148 ( .A1(n11696), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11519), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17002) );
  AOI22_X1 U20149 ( .A1(n11534), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9834), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17001) );
  AOI22_X1 U20150 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17000) );
  NAND4_X1 U20151 ( .A1(n17003), .A2(n17002), .A3(n17001), .A4(n17000), .ZN(
        n17010) );
  AOI22_X1 U20152 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17008) );
  AOI22_X1 U20153 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9831), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17007) );
  AOI22_X1 U20154 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17107), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17006) );
  AOI22_X1 U20155 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17005) );
  NAND4_X1 U20156 ( .A1(n17008), .A2(n17007), .A3(n17006), .A4(n17005), .ZN(
        n17009) );
  NOR2_X1 U20157 ( .A1(n17010), .A2(n17009), .ZN(n17261) );
  OAI21_X1 U20158 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17023), .A(n17011), .ZN(
        n17012) );
  AOI22_X1 U20159 ( .A1(n17188), .A2(n17261), .B1(n17012), .B2(n17178), .ZN(
        P3_U2684) );
  NOR3_X1 U20160 ( .A1(n17160), .A2(n17053), .A3(n17050), .ZN(n17038) );
  NAND2_X1 U20161 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17038), .ZN(n17037) );
  AOI22_X1 U20162 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11534), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17022) );
  AOI22_X1 U20163 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17107), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17021) );
  AOI22_X1 U20164 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17020) );
  AND2_X1 U20165 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n17018) );
  AOI22_X1 U20166 ( .A1(n17128), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9831), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17016) );
  AOI22_X1 U20167 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17015) );
  AOI22_X1 U20168 ( .A1(n9834), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17094), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17014) );
  AOI22_X1 U20169 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11696), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17013) );
  NAND4_X1 U20170 ( .A1(n17016), .A2(n17015), .A3(n17014), .A4(n17013), .ZN(
        n17017) );
  AOI211_X1 U20171 ( .C1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .C2(n9830), .A(
        n17018), .B(n17017), .ZN(n17019) );
  NAND4_X1 U20172 ( .A1(n17022), .A2(n17021), .A3(n17020), .A4(n17019), .ZN(
        n17262) );
  OAI21_X1 U20173 ( .B1(n17024), .B2(n17023), .A(n17178), .ZN(n17025) );
  OAI21_X1 U20174 ( .B1(n17184), .B2(n17262), .A(n17025), .ZN(n17026) );
  OAI21_X1 U20175 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17037), .A(n17026), .ZN(
        P3_U2685) );
  AOI22_X1 U20176 ( .A1(n11534), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17030) );
  AOI22_X1 U20177 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17128), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17029) );
  AOI22_X1 U20178 ( .A1(n11696), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17028) );
  AOI22_X1 U20179 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9832), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17027) );
  NAND4_X1 U20180 ( .A1(n17030), .A2(n17029), .A3(n17028), .A4(n17027), .ZN(
        n17036) );
  AOI22_X1 U20181 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17034) );
  AOI22_X1 U20182 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17033) );
  AOI22_X1 U20183 ( .A1(n9831), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9834), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17032) );
  AOI22_X1 U20184 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17031) );
  NAND4_X1 U20185 ( .A1(n17034), .A2(n17033), .A3(n17032), .A4(n17031), .ZN(
        n17035) );
  NOR2_X1 U20186 ( .A1(n17036), .A2(n17035), .ZN(n17274) );
  OAI211_X1 U20187 ( .C1(n17038), .C2(P3_EBX_REG_17__SCAN_IN), .A(n17178), .B(
        n17037), .ZN(n17039) );
  OAI21_X1 U20188 ( .B1(n17274), .B2(n17178), .A(n17039), .ZN(P3_U2686) );
  NAND2_X1 U20189 ( .A1(n17184), .A2(n17050), .ZN(n17066) );
  AOI22_X1 U20190 ( .A1(n9831), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17049) );
  AOI22_X1 U20191 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9832), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17048) );
  AOI22_X1 U20192 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17047) );
  AND2_X1 U20193 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n17045) );
  AOI22_X1 U20194 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17043) );
  AOI22_X1 U20195 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17094), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17042) );
  AOI22_X1 U20196 ( .A1(n17128), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11696), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17041) );
  AOI22_X1 U20197 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9834), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17040) );
  NAND4_X1 U20198 ( .A1(n17043), .A2(n17042), .A3(n17041), .A4(n17040), .ZN(
        n17044) );
  AOI211_X1 U20199 ( .C1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .C2(n9830), .A(
        n17045), .B(n17044), .ZN(n17046) );
  NAND4_X1 U20200 ( .A1(n17049), .A2(n17048), .A3(n17047), .A4(n17046), .ZN(
        n17275) );
  NOR2_X1 U20201 ( .A1(n17160), .A2(n17050), .ZN(n17051) );
  AOI22_X1 U20202 ( .A1(n17188), .A2(n17275), .B1(n17051), .B2(n17053), .ZN(
        n17052) );
  OAI21_X1 U20203 ( .B1(n17053), .B2(n17066), .A(n17052), .ZN(P3_U2687) );
  AOI22_X1 U20204 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n9834), .B1(
        n17153), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17058) );
  AOI22_X1 U20205 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n9832), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17057) );
  AOI22_X1 U20206 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__7__SCAN_IN), .B2(n17094), .ZN(n17056) );
  AOI22_X1 U20207 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n17054), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17055) );
  NAND4_X1 U20208 ( .A1(n17058), .A2(n17057), .A3(n17056), .A4(n17055), .ZN(
        n17064) );
  AOI22_X1 U20209 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17062) );
  AOI22_X1 U20210 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n17144), .B1(
        n9831), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17061) );
  AOI22_X1 U20211 ( .A1(n11696), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n17108), .ZN(n17060) );
  AOI22_X1 U20212 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n17145), .B1(
        P3_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n17146), .ZN(n17059) );
  NAND4_X1 U20213 ( .A1(n17062), .A2(n17061), .A3(n17060), .A4(n17059), .ZN(
        n17063) );
  NOR2_X1 U20214 ( .A1(n17064), .A2(n17063), .ZN(n17285) );
  NOR2_X1 U20215 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17065), .ZN(n17067) );
  OAI22_X1 U20216 ( .A1(n17285), .A2(n17178), .B1(n17067), .B2(n17066), .ZN(
        P3_U2688) );
  NAND2_X1 U20217 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17068), .ZN(n17080) );
  AOI22_X1 U20218 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17072) );
  AOI22_X1 U20219 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11696), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17071) );
  AOI22_X1 U20220 ( .A1(n9834), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17070) );
  AOI22_X1 U20221 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9831), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17069) );
  NAND4_X1 U20222 ( .A1(n17072), .A2(n17071), .A3(n17070), .A4(n17069), .ZN(
        n17078) );
  AOI22_X1 U20223 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17076) );
  AOI22_X1 U20224 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17153), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17075) );
  AOI22_X1 U20225 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17074) );
  AOI22_X1 U20226 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17073) );
  NAND4_X1 U20227 ( .A1(n17076), .A2(n17075), .A3(n17074), .A4(n17073), .ZN(
        n17077) );
  NOR2_X1 U20228 ( .A1(n17078), .A2(n17077), .ZN(n17291) );
  NAND3_X1 U20229 ( .A1(n17080), .A2(P3_EBX_REG_14__SCAN_IN), .A3(n17184), 
        .ZN(n17079) );
  OAI221_X1 U20230 ( .B1(n17080), .B2(P3_EBX_REG_14__SCAN_IN), .C1(n17184), 
        .C2(n17291), .A(n17079), .ZN(P3_U2689) );
  AOI22_X1 U20231 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11696), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17084) );
  AOI22_X1 U20232 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17083) );
  AOI22_X1 U20233 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17082) );
  AOI22_X1 U20234 ( .A1(n9831), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17081) );
  NAND4_X1 U20235 ( .A1(n17084), .A2(n17083), .A3(n17082), .A4(n17081), .ZN(
        n17090) );
  AOI22_X1 U20236 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17088) );
  AOI22_X1 U20237 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17153), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17087) );
  AOI22_X1 U20238 ( .A1(n11534), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9834), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17086) );
  AOI22_X1 U20239 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17085) );
  NAND4_X1 U20240 ( .A1(n17088), .A2(n17087), .A3(n17086), .A4(n17085), .ZN(
        n17089) );
  NOR2_X1 U20241 ( .A1(n17090), .A2(n17089), .ZN(n17297) );
  OAI21_X1 U20242 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17106), .A(n17091), .ZN(
        n17092) );
  OAI21_X1 U20243 ( .B1(n17297), .B2(n17178), .A(n17092), .ZN(P3_U2691) );
  INV_X1 U20244 ( .A(n17119), .ZN(n17093) );
  OAI21_X1 U20245 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17093), .A(n17178), .ZN(
        n17105) );
  AOI22_X1 U20246 ( .A1(n11534), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17098) );
  AOI22_X1 U20247 ( .A1(n9831), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17094), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17097) );
  AOI22_X1 U20248 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9832), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17096) );
  AOI22_X1 U20249 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11696), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17095) );
  NAND4_X1 U20250 ( .A1(n17098), .A2(n17097), .A3(n17096), .A4(n17095), .ZN(
        n17104) );
  AOI22_X1 U20251 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17102) );
  AOI22_X1 U20252 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9834), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17101) );
  AOI22_X1 U20253 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17100) );
  AOI22_X1 U20254 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17099) );
  NAND4_X1 U20255 ( .A1(n17102), .A2(n17101), .A3(n17100), .A4(n17099), .ZN(
        n17103) );
  NOR2_X1 U20256 ( .A1(n17104), .A2(n17103), .ZN(n17302) );
  OAI22_X1 U20257 ( .A1(n17106), .A2(n17105), .B1(n17302), .B2(n17178), .ZN(
        P3_U2692) );
  AOI22_X1 U20258 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17112) );
  AOI22_X1 U20259 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17107), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17111) );
  AOI22_X1 U20260 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9834), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17110) );
  AOI22_X1 U20261 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17109) );
  NAND4_X1 U20262 ( .A1(n17112), .A2(n17111), .A3(n17110), .A4(n17109), .ZN(
        n17118) );
  AOI22_X1 U20263 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17116) );
  AOI22_X1 U20264 ( .A1(n9831), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11534), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17115) );
  AOI22_X1 U20265 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11696), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17114) );
  AOI22_X1 U20266 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17113) );
  NAND4_X1 U20267 ( .A1(n17116), .A2(n17115), .A3(n17114), .A4(n17113), .ZN(
        n17117) );
  NOR2_X1 U20268 ( .A1(n17118), .A2(n17117), .ZN(n17309) );
  OAI21_X1 U20269 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17136), .A(n17119), .ZN(
        n17120) );
  AOI22_X1 U20270 ( .A1(n17188), .A2(n17309), .B1(n17120), .B2(n17178), .ZN(
        P3_U2693) );
  INV_X1 U20271 ( .A(n17157), .ZN(n17121) );
  OAI21_X1 U20272 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17121), .A(n17178), .ZN(
        n17135) );
  AOI22_X1 U20273 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17127) );
  AOI22_X1 U20274 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11534), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17126) );
  AOI22_X1 U20275 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11519), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17125) );
  AOI22_X1 U20276 ( .A1(n9831), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9832), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17124) );
  NAND4_X1 U20277 ( .A1(n17127), .A2(n17126), .A3(n17125), .A4(n17124), .ZN(
        n17134) );
  AOI22_X1 U20278 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17132) );
  AOI22_X1 U20279 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17128), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17131) );
  AOI22_X1 U20280 ( .A1(n11696), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9834), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17130) );
  AOI22_X1 U20281 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17129) );
  NAND4_X1 U20282 ( .A1(n17132), .A2(n17131), .A3(n17130), .A4(n17129), .ZN(
        n17133) );
  NOR2_X1 U20283 ( .A1(n17134), .A2(n17133), .ZN(n17311) );
  OAI22_X1 U20284 ( .A1(n17136), .A2(n17135), .B1(n17311), .B2(n17178), .ZN(
        P3_U2694) );
  AOI22_X1 U20285 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17137), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17156) );
  AOI22_X1 U20286 ( .A1(n17140), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11696), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17155) );
  AOI22_X1 U20287 ( .A1(n9831), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9832), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17141) );
  OAI21_X1 U20288 ( .B1(n17142), .B2(n21041), .A(n17141), .ZN(n17152) );
  AOI22_X1 U20289 ( .A1(n11630), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17150) );
  AOI22_X1 U20290 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17122), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17149) );
  AOI22_X1 U20291 ( .A1(n9834), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11519), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17148) );
  AOI22_X1 U20292 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17145), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17147) );
  NAND4_X1 U20293 ( .A1(n17150), .A2(n17149), .A3(n17148), .A4(n17147), .ZN(
        n17151) );
  AOI211_X1 U20294 ( .C1(n17153), .C2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A(
        n17152), .B(n17151), .ZN(n17154) );
  NAND3_X1 U20295 ( .A1(n17156), .A2(n17155), .A3(n17154), .ZN(n17316) );
  INV_X1 U20296 ( .A(n17316), .ZN(n17159) );
  OAI21_X1 U20297 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17163), .A(n17157), .ZN(
        n17158) );
  AOI22_X1 U20298 ( .A1(n17188), .A2(n17159), .B1(n17158), .B2(n17178), .ZN(
        P3_U2695) );
  NOR2_X1 U20299 ( .A1(n17160), .A2(n17164), .ZN(n17165) );
  AOI22_X1 U20300 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n17178), .B1(
        P3_EBX_REG_6__SCAN_IN), .B2(n17165), .ZN(n17162) );
  INV_X1 U20301 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17161) );
  OAI22_X1 U20302 ( .A1(n17163), .A2(n17162), .B1(n17161), .B2(n17178), .ZN(
        P3_U2696) );
  NAND2_X1 U20303 ( .A1(n17184), .A2(n17164), .ZN(n17169) );
  AOI22_X1 U20304 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n17188), .B1(
        n17165), .B2(n17167), .ZN(n17166) );
  OAI21_X1 U20305 ( .B1(n17167), .B2(n17169), .A(n17166), .ZN(P3_U2697) );
  NOR2_X1 U20306 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17174), .ZN(n17170) );
  INV_X1 U20307 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17168) );
  OAI22_X1 U20308 ( .A1(n17170), .A2(n17169), .B1(n17168), .B2(n17178), .ZN(
        P3_U2698) );
  OAI21_X1 U20309 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17171), .A(n17178), .ZN(
        n17173) );
  INV_X1 U20310 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17172) );
  OAI22_X1 U20311 ( .A1(n17174), .A2(n17173), .B1(n17172), .B2(n17178), .ZN(
        P3_U2699) );
  NOR2_X1 U20312 ( .A1(n17188), .A2(n17176), .ZN(n17180) );
  OAI222_X1 U20313 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n18188), .B1(
        P3_EBX_REG_3__SCAN_IN), .B2(n17176), .C1(n17180), .C2(n17175), .ZN(
        n17177) );
  OAI21_X1 U20314 ( .B1(n17179), .B2(n17178), .A(n17177), .ZN(P3_U2700) );
  OAI21_X1 U20315 ( .B1(P3_EBX_REG_2__SCAN_IN), .B2(n17181), .A(n17180), .ZN(
        n17182) );
  OAI21_X1 U20316 ( .B1(n17184), .B2(n17183), .A(n17182), .ZN(P3_U2701) );
  INV_X1 U20317 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17185) );
  OAI222_X1 U20318 ( .A1(n17187), .A2(n17192), .B1(n17186), .B2(n17190), .C1(
        n17185), .C2(n17184), .ZN(P3_U2702) );
  NAND2_X1 U20319 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17188), .ZN(
        n17189) );
  OAI221_X1 U20320 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17192), .C1(n17191), 
        .C2(n17190), .A(n17189), .ZN(P3_U2703) );
  NAND2_X1 U20321 ( .A1(n17319), .A2(n17193), .ZN(n17281) );
  INV_X1 U20322 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17416) );
  INV_X1 U20323 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17412) );
  INV_X1 U20324 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17410) );
  INV_X1 U20325 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n21079) );
  INV_X1 U20326 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17395) );
  NAND2_X1 U20327 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .ZN(n17346) );
  INV_X1 U20328 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17434) );
  INV_X1 U20329 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17432) );
  NAND4_X1 U20330 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n17194) );
  NOR4_X1 U20331 ( .A1(n17346), .A2(n17434), .A3(n17432), .A4(n17194), .ZN(
        n17286) );
  NAND2_X1 U20332 ( .A1(n17286), .A2(n17195), .ZN(n17315) );
  INV_X1 U20333 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17444) );
  NAND2_X1 U20334 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .ZN(n17287) );
  NAND4_X1 U20335 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(P3_EAX_REG_13__SCAN_IN), 
        .A3(P3_EAX_REG_12__SCAN_IN), .A4(P3_EAX_REG_11__SCAN_IN), .ZN(n17196)
         );
  NAND2_X1 U20336 ( .A1(P3_EAX_REG_15__SCAN_IN), .A2(n17288), .ZN(n17282) );
  NOR2_X2 U20337 ( .A1(n17395), .A2(n17282), .ZN(n17277) );
  INV_X1 U20338 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17403) );
  INV_X1 U20339 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17401) );
  INV_X1 U20340 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17399) );
  INV_X1 U20341 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17397) );
  NOR4_X1 U20342 ( .A1(n17403), .A2(n17401), .A3(n17399), .A4(n17397), .ZN(
        n17197) );
  NAND4_X1 U20343 ( .A1(n17277), .A2(P3_EAX_REG_22__SCAN_IN), .A3(
        P3_EAX_REG_21__SCAN_IN), .A4(n17197), .ZN(n17238) );
  NAND2_X1 U20344 ( .A1(n18188), .A2(n17237), .ZN(n17231) );
  OR2_X2 U20345 ( .A1(n17410), .A2(n17231), .ZN(n17232) );
  NOR2_X2 U20346 ( .A1(n17412), .A2(n17232), .ZN(n17226) );
  NAND2_X1 U20347 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17218), .ZN(n17214) );
  NAND2_X1 U20348 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17209), .ZN(n17208) );
  NOR2_X1 U20349 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(n17208), .ZN(n17199) );
  NAND2_X1 U20350 ( .A1(n17339), .A2(n17208), .ZN(n17206) );
  OAI21_X1 U20351 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17337), .A(n17206), .ZN(
        n17198) );
  AOI22_X1 U20352 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17199), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17198), .ZN(n17200) );
  OAI21_X1 U20353 ( .B1(n20974), .B2(n17281), .A(n17200), .ZN(P3_U2704) );
  INV_X1 U20354 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17422) );
  NOR2_X2 U20355 ( .A1(n17201), .A2(n17339), .ZN(n17276) );
  OAI22_X1 U20356 ( .A1(n17203), .A2(n17350), .B1(n17202), .B2(n17281), .ZN(
        n17204) );
  AOI21_X1 U20357 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n17276), .A(n17204), .ZN(
        n17205) );
  OAI221_X1 U20358 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17208), .C1(n17422), 
        .C2(n17206), .A(n17205), .ZN(P3_U2705) );
  AOI22_X1 U20359 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17276), .B1(n17207), .B2(
        n17317), .ZN(n17211) );
  OAI211_X1 U20360 ( .C1(n17209), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17339), .B(
        n17208), .ZN(n17210) );
  OAI211_X1 U20361 ( .C1(n17281), .C2(n17212), .A(n17211), .B(n17210), .ZN(
        P3_U2706) );
  AOI22_X1 U20362 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17276), .B1(n17213), .B2(
        n17317), .ZN(n17216) );
  OAI211_X1 U20363 ( .C1(n17218), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17339), .B(
        n17214), .ZN(n17215) );
  OAI211_X1 U20364 ( .C1(n17281), .C2(n21025), .A(n17216), .B(n17215), .ZN(
        P3_U2707) );
  AOI22_X1 U20365 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17276), .B1(n17217), .B2(
        n17317), .ZN(n17221) );
  AOI211_X1 U20366 ( .C1(n17416), .C2(n17222), .A(n17218), .B(n17319), .ZN(
        n17219) );
  INV_X1 U20367 ( .A(n17219), .ZN(n17220) );
  OAI211_X1 U20368 ( .C1(n17281), .C2(n19178), .A(n17221), .B(n17220), .ZN(
        P3_U2708) );
  AOI22_X1 U20369 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17276), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17268), .ZN(n17224) );
  OAI211_X1 U20370 ( .C1(n17226), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17339), .B(
        n17222), .ZN(n17223) );
  OAI211_X1 U20371 ( .C1(n17350), .C2(n17225), .A(n17224), .B(n17223), .ZN(
        P3_U2709) );
  AOI22_X1 U20372 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17276), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17268), .ZN(n17229) );
  AOI211_X1 U20373 ( .C1(n17412), .C2(n17232), .A(n17226), .B(n17319), .ZN(
        n17227) );
  INV_X1 U20374 ( .A(n17227), .ZN(n17228) );
  OAI211_X1 U20375 ( .C1(n17350), .C2(n17230), .A(n17229), .B(n17228), .ZN(
        P3_U2710) );
  AOI22_X1 U20376 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17276), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17268), .ZN(n17235) );
  OAI21_X1 U20377 ( .B1(n17410), .B2(n17319), .A(n17231), .ZN(n17233) );
  NAND2_X1 U20378 ( .A1(n17233), .A2(n17232), .ZN(n17234) );
  OAI211_X1 U20379 ( .C1(n17350), .C2(n17236), .A(n17235), .B(n17234), .ZN(
        P3_U2711) );
  AOI211_X1 U20380 ( .C1(n21079), .C2(n17238), .A(n17319), .B(n17237), .ZN(
        n17241) );
  INV_X1 U20381 ( .A(n17276), .ZN(n17267) );
  OAI22_X1 U20382 ( .A1(n18185), .A2(n17267), .B1(n17350), .B2(n17239), .ZN(
        n17240) );
  AOI211_X1 U20383 ( .C1(n17268), .C2(BUF2_REG_23__SCAN_IN), .A(n17241), .B(
        n17240), .ZN(n17242) );
  INV_X1 U20384 ( .A(n17242), .ZN(P3_U2712) );
  NAND2_X1 U20385 ( .A1(n18188), .A2(n17277), .ZN(n17269) );
  NAND2_X1 U20386 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17263), .ZN(n17258) );
  NOR2_X1 U20387 ( .A1(n17403), .A2(n17258), .ZN(n17249) );
  INV_X1 U20388 ( .A(n17249), .ZN(n17253) );
  NAND2_X1 U20389 ( .A1(n17339), .A2(n17253), .ZN(n17252) );
  OAI21_X1 U20390 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17337), .A(n17252), .ZN(
        n17246) );
  INV_X1 U20391 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17405) );
  NOR3_X1 U20392 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17405), .A3(n17253), .ZN(
        n17245) );
  OAI22_X1 U20393 ( .A1(n17243), .A2(n17350), .B1(n15303), .B2(n17281), .ZN(
        n17244) );
  AOI211_X1 U20394 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n17246), .A(n17245), .B(
        n17244), .ZN(n17247) );
  OAI21_X1 U20395 ( .B1(n18181), .B2(n17267), .A(n17247), .ZN(P3_U2713) );
  AOI22_X1 U20396 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n17268), .B1(n17317), .B2(
        n17248), .ZN(n17251) );
  AOI22_X1 U20397 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17276), .B1(n17249), .B2(
        n17405), .ZN(n17250) );
  OAI211_X1 U20398 ( .C1(n17405), .C2(n17252), .A(n17251), .B(n17250), .ZN(
        P3_U2714) );
  AOI22_X1 U20399 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17276), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17268), .ZN(n17256) );
  INV_X1 U20400 ( .A(n17258), .ZN(n17254) );
  OAI211_X1 U20401 ( .C1(n17254), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17339), .B(
        n17253), .ZN(n17255) );
  OAI211_X1 U20402 ( .C1(n17257), .C2(n17350), .A(n17256), .B(n17255), .ZN(
        P3_U2715) );
  AOI22_X1 U20403 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17276), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17268), .ZN(n17260) );
  OAI211_X1 U20404 ( .C1(n17263), .C2(P3_EAX_REG_19__SCAN_IN), .A(n17339), .B(
        n17258), .ZN(n17259) );
  OAI211_X1 U20405 ( .C1(n17261), .C2(n17350), .A(n17260), .B(n17259), .ZN(
        P3_U2716) );
  AOI22_X1 U20406 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n17268), .B1(n17317), .B2(
        n17262), .ZN(n17266) );
  AOI211_X1 U20407 ( .C1(n17399), .C2(n17270), .A(n17263), .B(n17319), .ZN(
        n17264) );
  INV_X1 U20408 ( .A(n17264), .ZN(n17265) );
  OAI211_X1 U20409 ( .C1(n17267), .C2(n18166), .A(n17266), .B(n17265), .ZN(
        P3_U2717) );
  AOI22_X1 U20410 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17276), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17268), .ZN(n17273) );
  OAI21_X1 U20411 ( .B1(n17397), .B2(n17319), .A(n17269), .ZN(n17271) );
  NAND2_X1 U20412 ( .A1(n17271), .A2(n17270), .ZN(n17272) );
  OAI211_X1 U20413 ( .C1(n17274), .C2(n17350), .A(n17273), .B(n17272), .ZN(
        P3_U2718) );
  AOI22_X1 U20414 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17276), .B1(n17317), .B2(
        n17275), .ZN(n17280) );
  AOI211_X1 U20415 ( .C1(n17395), .C2(n17282), .A(n17319), .B(n17277), .ZN(
        n17278) );
  INV_X1 U20416 ( .A(n17278), .ZN(n17279) );
  OAI211_X1 U20417 ( .C1(n17281), .C2(n14135), .A(n17280), .B(n17279), .ZN(
        P3_U2719) );
  OAI211_X1 U20418 ( .C1(P3_EAX_REG_15__SCAN_IN), .C2(n17288), .A(n17339), .B(
        n17282), .ZN(n17284) );
  NAND2_X1 U20419 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17345), .ZN(n17283) );
  OAI211_X1 U20420 ( .C1(n17285), .C2(n17350), .A(n17284), .B(n17283), .ZN(
        P3_U2720) );
  INV_X1 U20421 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17451) );
  INV_X1 U20422 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17446) );
  INV_X1 U20423 ( .A(n17337), .ZN(n17347) );
  NAND2_X1 U20424 ( .A1(n17286), .A2(n17347), .ZN(n17310) );
  NOR2_X1 U20425 ( .A1(n17287), .A2(n17310), .ZN(n17313) );
  NAND2_X1 U20426 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17313), .ZN(n17306) );
  NOR2_X1 U20427 ( .A1(n17446), .A2(n17306), .ZN(n17304) );
  NAND2_X1 U20428 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17304), .ZN(n17292) );
  NOR2_X1 U20429 ( .A1(n17451), .A2(n17292), .ZN(n17295) );
  INV_X1 U20430 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17453) );
  AOI22_X1 U20431 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17345), .B1(n17295), .B2(
        n17453), .ZN(n17290) );
  OR3_X1 U20432 ( .A1(n17453), .A2(n17319), .A3(n17288), .ZN(n17289) );
  OAI211_X1 U20433 ( .C1(n17291), .C2(n17350), .A(n17290), .B(n17289), .ZN(
        P3_U2721) );
  INV_X1 U20434 ( .A(n17292), .ZN(n17299) );
  AOI21_X1 U20435 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17339), .A(n17299), .ZN(
        n17294) );
  OAI222_X1 U20436 ( .A1(n17343), .A2(n17296), .B1(n17295), .B2(n17294), .C1(
        n17350), .C2(n17293), .ZN(P3_U2722) );
  AOI21_X1 U20437 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17339), .A(n17304), .ZN(
        n17298) );
  OAI222_X1 U20438 ( .A1(n17343), .A2(n17300), .B1(n17299), .B2(n17298), .C1(
        n17350), .C2(n17297), .ZN(P3_U2723) );
  INV_X1 U20439 ( .A(n17306), .ZN(n17301) );
  AOI21_X1 U20440 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17339), .A(n17301), .ZN(
        n17303) );
  OAI222_X1 U20441 ( .A1(n17343), .A2(n17305), .B1(n17304), .B2(n17303), .C1(
        n17350), .C2(n17302), .ZN(P3_U2724) );
  NAND2_X1 U20442 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17345), .ZN(n17308) );
  OAI211_X1 U20443 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n17313), .A(n17339), .B(
        n17306), .ZN(n17307) );
  OAI211_X1 U20444 ( .C1(n17309), .C2(n17350), .A(n17308), .B(n17307), .ZN(
        P3_U2725) );
  INV_X1 U20445 ( .A(n17310), .ZN(n17323) );
  AOI22_X1 U20446 ( .A1(n17323), .A2(P3_EAX_REG_8__SCAN_IN), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n17339), .ZN(n17312) );
  OAI222_X1 U20447 ( .A1(n17343), .A2(n17314), .B1(n17313), .B2(n17312), .C1(
        n17350), .C2(n17311), .ZN(P3_U2726) );
  XOR2_X1 U20448 ( .A(n17315), .B(P3_EAX_REG_8__SCAN_IN), .Z(n17320) );
  AOI22_X1 U20449 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17345), .B1(n17317), .B2(
        n17316), .ZN(n17318) );
  OAI21_X1 U20450 ( .B1(n17320), .B2(n17319), .A(n17318), .ZN(P3_U2727) );
  INV_X1 U20451 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17436) );
  INV_X1 U20452 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17428) );
  NOR3_X1 U20453 ( .A1(n17346), .A2(n17428), .A3(n17337), .ZN(n17342) );
  NAND2_X1 U20454 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17342), .ZN(n17330) );
  NOR2_X1 U20455 ( .A1(n17432), .A2(n17330), .ZN(n17333) );
  NAND2_X1 U20456 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17333), .ZN(n17324) );
  NOR2_X1 U20457 ( .A1(n17436), .A2(n17324), .ZN(n17326) );
  AOI21_X1 U20458 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17339), .A(n17326), .ZN(
        n17322) );
  OAI222_X1 U20459 ( .A1(n18185), .A2(n17343), .B1(n17323), .B2(n17322), .C1(
        n17350), .C2(n17321), .ZN(P3_U2728) );
  INV_X1 U20460 ( .A(n17324), .ZN(n17329) );
  AOI21_X1 U20461 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17339), .A(n17329), .ZN(
        n17325) );
  OAI222_X1 U20462 ( .A1(n18181), .A2(n17343), .B1(n17326), .B2(n17325), .C1(
        n17350), .C2(n17746), .ZN(P3_U2729) );
  AOI21_X1 U20463 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17339), .A(n17333), .ZN(
        n17328) );
  OAI222_X1 U20464 ( .A1(n21103), .A2(n17343), .B1(n17329), .B2(n17328), .C1(
        n17350), .C2(n17327), .ZN(P3_U2730) );
  INV_X1 U20465 ( .A(n17330), .ZN(n17336) );
  AOI21_X1 U20466 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17339), .A(n17336), .ZN(
        n17332) );
  OAI222_X1 U20467 ( .A1(n18174), .A2(n17343), .B1(n17333), .B2(n17332), .C1(
        n17350), .C2(n17331), .ZN(P3_U2731) );
  AOI21_X1 U20468 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17339), .A(n17342), .ZN(
        n17335) );
  OAI222_X1 U20469 ( .A1(n18170), .A2(n17343), .B1(n17336), .B2(n17335), .C1(
        n17350), .C2(n17334), .ZN(P3_U2732) );
  NOR2_X1 U20470 ( .A1(n17346), .A2(n17337), .ZN(n17338) );
  AOI21_X1 U20471 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17339), .A(n17338), .ZN(
        n17341) );
  OAI222_X1 U20472 ( .A1(n18166), .A2(n17343), .B1(n17342), .B2(n17341), .C1(
        n17350), .C2(n17340), .ZN(P3_U2733) );
  AOI22_X1 U20473 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17345), .B1(n17344), .B2(
        P3_EAX_REG_1__SCAN_IN), .ZN(n17349) );
  OAI211_X1 U20474 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(P3_EAX_REG_0__SCAN_IN), 
        .A(n17347), .B(n17346), .ZN(n17348) );
  OAI211_X1 U20475 ( .C1(n11589), .C2(n17350), .A(n17349), .B(n17348), .ZN(
        P3_U2734) );
  INV_X1 U20476 ( .A(n17652), .ZN(n17818) );
  NOR2_X1 U20477 ( .A1(n18757), .A2(n17818), .ZN(n18804) );
  AND2_X1 U20478 ( .A1(n17379), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NAND2_X1 U20479 ( .A1(n17369), .A2(n17352), .ZN(n17368) );
  AOI22_X1 U20480 ( .A1(n18804), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17386), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17353) );
  OAI21_X1 U20481 ( .B1(n17422), .B2(n17368), .A(n17353), .ZN(P3_U2737) );
  INV_X1 U20482 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17420) );
  AOI22_X1 U20483 ( .A1(n18804), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17386), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17354) );
  OAI21_X1 U20484 ( .B1(n17420), .B2(n17368), .A(n17354), .ZN(P3_U2738) );
  INV_X1 U20485 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17418) );
  AOI22_X1 U20486 ( .A1(n18804), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17386), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17355) );
  OAI21_X1 U20487 ( .B1(n17418), .B2(n17368), .A(n17355), .ZN(P3_U2739) );
  AOI22_X1 U20488 ( .A1(n18804), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17379), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17356) );
  OAI21_X1 U20489 ( .B1(n17416), .B2(n17368), .A(n17356), .ZN(P3_U2740) );
  INV_X1 U20490 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17414) );
  AOI22_X1 U20491 ( .A1(n18804), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17379), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17357) );
  OAI21_X1 U20492 ( .B1(n17414), .B2(n17368), .A(n17357), .ZN(P3_U2741) );
  AOI22_X1 U20493 ( .A1(n18804), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17379), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17358) );
  OAI21_X1 U20494 ( .B1(n17412), .B2(n17368), .A(n17358), .ZN(P3_U2742) );
  AOI22_X1 U20495 ( .A1(n18804), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17379), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17359) );
  OAI21_X1 U20496 ( .B1(n17410), .B2(n17368), .A(n17359), .ZN(P3_U2743) );
  CLKBUF_X1 U20497 ( .A(n18804), .Z(n17387) );
  AOI22_X1 U20498 ( .A1(n17387), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17386), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17360) );
  OAI21_X1 U20499 ( .B1(n21079), .B2(n17368), .A(n17360), .ZN(P3_U2744) );
  INV_X1 U20500 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17407) );
  AOI22_X1 U20501 ( .A1(n17387), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17386), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17361) );
  OAI21_X1 U20502 ( .B1(n17407), .B2(n17368), .A(n17361), .ZN(P3_U2745) );
  AOI22_X1 U20503 ( .A1(n17387), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17386), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17362) );
  OAI21_X1 U20504 ( .B1(n17405), .B2(n17368), .A(n17362), .ZN(P3_U2746) );
  AOI22_X1 U20505 ( .A1(n17387), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17386), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17363) );
  OAI21_X1 U20506 ( .B1(n17403), .B2(n17368), .A(n17363), .ZN(P3_U2747) );
  AOI22_X1 U20507 ( .A1(n17387), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17386), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17364) );
  OAI21_X1 U20508 ( .B1(n17401), .B2(n17368), .A(n17364), .ZN(P3_U2748) );
  AOI22_X1 U20509 ( .A1(n17387), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17386), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17365) );
  OAI21_X1 U20510 ( .B1(n17399), .B2(n17368), .A(n17365), .ZN(P3_U2749) );
  AOI22_X1 U20511 ( .A1(n17387), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17386), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17366) );
  OAI21_X1 U20512 ( .B1(n17397), .B2(n17368), .A(n17366), .ZN(P3_U2750) );
  AOI22_X1 U20513 ( .A1(n17387), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17386), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17367) );
  OAI21_X1 U20514 ( .B1(n17395), .B2(n17368), .A(n17367), .ZN(P3_U2751) );
  INV_X1 U20515 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17458) );
  AOI22_X1 U20516 ( .A1(n17387), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17386), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17370) );
  OAI21_X1 U20517 ( .B1(n17458), .B2(n17389), .A(n17370), .ZN(P3_U2752) );
  AOI22_X1 U20518 ( .A1(n17387), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17386), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17371) );
  OAI21_X1 U20519 ( .B1(n17453), .B2(n17389), .A(n17371), .ZN(P3_U2753) );
  AOI22_X1 U20520 ( .A1(n17387), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17386), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17372) );
  OAI21_X1 U20521 ( .B1(n17451), .B2(n17389), .A(n17372), .ZN(P3_U2754) );
  INV_X1 U20522 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17449) );
  AOI22_X1 U20523 ( .A1(n17387), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17386), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17373) );
  OAI21_X1 U20524 ( .B1(n17449), .B2(n17389), .A(n17373), .ZN(P3_U2755) );
  AOI22_X1 U20525 ( .A1(n17387), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17379), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17374) );
  OAI21_X1 U20526 ( .B1(n17446), .B2(n17389), .A(n17374), .ZN(P3_U2756) );
  AOI22_X1 U20527 ( .A1(n17387), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17379), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17375) );
  OAI21_X1 U20528 ( .B1(n17444), .B2(n17389), .A(n17375), .ZN(P3_U2757) );
  INV_X1 U20529 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17442) );
  AOI22_X1 U20530 ( .A1(n17387), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17379), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17376) );
  OAI21_X1 U20531 ( .B1(n17442), .B2(n17389), .A(n17376), .ZN(P3_U2758) );
  INV_X1 U20532 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17440) );
  AOI22_X1 U20533 ( .A1(n17387), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17379), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17377) );
  OAI21_X1 U20534 ( .B1(n17440), .B2(n17389), .A(n17377), .ZN(P3_U2759) );
  INV_X1 U20535 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17438) );
  AOI22_X1 U20536 ( .A1(n17387), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17379), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17378) );
  OAI21_X1 U20537 ( .B1(n17438), .B2(n17389), .A(n17378), .ZN(P3_U2760) );
  AOI22_X1 U20538 ( .A1(n17387), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17379), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17380) );
  OAI21_X1 U20539 ( .B1(n17436), .B2(n17389), .A(n17380), .ZN(P3_U2761) );
  AOI22_X1 U20540 ( .A1(n17387), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17386), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17381) );
  OAI21_X1 U20541 ( .B1(n17434), .B2(n17389), .A(n17381), .ZN(P3_U2762) );
  AOI22_X1 U20542 ( .A1(n17387), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17386), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17382) );
  OAI21_X1 U20543 ( .B1(n17432), .B2(n17389), .A(n17382), .ZN(P3_U2763) );
  INV_X1 U20544 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17430) );
  AOI22_X1 U20545 ( .A1(n17387), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17386), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17383) );
  OAI21_X1 U20546 ( .B1(n17430), .B2(n17389), .A(n17383), .ZN(P3_U2764) );
  AOI22_X1 U20547 ( .A1(n17387), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17386), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17384) );
  OAI21_X1 U20548 ( .B1(n17428), .B2(n17389), .A(n17384), .ZN(P3_U2765) );
  INV_X1 U20549 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17426) );
  AOI22_X1 U20550 ( .A1(n17387), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17386), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17385) );
  OAI21_X1 U20551 ( .B1(n17426), .B2(n17389), .A(n17385), .ZN(P3_U2766) );
  AOI22_X1 U20552 ( .A1(n17387), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17386), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17388) );
  OAI21_X1 U20553 ( .B1(n17424), .B2(n17389), .A(n17388), .ZN(P3_U2767) );
  INV_X1 U20554 ( .A(n17390), .ZN(n17392) );
  INV_X2 U20555 ( .A(n17393), .ZN(n17454) );
  AOI22_X1 U20556 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17454), .ZN(n17394) );
  OAI21_X1 U20557 ( .B1(n17395), .B2(n17457), .A(n17394), .ZN(P3_U2768) );
  AOI22_X1 U20558 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17454), .ZN(n17396) );
  OAI21_X1 U20559 ( .B1(n17397), .B2(n17457), .A(n17396), .ZN(P3_U2769) );
  AOI22_X1 U20560 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17454), .ZN(n17398) );
  OAI21_X1 U20561 ( .B1(n17399), .B2(n17457), .A(n17398), .ZN(P3_U2770) );
  AOI22_X1 U20562 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17447), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17454), .ZN(n17400) );
  OAI21_X1 U20563 ( .B1(n17401), .B2(n17457), .A(n17400), .ZN(P3_U2771) );
  AOI22_X1 U20564 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17447), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17454), .ZN(n17402) );
  OAI21_X1 U20565 ( .B1(n17403), .B2(n17457), .A(n17402), .ZN(P3_U2772) );
  AOI22_X1 U20566 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17447), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17454), .ZN(n17404) );
  OAI21_X1 U20567 ( .B1(n17405), .B2(n17457), .A(n17404), .ZN(P3_U2773) );
  AOI22_X1 U20568 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17447), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17454), .ZN(n17406) );
  OAI21_X1 U20569 ( .B1(n17407), .B2(n17457), .A(n17406), .ZN(P3_U2774) );
  AOI22_X1 U20570 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17447), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17454), .ZN(n17408) );
  OAI21_X1 U20571 ( .B1(n21079), .B2(n17457), .A(n17408), .ZN(P3_U2775) );
  AOI22_X1 U20572 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17447), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17454), .ZN(n17409) );
  OAI21_X1 U20573 ( .B1(n17410), .B2(n17457), .A(n17409), .ZN(P3_U2776) );
  AOI22_X1 U20574 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17447), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17454), .ZN(n17411) );
  OAI21_X1 U20575 ( .B1(n17412), .B2(n17457), .A(n17411), .ZN(P3_U2777) );
  AOI22_X1 U20576 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17447), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17454), .ZN(n17413) );
  OAI21_X1 U20577 ( .B1(n17414), .B2(n17457), .A(n17413), .ZN(P3_U2778) );
  AOI22_X1 U20578 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17447), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17454), .ZN(n17415) );
  OAI21_X1 U20579 ( .B1(n17416), .B2(n17457), .A(n17415), .ZN(P3_U2779) );
  AOI22_X1 U20580 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17454), .ZN(n17417) );
  OAI21_X1 U20581 ( .B1(n17418), .B2(n17457), .A(n17417), .ZN(P3_U2780) );
  AOI22_X1 U20582 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17454), .ZN(n17419) );
  OAI21_X1 U20583 ( .B1(n17420), .B2(n17457), .A(n17419), .ZN(P3_U2781) );
  AOI22_X1 U20584 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17454), .ZN(n17421) );
  OAI21_X1 U20585 ( .B1(n17422), .B2(n17457), .A(n17421), .ZN(P3_U2782) );
  AOI22_X1 U20586 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17454), .ZN(n17423) );
  OAI21_X1 U20587 ( .B1(n17424), .B2(n17457), .A(n17423), .ZN(P3_U2783) );
  AOI22_X1 U20588 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17454), .ZN(n17425) );
  OAI21_X1 U20589 ( .B1(n17426), .B2(n17457), .A(n17425), .ZN(P3_U2784) );
  AOI22_X1 U20590 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17454), .ZN(n17427) );
  OAI21_X1 U20591 ( .B1(n17428), .B2(n17457), .A(n17427), .ZN(P3_U2785) );
  AOI22_X1 U20592 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17454), .ZN(n17429) );
  OAI21_X1 U20593 ( .B1(n17430), .B2(n17457), .A(n17429), .ZN(P3_U2786) );
  AOI22_X1 U20594 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17454), .ZN(n17431) );
  OAI21_X1 U20595 ( .B1(n17432), .B2(n17457), .A(n17431), .ZN(P3_U2787) );
  AOI22_X1 U20596 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17454), .ZN(n17433) );
  OAI21_X1 U20597 ( .B1(n17434), .B2(n17457), .A(n17433), .ZN(P3_U2788) );
  AOI22_X1 U20598 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17454), .ZN(n17435) );
  OAI21_X1 U20599 ( .B1(n17436), .B2(n17457), .A(n17435), .ZN(P3_U2789) );
  AOI22_X1 U20600 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17454), .ZN(n17437) );
  OAI21_X1 U20601 ( .B1(n17438), .B2(n17457), .A(n17437), .ZN(P3_U2790) );
  AOI22_X1 U20602 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17454), .ZN(n17439) );
  OAI21_X1 U20603 ( .B1(n17440), .B2(n17457), .A(n17439), .ZN(P3_U2791) );
  AOI22_X1 U20604 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17454), .ZN(n17441) );
  OAI21_X1 U20605 ( .B1(n17442), .B2(n17457), .A(n17441), .ZN(P3_U2792) );
  AOI22_X1 U20606 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17447), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17454), .ZN(n17443) );
  OAI21_X1 U20607 ( .B1(n17444), .B2(n17457), .A(n17443), .ZN(P3_U2793) );
  AOI22_X1 U20608 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17454), .ZN(n17445) );
  OAI21_X1 U20609 ( .B1(n17446), .B2(n17457), .A(n17445), .ZN(P3_U2794) );
  AOI22_X1 U20610 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17447), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17454), .ZN(n17448) );
  OAI21_X1 U20611 ( .B1(n17449), .B2(n17457), .A(n17448), .ZN(P3_U2795) );
  AOI22_X1 U20612 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17454), .ZN(n17450) );
  OAI21_X1 U20613 ( .B1(n17451), .B2(n17457), .A(n17450), .ZN(P3_U2796) );
  AOI22_X1 U20614 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17454), .ZN(n17452) );
  OAI21_X1 U20615 ( .B1(n17453), .B2(n17457), .A(n17452), .ZN(P3_U2797) );
  AOI22_X1 U20616 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17454), .ZN(n17456) );
  OAI21_X1 U20617 ( .B1(n17458), .B2(n17457), .A(n17456), .ZN(P3_U2798) );
  INV_X1 U20618 ( .A(n17459), .ZN(n17480) );
  OAI21_X1 U20619 ( .B1(n17460), .B2(n17715), .A(n17817), .ZN(n17461) );
  AOI21_X1 U20620 ( .B1(n17652), .B2(n17462), .A(n17461), .ZN(n17498) );
  OAI21_X1 U20621 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17603), .A(
        n17498), .ZN(n17482) );
  NOR2_X1 U20622 ( .A1(n17685), .A2(n17806), .ZN(n17575) );
  OAI22_X1 U20623 ( .A1(n17464), .A2(n17725), .B1(n17463), .B2(n17822), .ZN(
        n17500) );
  NOR2_X1 U20624 ( .A1(n20889), .A2(n17500), .ZN(n17466) );
  NOR3_X1 U20625 ( .A1(n17575), .A2(n17466), .A3(n17465), .ZN(n17474) );
  NAND2_X1 U20626 ( .A1(n18126), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17471) );
  NOR2_X1 U20627 ( .A1(n17661), .A2(n17468), .ZN(n17487) );
  NAND2_X1 U20628 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17469) );
  OAI211_X1 U20629 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17487), .B(n17469), .ZN(n17470) );
  OAI211_X1 U20630 ( .C1(n17667), .C2(n17472), .A(n17471), .B(n17470), .ZN(
        n17473) );
  AOI211_X1 U20631 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n17482), .A(
        n17474), .B(n17473), .ZN(n17479) );
  OAI211_X1 U20632 ( .C1(n17477), .C2(n17476), .A(n17697), .B(n17475), .ZN(
        n17478) );
  OAI211_X1 U20633 ( .C1(n17480), .C2(n17625), .A(n17479), .B(n17478), .ZN(
        P3_U2802) );
  AOI22_X1 U20634 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17482), .B1(
        n17655), .B2(n17481), .ZN(n17491) );
  NAND2_X1 U20635 ( .A1(n17484), .A2(n17483), .ZN(n17485) );
  XNOR2_X1 U20636 ( .A(n10101), .B(n17485), .ZN(n17833) );
  AOI22_X1 U20637 ( .A1(n17697), .A2(n17833), .B1(n17487), .B2(n17486), .ZN(
        n17490) );
  AOI22_X1 U20638 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17500), .B1(
        n17488), .B2(n20889), .ZN(n17489) );
  NAND2_X1 U20639 ( .A1(n18126), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17834) );
  NAND4_X1 U20640 ( .A1(n17491), .A2(n17490), .A3(n17489), .A4(n17834), .ZN(
        P3_U2803) );
  AOI21_X1 U20641 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17493), .A(
        n17492), .ZN(n17844) );
  NAND2_X1 U20642 ( .A1(n17512), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17838) );
  NOR2_X1 U20643 ( .A1(n17625), .A2(n17838), .ZN(n17501) );
  INV_X2 U20644 ( .A(n18499), .ZN(n18471) );
  AOI21_X1 U20645 ( .B1(n17494), .B2(n18471), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17497) );
  OAI21_X1 U20646 ( .B1(n17655), .B2(n17573), .A(n17495), .ZN(n17496) );
  NAND2_X1 U20647 ( .A1(n18126), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17842) );
  OAI211_X1 U20648 ( .C1(n17498), .C2(n17497), .A(n17496), .B(n17842), .ZN(
        n17499) );
  AOI221_X1 U20649 ( .B1(n17501), .B2(n17831), .C1(n17500), .C2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(n17499), .ZN(n17502) );
  OAI21_X1 U20650 ( .B1(n17844), .B2(n17726), .A(n17502), .ZN(P3_U2804) );
  NAND2_X1 U20651 ( .A1(n17512), .A2(n17953), .ZN(n17503) );
  XNOR2_X1 U20652 ( .A(n17503), .B(n17850), .ZN(n17857) );
  AOI21_X1 U20653 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17532), .A(
        n17818), .ZN(n17504) );
  AOI211_X1 U20654 ( .C1(n18471), .C2(n17505), .A(n17774), .B(n17504), .ZN(
        n17536) );
  OAI21_X1 U20655 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17603), .A(
        n17536), .ZN(n17521) );
  NAND2_X1 U20656 ( .A1(n18126), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n17849) );
  NOR2_X1 U20657 ( .A1(n17661), .A2(n17505), .ZN(n17523) );
  OAI211_X1 U20658 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17523), .B(n17506), .ZN(n17507) );
  OAI211_X1 U20659 ( .C1(n17667), .C2(n17508), .A(n17849), .B(n17507), .ZN(
        n17515) );
  OAI21_X1 U20660 ( .B1(n10101), .B2(n17510), .A(n17509), .ZN(n17511) );
  XNOR2_X1 U20661 ( .A(n17511), .B(n17850), .ZN(n17851) );
  INV_X1 U20662 ( .A(n17878), .ZN(n17952) );
  AND2_X1 U20663 ( .A1(n17512), .A2(n17952), .ZN(n17513) );
  OAI22_X1 U20664 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17513), .B1(
        n17838), .B2(n17878), .ZN(n17852) );
  OAI22_X1 U20665 ( .A1(n17726), .A2(n17851), .B1(n17822), .B2(n17852), .ZN(
        n17514) );
  AOI211_X1 U20666 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17521), .A(
        n17515), .B(n17514), .ZN(n17516) );
  OAI21_X1 U20667 ( .B1(n17725), .B2(n17857), .A(n17516), .ZN(P3_U2805) );
  AOI21_X1 U20668 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17518), .A(
        n17517), .ZN(n17870) );
  OAI22_X1 U20669 ( .A1(n18138), .A2(n18716), .B1(n17667), .B2(n17519), .ZN(
        n17520) );
  AOI221_X1 U20670 ( .B1(n17523), .B2(n17522), .C1(n17521), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17520), .ZN(n17527) );
  NOR2_X1 U20671 ( .A1(n17524), .A2(n17878), .ZN(n17859) );
  OAI22_X1 U20672 ( .A1(n17860), .A2(n17725), .B1(n17859), .B2(n17822), .ZN(
        n17538) );
  INV_X1 U20673 ( .A(n17625), .ZN(n17525) );
  NOR2_X1 U20674 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17524), .ZN(
        n17858) );
  AOI22_X1 U20675 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17538), .B1(
        n17525), .B2(n17858), .ZN(n17526) );
  OAI211_X1 U20676 ( .C1(n17870), .C2(n17726), .A(n17527), .B(n17526), .ZN(
        P3_U2806) );
  AOI22_X1 U20677 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n10101), .B1(
        n17529), .B2(n17542), .ZN(n17530) );
  NAND2_X1 U20678 ( .A1(n17528), .A2(n17530), .ZN(n17531) );
  XNOR2_X1 U20679 ( .A(n17531), .B(n17863), .ZN(n17876) );
  NOR2_X1 U20680 ( .A1(n17871), .A2(n17625), .ZN(n17539) );
  AOI21_X1 U20681 ( .B1(n17532), .B2(n18471), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17535) );
  OAI21_X1 U20682 ( .B1(n17655), .B2(n17573), .A(n17533), .ZN(n17534) );
  NAND2_X1 U20683 ( .A1(n18140), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17875) );
  OAI211_X1 U20684 ( .C1(n17536), .C2(n17535), .A(n17534), .B(n17875), .ZN(
        n17537) );
  AOI221_X1 U20685 ( .B1(n17539), .B2(n17863), .C1(n17538), .C2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n17537), .ZN(n17540) );
  OAI21_X1 U20686 ( .B1(n17726), .B2(n17876), .A(n17540), .ZN(P3_U2807) );
  INV_X1 U20687 ( .A(n17528), .ZN(n17541) );
  AOI221_X1 U20688 ( .B1(n17886), .B2(n17542), .C1(n11609), .C2(n17542), .A(
        n17541), .ZN(n17543) );
  XNOR2_X1 U20689 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n17543), .ZN(
        n17893) );
  NOR2_X1 U20690 ( .A1(n17886), .A2(n17625), .ZN(n17553) );
  INV_X1 U20691 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17885) );
  AOI22_X1 U20692 ( .A1(n17685), .A2(n11609), .B1(n17806), .B2(n17878), .ZN(
        n17624) );
  OAI21_X1 U20693 ( .B1(n17544), .B2(n17575), .A(n17624), .ZN(n17565) );
  OAI21_X1 U20694 ( .B1(n17545), .B2(n17818), .A(n17817), .ZN(n17546) );
  AOI21_X1 U20695 ( .B1(n17776), .B2(n17548), .A(n17546), .ZN(n17571) );
  OAI21_X1 U20696 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17603), .A(
        n17571), .ZN(n17558) );
  AOI22_X1 U20697 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17558), .B1(
        n17655), .B2(n17547), .ZN(n17551) );
  NOR2_X1 U20698 ( .A1(n17661), .A2(n17548), .ZN(n17560) );
  OAI211_X1 U20699 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17560), .B(n17549), .ZN(n17550) );
  OAI211_X1 U20700 ( .C1(n18712), .C2(n18138), .A(n17551), .B(n17550), .ZN(
        n17552) );
  AOI221_X1 U20701 ( .B1(n17553), .B2(n17885), .C1(n17565), .C2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n17552), .ZN(n17554) );
  OAI21_X1 U20702 ( .B1(n17726), .B2(n17893), .A(n17554), .ZN(P3_U2808) );
  NAND3_X1 U20703 ( .A1(n17585), .A2(n17898), .A3(n17555), .ZN(n17902) );
  OAI22_X1 U20704 ( .A1(n18138), .A2(n18711), .B1(n17667), .B2(n9962), .ZN(
        n17557) );
  AOI221_X1 U20705 ( .B1(n17560), .B2(n17559), .C1(n17558), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17557), .ZN(n17567) );
  INV_X1 U20706 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17882) );
  NOR3_X1 U20707 ( .A1(n10101), .A2(n17882), .A3(n17561), .ZN(n17581) );
  INV_X1 U20708 ( .A(n17562), .ZN(n17582) );
  AOI22_X1 U20709 ( .A1(n17898), .A2(n17581), .B1(n17582), .B2(n17563), .ZN(
        n17564) );
  XNOR2_X1 U20710 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17564), .ZN(
        n17894) );
  AOI22_X1 U20711 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17565), .B1(
        n17697), .B2(n17894), .ZN(n17566) );
  OAI211_X1 U20712 ( .C1(n17625), .C2(n17902), .A(n17567), .B(n17566), .ZN(
        P3_U2809) );
  NOR2_X1 U20713 ( .A1(n17896), .A2(n17584), .ZN(n17906) );
  NAND2_X1 U20714 ( .A1(n17906), .A2(n17568), .ZN(n17912) );
  INV_X1 U20715 ( .A(n17603), .ZN(n17573) );
  AOI21_X1 U20716 ( .B1(n17569), .B2(n18471), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17570) );
  OAI22_X1 U20717 ( .A1(n17571), .A2(n17570), .B1(n18138), .B2(n18708), .ZN(
        n17572) );
  AOI221_X1 U20718 ( .B1(n17655), .B2(n17574), .C1(n17573), .C2(n17574), .A(
        n17572), .ZN(n17578) );
  OAI21_X1 U20719 ( .B1(n17575), .B2(n17906), .A(n17624), .ZN(n17587) );
  OAI221_X1 U20720 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17598), 
        .C1(n17584), .C2(n17581), .A(n17528), .ZN(n17576) );
  XNOR2_X1 U20721 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17576), .ZN(
        n17903) );
  AOI22_X1 U20722 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17587), .B1(
        n17697), .B2(n17903), .ZN(n17577) );
  OAI211_X1 U20723 ( .C1(n17625), .C2(n17912), .A(n17578), .B(n17577), .ZN(
        P3_U2810) );
  AOI21_X1 U20724 ( .B1(n17776), .B2(n17588), .A(n17774), .ZN(n17605) );
  OAI21_X1 U20725 ( .B1(n17579), .B2(n17818), .A(n17605), .ZN(n17595) );
  AOI22_X1 U20726 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n17595), .B1(
        n17655), .B2(n17580), .ZN(n17592) );
  AOI21_X1 U20727 ( .B1(n17582), .B2(n17598), .A(n17581), .ZN(n17583) );
  XNOR2_X1 U20728 ( .A(n17583), .B(n17584), .ZN(n17918) );
  NAND2_X1 U20729 ( .A1(n17585), .A2(n17584), .ZN(n17913) );
  OAI22_X1 U20730 ( .A1(n17918), .A2(n17726), .B1(n17625), .B2(n17913), .ZN(
        n17586) );
  AOI21_X1 U20731 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17587), .A(
        n17586), .ZN(n17591) );
  NAND2_X1 U20732 ( .A1(n18140), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n17916) );
  NOR2_X1 U20733 ( .A1(n17661), .A2(n17588), .ZN(n17597) );
  OAI211_X1 U20734 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17597), .B(n17589), .ZN(n17590) );
  NAND4_X1 U20735 ( .A1(n17592), .A2(n17591), .A3(n17916), .A4(n17590), .ZN(
        P3_U2811) );
  NAND2_X1 U20736 ( .A1(n17923), .A2(n17882), .ZN(n17930) );
  OAI22_X1 U20737 ( .A1(n18138), .A2(n18704), .B1(n17667), .B2(n17593), .ZN(
        n17594) );
  AOI221_X1 U20738 ( .B1(n17597), .B2(n17596), .C1(n17595), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17594), .ZN(n17601) );
  OAI21_X1 U20739 ( .B1(n17923), .B2(n17625), .A(n17624), .ZN(n17610) );
  AOI21_X1 U20740 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n17724), .A(
        n17598), .ZN(n17599) );
  XNOR2_X1 U20741 ( .A(n17599), .B(n17562), .ZN(n17926) );
  AOI22_X1 U20742 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17610), .B1(
        n17697), .B2(n17926), .ZN(n17600) );
  OAI211_X1 U20743 ( .C1(n17625), .C2(n17930), .A(n17601), .B(n17600), .ZN(
        P3_U2812) );
  NAND2_X1 U20744 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17931), .ZN(
        n17937) );
  AOI21_X1 U20745 ( .B1(n17602), .B2(n18471), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17606) );
  OAI22_X1 U20746 ( .A1(n17606), .A2(n17605), .B1(n17800), .B2(n17604), .ZN(
        n17607) );
  AOI21_X1 U20747 ( .B1(n18126), .B2(P3_REIP_REG_17__SCAN_IN), .A(n17607), 
        .ZN(n17612) );
  OAI21_X1 U20748 ( .B1(n17609), .B2(n17931), .A(n17608), .ZN(n17935) );
  AOI22_X1 U20749 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17610), .B1(
        n17697), .B2(n17935), .ZN(n17611) );
  OAI211_X1 U20750 ( .C1(n17625), .C2(n17937), .A(n17612), .B(n17611), .ZN(
        P3_U2813) );
  NAND2_X1 U20751 ( .A1(n17724), .A2(n18011), .ZN(n17702) );
  OAI21_X1 U20752 ( .B1(n10088), .B2(n17702), .A(n17614), .ZN(n17615) );
  XNOR2_X1 U20753 ( .A(n17615), .B(n17947), .ZN(n17944) );
  AOI21_X1 U20754 ( .B1(n17776), .B2(n17618), .A(n17774), .ZN(n17643) );
  OAI21_X1 U20755 ( .B1(n17616), .B2(n17818), .A(n17643), .ZN(n17631) );
  AOI22_X1 U20756 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17631), .B1(
        n17655), .B2(n17617), .ZN(n17621) );
  NOR2_X1 U20757 ( .A1(n17661), .A2(n17618), .ZN(n17628) );
  OAI211_X1 U20758 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17628), .B(n17619), .ZN(n17620) );
  OAI211_X1 U20759 ( .C1(n20890), .C2(n18138), .A(n17621), .B(n17620), .ZN(
        n17622) );
  AOI21_X1 U20760 ( .B1(n17697), .B2(n17944), .A(n17622), .ZN(n17623) );
  OAI221_X1 U20761 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17625), 
        .C1(n17947), .C2(n17624), .A(n17623), .ZN(P3_U2814) );
  NOR2_X1 U20762 ( .A1(n17952), .A2(n17822), .ZN(n17629) );
  NAND3_X1 U20763 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17637), .A3(
        n17626), .ZN(n17646) );
  NAND2_X1 U20764 ( .A1(n17950), .A2(n17646), .ZN(n17957) );
  AOI22_X1 U20765 ( .A1(n17629), .A2(n17957), .B1(n17628), .B2(n17627), .ZN(
        n17636) );
  AOI22_X1 U20766 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17631), .B1(
        n17655), .B2(n17630), .ZN(n17635) );
  INV_X1 U20767 ( .A(n17658), .ZN(n17984) );
  NOR3_X1 U20768 ( .A1(n21186), .A2(n17984), .A3(n17702), .ZN(n17644) );
  NAND2_X1 U20769 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17991), .ZN(
        n17980) );
  OAI221_X1 U20770 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n9865), .C1(
        n17971), .C2(n17644), .A(n17980), .ZN(n17632) );
  XNOR2_X1 U20771 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17632), .ZN(
        n17960) );
  NOR2_X1 U20772 ( .A1(n17953), .A2(n17725), .ZN(n17633) );
  NAND3_X1 U20773 ( .A1(n18011), .A2(n17637), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17638) );
  NAND2_X1 U20774 ( .A1(n17950), .A2(n17638), .ZN(n17955) );
  AOI22_X1 U20775 ( .A1(n17697), .A2(n17960), .B1(n17633), .B2(n17955), .ZN(
        n17634) );
  NAND2_X1 U20776 ( .A1(n18126), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n17961) );
  NAND4_X1 U20777 ( .A1(n17636), .A2(n17635), .A3(n17634), .A4(n17961), .ZN(
        P3_U2815) );
  INV_X1 U20778 ( .A(n17637), .ZN(n17970) );
  NOR2_X1 U20779 ( .A1(n17723), .A2(n17970), .ZN(n17639) );
  OAI21_X1 U20780 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17639), .A(
        n17638), .ZN(n17978) );
  AOI21_X1 U20781 ( .B1(n18471), .B2(n17640), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17642) );
  OAI22_X1 U20782 ( .A1(n17643), .A2(n17642), .B1(n17800), .B2(n17641), .ZN(
        n17649) );
  OAI21_X1 U20783 ( .B1(n9865), .B2(n17644), .A(n17980), .ZN(n17645) );
  XNOR2_X1 U20784 ( .A(n17645), .B(n17971), .ZN(n17972) );
  NOR2_X1 U20785 ( .A1(n18008), .A2(n17970), .ZN(n17647) );
  OAI21_X1 U20786 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17647), .A(
        n17646), .ZN(n17973) );
  OAI22_X1 U20787 ( .A1(n17726), .A2(n17972), .B1(n17822), .B2(n17973), .ZN(
        n17648) );
  AOI211_X1 U20788 ( .C1(n18126), .C2(P3_REIP_REG_14__SCAN_IN), .A(n17649), 
        .B(n17648), .ZN(n17650) );
  OAI21_X1 U20789 ( .B1(n17725), .B2(n17978), .A(n17650), .ZN(P3_U2816) );
  AOI22_X1 U20790 ( .A1(n17652), .A2(n17651), .B1(n17776), .B2(n17660), .ZN(
        n17653) );
  NAND2_X1 U20791 ( .A1(n17653), .A2(n17817), .ZN(n17669) );
  AOI22_X1 U20792 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17669), .B1(
        n17655), .B2(n17654), .ZN(n17665) );
  NOR2_X1 U20793 ( .A1(n17723), .A2(n17965), .ZN(n17983) );
  NOR2_X1 U20794 ( .A1(n18008), .A2(n17965), .ZN(n17986) );
  OAI22_X1 U20795 ( .A1(n17983), .A2(n17725), .B1(n17986), .B2(n17822), .ZN(
        n17674) );
  AOI21_X1 U20796 ( .B1(n21186), .B2(n10101), .A(n17983), .ZN(n17656) );
  AOI21_X1 U20797 ( .B1(n10101), .B2(n17672), .A(n17656), .ZN(n17657) );
  XNOR2_X1 U20798 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n17657), .ZN(
        n17997) );
  NAND2_X1 U20799 ( .A1(n17658), .A2(n17713), .ZN(n17677) );
  OAI22_X1 U20800 ( .A1(n17726), .A2(n17997), .B1(n17980), .B2(n17677), .ZN(
        n17659) );
  AOI21_X1 U20801 ( .B1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n17674), .A(
        n17659), .ZN(n17664) );
  NAND2_X1 U20802 ( .A1(n18126), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n17995) );
  NOR2_X1 U20803 ( .A1(n17661), .A2(n17660), .ZN(n17671) );
  OAI211_X1 U20804 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17671), .B(n17662), .ZN(n17663) );
  NAND4_X1 U20805 ( .A1(n17665), .A2(n17664), .A3(n17995), .A4(n17663), .ZN(
        P3_U2817) );
  INV_X1 U20806 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17670) );
  NAND2_X1 U20807 ( .A1(n18140), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18002) );
  OAI21_X1 U20808 ( .B1(n17667), .B2(n17666), .A(n18002), .ZN(n17668) );
  AOI221_X1 U20809 ( .B1(n17671), .B2(n17670), .C1(n17669), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n17668), .ZN(n17676) );
  OAI21_X1 U20810 ( .B1(n17984), .B2(n17702), .A(n17672), .ZN(n17673) );
  XNOR2_X1 U20811 ( .A(n17673), .B(n21186), .ZN(n18001) );
  AOI22_X1 U20812 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17674), .B1(
        n17697), .B2(n18001), .ZN(n17675) );
  OAI211_X1 U20813 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n17677), .A(
        n17676), .B(n17675), .ZN(P3_U2818) );
  NOR2_X1 U20814 ( .A1(n18021), .A2(n17702), .ZN(n17693) );
  AOI21_X1 U20815 ( .B1(n17693), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n17678), .ZN(n17680) );
  XNOR2_X1 U20816 ( .A(n17680), .B(n17679), .ZN(n18019) );
  NAND3_X1 U20817 ( .A1(n18471), .A2(n17716), .A3(n17681), .ZN(n17690) );
  AND2_X1 U20818 ( .A1(n17804), .A2(n17690), .ZN(n17691) );
  NOR2_X1 U20819 ( .A1(n18138), .A2(n20924), .ZN(n17684) );
  OAI22_X1 U20820 ( .A1(n17800), .A2(n17682), .B1(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17690), .ZN(n17683) );
  AOI211_X1 U20821 ( .C1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n17691), .A(
        n17684), .B(n17683), .ZN(n17688) );
  AOI22_X1 U20822 ( .A1(n17685), .A2(n17723), .B1(n17806), .B2(n18008), .ZN(
        n17710) );
  NAND2_X1 U20823 ( .A1(n18014), .A2(n17713), .ZN(n17686) );
  NAND2_X1 U20824 ( .A1(n17710), .A2(n17686), .ZN(n17698) );
  NOR2_X1 U20825 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18014), .ZN(
        n18006) );
  AOI22_X1 U20826 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17698), .B1(
        n18006), .B2(n17713), .ZN(n17687) );
  OAI211_X1 U20827 ( .C1(n18019), .C2(n17726), .A(n17688), .B(n17687), .ZN(
        P3_U2819) );
  INV_X1 U20828 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17689) );
  NAND2_X1 U20829 ( .A1(n18471), .A2(n17716), .ZN(n17734) );
  NOR3_X1 U20830 ( .A1(n17719), .A2(n17689), .A3(n17734), .ZN(n17709) );
  AOI22_X1 U20831 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17691), .B1(
        n17709), .B2(n17690), .ZN(n17701) );
  INV_X1 U20832 ( .A(n17692), .ZN(n17694) );
  NOR2_X1 U20833 ( .A1(n17694), .A2(n17693), .ZN(n17695) );
  XNOR2_X1 U20834 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n17695), .ZN(
        n18023) );
  AOI22_X1 U20835 ( .A1(n17697), .A2(n18023), .B1(n17696), .B2(n17808), .ZN(
        n17700) );
  OAI221_X1 U20836 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n17713), .A(n17698), .ZN(
        n17699) );
  NAND2_X1 U20837 ( .A1(n18140), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n18030) );
  NAND4_X1 U20838 ( .A1(n17701), .A2(n17700), .A3(n17699), .A4(n18030), .ZN(
        P3_U2820) );
  INV_X1 U20839 ( .A(n17702), .ZN(n17704) );
  NOR2_X1 U20840 ( .A1(n17704), .A2(n17703), .ZN(n17705) );
  XNOR2_X1 U20841 ( .A(n17705), .B(n18021), .ZN(n18042) );
  NAND2_X1 U20842 ( .A1(n18140), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n18040) );
  OAI21_X1 U20843 ( .B1(n17800), .B2(n17706), .A(n18040), .ZN(n17712) );
  NOR2_X1 U20844 ( .A1(n17719), .A2(n17734), .ZN(n17707) );
  AOI21_X1 U20845 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17804), .A(
        n17707), .ZN(n17708) );
  OAI22_X1 U20846 ( .A1(n17710), .A2(n18021), .B1(n17709), .B2(n17708), .ZN(
        n17711) );
  AOI211_X1 U20847 ( .C1(n18021), .C2(n17713), .A(n17712), .B(n17711), .ZN(
        n17714) );
  OAI21_X1 U20848 ( .B1(n18042), .B2(n17726), .A(n17714), .ZN(P3_U2821) );
  OAI21_X1 U20849 ( .B1(n17716), .B2(n17715), .A(n17817), .ZN(n17738) );
  OAI21_X1 U20850 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17718), .A(
        n17717), .ZN(n18044) );
  NAND2_X1 U20851 ( .A1(n18126), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n18061) );
  OAI211_X1 U20852 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17720), .A(
        n18471), .B(n17719), .ZN(n17721) );
  OAI211_X1 U20853 ( .C1(n17822), .C2(n18044), .A(n18061), .B(n17721), .ZN(
        n17728) );
  NAND2_X1 U20854 ( .A1(n17723), .A2(n17722), .ZN(n18043) );
  XNOR2_X1 U20855 ( .A(n17724), .B(n18043), .ZN(n18046) );
  OAI22_X1 U20856 ( .A1(n18046), .A2(n17726), .B1(n17725), .B2(n18043), .ZN(
        n17727) );
  AOI211_X1 U20857 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17738), .A(
        n17728), .B(n17727), .ZN(n17729) );
  OAI21_X1 U20858 ( .B1(n17800), .B2(n17730), .A(n17729), .ZN(P3_U2822) );
  NOR2_X1 U20859 ( .A1(n17732), .A2(n17731), .ZN(n17733) );
  XNOR2_X1 U20860 ( .A(n17733), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18066) );
  OAI22_X1 U20861 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n17734), .B1(
        n18066), .B2(n17822), .ZN(n17735) );
  AOI21_X1 U20862 ( .B1(n18126), .B2(P3_REIP_REG_7__SCAN_IN), .A(n17735), .ZN(
        n17740) );
  AOI21_X1 U20863 ( .B1(n18071), .B2(n17737), .A(n17736), .ZN(n18069) );
  AOI22_X1 U20864 ( .A1(n9848), .A2(n18069), .B1(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17738), .ZN(n17739) );
  OAI211_X1 U20865 ( .C1(n17800), .C2(n17741), .A(n17740), .B(n17739), .ZN(
        P3_U2823) );
  OAI21_X1 U20866 ( .B1(n17742), .B2(n18499), .A(n17804), .ZN(n17767) );
  OR2_X1 U20867 ( .A1(n18499), .A2(n17742), .ZN(n17750) );
  INV_X1 U20868 ( .A(n17745), .ZN(n17743) );
  AOI22_X1 U20869 ( .A1(n17745), .A2(n17761), .B1(n17744), .B2(n17743), .ZN(
        n17749) );
  AOI22_X1 U20870 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17747), .B1(
        n17746), .B2(n18064), .ZN(n17748) );
  XNOR2_X1 U20871 ( .A(n17749), .B(n17748), .ZN(n18079) );
  OAI22_X1 U20872 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17750), .B1(
        n18079), .B2(n17822), .ZN(n17751) );
  AOI21_X1 U20873 ( .B1(n18126), .B2(P3_REIP_REG_6__SCAN_IN), .A(n17751), .ZN(
        n17756) );
  AOI21_X1 U20874 ( .B1(n9934), .B2(n17753), .A(n17752), .ZN(n18076) );
  AOI22_X1 U20875 ( .A1(n9848), .A2(n18076), .B1(n17754), .B2(n17808), .ZN(
        n17755) );
  OAI211_X1 U20876 ( .C1(n17757), .C2(n17767), .A(n17756), .B(n17755), .ZN(
        P3_U2824) );
  AOI21_X1 U20877 ( .B1(n17758), .B2(n17817), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17768) );
  AOI21_X1 U20878 ( .B1(n18088), .B2(n17760), .A(n17759), .ZN(n18081) );
  AOI22_X1 U20879 ( .A1(n9848), .A2(n18081), .B1(n18140), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17766) );
  AOI21_X1 U20880 ( .B1(n17763), .B2(n17762), .A(n17761), .ZN(n18085) );
  AOI22_X1 U20881 ( .A1(n17806), .A2(n18085), .B1(n17764), .B2(n17808), .ZN(
        n17765) );
  OAI211_X1 U20882 ( .C1(n17768), .C2(n17767), .A(n17766), .B(n17765), .ZN(
        P3_U2825) );
  AOI21_X1 U20883 ( .B1(n17771), .B2(n17770), .A(n17769), .ZN(n18090) );
  AOI22_X1 U20884 ( .A1(n18126), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n17806), 
        .B2(n18090), .ZN(n17781) );
  AOI21_X1 U20885 ( .B1(n9939), .B2(n17773), .A(n17772), .ZN(n18093) );
  AOI21_X1 U20886 ( .B1(n17776), .B2(n17775), .A(n17774), .ZN(n17792) );
  OAI22_X1 U20887 ( .A1(n17800), .A2(n17778), .B1(n17777), .B2(n17792), .ZN(
        n17779) );
  AOI21_X1 U20888 ( .B1(n9848), .B2(n18093), .A(n17779), .ZN(n17780) );
  OAI211_X1 U20889 ( .C1(n18499), .C2(n17782), .A(n17781), .B(n17780), .ZN(
        P3_U2826) );
  AOI21_X1 U20890 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17817), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17793) );
  AOI21_X1 U20891 ( .B1(n17785), .B2(n17784), .A(n17783), .ZN(n18098) );
  AOI22_X1 U20892 ( .A1(n18126), .A2(P3_REIP_REG_3__SCAN_IN), .B1(n17806), 
        .B2(n18098), .ZN(n17791) );
  AOI21_X1 U20893 ( .B1(n17788), .B2(n17787), .A(n17786), .ZN(n18100) );
  AOI22_X1 U20894 ( .A1(n9848), .A2(n18100), .B1(n17789), .B2(n17808), .ZN(
        n17790) );
  OAI211_X1 U20895 ( .C1(n17793), .C2(n17792), .A(n17791), .B(n17790), .ZN(
        P3_U2827) );
  INV_X1 U20896 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17803) );
  AOI21_X1 U20897 ( .B1(n17796), .B2(n17795), .A(n17794), .ZN(n18112) );
  NOR2_X1 U20898 ( .A1(n18138), .A2(n21028), .ZN(n18118) );
  INV_X1 U20899 ( .A(n9848), .ZN(n17821) );
  XNOR2_X1 U20900 ( .A(n17798), .B(n17797), .ZN(n18117) );
  OAI22_X1 U20901 ( .A1(n17800), .A2(n17799), .B1(n17821), .B2(n18117), .ZN(
        n17801) );
  AOI211_X1 U20902 ( .C1(n17806), .C2(n18112), .A(n18118), .B(n17801), .ZN(
        n17802) );
  OAI221_X1 U20903 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18499), .C1(
        n17803), .C2(n17817), .A(n17802), .ZN(P3_U2828) );
  INV_X1 U20904 ( .A(n17804), .ZN(n17813) );
  OAI21_X1 U20905 ( .B1(n17814), .B2(n11774), .A(n17805), .ZN(n18124) );
  AOI22_X1 U20906 ( .A1(n18126), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n17806), 
        .B2(n18124), .ZN(n17811) );
  AOI21_X1 U20907 ( .B1(n17816), .B2(n11774), .A(n17807), .ZN(n18123) );
  AOI22_X1 U20908 ( .A1(n9848), .A2(n18123), .B1(n17812), .B2(n17808), .ZN(
        n17810) );
  OAI211_X1 U20909 ( .C1(n17813), .C2(n17812), .A(n17811), .B(n17810), .ZN(
        P3_U2829) );
  INV_X1 U20910 ( .A(n17814), .ZN(n17815) );
  NAND2_X1 U20911 ( .A1(n17816), .A2(n17815), .ZN(n18143) );
  INV_X1 U20912 ( .A(n18143), .ZN(n18145) );
  NAND3_X1 U20913 ( .A1(n18757), .A2(n17818), .A3(n17817), .ZN(n17819) );
  AOI22_X1 U20914 ( .A1(n18126), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17819), .ZN(n17820) );
  OAI221_X1 U20915 ( .B1(n18145), .B2(n17822), .C1(n18143), .C2(n17821), .A(
        n17820), .ZN(P3_U2830) );
  INV_X1 U20916 ( .A(n18113), .ZN(n18051) );
  OAI22_X1 U20917 ( .A1(n18615), .A2(n17885), .B1(n17871), .B2(n17940), .ZN(
        n17877) );
  OAI21_X1 U20918 ( .B1(n17886), .B2(n17920), .A(n18594), .ZN(n17823) );
  OAI21_X1 U20919 ( .B1(n18051), .B2(n17877), .A(n17823), .ZN(n17862) );
  AOI21_X1 U20920 ( .B1(n17824), .B2(n18113), .A(n17862), .ZN(n17847) );
  AOI22_X1 U20921 ( .A1(n18615), .A2(n17825), .B1(n17850), .B2(n18594), .ZN(
        n17830) );
  AOI22_X1 U20922 ( .A1(n9828), .A2(n17827), .B1(n17989), .B2(n17826), .ZN(
        n17829) );
  NAND4_X1 U20923 ( .A1(n17847), .A2(n17830), .A3(n17829), .A4(n17828), .ZN(
        n17839) );
  AOI211_X1 U20924 ( .C1(n17831), .C2(n18594), .A(n20889), .B(n17839), .ZN(
        n17837) );
  AOI21_X1 U20925 ( .B1(n18136), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n17832), .ZN(n17836) );
  AOI22_X1 U20926 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18130), .B1(
        n18024), .B2(n17833), .ZN(n17835) );
  OAI211_X1 U20927 ( .C1(n17837), .C2(n17836), .A(n17835), .B(n17834), .ZN(
        P3_U2835) );
  NOR2_X1 U20928 ( .A1(n17887), .A2(n17838), .ZN(n17840) );
  MUX2_X1 U20929 ( .A(n17840), .B(n17839), .S(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .Z(n17841) );
  AOI22_X1 U20930 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18130), .B1(
        n18136), .B2(n17841), .ZN(n17843) );
  OAI211_X1 U20931 ( .C1(n17844), .C2(n18045), .A(n17843), .B(n17842), .ZN(
        P3_U2836) );
  AOI21_X1 U20932 ( .B1(n18606), .B2(n17845), .A(n17850), .ZN(n17848) );
  AOI22_X1 U20933 ( .A1(n17848), .A2(n17847), .B1(n17850), .B2(n17846), .ZN(
        n17855) );
  OAI21_X1 U20934 ( .B1(n18121), .B2(n17850), .A(n17849), .ZN(n17854) );
  OAI22_X1 U20935 ( .A1(n18144), .A2(n17852), .B1(n18045), .B2(n17851), .ZN(
        n17853) );
  AOI211_X1 U20936 ( .C1(n18136), .C2(n17855), .A(n17854), .B(n17853), .ZN(
        n17856) );
  OAI21_X1 U20937 ( .B1(n17979), .B2(n17857), .A(n17856), .ZN(P3_U2837) );
  AOI22_X1 U20938 ( .A1(n18126), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n17919), 
        .B2(n17858), .ZN(n17869) );
  OAI22_X1 U20939 ( .A1(n17860), .A2(n18010), .B1(n17859), .B2(n18787), .ZN(
        n17861) );
  NOR3_X1 U20940 ( .A1(n18130), .A2(n17862), .A3(n17861), .ZN(n17866) );
  INV_X1 U20941 ( .A(n17866), .ZN(n17867) );
  AOI221_X1 U20942 ( .B1(n17871), .B2(n18606), .C1(n17864), .C2(n18606), .A(
        n17863), .ZN(n17865) );
  AOI21_X1 U20943 ( .B1(n17866), .B2(n17865), .A(n18140), .ZN(n17872) );
  OAI211_X1 U20944 ( .C1(n18091), .C2(n17867), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n17872), .ZN(n17868) );
  OAI211_X1 U20945 ( .C1(n17870), .C2(n18045), .A(n17869), .B(n17868), .ZN(
        P3_U2838) );
  NOR3_X1 U20946 ( .A1(n18130), .A2(n17887), .A3(n17871), .ZN(n17873) );
  OAI21_X1 U20947 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17873), .A(
        n17872), .ZN(n17874) );
  OAI211_X1 U20948 ( .C1(n17876), .C2(n18045), .A(n17875), .B(n17874), .ZN(
        P3_U2839) );
  AOI22_X1 U20949 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18130), .B1(
        n18140), .B2(P3_REIP_REG_22__SCAN_IN), .ZN(n17892) );
  INV_X1 U20950 ( .A(n17877), .ZN(n17890) );
  INV_X1 U20951 ( .A(n17990), .ZN(n18026) );
  AOI22_X1 U20952 ( .A1(n9828), .A2(n17878), .B1(n17989), .B2(n11609), .ZN(
        n17895) );
  NAND2_X1 U20953 ( .A1(n18787), .A2(n18010), .ZN(n18013) );
  AOI21_X1 U20954 ( .B1(n17923), .B2(n17879), .A(n18629), .ZN(n17925) );
  INV_X1 U20955 ( .A(n17920), .ZN(n17880) );
  AOI21_X1 U20956 ( .B1(n17880), .B2(n17906), .A(n18617), .ZN(n17881) );
  AOI211_X1 U20957 ( .C1(n18606), .C2(n17882), .A(n17925), .B(n17881), .ZN(
        n17904) );
  OAI21_X1 U20958 ( .B1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n18617), .A(
        n17904), .ZN(n17883) );
  AOI21_X1 U20959 ( .B1(n17886), .B2(n18013), .A(n17883), .ZN(n17897) );
  OAI211_X1 U20960 ( .C1(n17884), .C2(n18026), .A(n17895), .B(n17897), .ZN(
        n17889) );
  OAI21_X1 U20961 ( .B1(n17887), .B2(n17886), .A(n17885), .ZN(n17888) );
  OAI211_X1 U20962 ( .C1(n17890), .C2(n17889), .A(n18136), .B(n17888), .ZN(
        n17891) );
  OAI211_X1 U20963 ( .C1(n17893), .C2(n18045), .A(n17892), .B(n17891), .ZN(
        P3_U2840) );
  AOI22_X1 U20964 ( .A1(n18126), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18024), 
        .B2(n17894), .ZN(n17901) );
  NAND2_X1 U20965 ( .A1(n18136), .A2(n17895), .ZN(n17943) );
  AOI221_X1 U20966 ( .B1(n17896), .B2(n18615), .C1(n17940), .C2(n18615), .A(
        n17943), .ZN(n17905) );
  OAI211_X1 U20967 ( .C1(n18129), .C2(n17898), .A(n17905), .B(n17897), .ZN(
        n17899) );
  NAND3_X1 U20968 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18138), .A3(
        n17899), .ZN(n17900) );
  OAI211_X1 U20969 ( .C1(n17902), .C2(n17911), .A(n17901), .B(n17900), .ZN(
        P3_U2841) );
  AOI22_X1 U20970 ( .A1(n18126), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n18024), 
        .B2(n17903), .ZN(n17910) );
  INV_X1 U20971 ( .A(n18013), .ZN(n17922) );
  OAI211_X1 U20972 ( .C1(n17906), .C2(n17922), .A(n17905), .B(n17904), .ZN(
        n17907) );
  AND2_X1 U20973 ( .A1(n18138), .A2(n17907), .ZN(n17915) );
  NOR3_X1 U20974 ( .A1(n18129), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n18809), .ZN(n17908) );
  OAI21_X1 U20975 ( .B1(n17915), .B2(n17908), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17909) );
  OAI211_X1 U20976 ( .C1(n17912), .C2(n17911), .A(n17910), .B(n17909), .ZN(
        P3_U2842) );
  INV_X1 U20977 ( .A(n17913), .ZN(n17914) );
  AOI22_X1 U20978 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17915), .B1(
        n17919), .B2(n17914), .ZN(n17917) );
  OAI211_X1 U20979 ( .C1(n17918), .C2(n18045), .A(n17917), .B(n17916), .ZN(
        P3_U2843) );
  NOR2_X1 U20980 ( .A1(n18033), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18114) );
  NOR3_X1 U20981 ( .A1(n18114), .A2(n17920), .A3(n17947), .ZN(n17921) );
  OAI22_X1 U20982 ( .A1(n17923), .A2(n17922), .B1(n18051), .B2(n17921), .ZN(
        n17924) );
  NOR3_X1 U20983 ( .A1(n17925), .A2(n17943), .A3(n17924), .ZN(n17932) );
  AOI221_X1 U20984 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17932), 
        .C1(n18051), .C2(n17932), .A(n18126), .ZN(n17927) );
  AOI22_X1 U20985 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17927), .B1(
        n18024), .B2(n17926), .ZN(n17929) );
  NAND2_X1 U20986 ( .A1(n18126), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n17928) );
  OAI211_X1 U20987 ( .C1(n17930), .C2(n17911), .A(n17929), .B(n17928), .ZN(
        P3_U2844) );
  NOR2_X1 U20988 ( .A1(n18138), .A2(n18702), .ZN(n17934) );
  NOR3_X1 U20989 ( .A1(n18126), .A2(n17932), .A3(n17931), .ZN(n17933) );
  AOI211_X1 U20990 ( .C1(n18024), .C2(n17935), .A(n17934), .B(n17933), .ZN(
        n17936) );
  OAI21_X1 U20991 ( .B1(n17911), .B2(n17937), .A(n17936), .ZN(P3_U2845) );
  INV_X1 U20992 ( .A(n17951), .ZN(n17942) );
  NOR2_X1 U20993 ( .A1(n17938), .A2(n18629), .ZN(n18007) );
  NOR2_X1 U20994 ( .A1(n18617), .A2(n17939), .ZN(n18028) );
  NOR2_X1 U20995 ( .A1(n18007), .A2(n18028), .ZN(n17966) );
  OAI21_X1 U20996 ( .B1(n17950), .B2(n18615), .A(n17940), .ZN(n17941) );
  OAI211_X1 U20997 ( .C1(n17942), .C2(n18026), .A(n17966), .B(n17941), .ZN(
        n17958) );
  OAI221_X1 U20998 ( .B1(n17943), .B2(n18091), .C1(n17943), .C2(n17958), .A(
        n18138), .ZN(n17946) );
  AOI22_X1 U20999 ( .A1(n18126), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n18024), 
        .B2(n17944), .ZN(n17945) );
  OAI221_X1 U21000 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17911), 
        .C1(n17947), .C2(n17946), .A(n17945), .ZN(P3_U2846) );
  INV_X1 U21001 ( .A(n18053), .ZN(n18108) );
  INV_X1 U21002 ( .A(n18106), .ZN(n17948) );
  AOI22_X1 U21003 ( .A1(n18108), .A2(n18606), .B1(n17948), .B2(n18050), .ZN(
        n18105) );
  NOR2_X1 U21004 ( .A1(n17949), .A2(n18105), .ZN(n17981) );
  INV_X1 U21005 ( .A(n17981), .ZN(n17969) );
  OAI21_X1 U21006 ( .B1(n17951), .B2(n17969), .A(n17950), .ZN(n17959) );
  NOR2_X1 U21007 ( .A1(n17952), .A2(n18787), .ZN(n17956) );
  NOR2_X1 U21008 ( .A1(n17953), .A2(n18010), .ZN(n17954) );
  AOI222_X1 U21009 ( .A1(n17959), .A2(n17958), .B1(n17957), .B2(n17956), .C1(
        n17955), .C2(n17954), .ZN(n17963) );
  AOI22_X1 U21010 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18130), .B1(
        n18024), .B2(n17960), .ZN(n17962) );
  OAI211_X1 U21011 ( .C1(n17963), .C2(n18128), .A(n17962), .B(n17961), .ZN(
        P3_U2847) );
  OAI21_X1 U21012 ( .B1(n17965), .B2(n17964), .A(n18615), .ZN(n17985) );
  OAI211_X1 U21013 ( .C1(n18129), .C2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n17966), .B(n17985), .ZN(n17967) );
  AOI211_X1 U21014 ( .C1(n17970), .C2(n17990), .A(n17971), .B(n17967), .ZN(
        n17968) );
  AOI221_X1 U21015 ( .B1(n17970), .B2(n17971), .C1(n17969), .C2(n17971), .A(
        n17968), .ZN(n17976) );
  OAI22_X1 U21016 ( .A1(n17971), .A2(n18121), .B1(n18138), .B2(n18698), .ZN(
        n17975) );
  OAI22_X1 U21017 ( .A1(n18144), .A2(n17973), .B1(n18045), .B2(n17972), .ZN(
        n17974) );
  AOI211_X1 U21018 ( .C1(n18136), .C2(n17976), .A(n17975), .B(n17974), .ZN(
        n17977) );
  OAI21_X1 U21019 ( .B1(n17979), .B2(n17978), .A(n17977), .ZN(P3_U2848) );
  INV_X1 U21020 ( .A(n17980), .ZN(n17994) );
  OAI21_X1 U21021 ( .B1(n17982), .B2(n17981), .A(n18136), .ZN(n18020) );
  NOR2_X1 U21022 ( .A1(n17984), .A2(n18020), .ZN(n17998) );
  INV_X1 U21023 ( .A(n17983), .ZN(n17988) );
  AOI21_X1 U21024 ( .B1(n17984), .B2(n17990), .A(n18028), .ZN(n18015) );
  OAI211_X1 U21025 ( .C1(n17986), .C2(n18787), .A(n18015), .B(n17985), .ZN(
        n17987) );
  AOI21_X1 U21026 ( .B1(n17989), .B2(n17988), .A(n17987), .ZN(n17999) );
  AOI211_X1 U21027 ( .C1(n21186), .C2(n17990), .A(n18007), .B(n18128), .ZN(
        n17992) );
  AOI211_X1 U21028 ( .C1(n17999), .C2(n17992), .A(n18126), .B(n17991), .ZN(
        n17993) );
  AOI21_X1 U21029 ( .B1(n17994), .B2(n17998), .A(n17993), .ZN(n17996) );
  OAI211_X1 U21030 ( .C1(n17997), .C2(n18045), .A(n17996), .B(n17995), .ZN(
        P3_U2849) );
  AOI21_X1 U21031 ( .B1(n18136), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n17998), .ZN(n18005) );
  INV_X1 U21032 ( .A(n17999), .ZN(n18000) );
  NOR3_X1 U21033 ( .A1(n18007), .A2(n21186), .A3(n18000), .ZN(n18004) );
  AOI22_X1 U21034 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18130), .B1(
        n18024), .B2(n18001), .ZN(n18003) );
  OAI211_X1 U21035 ( .C1(n18005), .C2(n18004), .A(n18003), .B(n18002), .ZN(
        P3_U2850) );
  INV_X1 U21036 ( .A(n18020), .ZN(n18039) );
  AOI22_X1 U21037 ( .A1(n18126), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18039), 
        .B2(n18006), .ZN(n18018) );
  AOI21_X1 U21038 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18032), .A(
        n18033), .ZN(n18012) );
  AOI211_X1 U21039 ( .C1(n18008), .C2(n9828), .A(n18007), .B(n18128), .ZN(
        n18009) );
  OAI21_X1 U21040 ( .B1(n18011), .B2(n18010), .A(n18009), .ZN(n18034) );
  AOI211_X1 U21041 ( .C1(n18014), .C2(n18013), .A(n18012), .B(n18034), .ZN(
        n18025) );
  OAI211_X1 U21042 ( .C1(n18033), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18015), .B(n18025), .ZN(n18016) );
  NAND3_X1 U21043 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18138), .A3(
        n18016), .ZN(n18017) );
  OAI211_X1 U21044 ( .C1(n18019), .C2(n18045), .A(n18018), .B(n18017), .ZN(
        P3_U2851) );
  NOR3_X1 U21045 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18021), .A3(
        n18020), .ZN(n18022) );
  AOI21_X1 U21046 ( .B1(n18024), .B2(n18023), .A(n18022), .ZN(n18031) );
  OAI21_X1 U21047 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18026), .A(
        n18025), .ZN(n18027) );
  OAI211_X1 U21048 ( .C1(n18028), .C2(n18027), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n18138), .ZN(n18029) );
  NAND3_X1 U21049 ( .A1(n18031), .A2(n18030), .A3(n18029), .ZN(P3_U2852) );
  AOI221_X1 U21050 ( .B1(n18593), .B2(n18033), .C1(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n18033), .A(n18032), .ZN(
        n18035) );
  AOI211_X1 U21051 ( .C1(n18594), .C2(n18036), .A(n18035), .B(n18034), .ZN(
        n18037) );
  OAI21_X1 U21052 ( .B1(n18140), .B2(n18037), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18038) );
  OAI21_X1 U21053 ( .B1(n18039), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n18038), .ZN(n18041) );
  OAI211_X1 U21054 ( .C1(n18042), .C2(n18045), .A(n18041), .B(n18040), .ZN(
        P3_U2853) );
  INV_X1 U21055 ( .A(n18043), .ZN(n18048) );
  OAI22_X1 U21056 ( .A1(n18046), .A2(n18045), .B1(n18144), .B2(n18044), .ZN(
        n18047) );
  AOI21_X1 U21057 ( .B1(n18049), .B2(n18048), .A(n18047), .ZN(n18062) );
  INV_X1 U21058 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18083) );
  NOR2_X1 U21059 ( .A1(n18083), .A2(n18088), .ZN(n18054) );
  OAI21_X1 U21060 ( .B1(n18051), .B2(n18050), .A(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18052) );
  AOI211_X1 U21061 ( .C1(n18053), .C2(n18606), .A(n18114), .B(n18052), .ZN(
        n18099) );
  AOI21_X1 U21062 ( .B1(n18054), .B2(n18099), .A(n18055), .ZN(n18080) );
  OAI22_X1 U21063 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18128), .B1(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18055), .ZN(n18056) );
  NOR2_X1 U21064 ( .A1(n18080), .A2(n18056), .ZN(n18065) );
  NAND2_X1 U21065 ( .A1(n18065), .A2(n18121), .ZN(n18063) );
  OAI211_X1 U21066 ( .C1(n18130), .C2(n18091), .A(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n18063), .ZN(n18060) );
  INV_X1 U21067 ( .A(n18105), .ZN(n18082) );
  NAND4_X1 U21068 ( .A1(n18136), .A2(n18058), .A3(n18057), .A4(n18082), .ZN(
        n18059) );
  NAND4_X1 U21069 ( .A1(n18062), .A2(n18061), .A3(n18060), .A4(n18059), .ZN(
        P3_U2854) );
  INV_X1 U21070 ( .A(n18063), .ZN(n18072) );
  NOR4_X1 U21071 ( .A1(n18105), .A2(n18065), .A3(n18073), .A4(n18064), .ZN(
        n18068) );
  OAI22_X1 U21072 ( .A1(n18138), .A2(n18686), .B1(n18144), .B2(n18066), .ZN(
        n18067) );
  AOI211_X1 U21073 ( .C1(n18069), .C2(n18135), .A(n18068), .B(n18067), .ZN(
        n18070) );
  OAI21_X1 U21074 ( .B1(n18072), .B2(n18071), .A(n18070), .ZN(P3_U2855) );
  NOR2_X1 U21075 ( .A1(n18138), .A2(n20952), .ZN(n18075) );
  NOR4_X1 U21076 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18105), .A3(
        n18128), .A4(n18073), .ZN(n18074) );
  AOI211_X1 U21077 ( .C1(n18076), .C2(n18135), .A(n18075), .B(n18074), .ZN(
        n18078) );
  OAI21_X1 U21078 ( .B1(n18130), .B2(n18080), .A(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18077) );
  OAI211_X1 U21079 ( .C1(n18079), .C2(n18144), .A(n18078), .B(n18077), .ZN(
        P3_U2856) );
  NOR2_X1 U21080 ( .A1(n18130), .A2(n18080), .ZN(n18089) );
  AOI22_X1 U21081 ( .A1(n18126), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18135), 
        .B2(n18081), .ZN(n18087) );
  NAND3_X1 U21082 ( .A1(n18136), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n18082), .ZN(n18097) );
  NOR3_X1 U21083 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18083), .A3(
        n18097), .ZN(n18084) );
  AOI21_X1 U21084 ( .B1(n18085), .B2(n18125), .A(n18084), .ZN(n18086) );
  OAI211_X1 U21085 ( .C1(n18089), .C2(n18088), .A(n18087), .B(n18086), .ZN(
        P3_U2857) );
  AOI22_X1 U21086 ( .A1(n18126), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18125), 
        .B2(n18090), .ZN(n18096) );
  INV_X1 U21087 ( .A(n18091), .ZN(n18092) );
  OR2_X1 U21088 ( .A1(n18099), .A2(n18128), .ZN(n18104) );
  OAI21_X1 U21089 ( .B1(n18092), .B2(n18104), .A(n18121), .ZN(n18094) );
  AOI22_X1 U21090 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18094), .B1(
        n18135), .B2(n18093), .ZN(n18095) );
  OAI211_X1 U21091 ( .C1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n18097), .A(
        n18096), .B(n18095), .ZN(P3_U2858) );
  AOI22_X1 U21092 ( .A1(n18126), .A2(P3_REIP_REG_3__SCAN_IN), .B1(n18125), 
        .B2(n18098), .ZN(n18103) );
  OAI21_X1 U21093 ( .B1(n18099), .B2(n18128), .A(n18121), .ZN(n18101) );
  AOI22_X1 U21094 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18101), .B1(
        n18135), .B2(n18100), .ZN(n18102) );
  OAI211_X1 U21095 ( .C1(n18105), .C2(n18104), .A(n18103), .B(n18102), .ZN(
        P3_U2859) );
  NOR3_X1 U21096 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n21073), .A3(
        n18106), .ZN(n18110) );
  NAND2_X1 U21097 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18107) );
  AOI221_X1 U21098 ( .B1(n18122), .B2(n18108), .C1(n18107), .C2(n18108), .A(
        n18629), .ZN(n18109) );
  AOI211_X1 U21099 ( .C1(n18112), .C2(n9828), .A(n18110), .B(n18109), .ZN(
        n18116) );
  OAI211_X1 U21100 ( .C1(n18114), .C2(n21073), .A(n18113), .B(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18115) );
  OAI211_X1 U21101 ( .C1(n18117), .C2(n18785), .A(n18116), .B(n18115), .ZN(
        n18119) );
  AOI21_X1 U21102 ( .B1(n18136), .B2(n18119), .A(n18118), .ZN(n18120) );
  OAI21_X1 U21103 ( .B1(n18122), .B2(n18121), .A(n18120), .ZN(P3_U2860) );
  AOI22_X1 U21104 ( .A1(n18125), .A2(n18124), .B1(n18135), .B2(n18123), .ZN(
        n18134) );
  NAND2_X1 U21105 ( .A1(n18126), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18133) );
  OAI211_X1 U21106 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n18594), .A(
        n18127), .B(n21073), .ZN(n18132) );
  NOR3_X1 U21107 ( .A1(n18129), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n18128), .ZN(n18137) );
  OAI21_X1 U21108 ( .B1(n18130), .B2(n18137), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18131) );
  NAND4_X1 U21109 ( .A1(n18134), .A2(n18133), .A3(n18132), .A4(n18131), .ZN(
        P3_U2861) );
  INV_X1 U21110 ( .A(n18135), .ZN(n18142) );
  INV_X1 U21111 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21053) );
  AOI21_X1 U21112 ( .B1(n18136), .B2(n18617), .A(n21053), .ZN(n18139) );
  AOI221_X1 U21113 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(n18140), .C1(n18139), 
        .C2(n18138), .A(n18137), .ZN(n18141) );
  OAI221_X1 U21114 ( .B1(n18145), .B2(n18144), .C1(n18143), .C2(n18142), .A(
        n18141), .ZN(P3_U2862) );
  AOI21_X1 U21115 ( .B1(n18148), .B2(n18147), .A(n18146), .ZN(n18646) );
  OAI21_X1 U21116 ( .B1(n18646), .B2(n18192), .A(n18153), .ZN(n18149) );
  OAI221_X1 U21117 ( .B1(n18392), .B2(n18801), .C1(n18392), .C2(n18153), .A(
        n18149), .ZN(P3_U2863) );
  NOR2_X1 U21118 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n21022), .ZN(
        n18371) );
  NOR2_X1 U21119 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18626), .ZN(
        n18325) );
  NOR2_X1 U21120 ( .A1(n18371), .A2(n18325), .ZN(n18151) );
  OAI22_X1 U21121 ( .A1(n18152), .A2(n21022), .B1(n18151), .B2(n18150), .ZN(
        P3_U2866) );
  NOR2_X1 U21122 ( .A1(n18154), .A2(n18153), .ZN(P3_U2867) );
  NOR2_X1 U21123 ( .A1(n18626), .A2(n21022), .ZN(n18469) );
  NOR2_X1 U21124 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18392), .ZN(
        n18370) );
  NAND2_X1 U21125 ( .A1(n18469), .A2(n18370), .ZN(n18575) );
  NAND2_X1 U21126 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18471), .ZN(n18537) );
  NOR2_X1 U21127 ( .A1(n21022), .A2(n18300), .ZN(n18532) );
  NAND2_X1 U21128 ( .A1(n18392), .A2(n18532), .ZN(n18498) );
  INV_X1 U21129 ( .A(n18498), .ZN(n18523) );
  NOR2_X2 U21130 ( .A1(n18499), .A2(n14135), .ZN(n18530) );
  NOR2_X2 U21131 ( .A1(n18441), .A2(n18155), .ZN(n18529) );
  NAND2_X1 U21132 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18621) );
  INV_X1 U21133 ( .A(n18469), .ZN(n18466) );
  NOR2_X2 U21134 ( .A1(n18621), .A2(n18466), .ZN(n18581) );
  NAND2_X1 U21135 ( .A1(n20915), .A2(n18392), .ZN(n18622) );
  NAND2_X1 U21136 ( .A1(n18626), .A2(n21022), .ZN(n18233) );
  NOR2_X1 U21137 ( .A1(n18622), .A2(n18233), .ZN(n18244) );
  CLKBUF_X1 U21138 ( .A(n18244), .Z(n18253) );
  NOR2_X1 U21139 ( .A1(n18581), .A2(n18253), .ZN(n18212) );
  NOR2_X1 U21140 ( .A1(n18654), .A2(n18212), .ZN(n18186) );
  AOI22_X1 U21141 ( .A1(n18523), .A2(n18530), .B1(n18529), .B2(n18186), .ZN(
        n18162) );
  AOI21_X1 U21142 ( .B1(n18575), .B2(n18498), .A(n18441), .ZN(n18502) );
  AOI211_X1 U21143 ( .C1(P3_STATE2_REG_3__SCAN_IN), .C2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n18212), .B(n18441), .ZN(
        n18156) );
  AOI21_X1 U21144 ( .B1(n18502), .B2(n18211), .A(n18156), .ZN(n18189) );
  INV_X1 U21145 ( .A(n18157), .ZN(n18158) );
  NAND2_X1 U21146 ( .A1(n18159), .A2(n18158), .ZN(n18187) );
  NOR2_X1 U21147 ( .A1(n18160), .A2(n18187), .ZN(n18534) );
  AOI22_X1 U21148 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18189), .B1(
        n18253), .B2(n18534), .ZN(n18161) );
  OAI211_X1 U21149 ( .C1(n18575), .C2(n18537), .A(n18162), .B(n18161), .ZN(
        P3_U2868) );
  NAND2_X1 U21150 ( .A1(n18471), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18543) );
  INV_X1 U21151 ( .A(n18575), .ZN(n18579) );
  NAND2_X1 U21152 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18471), .ZN(n18448) );
  INV_X1 U21153 ( .A(n18448), .ZN(n18539) );
  AND2_X1 U21154 ( .A1(n18393), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18538) );
  AOI22_X1 U21155 ( .A1(n18579), .A2(n18539), .B1(n18186), .B2(n18538), .ZN(
        n18165) );
  NOR2_X2 U21156 ( .A1(n18163), .A2(n18187), .ZN(n18540) );
  AOI22_X1 U21157 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18189), .B1(
        n18253), .B2(n18540), .ZN(n18164) );
  OAI211_X1 U21158 ( .C1(n18498), .C2(n18543), .A(n18165), .B(n18164), .ZN(
        P3_U2869) );
  NAND2_X1 U21159 ( .A1(n18471), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18549) );
  NAND2_X1 U21160 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18471), .ZN(n18510) );
  INV_X1 U21161 ( .A(n18510), .ZN(n18545) );
  NOR2_X2 U21162 ( .A1(n18441), .A2(n18166), .ZN(n18544) );
  AOI22_X1 U21163 ( .A1(n18579), .A2(n18545), .B1(n18186), .B2(n18544), .ZN(
        n18169) );
  NOR2_X2 U21164 ( .A1(n18167), .A2(n18187), .ZN(n18546) );
  AOI22_X1 U21165 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18189), .B1(
        n18244), .B2(n18546), .ZN(n18168) );
  OAI211_X1 U21166 ( .C1(n18498), .C2(n18549), .A(n18169), .B(n18168), .ZN(
        P3_U2870) );
  NAND2_X1 U21167 ( .A1(n18471), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18555) );
  NOR2_X1 U21168 ( .A1(n19178), .A2(n18499), .ZN(n18550) );
  NOR2_X2 U21169 ( .A1(n18441), .A2(n18170), .ZN(n18551) );
  AOI22_X1 U21170 ( .A1(n18579), .A2(n18550), .B1(n18186), .B2(n18551), .ZN(
        n18173) );
  NOR2_X2 U21171 ( .A1(n18171), .A2(n18187), .ZN(n18552) );
  AOI22_X1 U21172 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18189), .B1(
        n18244), .B2(n18552), .ZN(n18172) );
  OAI211_X1 U21173 ( .C1(n18498), .C2(n18555), .A(n18173), .B(n18172), .ZN(
        P3_U2871) );
  NAND2_X1 U21174 ( .A1(n18471), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18561) );
  NOR2_X1 U21175 ( .A1(n21025), .A2(n18499), .ZN(n18556) );
  NOR2_X2 U21176 ( .A1(n18441), .A2(n18174), .ZN(n18557) );
  AOI22_X1 U21177 ( .A1(n18579), .A2(n18556), .B1(n18186), .B2(n18557), .ZN(
        n18177) );
  NOR2_X2 U21178 ( .A1(n18175), .A2(n18187), .ZN(n18558) );
  AOI22_X1 U21179 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18189), .B1(
        n18253), .B2(n18558), .ZN(n18176) );
  OAI211_X1 U21180 ( .C1(n18498), .C2(n18561), .A(n18177), .B(n18176), .ZN(
        P3_U2872) );
  NAND2_X1 U21181 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18471), .ZN(n18567) );
  NOR2_X2 U21182 ( .A1(n18499), .A2(n15309), .ZN(n18563) );
  NOR2_X2 U21183 ( .A1(n18441), .A2(n21103), .ZN(n18562) );
  AOI22_X1 U21184 ( .A1(n18523), .A2(n18563), .B1(n18186), .B2(n18562), .ZN(
        n18180) );
  NOR2_X1 U21185 ( .A1(n18178), .A2(n18187), .ZN(n18564) );
  AOI22_X1 U21186 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18189), .B1(
        n18253), .B2(n18564), .ZN(n18179) );
  OAI211_X1 U21187 ( .C1(n18575), .C2(n18567), .A(n18180), .B(n18179), .ZN(
        P3_U2873) );
  NAND2_X1 U21188 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18471), .ZN(n18493) );
  NOR2_X1 U21189 ( .A1(n18499), .A2(n15303), .ZN(n18490) );
  NOR2_X2 U21190 ( .A1(n18441), .A2(n18181), .ZN(n18568) );
  AOI22_X1 U21191 ( .A1(n18523), .A2(n18490), .B1(n18186), .B2(n18568), .ZN(
        n18184) );
  NOR2_X2 U21192 ( .A1(n18182), .A2(n18187), .ZN(n18571) );
  AOI22_X1 U21193 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18189), .B1(
        n18244), .B2(n18571), .ZN(n18183) );
  OAI211_X1 U21194 ( .C1(n18575), .C2(n18493), .A(n18184), .B(n18183), .ZN(
        P3_U2874) );
  NAND2_X1 U21195 ( .A1(n18471), .A2(BUF2_REG_23__SCAN_IN), .ZN(n18369) );
  NOR2_X1 U21196 ( .A1(n18499), .A2(n20974), .ZN(n18364) );
  NOR2_X2 U21197 ( .A1(n18441), .A2(n18185), .ZN(n18577) );
  AOI22_X1 U21198 ( .A1(n18579), .A2(n18364), .B1(n18186), .B2(n18577), .ZN(
        n18191) );
  NOR2_X2 U21199 ( .A1(n18188), .A2(n18187), .ZN(n18580) );
  AOI22_X1 U21200 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18189), .B1(
        n18253), .B2(n18580), .ZN(n18190) );
  OAI211_X1 U21201 ( .C1(n18498), .C2(n18369), .A(n18191), .B(n18190), .ZN(
        P3_U2875) );
  INV_X1 U21202 ( .A(n18233), .ZN(n18235) );
  NAND2_X1 U21203 ( .A1(n18370), .A2(n18235), .ZN(n18278) );
  INV_X1 U21204 ( .A(n18537), .ZN(n18467) );
  INV_X1 U21205 ( .A(n18654), .ZN(n18528) );
  NAND2_X1 U21206 ( .A1(n20915), .A2(n18528), .ZN(n18465) );
  NOR2_X1 U21207 ( .A1(n18233), .A2(n18465), .ZN(n18207) );
  AOI22_X1 U21208 ( .A1(n18467), .A2(n18523), .B1(n18529), .B2(n18207), .ZN(
        n18194) );
  NOR2_X1 U21209 ( .A1(n18441), .A2(n18192), .ZN(n18531) );
  INV_X1 U21210 ( .A(n18531), .ZN(n18234) );
  NOR2_X1 U21211 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18234), .ZN(
        n18468) );
  AOI22_X1 U21212 ( .A1(n18471), .A2(n18532), .B1(n18235), .B2(n18468), .ZN(
        n18208) );
  AOI22_X1 U21213 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18208), .B1(
        n18581), .B2(n18530), .ZN(n18193) );
  OAI211_X1 U21214 ( .C1(n18474), .C2(n18278), .A(n18194), .B(n18193), .ZN(
        P3_U2876) );
  INV_X1 U21215 ( .A(n18581), .ZN(n18228) );
  AOI22_X1 U21216 ( .A1(n18523), .A2(n18539), .B1(n18538), .B2(n18207), .ZN(
        n18196) );
  INV_X1 U21217 ( .A(n18278), .ZN(n18271) );
  AOI22_X1 U21218 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18208), .B1(
        n18540), .B2(n18271), .ZN(n18195) );
  OAI211_X1 U21219 ( .C1(n18228), .C2(n18543), .A(n18196), .B(n18195), .ZN(
        P3_U2877) );
  AOI22_X1 U21220 ( .A1(n18523), .A2(n18545), .B1(n18544), .B2(n18207), .ZN(
        n18198) );
  AOI22_X1 U21221 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18208), .B1(
        n18546), .B2(n18271), .ZN(n18197) );
  OAI211_X1 U21222 ( .C1(n18228), .C2(n18549), .A(n18198), .B(n18197), .ZN(
        P3_U2878) );
  AOI22_X1 U21223 ( .A1(n18523), .A2(n18550), .B1(n18551), .B2(n18207), .ZN(
        n18200) );
  AOI22_X1 U21224 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18208), .B1(
        n18552), .B2(n18271), .ZN(n18199) );
  OAI211_X1 U21225 ( .C1(n18228), .C2(n18555), .A(n18200), .B(n18199), .ZN(
        P3_U2879) );
  AOI22_X1 U21226 ( .A1(n18523), .A2(n18556), .B1(n18557), .B2(n18207), .ZN(
        n18202) );
  AOI22_X1 U21227 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18208), .B1(
        n18558), .B2(n18271), .ZN(n18201) );
  OAI211_X1 U21228 ( .C1(n18228), .C2(n18561), .A(n18202), .B(n18201), .ZN(
        P3_U2880) );
  AOI22_X1 U21229 ( .A1(n18581), .A2(n18563), .B1(n18562), .B2(n18207), .ZN(
        n18204) );
  AOI22_X1 U21230 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18208), .B1(
        n18564), .B2(n18271), .ZN(n18203) );
  OAI211_X1 U21231 ( .C1(n18498), .C2(n18567), .A(n18204), .B(n18203), .ZN(
        P3_U2881) );
  AOI22_X1 U21232 ( .A1(n18581), .A2(n18490), .B1(n18568), .B2(n18207), .ZN(
        n18206) );
  AOI22_X1 U21233 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18208), .B1(
        n18571), .B2(n18271), .ZN(n18205) );
  OAI211_X1 U21234 ( .C1(n18498), .C2(n18493), .A(n18206), .B(n18205), .ZN(
        P3_U2882) );
  AOI22_X1 U21235 ( .A1(n18523), .A2(n18364), .B1(n18577), .B2(n18207), .ZN(
        n18210) );
  AOI22_X1 U21236 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18208), .B1(
        n18580), .B2(n18271), .ZN(n18209) );
  OAI211_X1 U21237 ( .C1(n18228), .C2(n18369), .A(n18210), .B(n18209), .ZN(
        P3_U2883) );
  NOR2_X1 U21238 ( .A1(n20915), .A2(n18233), .ZN(n18279) );
  NAND2_X1 U21239 ( .A1(n18392), .A2(n18279), .ZN(n18299) );
  INV_X1 U21240 ( .A(n18211), .ZN(n18440) );
  NOR2_X1 U21241 ( .A1(n18271), .A2(n18290), .ZN(n18257) );
  OAI21_X1 U21242 ( .B1(n18212), .B2(n18440), .A(n18257), .ZN(n18213) );
  OAI211_X1 U21243 ( .C1(n18290), .C2(n18748), .A(n18393), .B(n18213), .ZN(
        n18230) );
  NOR2_X1 U21244 ( .A1(n18654), .A2(n18257), .ZN(n18229) );
  AOI22_X1 U21245 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18230), .B1(
        n18529), .B2(n18229), .ZN(n18215) );
  AOI22_X1 U21246 ( .A1(n18244), .A2(n18530), .B1(n18534), .B2(n18290), .ZN(
        n18214) );
  OAI211_X1 U21247 ( .C1(n18537), .C2(n18228), .A(n18215), .B(n18214), .ZN(
        P3_U2884) );
  INV_X1 U21248 ( .A(n18543), .ZN(n18445) );
  AOI22_X1 U21249 ( .A1(n18253), .A2(n18445), .B1(n18538), .B2(n18229), .ZN(
        n18217) );
  AOI22_X1 U21250 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18230), .B1(
        n18540), .B2(n18290), .ZN(n18216) );
  OAI211_X1 U21251 ( .C1(n18228), .C2(n18448), .A(n18217), .B(n18216), .ZN(
        P3_U2885) );
  INV_X1 U21252 ( .A(n18549), .ZN(n18507) );
  AOI22_X1 U21253 ( .A1(n18253), .A2(n18507), .B1(n18544), .B2(n18229), .ZN(
        n18219) );
  AOI22_X1 U21254 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18230), .B1(
        n18546), .B2(n18290), .ZN(n18218) );
  OAI211_X1 U21255 ( .C1(n18228), .C2(n18510), .A(n18219), .B(n18218), .ZN(
        P3_U2886) );
  INV_X1 U21256 ( .A(n18550), .ZN(n18514) );
  INV_X1 U21257 ( .A(n18555), .ZN(n18511) );
  AOI22_X1 U21258 ( .A1(n18244), .A2(n18511), .B1(n18551), .B2(n18229), .ZN(
        n18221) );
  AOI22_X1 U21259 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18230), .B1(
        n18552), .B2(n18290), .ZN(n18220) );
  OAI211_X1 U21260 ( .C1(n18228), .C2(n18514), .A(n18221), .B(n18220), .ZN(
        P3_U2887) );
  INV_X1 U21261 ( .A(n18556), .ZN(n18484) );
  INV_X1 U21262 ( .A(n18561), .ZN(n18481) );
  AOI22_X1 U21263 ( .A1(n18244), .A2(n18481), .B1(n18557), .B2(n18229), .ZN(
        n18223) );
  AOI22_X1 U21264 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18230), .B1(
        n18558), .B2(n18290), .ZN(n18222) );
  OAI211_X1 U21265 ( .C1(n18228), .C2(n18484), .A(n18223), .B(n18222), .ZN(
        P3_U2888) );
  INV_X1 U21266 ( .A(n18564), .ZN(n18489) );
  INV_X1 U21267 ( .A(n18567), .ZN(n18486) );
  AOI22_X1 U21268 ( .A1(n18581), .A2(n18486), .B1(n18562), .B2(n18229), .ZN(
        n18225) );
  AOI22_X1 U21269 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18230), .B1(
        n18253), .B2(n18563), .ZN(n18224) );
  OAI211_X1 U21270 ( .C1(n18489), .C2(n18299), .A(n18225), .B(n18224), .ZN(
        P3_U2889) );
  AOI22_X1 U21271 ( .A1(n18253), .A2(n18490), .B1(n18568), .B2(n18229), .ZN(
        n18227) );
  AOI22_X1 U21272 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18230), .B1(
        n18571), .B2(n18290), .ZN(n18226) );
  OAI211_X1 U21273 ( .C1(n18228), .C2(n18493), .A(n18227), .B(n18226), .ZN(
        P3_U2890) );
  INV_X1 U21274 ( .A(n18244), .ZN(n18251) );
  AOI22_X1 U21275 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18230), .B1(
        n18577), .B2(n18229), .ZN(n18232) );
  AOI22_X1 U21276 ( .A1(n18581), .A2(n18364), .B1(n18580), .B2(n18290), .ZN(
        n18231) );
  OAI211_X1 U21277 ( .C1(n18251), .C2(n18369), .A(n18232), .B(n18231), .ZN(
        P3_U2891) );
  NOR2_X2 U21278 ( .A1(n18621), .A2(n18233), .ZN(n18315) );
  INV_X1 U21279 ( .A(n18315), .ZN(n18322) );
  AND2_X1 U21280 ( .A1(n18528), .A2(n18279), .ZN(n18252) );
  AOI22_X1 U21281 ( .A1(n18467), .A2(n18244), .B1(n18529), .B2(n18252), .ZN(
        n18237) );
  AOI21_X1 U21282 ( .B1(n20915), .B2(n18440), .A(n18234), .ZN(n18324) );
  NAND2_X1 U21283 ( .A1(n18235), .A2(n18324), .ZN(n18254) );
  AOI22_X1 U21284 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18254), .B1(
        n18530), .B2(n18271), .ZN(n18236) );
  OAI211_X1 U21285 ( .C1(n18474), .C2(n18322), .A(n18237), .B(n18236), .ZN(
        P3_U2892) );
  AOI22_X1 U21286 ( .A1(n18253), .A2(n18539), .B1(n18538), .B2(n18252), .ZN(
        n18239) );
  AOI22_X1 U21287 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18254), .B1(
        n18540), .B2(n18315), .ZN(n18238) );
  OAI211_X1 U21288 ( .C1(n18543), .C2(n18278), .A(n18239), .B(n18238), .ZN(
        P3_U2893) );
  AOI22_X1 U21289 ( .A1(n18244), .A2(n18545), .B1(n18544), .B2(n18252), .ZN(
        n18241) );
  AOI22_X1 U21290 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18254), .B1(
        n18546), .B2(n18315), .ZN(n18240) );
  OAI211_X1 U21291 ( .C1(n18549), .C2(n18278), .A(n18241), .B(n18240), .ZN(
        P3_U2894) );
  AOI22_X1 U21292 ( .A1(n18511), .A2(n18271), .B1(n18551), .B2(n18252), .ZN(
        n18243) );
  AOI22_X1 U21293 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18254), .B1(
        n18552), .B2(n18315), .ZN(n18242) );
  OAI211_X1 U21294 ( .C1(n18251), .C2(n18514), .A(n18243), .B(n18242), .ZN(
        P3_U2895) );
  AOI22_X1 U21295 ( .A1(n18244), .A2(n18556), .B1(n18557), .B2(n18252), .ZN(
        n18246) );
  AOI22_X1 U21296 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18254), .B1(
        n18558), .B2(n18315), .ZN(n18245) );
  OAI211_X1 U21297 ( .C1(n18561), .C2(n18278), .A(n18246), .B(n18245), .ZN(
        P3_U2896) );
  AOI22_X1 U21298 ( .A1(n18562), .A2(n18252), .B1(n18563), .B2(n18271), .ZN(
        n18248) );
  AOI22_X1 U21299 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18254), .B1(
        n18564), .B2(n18315), .ZN(n18247) );
  OAI211_X1 U21300 ( .C1(n18251), .C2(n18567), .A(n18248), .B(n18247), .ZN(
        P3_U2897) );
  AOI22_X1 U21301 ( .A1(n18490), .A2(n18271), .B1(n18568), .B2(n18252), .ZN(
        n18250) );
  AOI22_X1 U21302 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18254), .B1(
        n18571), .B2(n18315), .ZN(n18249) );
  OAI211_X1 U21303 ( .C1(n18251), .C2(n18493), .A(n18250), .B(n18249), .ZN(
        P3_U2898) );
  AOI22_X1 U21304 ( .A1(n18253), .A2(n18364), .B1(n18577), .B2(n18252), .ZN(
        n18256) );
  AOI22_X1 U21305 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18254), .B1(
        n18580), .B2(n18315), .ZN(n18255) );
  OAI211_X1 U21306 ( .C1(n18369), .C2(n18278), .A(n18256), .B(n18255), .ZN(
        P3_U2899) );
  INV_X1 U21307 ( .A(n18622), .ZN(n18438) );
  NAND2_X1 U21308 ( .A1(n18438), .A2(n18325), .ZN(n18340) );
  AOI21_X1 U21309 ( .B1(n18322), .B2(n18340), .A(n18654), .ZN(n18274) );
  AOI22_X1 U21310 ( .A1(n18467), .A2(n18271), .B1(n18529), .B2(n18274), .ZN(
        n18260) );
  INV_X1 U21311 ( .A(n18340), .ZN(n18341) );
  OAI21_X1 U21312 ( .B1(n18315), .B2(n18341), .A(n18393), .ZN(n18301) );
  OAI21_X1 U21313 ( .B1(n18257), .B2(n18499), .A(n18301), .ZN(n18258) );
  OAI21_X1 U21314 ( .B1(n18341), .B2(n18748), .A(n18258), .ZN(n18275) );
  AOI22_X1 U21315 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18275), .B1(
        n18530), .B2(n18290), .ZN(n18259) );
  OAI211_X1 U21316 ( .C1(n18474), .C2(n18340), .A(n18260), .B(n18259), .ZN(
        P3_U2900) );
  AOI22_X1 U21317 ( .A1(n18445), .A2(n18290), .B1(n18538), .B2(n18274), .ZN(
        n18262) );
  AOI22_X1 U21318 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18275), .B1(
        n18540), .B2(n18341), .ZN(n18261) );
  OAI211_X1 U21319 ( .C1(n18448), .C2(n18278), .A(n18262), .B(n18261), .ZN(
        P3_U2901) );
  AOI22_X1 U21320 ( .A1(n18507), .A2(n18290), .B1(n18544), .B2(n18274), .ZN(
        n18264) );
  AOI22_X1 U21321 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18275), .B1(
        n18546), .B2(n18341), .ZN(n18263) );
  OAI211_X1 U21322 ( .C1(n18510), .C2(n18278), .A(n18264), .B(n18263), .ZN(
        P3_U2902) );
  AOI22_X1 U21323 ( .A1(n18551), .A2(n18274), .B1(n18550), .B2(n18271), .ZN(
        n18266) );
  AOI22_X1 U21324 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18275), .B1(
        n18552), .B2(n18341), .ZN(n18265) );
  OAI211_X1 U21325 ( .C1(n18555), .C2(n18299), .A(n18266), .B(n18265), .ZN(
        P3_U2903) );
  AOI22_X1 U21326 ( .A1(n18557), .A2(n18274), .B1(n18556), .B2(n18271), .ZN(
        n18268) );
  AOI22_X1 U21327 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18275), .B1(
        n18558), .B2(n18341), .ZN(n18267) );
  OAI211_X1 U21328 ( .C1(n18561), .C2(n18299), .A(n18268), .B(n18267), .ZN(
        P3_U2904) );
  AOI22_X1 U21329 ( .A1(n18486), .A2(n18271), .B1(n18562), .B2(n18274), .ZN(
        n18270) );
  AOI22_X1 U21330 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18275), .B1(
        n18563), .B2(n18290), .ZN(n18269) );
  OAI211_X1 U21331 ( .C1(n18489), .C2(n18340), .A(n18270), .B(n18269), .ZN(
        P3_U2905) );
  INV_X1 U21332 ( .A(n18490), .ZN(n18574) );
  INV_X1 U21333 ( .A(n18493), .ZN(n18570) );
  AOI22_X1 U21334 ( .A1(n18570), .A2(n18271), .B1(n18568), .B2(n18274), .ZN(
        n18273) );
  AOI22_X1 U21335 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18275), .B1(
        n18571), .B2(n18341), .ZN(n18272) );
  OAI211_X1 U21336 ( .C1(n18574), .C2(n18299), .A(n18273), .B(n18272), .ZN(
        P3_U2906) );
  INV_X1 U21337 ( .A(n18364), .ZN(n18586) );
  INV_X1 U21338 ( .A(n18369), .ZN(n18578) );
  AOI22_X1 U21339 ( .A1(n18578), .A2(n18290), .B1(n18577), .B2(n18274), .ZN(
        n18277) );
  AOI22_X1 U21340 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18275), .B1(
        n18580), .B2(n18341), .ZN(n18276) );
  OAI211_X1 U21341 ( .C1(n18586), .C2(n18278), .A(n18277), .B(n18276), .ZN(
        P3_U2907) );
  NAND2_X1 U21342 ( .A1(n18325), .A2(n18370), .ZN(n18362) );
  INV_X1 U21343 ( .A(n18325), .ZN(n18323) );
  NOR2_X1 U21344 ( .A1(n18323), .A2(n18465), .ZN(n18295) );
  AOI22_X1 U21345 ( .A1(n18467), .A2(n18290), .B1(n18529), .B2(n18295), .ZN(
        n18281) );
  AOI22_X1 U21346 ( .A1(n18471), .A2(n18279), .B1(n18325), .B2(n18468), .ZN(
        n18296) );
  AOI22_X1 U21347 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18296), .B1(
        n18530), .B2(n18315), .ZN(n18280) );
  OAI211_X1 U21348 ( .C1(n18474), .C2(n18362), .A(n18281), .B(n18280), .ZN(
        P3_U2908) );
  AOI22_X1 U21349 ( .A1(n18445), .A2(n18315), .B1(n18538), .B2(n18295), .ZN(
        n18283) );
  INV_X1 U21350 ( .A(n18362), .ZN(n18363) );
  AOI22_X1 U21351 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18296), .B1(
        n18540), .B2(n18363), .ZN(n18282) );
  OAI211_X1 U21352 ( .C1(n18448), .C2(n18299), .A(n18283), .B(n18282), .ZN(
        P3_U2909) );
  AOI22_X1 U21353 ( .A1(n18507), .A2(n18315), .B1(n18544), .B2(n18295), .ZN(
        n18285) );
  AOI22_X1 U21354 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18296), .B1(
        n18546), .B2(n18363), .ZN(n18284) );
  OAI211_X1 U21355 ( .C1(n18510), .C2(n18299), .A(n18285), .B(n18284), .ZN(
        P3_U2910) );
  AOI22_X1 U21356 ( .A1(n18551), .A2(n18295), .B1(n18550), .B2(n18290), .ZN(
        n18287) );
  AOI22_X1 U21357 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18296), .B1(
        n18552), .B2(n18363), .ZN(n18286) );
  OAI211_X1 U21358 ( .C1(n18555), .C2(n18322), .A(n18287), .B(n18286), .ZN(
        P3_U2911) );
  AOI22_X1 U21359 ( .A1(n18557), .A2(n18295), .B1(n18556), .B2(n18290), .ZN(
        n18289) );
  AOI22_X1 U21360 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18296), .B1(
        n18558), .B2(n18363), .ZN(n18288) );
  OAI211_X1 U21361 ( .C1(n18561), .C2(n18322), .A(n18289), .B(n18288), .ZN(
        P3_U2912) );
  AOI22_X1 U21362 ( .A1(n18486), .A2(n18290), .B1(n18562), .B2(n18295), .ZN(
        n18292) );
  AOI22_X1 U21363 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18296), .B1(
        n18563), .B2(n18315), .ZN(n18291) );
  OAI211_X1 U21364 ( .C1(n18489), .C2(n18362), .A(n18292), .B(n18291), .ZN(
        P3_U2913) );
  AOI22_X1 U21365 ( .A1(n18490), .A2(n18315), .B1(n18568), .B2(n18295), .ZN(
        n18294) );
  AOI22_X1 U21366 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18296), .B1(
        n18571), .B2(n18363), .ZN(n18293) );
  OAI211_X1 U21367 ( .C1(n18493), .C2(n18299), .A(n18294), .B(n18293), .ZN(
        P3_U2914) );
  AOI22_X1 U21368 ( .A1(n18578), .A2(n18315), .B1(n18577), .B2(n18295), .ZN(
        n18298) );
  AOI22_X1 U21369 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18296), .B1(
        n18580), .B2(n18363), .ZN(n18297) );
  OAI211_X1 U21370 ( .C1(n18586), .C2(n18299), .A(n18298), .B(n18297), .ZN(
        P3_U2915) );
  NOR2_X1 U21371 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18300), .ZN(
        n18372) );
  NAND2_X1 U21372 ( .A1(n18372), .A2(n18392), .ZN(n18391) );
  INV_X1 U21373 ( .A(n18391), .ZN(n18385) );
  NOR2_X1 U21374 ( .A1(n18363), .A2(n18385), .ZN(n18346) );
  NOR2_X1 U21375 ( .A1(n18654), .A2(n18346), .ZN(n18318) );
  AOI22_X1 U21376 ( .A1(n18467), .A2(n18315), .B1(n18529), .B2(n18318), .ZN(
        n18304) );
  OAI22_X1 U21377 ( .A1(n18346), .A2(n18441), .B1(n18440), .B2(n18301), .ZN(
        n18302) );
  OAI21_X1 U21378 ( .B1(n18385), .B2(n18748), .A(n18302), .ZN(n18319) );
  AOI22_X1 U21379 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18319), .B1(
        n18530), .B2(n18341), .ZN(n18303) );
  OAI211_X1 U21380 ( .C1(n18474), .C2(n18391), .A(n18304), .B(n18303), .ZN(
        P3_U2916) );
  AOI22_X1 U21381 ( .A1(n18539), .A2(n18315), .B1(n18538), .B2(n18318), .ZN(
        n18306) );
  AOI22_X1 U21382 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18319), .B1(
        n18540), .B2(n18385), .ZN(n18305) );
  OAI211_X1 U21383 ( .C1(n18543), .C2(n18340), .A(n18306), .B(n18305), .ZN(
        P3_U2917) );
  AOI22_X1 U21384 ( .A1(n18507), .A2(n18341), .B1(n18544), .B2(n18318), .ZN(
        n18308) );
  AOI22_X1 U21385 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18319), .B1(
        n18546), .B2(n18385), .ZN(n18307) );
  OAI211_X1 U21386 ( .C1(n18510), .C2(n18322), .A(n18308), .B(n18307), .ZN(
        P3_U2918) );
  AOI22_X1 U21387 ( .A1(n18511), .A2(n18341), .B1(n18551), .B2(n18318), .ZN(
        n18310) );
  AOI22_X1 U21388 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18319), .B1(
        n18552), .B2(n18385), .ZN(n18309) );
  OAI211_X1 U21389 ( .C1(n18514), .C2(n18322), .A(n18310), .B(n18309), .ZN(
        P3_U2919) );
  AOI22_X1 U21390 ( .A1(n18481), .A2(n18341), .B1(n18557), .B2(n18318), .ZN(
        n18312) );
  AOI22_X1 U21391 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18319), .B1(
        n18558), .B2(n18385), .ZN(n18311) );
  OAI211_X1 U21392 ( .C1(n18484), .C2(n18322), .A(n18312), .B(n18311), .ZN(
        P3_U2920) );
  AOI22_X1 U21393 ( .A1(n18562), .A2(n18318), .B1(n18563), .B2(n18341), .ZN(
        n18314) );
  AOI22_X1 U21394 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18319), .B1(
        n18564), .B2(n18385), .ZN(n18313) );
  OAI211_X1 U21395 ( .C1(n18567), .C2(n18322), .A(n18314), .B(n18313), .ZN(
        P3_U2921) );
  AOI22_X1 U21396 ( .A1(n18570), .A2(n18315), .B1(n18568), .B2(n18318), .ZN(
        n18317) );
  AOI22_X1 U21397 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18319), .B1(
        n18571), .B2(n18385), .ZN(n18316) );
  OAI211_X1 U21398 ( .C1(n18574), .C2(n18340), .A(n18317), .B(n18316), .ZN(
        P3_U2922) );
  AOI22_X1 U21399 ( .A1(n18578), .A2(n18341), .B1(n18577), .B2(n18318), .ZN(
        n18321) );
  AOI22_X1 U21400 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18319), .B1(
        n18580), .B2(n18385), .ZN(n18320) );
  OAI211_X1 U21401 ( .C1(n18586), .C2(n18322), .A(n18321), .B(n18320), .ZN(
        P3_U2923) );
  NOR2_X2 U21402 ( .A1(n18621), .A2(n18323), .ZN(n18408) );
  INV_X1 U21403 ( .A(n18408), .ZN(n18415) );
  AND2_X1 U21404 ( .A1(n18528), .A2(n18372), .ZN(n18342) );
  AOI22_X1 U21405 ( .A1(n18467), .A2(n18341), .B1(n18529), .B2(n18342), .ZN(
        n18327) );
  NAND2_X1 U21406 ( .A1(n18325), .A2(n18324), .ZN(n18343) );
  AOI22_X1 U21407 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18343), .B1(
        n18530), .B2(n18363), .ZN(n18326) );
  OAI211_X1 U21408 ( .C1(n18474), .C2(n18415), .A(n18327), .B(n18326), .ZN(
        P3_U2924) );
  AOI22_X1 U21409 ( .A1(n18445), .A2(n18363), .B1(n18538), .B2(n18342), .ZN(
        n18329) );
  AOI22_X1 U21410 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18343), .B1(
        n18540), .B2(n18408), .ZN(n18328) );
  OAI211_X1 U21411 ( .C1(n18448), .C2(n18340), .A(n18329), .B(n18328), .ZN(
        P3_U2925) );
  AOI22_X1 U21412 ( .A1(n18507), .A2(n18363), .B1(n18544), .B2(n18342), .ZN(
        n18331) );
  AOI22_X1 U21413 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18343), .B1(
        n18546), .B2(n18408), .ZN(n18330) );
  OAI211_X1 U21414 ( .C1(n18510), .C2(n18340), .A(n18331), .B(n18330), .ZN(
        P3_U2926) );
  AOI22_X1 U21415 ( .A1(n18551), .A2(n18342), .B1(n18550), .B2(n18341), .ZN(
        n18333) );
  AOI22_X1 U21416 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18343), .B1(
        n18552), .B2(n18408), .ZN(n18332) );
  OAI211_X1 U21417 ( .C1(n18555), .C2(n18362), .A(n18333), .B(n18332), .ZN(
        P3_U2927) );
  AOI22_X1 U21418 ( .A1(n18481), .A2(n18363), .B1(n18557), .B2(n18342), .ZN(
        n18335) );
  AOI22_X1 U21419 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18343), .B1(
        n18558), .B2(n18408), .ZN(n18334) );
  OAI211_X1 U21420 ( .C1(n18484), .C2(n18340), .A(n18335), .B(n18334), .ZN(
        P3_U2928) );
  AOI22_X1 U21421 ( .A1(n18562), .A2(n18342), .B1(n18563), .B2(n18363), .ZN(
        n18337) );
  AOI22_X1 U21422 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18343), .B1(
        n18564), .B2(n18408), .ZN(n18336) );
  OAI211_X1 U21423 ( .C1(n18567), .C2(n18340), .A(n18337), .B(n18336), .ZN(
        P3_U2929) );
  AOI22_X1 U21424 ( .A1(n18490), .A2(n18363), .B1(n18568), .B2(n18342), .ZN(
        n18339) );
  AOI22_X1 U21425 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18343), .B1(
        n18571), .B2(n18408), .ZN(n18338) );
  OAI211_X1 U21426 ( .C1(n18493), .C2(n18340), .A(n18339), .B(n18338), .ZN(
        P3_U2930) );
  AOI22_X1 U21427 ( .A1(n18577), .A2(n18342), .B1(n18364), .B2(n18341), .ZN(
        n18345) );
  AOI22_X1 U21428 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18343), .B1(
        n18580), .B2(n18408), .ZN(n18344) );
  OAI211_X1 U21429 ( .C1(n18369), .C2(n18362), .A(n18345), .B(n18344), .ZN(
        P3_U2931) );
  NAND2_X1 U21430 ( .A1(n18438), .A2(n18371), .ZN(n18437) );
  INV_X1 U21431 ( .A(n18437), .ZN(n18428) );
  NOR2_X1 U21432 ( .A1(n18408), .A2(n18428), .ZN(n18394) );
  NOR2_X1 U21433 ( .A1(n18654), .A2(n18394), .ZN(n18365) );
  AOI22_X1 U21434 ( .A1(n18530), .A2(n18385), .B1(n18529), .B2(n18365), .ZN(
        n18349) );
  OAI21_X1 U21435 ( .B1(n18346), .B2(n18440), .A(n18394), .ZN(n18347) );
  OAI211_X1 U21436 ( .C1(n18428), .C2(n18748), .A(n18393), .B(n18347), .ZN(
        n18366) );
  AOI22_X1 U21437 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18366), .B1(
        n18467), .B2(n18363), .ZN(n18348) );
  OAI211_X1 U21438 ( .C1(n18474), .C2(n18437), .A(n18349), .B(n18348), .ZN(
        P3_U2932) );
  AOI22_X1 U21439 ( .A1(n18445), .A2(n18385), .B1(n18538), .B2(n18365), .ZN(
        n18351) );
  AOI22_X1 U21440 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18366), .B1(
        n18540), .B2(n18428), .ZN(n18350) );
  OAI211_X1 U21441 ( .C1(n18448), .C2(n18362), .A(n18351), .B(n18350), .ZN(
        P3_U2933) );
  AOI22_X1 U21442 ( .A1(n18507), .A2(n18385), .B1(n18544), .B2(n18365), .ZN(
        n18353) );
  AOI22_X1 U21443 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18366), .B1(
        n18546), .B2(n18428), .ZN(n18352) );
  OAI211_X1 U21444 ( .C1(n18510), .C2(n18362), .A(n18353), .B(n18352), .ZN(
        P3_U2934) );
  AOI22_X1 U21445 ( .A1(n18551), .A2(n18365), .B1(n18550), .B2(n18363), .ZN(
        n18355) );
  AOI22_X1 U21446 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18366), .B1(
        n18552), .B2(n18428), .ZN(n18354) );
  OAI211_X1 U21447 ( .C1(n18555), .C2(n18391), .A(n18355), .B(n18354), .ZN(
        P3_U2935) );
  AOI22_X1 U21448 ( .A1(n18557), .A2(n18365), .B1(n18556), .B2(n18363), .ZN(
        n18357) );
  AOI22_X1 U21449 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18366), .B1(
        n18558), .B2(n18428), .ZN(n18356) );
  OAI211_X1 U21450 ( .C1(n18561), .C2(n18391), .A(n18357), .B(n18356), .ZN(
        P3_U2936) );
  AOI22_X1 U21451 ( .A1(n18562), .A2(n18365), .B1(n18563), .B2(n18385), .ZN(
        n18359) );
  AOI22_X1 U21452 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18366), .B1(
        n18564), .B2(n18428), .ZN(n18358) );
  OAI211_X1 U21453 ( .C1(n18567), .C2(n18362), .A(n18359), .B(n18358), .ZN(
        P3_U2937) );
  AOI22_X1 U21454 ( .A1(n18490), .A2(n18385), .B1(n18568), .B2(n18365), .ZN(
        n18361) );
  AOI22_X1 U21455 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18366), .B1(
        n18571), .B2(n18428), .ZN(n18360) );
  OAI211_X1 U21456 ( .C1(n18493), .C2(n18362), .A(n18361), .B(n18360), .ZN(
        P3_U2938) );
  AOI22_X1 U21457 ( .A1(n18577), .A2(n18365), .B1(n18364), .B2(n18363), .ZN(
        n18368) );
  AOI22_X1 U21458 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18366), .B1(
        n18580), .B2(n18428), .ZN(n18367) );
  OAI211_X1 U21459 ( .C1(n18369), .C2(n18391), .A(n18368), .B(n18367), .ZN(
        P3_U2939) );
  NAND2_X1 U21460 ( .A1(n18371), .A2(n18370), .ZN(n18464) );
  INV_X1 U21461 ( .A(n18371), .ZN(n18416) );
  NOR2_X1 U21462 ( .A1(n18416), .A2(n18465), .ZN(n18417) );
  AOI22_X1 U21463 ( .A1(n18467), .A2(n18385), .B1(n18529), .B2(n18417), .ZN(
        n18374) );
  AOI22_X1 U21464 ( .A1(n18471), .A2(n18372), .B1(n18371), .B2(n18468), .ZN(
        n18388) );
  AOI22_X1 U21465 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18388), .B1(
        n18530), .B2(n18408), .ZN(n18373) );
  OAI211_X1 U21466 ( .C1(n18474), .C2(n18464), .A(n18374), .B(n18373), .ZN(
        P3_U2940) );
  AOI22_X1 U21467 ( .A1(n18539), .A2(n18385), .B1(n18538), .B2(n18417), .ZN(
        n18376) );
  INV_X1 U21468 ( .A(n18464), .ZN(n18455) );
  AOI22_X1 U21469 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18388), .B1(
        n18540), .B2(n18455), .ZN(n18375) );
  OAI211_X1 U21470 ( .C1(n18543), .C2(n18415), .A(n18376), .B(n18375), .ZN(
        P3_U2941) );
  AOI22_X1 U21471 ( .A1(n18545), .A2(n18385), .B1(n18544), .B2(n18417), .ZN(
        n18378) );
  AOI22_X1 U21472 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18388), .B1(
        n18546), .B2(n18455), .ZN(n18377) );
  OAI211_X1 U21473 ( .C1(n18549), .C2(n18415), .A(n18378), .B(n18377), .ZN(
        P3_U2942) );
  AOI22_X1 U21474 ( .A1(n18551), .A2(n18417), .B1(n18550), .B2(n18385), .ZN(
        n18380) );
  AOI22_X1 U21475 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18388), .B1(
        n18552), .B2(n18455), .ZN(n18379) );
  OAI211_X1 U21476 ( .C1(n18555), .C2(n18415), .A(n18380), .B(n18379), .ZN(
        P3_U2943) );
  AOI22_X1 U21477 ( .A1(n18557), .A2(n18417), .B1(n18556), .B2(n18385), .ZN(
        n18382) );
  AOI22_X1 U21478 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18388), .B1(
        n18558), .B2(n18455), .ZN(n18381) );
  OAI211_X1 U21479 ( .C1(n18561), .C2(n18415), .A(n18382), .B(n18381), .ZN(
        P3_U2944) );
  AOI22_X1 U21480 ( .A1(n18562), .A2(n18417), .B1(n18563), .B2(n18408), .ZN(
        n18384) );
  AOI22_X1 U21481 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18388), .B1(
        n18564), .B2(n18455), .ZN(n18383) );
  OAI211_X1 U21482 ( .C1(n18567), .C2(n18391), .A(n18384), .B(n18383), .ZN(
        P3_U2945) );
  AOI22_X1 U21483 ( .A1(n18570), .A2(n18385), .B1(n18568), .B2(n18417), .ZN(
        n18387) );
  AOI22_X1 U21484 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18388), .B1(
        n18571), .B2(n18455), .ZN(n18386) );
  OAI211_X1 U21485 ( .C1(n18574), .C2(n18415), .A(n18387), .B(n18386), .ZN(
        P3_U2946) );
  AOI22_X1 U21486 ( .A1(n18578), .A2(n18408), .B1(n18577), .B2(n18417), .ZN(
        n18390) );
  AOI22_X1 U21487 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18388), .B1(
        n18580), .B2(n18455), .ZN(n18389) );
  OAI211_X1 U21488 ( .C1(n18586), .C2(n18391), .A(n18390), .B(n18389), .ZN(
        P3_U2947) );
  NOR2_X1 U21489 ( .A1(n20915), .A2(n18416), .ZN(n18470) );
  NAND2_X1 U21490 ( .A1(n18470), .A2(n18392), .ZN(n18497) );
  AOI21_X1 U21491 ( .B1(n18464), .B2(n18497), .A(n18654), .ZN(n18411) );
  AOI22_X1 U21492 ( .A1(n18467), .A2(n18408), .B1(n18529), .B2(n18411), .ZN(
        n18397) );
  OAI21_X1 U21493 ( .B1(n18455), .B2(n18485), .A(n18393), .ZN(n18439) );
  OAI21_X1 U21494 ( .B1(n18394), .B2(n18499), .A(n18439), .ZN(n18395) );
  OAI21_X1 U21495 ( .B1(n18485), .B2(n18748), .A(n18395), .ZN(n18412) );
  AOI22_X1 U21496 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18412), .B1(
        n18530), .B2(n18428), .ZN(n18396) );
  OAI211_X1 U21497 ( .C1(n18474), .C2(n18497), .A(n18397), .B(n18396), .ZN(
        P3_U2948) );
  AOI22_X1 U21498 ( .A1(n18445), .A2(n18428), .B1(n18538), .B2(n18411), .ZN(
        n18399) );
  AOI22_X1 U21499 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18412), .B1(
        n18540), .B2(n18485), .ZN(n18398) );
  OAI211_X1 U21500 ( .C1(n18448), .C2(n18415), .A(n18399), .B(n18398), .ZN(
        P3_U2949) );
  AOI22_X1 U21501 ( .A1(n18507), .A2(n18428), .B1(n18544), .B2(n18411), .ZN(
        n18401) );
  AOI22_X1 U21502 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18412), .B1(
        n18546), .B2(n18485), .ZN(n18400) );
  OAI211_X1 U21503 ( .C1(n18510), .C2(n18415), .A(n18401), .B(n18400), .ZN(
        P3_U2950) );
  AOI22_X1 U21504 ( .A1(n18551), .A2(n18411), .B1(n18550), .B2(n18408), .ZN(
        n18403) );
  AOI22_X1 U21505 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18412), .B1(
        n18552), .B2(n18485), .ZN(n18402) );
  OAI211_X1 U21506 ( .C1(n18555), .C2(n18437), .A(n18403), .B(n18402), .ZN(
        P3_U2951) );
  AOI22_X1 U21507 ( .A1(n18557), .A2(n18411), .B1(n18556), .B2(n18408), .ZN(
        n18405) );
  AOI22_X1 U21508 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18412), .B1(
        n18558), .B2(n18485), .ZN(n18404) );
  OAI211_X1 U21509 ( .C1(n18561), .C2(n18437), .A(n18405), .B(n18404), .ZN(
        P3_U2952) );
  AOI22_X1 U21510 ( .A1(n18486), .A2(n18408), .B1(n18562), .B2(n18411), .ZN(
        n18407) );
  AOI22_X1 U21511 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18412), .B1(
        n18563), .B2(n18428), .ZN(n18406) );
  OAI211_X1 U21512 ( .C1(n18489), .C2(n18497), .A(n18407), .B(n18406), .ZN(
        P3_U2953) );
  AOI22_X1 U21513 ( .A1(n18570), .A2(n18408), .B1(n18568), .B2(n18411), .ZN(
        n18410) );
  AOI22_X1 U21514 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18412), .B1(
        n18571), .B2(n18485), .ZN(n18409) );
  OAI211_X1 U21515 ( .C1(n18574), .C2(n18437), .A(n18410), .B(n18409), .ZN(
        P3_U2954) );
  AOI22_X1 U21516 ( .A1(n18578), .A2(n18428), .B1(n18577), .B2(n18411), .ZN(
        n18414) );
  AOI22_X1 U21517 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18412), .B1(
        n18580), .B2(n18485), .ZN(n18413) );
  OAI211_X1 U21518 ( .C1(n18586), .C2(n18415), .A(n18414), .B(n18413), .ZN(
        P3_U2955) );
  NOR2_X2 U21519 ( .A1(n18621), .A2(n18416), .ZN(n18519) );
  INV_X1 U21520 ( .A(n18519), .ZN(n18527) );
  AND2_X1 U21521 ( .A1(n18528), .A2(n18470), .ZN(n18433) );
  AOI22_X1 U21522 ( .A1(n18467), .A2(n18428), .B1(n18529), .B2(n18433), .ZN(
        n18419) );
  AOI22_X1 U21523 ( .A1(n18471), .A2(n18417), .B1(n18531), .B2(n18470), .ZN(
        n18434) );
  AOI22_X1 U21524 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18434), .B1(
        n18530), .B2(n18455), .ZN(n18418) );
  OAI211_X1 U21525 ( .C1(n18474), .C2(n18527), .A(n18419), .B(n18418), .ZN(
        P3_U2956) );
  AOI22_X1 U21526 ( .A1(n18445), .A2(n18455), .B1(n18538), .B2(n18433), .ZN(
        n18421) );
  AOI22_X1 U21527 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18434), .B1(
        n18540), .B2(n18519), .ZN(n18420) );
  OAI211_X1 U21528 ( .C1(n18448), .C2(n18437), .A(n18421), .B(n18420), .ZN(
        P3_U2957) );
  AOI22_X1 U21529 ( .A1(n18507), .A2(n18455), .B1(n18544), .B2(n18433), .ZN(
        n18423) );
  AOI22_X1 U21530 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18434), .B1(
        n18546), .B2(n18519), .ZN(n18422) );
  OAI211_X1 U21531 ( .C1(n18510), .C2(n18437), .A(n18423), .B(n18422), .ZN(
        P3_U2958) );
  AOI22_X1 U21532 ( .A1(n18551), .A2(n18433), .B1(n18550), .B2(n18428), .ZN(
        n18425) );
  AOI22_X1 U21533 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18434), .B1(
        n18552), .B2(n18519), .ZN(n18424) );
  OAI211_X1 U21534 ( .C1(n18555), .C2(n18464), .A(n18425), .B(n18424), .ZN(
        P3_U2959) );
  AOI22_X1 U21535 ( .A1(n18557), .A2(n18433), .B1(n18556), .B2(n18428), .ZN(
        n18427) );
  AOI22_X1 U21536 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18434), .B1(
        n18558), .B2(n18519), .ZN(n18426) );
  OAI211_X1 U21537 ( .C1(n18561), .C2(n18464), .A(n18427), .B(n18426), .ZN(
        P3_U2960) );
  AOI22_X1 U21538 ( .A1(n18486), .A2(n18428), .B1(n18562), .B2(n18433), .ZN(
        n18430) );
  AOI22_X1 U21539 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18434), .B1(
        n18563), .B2(n18455), .ZN(n18429) );
  OAI211_X1 U21540 ( .C1(n18489), .C2(n18527), .A(n18430), .B(n18429), .ZN(
        P3_U2961) );
  AOI22_X1 U21541 ( .A1(n18490), .A2(n18455), .B1(n18568), .B2(n18433), .ZN(
        n18432) );
  AOI22_X1 U21542 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18434), .B1(
        n18571), .B2(n18519), .ZN(n18431) );
  OAI211_X1 U21543 ( .C1(n18493), .C2(n18437), .A(n18432), .B(n18431), .ZN(
        P3_U2962) );
  AOI22_X1 U21544 ( .A1(n18578), .A2(n18455), .B1(n18577), .B2(n18433), .ZN(
        n18436) );
  AOI22_X1 U21545 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18434), .B1(
        n18580), .B2(n18519), .ZN(n18435) );
  OAI211_X1 U21546 ( .C1(n18586), .C2(n18437), .A(n18436), .B(n18435), .ZN(
        P3_U2963) );
  NAND2_X1 U21547 ( .A1(n18438), .A2(n18469), .ZN(n18585) );
  INV_X1 U21548 ( .A(n18585), .ZN(n18569) );
  NOR2_X1 U21549 ( .A1(n18519), .A2(n18569), .ZN(n18500) );
  NOR2_X1 U21550 ( .A1(n18654), .A2(n18500), .ZN(n18460) );
  AOI22_X1 U21551 ( .A1(n18467), .A2(n18455), .B1(n18529), .B2(n18460), .ZN(
        n18444) );
  OAI22_X1 U21552 ( .A1(n18500), .A2(n18441), .B1(n18440), .B2(n18439), .ZN(
        n18442) );
  OAI21_X1 U21553 ( .B1(n18569), .B2(n18748), .A(n18442), .ZN(n18461) );
  AOI22_X1 U21554 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18461), .B1(
        n18530), .B2(n18485), .ZN(n18443) );
  OAI211_X1 U21555 ( .C1(n18474), .C2(n18585), .A(n18444), .B(n18443), .ZN(
        P3_U2964) );
  AOI22_X1 U21556 ( .A1(n18445), .A2(n18485), .B1(n18538), .B2(n18460), .ZN(
        n18447) );
  AOI22_X1 U21557 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18461), .B1(
        n18540), .B2(n18569), .ZN(n18446) );
  OAI211_X1 U21558 ( .C1(n18448), .C2(n18464), .A(n18447), .B(n18446), .ZN(
        P3_U2965) );
  AOI22_X1 U21559 ( .A1(n18545), .A2(n18455), .B1(n18544), .B2(n18460), .ZN(
        n18450) );
  AOI22_X1 U21560 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18461), .B1(
        n18546), .B2(n18569), .ZN(n18449) );
  OAI211_X1 U21561 ( .C1(n18549), .C2(n18497), .A(n18450), .B(n18449), .ZN(
        P3_U2966) );
  AOI22_X1 U21562 ( .A1(n18511), .A2(n18485), .B1(n18551), .B2(n18460), .ZN(
        n18452) );
  AOI22_X1 U21563 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18461), .B1(
        n18552), .B2(n18569), .ZN(n18451) );
  OAI211_X1 U21564 ( .C1(n18514), .C2(n18464), .A(n18452), .B(n18451), .ZN(
        P3_U2967) );
  AOI22_X1 U21565 ( .A1(n18481), .A2(n18485), .B1(n18557), .B2(n18460), .ZN(
        n18454) );
  AOI22_X1 U21566 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18461), .B1(
        n18558), .B2(n18569), .ZN(n18453) );
  OAI211_X1 U21567 ( .C1(n18484), .C2(n18464), .A(n18454), .B(n18453), .ZN(
        P3_U2968) );
  AOI22_X1 U21568 ( .A1(n18486), .A2(n18455), .B1(n18562), .B2(n18460), .ZN(
        n18457) );
  AOI22_X1 U21569 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18461), .B1(
        n18563), .B2(n18485), .ZN(n18456) );
  OAI211_X1 U21570 ( .C1(n18489), .C2(n18585), .A(n18457), .B(n18456), .ZN(
        P3_U2969) );
  AOI22_X1 U21571 ( .A1(n18490), .A2(n18485), .B1(n18568), .B2(n18460), .ZN(
        n18459) );
  AOI22_X1 U21572 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18461), .B1(
        n18571), .B2(n18569), .ZN(n18458) );
  OAI211_X1 U21573 ( .C1(n18493), .C2(n18464), .A(n18459), .B(n18458), .ZN(
        P3_U2970) );
  AOI22_X1 U21574 ( .A1(n18578), .A2(n18485), .B1(n18577), .B2(n18460), .ZN(
        n18463) );
  AOI22_X1 U21575 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18461), .B1(
        n18580), .B2(n18569), .ZN(n18462) );
  OAI211_X1 U21576 ( .C1(n18586), .C2(n18464), .A(n18463), .B(n18462), .ZN(
        P3_U2971) );
  NOR2_X1 U21577 ( .A1(n18466), .A2(n18465), .ZN(n18533) );
  AOI22_X1 U21578 ( .A1(n18467), .A2(n18485), .B1(n18529), .B2(n18533), .ZN(
        n18473) );
  AOI22_X1 U21579 ( .A1(n18471), .A2(n18470), .B1(n18469), .B2(n18468), .ZN(
        n18494) );
  AOI22_X1 U21580 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18494), .B1(
        n18530), .B2(n18519), .ZN(n18472) );
  OAI211_X1 U21581 ( .C1(n18575), .C2(n18474), .A(n18473), .B(n18472), .ZN(
        P3_U2972) );
  AOI22_X1 U21582 ( .A1(n18539), .A2(n18485), .B1(n18538), .B2(n18533), .ZN(
        n18476) );
  AOI22_X1 U21583 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18494), .B1(
        n18579), .B2(n18540), .ZN(n18475) );
  OAI211_X1 U21584 ( .C1(n18543), .C2(n18527), .A(n18476), .B(n18475), .ZN(
        P3_U2973) );
  AOI22_X1 U21585 ( .A1(n18545), .A2(n18485), .B1(n18544), .B2(n18533), .ZN(
        n18478) );
  AOI22_X1 U21586 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18494), .B1(
        n18579), .B2(n18546), .ZN(n18477) );
  OAI211_X1 U21587 ( .C1(n18549), .C2(n18527), .A(n18478), .B(n18477), .ZN(
        P3_U2974) );
  AOI22_X1 U21588 ( .A1(n18551), .A2(n18533), .B1(n18550), .B2(n18485), .ZN(
        n18480) );
  AOI22_X1 U21589 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18494), .B1(
        n18579), .B2(n18552), .ZN(n18479) );
  OAI211_X1 U21590 ( .C1(n18555), .C2(n18527), .A(n18480), .B(n18479), .ZN(
        P3_U2975) );
  AOI22_X1 U21591 ( .A1(n18481), .A2(n18519), .B1(n18557), .B2(n18533), .ZN(
        n18483) );
  AOI22_X1 U21592 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18494), .B1(
        n18579), .B2(n18558), .ZN(n18482) );
  OAI211_X1 U21593 ( .C1(n18484), .C2(n18497), .A(n18483), .B(n18482), .ZN(
        P3_U2976) );
  AOI22_X1 U21594 ( .A1(n18486), .A2(n18485), .B1(n18562), .B2(n18533), .ZN(
        n18488) );
  AOI22_X1 U21595 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18494), .B1(
        n18563), .B2(n18519), .ZN(n18487) );
  OAI211_X1 U21596 ( .C1(n18575), .C2(n18489), .A(n18488), .B(n18487), .ZN(
        P3_U2977) );
  AOI22_X1 U21597 ( .A1(n18490), .A2(n18519), .B1(n18568), .B2(n18533), .ZN(
        n18492) );
  AOI22_X1 U21598 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18494), .B1(
        n18579), .B2(n18571), .ZN(n18491) );
  OAI211_X1 U21599 ( .C1(n18493), .C2(n18497), .A(n18492), .B(n18491), .ZN(
        P3_U2978) );
  AOI22_X1 U21600 ( .A1(n18578), .A2(n18519), .B1(n18577), .B2(n18533), .ZN(
        n18496) );
  AOI22_X1 U21601 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18494), .B1(
        n18579), .B2(n18580), .ZN(n18495) );
  OAI211_X1 U21602 ( .C1(n18586), .C2(n18497), .A(n18496), .B(n18495), .ZN(
        P3_U2979) );
  AOI21_X1 U21603 ( .B1(n18575), .B2(n18498), .A(n18654), .ZN(n18522) );
  AOI22_X1 U21604 ( .A1(n18530), .A2(n18569), .B1(n18529), .B2(n18522), .ZN(
        n18504) );
  NOR2_X1 U21605 ( .A1(n18500), .A2(n18499), .ZN(n18501) );
  OAI22_X1 U21606 ( .A1(n18523), .A2(n18748), .B1(n18502), .B2(n18501), .ZN(
        n18524) );
  AOI22_X1 U21607 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18524), .B1(
        n18523), .B2(n18534), .ZN(n18503) );
  OAI211_X1 U21608 ( .C1(n18537), .C2(n18527), .A(n18504), .B(n18503), .ZN(
        P3_U2980) );
  AOI22_X1 U21609 ( .A1(n18539), .A2(n18519), .B1(n18538), .B2(n18522), .ZN(
        n18506) );
  AOI22_X1 U21610 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18524), .B1(
        n18523), .B2(n18540), .ZN(n18505) );
  OAI211_X1 U21611 ( .C1(n18543), .C2(n18585), .A(n18506), .B(n18505), .ZN(
        P3_U2981) );
  AOI22_X1 U21612 ( .A1(n18507), .A2(n18569), .B1(n18544), .B2(n18522), .ZN(
        n18509) );
  AOI22_X1 U21613 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18524), .B1(
        n18523), .B2(n18546), .ZN(n18508) );
  OAI211_X1 U21614 ( .C1(n18510), .C2(n18527), .A(n18509), .B(n18508), .ZN(
        P3_U2982) );
  AOI22_X1 U21615 ( .A1(n18511), .A2(n18569), .B1(n18551), .B2(n18522), .ZN(
        n18513) );
  AOI22_X1 U21616 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18524), .B1(
        n18523), .B2(n18552), .ZN(n18512) );
  OAI211_X1 U21617 ( .C1(n18514), .C2(n18527), .A(n18513), .B(n18512), .ZN(
        P3_U2983) );
  AOI22_X1 U21618 ( .A1(n18557), .A2(n18522), .B1(n18556), .B2(n18519), .ZN(
        n18516) );
  AOI22_X1 U21619 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18524), .B1(
        n18523), .B2(n18558), .ZN(n18515) );
  OAI211_X1 U21620 ( .C1(n18561), .C2(n18585), .A(n18516), .B(n18515), .ZN(
        P3_U2984) );
  AOI22_X1 U21621 ( .A1(n18562), .A2(n18522), .B1(n18563), .B2(n18569), .ZN(
        n18518) );
  AOI22_X1 U21622 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18524), .B1(
        n18523), .B2(n18564), .ZN(n18517) );
  OAI211_X1 U21623 ( .C1(n18567), .C2(n18527), .A(n18518), .B(n18517), .ZN(
        P3_U2985) );
  AOI22_X1 U21624 ( .A1(n18570), .A2(n18519), .B1(n18568), .B2(n18522), .ZN(
        n18521) );
  AOI22_X1 U21625 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18524), .B1(
        n18523), .B2(n18571), .ZN(n18520) );
  OAI211_X1 U21626 ( .C1(n18574), .C2(n18585), .A(n18521), .B(n18520), .ZN(
        P3_U2986) );
  AOI22_X1 U21627 ( .A1(n18578), .A2(n18569), .B1(n18577), .B2(n18522), .ZN(
        n18526) );
  AOI22_X1 U21628 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18524), .B1(
        n18523), .B2(n18580), .ZN(n18525) );
  OAI211_X1 U21629 ( .C1(n18586), .C2(n18527), .A(n18526), .B(n18525), .ZN(
        P3_U2987) );
  AND2_X1 U21630 ( .A1(n18528), .A2(n18532), .ZN(n18576) );
  AOI22_X1 U21631 ( .A1(n18579), .A2(n18530), .B1(n18529), .B2(n18576), .ZN(
        n18536) );
  AOI22_X1 U21632 ( .A1(n18471), .A2(n18533), .B1(n18532), .B2(n18531), .ZN(
        n18582) );
  AOI22_X1 U21633 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18582), .B1(
        n18581), .B2(n18534), .ZN(n18535) );
  OAI211_X1 U21634 ( .C1(n18537), .C2(n18585), .A(n18536), .B(n18535), .ZN(
        P3_U2988) );
  AOI22_X1 U21635 ( .A1(n18539), .A2(n18569), .B1(n18538), .B2(n18576), .ZN(
        n18542) );
  AOI22_X1 U21636 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18582), .B1(
        n18581), .B2(n18540), .ZN(n18541) );
  OAI211_X1 U21637 ( .C1(n18575), .C2(n18543), .A(n18542), .B(n18541), .ZN(
        P3_U2989) );
  AOI22_X1 U21638 ( .A1(n18545), .A2(n18569), .B1(n18544), .B2(n18576), .ZN(
        n18548) );
  AOI22_X1 U21639 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18582), .B1(
        n18581), .B2(n18546), .ZN(n18547) );
  OAI211_X1 U21640 ( .C1(n18575), .C2(n18549), .A(n18548), .B(n18547), .ZN(
        P3_U2990) );
  AOI22_X1 U21641 ( .A1(n18551), .A2(n18576), .B1(n18550), .B2(n18569), .ZN(
        n18554) );
  AOI22_X1 U21642 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18582), .B1(
        n18581), .B2(n18552), .ZN(n18553) );
  OAI211_X1 U21643 ( .C1(n18575), .C2(n18555), .A(n18554), .B(n18553), .ZN(
        P3_U2991) );
  AOI22_X1 U21644 ( .A1(n18557), .A2(n18576), .B1(n18556), .B2(n18569), .ZN(
        n18560) );
  AOI22_X1 U21645 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18582), .B1(
        n18581), .B2(n18558), .ZN(n18559) );
  OAI211_X1 U21646 ( .C1(n18575), .C2(n18561), .A(n18560), .B(n18559), .ZN(
        P3_U2992) );
  AOI22_X1 U21647 ( .A1(n18579), .A2(n18563), .B1(n18562), .B2(n18576), .ZN(
        n18566) );
  AOI22_X1 U21648 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18582), .B1(
        n18581), .B2(n18564), .ZN(n18565) );
  OAI211_X1 U21649 ( .C1(n18567), .C2(n18585), .A(n18566), .B(n18565), .ZN(
        P3_U2993) );
  AOI22_X1 U21650 ( .A1(n18570), .A2(n18569), .B1(n18568), .B2(n18576), .ZN(
        n18573) );
  AOI22_X1 U21651 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18582), .B1(
        n18581), .B2(n18571), .ZN(n18572) );
  OAI211_X1 U21652 ( .C1(n18575), .C2(n18574), .A(n18573), .B(n18572), .ZN(
        P3_U2994) );
  AOI22_X1 U21653 ( .A1(n18579), .A2(n18578), .B1(n18577), .B2(n18576), .ZN(
        n18584) );
  AOI22_X1 U21654 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18582), .B1(
        n18581), .B2(n18580), .ZN(n18583) );
  OAI211_X1 U21655 ( .C1(n18586), .C2(n18585), .A(n18584), .B(n18583), .ZN(
        P3_U2995) );
  INV_X1 U21656 ( .A(n18587), .ZN(n18590) );
  OAI21_X1 U21657 ( .B1(n18590), .B2(n18589), .A(n18588), .ZN(n18599) );
  AOI22_X1 U21658 ( .A1(n18762), .A2(n18601), .B1(n18591), .B2(n18599), .ZN(
        n18592) );
  OAI21_X1 U21659 ( .B1(n18593), .B2(n18595), .A(n18592), .ZN(n18753) );
  NOR2_X1 U21660 ( .A1(n18633), .A2(n18753), .ZN(n18598) );
  NOR2_X1 U21661 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18594), .ZN(
        n18618) );
  INV_X1 U21662 ( .A(n18595), .ZN(n18607) );
  OAI22_X1 U21663 ( .A1(n18596), .A2(n18629), .B1(n18618), .B2(n18607), .ZN(
        n18750) );
  NAND2_X1 U21664 ( .A1(n18754), .A2(n18750), .ZN(n18597) );
  OAI22_X1 U21665 ( .A1(n18598), .A2(n18754), .B1(n18633), .B2(n18597), .ZN(
        n18640) );
  AOI21_X1 U21666 ( .B1(n18769), .B2(n18600), .A(n18599), .ZN(n18612) );
  NAND2_X1 U21667 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18601), .ZN(
        n18611) );
  INV_X1 U21668 ( .A(n18759), .ZN(n18605) );
  NAND2_X1 U21669 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18615), .ZN(
        n18602) );
  AOI211_X1 U21670 ( .C1(n18603), .C2(n18602), .A(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n18769), .ZN(n18604) );
  AOI21_X1 U21671 ( .B1(n18606), .B2(n18605), .A(n18604), .ZN(n18610) );
  OAI211_X1 U21672 ( .C1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n18608), .B(n18607), .ZN(
        n18609) );
  OAI211_X1 U21673 ( .C1(n18612), .C2(n18611), .A(n18610), .B(n18609), .ZN(
        n18760) );
  AOI22_X1 U21674 ( .A1(n18633), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n18760), .B2(n18613), .ZN(n18614) );
  OAI21_X1 U21675 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n18614), .ZN(n18639) );
  INV_X1 U21676 ( .A(n18640), .ZN(n18628) );
  INV_X1 U21677 ( .A(n18614), .ZN(n18625) );
  NOR2_X1 U21678 ( .A1(n18616), .A2(n18615), .ZN(n18620) );
  AOI22_X1 U21679 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18617), .B1(
        n18620), .B2(n18774), .ZN(n18771) );
  OAI22_X1 U21680 ( .A1(n18620), .A2(n18619), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18618), .ZN(n18767) );
  AOI222_X1 U21681 ( .A1(n18771), .A2(n18767), .B1(n18771), .B2(n20915), .C1(
        n18767), .C2(n18621), .ZN(n18623) );
  OAI21_X1 U21682 ( .B1(n18633), .B2(n18623), .A(n18622), .ZN(n18624) );
  AOI222_X1 U21683 ( .A1(n18626), .A2(n18625), .B1(n18626), .B2(n18624), .C1(
        n18625), .C2(n18624), .ZN(n18627) );
  AOI211_X1 U21684 ( .C1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n18628), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B(n18627), .ZN(n18638) );
  OAI22_X1 U21685 ( .A1(n18631), .A2(n18630), .B1(n18788), .B2(n18629), .ZN(
        n18789) );
  AOI211_X1 U21686 ( .C1(n18633), .C2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n18632), .B(n18789), .ZN(n18636) );
  OAI21_X1 U21687 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18634), .ZN(n18635) );
  NAND4_X1 U21688 ( .A1(n18636), .A2(n18785), .A3(n18787), .A4(n18635), .ZN(
        n18637) );
  AOI211_X1 U21689 ( .C1(n18640), .C2(n18639), .A(n18638), .B(n18637), .ZN(
        n18652) );
  INV_X1 U21690 ( .A(n18798), .ZN(n18641) );
  AOI22_X1 U21691 ( .A1(n18770), .A2(n18641), .B1(n18796), .B2(n18804), .ZN(
        n18642) );
  INV_X1 U21692 ( .A(n18642), .ZN(n18648) );
  OAI211_X1 U21693 ( .C1(n18645), .C2(n18644), .A(n18643), .B(n18652), .ZN(
        n18747) );
  OAI21_X1 U21694 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18803), .A(n18747), 
        .ZN(n18653) );
  NOR2_X1 U21695 ( .A1(n18646), .A2(n18653), .ZN(n18647) );
  MUX2_X1 U21696 ( .A(n18648), .B(n18647), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18650) );
  OAI211_X1 U21697 ( .C1(n18652), .C2(n18651), .A(n18650), .B(n18649), .ZN(
        P3_U2996) );
  NAND3_X1 U21698 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18796), .A3(n18809), 
        .ZN(n18659) );
  NOR2_X1 U21699 ( .A1(n18654), .A2(n18653), .ZN(n18655) );
  AOI22_X1 U21700 ( .A1(n18796), .A2(n18804), .B1(n18656), .B2(n18655), .ZN(
        n18658) );
  OAI211_X1 U21701 ( .C1(n18757), .C2(n18659), .A(n18658), .B(n18657), .ZN(
        P3_U2997) );
  AND4_X1 U21702 ( .A1(n18798), .A2(n18660), .A3(n18659), .A4(n18746), .ZN(
        P3_U2998) );
  AND2_X1 U21703 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18742), .ZN(
        P3_U2999) );
  INV_X1 U21704 ( .A(P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n20989) );
  NOR2_X1 U21705 ( .A1(n20989), .A2(n18745), .ZN(P3_U3000) );
  INV_X1 U21706 ( .A(P3_DATAWIDTH_REG_29__SCAN_IN), .ZN(n21031) );
  NOR2_X1 U21707 ( .A1(n21031), .A2(n18745), .ZN(P3_U3001) );
  AND2_X1 U21708 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18742), .ZN(
        P3_U3002) );
  AND2_X1 U21709 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18742), .ZN(
        P3_U3003) );
  AND2_X1 U21710 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18742), .ZN(
        P3_U3004) );
  AND2_X1 U21711 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18742), .ZN(
        P3_U3005) );
  AND2_X1 U21712 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18742), .ZN(
        P3_U3006) );
  AND2_X1 U21713 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18742), .ZN(
        P3_U3007) );
  AND2_X1 U21714 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18742), .ZN(
        P3_U3008) );
  AND2_X1 U21715 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18742), .ZN(
        P3_U3009) );
  AND2_X1 U21716 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18742), .ZN(
        P3_U3010) );
  AND2_X1 U21717 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18742), .ZN(
        P3_U3011) );
  AND2_X1 U21718 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18742), .ZN(
        P3_U3012) );
  INV_X1 U21719 ( .A(P3_DATAWIDTH_REG_17__SCAN_IN), .ZN(n21078) );
  NOR2_X1 U21720 ( .A1(n21078), .A2(n18745), .ZN(P3_U3013) );
  AND2_X1 U21721 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18742), .ZN(
        P3_U3014) );
  AND2_X1 U21722 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18742), .ZN(
        P3_U3015) );
  AND2_X1 U21723 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18742), .ZN(
        P3_U3016) );
  AND2_X1 U21724 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18742), .ZN(
        P3_U3017) );
  AND2_X1 U21725 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18742), .ZN(
        P3_U3018) );
  AND2_X1 U21726 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18742), .ZN(
        P3_U3019) );
  AND2_X1 U21727 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18742), .ZN(
        P3_U3020) );
  AND2_X1 U21728 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18742), .ZN(P3_U3021) );
  INV_X1 U21729 ( .A(P3_DATAWIDTH_REG_8__SCAN_IN), .ZN(n20979) );
  NOR2_X1 U21730 ( .A1(n20979), .A2(n18745), .ZN(P3_U3022) );
  AND2_X1 U21731 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18742), .ZN(P3_U3023) );
  AND2_X1 U21732 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18742), .ZN(P3_U3024) );
  AND2_X1 U21733 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18742), .ZN(P3_U3025) );
  AND2_X1 U21734 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18742), .ZN(P3_U3026) );
  AND2_X1 U21735 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18742), .ZN(P3_U3027) );
  AND2_X1 U21736 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18742), .ZN(P3_U3028) );
  NAND2_X1 U21737 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n18666) );
  INV_X1 U21738 ( .A(n18666), .ZN(n18661) );
  NOR2_X1 U21739 ( .A1(n18677), .A2(n20723), .ZN(n18672) );
  INV_X1 U21740 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18665) );
  NOR3_X1 U21741 ( .A1(n18661), .A2(n18672), .A3(n18665), .ZN(n18664) );
  AOI21_X1 U21742 ( .B1(n18796), .B2(P3_STATE_REG_1__SCAN_IN), .A(n18674), 
        .ZN(n18676) );
  INV_X1 U21743 ( .A(NA), .ZN(n20718) );
  OAI21_X1 U21744 ( .B1(n20718), .B2(n18662), .A(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18675) );
  INV_X1 U21745 ( .A(n18675), .ZN(n18663) );
  OAI22_X1 U21746 ( .A1(n18739), .A2(n18664), .B1(n18676), .B2(n18663), .ZN(
        P3_U3029) );
  OAI22_X1 U21747 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n18666), .B1(n18672), 
        .B2(n18665), .ZN(n18667) );
  AOI22_X1 U21748 ( .A1(n18796), .A2(P3_STATE_REG_1__SCAN_IN), .B1(
        P3_STATE_REG_0__SCAN_IN), .B2(n18667), .ZN(n18669) );
  NAND2_X1 U21749 ( .A1(n18669), .A2(n18668), .ZN(P3_U3030) );
  NAND2_X1 U21750 ( .A1(n18796), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18670) );
  OAI22_X1 U21751 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18670), .ZN(n18671) );
  OAI22_X1 U21752 ( .A1(n18672), .A2(n18671), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18673) );
  OAI22_X1 U21753 ( .A1(n18676), .A2(n18675), .B1(n18674), .B2(n18673), .ZN(
        P3_U3031) );
  OAI222_X1 U21754 ( .A1(n18720), .A2(n21028), .B1(n18678), .B2(n18739), .C1(
        n18776), .C2(n18732), .ZN(P3_U3032) );
  INV_X1 U21755 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18680) );
  OAI222_X1 U21756 ( .A1(n18720), .A2(n18680), .B1(n18679), .B2(n18739), .C1(
        n21028), .C2(n18732), .ZN(P3_U3033) );
  OAI222_X1 U21757 ( .A1(n18720), .A2(n18681), .B1(n21038), .B2(n18739), .C1(
        n18680), .C2(n18732), .ZN(P3_U3034) );
  OAI222_X1 U21758 ( .A1(n18720), .A2(n18683), .B1(n18682), .B2(n18739), .C1(
        n18681), .C2(n18732), .ZN(P3_U3035) );
  OAI222_X1 U21759 ( .A1(n18720), .A2(n20952), .B1(n18684), .B2(n18739), .C1(
        n18683), .C2(n18732), .ZN(P3_U3036) );
  OAI222_X1 U21760 ( .A1(n18720), .A2(n18686), .B1(n18685), .B2(n18739), .C1(
        n20952), .C2(n18732), .ZN(P3_U3037) );
  OAI222_X1 U21761 ( .A1(n18720), .A2(n21043), .B1(n18687), .B2(n18739), .C1(
        n18686), .C2(n18732), .ZN(P3_U3038) );
  OAI222_X1 U21762 ( .A1(n21043), .A2(n18732), .B1(n18688), .B2(n18739), .C1(
        n18689), .C2(n18720), .ZN(P3_U3039) );
  INV_X1 U21763 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18691) );
  OAI222_X1 U21764 ( .A1(n18720), .A2(n18691), .B1(n18690), .B2(n18739), .C1(
        n18689), .C2(n18732), .ZN(P3_U3040) );
  OAI222_X1 U21765 ( .A1(n18720), .A2(n20924), .B1(n18692), .B2(n18739), .C1(
        n18691), .C2(n18732), .ZN(P3_U3041) );
  INV_X1 U21766 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18693) );
  OAI222_X1 U21767 ( .A1(n18720), .A2(n18693), .B1(n20957), .B2(n18739), .C1(
        n20924), .C2(n18732), .ZN(P3_U3042) );
  OAI222_X1 U21768 ( .A1(n18720), .A2(n18696), .B1(n18694), .B2(n18739), .C1(
        n18693), .C2(n18732), .ZN(P3_U3043) );
  OAI222_X1 U21769 ( .A1(n18696), .A2(n18732), .B1(n18695), .B2(n18739), .C1(
        n18698), .C2(n18720), .ZN(P3_U3044) );
  OAI222_X1 U21770 ( .A1(n18698), .A2(n18732), .B1(n18697), .B2(n18739), .C1(
        n18699), .C2(n18720), .ZN(P3_U3045) );
  OAI222_X1 U21771 ( .A1(n18720), .A2(n20890), .B1(n18700), .B2(n18739), .C1(
        n18699), .C2(n18732), .ZN(P3_U3046) );
  OAI222_X1 U21772 ( .A1(n18720), .A2(n18702), .B1(n18701), .B2(n18739), .C1(
        n20890), .C2(n18732), .ZN(P3_U3047) );
  OAI222_X1 U21773 ( .A1(n18720), .A2(n18704), .B1(n18703), .B2(n18739), .C1(
        n18702), .C2(n18732), .ZN(P3_U3048) );
  INV_X1 U21774 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18707) );
  OAI222_X1 U21775 ( .A1(n18720), .A2(n18707), .B1(n18705), .B2(n18739), .C1(
        n18704), .C2(n18732), .ZN(P3_U3049) );
  OAI222_X1 U21776 ( .A1(n18707), .A2(n18732), .B1(n18706), .B2(n18739), .C1(
        n18708), .C2(n18720), .ZN(P3_U3050) );
  OAI222_X1 U21777 ( .A1(n18720), .A2(n18711), .B1(n18709), .B2(n18739), .C1(
        n18708), .C2(n18732), .ZN(P3_U3051) );
  OAI222_X1 U21778 ( .A1(n18711), .A2(n18732), .B1(n18710), .B2(n18739), .C1(
        n18712), .C2(n18720), .ZN(P3_U3052) );
  INV_X1 U21779 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18715) );
  OAI222_X1 U21780 ( .A1(n18720), .A2(n18715), .B1(n18713), .B2(n18739), .C1(
        n18712), .C2(n18732), .ZN(P3_U3053) );
  OAI222_X1 U21781 ( .A1(n18715), .A2(n18732), .B1(n18714), .B2(n18739), .C1(
        n18716), .C2(n18720), .ZN(P3_U3054) );
  INV_X1 U21782 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18718) );
  OAI222_X1 U21783 ( .A1(n18720), .A2(n18718), .B1(n18717), .B2(n18739), .C1(
        n18716), .C2(n18732), .ZN(P3_U3055) );
  INV_X1 U21784 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18721) );
  OAI222_X1 U21785 ( .A1(n18720), .A2(n18721), .B1(n18719), .B2(n18739), .C1(
        n18718), .C2(n18732), .ZN(P3_U3056) );
  OAI222_X1 U21786 ( .A1(n18720), .A2(n18723), .B1(n18722), .B2(n18739), .C1(
        n18721), .C2(n18732), .ZN(P3_U3057) );
  INV_X1 U21787 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18726) );
  OAI222_X1 U21788 ( .A1(n18720), .A2(n18726), .B1(n18724), .B2(n18739), .C1(
        n18723), .C2(n18732), .ZN(P3_U3058) );
  INV_X1 U21789 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18727) );
  OAI222_X1 U21790 ( .A1(n18726), .A2(n18732), .B1(n18725), .B2(n18739), .C1(
        n18727), .C2(n18720), .ZN(P3_U3059) );
  OAI222_X1 U21791 ( .A1(n18720), .A2(n18731), .B1(n18728), .B2(n18739), .C1(
        n18727), .C2(n18732), .ZN(P3_U3060) );
  OAI222_X1 U21792 ( .A1(n18732), .A2(n18731), .B1(n18730), .B2(n18739), .C1(
        n18729), .C2(n18720), .ZN(P3_U3061) );
  INV_X1 U21793 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n18733) );
  AOI22_X1 U21794 ( .A1(n18739), .A2(n18734), .B1(n18733), .B2(n18807), .ZN(
        P3_U3274) );
  INV_X1 U21795 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18779) );
  INV_X1 U21796 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n18735) );
  AOI22_X1 U21797 ( .A1(n18739), .A2(n18779), .B1(n18735), .B2(n18807), .ZN(
        P3_U3275) );
  INV_X1 U21798 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n18736) );
  AOI22_X1 U21799 ( .A1(n18739), .A2(n18737), .B1(n18736), .B2(n18807), .ZN(
        P3_U3276) );
  INV_X1 U21800 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18782) );
  INV_X1 U21801 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n18738) );
  AOI22_X1 U21802 ( .A1(n18739), .A2(n18782), .B1(n18738), .B2(n18807), .ZN(
        P3_U3277) );
  INV_X1 U21803 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18741) );
  AOI21_X1 U21804 ( .B1(n18742), .B2(n18741), .A(n18740), .ZN(P3_U3280) );
  OAI21_X1 U21805 ( .B1(n18745), .B2(n18744), .A(n18743), .ZN(P3_U3281) );
  OAI221_X1 U21806 ( .B1(n18748), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18748), 
        .C2(n18747), .A(n18746), .ZN(P3_U3282) );
  NOR2_X1 U21807 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18749), .ZN(
        n18751) );
  AOI22_X1 U21808 ( .A1(n18770), .A2(n18752), .B1(n18751), .B2(n18750), .ZN(
        n18756) );
  AOI21_X1 U21809 ( .B1(n18810), .B2(n18753), .A(n18775), .ZN(n18755) );
  OAI22_X1 U21810 ( .A1(n18775), .A2(n18756), .B1(n18755), .B2(n18754), .ZN(
        P3_U3285) );
  NOR2_X1 U21811 ( .A1(n18757), .A2(n21053), .ZN(n18764) );
  AOI22_X1 U21812 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n21073), .B2(n18758), .ZN(
        n18763) );
  AOI222_X1 U21813 ( .A1(n18760), .A2(n18810), .B1(n18764), .B2(n18763), .C1(
        n18770), .C2(n18759), .ZN(n18761) );
  AOI22_X1 U21814 ( .A1(n18775), .A2(n18762), .B1(n18761), .B2(n18772), .ZN(
        P3_U3288) );
  INV_X1 U21815 ( .A(n18763), .ZN(n18765) );
  AOI222_X1 U21816 ( .A1(n18767), .A2(n18810), .B1(n18770), .B2(n18766), .C1(
        n18765), .C2(n18764), .ZN(n18768) );
  AOI22_X1 U21817 ( .A1(n18775), .A2(n18769), .B1(n18768), .B2(n18772), .ZN(
        P3_U3289) );
  AOI222_X1 U21818 ( .A1(n21053), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18810), 
        .B2(n18771), .C1(n18774), .C2(n18770), .ZN(n18773) );
  AOI22_X1 U21819 ( .A1(n18775), .A2(n18774), .B1(n18773), .B2(n18772), .ZN(
        P3_U3290) );
  AOI21_X1 U21820 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18777) );
  AOI22_X1 U21821 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18777), .B2(n18776), .ZN(n18780) );
  AOI22_X1 U21822 ( .A1(n18783), .A2(n18780), .B1(n18779), .B2(n18778), .ZN(
        P3_U3292) );
  OAI21_X1 U21823 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18783), .ZN(n18781) );
  OAI21_X1 U21824 ( .B1(n18783), .B2(n18782), .A(n18781), .ZN(P3_U3293) );
  INV_X1 U21825 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18784) );
  AOI22_X1 U21826 ( .A1(n18739), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18784), 
        .B2(n18807), .ZN(P3_U3294) );
  INV_X1 U21827 ( .A(P3_MORE_REG_SCAN_IN), .ZN(n18792) );
  OAI22_X1 U21828 ( .A1(n18788), .A2(n18787), .B1(n18786), .B2(n18785), .ZN(
        n18790) );
  OAI21_X1 U21829 ( .B1(n18790), .B2(n18789), .A(n18793), .ZN(n18791) );
  OAI21_X1 U21830 ( .B1(n18793), .B2(n18792), .A(n18791), .ZN(P3_U3295) );
  OAI21_X1 U21831 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n18795), .A(n18794), 
        .ZN(n18797) );
  AOI211_X1 U21832 ( .C1(n18811), .C2(n18797), .A(n18796), .B(n18809), .ZN(
        n18800) );
  OAI21_X1 U21833 ( .B1(n18800), .B2(n18799), .A(n18798), .ZN(n18806) );
  AOI21_X1 U21834 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_2__SCAN_IN), .A(n18801), .ZN(n18802) );
  AOI211_X1 U21835 ( .C1(n18804), .C2(n18803), .A(n18802), .B(n18812), .ZN(
        n18805) );
  MUX2_X1 U21836 ( .A(n18806), .B(P3_REQUESTPENDING_REG_SCAN_IN), .S(n18805), 
        .Z(P3_U3296) );
  INV_X1 U21837 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18815) );
  INV_X1 U21838 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n18808) );
  AOI22_X1 U21839 ( .A1(n18739), .A2(n18815), .B1(n18808), .B2(n18807), .ZN(
        P3_U3297) );
  AOI21_X1 U21840 ( .B1(n18810), .B2(n18809), .A(n18812), .ZN(n18816) );
  INV_X1 U21841 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18813) );
  AOI22_X1 U21842 ( .A1(n18816), .A2(n18813), .B1(n18812), .B2(n18811), .ZN(
        P3_U3298) );
  AOI21_X1 U21843 ( .B1(n18816), .B2(n18815), .A(n18814), .ZN(P3_U3299) );
  INV_X1 U21844 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n18817) );
  NAND2_X1 U21845 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19752), .ZN(n19743) );
  NAND2_X1 U21846 ( .A1(n18818), .A2(n19736), .ZN(n19744) );
  OAI21_X1 U21847 ( .B1(n18818), .B2(n19743), .A(n19744), .ZN(n19807) );
  OAI21_X1 U21848 ( .B1(n18818), .B2(n18817), .A(n19804), .ZN(P2_U2815) );
  INV_X1 U21849 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18820) );
  OAI22_X1 U21850 ( .A1(n19854), .A2(n18820), .B1(n19859), .B2(n18819), .ZN(
        P2_U2816) );
  AOI22_X1 U21851 ( .A1(n19792), .A2(n18820), .B1(P2_D_C_N_REG_SCAN_IN), .B2(
        n19869), .ZN(n18821) );
  OAI21_X1 U21852 ( .B1(P2_STATE_REG_2__SCAN_IN), .B2(n19744), .A(n18821), 
        .ZN(P2_U2817) );
  AOI21_X1 U21853 ( .B1(n19748), .B2(n18822), .A(n19804), .ZN(n19802) );
  INV_X1 U21854 ( .A(n19802), .ZN(n19805) );
  OAI21_X1 U21855 ( .B1(n19807), .B2(n19626), .A(n19805), .ZN(P2_U2818) );
  NOR4_X1 U21856 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18832) );
  NOR4_X1 U21857 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18831) );
  NOR4_X1 U21858 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18823) );
  INV_X1 U21859 ( .A(P2_DATAWIDTH_REG_21__SCAN_IN), .ZN(n21037) );
  INV_X1 U21860 ( .A(P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n21006) );
  NAND3_X1 U21861 ( .A1(n18823), .A2(n21037), .A3(n21006), .ZN(n18829) );
  NOR4_X1 U21862 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18827) );
  NOR4_X1 U21863 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18826) );
  NOR4_X1 U21864 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18825) );
  NOR4_X1 U21865 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18824) );
  NAND4_X1 U21866 ( .A1(n18827), .A2(n18826), .A3(n18825), .A4(n18824), .ZN(
        n18828) );
  AOI211_X1 U21867 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(n18829), .B(n18828), .ZN(n18830) );
  NAND3_X1 U21868 ( .A1(n18832), .A2(n18831), .A3(n18830), .ZN(n18833) );
  NOR2_X1 U21869 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18833), .ZN(n18835) );
  INV_X1 U21870 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19801) );
  AOI22_X1 U21871 ( .A1(n18835), .A2(n18836), .B1(n18833), .B2(n19801), .ZN(
        P2_U2820) );
  INV_X1 U21872 ( .A(n18833), .ZN(n18841) );
  NOR2_X1 U21873 ( .A1(n18841), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18834)
         );
  INV_X1 U21874 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19806) );
  INV_X1 U21875 ( .A(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19803) );
  NAND4_X1 U21876 ( .A1(n18841), .A2(n18836), .A3(n19806), .A4(n19803), .ZN(
        n18840) );
  OAI21_X1 U21877 ( .B1(n18835), .B2(n18834), .A(n18840), .ZN(P2_U2821) );
  NAND2_X1 U21878 ( .A1(n18835), .A2(n19806), .ZN(n18839) );
  OAI21_X1 U21879 ( .B1(n18836), .B2(n19754), .A(n18841), .ZN(n18837) );
  OAI21_X1 U21880 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18841), .A(n18837), 
        .ZN(n18838) );
  OAI221_X1 U21881 ( .B1(n18839), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18839), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18838), .ZN(P2_U2822) );
  INV_X1 U21882 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19799) );
  OAI211_X1 U21883 ( .C1(n18841), .C2(n19799), .A(n18840), .B(n18839), .ZN(
        P2_U2823) );
  AOI22_X1 U21884 ( .A1(P2_REIP_REG_20__SCAN_IN), .A2(n18993), .B1(
        P2_EBX_REG_20__SCAN_IN), .B2(n18978), .ZN(n18853) );
  AOI22_X1 U21885 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18968), .B1(
        n18928), .B2(n18842), .ZN(n18852) );
  INV_X1 U21886 ( .A(n18843), .ZN(n18845) );
  AOI22_X1 U21887 ( .A1(n18845), .A2(n18984), .B1(n18844), .B2(n18979), .ZN(
        n18851) );
  AOI21_X1 U21888 ( .B1(n18848), .B2(n18846), .A(n18847), .ZN(n18849) );
  NAND2_X1 U21889 ( .A1(n18961), .A2(n18849), .ZN(n18850) );
  NAND4_X1 U21890 ( .A1(n18853), .A2(n18852), .A3(n18851), .A4(n18850), .ZN(
        P2_U2835) );
  OAI22_X1 U21891 ( .A1(n19776), .A2(n18938), .B1(n18854), .B2(n18982), .ZN(
        n18855) );
  AOI211_X1 U21892 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n18978), .A(n19138), .B(
        n18855), .ZN(n18864) );
  AOI211_X1 U21893 ( .C1(n18858), .C2(n18857), .A(n18856), .B(n19732), .ZN(
        n18862) );
  OAI22_X1 U21894 ( .A1(n18860), .A2(n18973), .B1(n18859), .B2(n18958), .ZN(
        n18861) );
  NOR2_X1 U21895 ( .A1(n18862), .A2(n18861), .ZN(n18863) );
  OAI211_X1 U21896 ( .C1(n18865), .C2(n18990), .A(n18864), .B(n18863), .ZN(
        P2_U2836) );
  NOR2_X1 U21897 ( .A1(n18966), .A2(n18866), .ZN(n18868) );
  XOR2_X1 U21898 ( .A(n18868), .B(n18867), .Z(n18877) );
  INV_X1 U21899 ( .A(n18869), .ZN(n18871) );
  AOI22_X1 U21900 ( .A1(P2_REIP_REG_16__SCAN_IN), .A2(n18993), .B1(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n18968), .ZN(n18870) );
  OAI21_X1 U21901 ( .B1(n18871), .B2(n18982), .A(n18870), .ZN(n18872) );
  AOI211_X1 U21902 ( .C1(P2_EBX_REG_16__SCAN_IN), .C2(n18978), .A(n19138), .B(
        n18872), .ZN(n18876) );
  AOI22_X1 U21903 ( .A1(n18874), .A2(n18984), .B1(n18979), .B2(n18873), .ZN(
        n18875) );
  OAI211_X1 U21904 ( .C1(n19732), .C2(n18877), .A(n18876), .B(n18875), .ZN(
        P2_U2839) );
  OAI21_X1 U21905 ( .B1(n11400), .B2(n18938), .A(n18878), .ZN(n18881) );
  OAI22_X1 U21906 ( .A1(n10870), .A2(n18950), .B1(n18879), .B2(n18982), .ZN(
        n18880) );
  AOI211_X1 U21907 ( .C1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .C2(n18968), .A(
        n18881), .B(n18880), .ZN(n18888) );
  NOR2_X1 U21908 ( .A1(n18966), .A2(n18882), .ZN(n18884) );
  XNOR2_X1 U21909 ( .A(n18884), .B(n18883), .ZN(n18886) );
  AOI22_X1 U21910 ( .A1(n18886), .A2(n18961), .B1(n18984), .B2(n18885), .ZN(
        n18887) );
  OAI211_X1 U21911 ( .C1(n19004), .C2(n18958), .A(n18888), .B(n18887), .ZN(
        P2_U2841) );
  OAI22_X1 U21912 ( .A1(n18890), .A2(n18990), .B1(n18889), .B2(n18982), .ZN(
        n18891) );
  AOI211_X1 U21913 ( .C1(P2_EBX_REG_13__SCAN_IN), .C2(n18978), .A(n19138), .B(
        n18891), .ZN(n18900) );
  NAND2_X1 U21914 ( .A1(n18954), .A2(n18892), .ZN(n18893) );
  XNOR2_X1 U21915 ( .A(n18894), .B(n18893), .ZN(n18898) );
  OAI22_X1 U21916 ( .A1(n18896), .A2(n18973), .B1(n18958), .B2(n18895), .ZN(
        n18897) );
  AOI21_X1 U21917 ( .B1(n18961), .B2(n18898), .A(n18897), .ZN(n18899) );
  OAI211_X1 U21918 ( .C1(n11397), .C2(n18938), .A(n18900), .B(n18899), .ZN(
        P2_U2842) );
  AOI22_X1 U21919 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n18968), .B1(
        P2_EBX_REG_11__SCAN_IN), .B2(n18978), .ZN(n18913) );
  OAI22_X1 U21920 ( .A1(n18902), .A2(n18982), .B1(n18901), .B2(n18958), .ZN(
        n18903) );
  AOI211_X1 U21921 ( .C1(P2_REIP_REG_11__SCAN_IN), .C2(n18993), .A(n19138), 
        .B(n18903), .ZN(n18912) );
  INV_X1 U21922 ( .A(n18989), .ZN(n18904) );
  AOI22_X1 U21923 ( .A1(n18905), .A2(n18984), .B1(n18907), .B2(n18904), .ZN(
        n18911) );
  AOI211_X1 U21924 ( .C1(n18908), .C2(n18907), .A(n19732), .B(n18906), .ZN(
        n18909) );
  INV_X1 U21925 ( .A(n18909), .ZN(n18910) );
  NAND4_X1 U21926 ( .A1(n18913), .A2(n18912), .A3(n18911), .A4(n18910), .ZN(
        P2_U2844) );
  NAND2_X1 U21927 ( .A1(n18954), .A2(n18914), .ZN(n18916) );
  XOR2_X1 U21928 ( .A(n18916), .B(n18915), .Z(n18924) );
  AOI22_X1 U21929 ( .A1(P2_EBX_REG_9__SCAN_IN), .A2(n18978), .B1(n18928), .B2(
        n18917), .ZN(n18918) );
  OAI211_X1 U21930 ( .C1(n11312), .C2(n18938), .A(n18918), .B(n18878), .ZN(
        n18922) );
  OAI22_X1 U21931 ( .A1(n18920), .A2(n18973), .B1(n18958), .B2(n18919), .ZN(
        n18921) );
  AOI211_X1 U21932 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n18968), .A(
        n18922), .B(n18921), .ZN(n18923) );
  OAI21_X1 U21933 ( .B1(n18924), .B2(n19732), .A(n18923), .ZN(P2_U2846) );
  NAND2_X1 U21934 ( .A1(n18954), .A2(n18925), .ZN(n18927) );
  XOR2_X1 U21935 ( .A(n18927), .B(n18926), .Z(n18936) );
  AOI22_X1 U21936 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n18968), .B1(
        n18929), .B2(n18928), .ZN(n18930) );
  OAI211_X1 U21937 ( .C1(n11057), .C2(n18950), .A(n18930), .B(n18878), .ZN(
        n18934) );
  OAI22_X1 U21938 ( .A1(n18932), .A2(n18958), .B1(n18973), .B2(n18931), .ZN(
        n18933) );
  AOI211_X1 U21939 ( .C1(P2_REIP_REG_7__SCAN_IN), .C2(n18993), .A(n18934), .B(
        n18933), .ZN(n18935) );
  OAI21_X1 U21940 ( .B1(n18936), .B2(n19732), .A(n18935), .ZN(P2_U2848) );
  OAI21_X1 U21941 ( .B1(n13686), .B2(n18950), .A(n18878), .ZN(n18940) );
  OAI22_X1 U21942 ( .A1(n19760), .A2(n18938), .B1(n18937), .B2(n18982), .ZN(
        n18939) );
  AOI211_X1 U21943 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n18968), .A(
        n18940), .B(n18939), .ZN(n18947) );
  NOR2_X1 U21944 ( .A1(n18966), .A2(n18941), .ZN(n18943) );
  XNOR2_X1 U21945 ( .A(n18943), .B(n18942), .ZN(n18945) );
  AOI22_X1 U21946 ( .A1(n18945), .A2(n18961), .B1(n18984), .B2(n18944), .ZN(
        n18946) );
  OAI211_X1 U21947 ( .C1(n18958), .C2(n18948), .A(n18947), .B(n18946), .ZN(
        P2_U2849) );
  OAI22_X1 U21948 ( .A1(n18951), .A2(n18950), .B1(n18949), .B2(n18982), .ZN(
        n18952) );
  AOI211_X1 U21949 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n18993), .A(n19138), .B(
        n18952), .ZN(n18963) );
  NAND2_X1 U21950 ( .A1(n18954), .A2(n18953), .ZN(n18955) );
  XNOR2_X1 U21951 ( .A(n18956), .B(n18955), .ZN(n18960) );
  OAI22_X1 U21952 ( .A1(n19020), .A2(n18958), .B1(n18973), .B2(n18957), .ZN(
        n18959) );
  AOI21_X1 U21953 ( .B1(n18961), .B2(n18960), .A(n18959), .ZN(n18962) );
  OAI211_X1 U21954 ( .C1(n18964), .C2(n18990), .A(n18963), .B(n18962), .ZN(
        P2_U2850) );
  NOR2_X1 U21955 ( .A1(n18966), .A2(n18965), .ZN(n18967) );
  XOR2_X1 U21956 ( .A(n19149), .B(n18967), .Z(n18977) );
  AOI21_X1 U21957 ( .B1(P2_REIP_REG_4__SCAN_IN), .B2(n18993), .A(n19138), .ZN(
        n18970) );
  AOI22_X1 U21958 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18968), .B1(
        P2_EBX_REG_4__SCAN_IN), .B2(n18978), .ZN(n18969) );
  OAI211_X1 U21959 ( .C1(n18971), .C2(n18982), .A(n18970), .B(n18969), .ZN(
        n18975) );
  OAI22_X1 U21960 ( .A1(n19023), .A2(n18987), .B1(n18973), .B2(n18972), .ZN(
        n18974) );
  AOI211_X1 U21961 ( .C1(n18979), .C2(n19022), .A(n18975), .B(n18974), .ZN(
        n18976) );
  OAI21_X1 U21962 ( .B1(n19732), .B2(n18977), .A(n18976), .ZN(P2_U2851) );
  AOI22_X1 U21963 ( .A1(n18979), .A2(n19054), .B1(n18978), .B2(
        P2_EBX_REG_0__SCAN_IN), .ZN(n18980) );
  OAI21_X1 U21964 ( .B1(n18982), .B2(n18981), .A(n18980), .ZN(n18983) );
  AOI21_X1 U21965 ( .B1(n18985), .B2(n18984), .A(n18983), .ZN(n18986) );
  OAI21_X1 U21966 ( .B1(n19837), .B2(n18987), .A(n18986), .ZN(n18992) );
  AOI21_X1 U21967 ( .B1(n18990), .B2(n18989), .A(n18988), .ZN(n18991) );
  AOI211_X1 U21968 ( .C1(n18993), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18992), .B(
        n18991), .ZN(n18994) );
  OAI21_X1 U21969 ( .B1(n18996), .B2(n18995), .A(n18994), .ZN(P2_U2855) );
  AOI22_X1 U21970 ( .A1(n18998), .A2(BUF1_REG_31__SCAN_IN), .B1(n19051), .B2(
        n18997), .ZN(n19001) );
  AOI22_X1 U21971 ( .A1(n18999), .A2(BUF2_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n19050), .ZN(n19000) );
  NAND2_X1 U21972 ( .A1(n19001), .A2(n19000), .ZN(P2_U2888) );
  INV_X1 U21973 ( .A(n19057), .ZN(n19010) );
  INV_X1 U21974 ( .A(n19002), .ZN(n19131) );
  AOI22_X1 U21975 ( .A1(n19010), .A2(n19131), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n19050), .ZN(n19003) );
  OAI21_X1 U21976 ( .B1(n19021), .B2(n19004), .A(n19003), .ZN(P2_U2905) );
  INV_X1 U21977 ( .A(n19005), .ZN(n19008) );
  AOI22_X1 U21978 ( .A1(n19010), .A2(n19006), .B1(P2_EAX_REG_8__SCAN_IN), .B2(
        n19050), .ZN(n19007) );
  OAI21_X1 U21979 ( .B1(n19021), .B2(n19008), .A(n19007), .ZN(P2_U2911) );
  AOI22_X1 U21980 ( .A1(n19010), .A2(n19009), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n19050), .ZN(n19019) );
  XNOR2_X1 U21981 ( .A(n19449), .B(n19814), .ZN(n19030) );
  INV_X1 U21982 ( .A(n19820), .ZN(n19011) );
  NAND2_X1 U21983 ( .A1(n19817), .A2(n19011), .ZN(n19014) );
  XNOR2_X1 U21984 ( .A(n19817), .B(n19820), .ZN(n19041) );
  NAND2_X1 U21985 ( .A1(n19824), .A2(n19012), .ZN(n19013) );
  XNOR2_X1 U21986 ( .A(n19824), .B(n19829), .ZN(n19046) );
  NAND2_X1 U21987 ( .A1(n19417), .A2(n19054), .ZN(n19053) );
  NAND2_X1 U21988 ( .A1(n19046), .A2(n19053), .ZN(n19045) );
  NAND2_X1 U21989 ( .A1(n19013), .A2(n19045), .ZN(n19040) );
  NAND2_X1 U21990 ( .A1(n19041), .A2(n19040), .ZN(n19039) );
  NAND2_X1 U21991 ( .A1(n19014), .A2(n19039), .ZN(n19029) );
  NAND2_X1 U21992 ( .A1(n19030), .A2(n19029), .ZN(n19028) );
  OAI21_X1 U21993 ( .B1(n19815), .B2(n19814), .A(n19028), .ZN(n19016) );
  NAND2_X1 U21994 ( .A1(n19016), .A2(n19015), .ZN(n19024) );
  INV_X1 U21995 ( .A(n19023), .ZN(n19017) );
  NAND3_X1 U21996 ( .A1(n19024), .A2(n19017), .A3(n19052), .ZN(n19018) );
  OAI211_X1 U21997 ( .C1(n19021), .C2(n19020), .A(n19019), .B(n19018), .ZN(
        P2_U2914) );
  AOI22_X1 U21998 ( .A1(n19051), .A2(n19022), .B1(n19050), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n19027) );
  XNOR2_X1 U21999 ( .A(n19024), .B(n19023), .ZN(n19025) );
  NAND2_X1 U22000 ( .A1(n19025), .A2(n19052), .ZN(n19026) );
  OAI211_X1 U22001 ( .C1(n19185), .C2(n19057), .A(n19027), .B(n19026), .ZN(
        P2_U2915) );
  OAI21_X1 U22002 ( .B1(n19030), .B2(n19029), .A(n19028), .ZN(n19031) );
  NAND2_X1 U22003 ( .A1(n19031), .A2(n19052), .ZN(n19038) );
  INV_X1 U22004 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19032) );
  OAI22_X1 U22005 ( .A1(n19035), .A2(n19034), .B1(n19033), .B2(n19032), .ZN(
        n19036) );
  INV_X1 U22006 ( .A(n19036), .ZN(n19037) );
  OAI211_X1 U22007 ( .C1(n19181), .C2(n19057), .A(n19038), .B(n19037), .ZN(
        P2_U2916) );
  AOI22_X1 U22008 ( .A1(n19820), .A2(n19051), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19050), .ZN(n19044) );
  OAI21_X1 U22009 ( .B1(n19041), .B2(n19040), .A(n19039), .ZN(n19042) );
  NAND2_X1 U22010 ( .A1(n19042), .A2(n19052), .ZN(n19043) );
  OAI211_X1 U22011 ( .C1(n19175), .C2(n19057), .A(n19044), .B(n19043), .ZN(
        P2_U2917) );
  AOI22_X1 U22012 ( .A1(n19051), .A2(n19829), .B1(n19050), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19049) );
  OAI21_X1 U22013 ( .B1(n19046), .B2(n19053), .A(n19045), .ZN(n19047) );
  NAND2_X1 U22014 ( .A1(n19047), .A2(n19052), .ZN(n19048) );
  OAI211_X1 U22015 ( .C1(n19170), .C2(n19057), .A(n19049), .B(n19048), .ZN(
        P2_U2918) );
  AOI22_X1 U22016 ( .A1(n19051), .A2(n19054), .B1(n19050), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n19056) );
  OAI211_X1 U22017 ( .C1(n19417), .C2(n19054), .A(n19053), .B(n19052), .ZN(
        n19055) );
  OAI211_X1 U22018 ( .C1(n19161), .C2(n19057), .A(n19056), .B(n19055), .ZN(
        P2_U2919) );
  INV_X1 U22019 ( .A(n19058), .ZN(n19060) );
  NAND2_X1 U22020 ( .A1(n19060), .A2(n19059), .ZN(n19063) );
  INV_X1 U22021 ( .A(n19861), .ZN(n19061) );
  NOR2_X1 U22022 ( .A1(n19834), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19087) );
  NOR2_X1 U22023 ( .A1(n19094), .A2(n19064), .ZN(P2_U2920) );
  AND2_X1 U22024 ( .A1(n19100), .A2(n19065), .ZN(n19068) );
  AOI22_X1 U22025 ( .A1(P2_EAX_REG_30__SCAN_IN), .A2(n19068), .B1(n19087), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n19066) );
  OAI21_X1 U22026 ( .B1(n19094), .B2(n19067), .A(n19066), .ZN(P2_U2921) );
  INV_X2 U22027 ( .A(n19094), .ZN(n19126) );
  AOI22_X1 U22028 ( .A1(n19087), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n19069) );
  OAI21_X1 U22029 ( .B1(n19070), .B2(n19098), .A(n19069), .ZN(P2_U2922) );
  AOI22_X1 U22030 ( .A1(n19087), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n19071) );
  OAI21_X1 U22031 ( .B1(n19072), .B2(n19098), .A(n19071), .ZN(P2_U2923) );
  AOI22_X1 U22032 ( .A1(n19087), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n19073) );
  OAI21_X1 U22033 ( .B1(n19074), .B2(n19098), .A(n19073), .ZN(P2_U2924) );
  AOI22_X1 U22034 ( .A1(n19087), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n19075) );
  OAI21_X1 U22035 ( .B1(n19076), .B2(n19098), .A(n19075), .ZN(P2_U2925) );
  AOI22_X1 U22036 ( .A1(n19087), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n19077) );
  OAI21_X1 U22037 ( .B1(n19078), .B2(n19098), .A(n19077), .ZN(P2_U2926) );
  AOI22_X1 U22038 ( .A1(n19087), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n19079) );
  OAI21_X1 U22039 ( .B1(n19080), .B2(n19098), .A(n19079), .ZN(P2_U2927) );
  AOI22_X1 U22040 ( .A1(n19087), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n19081) );
  OAI21_X1 U22041 ( .B1(n19082), .B2(n19098), .A(n19081), .ZN(P2_U2928) );
  AOI22_X1 U22042 ( .A1(n19087), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n19083) );
  OAI21_X1 U22043 ( .B1(n19084), .B2(n19098), .A(n19083), .ZN(P2_U2929) );
  AOI22_X1 U22044 ( .A1(n19087), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n19085) );
  OAI21_X1 U22045 ( .B1(n19086), .B2(n19098), .A(n19085), .ZN(P2_U2930) );
  AOI22_X1 U22046 ( .A1(n19087), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n19088) );
  OAI21_X1 U22047 ( .B1(n19089), .B2(n19098), .A(n19088), .ZN(P2_U2931) );
  AOI22_X1 U22048 ( .A1(n19856), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n19090) );
  OAI21_X1 U22049 ( .B1(n19091), .B2(n19098), .A(n19090), .ZN(P2_U2932) );
  AOI22_X1 U22050 ( .A1(n19856), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n19092) );
  OAI21_X1 U22051 ( .B1(n19093), .B2(n19098), .A(n19092), .ZN(P2_U2933) );
  AOI22_X1 U22052 ( .A1(n19856), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n19095) );
  OAI21_X1 U22053 ( .B1(n19096), .B2(n19098), .A(n19095), .ZN(P2_U2934) );
  AOI22_X1 U22054 ( .A1(n19856), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n19097) );
  OAI21_X1 U22055 ( .B1(n19099), .B2(n19098), .A(n19097), .ZN(P2_U2935) );
  AOI22_X1 U22056 ( .A1(n19856), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19101) );
  OAI21_X1 U22057 ( .B1(n13360), .B2(n19130), .A(n19101), .ZN(P2_U2936) );
  INV_X1 U22058 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19103) );
  AOI22_X1 U22059 ( .A1(n19856), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19102) );
  OAI21_X1 U22060 ( .B1(n19103), .B2(n19130), .A(n19102), .ZN(P2_U2937) );
  AOI22_X1 U22061 ( .A1(n19856), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19104) );
  OAI21_X1 U22062 ( .B1(n19105), .B2(n19130), .A(n19104), .ZN(P2_U2938) );
  AOI22_X1 U22063 ( .A1(n19856), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19106) );
  OAI21_X1 U22064 ( .B1(n19107), .B2(n19130), .A(n19106), .ZN(P2_U2939) );
  AOI22_X1 U22065 ( .A1(n19856), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19108) );
  OAI21_X1 U22066 ( .B1(n19109), .B2(n19130), .A(n19108), .ZN(P2_U2940) );
  AOI22_X1 U22067 ( .A1(n19856), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19110) );
  OAI21_X1 U22068 ( .B1(n19111), .B2(n19130), .A(n19110), .ZN(P2_U2941) );
  AOI22_X1 U22069 ( .A1(n19856), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19112) );
  OAI21_X1 U22070 ( .B1(n19113), .B2(n19130), .A(n19112), .ZN(P2_U2942) );
  AOI22_X1 U22071 ( .A1(n19856), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19114) );
  OAI21_X1 U22072 ( .B1(n19115), .B2(n19130), .A(n19114), .ZN(P2_U2943) );
  AOI22_X1 U22073 ( .A1(n19856), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19116) );
  OAI21_X1 U22074 ( .B1(n19117), .B2(n19130), .A(n19116), .ZN(P2_U2944) );
  AOI22_X1 U22075 ( .A1(n19856), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19118) );
  OAI21_X1 U22076 ( .B1(n19119), .B2(n19130), .A(n19118), .ZN(P2_U2945) );
  INV_X1 U22077 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19121) );
  AOI22_X1 U22078 ( .A1(n19856), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19120) );
  OAI21_X1 U22079 ( .B1(n19121), .B2(n19130), .A(n19120), .ZN(P2_U2946) );
  INV_X1 U22080 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19123) );
  AOI22_X1 U22081 ( .A1(n19856), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19122) );
  OAI21_X1 U22082 ( .B1(n19123), .B2(n19130), .A(n19122), .ZN(P2_U2947) );
  AOI22_X1 U22083 ( .A1(n19856), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19124) );
  OAI21_X1 U22084 ( .B1(n19032), .B2(n19130), .A(n19124), .ZN(P2_U2948) );
  INV_X1 U22085 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n20953) );
  AOI22_X1 U22086 ( .A1(n19856), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19125) );
  OAI21_X1 U22087 ( .B1(n20953), .B2(n19130), .A(n19125), .ZN(P2_U2949) );
  INV_X1 U22088 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19128) );
  AOI22_X1 U22089 ( .A1(n19856), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19127) );
  OAI21_X1 U22090 ( .B1(n19128), .B2(n19130), .A(n19127), .ZN(P2_U2950) );
  AOI22_X1 U22091 ( .A1(n19856), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19129) );
  OAI21_X1 U22092 ( .B1(n11229), .B2(n19130), .A(n19129), .ZN(P2_U2951) );
  AOI22_X1 U22093 ( .A1(n19134), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_30__SCAN_IN), .B2(n13451), .ZN(n19133) );
  NAND2_X1 U22094 ( .A1(n19132), .A2(n19131), .ZN(n19135) );
  NAND2_X1 U22095 ( .A1(n19133), .A2(n19135), .ZN(P2_U2966) );
  AOI22_X1 U22096 ( .A1(n19134), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_14__SCAN_IN), .B2(n13451), .ZN(n19136) );
  NAND2_X1 U22097 ( .A1(n19136), .A2(n19135), .ZN(P2_U2981) );
  AOI22_X1 U22098 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19138), .B1(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n19137), .ZN(n19148) );
  INV_X1 U22099 ( .A(n19139), .ZN(n19143) );
  OAI22_X1 U22100 ( .A1(n19143), .A2(n19142), .B1(n19141), .B2(n19140), .ZN(
        n19144) );
  AOI21_X1 U22101 ( .B1(n19146), .B2(n19145), .A(n19144), .ZN(n19147) );
  OAI211_X1 U22102 ( .C1(n19150), .C2(n19149), .A(n19148), .B(n19147), .ZN(
        P2_U3010) );
  INV_X1 U22103 ( .A(n19232), .ZN(n19151) );
  NAND3_X1 U22104 ( .A1(n19159), .A2(n19813), .A3(n19151), .ZN(n19152) );
  NAND2_X1 U22105 ( .A1(n19813), .A2(n19626), .ZN(n19808) );
  NAND2_X1 U22106 ( .A1(n19152), .A2(n19808), .ZN(n19162) );
  NOR2_X1 U22107 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19236) );
  NAND2_X1 U22108 ( .A1(n19236), .A2(n19831), .ZN(n19211) );
  NOR2_X1 U22109 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19211), .ZN(
        n19200) );
  INV_X1 U22110 ( .A(n19200), .ZN(n19153) );
  AND2_X1 U22111 ( .A1(n19667), .A2(n19153), .ZN(n19165) );
  INV_X1 U22112 ( .A(n19154), .ZN(n19163) );
  AOI211_X1 U22113 ( .C1(n19163), .C2(n20990), .A(n19200), .B(n19813), .ZN(
        n19155) );
  AOI22_X1 U22114 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19203), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n9822), .ZN(n19680) );
  NOR2_X2 U22115 ( .A1(n19160), .A2(n19184), .ZN(n19668) );
  AOI22_X1 U22116 ( .A1(n19625), .A2(n19722), .B1(n19668), .B2(n19200), .ZN(
        n19168) );
  NOR2_X2 U22117 ( .A1(n19161), .A2(n19585), .ZN(n19669) );
  INV_X1 U22118 ( .A(n19162), .ZN(n19166) );
  OAI21_X1 U22119 ( .B1(n19163), .B2(n19200), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19164) );
  AOI22_X1 U22120 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n9822), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19203), .ZN(n19638) );
  AOI22_X1 U22121 ( .A1(n19669), .A2(n19204), .B1(n19232), .B2(n19677), .ZN(
        n19167) );
  OAI211_X1 U22122 ( .C1(n19208), .C2(n11284), .A(n19168), .B(n19167), .ZN(
        P2_U3048) );
  AOI22_X1 U22123 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n9822), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19203), .ZN(n19686) );
  INV_X1 U22124 ( .A(n19686), .ZN(n19593) );
  AOI22_X1 U22125 ( .A1(n19593), .A2(n19722), .B1(n19681), .B2(n19200), .ZN(
        n19172) );
  NOR2_X2 U22126 ( .A1(n19170), .A2(n19585), .ZN(n19682) );
  OAI22_X2 U22127 ( .A1(n15341), .A2(n19202), .B1(n15343), .B2(n19195), .ZN(
        n19683) );
  AOI22_X1 U22128 ( .A1(n19682), .A2(n19204), .B1(n19232), .B2(n19683), .ZN(
        n19171) );
  OAI211_X1 U22129 ( .C1(n19208), .C2(n19173), .A(n19172), .B(n19171), .ZN(
        P2_U3049) );
  AOI22_X1 U22130 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n9822), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19203), .ZN(n19692) );
  INV_X1 U22131 ( .A(n19692), .ZN(n19597) );
  NOR2_X2 U22132 ( .A1(n19174), .A2(n19184), .ZN(n19687) );
  AOI22_X1 U22133 ( .A1(n19597), .A2(n19722), .B1(n19687), .B2(n19200), .ZN(
        n19177) );
  NOR2_X2 U22134 ( .A1(n19175), .A2(n19585), .ZN(n19688) );
  AOI22_X1 U22135 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n9822), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19203), .ZN(n19600) );
  AOI22_X1 U22136 ( .A1(n19688), .A2(n19204), .B1(n19232), .B2(n19689), .ZN(
        n19176) );
  OAI211_X1 U22137 ( .C1(n19208), .C2(n11920), .A(n19177), .B(n19176), .ZN(
        P2_U3050) );
  OAI22_X2 U22138 ( .A1(n19179), .A2(n19202), .B1(n19178), .B2(n19195), .ZN(
        n19643) );
  AOI22_X1 U22139 ( .A1(n19643), .A2(n19722), .B1(n19693), .B2(n19200), .ZN(
        n19183) );
  NOR2_X2 U22140 ( .A1(n19181), .A2(n19585), .ZN(n19694) );
  AOI22_X1 U22141 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n9822), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19203), .ZN(n19646) );
  INV_X1 U22142 ( .A(n19646), .ZN(n19695) );
  AOI22_X1 U22143 ( .A1(n19694), .A2(n19204), .B1(n19232), .B2(n19695), .ZN(
        n19182) );
  OAI211_X1 U22144 ( .C1(n19208), .C2(n11939), .A(n19183), .B(n19182), .ZN(
        P2_U3051) );
  AOI22_X1 U22145 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19203), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n9822), .ZN(n19704) );
  INV_X1 U22146 ( .A(n19704), .ZN(n19648) );
  NOR2_X2 U22147 ( .A1(n10441), .A2(n19184), .ZN(n19699) );
  AOI22_X1 U22148 ( .A1(n19648), .A2(n19722), .B1(n19699), .B2(n19200), .ZN(
        n19187) );
  NOR2_X2 U22149 ( .A1(n19185), .A2(n19585), .ZN(n19700) );
  OAI22_X2 U22150 ( .A1(n15318), .A2(n19202), .B1(n15319), .B2(n19195), .ZN(
        n19701) );
  AOI22_X1 U22151 ( .A1(n19700), .A2(n19204), .B1(n19232), .B2(n19701), .ZN(
        n19186) );
  OAI211_X1 U22152 ( .C1(n19208), .C2(n11368), .A(n19187), .B(n19186), .ZN(
        P2_U3052) );
  AOI22_X1 U22153 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19203), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n9822), .ZN(n19710) );
  INV_X1 U22154 ( .A(n19710), .ZN(n19605) );
  AOI22_X1 U22155 ( .A1(n19605), .A2(n19722), .B1(n19705), .B2(n19200), .ZN(
        n19190) );
  NOR2_X2 U22156 ( .A1(n19188), .A2(n19585), .ZN(n19706) );
  OAI22_X2 U22157 ( .A1(n15308), .A2(n19202), .B1(n15309), .B2(n19195), .ZN(
        n19707) );
  AOI22_X1 U22158 ( .A1(n19706), .A2(n19204), .B1(n19232), .B2(n19707), .ZN(
        n19189) );
  OAI211_X1 U22159 ( .C1(n19208), .C2(n13679), .A(n19190), .B(n19189), .ZN(
        P2_U3053) );
  AOI22_X1 U22160 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n9822), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19203), .ZN(n19716) );
  INV_X1 U22161 ( .A(n19716), .ZN(n19609) );
  AND2_X1 U22162 ( .A1(n10425), .A2(n19198), .ZN(n19711) );
  AOI22_X1 U22163 ( .A1(n19609), .A2(n19722), .B1(n19711), .B2(n19200), .ZN(
        n19193) );
  NOR2_X2 U22164 ( .A1(n19191), .A2(n19585), .ZN(n19712) );
  AOI22_X1 U22165 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n9822), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19203), .ZN(n19612) );
  AOI22_X1 U22166 ( .A1(n19712), .A2(n19204), .B1(n19232), .B2(n19713), .ZN(
        n19192) );
  OAI211_X1 U22167 ( .C1(n19208), .C2(n19194), .A(n19193), .B(n19192), .ZN(
        P2_U3054) );
  AND2_X1 U22168 ( .A1(n19199), .A2(n19198), .ZN(n19717) );
  AOI22_X1 U22169 ( .A1(n19615), .A2(n19722), .B1(n19717), .B2(n19200), .ZN(
        n19206) );
  NOR2_X2 U22170 ( .A1(n19201), .A2(n19585), .ZN(n19719) );
  AOI22_X1 U22171 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19203), .B1(
        BUF1_REG_23__SCAN_IN), .B2(n9822), .ZN(n19620) );
  AOI22_X1 U22172 ( .A1(n19719), .A2(n19204), .B1(n19232), .B2(n19721), .ZN(
        n19205) );
  OAI211_X1 U22173 ( .C1(n19208), .C2(n19207), .A(n19206), .B(n19205), .ZN(
        P2_U3055) );
  INV_X1 U22174 ( .A(n19460), .ZN(n19209) );
  INV_X1 U22175 ( .A(n19728), .ZN(n19581) );
  INV_X1 U22176 ( .A(n19236), .ZN(n19264) );
  NOR2_X1 U22177 ( .A1(n19577), .A2(n19264), .ZN(n19230) );
  NOR3_X1 U22178 ( .A1(n19210), .A2(n19230), .A3(n21095), .ZN(n19212) );
  AOI211_X2 U22179 ( .C1(n19211), .C2(n21095), .A(n19581), .B(n19212), .ZN(
        n19231) );
  AOI22_X1 U22180 ( .A1(n19231), .A2(n19669), .B1(n19668), .B2(n19230), .ZN(
        n19217) );
  NAND2_X1 U22181 ( .A1(n19449), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19385) );
  OAI21_X1 U22182 ( .B1(n19385), .B2(n19460), .A(n19211), .ZN(n19215) );
  INV_X1 U22183 ( .A(n19230), .ZN(n19213) );
  AOI211_X1 U22184 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19213), .A(n19585), 
        .B(n19212), .ZN(n19214) );
  NAND2_X1 U22185 ( .A1(n19215), .A2(n19214), .ZN(n19233) );
  AOI22_X1 U22186 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19233), .B1(
        n19232), .B2(n19625), .ZN(n19216) );
  OAI211_X1 U22187 ( .C1(n19638), .C2(n19263), .A(n19217), .B(n19216), .ZN(
        P2_U3056) );
  INV_X1 U22188 ( .A(n19683), .ZN(n19596) );
  AOI22_X1 U22189 ( .A1(n19231), .A2(n19682), .B1(n19681), .B2(n19230), .ZN(
        n19219) );
  AOI22_X1 U22190 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19233), .B1(
        n19232), .B2(n19593), .ZN(n19218) );
  OAI211_X1 U22191 ( .C1(n19596), .C2(n19263), .A(n19219), .B(n19218), .ZN(
        P2_U3057) );
  AOI22_X1 U22192 ( .A1(n19231), .A2(n19688), .B1(n19687), .B2(n19230), .ZN(
        n19221) );
  AOI22_X1 U22193 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19233), .B1(
        n19232), .B2(n19597), .ZN(n19220) );
  OAI211_X1 U22194 ( .C1(n19600), .C2(n19263), .A(n19221), .B(n19220), .ZN(
        P2_U3058) );
  AOI22_X1 U22195 ( .A1(n19231), .A2(n19694), .B1(n19693), .B2(n19230), .ZN(
        n19223) );
  AOI22_X1 U22196 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19233), .B1(
        n19232), .B2(n19643), .ZN(n19222) );
  OAI211_X1 U22197 ( .C1(n19646), .C2(n19263), .A(n19223), .B(n19222), .ZN(
        P2_U3059) );
  AOI22_X1 U22198 ( .A1(n19231), .A2(n19700), .B1(n19699), .B2(n19230), .ZN(
        n19225) );
  AOI22_X1 U22199 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19233), .B1(
        n19232), .B2(n19648), .ZN(n19224) );
  OAI211_X1 U22200 ( .C1(n19651), .C2(n19263), .A(n19225), .B(n19224), .ZN(
        P2_U3060) );
  INV_X1 U22201 ( .A(n19707), .ZN(n19608) );
  AOI22_X1 U22202 ( .A1(n19231), .A2(n19706), .B1(n19705), .B2(n19230), .ZN(
        n19227) );
  AOI22_X1 U22203 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19233), .B1(
        n19232), .B2(n19605), .ZN(n19226) );
  OAI211_X1 U22204 ( .C1(n19608), .C2(n19263), .A(n19227), .B(n19226), .ZN(
        P2_U3061) );
  AOI22_X1 U22205 ( .A1(n19231), .A2(n19712), .B1(n19711), .B2(n19230), .ZN(
        n19229) );
  AOI22_X1 U22206 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19233), .B1(
        n19232), .B2(n19609), .ZN(n19228) );
  OAI211_X1 U22207 ( .C1(n19612), .C2(n19263), .A(n19229), .B(n19228), .ZN(
        P2_U3062) );
  AOI22_X1 U22208 ( .A1(n19231), .A2(n19719), .B1(n19717), .B2(n19230), .ZN(
        n19235) );
  AOI22_X1 U22209 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19233), .B1(
        n19232), .B2(n19615), .ZN(n19234) );
  OAI211_X1 U22210 ( .C1(n19620), .C2(n19263), .A(n19235), .B(n19234), .ZN(
        P2_U3063) );
  NOR2_X1 U22211 ( .A1(n19623), .A2(n19264), .ZN(n19258) );
  INV_X1 U22212 ( .A(n19258), .ZN(n19239) );
  AND2_X1 U22213 ( .A1(n19240), .A2(n19239), .ZN(n19237) );
  NAND3_X1 U22214 ( .A1(n19813), .A2(n19236), .A3(n19628), .ZN(n19238) );
  OAI21_X1 U22215 ( .B1(n19237), .B2(n21095), .A(n19238), .ZN(n19259) );
  AOI22_X1 U22216 ( .A1(n19259), .A2(n19669), .B1(n19668), .B2(n19258), .ZN(
        n19245) );
  OAI221_X1 U22217 ( .B1(n19626), .B2(n19263), .C1(n19626), .C2(n19293), .A(
        n19238), .ZN(n19242) );
  OAI21_X1 U22218 ( .B1(n19240), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19239), 
        .ZN(n19241) );
  MUX2_X1 U22219 ( .A(n19242), .B(n19241), .S(n19810), .Z(n19243) );
  NAND2_X1 U22220 ( .A1(n19243), .A2(n19672), .ZN(n19260) );
  AOI22_X1 U22221 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19260), .B1(
        n19281), .B2(n19677), .ZN(n19244) );
  OAI211_X1 U22222 ( .C1(n19680), .C2(n19263), .A(n19245), .B(n19244), .ZN(
        P2_U3064) );
  AOI22_X1 U22223 ( .A1(n19259), .A2(n19682), .B1(n19681), .B2(n19258), .ZN(
        n19247) );
  AOI22_X1 U22224 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19260), .B1(
        n19281), .B2(n19683), .ZN(n19246) );
  OAI211_X1 U22225 ( .C1(n19686), .C2(n19263), .A(n19247), .B(n19246), .ZN(
        P2_U3065) );
  AOI22_X1 U22226 ( .A1(n19259), .A2(n19688), .B1(n19687), .B2(n19258), .ZN(
        n19249) );
  AOI22_X1 U22227 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19260), .B1(
        n19281), .B2(n19689), .ZN(n19248) );
  OAI211_X1 U22228 ( .C1(n19692), .C2(n19263), .A(n19249), .B(n19248), .ZN(
        P2_U3066) );
  AOI22_X1 U22229 ( .A1(n19259), .A2(n19694), .B1(n19693), .B2(n19258), .ZN(
        n19251) );
  AOI22_X1 U22230 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19260), .B1(
        n19281), .B2(n19695), .ZN(n19250) );
  OAI211_X1 U22231 ( .C1(n19698), .C2(n19263), .A(n19251), .B(n19250), .ZN(
        P2_U3067) );
  AOI22_X1 U22232 ( .A1(n19259), .A2(n19700), .B1(n19699), .B2(n19258), .ZN(
        n19253) );
  AOI22_X1 U22233 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19260), .B1(
        n19281), .B2(n19701), .ZN(n19252) );
  OAI211_X1 U22234 ( .C1(n19704), .C2(n19263), .A(n19253), .B(n19252), .ZN(
        P2_U3068) );
  AOI22_X1 U22235 ( .A1(n19259), .A2(n19706), .B1(n19705), .B2(n19258), .ZN(
        n19255) );
  AOI22_X1 U22236 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19260), .B1(
        n19281), .B2(n19707), .ZN(n19254) );
  OAI211_X1 U22237 ( .C1(n19710), .C2(n19263), .A(n19255), .B(n19254), .ZN(
        P2_U3069) );
  AOI22_X1 U22238 ( .A1(n19259), .A2(n19712), .B1(n19711), .B2(n19258), .ZN(
        n19257) );
  AOI22_X1 U22239 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19260), .B1(
        n19281), .B2(n19713), .ZN(n19256) );
  OAI211_X1 U22240 ( .C1(n19716), .C2(n19263), .A(n19257), .B(n19256), .ZN(
        P2_U3070) );
  INV_X1 U22241 ( .A(n19615), .ZN(n19727) );
  AOI22_X1 U22242 ( .A1(n19259), .A2(n19719), .B1(n19717), .B2(n19258), .ZN(
        n19262) );
  AOI22_X1 U22243 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19260), .B1(
        n19281), .B2(n19721), .ZN(n19261) );
  OAI211_X1 U22244 ( .C1(n19727), .C2(n19263), .A(n19262), .B(n19261), .ZN(
        P2_U3071) );
  INV_X1 U22245 ( .A(n19522), .ZN(n19517) );
  NOR2_X1 U22246 ( .A1(n19387), .A2(n19264), .ZN(n19288) );
  AOI22_X1 U22247 ( .A1(n19677), .A2(n19319), .B1(n19288), .B2(n19668), .ZN(
        n19274) );
  OAI21_X1 U22248 ( .B1(n19385), .B2(n19522), .A(n19813), .ZN(n19272) );
  NOR2_X1 U22249 ( .A1(n19831), .A2(n19264), .ZN(n19268) );
  NAND2_X1 U22250 ( .A1(n19269), .A2(n20990), .ZN(n19266) );
  INV_X1 U22251 ( .A(n19288), .ZN(n19265) );
  NAND3_X1 U22252 ( .A1(n19266), .A2(n19810), .A3(n19265), .ZN(n19267) );
  OAI211_X1 U22253 ( .C1(n19272), .C2(n19268), .A(n19672), .B(n19267), .ZN(
        n19290) );
  INV_X1 U22254 ( .A(n19268), .ZN(n19271) );
  OAI21_X1 U22255 ( .B1(n19269), .B2(n19288), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19270) );
  OAI21_X1 U22256 ( .B1(n19272), .B2(n19271), .A(n19270), .ZN(n19289) );
  AOI22_X1 U22257 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19290), .B1(
        n19669), .B2(n19289), .ZN(n19273) );
  OAI211_X1 U22258 ( .C1(n19680), .C2(n19293), .A(n19274), .B(n19273), .ZN(
        P2_U3072) );
  AOI22_X1 U22259 ( .A1(n19683), .A2(n19319), .B1(n19288), .B2(n19681), .ZN(
        n19276) );
  AOI22_X1 U22260 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19290), .B1(
        n19682), .B2(n19289), .ZN(n19275) );
  OAI211_X1 U22261 ( .C1(n19686), .C2(n19293), .A(n19276), .B(n19275), .ZN(
        P2_U3073) );
  AOI22_X1 U22262 ( .A1(n19597), .A2(n19281), .B1(n19288), .B2(n19687), .ZN(
        n19278) );
  AOI22_X1 U22263 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19290), .B1(
        n19688), .B2(n19289), .ZN(n19277) );
  OAI211_X1 U22264 ( .C1(n19600), .C2(n19316), .A(n19278), .B(n19277), .ZN(
        P2_U3074) );
  AOI22_X1 U22265 ( .A1(n19643), .A2(n19281), .B1(n19288), .B2(n19693), .ZN(
        n19280) );
  AOI22_X1 U22266 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19290), .B1(
        n19694), .B2(n19289), .ZN(n19279) );
  OAI211_X1 U22267 ( .C1(n19646), .C2(n19316), .A(n19280), .B(n19279), .ZN(
        P2_U3075) );
  AOI22_X1 U22268 ( .A1(n19648), .A2(n19281), .B1(n19288), .B2(n19699), .ZN(
        n19283) );
  AOI22_X1 U22269 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19290), .B1(
        n19700), .B2(n19289), .ZN(n19282) );
  OAI211_X1 U22270 ( .C1(n19651), .C2(n19316), .A(n19283), .B(n19282), .ZN(
        P2_U3076) );
  AOI22_X1 U22271 ( .A1(n19707), .A2(n19319), .B1(n19288), .B2(n19705), .ZN(
        n19285) );
  AOI22_X1 U22272 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19290), .B1(
        n19706), .B2(n19289), .ZN(n19284) );
  OAI211_X1 U22273 ( .C1(n19710), .C2(n19293), .A(n19285), .B(n19284), .ZN(
        P2_U3077) );
  AOI22_X1 U22274 ( .A1(n19713), .A2(n19319), .B1(n19288), .B2(n19711), .ZN(
        n19287) );
  AOI22_X1 U22275 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19290), .B1(
        n19712), .B2(n19289), .ZN(n19286) );
  OAI211_X1 U22276 ( .C1(n19716), .C2(n19293), .A(n19287), .B(n19286), .ZN(
        P2_U3078) );
  AOI22_X1 U22277 ( .A1(n19721), .A2(n19319), .B1(n19288), .B2(n19717), .ZN(
        n19292) );
  AOI22_X1 U22278 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19290), .B1(
        n19719), .B2(n19289), .ZN(n19291) );
  OAI211_X1 U22279 ( .C1(n19727), .C2(n19293), .A(n19292), .B(n19291), .ZN(
        P2_U3079) );
  NOR2_X1 U22280 ( .A1(n19294), .A2(n19628), .ZN(n19543) );
  NAND2_X1 U22281 ( .A1(n19543), .A2(n11933), .ZN(n19300) );
  NOR2_X1 U22282 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19822), .ZN(
        n19357) );
  NAND2_X1 U22283 ( .A1(n19357), .A2(n19831), .ZN(n19331) );
  NOR2_X1 U22284 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19331), .ZN(
        n19317) );
  OAI21_X1 U22285 ( .B1(n10603), .B2(n19317), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19295) );
  OAI21_X1 U22286 ( .B1(n19300), .B2(n19810), .A(n19295), .ZN(n19318) );
  AOI22_X1 U22287 ( .A1(n19318), .A2(n19669), .B1(n19668), .B2(n19317), .ZN(
        n19303) );
  OAI21_X1 U22288 ( .B1(n19319), .B2(n19351), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19299) );
  AOI211_X1 U22289 ( .C1(n19300), .C2(n19299), .A(n19585), .B(n19298), .ZN(
        n19301) );
  AOI22_X1 U22290 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19320), .B1(
        n19351), .B2(n19677), .ZN(n19302) );
  OAI211_X1 U22291 ( .C1(n19680), .C2(n19316), .A(n19303), .B(n19302), .ZN(
        P2_U3080) );
  AOI22_X1 U22292 ( .A1(n19318), .A2(n19682), .B1(n19681), .B2(n19317), .ZN(
        n19305) );
  AOI22_X1 U22293 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19320), .B1(
        n19351), .B2(n19683), .ZN(n19304) );
  OAI211_X1 U22294 ( .C1(n19686), .C2(n19316), .A(n19305), .B(n19304), .ZN(
        P2_U3081) );
  AOI22_X1 U22295 ( .A1(n19318), .A2(n19688), .B1(n19687), .B2(n19317), .ZN(
        n19307) );
  AOI22_X1 U22296 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19320), .B1(
        n19351), .B2(n19689), .ZN(n19306) );
  OAI211_X1 U22297 ( .C1(n19692), .C2(n19316), .A(n19307), .B(n19306), .ZN(
        P2_U3082) );
  AOI22_X1 U22298 ( .A1(n19318), .A2(n19694), .B1(n19693), .B2(n19317), .ZN(
        n19309) );
  AOI22_X1 U22299 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19320), .B1(
        n19319), .B2(n19643), .ZN(n19308) );
  OAI211_X1 U22300 ( .C1(n19646), .C2(n19297), .A(n19309), .B(n19308), .ZN(
        P2_U3083) );
  AOI22_X1 U22301 ( .A1(n19318), .A2(n19700), .B1(n19699), .B2(n19317), .ZN(
        n19311) );
  AOI22_X1 U22302 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19320), .B1(
        n19319), .B2(n19648), .ZN(n19310) );
  OAI211_X1 U22303 ( .C1(n19651), .C2(n19297), .A(n19311), .B(n19310), .ZN(
        P2_U3084) );
  AOI22_X1 U22304 ( .A1(n19318), .A2(n19706), .B1(n19705), .B2(n19317), .ZN(
        n19313) );
  AOI22_X1 U22305 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19320), .B1(
        n19319), .B2(n19605), .ZN(n19312) );
  OAI211_X1 U22306 ( .C1(n19608), .C2(n19297), .A(n19313), .B(n19312), .ZN(
        P2_U3085) );
  AOI22_X1 U22307 ( .A1(n19318), .A2(n19712), .B1(n19711), .B2(n19317), .ZN(
        n19315) );
  AOI22_X1 U22308 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19320), .B1(
        n19351), .B2(n19713), .ZN(n19314) );
  OAI211_X1 U22309 ( .C1(n19716), .C2(n19316), .A(n19315), .B(n19314), .ZN(
        P2_U3086) );
  AOI22_X1 U22310 ( .A1(n19318), .A2(n19719), .B1(n19717), .B2(n19317), .ZN(
        n19322) );
  AOI22_X1 U22311 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19320), .B1(
        n19319), .B2(n19615), .ZN(n19321) );
  OAI211_X1 U22312 ( .C1(n19620), .C2(n19297), .A(n19322), .B(n19321), .ZN(
        P2_U3087) );
  OR2_X1 U22313 ( .A1(n19385), .A2(n19575), .ZN(n19323) );
  NAND2_X1 U22314 ( .A1(n19323), .A2(n19813), .ZN(n19332) );
  INV_X1 U22315 ( .A(n19331), .ZN(n19324) );
  OR2_X1 U22316 ( .A1(n19332), .A2(n19324), .ZN(n19328) );
  INV_X1 U22317 ( .A(n19357), .ZN(n19386) );
  NOR2_X1 U22318 ( .A1(n19577), .A2(n19386), .ZN(n19350) );
  OR2_X1 U22319 ( .A1(n19350), .A2(n19813), .ZN(n19325) );
  AOI21_X1 U22320 ( .B1(n19329), .B2(n20990), .A(n19325), .ZN(n19326) );
  NOR2_X1 U22321 ( .A1(n19585), .A2(n19326), .ZN(n19327) );
  INV_X1 U22322 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n19335) );
  AOI22_X1 U22323 ( .A1(n19625), .A2(n19351), .B1(n19668), .B2(n19350), .ZN(
        n19334) );
  OAI21_X1 U22324 ( .B1(n19329), .B2(n19350), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19330) );
  OAI21_X1 U22325 ( .B1(n19332), .B2(n19331), .A(n19330), .ZN(n19352) );
  AOI22_X1 U22326 ( .A1(n19669), .A2(n19352), .B1(n19381), .B2(n19677), .ZN(
        n19333) );
  OAI211_X1 U22327 ( .C1(n19343), .C2(n19335), .A(n19334), .B(n19333), .ZN(
        P2_U3088) );
  INV_X1 U22328 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n19338) );
  AOI22_X1 U22329 ( .A1(n19683), .A2(n19381), .B1(n19350), .B2(n19681), .ZN(
        n19337) );
  AOI22_X1 U22330 ( .A1(n19682), .A2(n19352), .B1(n19351), .B2(n19593), .ZN(
        n19336) );
  OAI211_X1 U22331 ( .C1(n19343), .C2(n19338), .A(n19337), .B(n19336), .ZN(
        P2_U3089) );
  AOI22_X1 U22332 ( .A1(n19689), .A2(n19381), .B1(n19350), .B2(n19687), .ZN(
        n19340) );
  AOI22_X1 U22333 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19353), .B1(
        n19688), .B2(n19352), .ZN(n19339) );
  OAI211_X1 U22334 ( .C1(n19692), .C2(n19297), .A(n19340), .B(n19339), .ZN(
        P2_U3090) );
  AOI22_X1 U22335 ( .A1(n19643), .A2(n19351), .B1(n19350), .B2(n19693), .ZN(
        n19342) );
  AOI22_X1 U22336 ( .A1(n19694), .A2(n19352), .B1(n19381), .B2(n19695), .ZN(
        n19341) );
  OAI211_X1 U22337 ( .C1(n19343), .C2(n10612), .A(n19342), .B(n19341), .ZN(
        P2_U3091) );
  AOI22_X1 U22338 ( .A1(n19648), .A2(n19351), .B1(n19350), .B2(n19699), .ZN(
        n19345) );
  AOI22_X1 U22339 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19353), .B1(
        n19700), .B2(n19352), .ZN(n19344) );
  OAI211_X1 U22340 ( .C1(n19651), .C2(n19378), .A(n19345), .B(n19344), .ZN(
        P2_U3092) );
  AOI22_X1 U22341 ( .A1(n19707), .A2(n19381), .B1(n19350), .B2(n19705), .ZN(
        n19347) );
  AOI22_X1 U22342 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19353), .B1(
        n19706), .B2(n19352), .ZN(n19346) );
  OAI211_X1 U22343 ( .C1(n19710), .C2(n19297), .A(n19347), .B(n19346), .ZN(
        P2_U3093) );
  AOI22_X1 U22344 ( .A1(n19609), .A2(n19351), .B1(n19350), .B2(n19711), .ZN(
        n19349) );
  AOI22_X1 U22345 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19353), .B1(
        n19712), .B2(n19352), .ZN(n19348) );
  OAI211_X1 U22346 ( .C1(n19612), .C2(n19378), .A(n19349), .B(n19348), .ZN(
        P2_U3094) );
  AOI22_X1 U22347 ( .A1(n19615), .A2(n19351), .B1(n19350), .B2(n19717), .ZN(
        n19355) );
  AOI22_X1 U22348 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19353), .B1(
        n19719), .B2(n19352), .ZN(n19354) );
  OAI211_X1 U22349 ( .C1(n19620), .C2(n19378), .A(n19355), .B(n19354), .ZN(
        P2_U3095) );
  NAND2_X1 U22350 ( .A1(n19628), .A2(n19357), .ZN(n19361) );
  OR2_X1 U22351 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19361), .ZN(n19359) );
  NOR2_X1 U22352 ( .A1(n19623), .A2(n19386), .ZN(n19379) );
  NOR3_X1 U22353 ( .A1(n19358), .A2(n19379), .A3(n21095), .ZN(n19360) );
  AOI21_X1 U22354 ( .B1(n21095), .B2(n19359), .A(n19360), .ZN(n19380) );
  AOI22_X1 U22355 ( .A1(n19380), .A2(n19669), .B1(n19668), .B2(n19379), .ZN(
        n19365) );
  OAI21_X1 U22356 ( .B1(n19381), .B2(n19404), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19362) );
  AOI211_X1 U22357 ( .C1(n19362), .C2(n19361), .A(n19585), .B(n19360), .ZN(
        n19363) );
  AOI22_X1 U22358 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19382), .B1(
        n19381), .B2(n19625), .ZN(n19364) );
  OAI211_X1 U22359 ( .C1(n19638), .C2(n19416), .A(n19365), .B(n19364), .ZN(
        P2_U3096) );
  AOI22_X1 U22360 ( .A1(n19380), .A2(n19682), .B1(n19681), .B2(n19379), .ZN(
        n19367) );
  AOI22_X1 U22361 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19382), .B1(
        n19404), .B2(n19683), .ZN(n19366) );
  OAI211_X1 U22362 ( .C1(n19686), .C2(n19378), .A(n19367), .B(n19366), .ZN(
        P2_U3097) );
  AOI22_X1 U22363 ( .A1(n19380), .A2(n19688), .B1(n19687), .B2(n19379), .ZN(
        n19369) );
  AOI22_X1 U22364 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19382), .B1(
        n19404), .B2(n19689), .ZN(n19368) );
  OAI211_X1 U22365 ( .C1(n19692), .C2(n19378), .A(n19369), .B(n19368), .ZN(
        P2_U3098) );
  AOI22_X1 U22366 ( .A1(n19380), .A2(n19694), .B1(n19693), .B2(n19379), .ZN(
        n19371) );
  AOI22_X1 U22367 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19382), .B1(
        n19381), .B2(n19643), .ZN(n19370) );
  OAI211_X1 U22368 ( .C1(n19646), .C2(n19416), .A(n19371), .B(n19370), .ZN(
        P2_U3099) );
  AOI22_X1 U22369 ( .A1(n19380), .A2(n19700), .B1(n19699), .B2(n19379), .ZN(
        n19373) );
  AOI22_X1 U22370 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19382), .B1(
        n19404), .B2(n19701), .ZN(n19372) );
  OAI211_X1 U22371 ( .C1(n19704), .C2(n19378), .A(n19373), .B(n19372), .ZN(
        P2_U3100) );
  AOI22_X1 U22372 ( .A1(n19380), .A2(n19706), .B1(n19705), .B2(n19379), .ZN(
        n19375) );
  AOI22_X1 U22373 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19382), .B1(
        n19404), .B2(n19707), .ZN(n19374) );
  OAI211_X1 U22374 ( .C1(n19710), .C2(n19378), .A(n19375), .B(n19374), .ZN(
        P2_U3101) );
  AOI22_X1 U22375 ( .A1(n19380), .A2(n19712), .B1(n19711), .B2(n19379), .ZN(
        n19377) );
  AOI22_X1 U22376 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19382), .B1(
        n19404), .B2(n19713), .ZN(n19376) );
  OAI211_X1 U22377 ( .C1(n19716), .C2(n19378), .A(n19377), .B(n19376), .ZN(
        P2_U3102) );
  AOI22_X1 U22378 ( .A1(n19380), .A2(n19719), .B1(n19717), .B2(n19379), .ZN(
        n19384) );
  AOI22_X1 U22379 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19382), .B1(
        n19381), .B2(n19615), .ZN(n19383) );
  OAI211_X1 U22380 ( .C1(n19620), .C2(n19416), .A(n19384), .B(n19383), .ZN(
        P2_U3103) );
  NOR2_X1 U22381 ( .A1(n19385), .A2(n19621), .ZN(n19812) );
  NOR2_X1 U22382 ( .A1(n19831), .A2(n19386), .ZN(n19391) );
  OAI21_X1 U22383 ( .B1(n19812), .B2(n19391), .A(n19672), .ZN(n19390) );
  NOR2_X1 U22384 ( .A1(n19387), .A2(n19386), .ZN(n19424) );
  OR3_X1 U22385 ( .A1(n19388), .A2(n19424), .A3(n21095), .ZN(n19394) );
  OAI21_X1 U22386 ( .B1(n19424), .B2(n20990), .A(n19394), .ZN(n19389) );
  INV_X1 U22387 ( .A(n19413), .ZN(n19407) );
  INV_X1 U22388 ( .A(n19391), .ZN(n19392) );
  OAI21_X1 U22389 ( .B1(n19392), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n21095), 
        .ZN(n19393) );
  AND2_X1 U22390 ( .A1(n19394), .A2(n19393), .ZN(n19412) );
  AOI22_X1 U22391 ( .A1(n19412), .A2(n19669), .B1(n19424), .B2(n19668), .ZN(
        n19397) );
  AOI22_X1 U22392 ( .A1(n19444), .A2(n19677), .B1(n19404), .B2(n19625), .ZN(
        n19396) );
  OAI211_X1 U22393 ( .C1(n19407), .C2(n21089), .A(n19397), .B(n19396), .ZN(
        P2_U3104) );
  AOI22_X1 U22394 ( .A1(n19412), .A2(n19682), .B1(n19424), .B2(n19681), .ZN(
        n19399) );
  AOI22_X1 U22395 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19413), .B1(
        n19404), .B2(n19593), .ZN(n19398) );
  OAI211_X1 U22396 ( .C1(n19596), .C2(n19440), .A(n19399), .B(n19398), .ZN(
        P2_U3105) );
  AOI22_X1 U22397 ( .A1(n19412), .A2(n19688), .B1(n19424), .B2(n19687), .ZN(
        n19401) );
  AOI22_X1 U22398 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19413), .B1(
        n19404), .B2(n19597), .ZN(n19400) );
  OAI211_X1 U22399 ( .C1(n19600), .C2(n19440), .A(n19401), .B(n19400), .ZN(
        P2_U3106) );
  AOI22_X1 U22400 ( .A1(n19412), .A2(n19694), .B1(n19424), .B2(n19693), .ZN(
        n19403) );
  AOI22_X1 U22401 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19413), .B1(
        n19444), .B2(n19695), .ZN(n19402) );
  OAI211_X1 U22402 ( .C1(n19698), .C2(n19416), .A(n19403), .B(n19402), .ZN(
        P2_U3107) );
  AOI22_X1 U22403 ( .A1(n19412), .A2(n19700), .B1(n19424), .B2(n19699), .ZN(
        n19406) );
  AOI22_X1 U22404 ( .A1(n19444), .A2(n19701), .B1(n19404), .B2(n19648), .ZN(
        n19405) );
  OAI211_X1 U22405 ( .C1(n19407), .C2(n10721), .A(n19406), .B(n19405), .ZN(
        P2_U3108) );
  AOI22_X1 U22406 ( .A1(n19412), .A2(n19706), .B1(n19424), .B2(n19705), .ZN(
        n19409) );
  AOI22_X1 U22407 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19413), .B1(
        n19444), .B2(n19707), .ZN(n19408) );
  OAI211_X1 U22408 ( .C1(n19710), .C2(n19416), .A(n19409), .B(n19408), .ZN(
        P2_U3109) );
  AOI22_X1 U22409 ( .A1(n19412), .A2(n19712), .B1(n19424), .B2(n19711), .ZN(
        n19411) );
  AOI22_X1 U22410 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19413), .B1(
        n19444), .B2(n19713), .ZN(n19410) );
  OAI211_X1 U22411 ( .C1(n19716), .C2(n19416), .A(n19411), .B(n19410), .ZN(
        P2_U3110) );
  AOI22_X1 U22412 ( .A1(n19412), .A2(n19719), .B1(n19424), .B2(n19717), .ZN(
        n19415) );
  AOI22_X1 U22413 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19413), .B1(
        n19444), .B2(n19721), .ZN(n19414) );
  OAI211_X1 U22414 ( .C1(n19727), .C2(n19416), .A(n19415), .B(n19414), .ZN(
        P2_U3111) );
  NOR2_X1 U22415 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n11933), .ZN(
        n19513) );
  NAND2_X1 U22416 ( .A1(n19513), .A2(n19831), .ZN(n19458) );
  NOR2_X1 U22417 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19458), .ZN(
        n19443) );
  AOI22_X1 U22418 ( .A1(n19677), .A2(n19474), .B1(n19668), .B2(n19443), .ZN(
        n19429) );
  NAND3_X1 U22419 ( .A1(n19440), .A2(n19813), .A3(n19418), .ZN(n19419) );
  NAND2_X1 U22420 ( .A1(n19419), .A2(n19808), .ZN(n19423) );
  INV_X1 U22421 ( .A(n19424), .ZN(n19421) );
  OAI21_X1 U22422 ( .B1(n19425), .B2(n21095), .A(n20990), .ZN(n19420) );
  AOI21_X1 U22423 ( .B1(n19423), .B2(n19421), .A(n19420), .ZN(n19422) );
  OAI21_X1 U22424 ( .B1(n19424), .B2(n19443), .A(n19423), .ZN(n19427) );
  OAI21_X1 U22425 ( .B1(n19425), .B2(n19443), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19426) );
  NAND2_X1 U22426 ( .A1(n19427), .A2(n19426), .ZN(n19445) );
  AOI22_X1 U22427 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19446), .B1(
        n19669), .B2(n19445), .ZN(n19428) );
  OAI211_X1 U22428 ( .C1(n19680), .C2(n19440), .A(n19429), .B(n19428), .ZN(
        P2_U3112) );
  AOI22_X1 U22429 ( .A1(n19683), .A2(n19474), .B1(n19681), .B2(n19443), .ZN(
        n19431) );
  AOI22_X1 U22430 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19446), .B1(
        n19445), .B2(n19682), .ZN(n19430) );
  OAI211_X1 U22431 ( .C1(n19686), .C2(n19440), .A(n19431), .B(n19430), .ZN(
        P2_U3113) );
  AOI22_X1 U22432 ( .A1(n19597), .A2(n19444), .B1(n19687), .B2(n19443), .ZN(
        n19433) );
  AOI22_X1 U22433 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19446), .B1(
        n19445), .B2(n19688), .ZN(n19432) );
  OAI211_X1 U22434 ( .C1(n19600), .C2(n19418), .A(n19433), .B(n19432), .ZN(
        P2_U3114) );
  AOI22_X1 U22435 ( .A1(n19643), .A2(n19444), .B1(n19693), .B2(n19443), .ZN(
        n19435) );
  AOI22_X1 U22436 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19446), .B1(
        n19445), .B2(n19694), .ZN(n19434) );
  OAI211_X1 U22437 ( .C1(n19646), .C2(n19418), .A(n19435), .B(n19434), .ZN(
        P2_U3115) );
  AOI22_X1 U22438 ( .A1(n19701), .A2(n19474), .B1(n19699), .B2(n19443), .ZN(
        n19437) );
  AOI22_X1 U22439 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19446), .B1(
        n19445), .B2(n19700), .ZN(n19436) );
  OAI211_X1 U22440 ( .C1(n19704), .C2(n19440), .A(n19437), .B(n19436), .ZN(
        P2_U3116) );
  AOI22_X1 U22441 ( .A1(n19707), .A2(n19474), .B1(n19705), .B2(n19443), .ZN(
        n19439) );
  AOI22_X1 U22442 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19446), .B1(
        n19445), .B2(n19706), .ZN(n19438) );
  OAI211_X1 U22443 ( .C1(n19710), .C2(n19440), .A(n19439), .B(n19438), .ZN(
        P2_U3117) );
  AOI22_X1 U22444 ( .A1(n19609), .A2(n19444), .B1(n19711), .B2(n19443), .ZN(
        n19442) );
  AOI22_X1 U22445 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19446), .B1(
        n19445), .B2(n19712), .ZN(n19441) );
  OAI211_X1 U22446 ( .C1(n19612), .C2(n19418), .A(n19442), .B(n19441), .ZN(
        P2_U3118) );
  AOI22_X1 U22447 ( .A1(n19615), .A2(n19444), .B1(n19717), .B2(n19443), .ZN(
        n19448) );
  AOI22_X1 U22448 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19446), .B1(
        n19445), .B2(n19719), .ZN(n19447) );
  OAI211_X1 U22449 ( .C1(n19620), .C2(n19418), .A(n19448), .B(n19447), .ZN(
        P2_U3119) );
  OR2_X1 U22450 ( .A1(n19449), .A2(n19626), .ZN(n19516) );
  OAI21_X1 U22451 ( .B1(n19516), .B2(n19460), .A(n19813), .ZN(n19459) );
  INV_X1 U22452 ( .A(n19458), .ZN(n19450) );
  OR2_X1 U22453 ( .A1(n19459), .A2(n19450), .ZN(n19455) );
  INV_X1 U22454 ( .A(n19513), .ZN(n19482) );
  NOR2_X1 U22455 ( .A1(n19577), .A2(n19482), .ZN(n19477) );
  INV_X1 U22456 ( .A(n19477), .ZN(n19452) );
  OAI211_X1 U22457 ( .C1(n19451), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19452), 
        .B(n19810), .ZN(n19453) );
  AND2_X1 U22458 ( .A1(n19672), .A2(n19453), .ZN(n19454) );
  AOI22_X1 U22459 ( .A1(n19625), .A2(n19474), .B1(n19668), .B2(n19477), .ZN(
        n19462) );
  OAI21_X1 U22460 ( .B1(n19456), .B2(n19477), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19457) );
  OAI21_X1 U22461 ( .B1(n19459), .B2(n19458), .A(n19457), .ZN(n19478) );
  AOI22_X1 U22462 ( .A1(n19669), .A2(n19478), .B1(n19501), .B2(n19677), .ZN(
        n19461) );
  OAI211_X1 U22463 ( .C1(n19465), .C2(n20926), .A(n19462), .B(n19461), .ZN(
        P2_U3120) );
  AOI22_X1 U22464 ( .A1(n19683), .A2(n19501), .B1(n19681), .B2(n19477), .ZN(
        n19464) );
  AOI22_X1 U22465 ( .A1(n19474), .A2(n19593), .B1(n19682), .B2(n19478), .ZN(
        n19463) );
  OAI211_X1 U22466 ( .C1(n19465), .C2(n20917), .A(n19464), .B(n19463), .ZN(
        P2_U3121) );
  AOI22_X1 U22467 ( .A1(n19597), .A2(n19474), .B1(n19687), .B2(n19477), .ZN(
        n19467) );
  AOI22_X1 U22468 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19479), .B1(
        n19688), .B2(n19478), .ZN(n19466) );
  OAI211_X1 U22469 ( .C1(n19600), .C2(n19510), .A(n19467), .B(n19466), .ZN(
        P2_U3122) );
  AOI22_X1 U22470 ( .A1(n19695), .A2(n19501), .B1(n19693), .B2(n19477), .ZN(
        n19469) );
  AOI22_X1 U22471 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19479), .B1(
        n19694), .B2(n19478), .ZN(n19468) );
  OAI211_X1 U22472 ( .C1(n19698), .C2(n19418), .A(n19469), .B(n19468), .ZN(
        P2_U3123) );
  AOI22_X1 U22473 ( .A1(n19701), .A2(n19501), .B1(n19699), .B2(n19477), .ZN(
        n19471) );
  AOI22_X1 U22474 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19479), .B1(
        n19700), .B2(n19478), .ZN(n19470) );
  OAI211_X1 U22475 ( .C1(n19704), .C2(n19418), .A(n19471), .B(n19470), .ZN(
        P2_U3124) );
  AOI22_X1 U22476 ( .A1(n19605), .A2(n19474), .B1(n19705), .B2(n19477), .ZN(
        n19473) );
  AOI22_X1 U22477 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19479), .B1(
        n19706), .B2(n19478), .ZN(n19472) );
  OAI211_X1 U22478 ( .C1(n19608), .C2(n19510), .A(n19473), .B(n19472), .ZN(
        P2_U3125) );
  AOI22_X1 U22479 ( .A1(n19609), .A2(n19474), .B1(n19711), .B2(n19477), .ZN(
        n19476) );
  AOI22_X1 U22480 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19479), .B1(
        n19712), .B2(n19478), .ZN(n19475) );
  OAI211_X1 U22481 ( .C1(n19612), .C2(n19510), .A(n19476), .B(n19475), .ZN(
        P2_U3126) );
  AOI22_X1 U22482 ( .A1(n19721), .A2(n19501), .B1(n19717), .B2(n19477), .ZN(
        n19481) );
  AOI22_X1 U22483 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19479), .B1(
        n19719), .B2(n19478), .ZN(n19480) );
  OAI211_X1 U22484 ( .C1(n19727), .C2(n19418), .A(n19481), .B(n19480), .ZN(
        P2_U3127) );
  NOR2_X1 U22485 ( .A1(n19623), .A2(n19482), .ZN(n19504) );
  AOI22_X1 U22486 ( .A1(n19625), .A2(n19501), .B1(n19668), .B2(n19504), .ZN(
        n19490) );
  NAND3_X1 U22487 ( .A1(n19542), .A2(n19510), .A3(n19813), .ZN(n19483) );
  NAND2_X1 U22488 ( .A1(n19483), .A2(n19808), .ZN(n19485) );
  NAND2_X1 U22489 ( .A1(n19628), .A2(n19513), .ZN(n19487) );
  NOR2_X1 U22490 ( .A1(n10753), .A2(n19504), .ZN(n19486) );
  AOI22_X1 U22491 ( .A1(n19485), .A2(n19487), .B1(P2_STATE2_REG_2__SCAN_IN), 
        .B2(n19486), .ZN(n19484) );
  OAI211_X1 U22492 ( .C1(n19504), .C2(n20990), .A(n19484), .B(n19672), .ZN(
        n19507) );
  INV_X1 U22493 ( .A(n19485), .ZN(n19488) );
  AOI22_X1 U22494 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19507), .B1(
        n19669), .B2(n19506), .ZN(n19489) );
  OAI211_X1 U22495 ( .C1(n19638), .C2(n19542), .A(n19490), .B(n19489), .ZN(
        P2_U3128) );
  INV_X1 U22496 ( .A(n19542), .ZN(n19505) );
  AOI22_X1 U22497 ( .A1(n19683), .A2(n19505), .B1(n19681), .B2(n19504), .ZN(
        n19492) );
  AOI22_X1 U22498 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19507), .B1(
        n19682), .B2(n19506), .ZN(n19491) );
  OAI211_X1 U22499 ( .C1(n19686), .C2(n19510), .A(n19492), .B(n19491), .ZN(
        P2_U3129) );
  AOI22_X1 U22500 ( .A1(n19689), .A2(n19505), .B1(n19687), .B2(n19504), .ZN(
        n19494) );
  AOI22_X1 U22501 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19507), .B1(
        n19688), .B2(n19506), .ZN(n19493) );
  OAI211_X1 U22502 ( .C1(n19692), .C2(n19510), .A(n19494), .B(n19493), .ZN(
        P2_U3130) );
  AOI22_X1 U22503 ( .A1(n19695), .A2(n19505), .B1(n19693), .B2(n19504), .ZN(
        n19496) );
  AOI22_X1 U22504 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19507), .B1(
        n19694), .B2(n19506), .ZN(n19495) );
  OAI211_X1 U22505 ( .C1(n19698), .C2(n19510), .A(n19496), .B(n19495), .ZN(
        P2_U3131) );
  AOI22_X1 U22506 ( .A1(n19701), .A2(n19505), .B1(n19699), .B2(n19504), .ZN(
        n19498) );
  AOI22_X1 U22507 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19507), .B1(
        n19700), .B2(n19506), .ZN(n19497) );
  OAI211_X1 U22508 ( .C1(n19704), .C2(n19510), .A(n19498), .B(n19497), .ZN(
        P2_U3132) );
  AOI22_X1 U22509 ( .A1(n19605), .A2(n19501), .B1(n19705), .B2(n19504), .ZN(
        n19500) );
  AOI22_X1 U22510 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19507), .B1(
        n19706), .B2(n19506), .ZN(n19499) );
  OAI211_X1 U22511 ( .C1(n19608), .C2(n19542), .A(n19500), .B(n19499), .ZN(
        P2_U3133) );
  AOI22_X1 U22512 ( .A1(n19609), .A2(n19501), .B1(n19711), .B2(n19504), .ZN(
        n19503) );
  AOI22_X1 U22513 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19507), .B1(
        n19712), .B2(n19506), .ZN(n19502) );
  OAI211_X1 U22514 ( .C1(n19612), .C2(n19542), .A(n19503), .B(n19502), .ZN(
        P2_U3134) );
  AOI22_X1 U22515 ( .A1(n19721), .A2(n19505), .B1(n19717), .B2(n19504), .ZN(
        n19509) );
  AOI22_X1 U22516 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19507), .B1(
        n19719), .B2(n19506), .ZN(n19508) );
  OAI211_X1 U22517 ( .C1(n19727), .C2(n19510), .A(n19509), .B(n19508), .ZN(
        P2_U3135) );
  NAND2_X1 U22518 ( .A1(n19511), .A2(n19513), .ZN(n19515) );
  AND2_X1 U22519 ( .A1(n19515), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19512) );
  NAND2_X1 U22520 ( .A1(n10754), .A2(n19512), .ZN(n19520) );
  NAND2_X1 U22521 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19513), .ZN(
        n19519) );
  OAI21_X1 U22522 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19519), .A(n21095), 
        .ZN(n19514) );
  INV_X1 U22523 ( .A(n19515), .ZN(n19537) );
  AOI22_X1 U22524 ( .A1(n19538), .A2(n19669), .B1(n19537), .B2(n19668), .ZN(
        n19524) );
  NOR2_X1 U22525 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20990), .ZN(
        n19838) );
  NAND3_X1 U22526 ( .A1(n19517), .A2(n19675), .A3(n20990), .ZN(n19518) );
  OAI21_X1 U22527 ( .B1(n19838), .B2(n19519), .A(n19518), .ZN(n19521) );
  NAND3_X1 U22528 ( .A1(n19521), .A2(n19672), .A3(n19520), .ZN(n19539) );
  NOR2_X2 U22529 ( .A1(n19576), .A2(n19522), .ZN(n19570) );
  AOI22_X1 U22530 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19539), .B1(
        n19570), .B2(n19677), .ZN(n19523) );
  OAI211_X1 U22531 ( .C1(n19680), .C2(n19542), .A(n19524), .B(n19523), .ZN(
        P2_U3136) );
  AOI22_X1 U22532 ( .A1(n19538), .A2(n19682), .B1(n19537), .B2(n19681), .ZN(
        n19526) );
  AOI22_X1 U22533 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19539), .B1(
        n19570), .B2(n19683), .ZN(n19525) );
  OAI211_X1 U22534 ( .C1(n19686), .C2(n19542), .A(n19526), .B(n19525), .ZN(
        P2_U3137) );
  AOI22_X1 U22535 ( .A1(n19538), .A2(n19688), .B1(n19537), .B2(n19687), .ZN(
        n19528) );
  AOI22_X1 U22536 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19539), .B1(
        n19570), .B2(n19689), .ZN(n19527) );
  OAI211_X1 U22537 ( .C1(n19692), .C2(n19542), .A(n19528), .B(n19527), .ZN(
        P2_U3138) );
  AOI22_X1 U22538 ( .A1(n19538), .A2(n19694), .B1(n19537), .B2(n19693), .ZN(
        n19530) );
  AOI22_X1 U22539 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19539), .B1(
        n19570), .B2(n19695), .ZN(n19529) );
  OAI211_X1 U22540 ( .C1(n19698), .C2(n19542), .A(n19530), .B(n19529), .ZN(
        P2_U3139) );
  AOI22_X1 U22541 ( .A1(n19538), .A2(n19700), .B1(n19537), .B2(n19699), .ZN(
        n19532) );
  AOI22_X1 U22542 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19539), .B1(
        n19570), .B2(n19701), .ZN(n19531) );
  OAI211_X1 U22543 ( .C1(n19704), .C2(n19542), .A(n19532), .B(n19531), .ZN(
        P2_U3140) );
  AOI22_X1 U22544 ( .A1(n19538), .A2(n19706), .B1(n19537), .B2(n19705), .ZN(
        n19534) );
  AOI22_X1 U22545 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19539), .B1(
        n19570), .B2(n19707), .ZN(n19533) );
  OAI211_X1 U22546 ( .C1(n19710), .C2(n19542), .A(n19534), .B(n19533), .ZN(
        P2_U3141) );
  AOI22_X1 U22547 ( .A1(n19538), .A2(n19712), .B1(n19537), .B2(n19711), .ZN(
        n19536) );
  AOI22_X1 U22548 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19539), .B1(
        n19570), .B2(n19713), .ZN(n19535) );
  OAI211_X1 U22549 ( .C1(n19716), .C2(n19542), .A(n19536), .B(n19535), .ZN(
        P2_U3142) );
  AOI22_X1 U22550 ( .A1(n19538), .A2(n19719), .B1(n19537), .B2(n19717), .ZN(
        n19541) );
  AOI22_X1 U22551 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19539), .B1(
        n19570), .B2(n19721), .ZN(n19540) );
  OAI211_X1 U22552 ( .C1(n19727), .C2(n19542), .A(n19541), .B(n19540), .ZN(
        P2_U3143) );
  NOR2_X2 U22553 ( .A1(n19622), .A2(n19575), .ZN(n19616) );
  OAI21_X1 U22554 ( .B1(n19616), .B2(n19570), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19549) );
  NAND2_X1 U22555 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19543), .ZN(
        n19550) );
  NOR2_X1 U22556 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19544) );
  NAND2_X1 U22557 ( .A1(n19665), .A2(n19544), .ZN(n19545) );
  INV_X1 U22558 ( .A(n19545), .ZN(n19568) );
  AND2_X1 U22559 ( .A1(n19545), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19546) );
  NAND2_X1 U22560 ( .A1(n19547), .A2(n19546), .ZN(n19552) );
  OAI211_X1 U22561 ( .C1(n19568), .C2(n20990), .A(n19672), .B(n19552), .ZN(
        n19548) );
  OAI21_X1 U22562 ( .B1(n19550), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n21095), 
        .ZN(n19551) );
  AND2_X1 U22563 ( .A1(n19552), .A2(n19551), .ZN(n19569) );
  AOI22_X1 U22564 ( .A1(n19569), .A2(n19669), .B1(n19568), .B2(n19668), .ZN(
        n19554) );
  AOI22_X1 U22565 ( .A1(n19616), .A2(n19677), .B1(n19570), .B2(n19625), .ZN(
        n19553) );
  OAI211_X1 U22566 ( .C1(n19574), .C2(n19555), .A(n19554), .B(n19553), .ZN(
        P2_U3144) );
  AOI22_X1 U22567 ( .A1(n19569), .A2(n19682), .B1(n19568), .B2(n19681), .ZN(
        n19557) );
  AOI22_X1 U22568 ( .A1(n19616), .A2(n19683), .B1(n19570), .B2(n19593), .ZN(
        n19556) );
  OAI211_X1 U22569 ( .C1(n19574), .C2(n11967), .A(n19557), .B(n19556), .ZN(
        P2_U3145) );
  AOI22_X1 U22570 ( .A1(n19569), .A2(n19688), .B1(n19568), .B2(n19687), .ZN(
        n19559) );
  AOI22_X1 U22571 ( .A1(n19570), .A2(n19597), .B1(n19616), .B2(n19689), .ZN(
        n19558) );
  OAI211_X1 U22572 ( .C1(n19574), .C2(n12011), .A(n19559), .B(n19558), .ZN(
        P2_U3146) );
  AOI22_X1 U22573 ( .A1(n19569), .A2(n19694), .B1(n19568), .B2(n19693), .ZN(
        n19561) );
  AOI22_X1 U22574 ( .A1(n19570), .A2(n19643), .B1(n19616), .B2(n19695), .ZN(
        n19560) );
  OAI211_X1 U22575 ( .C1(n19574), .C2(n11998), .A(n19561), .B(n19560), .ZN(
        P2_U3147) );
  AOI22_X1 U22576 ( .A1(n19569), .A2(n19700), .B1(n19568), .B2(n19699), .ZN(
        n19563) );
  AOI22_X1 U22577 ( .A1(n19616), .A2(n19701), .B1(n19570), .B2(n19648), .ZN(
        n19562) );
  OAI211_X1 U22578 ( .C1(n19574), .C2(n11985), .A(n19563), .B(n19562), .ZN(
        P2_U3148) );
  AOI22_X1 U22579 ( .A1(n19569), .A2(n19706), .B1(n19568), .B2(n19705), .ZN(
        n19565) );
  AOI22_X1 U22580 ( .A1(n19616), .A2(n19707), .B1(n19570), .B2(n19605), .ZN(
        n19564) );
  OAI211_X1 U22581 ( .C1(n19574), .C2(n12027), .A(n19565), .B(n19564), .ZN(
        P2_U3149) );
  AOI22_X1 U22582 ( .A1(n19569), .A2(n19712), .B1(n19568), .B2(n19711), .ZN(
        n19567) );
  AOI22_X1 U22583 ( .A1(n19570), .A2(n19609), .B1(n19616), .B2(n19713), .ZN(
        n19566) );
  OAI211_X1 U22584 ( .C1(n19574), .C2(n12047), .A(n19567), .B(n19566), .ZN(
        P2_U3150) );
  INV_X1 U22585 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n19573) );
  AOI22_X1 U22586 ( .A1(n19569), .A2(n19719), .B1(n19568), .B2(n19717), .ZN(
        n19572) );
  AOI22_X1 U22587 ( .A1(n19570), .A2(n19615), .B1(n19616), .B2(n19721), .ZN(
        n19571) );
  OAI211_X1 U22588 ( .C1(n19574), .C2(n19573), .A(n19572), .B(n19571), .ZN(
        P2_U3151) );
  NAND2_X1 U22589 ( .A1(n19665), .A2(n19831), .ZN(n19582) );
  INV_X1 U22590 ( .A(n19577), .ZN(n19578) );
  NAND2_X1 U22591 ( .A1(n19665), .A2(n19578), .ZN(n19583) );
  AND2_X1 U22592 ( .A1(n19583), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19579) );
  AOI211_X2 U22593 ( .C1(n21095), .C2(n19582), .A(n19581), .B(n19587), .ZN(
        n19614) );
  INV_X1 U22594 ( .A(n19583), .ZN(n19613) );
  AOI22_X1 U22595 ( .A1(n19614), .A2(n19669), .B1(n19668), .B2(n19613), .ZN(
        n19592) );
  INV_X1 U22596 ( .A(n19582), .ZN(n19590) );
  AND2_X1 U22597 ( .A1(n19583), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19584) );
  OR2_X1 U22598 ( .A1(n19585), .A2(n19584), .ZN(n19586) );
  NOR2_X1 U22599 ( .A1(n19587), .A2(n19586), .ZN(n19588) );
  OAI221_X1 U22600 ( .B1(n19590), .B2(n19589), .C1(n19590), .C2(n19675), .A(
        n19588), .ZN(n19617) );
  AOI22_X1 U22601 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19617), .B1(
        n19616), .B2(n19625), .ZN(n19591) );
  OAI211_X1 U22602 ( .C1(n19638), .C2(n19662), .A(n19592), .B(n19591), .ZN(
        P2_U3152) );
  AOI22_X1 U22603 ( .A1(n19614), .A2(n19682), .B1(n19681), .B2(n19613), .ZN(
        n19595) );
  AOI22_X1 U22604 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19617), .B1(
        n19616), .B2(n19593), .ZN(n19594) );
  OAI211_X1 U22605 ( .C1(n19596), .C2(n19662), .A(n19595), .B(n19594), .ZN(
        P2_U3153) );
  AOI22_X1 U22606 ( .A1(n19614), .A2(n19688), .B1(n19687), .B2(n19613), .ZN(
        n19599) );
  AOI22_X1 U22607 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19617), .B1(
        n19616), .B2(n19597), .ZN(n19598) );
  OAI211_X1 U22608 ( .C1(n19600), .C2(n19662), .A(n19599), .B(n19598), .ZN(
        P2_U3154) );
  AOI22_X1 U22609 ( .A1(n19614), .A2(n19694), .B1(n19693), .B2(n19613), .ZN(
        n19602) );
  AOI22_X1 U22610 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19617), .B1(
        n19616), .B2(n19643), .ZN(n19601) );
  OAI211_X1 U22611 ( .C1(n19646), .C2(n19662), .A(n19602), .B(n19601), .ZN(
        P2_U3155) );
  AOI22_X1 U22612 ( .A1(n19614), .A2(n19700), .B1(n19699), .B2(n19613), .ZN(
        n19604) );
  AOI22_X1 U22613 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19617), .B1(
        n19616), .B2(n19648), .ZN(n19603) );
  OAI211_X1 U22614 ( .C1(n19651), .C2(n19662), .A(n19604), .B(n19603), .ZN(
        P2_U3156) );
  AOI22_X1 U22615 ( .A1(n19614), .A2(n19706), .B1(n19705), .B2(n19613), .ZN(
        n19607) );
  AOI22_X1 U22616 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19617), .B1(
        n19616), .B2(n19605), .ZN(n19606) );
  OAI211_X1 U22617 ( .C1(n19608), .C2(n19662), .A(n19607), .B(n19606), .ZN(
        P2_U3157) );
  AOI22_X1 U22618 ( .A1(n19614), .A2(n19712), .B1(n19711), .B2(n19613), .ZN(
        n19611) );
  AOI22_X1 U22619 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19617), .B1(
        n19616), .B2(n19609), .ZN(n19610) );
  OAI211_X1 U22620 ( .C1(n19612), .C2(n19662), .A(n19611), .B(n19610), .ZN(
        P2_U3158) );
  AOI22_X1 U22621 ( .A1(n19614), .A2(n19719), .B1(n19717), .B2(n19613), .ZN(
        n19619) );
  AOI22_X1 U22622 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19617), .B1(
        n19616), .B2(n19615), .ZN(n19618) );
  OAI211_X1 U22623 ( .C1(n19620), .C2(n19662), .A(n19619), .B(n19618), .ZN(
        P2_U3159) );
  INV_X1 U22624 ( .A(n19623), .ZN(n19624) );
  AND2_X1 U22625 ( .A1(n19665), .A2(n19624), .ZN(n19656) );
  AOI22_X1 U22626 ( .A1(n19625), .A2(n19647), .B1(n19656), .B2(n19668), .ZN(
        n19637) );
  NOR2_X1 U22627 ( .A1(n19657), .A2(n19647), .ZN(n19627) );
  OAI21_X1 U22628 ( .B1(n19627), .B2(n19626), .A(n19813), .ZN(n19635) );
  AND2_X1 U22629 ( .A1(n19665), .A2(n19628), .ZN(n19632) );
  INV_X1 U22630 ( .A(n19656), .ZN(n19629) );
  OAI211_X1 U22631 ( .C1(n19630), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19629), 
        .B(n19810), .ZN(n19631) );
  OAI211_X1 U22632 ( .C1(n19635), .C2(n19632), .A(n19672), .B(n19631), .ZN(
        n19659) );
  INV_X1 U22633 ( .A(n19632), .ZN(n19634) );
  OAI21_X1 U22634 ( .B1(n10741), .B2(n19656), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19633) );
  AOI22_X1 U22635 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19659), .B1(
        n19669), .B2(n19658), .ZN(n19636) );
  OAI211_X1 U22636 ( .C1(n19638), .C2(n19726), .A(n19637), .B(n19636), .ZN(
        P2_U3160) );
  AOI22_X1 U22637 ( .A1(n19683), .A2(n19657), .B1(n19656), .B2(n19681), .ZN(
        n19640) );
  AOI22_X1 U22638 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19659), .B1(
        n19682), .B2(n19658), .ZN(n19639) );
  OAI211_X1 U22639 ( .C1(n19686), .C2(n19662), .A(n19640), .B(n19639), .ZN(
        P2_U3161) );
  AOI22_X1 U22640 ( .A1(n19689), .A2(n19657), .B1(n19656), .B2(n19687), .ZN(
        n19642) );
  AOI22_X1 U22641 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19659), .B1(
        n19688), .B2(n19658), .ZN(n19641) );
  OAI211_X1 U22642 ( .C1(n19692), .C2(n19662), .A(n19642), .B(n19641), .ZN(
        P2_U3162) );
  AOI22_X1 U22643 ( .A1(n19643), .A2(n19647), .B1(n19656), .B2(n19693), .ZN(
        n19645) );
  AOI22_X1 U22644 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19659), .B1(
        n19694), .B2(n19658), .ZN(n19644) );
  OAI211_X1 U22645 ( .C1(n19646), .C2(n19726), .A(n19645), .B(n19644), .ZN(
        P2_U3163) );
  AOI22_X1 U22646 ( .A1(n19648), .A2(n19647), .B1(n19656), .B2(n19699), .ZN(
        n19650) );
  AOI22_X1 U22647 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19659), .B1(
        n19700), .B2(n19658), .ZN(n19649) );
  OAI211_X1 U22648 ( .C1(n19651), .C2(n19726), .A(n19650), .B(n19649), .ZN(
        P2_U3164) );
  AOI22_X1 U22649 ( .A1(n19707), .A2(n19657), .B1(n19656), .B2(n19705), .ZN(
        n19653) );
  AOI22_X1 U22650 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19659), .B1(
        n19706), .B2(n19658), .ZN(n19652) );
  OAI211_X1 U22651 ( .C1(n19710), .C2(n19662), .A(n19653), .B(n19652), .ZN(
        P2_U3165) );
  AOI22_X1 U22652 ( .A1(n19713), .A2(n19657), .B1(n19656), .B2(n19711), .ZN(
        n19655) );
  AOI22_X1 U22653 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19659), .B1(
        n19712), .B2(n19658), .ZN(n19654) );
  OAI211_X1 U22654 ( .C1(n19716), .C2(n19662), .A(n19655), .B(n19654), .ZN(
        P2_U3166) );
  AOI22_X1 U22655 ( .A1(n19721), .A2(n19657), .B1(n19656), .B2(n19717), .ZN(
        n19661) );
  AOI22_X1 U22656 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19659), .B1(
        n19719), .B2(n19658), .ZN(n19660) );
  OAI211_X1 U22657 ( .C1(n19727), .C2(n19662), .A(n19661), .B(n19660), .ZN(
        P2_U3167) );
  AND2_X1 U22658 ( .A1(n19667), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19663) );
  NAND2_X1 U22659 ( .A1(n19664), .A2(n19663), .ZN(n19671) );
  NAND2_X1 U22660 ( .A1(n19665), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19670) );
  OAI21_X1 U22661 ( .B1(n19670), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n21095), 
        .ZN(n19666) );
  AND2_X1 U22662 ( .A1(n19671), .A2(n19666), .ZN(n19720) );
  INV_X1 U22663 ( .A(n19667), .ZN(n19718) );
  AOI22_X1 U22664 ( .A1(n19720), .A2(n19669), .B1(n19718), .B2(n19668), .ZN(
        n19679) );
  INV_X1 U22665 ( .A(n19670), .ZN(n19676) );
  OAI211_X1 U22666 ( .C1(n19718), .C2(n20990), .A(n19672), .B(n19671), .ZN(
        n19673) );
  INV_X1 U22667 ( .A(n19673), .ZN(n19674) );
  OAI221_X1 U22668 ( .B1(n19676), .B2(n19811), .C1(n19676), .C2(n19675), .A(
        n19674), .ZN(n19723) );
  AOI22_X1 U22669 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19723), .B1(
        n19722), .B2(n19677), .ZN(n19678) );
  OAI211_X1 U22670 ( .C1(n19680), .C2(n19726), .A(n19679), .B(n19678), .ZN(
        P2_U3168) );
  AOI22_X1 U22671 ( .A1(n19720), .A2(n19682), .B1(n19718), .B2(n19681), .ZN(
        n19685) );
  AOI22_X1 U22672 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19723), .B1(
        n19722), .B2(n19683), .ZN(n19684) );
  OAI211_X1 U22673 ( .C1(n19686), .C2(n19726), .A(n19685), .B(n19684), .ZN(
        P2_U3169) );
  AOI22_X1 U22674 ( .A1(n19720), .A2(n19688), .B1(n19718), .B2(n19687), .ZN(
        n19691) );
  AOI22_X1 U22675 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19723), .B1(
        n19722), .B2(n19689), .ZN(n19690) );
  OAI211_X1 U22676 ( .C1(n19692), .C2(n19726), .A(n19691), .B(n19690), .ZN(
        P2_U3170) );
  AOI22_X1 U22677 ( .A1(n19720), .A2(n19694), .B1(n19718), .B2(n19693), .ZN(
        n19697) );
  AOI22_X1 U22678 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19723), .B1(
        n19722), .B2(n19695), .ZN(n19696) );
  OAI211_X1 U22679 ( .C1(n19698), .C2(n19726), .A(n19697), .B(n19696), .ZN(
        P2_U3171) );
  AOI22_X1 U22680 ( .A1(n19720), .A2(n19700), .B1(n19718), .B2(n19699), .ZN(
        n19703) );
  AOI22_X1 U22681 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19723), .B1(
        n19722), .B2(n19701), .ZN(n19702) );
  OAI211_X1 U22682 ( .C1(n19704), .C2(n19726), .A(n19703), .B(n19702), .ZN(
        P2_U3172) );
  AOI22_X1 U22683 ( .A1(n19720), .A2(n19706), .B1(n19718), .B2(n19705), .ZN(
        n19709) );
  AOI22_X1 U22684 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19723), .B1(
        n19722), .B2(n19707), .ZN(n19708) );
  OAI211_X1 U22685 ( .C1(n19710), .C2(n19726), .A(n19709), .B(n19708), .ZN(
        P2_U3173) );
  AOI22_X1 U22686 ( .A1(n19720), .A2(n19712), .B1(n19718), .B2(n19711), .ZN(
        n19715) );
  AOI22_X1 U22687 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19723), .B1(
        n19722), .B2(n19713), .ZN(n19714) );
  OAI211_X1 U22688 ( .C1(n19716), .C2(n19726), .A(n19715), .B(n19714), .ZN(
        P2_U3174) );
  AOI22_X1 U22689 ( .A1(n19720), .A2(n19719), .B1(n19718), .B2(n19717), .ZN(
        n19725) );
  AOI22_X1 U22690 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19723), .B1(
        n19722), .B2(n19721), .ZN(n19724) );
  OAI211_X1 U22691 ( .C1(n19727), .C2(n19726), .A(n19725), .B(n19724), .ZN(
        P2_U3175) );
  OAI211_X1 U22692 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19858), .A(n19729), 
        .B(n19728), .ZN(n19734) );
  OAI21_X1 U22693 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n19859), .A(n19729), 
        .ZN(n19730) );
  NAND3_X1 U22694 ( .A1(n19731), .A2(P2_STATE2_REG_1__SCAN_IN), .A3(n19730), 
        .ZN(n19733) );
  OAI211_X1 U22695 ( .C1(n19735), .C2(n19734), .A(n19733), .B(n19732), .ZN(
        P2_U3177) );
  AND2_X1 U22696 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19804), .ZN(
        P2_U3179) );
  AND2_X1 U22697 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19804), .ZN(
        P2_U3180) );
  AND2_X1 U22698 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19804), .ZN(
        P2_U3181) );
  AND2_X1 U22699 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19804), .ZN(
        P2_U3182) );
  AND2_X1 U22700 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19804), .ZN(
        P2_U3183) );
  AND2_X1 U22701 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19804), .ZN(
        P2_U3184) );
  AND2_X1 U22702 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19804), .ZN(
        P2_U3185) );
  AND2_X1 U22703 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19804), .ZN(
        P2_U3186) );
  AND2_X1 U22704 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19804), .ZN(
        P2_U3187) );
  AND2_X1 U22705 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19804), .ZN(
        P2_U3188) );
  NOR2_X1 U22706 ( .A1(n21037), .A2(n19807), .ZN(P2_U3189) );
  AND2_X1 U22707 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19804), .ZN(
        P2_U3190) );
  AND2_X1 U22708 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19804), .ZN(
        P2_U3191) );
  AND2_X1 U22709 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19804), .ZN(
        P2_U3192) );
  AND2_X1 U22710 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19804), .ZN(
        P2_U3193) );
  AND2_X1 U22711 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19804), .ZN(
        P2_U3194) );
  AND2_X1 U22712 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19804), .ZN(
        P2_U3195) );
  AND2_X1 U22713 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19804), .ZN(
        P2_U3196) );
  AND2_X1 U22714 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19804), .ZN(
        P2_U3197) );
  AND2_X1 U22715 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19804), .ZN(
        P2_U3198) );
  AND2_X1 U22716 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19804), .ZN(
        P2_U3199) );
  AND2_X1 U22717 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19804), .ZN(
        P2_U3200) );
  AND2_X1 U22718 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19804), .ZN(P2_U3201) );
  AND2_X1 U22719 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19804), .ZN(P2_U3202) );
  AND2_X1 U22720 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19804), .ZN(P2_U3203) );
  AND2_X1 U22721 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19804), .ZN(P2_U3204) );
  AND2_X1 U22722 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19804), .ZN(P2_U3205) );
  AND2_X1 U22723 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19804), .ZN(P2_U3206) );
  NOR2_X1 U22724 ( .A1(n21006), .A2(n19807), .ZN(P2_U3207) );
  AND2_X1 U22725 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19804), .ZN(P2_U3208) );
  NOR2_X1 U22726 ( .A1(n19736), .A2(n19858), .ZN(n19746) );
  NAND2_X1 U22727 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(
        P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19737) );
  OAI21_X1 U22728 ( .B1(n19746), .B2(n19737), .A(n19752), .ZN(n19739) );
  INV_X1 U22729 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19740) );
  OAI211_X1 U22730 ( .C1(HOLD), .C2(n19740), .A(n19869), .B(n19748), .ZN(
        n19738) );
  OAI211_X1 U22731 ( .C1(n19744), .C2(n20718), .A(n19739), .B(n19738), .ZN(
        P2_U3209) );
  NAND2_X1 U22732 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20723), .ZN(n19745) );
  AOI21_X1 U22733 ( .B1(P2_STATE_REG_2__SCAN_IN), .B2(n19745), .A(n19740), 
        .ZN(n19741) );
  AOI211_X1 U22734 ( .C1(n19741), .C2(n19744), .A(n19861), .B(n19746), .ZN(
        n19742) );
  OAI21_X1 U22735 ( .B1(n20723), .B2(n19743), .A(n19742), .ZN(P2_U3210) );
  OAI22_X1 U22736 ( .A1(n19746), .A2(n19745), .B1(n20718), .B2(n19744), .ZN(
        n19751) );
  INV_X1 U22737 ( .A(n19746), .ZN(n19747) );
  OAI22_X1 U22738 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19748), .B1(NA), 
        .B2(n19747), .ZN(n19749) );
  OAI211_X1 U22739 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19749), .ZN(n19750) );
  OAI21_X1 U22740 ( .B1(n19752), .B2(n19751), .A(n19750), .ZN(P2_U3211) );
  NAND2_X1 U22741 ( .A1(n19792), .A2(n19752), .ZN(n19797) );
  CLKBUF_X1 U22742 ( .A(n19797), .Z(n19793) );
  OAI222_X1 U22743 ( .A1(n19794), .A2(n19754), .B1(n19753), .B2(n19792), .C1(
        n19756), .C2(n19793), .ZN(P2_U3212) );
  OAI222_X1 U22744 ( .A1(n19794), .A2(n19756), .B1(n19755), .B2(n19792), .C1(
        n13887), .C2(n19793), .ZN(P2_U3213) );
  OAI222_X1 U22745 ( .A1(n19794), .A2(n13887), .B1(n19757), .B2(n19792), .C1(
        n11256), .C2(n19793), .ZN(P2_U3214) );
  OAI222_X1 U22746 ( .A1(n19793), .A2(n19758), .B1(n21027), .B2(n19792), .C1(
        n11256), .C2(n19794), .ZN(P2_U3215) );
  OAI222_X1 U22747 ( .A1(n19797), .A2(n19760), .B1(n19759), .B2(n19792), .C1(
        n19758), .C2(n19794), .ZN(P2_U3216) );
  OAI222_X1 U22748 ( .A1(n19797), .A2(n19762), .B1(n19761), .B2(n19792), .C1(
        n19760), .C2(n19794), .ZN(P2_U3217) );
  OAI222_X1 U22749 ( .A1(n19797), .A2(n11271), .B1(n19763), .B2(n19792), .C1(
        n19762), .C2(n19794), .ZN(P2_U3218) );
  OAI222_X1 U22750 ( .A1(n19797), .A2(n11312), .B1(n19764), .B2(n19792), .C1(
        n11271), .C2(n19794), .ZN(P2_U3219) );
  OAI222_X1 U22751 ( .A1(n19797), .A2(n11318), .B1(n19765), .B2(n19792), .C1(
        n11312), .C2(n19794), .ZN(P2_U3220) );
  INV_X1 U22752 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n19767) );
  OAI222_X1 U22753 ( .A1(n19793), .A2(n19767), .B1(n19766), .B2(n19792), .C1(
        n11318), .C2(n19794), .ZN(P2_U3221) );
  OAI222_X1 U22754 ( .A1(n19793), .A2(n11358), .B1(n19768), .B2(n19792), .C1(
        n19767), .C2(n19794), .ZN(P2_U3222) );
  OAI222_X1 U22755 ( .A1(n19793), .A2(n11397), .B1(n19769), .B2(n19792), .C1(
        n11358), .C2(n19794), .ZN(P2_U3223) );
  OAI222_X1 U22756 ( .A1(n19793), .A2(n11400), .B1(n19770), .B2(n19792), .C1(
        n11397), .C2(n19794), .ZN(P2_U3224) );
  OAI222_X1 U22757 ( .A1(n19793), .A2(n11437), .B1(n19771), .B2(n19792), .C1(
        n11400), .C2(n19794), .ZN(P2_U3225) );
  OAI222_X1 U22758 ( .A1(n19793), .A2(n11442), .B1(n19772), .B2(n19792), .C1(
        n11437), .C2(n19794), .ZN(P2_U3226) );
  OAI222_X1 U22759 ( .A1(n19797), .A2(n19773), .B1(n20935), .B2(n19792), .C1(
        n11442), .C2(n19794), .ZN(P2_U3227) );
  OAI222_X1 U22760 ( .A1(n19797), .A2(n11447), .B1(n19774), .B2(n19792), .C1(
        n19773), .C2(n19794), .ZN(P2_U3228) );
  OAI222_X1 U22761 ( .A1(n19797), .A2(n19776), .B1(n19775), .B2(n19792), .C1(
        n11447), .C2(n19794), .ZN(P2_U3229) );
  OAI222_X1 U22762 ( .A1(n19797), .A2(n11452), .B1(n19777), .B2(n19792), .C1(
        n19776), .C2(n19794), .ZN(P2_U3230) );
  OAI222_X1 U22763 ( .A1(n19797), .A2(n19779), .B1(n19778), .B2(n19792), .C1(
        n11452), .C2(n19794), .ZN(P2_U3231) );
  OAI222_X1 U22764 ( .A1(n19797), .A2(n19781), .B1(n19780), .B2(n19792), .C1(
        n19779), .C2(n19794), .ZN(P2_U3232) );
  OAI222_X1 U22765 ( .A1(n19793), .A2(n19783), .B1(n19782), .B2(n19792), .C1(
        n19781), .C2(n19794), .ZN(P2_U3233) );
  OAI222_X1 U22766 ( .A1(n19793), .A2(n11461), .B1(n19784), .B2(n19792), .C1(
        n19783), .C2(n19794), .ZN(P2_U3234) );
  OAI222_X1 U22767 ( .A1(n19793), .A2(n19786), .B1(n19785), .B2(n19792), .C1(
        n11461), .C2(n19794), .ZN(P2_U3235) );
  OAI222_X1 U22768 ( .A1(n19793), .A2(n11464), .B1(n19787), .B2(n19792), .C1(
        n19786), .C2(n19794), .ZN(P2_U3236) );
  OAI222_X1 U22769 ( .A1(n19793), .A2(n19790), .B1(n19788), .B2(n19792), .C1(
        n11464), .C2(n19794), .ZN(P2_U3237) );
  OAI222_X1 U22770 ( .A1(n19794), .A2(n19790), .B1(n19789), .B2(n19792), .C1(
        n11469), .C2(n19793), .ZN(P2_U3238) );
  OAI222_X1 U22771 ( .A1(n19793), .A2(n21124), .B1(n19791), .B2(n19792), .C1(
        n11469), .C2(n19794), .ZN(P2_U3239) );
  OAI222_X1 U22772 ( .A1(n19793), .A2(n11474), .B1(n20955), .B2(n19792), .C1(
        n21124), .C2(n19794), .ZN(P2_U3240) );
  OAI222_X1 U22773 ( .A1(n19797), .A2(n19796), .B1(n19795), .B2(n19792), .C1(
        n11474), .C2(n19794), .ZN(P2_U3241) );
  INV_X1 U22774 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n19798) );
  AOI22_X1 U22775 ( .A1(n19792), .A2(n19799), .B1(n19798), .B2(n19869), .ZN(
        P2_U3585) );
  MUX2_X1 U22776 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n19792), .Z(P2_U3586) );
  MUX2_X1 U22777 ( .A(P2_BE_N_REG_1__SCAN_IN), .B(P2_BYTEENABLE_REG_1__SCAN_IN), .S(n19792), .Z(P2_U3587) );
  INV_X1 U22778 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n19800) );
  AOI22_X1 U22779 ( .A1(n19792), .A2(n19801), .B1(n19800), .B2(n19869), .ZN(
        P2_U3588) );
  AOI21_X1 U22780 ( .B1(n19804), .B2(n19803), .A(n19802), .ZN(P2_U3591) );
  OAI21_X1 U22781 ( .B1(n19807), .B2(n19806), .A(n19805), .ZN(P2_U3592) );
  INV_X1 U22782 ( .A(n19842), .ZN(n19832) );
  OAI211_X1 U22783 ( .C1(n19811), .C2(n19810), .A(n19809), .B(n19808), .ZN(
        n19819) );
  AOI222_X1 U22784 ( .A1(n19819), .A2(n19815), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n19814), .C1(n19813), .C2(n19812), .ZN(n19816) );
  AOI22_X1 U22785 ( .A1(n19832), .A2(n11933), .B1(n19816), .B2(n19842), .ZN(
        P2_U3602) );
  OAI21_X1 U22786 ( .B1(n19824), .B2(n19827), .A(n19817), .ZN(n19818) );
  AOI22_X1 U22787 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19820), .B1(n19819), 
        .B2(n19818), .ZN(n19821) );
  AOI22_X1 U22788 ( .A1(n19832), .A2(n19822), .B1(n19821), .B2(n19842), .ZN(
        P2_U3603) );
  INV_X1 U22789 ( .A(n19823), .ZN(n19836) );
  OR3_X1 U22790 ( .A1(n19824), .A2(n19836), .A3(n10320), .ZN(n19825) );
  OAI21_X1 U22791 ( .B1(n19827), .B2(n19826), .A(n19825), .ZN(n19828) );
  AOI21_X1 U22792 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19829), .A(n19828), 
        .ZN(n19830) );
  AOI22_X1 U22793 ( .A1(n19832), .A2(n19831), .B1(n19830), .B2(n19842), .ZN(
        P2_U3604) );
  INV_X1 U22794 ( .A(n19833), .ZN(n19835) );
  OAI22_X1 U22795 ( .A1(n19837), .A2(n19836), .B1(n19835), .B2(n19834), .ZN(
        n19839) );
  OAI21_X1 U22796 ( .B1(n19839), .B2(n19838), .A(n19842), .ZN(n19840) );
  OAI21_X1 U22797 ( .B1(n19842), .B2(n19841), .A(n19840), .ZN(P2_U3605) );
  INV_X1 U22798 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19843) );
  AOI22_X1 U22799 ( .A1(n19792), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19843), 
        .B2(n19869), .ZN(P2_U3608) );
  AOI22_X1 U22800 ( .A1(n19846), .A2(n19865), .B1(n19845), .B2(n19844), .ZN(
        n19850) );
  INV_X1 U22801 ( .A(n19847), .ZN(n19848) );
  OAI21_X1 U22802 ( .B1(n19850), .B2(n19849), .A(n19848), .ZN(n19852) );
  MUX2_X1 U22803 ( .A(P2_MORE_REG_SCAN_IN), .B(n19852), .S(n19851), .Z(
        P2_U3609) );
  AOI21_X1 U22804 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n19853), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19855) );
  AOI211_X1 U22805 ( .C1(n19856), .C2(n19858), .A(n19855), .B(n19854), .ZN(
        n19868) );
  AOI21_X1 U22806 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n19861), .A(n19859), 
        .ZN(n19864) );
  AOI22_X1 U22807 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19858), .B1(n19859), 
        .B2(n19857), .ZN(n19863) );
  NOR4_X1 U22808 ( .A1(n19861), .A2(n19860), .A3(n10512), .A4(n19859), .ZN(
        n19862) );
  AOI211_X1 U22809 ( .C1(n19865), .C2(n19864), .A(n19863), .B(n19862), .ZN(
        n19867) );
  NAND2_X1 U22810 ( .A1(n19868), .A2(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n19866) );
  OAI21_X1 U22811 ( .B1(n19868), .B2(n19867), .A(n19866), .ZN(P2_U3610) );
  INV_X1 U22812 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n19870) );
  AOI22_X1 U22813 ( .A1(n19792), .A2(n19871), .B1(n19870), .B2(n19869), .ZN(
        P2_U3611) );
  INV_X1 U22814 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n19872) );
  OAI21_X1 U22815 ( .B1(n19872), .B2(P1_STATE_REG_2__SCAN_IN), .A(
        P1_STATE_REG_0__SCAN_IN), .ZN(n19880) );
  OAI21_X1 U22816 ( .B1(n19880), .B2(P1_ADS_N_REG_SCAN_IN), .A(n20810), .ZN(
        n19873) );
  INV_X1 U22817 ( .A(n19873), .ZN(P1_U2802) );
  INV_X1 U22818 ( .A(n19874), .ZN(n19876) );
  OAI21_X1 U22819 ( .B1(n19876), .B2(n19875), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19877) );
  OAI21_X1 U22820 ( .B1(n19878), .B2(n20706), .A(n19877), .ZN(P1_U2803) );
  NOR2_X1 U22821 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19881) );
  OAI21_X1 U22822 ( .B1(n19881), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20810), .ZN(
        n19879) );
  OAI21_X1 U22823 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20810), .A(n19879), 
        .ZN(P1_U2804) );
  NAND2_X1 U22824 ( .A1(n20810), .A2(n19880), .ZN(n20783) );
  INV_X1 U22825 ( .A(n20783), .ZN(n20787) );
  OAI21_X1 U22826 ( .B1(BS16), .B2(n19881), .A(n20787), .ZN(n20785) );
  OAI21_X1 U22827 ( .B1(n20787), .B2(n20200), .A(n20785), .ZN(P1_U2805) );
  OAI21_X1 U22828 ( .B1(n19884), .B2(n19883), .A(n19882), .ZN(P1_U2806) );
  NOR4_X1 U22829 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_18__SCAN_IN), .A3(P1_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_20__SCAN_IN), .ZN(n19888) );
  NOR4_X1 U22830 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_14__SCAN_IN), .A3(P1_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_16__SCAN_IN), .ZN(n19887) );
  NOR4_X1 U22831 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_27__SCAN_IN), .A3(P1_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n19886) );
  NOR4_X1 U22832 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_23__SCAN_IN), .A3(P1_DATAWIDTH_REG_24__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_25__SCAN_IN), .ZN(n19885) );
  NAND4_X1 U22833 ( .A1(n19888), .A2(n19887), .A3(n19886), .A4(n19885), .ZN(
        n19894) );
  NOR4_X1 U22834 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_2__SCAN_IN), .A3(P1_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_4__SCAN_IN), .ZN(n19892) );
  AOI211_X1 U22835 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_22__SCAN_IN), .B(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19891) );
  NOR4_X1 U22836 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_10__SCAN_IN), .A3(P1_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_12__SCAN_IN), .ZN(n19890) );
  NOR4_X1 U22837 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_6__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_8__SCAN_IN), .ZN(n19889) );
  NAND4_X1 U22838 ( .A1(n19892), .A2(n19891), .A3(n19890), .A4(n19889), .ZN(
        n19893) );
  NOR2_X1 U22839 ( .A1(n19894), .A2(n19893), .ZN(n20806) );
  INV_X1 U22840 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20780) );
  NOR3_X1 U22841 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19896) );
  OAI21_X1 U22842 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19896), .A(n20806), .ZN(
        n19895) );
  OAI21_X1 U22843 ( .B1(n20806), .B2(n20780), .A(n19895), .ZN(P1_U2807) );
  INV_X1 U22844 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20786) );
  AOI21_X1 U22845 ( .B1(n13981), .B2(n20786), .A(n19896), .ZN(n19897) );
  INV_X1 U22846 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20777) );
  INV_X1 U22847 ( .A(n20806), .ZN(n20808) );
  AOI22_X1 U22848 ( .A1(n20806), .A2(n19897), .B1(n20777), .B2(n20808), .ZN(
        P1_U2808) );
  AOI22_X1 U22849 ( .A1(P1_EBX_REG_9__SCAN_IN), .A2(n19961), .B1(n19898), .B2(
        n20739), .ZN(n19909) );
  OAI22_X1 U22850 ( .A1(n19901), .A2(n20739), .B1(n19900), .B2(n19899), .ZN(
        n19902) );
  AOI211_X1 U22851 ( .C1(n19960), .C2(n19903), .A(n19948), .B(n19902), .ZN(
        n19908) );
  INV_X1 U22852 ( .A(n19904), .ZN(n19906) );
  AOI22_X1 U22853 ( .A1(n19906), .A2(n19928), .B1(n19971), .B2(n19905), .ZN(
        n19907) );
  NAND3_X1 U22854 ( .A1(n19909), .A2(n19908), .A3(n19907), .ZN(P1_U2831) );
  AOI21_X1 U22855 ( .B1(n19945), .B2(n19919), .A(n19932), .ZN(n19925) );
  AOI22_X1 U22856 ( .A1(P1_EBX_REG_7__SCAN_IN), .A2(n19961), .B1(n19960), .B2(
        n19910), .ZN(n19911) );
  OAI21_X1 U22857 ( .B1(n19912), .B2(n19959), .A(n19911), .ZN(n19916) );
  NOR3_X1 U22858 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19934), .A3(n19919), .ZN(
        n19913) );
  AOI211_X1 U22859 ( .C1(n19964), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n19948), .B(n19913), .ZN(n19914) );
  INV_X1 U22860 ( .A(n19914), .ZN(n19915) );
  AOI211_X1 U22861 ( .C1(n19928), .C2(n19917), .A(n19916), .B(n19915), .ZN(
        n19918) );
  OAI21_X1 U22862 ( .B1(n19925), .B2(n20735), .A(n19918), .ZN(P1_U2833) );
  AND2_X1 U22863 ( .A1(n19919), .A2(n19945), .ZN(n19920) );
  AOI22_X1 U22864 ( .A1(n19960), .A2(n19922), .B1(n19921), .B2(n19920), .ZN(
        n19930) );
  INV_X1 U22865 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20733) );
  AOI22_X1 U22866 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n19964), .B1(
        P1_EBX_REG_6__SCAN_IN), .B2(n19961), .ZN(n19924) );
  OAI211_X1 U22867 ( .C1(n19925), .C2(n20733), .A(n19924), .B(n19923), .ZN(
        n19926) );
  AOI21_X1 U22868 ( .B1(n19928), .B2(n19927), .A(n19926), .ZN(n19929) );
  OAI211_X1 U22869 ( .C1(n19931), .C2(n19959), .A(n19930), .B(n19929), .ZN(
        P1_U2834) );
  AOI21_X1 U22870 ( .B1(n19945), .B2(n19933), .A(n19932), .ZN(n19956) );
  NOR3_X1 U22871 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n19934), .A3(n19933), .ZN(
        n19935) );
  AOI211_X1 U22872 ( .C1(n19964), .C2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n19948), .B(n19935), .ZN(n19942) );
  AOI22_X1 U22873 ( .A1(P1_EBX_REG_5__SCAN_IN), .A2(n19961), .B1(n19960), .B2(
        n19936), .ZN(n19941) );
  INV_X1 U22874 ( .A(n19937), .ZN(n19938) );
  AOI22_X1 U22875 ( .A1(n19939), .A2(n19952), .B1(n19938), .B2(n19971), .ZN(
        n19940) );
  AND3_X1 U22876 ( .A1(n19942), .A2(n19941), .A3(n19940), .ZN(n19943) );
  OAI21_X1 U22877 ( .B1(n19956), .B2(n20732), .A(n19943), .ZN(P1_U2835) );
  AND3_X1 U22878 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n19944) );
  AOI21_X1 U22879 ( .B1(n19945), .B2(n19944), .A(P1_REIP_REG_4__SCAN_IN), .ZN(
        n19955) );
  INV_X1 U22880 ( .A(n19946), .ZN(n20080) );
  AOI22_X1 U22881 ( .A1(P1_EBX_REG_4__SCAN_IN), .A2(n19961), .B1(n19947), .B2(
        n19965), .ZN(n19950) );
  AOI21_X1 U22882 ( .B1(n19964), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n19948), .ZN(n19949) );
  NAND2_X1 U22883 ( .A1(n19950), .A2(n19949), .ZN(n19951) );
  AOI21_X1 U22884 ( .B1(n19960), .B2(n20080), .A(n19951), .ZN(n19954) );
  NAND2_X1 U22885 ( .A1(n20070), .A2(n19952), .ZN(n19953) );
  OAI211_X1 U22886 ( .C1(n19956), .C2(n19955), .A(n19954), .B(n19953), .ZN(
        n19957) );
  INV_X1 U22887 ( .A(n19957), .ZN(n19958) );
  OAI21_X1 U22888 ( .B1(n20075), .B2(n19959), .A(n19958), .ZN(P1_U2836) );
  AOI22_X1 U22889 ( .A1(P1_EBX_REG_3__SCAN_IN), .A2(n19961), .B1(n19960), .B2(
        n20086), .ZN(n19974) );
  NAND2_X1 U22890 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n19962) );
  OAI211_X1 U22891 ( .C1(P1_REIP_REG_3__SCAN_IN), .C2(P1_REIP_REG_2__SCAN_IN), 
        .A(n19963), .B(n19962), .ZN(n19967) );
  AOI22_X1 U22892 ( .A1(n20397), .A2(n19965), .B1(n19964), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n19966) );
  OAI211_X1 U22893 ( .C1(n19969), .C2(n19968), .A(n19967), .B(n19966), .ZN(
        n19970) );
  AOI21_X1 U22894 ( .B1(n19972), .B2(n19971), .A(n19970), .ZN(n19973) );
  OAI211_X1 U22895 ( .C1(n19975), .C2(n13791), .A(n19974), .B(n19973), .ZN(
        P1_U2837) );
  AOI22_X1 U22896 ( .A1(n20819), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n19977) );
  OAI21_X1 U22897 ( .B1(n20063), .B2(n20007), .A(n19977), .ZN(P1_U2921) );
  AOI22_X1 U22898 ( .A1(n20819), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n19978) );
  OAI21_X1 U22899 ( .B1(n19979), .B2(n20007), .A(n19978), .ZN(P1_U2922) );
  AOI22_X1 U22900 ( .A1(n20819), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n19980) );
  OAI21_X1 U22901 ( .B1(n19981), .B2(n20007), .A(n19980), .ZN(P1_U2923) );
  AOI22_X1 U22902 ( .A1(n20819), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n19982) );
  OAI21_X1 U22903 ( .B1(n19983), .B2(n20007), .A(n19982), .ZN(P1_U2924) );
  AOI22_X1 U22904 ( .A1(n20819), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n19984) );
  OAI21_X1 U22905 ( .B1(n19985), .B2(n20007), .A(n19984), .ZN(P1_U2925) );
  AOI22_X1 U22906 ( .A1(n20819), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n19986) );
  OAI21_X1 U22907 ( .B1(n19987), .B2(n20007), .A(n19986), .ZN(P1_U2926) );
  AOI22_X1 U22908 ( .A1(n20819), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n19988) );
  OAI21_X1 U22909 ( .B1(n19989), .B2(n20007), .A(n19988), .ZN(P1_U2927) );
  AOI22_X1 U22910 ( .A1(n20819), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n19990) );
  OAI21_X1 U22911 ( .B1(n19991), .B2(n20007), .A(n19990), .ZN(P1_U2928) );
  AOI22_X1 U22912 ( .A1(n20005), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n19992) );
  OAI21_X1 U22913 ( .B1(n12639), .B2(n20007), .A(n19992), .ZN(P1_U2929) );
  AOI22_X1 U22914 ( .A1(n20005), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n19993) );
  OAI21_X1 U22915 ( .B1(n12629), .B2(n20007), .A(n19993), .ZN(P1_U2930) );
  AOI22_X1 U22916 ( .A1(n20005), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n19994) );
  OAI21_X1 U22917 ( .B1(n19995), .B2(n20007), .A(n19994), .ZN(P1_U2931) );
  AOI22_X1 U22918 ( .A1(n20005), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n19996) );
  OAI21_X1 U22919 ( .B1(n19997), .B2(n20007), .A(n19996), .ZN(P1_U2932) );
  AOI22_X1 U22920 ( .A1(n20005), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n19998) );
  OAI21_X1 U22921 ( .B1(n19999), .B2(n20007), .A(n19998), .ZN(P1_U2933) );
  AOI22_X1 U22922 ( .A1(n20005), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20000) );
  OAI21_X1 U22923 ( .B1(n20001), .B2(n20007), .A(n20000), .ZN(P1_U2934) );
  AOI22_X1 U22924 ( .A1(n20005), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20002) );
  OAI21_X1 U22925 ( .B1(n20003), .B2(n20007), .A(n20002), .ZN(P1_U2935) );
  AOI22_X1 U22926 ( .A1(n20005), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n20004), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20006) );
  OAI21_X1 U22927 ( .B1(n20008), .B2(n20007), .A(n20006), .ZN(P1_U2936) );
  NOR2_X1 U22928 ( .A1(n20009), .A2(n20818), .ZN(n20010) );
  OR2_X2 U22929 ( .A1(n20011), .A2(n20010), .ZN(n20059) );
  OR2_X2 U22930 ( .A1(n20013), .A2(n20012), .ZN(n20062) );
  INV_X1 U22931 ( .A(n20062), .ZN(n20021) );
  AOI22_X1 U22932 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20059), .B1(n20021), 
        .B2(n20014), .ZN(n20015) );
  OAI21_X1 U22933 ( .B1(n20016), .B2(n20064), .A(n20015), .ZN(P1_U2937) );
  AOI22_X1 U22934 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20059), .B1(n20021), 
        .B2(n20017), .ZN(n20018) );
  OAI21_X1 U22935 ( .B1(n20019), .B2(n20064), .A(n20018), .ZN(P1_U2938) );
  AOI22_X1 U22936 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20059), .B1(n20021), 
        .B2(n20020), .ZN(n20022) );
  OAI21_X1 U22937 ( .B1(n20023), .B2(n20064), .A(n20022), .ZN(P1_U2939) );
  INV_X2 U22938 ( .A(n20064), .ZN(n20056) );
  AOI22_X1 U22939 ( .A1(P1_EAX_REG_19__SCAN_IN), .A2(n20056), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20059), .ZN(n20024) );
  OAI21_X1 U22940 ( .B1(n20147), .B2(n20062), .A(n20024), .ZN(P1_U2940) );
  AOI22_X1 U22941 ( .A1(P1_EAX_REG_20__SCAN_IN), .A2(n20056), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20059), .ZN(n20025) );
  OAI21_X1 U22942 ( .B1(n20151), .B2(n20062), .A(n20025), .ZN(P1_U2941) );
  AOI22_X1 U22943 ( .A1(P1_EAX_REG_21__SCAN_IN), .A2(n20056), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20059), .ZN(n20026) );
  OAI21_X1 U22944 ( .B1(n20155), .B2(n20062), .A(n20026), .ZN(P1_U2942) );
  AOI22_X1 U22945 ( .A1(P1_EAX_REG_22__SCAN_IN), .A2(n20056), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20059), .ZN(n20027) );
  OAI21_X1 U22946 ( .B1(n20159), .B2(n20062), .A(n20027), .ZN(P1_U2943) );
  AOI22_X1 U22947 ( .A1(P1_EAX_REG_23__SCAN_IN), .A2(n20056), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20059), .ZN(n20028) );
  OAI21_X1 U22948 ( .B1(n20165), .B2(n20062), .A(n20028), .ZN(P1_U2944) );
  AOI22_X1 U22949 ( .A1(P1_EAX_REG_24__SCAN_IN), .A2(n20056), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20059), .ZN(n20029) );
  OAI21_X1 U22950 ( .B1(n20045), .B2(n20062), .A(n20029), .ZN(P1_U2945) );
  AOI22_X1 U22951 ( .A1(P1_EAX_REG_25__SCAN_IN), .A2(n20056), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20059), .ZN(n20030) );
  OAI21_X1 U22952 ( .B1(n20047), .B2(n20062), .A(n20030), .ZN(P1_U2946) );
  AOI22_X1 U22953 ( .A1(P1_EAX_REG_26__SCAN_IN), .A2(n20056), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n20059), .ZN(n20031) );
  OAI21_X1 U22954 ( .B1(n20049), .B2(n20062), .A(n20031), .ZN(P1_U2947) );
  AOI22_X1 U22955 ( .A1(P1_EAX_REG_27__SCAN_IN), .A2(n20056), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n20059), .ZN(n20032) );
  OAI21_X1 U22956 ( .B1(n20051), .B2(n20062), .A(n20032), .ZN(P1_U2948) );
  AOI22_X1 U22957 ( .A1(P1_EAX_REG_28__SCAN_IN), .A2(n20056), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n20059), .ZN(n20033) );
  OAI21_X1 U22958 ( .B1(n20053), .B2(n20062), .A(n20033), .ZN(P1_U2949) );
  AOI22_X1 U22959 ( .A1(P1_EAX_REG_29__SCAN_IN), .A2(n20056), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n20059), .ZN(n20034) );
  OAI21_X1 U22960 ( .B1(n20055), .B2(n20062), .A(n20034), .ZN(P1_U2950) );
  AOI22_X1 U22961 ( .A1(P1_EAX_REG_30__SCAN_IN), .A2(n20056), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n20059), .ZN(n20035) );
  OAI21_X1 U22962 ( .B1(n20058), .B2(n20062), .A(n20035), .ZN(P1_U2951) );
  AOI22_X1 U22963 ( .A1(P1_EAX_REG_0__SCAN_IN), .A2(n20056), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20059), .ZN(n20036) );
  OAI21_X1 U22964 ( .B1(n20131), .B2(n20062), .A(n20036), .ZN(P1_U2952) );
  AOI22_X1 U22965 ( .A1(P1_EAX_REG_1__SCAN_IN), .A2(n20056), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20059), .ZN(n20037) );
  OAI21_X1 U22966 ( .B1(n20140), .B2(n20062), .A(n20037), .ZN(P1_U2953) );
  AOI22_X1 U22967 ( .A1(P1_EAX_REG_2__SCAN_IN), .A2(n20056), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20059), .ZN(n20038) );
  OAI21_X1 U22968 ( .B1(n20143), .B2(n20062), .A(n20038), .ZN(P1_U2954) );
  AOI22_X1 U22969 ( .A1(P1_EAX_REG_3__SCAN_IN), .A2(n20056), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20059), .ZN(n20039) );
  OAI21_X1 U22970 ( .B1(n20147), .B2(n20062), .A(n20039), .ZN(P1_U2955) );
  AOI22_X1 U22971 ( .A1(P1_EAX_REG_4__SCAN_IN), .A2(n20056), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20059), .ZN(n20040) );
  OAI21_X1 U22972 ( .B1(n20151), .B2(n20062), .A(n20040), .ZN(P1_U2956) );
  AOI22_X1 U22973 ( .A1(P1_EAX_REG_5__SCAN_IN), .A2(n20056), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20059), .ZN(n20041) );
  OAI21_X1 U22974 ( .B1(n20155), .B2(n20062), .A(n20041), .ZN(P1_U2957) );
  AOI22_X1 U22975 ( .A1(P1_EAX_REG_6__SCAN_IN), .A2(n20056), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20059), .ZN(n20042) );
  OAI21_X1 U22976 ( .B1(n20159), .B2(n20062), .A(n20042), .ZN(P1_U2958) );
  AOI22_X1 U22977 ( .A1(P1_EAX_REG_7__SCAN_IN), .A2(n20056), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20059), .ZN(n20043) );
  OAI21_X1 U22978 ( .B1(n20165), .B2(n20062), .A(n20043), .ZN(P1_U2959) );
  AOI22_X1 U22979 ( .A1(P1_EAX_REG_8__SCAN_IN), .A2(n20056), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n20059), .ZN(n20044) );
  OAI21_X1 U22980 ( .B1(n20045), .B2(n20062), .A(n20044), .ZN(P1_U2960) );
  AOI22_X1 U22981 ( .A1(P1_EAX_REG_9__SCAN_IN), .A2(n20056), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20059), .ZN(n20046) );
  OAI21_X1 U22982 ( .B1(n20047), .B2(n20062), .A(n20046), .ZN(P1_U2961) );
  AOI22_X1 U22983 ( .A1(P1_EAX_REG_10__SCAN_IN), .A2(n20056), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20059), .ZN(n20048) );
  OAI21_X1 U22984 ( .B1(n20049), .B2(n20062), .A(n20048), .ZN(P1_U2962) );
  AOI22_X1 U22985 ( .A1(P1_EAX_REG_11__SCAN_IN), .A2(n20056), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20059), .ZN(n20050) );
  OAI21_X1 U22986 ( .B1(n20051), .B2(n20062), .A(n20050), .ZN(P1_U2963) );
  AOI22_X1 U22987 ( .A1(P1_EAX_REG_12__SCAN_IN), .A2(n20056), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20059), .ZN(n20052) );
  OAI21_X1 U22988 ( .B1(n20053), .B2(n20062), .A(n20052), .ZN(P1_U2964) );
  AOI22_X1 U22989 ( .A1(P1_EAX_REG_13__SCAN_IN), .A2(n20056), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20059), .ZN(n20054) );
  OAI21_X1 U22990 ( .B1(n20055), .B2(n20062), .A(n20054), .ZN(P1_U2965) );
  AOI22_X1 U22991 ( .A1(P1_EAX_REG_14__SCAN_IN), .A2(n20056), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20059), .ZN(n20057) );
  OAI21_X1 U22992 ( .B1(n20058), .B2(n20062), .A(n20057), .ZN(P1_U2966) );
  INV_X1 U22993 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n21007) );
  INV_X1 U22994 ( .A(n20059), .ZN(n20060) );
  OAI222_X1 U22995 ( .A1(n20064), .A2(n20063), .B1(n20062), .B2(n20061), .C1(
        n21007), .C2(n20060), .ZN(P1_U2967) );
  AOI22_X1 U22996 ( .A1(n20065), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n13703), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20074) );
  OAI21_X1 U22997 ( .B1(n20068), .B2(n20067), .A(n20066), .ZN(n20069) );
  INV_X1 U22998 ( .A(n20069), .ZN(n20079) );
  AOI22_X1 U22999 ( .A1(n20079), .A2(n20072), .B1(n20071), .B2(n20070), .ZN(
        n20073) );
  OAI211_X1 U23000 ( .C1(n20076), .C2(n20075), .A(n20074), .B(n20073), .ZN(
        P1_U2995) );
  AOI21_X1 U23001 ( .B1(n20078), .B2(n20100), .A(n20077), .ZN(n20093) );
  AOI222_X1 U23002 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n13703), .B1(n20110), 
        .B2(n20080), .C1(n20087), .C2(n20079), .ZN(n20083) );
  OAI211_X1 U23003 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n20089), .B(n20081), .ZN(n20082) );
  OAI211_X1 U23004 ( .C1(n20093), .C2(n20084), .A(n20083), .B(n20082), .ZN(
        P1_U3027) );
  AOI21_X1 U23005 ( .B1(n20110), .B2(n20086), .A(n20085), .ZN(n20091) );
  AOI22_X1 U23006 ( .A1(n20089), .A2(n20092), .B1(n20088), .B2(n20087), .ZN(
        n20090) );
  OAI211_X1 U23007 ( .C1(n20093), .C2(n20092), .A(n20091), .B(n20090), .ZN(
        P1_U3028) );
  INV_X1 U23008 ( .A(n20094), .ZN(n20114) );
  AOI21_X1 U23009 ( .B1(n20098), .B2(n20096), .A(n20095), .ZN(n20112) );
  INV_X1 U23010 ( .A(n20097), .ZN(n20109) );
  NOR2_X1 U23011 ( .A1(n20099), .A2(n20098), .ZN(n20101) );
  AOI21_X1 U23012 ( .B1(n20101), .B2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n20100), .ZN(n20103) );
  OAI22_X1 U23013 ( .A1(n20104), .A2(n20103), .B1(n20727), .B2(n20102), .ZN(
        n20108) );
  NOR2_X1 U23014 ( .A1(n20106), .A2(n20105), .ZN(n20107) );
  AOI211_X1 U23015 ( .C1(n20110), .C2(n20109), .A(n20108), .B(n20107), .ZN(
        n20111) );
  OAI221_X1 U23016 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20114), .C1(
        n20113), .C2(n20112), .A(n20111), .ZN(P1_U3029) );
  NOR2_X1 U23017 ( .A1(n20116), .A2(n20115), .ZN(P1_U3032) );
  NOR2_X2 U23018 ( .A1(n20120), .A2(n20119), .ZN(n20162) );
  INV_X1 U23019 ( .A(n13164), .ZN(n20123) );
  AOI22_X1 U23020 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20162), .B1(DATAI_24_), 
        .B2(n20118), .ZN(n20544) );
  INV_X1 U23021 ( .A(n20544), .ZN(n20653) );
  NAND2_X1 U23022 ( .A1(n20453), .A2(n20398), .ZN(n20237) );
  OR2_X1 U23023 ( .A1(n20529), .A2(n20237), .ZN(n20129) );
  INV_X1 U23024 ( .A(n20129), .ZN(n20164) );
  OR2_X1 U23025 ( .A1(n20124), .A2(n20158), .ZN(n20448) );
  AOI22_X1 U23026 ( .A1(n20699), .A2(n20653), .B1(n20164), .B2(n20650), .ZN(
        n20138) );
  INV_X1 U23027 ( .A(n20454), .ZN(n20125) );
  NOR2_X1 U23028 ( .A1(n20399), .A2(n20125), .ZN(n20134) );
  NAND2_X1 U23029 ( .A1(n20133), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20593) );
  AND2_X1 U23030 ( .A1(n20172), .A2(n20593), .ZN(n20456) );
  INV_X1 U23031 ( .A(n20699), .ZN(n20126) );
  NAND3_X1 U23032 ( .A1(n20126), .A2(n20570), .A3(n20190), .ZN(n20127) );
  NAND2_X1 U23033 ( .A1(n20570), .A2(n20200), .ZN(n20531) );
  NAND2_X1 U23034 ( .A1(n20127), .A2(n20531), .ZN(n20132) );
  NAND2_X1 U23035 ( .A1(n9928), .A2(n20535), .ZN(n20135) );
  AOI22_X1 U23036 ( .A1(n20132), .A2(n20135), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20129), .ZN(n20130) );
  OAI211_X1 U23037 ( .C1(n20134), .C2(n20708), .A(n20456), .B(n20130), .ZN(
        n20167) );
  NOR2_X2 U23038 ( .A1(n20131), .A2(n20284), .ZN(n20651) );
  INV_X1 U23039 ( .A(n20132), .ZN(n20136) );
  OR2_X1 U23040 ( .A1(n20133), .A2(n20708), .ZN(n20459) );
  INV_X1 U23041 ( .A(n20134), .ZN(n20279) );
  OAI22_X1 U23042 ( .A1(n20136), .A2(n20135), .B1(n20459), .B2(n20279), .ZN(
        n20166) );
  AOI22_X1 U23043 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20167), .B1(
        n20651), .B2(n20166), .ZN(n20137) );
  OAI211_X1 U23044 ( .C1(n20603), .C2(n20190), .A(n20138), .B(n20137), .ZN(
        P1_U3033) );
  AOI22_X1 U23045 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20162), .B1(DATAI_17_), 
        .B2(n20118), .ZN(n20607) );
  AOI22_X1 U23046 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20162), .B1(DATAI_25_), 
        .B2(n20118), .ZN(n20663) );
  INV_X1 U23047 ( .A(n20663), .ZN(n20604) );
  NOR2_X2 U23048 ( .A1(n20139), .A2(n20158), .ZN(n20657) );
  AOI22_X1 U23049 ( .A1(n20699), .A2(n20604), .B1(n20164), .B2(n20657), .ZN(
        n20142) );
  NOR2_X2 U23050 ( .A1(n20140), .A2(n20284), .ZN(n20658) );
  AOI22_X1 U23051 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20167), .B1(
        n20658), .B2(n20166), .ZN(n20141) );
  OAI211_X1 U23052 ( .C1(n20607), .C2(n20190), .A(n20142), .B(n20141), .ZN(
        P1_U3034) );
  AOI22_X1 U23053 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20162), .B1(DATAI_18_), 
        .B2(n20118), .ZN(n20611) );
  INV_X1 U23054 ( .A(n20669), .ZN(n20608) );
  AOI22_X1 U23055 ( .A1(n20699), .A2(n20608), .B1(n20164), .B2(n20664), .ZN(
        n20145) );
  NOR2_X2 U23056 ( .A1(n20143), .A2(n20284), .ZN(n20665) );
  AOI22_X1 U23057 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20167), .B1(
        n20665), .B2(n20166), .ZN(n20144) );
  OAI211_X1 U23058 ( .C1(n20611), .C2(n20190), .A(n20145), .B(n20144), .ZN(
        P1_U3035) );
  AOI22_X1 U23059 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20162), .B1(DATAI_27_), 
        .B2(n20118), .ZN(n20675) );
  INV_X1 U23060 ( .A(n20675), .ZN(n20612) );
  AOI22_X1 U23061 ( .A1(n20699), .A2(n20612), .B1(n20164), .B2(n20670), .ZN(
        n20149) );
  NOR2_X2 U23062 ( .A1(n20147), .A2(n20284), .ZN(n20671) );
  AOI22_X1 U23063 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20167), .B1(
        n20671), .B2(n20166), .ZN(n20148) );
  OAI211_X1 U23064 ( .C1(n20615), .C2(n20190), .A(n20149), .B(n20148), .ZN(
        P1_U3036) );
  AOI22_X1 U23065 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20162), .B1(DATAI_20_), 
        .B2(n20118), .ZN(n20619) );
  AOI22_X1 U23066 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20162), .B1(DATAI_28_), 
        .B2(n20118), .ZN(n20681) );
  INV_X1 U23067 ( .A(n20681), .ZN(n20616) );
  OR2_X1 U23068 ( .A1(n20150), .A2(n20158), .ZN(n20475) );
  AOI22_X1 U23069 ( .A1(n20699), .A2(n20616), .B1(n20164), .B2(n20676), .ZN(
        n20153) );
  NOR2_X2 U23070 ( .A1(n20151), .A2(n20284), .ZN(n20677) );
  AOI22_X1 U23071 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20167), .B1(
        n20677), .B2(n20166), .ZN(n20152) );
  OAI211_X1 U23072 ( .C1(n20619), .C2(n20190), .A(n20153), .B(n20152), .ZN(
        P1_U3037) );
  AOI22_X1 U23073 ( .A1(DATAI_21_), .A2(n20118), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n20162), .ZN(n20623) );
  AOI22_X1 U23074 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20162), .B1(DATAI_29_), 
        .B2(n20118), .ZN(n20687) );
  INV_X1 U23075 ( .A(n20687), .ZN(n20620) );
  AOI22_X1 U23076 ( .A1(n20699), .A2(n20620), .B1(n20164), .B2(n20682), .ZN(
        n20157) );
  NOR2_X2 U23077 ( .A1(n20155), .A2(n20284), .ZN(n20683) );
  AOI22_X1 U23078 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20167), .B1(
        n20683), .B2(n20166), .ZN(n20156) );
  OAI211_X1 U23079 ( .C1(n20623), .C2(n20190), .A(n20157), .B(n20156), .ZN(
        P1_U3038) );
  AOI22_X1 U23080 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20162), .B1(DATAI_22_), 
        .B2(n20118), .ZN(n20627) );
  INV_X1 U23081 ( .A(n20693), .ZN(n20624) );
  OR2_X1 U23082 ( .A1(n12402), .A2(n20158), .ZN(n20483) );
  AOI22_X1 U23083 ( .A1(n20699), .A2(n20624), .B1(n20164), .B2(n20688), .ZN(
        n20161) );
  NOR2_X2 U23084 ( .A1(n20159), .A2(n20284), .ZN(n20689) );
  AOI22_X1 U23085 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20167), .B1(
        n20689), .B2(n20166), .ZN(n20160) );
  OAI211_X1 U23086 ( .C1(n20627), .C2(n20190), .A(n20161), .B(n20160), .ZN(
        P1_U3039) );
  AOI22_X1 U23087 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20162), .B1(DATAI_23_), 
        .B2(n20118), .ZN(n20635) );
  AOI22_X1 U23088 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n20162), .B1(DATAI_31_), 
        .B2(n20118), .ZN(n20704) );
  INV_X1 U23089 ( .A(n20704), .ZN(n20630) );
  AOI22_X1 U23090 ( .A1(n20699), .A2(n20630), .B1(n20164), .B2(n20695), .ZN(
        n20169) );
  NOR2_X2 U23091 ( .A1(n20165), .A2(n20284), .ZN(n20697) );
  AOI22_X1 U23092 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20167), .B1(
        n20697), .B2(n20166), .ZN(n20168) );
  OAI211_X1 U23093 ( .C1(n20635), .C2(n20190), .A(n20169), .B(n20168), .ZN(
        P1_U3040) );
  INV_X1 U23094 ( .A(n20170), .ZN(n20564) );
  NOR3_X2 U23095 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20563), .A3(
        n20237), .ZN(n20191) );
  AOI21_X1 U23096 ( .B1(n9928), .B2(n20564), .A(n20191), .ZN(n20173) );
  NOR2_X1 U23097 ( .A1(n20237), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20175) );
  INV_X1 U23098 ( .A(n20175), .ZN(n20171) );
  OAI22_X1 U23099 ( .A1(n20173), .A2(n20648), .B1(n20171), .B2(n20708), .ZN(
        n20192) );
  AOI22_X1 U23100 ( .A1(n20651), .A2(n20192), .B1(n20650), .B2(n20191), .ZN(
        n20177) );
  OAI21_X1 U23101 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n20537), .A(
        n20172), .ZN(n20241) );
  OAI211_X1 U23102 ( .C1(n20239), .C2(n20425), .A(n20570), .B(n20173), .ZN(
        n20174) );
  OAI211_X1 U23103 ( .C1(n20570), .C2(n20175), .A(n20640), .B(n20174), .ZN(
        n20194) );
  INV_X1 U23104 ( .A(n20190), .ZN(n20193) );
  AOI22_X1 U23105 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20194), .B1(
        n20193), .B2(n20653), .ZN(n20176) );
  OAI211_X1 U23106 ( .C1(n20603), .C2(n20233), .A(n20177), .B(n20176), .ZN(
        P1_U3041) );
  AOI22_X1 U23107 ( .A1(n20658), .A2(n20192), .B1(n20657), .B2(n20191), .ZN(
        n20179) );
  INV_X1 U23108 ( .A(n20233), .ZN(n20208) );
  INV_X1 U23109 ( .A(n20607), .ZN(n20660) );
  AOI22_X1 U23110 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20194), .B1(
        n20208), .B2(n20660), .ZN(n20178) );
  OAI211_X1 U23111 ( .C1(n20663), .C2(n20190), .A(n20179), .B(n20178), .ZN(
        P1_U3042) );
  AOI22_X1 U23112 ( .A1(n20665), .A2(n20192), .B1(n20664), .B2(n20191), .ZN(
        n20181) );
  INV_X1 U23113 ( .A(n20611), .ZN(n20666) );
  AOI22_X1 U23114 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20194), .B1(
        n20208), .B2(n20666), .ZN(n20180) );
  OAI211_X1 U23115 ( .C1(n20669), .C2(n20190), .A(n20181), .B(n20180), .ZN(
        P1_U3043) );
  AOI22_X1 U23116 ( .A1(n20671), .A2(n20192), .B1(n20670), .B2(n20191), .ZN(
        n20183) );
  INV_X1 U23117 ( .A(n20615), .ZN(n20672) );
  AOI22_X1 U23118 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20194), .B1(
        n20208), .B2(n20672), .ZN(n20182) );
  OAI211_X1 U23119 ( .C1(n20675), .C2(n20190), .A(n20183), .B(n20182), .ZN(
        P1_U3044) );
  AOI22_X1 U23120 ( .A1(n20677), .A2(n20192), .B1(n20676), .B2(n20191), .ZN(
        n20185) );
  AOI22_X1 U23121 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20194), .B1(
        n20193), .B2(n20616), .ZN(n20184) );
  OAI211_X1 U23122 ( .C1(n20619), .C2(n20233), .A(n20185), .B(n20184), .ZN(
        P1_U3045) );
  AOI22_X1 U23123 ( .A1(n20683), .A2(n20192), .B1(n20682), .B2(n20191), .ZN(
        n20187) );
  AOI22_X1 U23124 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20194), .B1(
        n20193), .B2(n20620), .ZN(n20186) );
  OAI211_X1 U23125 ( .C1(n20623), .C2(n20233), .A(n20187), .B(n20186), .ZN(
        P1_U3046) );
  AOI22_X1 U23126 ( .A1(n20689), .A2(n20192), .B1(n20688), .B2(n20191), .ZN(
        n20189) );
  INV_X1 U23127 ( .A(n20627), .ZN(n20690) );
  AOI22_X1 U23128 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20194), .B1(
        n20208), .B2(n20690), .ZN(n20188) );
  OAI211_X1 U23129 ( .C1(n20693), .C2(n20190), .A(n20189), .B(n20188), .ZN(
        P1_U3047) );
  AOI22_X1 U23130 ( .A1(n20697), .A2(n20192), .B1(n20695), .B2(n20191), .ZN(
        n20196) );
  AOI22_X1 U23131 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20194), .B1(
        n20193), .B2(n20630), .ZN(n20195) );
  OAI211_X1 U23132 ( .C1(n20635), .C2(n20233), .A(n20196), .B(n20195), .ZN(
        P1_U3048) );
  INV_X1 U23133 ( .A(n20591), .ZN(n20198) );
  NOR3_X1 U23134 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20638), .A3(
        n20237), .ZN(n20209) );
  INV_X1 U23135 ( .A(n20209), .ZN(n20227) );
  OAI22_X1 U23136 ( .A1(n20233), .A2(n20544), .B1(n20448), .B2(n20227), .ZN(
        n20199) );
  INV_X1 U23137 ( .A(n20199), .ZN(n20207) );
  AOI21_X1 U23138 ( .B1(n20269), .B2(n20233), .A(n20200), .ZN(n20201) );
  NOR2_X1 U23139 ( .A1(n20201), .A2(n20648), .ZN(n20203) );
  NAND2_X1 U23140 ( .A1(n9928), .A2(n20592), .ZN(n20204) );
  AOI22_X1 U23141 ( .A1(n20203), .A2(n20204), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20227), .ZN(n20202) );
  OR2_X1 U23142 ( .A1(n20454), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20337) );
  NAND2_X1 U23143 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20337), .ZN(n20334) );
  NAND3_X1 U23144 ( .A1(n20456), .A2(n20202), .A3(n20334), .ZN(n20230) );
  INV_X1 U23145 ( .A(n20203), .ZN(n20205) );
  AOI22_X1 U23146 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20230), .B1(
        n20651), .B2(n20229), .ZN(n20206) );
  OAI211_X1 U23147 ( .C1(n20603), .C2(n20269), .A(n20207), .B(n20206), .ZN(
        P1_U3049) );
  AOI22_X1 U23148 ( .A1(n20657), .A2(n20209), .B1(n20208), .B2(n20604), .ZN(
        n20211) );
  AOI22_X1 U23149 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20230), .B1(
        n20658), .B2(n20229), .ZN(n20210) );
  OAI211_X1 U23150 ( .C1(n20607), .C2(n20269), .A(n20211), .B(n20210), .ZN(
        P1_U3050) );
  INV_X1 U23151 ( .A(n20664), .ZN(n20467) );
  OAI22_X1 U23152 ( .A1(n20233), .A2(n20669), .B1(n20467), .B2(n20227), .ZN(
        n20212) );
  INV_X1 U23153 ( .A(n20212), .ZN(n20214) );
  AOI22_X1 U23154 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20230), .B1(
        n20665), .B2(n20229), .ZN(n20213) );
  OAI211_X1 U23155 ( .C1(n20611), .C2(n20269), .A(n20214), .B(n20213), .ZN(
        P1_U3051) );
  INV_X1 U23156 ( .A(n20670), .ZN(n20471) );
  OAI22_X1 U23157 ( .A1(n20269), .A2(n20615), .B1(n20471), .B2(n20227), .ZN(
        n20215) );
  INV_X1 U23158 ( .A(n20215), .ZN(n20217) );
  AOI22_X1 U23159 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20230), .B1(
        n20671), .B2(n20229), .ZN(n20216) );
  OAI211_X1 U23160 ( .C1(n20675), .C2(n20233), .A(n20217), .B(n20216), .ZN(
        P1_U3052) );
  OAI22_X1 U23161 ( .A1(n20233), .A2(n20681), .B1(n20475), .B2(n20227), .ZN(
        n20218) );
  INV_X1 U23162 ( .A(n20218), .ZN(n20220) );
  AOI22_X1 U23163 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20230), .B1(
        n20677), .B2(n20229), .ZN(n20219) );
  OAI211_X1 U23164 ( .C1(n20619), .C2(n20269), .A(n20220), .B(n20219), .ZN(
        P1_U3053) );
  INV_X1 U23165 ( .A(n20682), .ZN(n20479) );
  OAI22_X1 U23166 ( .A1(n20233), .A2(n20687), .B1(n20479), .B2(n20227), .ZN(
        n20221) );
  INV_X1 U23167 ( .A(n20221), .ZN(n20223) );
  AOI22_X1 U23168 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20230), .B1(
        n20683), .B2(n20229), .ZN(n20222) );
  OAI211_X1 U23169 ( .C1(n20623), .C2(n20269), .A(n20223), .B(n20222), .ZN(
        P1_U3054) );
  OAI22_X1 U23170 ( .A1(n20269), .A2(n20627), .B1(n20483), .B2(n20227), .ZN(
        n20224) );
  INV_X1 U23171 ( .A(n20224), .ZN(n20226) );
  AOI22_X1 U23172 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20230), .B1(
        n20689), .B2(n20229), .ZN(n20225) );
  OAI211_X1 U23173 ( .C1(n20693), .C2(n20233), .A(n20226), .B(n20225), .ZN(
        P1_U3055) );
  INV_X1 U23174 ( .A(n20695), .ZN(n20488) );
  OAI22_X1 U23175 ( .A1(n20269), .A2(n20635), .B1(n20488), .B2(n20227), .ZN(
        n20228) );
  INV_X1 U23176 ( .A(n20228), .ZN(n20232) );
  AOI22_X1 U23177 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20230), .B1(
        n20697), .B2(n20229), .ZN(n20231) );
  OAI211_X1 U23178 ( .C1(n20704), .C2(n20233), .A(n20232), .B(n20231), .ZN(
        P1_U3056) );
  INV_X1 U23179 ( .A(n20495), .ZN(n20234) );
  INV_X1 U23180 ( .A(n20237), .ZN(n20235) );
  AND2_X1 U23181 ( .A1(n20644), .A2(n20235), .ZN(n20250) );
  INV_X1 U23182 ( .A(n20250), .ZN(n20268) );
  OAI22_X1 U23183 ( .A1(n20269), .A2(n20544), .B1(n20448), .B2(n20268), .ZN(
        n20236) );
  INV_X1 U23184 ( .A(n20236), .ZN(n20249) );
  NOR2_X1 U23185 ( .A1(n20638), .A2(n20237), .ZN(n20244) );
  AND2_X1 U23186 ( .A1(n12524), .A2(n20238), .ZN(n20645) );
  AOI21_X1 U23187 ( .B1(n9928), .B2(n20645), .A(n20250), .ZN(n20247) );
  OR2_X1 U23188 ( .A1(n20239), .A2(n20502), .ZN(n20240) );
  AND2_X1 U23189 ( .A1(n20240), .A2(n20570), .ZN(n20243) );
  AOI21_X1 U23190 ( .B1(n20247), .B2(n20243), .A(n20241), .ZN(n20242) );
  OAI21_X1 U23191 ( .B1(n20570), .B2(n20244), .A(n20242), .ZN(n20272) );
  INV_X1 U23192 ( .A(n20243), .ZN(n20246) );
  INV_X1 U23193 ( .A(n20244), .ZN(n20245) );
  OAI22_X1 U23194 ( .A1(n20247), .A2(n20246), .B1(n20708), .B2(n20245), .ZN(
        n20271) );
  AOI22_X1 U23195 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20272), .B1(
        n20651), .B2(n20271), .ZN(n20248) );
  OAI211_X1 U23196 ( .C1(n20603), .C2(n20275), .A(n20249), .B(n20248), .ZN(
        P1_U3057) );
  AOI22_X1 U23197 ( .A1(n20250), .A2(n20657), .B1(n20301), .B2(n20660), .ZN(
        n20252) );
  AOI22_X1 U23198 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20272), .B1(
        n20658), .B2(n20271), .ZN(n20251) );
  OAI211_X1 U23199 ( .C1(n20663), .C2(n20269), .A(n20252), .B(n20251), .ZN(
        P1_U3058) );
  OAI22_X1 U23200 ( .A1(n20275), .A2(n20611), .B1(n20467), .B2(n20268), .ZN(
        n20253) );
  INV_X1 U23201 ( .A(n20253), .ZN(n20255) );
  AOI22_X1 U23202 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20272), .B1(
        n20665), .B2(n20271), .ZN(n20254) );
  OAI211_X1 U23203 ( .C1(n20669), .C2(n20269), .A(n20255), .B(n20254), .ZN(
        P1_U3059) );
  OAI22_X1 U23204 ( .A1(n20275), .A2(n20615), .B1(n20471), .B2(n20268), .ZN(
        n20256) );
  INV_X1 U23205 ( .A(n20256), .ZN(n20258) );
  AOI22_X1 U23206 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20272), .B1(
        n20671), .B2(n20271), .ZN(n20257) );
  OAI211_X1 U23207 ( .C1(n20675), .C2(n20269), .A(n20258), .B(n20257), .ZN(
        P1_U3060) );
  OAI22_X1 U23208 ( .A1(n20269), .A2(n20681), .B1(n20475), .B2(n20268), .ZN(
        n20259) );
  INV_X1 U23209 ( .A(n20259), .ZN(n20261) );
  AOI22_X1 U23210 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20272), .B1(
        n20677), .B2(n20271), .ZN(n20260) );
  OAI211_X1 U23211 ( .C1(n20619), .C2(n20275), .A(n20261), .B(n20260), .ZN(
        P1_U3061) );
  OAI22_X1 U23212 ( .A1(n20269), .A2(n20687), .B1(n20479), .B2(n20268), .ZN(
        n20262) );
  INV_X1 U23213 ( .A(n20262), .ZN(n20264) );
  AOI22_X1 U23214 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20272), .B1(
        n20683), .B2(n20271), .ZN(n20263) );
  OAI211_X1 U23215 ( .C1(n20623), .C2(n20275), .A(n20264), .B(n20263), .ZN(
        P1_U3062) );
  OAI22_X1 U23216 ( .A1(n20275), .A2(n20627), .B1(n20483), .B2(n20268), .ZN(
        n20265) );
  INV_X1 U23217 ( .A(n20265), .ZN(n20267) );
  AOI22_X1 U23218 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20272), .B1(
        n20689), .B2(n20271), .ZN(n20266) );
  OAI211_X1 U23219 ( .C1(n20693), .C2(n20269), .A(n20267), .B(n20266), .ZN(
        P1_U3063) );
  OAI22_X1 U23220 ( .A1(n20269), .A2(n20704), .B1(n20488), .B2(n20268), .ZN(
        n20270) );
  INV_X1 U23221 ( .A(n20270), .ZN(n20274) );
  AOI22_X1 U23222 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20272), .B1(
        n20697), .B2(n20271), .ZN(n20273) );
  OAI211_X1 U23223 ( .C1(n20635), .C2(n20275), .A(n20274), .B(n20273), .ZN(
        P1_U3064) );
  NOR2_X1 U23224 ( .A1(n20534), .A2(n20277), .ZN(n20368) );
  NAND3_X1 U23225 ( .A1(n20368), .A2(n20570), .A3(n20535), .ZN(n20278) );
  OAI21_X1 U23226 ( .B1(n20279), .B2(n20593), .A(n20278), .ZN(n20300) );
  AOI22_X1 U23227 ( .A1(n20651), .A2(n20300), .B1(n20650), .B2(n10300), .ZN(
        n20287) );
  INV_X1 U23228 ( .A(n20368), .ZN(n20282) );
  INV_X1 U23229 ( .A(n20330), .ZN(n20280) );
  OAI21_X1 U23230 ( .B1(n20301), .B2(n20280), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20281) );
  OAI21_X1 U23231 ( .B1(n20592), .B2(n20282), .A(n20281), .ZN(n20285) );
  INV_X1 U23232 ( .A(n20459), .ZN(n20283) );
  AOI22_X1 U23233 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20302), .B1(
        n20301), .B2(n20653), .ZN(n20286) );
  OAI211_X1 U23234 ( .C1(n20603), .C2(n20330), .A(n20287), .B(n20286), .ZN(
        P1_U3065) );
  AOI22_X1 U23235 ( .A1(n20658), .A2(n20300), .B1(n20657), .B2(n10300), .ZN(
        n20289) );
  AOI22_X1 U23236 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20302), .B1(
        n20301), .B2(n20604), .ZN(n20288) );
  OAI211_X1 U23237 ( .C1(n20607), .C2(n20330), .A(n20289), .B(n20288), .ZN(
        P1_U3066) );
  AOI22_X1 U23238 ( .A1(n20665), .A2(n20300), .B1(n20664), .B2(n10300), .ZN(
        n20291) );
  AOI22_X1 U23239 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20302), .B1(
        n20301), .B2(n20608), .ZN(n20290) );
  OAI211_X1 U23240 ( .C1(n20611), .C2(n20330), .A(n20291), .B(n20290), .ZN(
        P1_U3067) );
  AOI22_X1 U23241 ( .A1(n20671), .A2(n20300), .B1(n20670), .B2(n10300), .ZN(
        n20293) );
  AOI22_X1 U23242 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20302), .B1(
        n20301), .B2(n20612), .ZN(n20292) );
  OAI211_X1 U23243 ( .C1(n20615), .C2(n20330), .A(n20293), .B(n20292), .ZN(
        P1_U3068) );
  AOI22_X1 U23244 ( .A1(n20677), .A2(n20300), .B1(n20676), .B2(n10300), .ZN(
        n20295) );
  AOI22_X1 U23245 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20302), .B1(
        n20301), .B2(n20616), .ZN(n20294) );
  OAI211_X1 U23246 ( .C1(n20619), .C2(n20330), .A(n20295), .B(n20294), .ZN(
        P1_U3069) );
  AOI22_X1 U23247 ( .A1(n20683), .A2(n20300), .B1(n20682), .B2(n10300), .ZN(
        n20297) );
  AOI22_X1 U23248 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20302), .B1(
        n20301), .B2(n20620), .ZN(n20296) );
  OAI211_X1 U23249 ( .C1(n20623), .C2(n20330), .A(n20297), .B(n20296), .ZN(
        P1_U3070) );
  AOI22_X1 U23250 ( .A1(n20689), .A2(n20300), .B1(n20688), .B2(n10300), .ZN(
        n20299) );
  AOI22_X1 U23251 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20302), .B1(
        n20301), .B2(n20624), .ZN(n20298) );
  OAI211_X1 U23252 ( .C1(n20627), .C2(n20330), .A(n20299), .B(n20298), .ZN(
        P1_U3071) );
  AOI22_X1 U23253 ( .A1(n20697), .A2(n20300), .B1(n20695), .B2(n10300), .ZN(
        n20304) );
  AOI22_X1 U23254 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20302), .B1(
        n20301), .B2(n20630), .ZN(n20303) );
  OAI211_X1 U23255 ( .C1(n20635), .C2(n20330), .A(n20304), .B(n20303), .ZN(
        P1_U3072) );
  NOR2_X1 U23256 ( .A1(n20331), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20308) );
  INV_X1 U23257 ( .A(n20308), .ZN(n20305) );
  NOR2_X1 U23258 ( .A1(n20563), .A2(n20305), .ZN(n20325) );
  AOI21_X1 U23259 ( .B1(n20368), .B2(n20564), .A(n20325), .ZN(n20306) );
  OAI22_X1 U23260 ( .A1(n20306), .A2(n20648), .B1(n20305), .B2(n20708), .ZN(
        n20326) );
  AOI22_X1 U23261 ( .A1(n20651), .A2(n20326), .B1(n20650), .B2(n20325), .ZN(
        n20312) );
  INV_X1 U23262 ( .A(n20374), .ZN(n20307) );
  NOR3_X1 U23263 ( .A1(n20307), .A2(n20648), .A3(n20425), .ZN(n20309) );
  OAI21_X1 U23264 ( .B1(n20309), .B2(n20308), .A(n20640), .ZN(n20327) );
  NAND2_X1 U23265 ( .A1(n20374), .A2(n20562), .ZN(n20362) );
  INV_X1 U23266 ( .A(n20603), .ZN(n20652) );
  AOI22_X1 U23267 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20327), .B1(
        n20342), .B2(n20652), .ZN(n20311) );
  OAI211_X1 U23268 ( .C1(n20544), .C2(n20330), .A(n20312), .B(n20311), .ZN(
        P1_U3073) );
  AOI22_X1 U23269 ( .A1(n20658), .A2(n20326), .B1(n20657), .B2(n20325), .ZN(
        n20314) );
  AOI22_X1 U23270 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20327), .B1(
        n20342), .B2(n20660), .ZN(n20313) );
  OAI211_X1 U23271 ( .C1(n20663), .C2(n20330), .A(n20314), .B(n20313), .ZN(
        P1_U3074) );
  AOI22_X1 U23272 ( .A1(n20665), .A2(n20326), .B1(n20664), .B2(n20325), .ZN(
        n20316) );
  AOI22_X1 U23273 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20327), .B1(
        n20342), .B2(n20666), .ZN(n20315) );
  OAI211_X1 U23274 ( .C1(n20669), .C2(n20330), .A(n20316), .B(n20315), .ZN(
        P1_U3075) );
  AOI22_X1 U23275 ( .A1(n20671), .A2(n20326), .B1(n20670), .B2(n20325), .ZN(
        n20318) );
  AOI22_X1 U23276 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20327), .B1(
        n20342), .B2(n20672), .ZN(n20317) );
  OAI211_X1 U23277 ( .C1(n20675), .C2(n20330), .A(n20318), .B(n20317), .ZN(
        P1_U3076) );
  AOI22_X1 U23278 ( .A1(n20677), .A2(n20326), .B1(n20676), .B2(n20325), .ZN(
        n20320) );
  INV_X1 U23279 ( .A(n20619), .ZN(n20678) );
  AOI22_X1 U23280 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20327), .B1(
        n20342), .B2(n20678), .ZN(n20319) );
  OAI211_X1 U23281 ( .C1(n20681), .C2(n20330), .A(n20320), .B(n20319), .ZN(
        P1_U3077) );
  AOI22_X1 U23282 ( .A1(n20683), .A2(n20326), .B1(n20682), .B2(n20325), .ZN(
        n20322) );
  INV_X1 U23283 ( .A(n20623), .ZN(n20684) );
  AOI22_X1 U23284 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20327), .B1(
        n20342), .B2(n20684), .ZN(n20321) );
  OAI211_X1 U23285 ( .C1(n20687), .C2(n20330), .A(n20322), .B(n20321), .ZN(
        P1_U3078) );
  AOI22_X1 U23286 ( .A1(n20689), .A2(n20326), .B1(n20688), .B2(n20325), .ZN(
        n20324) );
  AOI22_X1 U23287 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20327), .B1(
        n20342), .B2(n20690), .ZN(n20323) );
  OAI211_X1 U23288 ( .C1(n20693), .C2(n20330), .A(n20324), .B(n20323), .ZN(
        P1_U3079) );
  AOI22_X1 U23289 ( .A1(n20697), .A2(n20326), .B1(n20695), .B2(n20325), .ZN(
        n20329) );
  INV_X1 U23290 ( .A(n20635), .ZN(n20698) );
  AOI22_X1 U23291 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20327), .B1(
        n20342), .B2(n20698), .ZN(n20328) );
  OAI211_X1 U23292 ( .C1(n20704), .C2(n20330), .A(n20329), .B(n20328), .ZN(
        P1_U3080) );
  NOR2_X1 U23293 ( .A1(n20638), .A2(n20331), .ZN(n20373) );
  INV_X1 U23294 ( .A(n20373), .ZN(n20369) );
  NOR2_X1 U23295 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20369), .ZN(
        n20343) );
  INV_X1 U23296 ( .A(n20343), .ZN(n20361) );
  OAI22_X1 U23297 ( .A1(n20362), .A2(n20544), .B1(n20448), .B2(n20361), .ZN(
        n20332) );
  INV_X1 U23298 ( .A(n20332), .ZN(n20341) );
  NAND3_X1 U23299 ( .A1(n20396), .A2(n20362), .A3(n20570), .ZN(n20333) );
  NAND2_X1 U23300 ( .A1(n20333), .A2(n20531), .ZN(n20336) );
  NAND2_X1 U23301 ( .A1(n20368), .A2(n20592), .ZN(n20338) );
  AOI22_X1 U23302 ( .A1(n20336), .A2(n20338), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20361), .ZN(n20335) );
  NAND3_X1 U23303 ( .A1(n20599), .A2(n20335), .A3(n20334), .ZN(n20365) );
  INV_X1 U23304 ( .A(n20336), .ZN(n20339) );
  OAI22_X1 U23305 ( .A1(n20339), .A2(n20338), .B1(n20337), .B2(n20593), .ZN(
        n20364) );
  AOI22_X1 U23306 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20365), .B1(
        n20651), .B2(n20364), .ZN(n20340) );
  OAI211_X1 U23307 ( .C1(n20603), .C2(n20396), .A(n20341), .B(n20340), .ZN(
        P1_U3081) );
  AOI22_X1 U23308 ( .A1(n20657), .A2(n20343), .B1(n20342), .B2(n20604), .ZN(
        n20345) );
  AOI22_X1 U23309 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20365), .B1(
        n20658), .B2(n20364), .ZN(n20344) );
  OAI211_X1 U23310 ( .C1(n20607), .C2(n20396), .A(n20345), .B(n20344), .ZN(
        P1_U3082) );
  OAI22_X1 U23311 ( .A1(n20396), .A2(n20611), .B1(n20467), .B2(n20361), .ZN(
        n20346) );
  INV_X1 U23312 ( .A(n20346), .ZN(n20348) );
  AOI22_X1 U23313 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20365), .B1(
        n20665), .B2(n20364), .ZN(n20347) );
  OAI211_X1 U23314 ( .C1(n20669), .C2(n20362), .A(n20348), .B(n20347), .ZN(
        P1_U3083) );
  OAI22_X1 U23315 ( .A1(n20396), .A2(n20615), .B1(n20471), .B2(n20361), .ZN(
        n20349) );
  INV_X1 U23316 ( .A(n20349), .ZN(n20351) );
  AOI22_X1 U23317 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20365), .B1(
        n20671), .B2(n20364), .ZN(n20350) );
  OAI211_X1 U23318 ( .C1(n20675), .C2(n20362), .A(n20351), .B(n20350), .ZN(
        P1_U3084) );
  OAI22_X1 U23319 ( .A1(n20396), .A2(n20619), .B1(n20475), .B2(n20361), .ZN(
        n20352) );
  INV_X1 U23320 ( .A(n20352), .ZN(n20354) );
  AOI22_X1 U23321 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20365), .B1(
        n20677), .B2(n20364), .ZN(n20353) );
  OAI211_X1 U23322 ( .C1(n20681), .C2(n20362), .A(n20354), .B(n20353), .ZN(
        P1_U3085) );
  OAI22_X1 U23323 ( .A1(n20362), .A2(n20687), .B1(n20479), .B2(n20361), .ZN(
        n20355) );
  INV_X1 U23324 ( .A(n20355), .ZN(n20357) );
  AOI22_X1 U23325 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20365), .B1(
        n20683), .B2(n20364), .ZN(n20356) );
  OAI211_X1 U23326 ( .C1(n20623), .C2(n20396), .A(n20357), .B(n20356), .ZN(
        P1_U3086) );
  OAI22_X1 U23327 ( .A1(n20396), .A2(n20627), .B1(n20483), .B2(n20361), .ZN(
        n20358) );
  INV_X1 U23328 ( .A(n20358), .ZN(n20360) );
  AOI22_X1 U23329 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20365), .B1(
        n20689), .B2(n20364), .ZN(n20359) );
  OAI211_X1 U23330 ( .C1(n20693), .C2(n20362), .A(n20360), .B(n20359), .ZN(
        P1_U3087) );
  OAI22_X1 U23331 ( .A1(n20362), .A2(n20704), .B1(n20488), .B2(n20361), .ZN(
        n20363) );
  INV_X1 U23332 ( .A(n20363), .ZN(n20367) );
  AOI22_X1 U23333 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20365), .B1(
        n20697), .B2(n20364), .ZN(n20366) );
  OAI211_X1 U23334 ( .C1(n20635), .C2(n20396), .A(n20367), .B(n20366), .ZN(
        P1_U3088) );
  AOI21_X1 U23335 ( .B1(n20368), .B2(n20645), .A(n20391), .ZN(n20370) );
  OAI22_X1 U23336 ( .A1(n20370), .A2(n20648), .B1(n20369), .B2(n20708), .ZN(
        n20392) );
  AOI22_X1 U23337 ( .A1(n20651), .A2(n20392), .B1(n20391), .B2(n20650), .ZN(
        n20376) );
  NAND2_X1 U23338 ( .A1(n20371), .A2(n20370), .ZN(n20372) );
  OAI221_X1 U23339 ( .B1(n20570), .B2(n20373), .C1(n20648), .C2(n20372), .A(
        n20640), .ZN(n20393) );
  NAND2_X1 U23340 ( .A1(n20374), .A2(n20495), .ZN(n20384) );
  AOI22_X1 U23341 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20393), .B1(
        n20419), .B2(n20652), .ZN(n20375) );
  OAI211_X1 U23342 ( .C1(n20544), .C2(n20396), .A(n20376), .B(n20375), .ZN(
        P1_U3089) );
  AOI22_X1 U23343 ( .A1(n20391), .A2(n20657), .B1(n20658), .B2(n20392), .ZN(
        n20378) );
  AOI22_X1 U23344 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20393), .B1(
        n20419), .B2(n20660), .ZN(n20377) );
  OAI211_X1 U23345 ( .C1(n20663), .C2(n20396), .A(n20378), .B(n20377), .ZN(
        P1_U3090) );
  AOI22_X1 U23346 ( .A1(n20665), .A2(n20392), .B1(n20391), .B2(n20664), .ZN(
        n20380) );
  AOI22_X1 U23347 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20393), .B1(
        n20419), .B2(n20666), .ZN(n20379) );
  OAI211_X1 U23348 ( .C1(n20669), .C2(n20396), .A(n20380), .B(n20379), .ZN(
        P1_U3091) );
  AOI22_X1 U23349 ( .A1(n20671), .A2(n20392), .B1(n20391), .B2(n20670), .ZN(
        n20383) );
  INV_X1 U23350 ( .A(n20396), .ZN(n20381) );
  AOI22_X1 U23351 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20393), .B1(
        n20381), .B2(n20612), .ZN(n20382) );
  OAI211_X1 U23352 ( .C1(n20615), .C2(n20384), .A(n20383), .B(n20382), .ZN(
        P1_U3092) );
  AOI22_X1 U23353 ( .A1(n20677), .A2(n20392), .B1(n20391), .B2(n20676), .ZN(
        n20386) );
  AOI22_X1 U23354 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20393), .B1(
        n20419), .B2(n20678), .ZN(n20385) );
  OAI211_X1 U23355 ( .C1(n20681), .C2(n20396), .A(n20386), .B(n20385), .ZN(
        P1_U3093) );
  AOI22_X1 U23356 ( .A1(n20683), .A2(n20392), .B1(n20391), .B2(n20682), .ZN(
        n20388) );
  AOI22_X1 U23357 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20393), .B1(
        n20419), .B2(n20684), .ZN(n20387) );
  OAI211_X1 U23358 ( .C1(n20687), .C2(n20396), .A(n20388), .B(n20387), .ZN(
        P1_U3094) );
  AOI22_X1 U23359 ( .A1(n20689), .A2(n20392), .B1(n20391), .B2(n20688), .ZN(
        n20390) );
  AOI22_X1 U23360 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20393), .B1(
        n20419), .B2(n20690), .ZN(n20389) );
  OAI211_X1 U23361 ( .C1(n20693), .C2(n20396), .A(n20390), .B(n20389), .ZN(
        P1_U3095) );
  AOI22_X1 U23362 ( .A1(n20697), .A2(n20392), .B1(n20391), .B2(n20695), .ZN(
        n20395) );
  AOI22_X1 U23363 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20393), .B1(
        n20419), .B2(n20698), .ZN(n20394) );
  OAI211_X1 U23364 ( .C1(n20704), .C2(n20396), .A(n20395), .B(n20394), .ZN(
        P1_U3096) );
  NAND2_X1 U23365 ( .A1(n20397), .A2(n20534), .ZN(n20452) );
  INV_X1 U23366 ( .A(n20452), .ZN(n20499) );
  NAND2_X1 U23367 ( .A1(n20398), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20497) );
  AOI21_X1 U23368 ( .B1(n20499), .B2(n20535), .A(n10305), .ZN(n20401) );
  NAND2_X1 U23369 ( .A1(n20399), .A2(n20454), .ZN(n20539) );
  OAI22_X1 U23370 ( .A1(n20401), .A2(n20648), .B1(n20459), .B2(n20539), .ZN(
        n20418) );
  AOI22_X1 U23371 ( .A1(n20651), .A2(n20418), .B1(n10305), .B2(n20650), .ZN(
        n20405) );
  INV_X1 U23372 ( .A(n20447), .ZN(n20400) );
  OAI21_X1 U23373 ( .B1(n20400), .B2(n20419), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20402) );
  NAND2_X1 U23374 ( .A1(n20402), .A2(n20401), .ZN(n20403) );
  AOI22_X1 U23375 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20420), .B1(
        n20419), .B2(n20653), .ZN(n20404) );
  OAI211_X1 U23376 ( .C1(n20603), .C2(n20447), .A(n20405), .B(n20404), .ZN(
        P1_U3097) );
  AOI22_X1 U23377 ( .A1(n20658), .A2(n20418), .B1(n20657), .B2(n10305), .ZN(
        n20407) );
  AOI22_X1 U23378 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20420), .B1(
        n20419), .B2(n20604), .ZN(n20406) );
  OAI211_X1 U23379 ( .C1(n20607), .C2(n20447), .A(n20407), .B(n20406), .ZN(
        P1_U3098) );
  AOI22_X1 U23380 ( .A1(n20665), .A2(n20418), .B1(n10305), .B2(n20664), .ZN(
        n20409) );
  AOI22_X1 U23381 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20420), .B1(
        n20419), .B2(n20608), .ZN(n20408) );
  OAI211_X1 U23382 ( .C1(n20611), .C2(n20447), .A(n20409), .B(n20408), .ZN(
        P1_U3099) );
  AOI22_X1 U23383 ( .A1(n20671), .A2(n20418), .B1(n10305), .B2(n20670), .ZN(
        n20411) );
  AOI22_X1 U23384 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20420), .B1(
        n20419), .B2(n20612), .ZN(n20410) );
  OAI211_X1 U23385 ( .C1(n20615), .C2(n20447), .A(n20411), .B(n20410), .ZN(
        P1_U3100) );
  AOI22_X1 U23386 ( .A1(n20677), .A2(n20418), .B1(n10305), .B2(n20676), .ZN(
        n20413) );
  AOI22_X1 U23387 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20420), .B1(
        n20419), .B2(n20616), .ZN(n20412) );
  OAI211_X1 U23388 ( .C1(n20619), .C2(n20447), .A(n20413), .B(n20412), .ZN(
        P1_U3101) );
  AOI22_X1 U23389 ( .A1(n20683), .A2(n20418), .B1(n10305), .B2(n20682), .ZN(
        n20415) );
  AOI22_X1 U23390 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20420), .B1(
        n20419), .B2(n20620), .ZN(n20414) );
  OAI211_X1 U23391 ( .C1(n20623), .C2(n20447), .A(n20415), .B(n20414), .ZN(
        P1_U3102) );
  AOI22_X1 U23392 ( .A1(n20689), .A2(n20418), .B1(n10305), .B2(n20688), .ZN(
        n20417) );
  AOI22_X1 U23393 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20420), .B1(
        n20419), .B2(n20624), .ZN(n20416) );
  OAI211_X1 U23394 ( .C1(n20627), .C2(n20447), .A(n20417), .B(n20416), .ZN(
        P1_U3103) );
  AOI22_X1 U23395 ( .A1(n20697), .A2(n20418), .B1(n10305), .B2(n20695), .ZN(
        n20422) );
  AOI22_X1 U23396 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20420), .B1(
        n20419), .B2(n20630), .ZN(n20421) );
  OAI211_X1 U23397 ( .C1(n20635), .C2(n20447), .A(n20422), .B(n20421), .ZN(
        P1_U3104) );
  NOR2_X1 U23398 ( .A1(n20497), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20427) );
  INV_X1 U23399 ( .A(n20427), .ZN(n20423) );
  NOR2_X1 U23400 ( .A1(n20563), .A2(n20423), .ZN(n20442) );
  AOI21_X1 U23401 ( .B1(n20499), .B2(n20564), .A(n20442), .ZN(n20424) );
  OAI22_X1 U23402 ( .A1(n20424), .A2(n20648), .B1(n20423), .B2(n20708), .ZN(
        n20443) );
  AOI22_X1 U23403 ( .A1(n20651), .A2(n20443), .B1(n20650), .B2(n20442), .ZN(
        n20429) );
  OAI211_X1 U23404 ( .C1(n20503), .C2(n20425), .A(n20570), .B(n20424), .ZN(
        n20426) );
  OAI211_X1 U23405 ( .C1(n20570), .C2(n20427), .A(n20640), .B(n20426), .ZN(
        n20444) );
  AOI22_X1 U23406 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20444), .B1(
        n20450), .B2(n20652), .ZN(n20428) );
  OAI211_X1 U23407 ( .C1(n20544), .C2(n20447), .A(n20429), .B(n20428), .ZN(
        P1_U3105) );
  AOI22_X1 U23408 ( .A1(n20658), .A2(n20443), .B1(n20657), .B2(n20442), .ZN(
        n20431) );
  AOI22_X1 U23409 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20444), .B1(
        n20450), .B2(n20660), .ZN(n20430) );
  OAI211_X1 U23410 ( .C1(n20663), .C2(n20447), .A(n20431), .B(n20430), .ZN(
        P1_U3106) );
  AOI22_X1 U23411 ( .A1(n20665), .A2(n20443), .B1(n20664), .B2(n20442), .ZN(
        n20433) );
  AOI22_X1 U23412 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20444), .B1(
        n20450), .B2(n20666), .ZN(n20432) );
  OAI211_X1 U23413 ( .C1(n20669), .C2(n20447), .A(n20433), .B(n20432), .ZN(
        P1_U3107) );
  AOI22_X1 U23414 ( .A1(n20671), .A2(n20443), .B1(n20670), .B2(n20442), .ZN(
        n20435) );
  AOI22_X1 U23415 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20444), .B1(
        n20450), .B2(n20672), .ZN(n20434) );
  OAI211_X1 U23416 ( .C1(n20675), .C2(n20447), .A(n20435), .B(n20434), .ZN(
        P1_U3108) );
  AOI22_X1 U23417 ( .A1(n20677), .A2(n20443), .B1(n20676), .B2(n20442), .ZN(
        n20437) );
  AOI22_X1 U23418 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20444), .B1(
        n20450), .B2(n20678), .ZN(n20436) );
  OAI211_X1 U23419 ( .C1(n20681), .C2(n20447), .A(n20437), .B(n20436), .ZN(
        P1_U3109) );
  AOI22_X1 U23420 ( .A1(n20683), .A2(n20443), .B1(n20682), .B2(n20442), .ZN(
        n20439) );
  AOI22_X1 U23421 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20444), .B1(
        n20450), .B2(n20684), .ZN(n20438) );
  OAI211_X1 U23422 ( .C1(n20687), .C2(n20447), .A(n20439), .B(n20438), .ZN(
        P1_U3110) );
  AOI22_X1 U23423 ( .A1(n20689), .A2(n20443), .B1(n20688), .B2(n20442), .ZN(
        n20441) );
  AOI22_X1 U23424 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20444), .B1(
        n20450), .B2(n20690), .ZN(n20440) );
  OAI211_X1 U23425 ( .C1(n20693), .C2(n20447), .A(n20441), .B(n20440), .ZN(
        P1_U3111) );
  AOI22_X1 U23426 ( .A1(n20697), .A2(n20443), .B1(n20695), .B2(n20442), .ZN(
        n20446) );
  AOI22_X1 U23427 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20444), .B1(
        n20450), .B2(n20698), .ZN(n20445) );
  OAI211_X1 U23428 ( .C1(n20704), .C2(n20447), .A(n20446), .B(n20445), .ZN(
        P1_U3112) );
  NOR2_X1 U23429 ( .A1(n20638), .A2(n20497), .ZN(n20505) );
  INV_X1 U23430 ( .A(n20505), .ZN(n20500) );
  NOR2_X1 U23431 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20500), .ZN(
        n20464) );
  INV_X1 U23432 ( .A(n20464), .ZN(n20487) );
  OAI22_X1 U23433 ( .A1(n20494), .A2(n20544), .B1(n20448), .B2(n20487), .ZN(
        n20449) );
  INV_X1 U23434 ( .A(n20449), .ZN(n20463) );
  OAI21_X1 U23435 ( .B1(n20512), .B2(n20450), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20451) );
  NAND2_X1 U23436 ( .A1(n20451), .A2(n20570), .ZN(n20461) );
  NOR2_X1 U23437 ( .A1(n20452), .A2(n20535), .ZN(n20458) );
  OR2_X1 U23438 ( .A1(n20454), .A2(n20453), .ZN(n20594) );
  NAND2_X1 U23439 ( .A1(n20594), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20598) );
  OAI21_X1 U23440 ( .B1(n20537), .B2(n20464), .A(n20598), .ZN(n20455) );
  INV_X1 U23441 ( .A(n20455), .ZN(n20457) );
  OAI211_X1 U23442 ( .C1(n20461), .C2(n20458), .A(n20457), .B(n20456), .ZN(
        n20491) );
  INV_X1 U23443 ( .A(n20458), .ZN(n20460) );
  AOI22_X1 U23444 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20491), .B1(
        n20651), .B2(n20490), .ZN(n20462) );
  OAI211_X1 U23445 ( .C1(n20603), .C2(n20527), .A(n20463), .B(n20462), .ZN(
        P1_U3113) );
  AOI22_X1 U23446 ( .A1(n20464), .A2(n20657), .B1(n20512), .B2(n20660), .ZN(
        n20466) );
  AOI22_X1 U23447 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20491), .B1(
        n20658), .B2(n20490), .ZN(n20465) );
  OAI211_X1 U23448 ( .C1(n20663), .C2(n20494), .A(n20466), .B(n20465), .ZN(
        P1_U3114) );
  OAI22_X1 U23449 ( .A1(n20527), .A2(n20611), .B1(n20467), .B2(n20487), .ZN(
        n20468) );
  INV_X1 U23450 ( .A(n20468), .ZN(n20470) );
  AOI22_X1 U23451 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20491), .B1(
        n20665), .B2(n20490), .ZN(n20469) );
  OAI211_X1 U23452 ( .C1(n20669), .C2(n20494), .A(n20470), .B(n20469), .ZN(
        P1_U3115) );
  OAI22_X1 U23453 ( .A1(n20494), .A2(n20675), .B1(n20471), .B2(n20487), .ZN(
        n20472) );
  INV_X1 U23454 ( .A(n20472), .ZN(n20474) );
  AOI22_X1 U23455 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20491), .B1(
        n20671), .B2(n20490), .ZN(n20473) );
  OAI211_X1 U23456 ( .C1(n20615), .C2(n20527), .A(n20474), .B(n20473), .ZN(
        P1_U3116) );
  OAI22_X1 U23457 ( .A1(n20494), .A2(n20681), .B1(n20475), .B2(n20487), .ZN(
        n20476) );
  INV_X1 U23458 ( .A(n20476), .ZN(n20478) );
  AOI22_X1 U23459 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20491), .B1(
        n20677), .B2(n20490), .ZN(n20477) );
  OAI211_X1 U23460 ( .C1(n20619), .C2(n20527), .A(n20478), .B(n20477), .ZN(
        P1_U3117) );
  OAI22_X1 U23461 ( .A1(n20527), .A2(n20623), .B1(n20479), .B2(n20487), .ZN(
        n20480) );
  INV_X1 U23462 ( .A(n20480), .ZN(n20482) );
  AOI22_X1 U23463 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20491), .B1(
        n20683), .B2(n20490), .ZN(n20481) );
  OAI211_X1 U23464 ( .C1(n20687), .C2(n20494), .A(n20482), .B(n20481), .ZN(
        P1_U3118) );
  OAI22_X1 U23465 ( .A1(n20494), .A2(n20693), .B1(n20483), .B2(n20487), .ZN(
        n20484) );
  INV_X1 U23466 ( .A(n20484), .ZN(n20486) );
  AOI22_X1 U23467 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20491), .B1(
        n20689), .B2(n20490), .ZN(n20485) );
  OAI211_X1 U23468 ( .C1(n20627), .C2(n20527), .A(n20486), .B(n20485), .ZN(
        P1_U3119) );
  OAI22_X1 U23469 ( .A1(n20527), .A2(n20635), .B1(n20488), .B2(n20487), .ZN(
        n20489) );
  INV_X1 U23470 ( .A(n20489), .ZN(n20493) );
  AOI22_X1 U23471 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20491), .B1(
        n20697), .B2(n20490), .ZN(n20492) );
  OAI211_X1 U23472 ( .C1(n20704), .C2(n20494), .A(n20493), .B(n20492), .ZN(
        P1_U3120) );
  INV_X1 U23473 ( .A(n20497), .ZN(n20498) );
  AND2_X1 U23474 ( .A1(n20644), .A2(n20498), .ZN(n20521) );
  AOI21_X1 U23475 ( .B1(n20499), .B2(n20645), .A(n20521), .ZN(n20501) );
  OAI22_X1 U23476 ( .A1(n20501), .A2(n20648), .B1(n20500), .B2(n20708), .ZN(
        n20522) );
  AOI22_X1 U23477 ( .A1(n20651), .A2(n20522), .B1(n20650), .B2(n20521), .ZN(
        n20507) );
  OAI211_X1 U23478 ( .C1(n20503), .C2(n20502), .A(n20570), .B(n20501), .ZN(
        n20504) );
  OAI211_X1 U23479 ( .C1(n20570), .C2(n20505), .A(n20640), .B(n20504), .ZN(
        n20524) );
  AOI22_X1 U23480 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20524), .B1(
        n20512), .B2(n20653), .ZN(n20506) );
  OAI211_X1 U23481 ( .C1(n20603), .C2(n20561), .A(n20507), .B(n20506), .ZN(
        P1_U3121) );
  AOI22_X1 U23482 ( .A1(n20658), .A2(n20522), .B1(n20657), .B2(n20521), .ZN(
        n20509) );
  INV_X1 U23483 ( .A(n20561), .ZN(n20523) );
  AOI22_X1 U23484 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20524), .B1(
        n20523), .B2(n20660), .ZN(n20508) );
  OAI211_X1 U23485 ( .C1(n20663), .C2(n20527), .A(n20509), .B(n20508), .ZN(
        P1_U3122) );
  AOI22_X1 U23486 ( .A1(n20665), .A2(n20522), .B1(n20664), .B2(n20521), .ZN(
        n20511) );
  AOI22_X1 U23487 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20524), .B1(
        n20523), .B2(n20666), .ZN(n20510) );
  OAI211_X1 U23488 ( .C1(n20669), .C2(n20527), .A(n20511), .B(n20510), .ZN(
        P1_U3123) );
  AOI22_X1 U23489 ( .A1(n20671), .A2(n20522), .B1(n20670), .B2(n20521), .ZN(
        n20514) );
  AOI22_X1 U23490 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20524), .B1(
        n20512), .B2(n20612), .ZN(n20513) );
  OAI211_X1 U23491 ( .C1(n20615), .C2(n20561), .A(n20514), .B(n20513), .ZN(
        P1_U3124) );
  AOI22_X1 U23492 ( .A1(n20677), .A2(n20522), .B1(n20676), .B2(n20521), .ZN(
        n20516) );
  AOI22_X1 U23493 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20524), .B1(
        n20523), .B2(n20678), .ZN(n20515) );
  OAI211_X1 U23494 ( .C1(n20681), .C2(n20527), .A(n20516), .B(n20515), .ZN(
        P1_U3125) );
  AOI22_X1 U23495 ( .A1(n20683), .A2(n20522), .B1(n20682), .B2(n20521), .ZN(
        n20518) );
  AOI22_X1 U23496 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20524), .B1(
        n20523), .B2(n20684), .ZN(n20517) );
  OAI211_X1 U23497 ( .C1(n20687), .C2(n20527), .A(n20518), .B(n20517), .ZN(
        P1_U3126) );
  AOI22_X1 U23498 ( .A1(n20689), .A2(n20522), .B1(n20688), .B2(n20521), .ZN(
        n20520) );
  AOI22_X1 U23499 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20524), .B1(
        n20523), .B2(n20690), .ZN(n20519) );
  OAI211_X1 U23500 ( .C1(n20693), .C2(n20527), .A(n20520), .B(n20519), .ZN(
        P1_U3127) );
  AOI22_X1 U23501 ( .A1(n20697), .A2(n20522), .B1(n20695), .B2(n20521), .ZN(
        n20526) );
  AOI22_X1 U23502 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20524), .B1(
        n20523), .B2(n20698), .ZN(n20525) );
  OAI211_X1 U23503 ( .C1(n20704), .C2(n20527), .A(n20526), .B(n20525), .ZN(
        P1_U3128) );
  NAND2_X1 U23504 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20642) );
  AOI22_X1 U23505 ( .A1(n20587), .A2(n20652), .B1(n20650), .B2(n10299), .ZN(
        n20543) );
  INV_X1 U23506 ( .A(n20587), .ZN(n20530) );
  NAND3_X1 U23507 ( .A1(n20561), .A2(n20530), .A3(n20570), .ZN(n20532) );
  NAND2_X1 U23508 ( .A1(n20532), .A2(n20531), .ZN(n20538) );
  NOR2_X1 U23509 ( .A1(n20534), .A2(n20533), .ZN(n20646) );
  NAND2_X1 U23510 ( .A1(n20646), .A2(n20535), .ZN(n20540) );
  AOI22_X1 U23511 ( .A1(n20538), .A2(n20540), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20539), .ZN(n20536) );
  OAI211_X1 U23512 ( .C1(n10299), .C2(n20537), .A(n20599), .B(n20536), .ZN(
        n20558) );
  INV_X1 U23513 ( .A(n20538), .ZN(n20541) );
  OAI22_X1 U23514 ( .A1(n20541), .A2(n20540), .B1(n20593), .B2(n20539), .ZN(
        n20557) );
  AOI22_X1 U23515 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20558), .B1(
        n20651), .B2(n20557), .ZN(n20542) );
  OAI211_X1 U23516 ( .C1(n20544), .C2(n20561), .A(n20543), .B(n20542), .ZN(
        P1_U3129) );
  AOI22_X1 U23517 ( .A1(n10299), .A2(n20657), .B1(n20587), .B2(n20660), .ZN(
        n20546) );
  AOI22_X1 U23518 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20558), .B1(
        n20658), .B2(n20557), .ZN(n20545) );
  OAI211_X1 U23519 ( .C1(n20663), .C2(n20561), .A(n20546), .B(n20545), .ZN(
        P1_U3130) );
  AOI22_X1 U23520 ( .A1(n20587), .A2(n20666), .B1(n20664), .B2(n10299), .ZN(
        n20548) );
  AOI22_X1 U23521 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20558), .B1(
        n20665), .B2(n20557), .ZN(n20547) );
  OAI211_X1 U23522 ( .C1(n20669), .C2(n20561), .A(n20548), .B(n20547), .ZN(
        P1_U3131) );
  AOI22_X1 U23523 ( .A1(n20587), .A2(n20672), .B1(n20670), .B2(n10299), .ZN(
        n20550) );
  AOI22_X1 U23524 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20558), .B1(
        n20671), .B2(n20557), .ZN(n20549) );
  OAI211_X1 U23525 ( .C1(n20675), .C2(n20561), .A(n20550), .B(n20549), .ZN(
        P1_U3132) );
  AOI22_X1 U23526 ( .A1(n20587), .A2(n20678), .B1(n20676), .B2(n10299), .ZN(
        n20552) );
  AOI22_X1 U23527 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20558), .B1(
        n20677), .B2(n20557), .ZN(n20551) );
  OAI211_X1 U23528 ( .C1(n20681), .C2(n20561), .A(n20552), .B(n20551), .ZN(
        P1_U3133) );
  AOI22_X1 U23529 ( .A1(n20587), .A2(n20684), .B1(n20682), .B2(n10299), .ZN(
        n20554) );
  AOI22_X1 U23530 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20558), .B1(
        n20683), .B2(n20557), .ZN(n20553) );
  OAI211_X1 U23531 ( .C1(n20687), .C2(n20561), .A(n20554), .B(n20553), .ZN(
        P1_U3134) );
  AOI22_X1 U23532 ( .A1(n20587), .A2(n20690), .B1(n20688), .B2(n10299), .ZN(
        n20556) );
  AOI22_X1 U23533 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20558), .B1(
        n20689), .B2(n20557), .ZN(n20555) );
  OAI211_X1 U23534 ( .C1(n20693), .C2(n20561), .A(n20556), .B(n20555), .ZN(
        P1_U3135) );
  AOI22_X1 U23535 ( .A1(n20587), .A2(n20698), .B1(n20695), .B2(n10299), .ZN(
        n20560) );
  AOI22_X1 U23536 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20558), .B1(
        n20697), .B2(n20557), .ZN(n20559) );
  OAI211_X1 U23537 ( .C1(n20704), .C2(n20561), .A(n20560), .B(n20559), .ZN(
        P1_U3136) );
  NOR3_X2 U23538 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20563), .A3(
        n20642), .ZN(n20585) );
  AOI21_X1 U23539 ( .B1(n20646), .B2(n20564), .A(n20585), .ZN(n20566) );
  NOR2_X1 U23540 ( .A1(n20642), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20569) );
  INV_X1 U23541 ( .A(n20569), .ZN(n20565) );
  OAI22_X1 U23542 ( .A1(n20566), .A2(n20648), .B1(n20565), .B2(n20708), .ZN(
        n20586) );
  AOI22_X1 U23543 ( .A1(n20651), .A2(n20586), .B1(n20650), .B2(n20585), .ZN(
        n20572) );
  NAND2_X1 U23544 ( .A1(n20567), .A2(n20566), .ZN(n20568) );
  OAI221_X1 U23545 ( .B1(n20570), .B2(n20569), .C1(n20648), .C2(n20568), .A(
        n20640), .ZN(n20588) );
  AOI22_X1 U23546 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20588), .B1(
        n20587), .B2(n20653), .ZN(n20571) );
  OAI211_X1 U23547 ( .C1(n20603), .C2(n20595), .A(n20572), .B(n20571), .ZN(
        P1_U3137) );
  AOI22_X1 U23548 ( .A1(n20658), .A2(n20586), .B1(n20657), .B2(n20585), .ZN(
        n20574) );
  AOI22_X1 U23549 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20588), .B1(
        n20587), .B2(n20604), .ZN(n20573) );
  OAI211_X1 U23550 ( .C1(n20607), .C2(n20595), .A(n20574), .B(n20573), .ZN(
        P1_U3138) );
  AOI22_X1 U23551 ( .A1(n20665), .A2(n20586), .B1(n20664), .B2(n20585), .ZN(
        n20576) );
  AOI22_X1 U23552 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20588), .B1(
        n20587), .B2(n20608), .ZN(n20575) );
  OAI211_X1 U23553 ( .C1(n20611), .C2(n20595), .A(n20576), .B(n20575), .ZN(
        P1_U3139) );
  AOI22_X1 U23554 ( .A1(n20671), .A2(n20586), .B1(n20670), .B2(n20585), .ZN(
        n20578) );
  AOI22_X1 U23555 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20588), .B1(
        n20587), .B2(n20612), .ZN(n20577) );
  OAI211_X1 U23556 ( .C1(n20615), .C2(n20595), .A(n20578), .B(n20577), .ZN(
        P1_U3140) );
  AOI22_X1 U23557 ( .A1(n20677), .A2(n20586), .B1(n20676), .B2(n20585), .ZN(
        n20580) );
  AOI22_X1 U23558 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20588), .B1(
        n20587), .B2(n20616), .ZN(n20579) );
  OAI211_X1 U23559 ( .C1(n20619), .C2(n20595), .A(n20580), .B(n20579), .ZN(
        P1_U3141) );
  AOI22_X1 U23560 ( .A1(n20683), .A2(n20586), .B1(n20682), .B2(n20585), .ZN(
        n20582) );
  AOI22_X1 U23561 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20588), .B1(
        n20587), .B2(n20620), .ZN(n20581) );
  OAI211_X1 U23562 ( .C1(n20623), .C2(n20595), .A(n20582), .B(n20581), .ZN(
        P1_U3142) );
  AOI22_X1 U23563 ( .A1(n20689), .A2(n20586), .B1(n20688), .B2(n20585), .ZN(
        n20584) );
  AOI22_X1 U23564 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20588), .B1(
        n20587), .B2(n20624), .ZN(n20583) );
  OAI211_X1 U23565 ( .C1(n20627), .C2(n20595), .A(n20584), .B(n20583), .ZN(
        P1_U3143) );
  AOI22_X1 U23566 ( .A1(n20697), .A2(n20586), .B1(n20695), .B2(n20585), .ZN(
        n20590) );
  AOI22_X1 U23567 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20588), .B1(
        n20587), .B2(n20630), .ZN(n20589) );
  OAI211_X1 U23568 ( .C1(n20635), .C2(n20595), .A(n20590), .B(n20589), .ZN(
        P1_U3144) );
  NAND2_X1 U23569 ( .A1(n20646), .A2(n20592), .ZN(n20596) );
  OAI22_X1 U23570 ( .A1(n20596), .A2(n20648), .B1(n20594), .B2(n20593), .ZN(
        n20629) );
  NOR3_X2 U23571 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20638), .A3(
        n20642), .ZN(n20628) );
  AOI22_X1 U23572 ( .A1(n20651), .A2(n20629), .B1(n20650), .B2(n20628), .ZN(
        n20602) );
  INV_X1 U23573 ( .A(n20703), .ZN(n20654) );
  OAI21_X1 U23574 ( .B1(n20654), .B2(n20631), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20597) );
  AOI21_X1 U23575 ( .B1(n20597), .B2(n20596), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20600) );
  AOI22_X1 U23576 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20632), .B1(
        n20631), .B2(n20653), .ZN(n20601) );
  OAI211_X1 U23577 ( .C1(n20603), .C2(n20703), .A(n20602), .B(n20601), .ZN(
        P1_U3145) );
  AOI22_X1 U23578 ( .A1(n20658), .A2(n20629), .B1(n20657), .B2(n20628), .ZN(
        n20606) );
  AOI22_X1 U23579 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20632), .B1(
        n20631), .B2(n20604), .ZN(n20605) );
  OAI211_X1 U23580 ( .C1(n20607), .C2(n20703), .A(n20606), .B(n20605), .ZN(
        P1_U3146) );
  AOI22_X1 U23581 ( .A1(n20665), .A2(n20629), .B1(n20664), .B2(n20628), .ZN(
        n20610) );
  AOI22_X1 U23582 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20632), .B1(
        n20631), .B2(n20608), .ZN(n20609) );
  OAI211_X1 U23583 ( .C1(n20611), .C2(n20703), .A(n20610), .B(n20609), .ZN(
        P1_U3147) );
  AOI22_X1 U23584 ( .A1(n20671), .A2(n20629), .B1(n20670), .B2(n20628), .ZN(
        n20614) );
  AOI22_X1 U23585 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20632), .B1(
        n20631), .B2(n20612), .ZN(n20613) );
  OAI211_X1 U23586 ( .C1(n20615), .C2(n20703), .A(n20614), .B(n20613), .ZN(
        P1_U3148) );
  AOI22_X1 U23587 ( .A1(n20677), .A2(n20629), .B1(n20676), .B2(n20628), .ZN(
        n20618) );
  AOI22_X1 U23588 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20632), .B1(
        n20631), .B2(n20616), .ZN(n20617) );
  OAI211_X1 U23589 ( .C1(n20619), .C2(n20703), .A(n20618), .B(n20617), .ZN(
        P1_U3149) );
  AOI22_X1 U23590 ( .A1(n20683), .A2(n20629), .B1(n20682), .B2(n20628), .ZN(
        n20622) );
  AOI22_X1 U23591 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20632), .B1(
        n20631), .B2(n20620), .ZN(n20621) );
  OAI211_X1 U23592 ( .C1(n20623), .C2(n20703), .A(n20622), .B(n20621), .ZN(
        P1_U3150) );
  AOI22_X1 U23593 ( .A1(n20689), .A2(n20629), .B1(n20688), .B2(n20628), .ZN(
        n20626) );
  AOI22_X1 U23594 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20632), .B1(
        n20631), .B2(n20624), .ZN(n20625) );
  OAI211_X1 U23595 ( .C1(n20627), .C2(n20703), .A(n20626), .B(n20625), .ZN(
        P1_U3151) );
  AOI22_X1 U23596 ( .A1(n20697), .A2(n20629), .B1(n20695), .B2(n20628), .ZN(
        n20634) );
  AOI22_X1 U23597 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20632), .B1(
        n20631), .B2(n20630), .ZN(n20633) );
  OAI211_X1 U23598 ( .C1(n20635), .C2(n20703), .A(n20634), .B(n20633), .ZN(
        P1_U3152) );
  NAND3_X1 U23599 ( .A1(n20637), .A2(n20570), .A3(n20636), .ZN(n20639) );
  OR2_X1 U23600 ( .A1(n20638), .A2(n20642), .ZN(n20647) );
  NAND2_X1 U23601 ( .A1(n20639), .A2(n20647), .ZN(n20641) );
  INV_X1 U23602 ( .A(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n21047) );
  INV_X1 U23603 ( .A(n20642), .ZN(n20643) );
  AND2_X1 U23604 ( .A1(n20644), .A2(n20643), .ZN(n20694) );
  AOI21_X1 U23605 ( .B1(n20646), .B2(n20645), .A(n20694), .ZN(n20649) );
  OAI22_X1 U23606 ( .A1(n20649), .A2(n20648), .B1(n20647), .B2(n20708), .ZN(
        n20696) );
  AOI22_X1 U23607 ( .A1(n20651), .A2(n20696), .B1(n20650), .B2(n20694), .ZN(
        n20656) );
  AOI22_X1 U23608 ( .A1(n20654), .A2(n20653), .B1(n20699), .B2(n20652), .ZN(
        n20655) );
  OAI211_X1 U23609 ( .C1(n20659), .C2(n21047), .A(n20656), .B(n20655), .ZN(
        P1_U3153) );
  AOI22_X1 U23610 ( .A1(n20658), .A2(n20696), .B1(n20657), .B2(n20694), .ZN(
        n20662) );
  INV_X1 U23611 ( .A(n20659), .ZN(n20700) );
  AOI22_X1 U23612 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20700), .B1(
        n20699), .B2(n20660), .ZN(n20661) );
  OAI211_X1 U23613 ( .C1(n20663), .C2(n20703), .A(n20662), .B(n20661), .ZN(
        P1_U3154) );
  AOI22_X1 U23614 ( .A1(n20665), .A2(n20696), .B1(n20664), .B2(n20694), .ZN(
        n20668) );
  AOI22_X1 U23615 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20700), .B1(
        n20699), .B2(n20666), .ZN(n20667) );
  OAI211_X1 U23616 ( .C1(n20669), .C2(n20703), .A(n20668), .B(n20667), .ZN(
        P1_U3155) );
  AOI22_X1 U23617 ( .A1(n20671), .A2(n20696), .B1(n20670), .B2(n20694), .ZN(
        n20674) );
  AOI22_X1 U23618 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20700), .B1(
        n20699), .B2(n20672), .ZN(n20673) );
  OAI211_X1 U23619 ( .C1(n20675), .C2(n20703), .A(n20674), .B(n20673), .ZN(
        P1_U3156) );
  AOI22_X1 U23620 ( .A1(n20677), .A2(n20696), .B1(n20676), .B2(n20694), .ZN(
        n20680) );
  AOI22_X1 U23621 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20700), .B1(
        n20699), .B2(n20678), .ZN(n20679) );
  OAI211_X1 U23622 ( .C1(n20681), .C2(n20703), .A(n20680), .B(n20679), .ZN(
        P1_U3157) );
  AOI22_X1 U23623 ( .A1(n20683), .A2(n20696), .B1(n20682), .B2(n20694), .ZN(
        n20686) );
  AOI22_X1 U23624 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20700), .B1(
        n20699), .B2(n20684), .ZN(n20685) );
  OAI211_X1 U23625 ( .C1(n20687), .C2(n20703), .A(n20686), .B(n20685), .ZN(
        P1_U3158) );
  AOI22_X1 U23626 ( .A1(n20689), .A2(n20696), .B1(n20688), .B2(n20694), .ZN(
        n20692) );
  AOI22_X1 U23627 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20700), .B1(
        n20699), .B2(n20690), .ZN(n20691) );
  OAI211_X1 U23628 ( .C1(n20693), .C2(n20703), .A(n20692), .B(n20691), .ZN(
        P1_U3159) );
  AOI22_X1 U23629 ( .A1(n20697), .A2(n20696), .B1(n20695), .B2(n20694), .ZN(
        n20702) );
  AOI22_X1 U23630 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20700), .B1(
        n20699), .B2(n20698), .ZN(n20701) );
  OAI211_X1 U23631 ( .C1(n20704), .C2(n20703), .A(n20702), .B(n20701), .ZN(
        P1_U3160) );
  NOR2_X1 U23632 ( .A1(n20706), .A2(n20705), .ZN(n20709) );
  OAI21_X1 U23633 ( .B1(n20709), .B2(n20708), .A(n20707), .ZN(P1_U3163) );
  INV_X1 U23634 ( .A(P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20940) );
  NOR2_X1 U23635 ( .A1(n20787), .A2(n20940), .ZN(P1_U3164) );
  AND2_X1 U23636 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20783), .ZN(
        P1_U3165) );
  AND2_X1 U23637 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20783), .ZN(
        P1_U3166) );
  INV_X1 U23638 ( .A(P1_DATAWIDTH_REG_28__SCAN_IN), .ZN(n20988) );
  NOR2_X1 U23639 ( .A1(n20787), .A2(n20988), .ZN(P1_U3167) );
  AND2_X1 U23640 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20783), .ZN(
        P1_U3168) );
  AND2_X1 U23641 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20783), .ZN(
        P1_U3169) );
  AND2_X1 U23642 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20783), .ZN(
        P1_U3170) );
  AND2_X1 U23643 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20783), .ZN(
        P1_U3171) );
  AND2_X1 U23644 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20783), .ZN(
        P1_U3172) );
  AND2_X1 U23645 ( .A1(n20783), .A2(P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(
        P1_U3173) );
  AND2_X1 U23646 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20783), .ZN(
        P1_U3174) );
  AND2_X1 U23647 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20783), .ZN(
        P1_U3175) );
  AND2_X1 U23648 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20783), .ZN(
        P1_U3176) );
  AND2_X1 U23649 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20783), .ZN(
        P1_U3177) );
  AND2_X1 U23650 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20783), .ZN(
        P1_U3178) );
  AND2_X1 U23651 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20783), .ZN(
        P1_U3179) );
  AND2_X1 U23652 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20783), .ZN(
        P1_U3180) );
  AND2_X1 U23653 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20783), .ZN(
        P1_U3181) );
  AND2_X1 U23654 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20783), .ZN(
        P1_U3182) );
  AND2_X1 U23655 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20783), .ZN(
        P1_U3183) );
  AND2_X1 U23656 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20783), .ZN(
        P1_U3184) );
  AND2_X1 U23657 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20783), .ZN(
        P1_U3185) );
  AND2_X1 U23658 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20783), .ZN(P1_U3186) );
  AND2_X1 U23659 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20783), .ZN(P1_U3187) );
  AND2_X1 U23660 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20783), .ZN(P1_U3188) );
  AND2_X1 U23661 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20783), .ZN(P1_U3189) );
  AND2_X1 U23662 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20783), .ZN(P1_U3190) );
  AND2_X1 U23663 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20783), .ZN(P1_U3191) );
  AND2_X1 U23664 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20783), .ZN(P1_U3192) );
  AND2_X1 U23665 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20783), .ZN(P1_U3193) );
  NAND2_X1 U23666 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20717), .ZN(n20716) );
  INV_X1 U23667 ( .A(n20716), .ZN(n20713) );
  INV_X2 U23668 ( .A(n20810), .ZN(n20823) );
  OAI21_X1 U23669 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20718), .A(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20710) );
  AOI211_X1 U23670 ( .C1(HOLD), .C2(P1_STATE_REG_1__SCAN_IN), .A(n20711), .B(
        n20710), .ZN(n20712) );
  OAI22_X1 U23671 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20713), .B1(n20823), 
        .B2(n20712), .ZN(P1_U3194) );
  INV_X1 U23672 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20715) );
  OAI211_X1 U23673 ( .C1(NA), .C2(n20818), .A(P1_STATE_REG_1__SCAN_IN), .B(
        n20724), .ZN(n20714) );
  OAI211_X1 U23674 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20715), .A(
        P1_STATE_REG_0__SCAN_IN), .B(n20714), .ZN(n20722) );
  OAI211_X1 U23675 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n20718), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n20716), .ZN(n20721) );
  INV_X1 U23676 ( .A(n20717), .ZN(n20719) );
  NAND4_X1 U23677 ( .A1(P1_REQUESTPENDING_REG_SCAN_IN), .A2(
        P1_STATE_REG_0__SCAN_IN), .A3(n20719), .A4(n20718), .ZN(n20720) );
  OAI211_X1 U23678 ( .C1(n20723), .C2(n20722), .A(n20721), .B(n20720), .ZN(
        P1_U3196) );
  NAND2_X1 U23679 ( .A1(n20823), .A2(n20724), .ZN(n20771) );
  INV_X1 U23680 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20725) );
  AND2_X1 U23681 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20823), .ZN(n20769) );
  OAI222_X1 U23682 ( .A1(n20771), .A2(n20727), .B1(n20725), .B2(n20823), .C1(
        n13981), .C2(n20775), .ZN(P1_U3197) );
  INV_X1 U23683 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n20726) );
  OAI222_X1 U23684 ( .A1(n20775), .A2(n20727), .B1(n20726), .B2(n20823), .C1(
        n13791), .C2(n20771), .ZN(P1_U3198) );
  INV_X1 U23685 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20730) );
  OAI222_X1 U23686 ( .A1(n20775), .A2(n13791), .B1(n20728), .B2(n20823), .C1(
        n20730), .C2(n20771), .ZN(P1_U3199) );
  INV_X1 U23687 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20729) );
  OAI222_X1 U23688 ( .A1(n20775), .A2(n20730), .B1(n20729), .B2(n20823), .C1(
        n20732), .C2(n20771), .ZN(P1_U3200) );
  INV_X1 U23689 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n20731) );
  OAI222_X1 U23690 ( .A1(n20775), .A2(n20732), .B1(n20731), .B2(n20823), .C1(
        n20733), .C2(n20771), .ZN(P1_U3201) );
  INV_X1 U23691 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n21108) );
  OAI222_X1 U23692 ( .A1(n20775), .A2(n20733), .B1(n21108), .B2(n20823), .C1(
        n20735), .C2(n20771), .ZN(P1_U3202) );
  INV_X1 U23693 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n20734) );
  OAI222_X1 U23694 ( .A1(n20775), .A2(n20735), .B1(n20734), .B2(n20823), .C1(
        n20737), .C2(n20771), .ZN(P1_U3203) );
  INV_X1 U23695 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20736) );
  OAI222_X1 U23696 ( .A1(n20775), .A2(n20737), .B1(n20736), .B2(n20823), .C1(
        n20739), .C2(n20771), .ZN(P1_U3204) );
  INV_X1 U23697 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n20738) );
  OAI222_X1 U23698 ( .A1(n20775), .A2(n20739), .B1(n20738), .B2(n20823), .C1(
        n20740), .C2(n20771), .ZN(P1_U3205) );
  INV_X1 U23699 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n20741) );
  OAI222_X1 U23700 ( .A1(n20771), .A2(n20743), .B1(n20741), .B2(n20823), .C1(
        n20740), .C2(n20775), .ZN(P1_U3206) );
  INV_X1 U23701 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n20742) );
  OAI222_X1 U23702 ( .A1(n20775), .A2(n20743), .B1(n20742), .B2(n20823), .C1(
        n20744), .C2(n20771), .ZN(P1_U3207) );
  INV_X1 U23703 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n20745) );
  OAI222_X1 U23704 ( .A1(n20771), .A2(n20746), .B1(n20745), .B2(n20823), .C1(
        n20744), .C2(n20775), .ZN(P1_U3208) );
  INV_X1 U23705 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n21111) );
  OAI222_X1 U23706 ( .A1(n20775), .A2(n20746), .B1(n21111), .B2(n20823), .C1(
        n14927), .C2(n20771), .ZN(P1_U3209) );
  INV_X1 U23707 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n20747) );
  OAI222_X1 U23708 ( .A1(n20771), .A2(n20749), .B1(n20747), .B2(n20823), .C1(
        n14927), .C2(n20775), .ZN(P1_U3210) );
  INV_X1 U23709 ( .A(n20771), .ZN(n20768) );
  AOI22_X1 U23710 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(n20810), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n20768), .ZN(n20748) );
  OAI21_X1 U23711 ( .B1(n20749), .B2(n20775), .A(n20748), .ZN(P1_U3211) );
  AOI22_X1 U23712 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20810), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n20769), .ZN(n20750) );
  OAI21_X1 U23713 ( .B1(n20752), .B2(n20771), .A(n20750), .ZN(P1_U3212) );
  AOI22_X1 U23714 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20810), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n20768), .ZN(n20751) );
  OAI21_X1 U23715 ( .B1(n20752), .B2(n20775), .A(n20751), .ZN(P1_U3213) );
  INV_X1 U23716 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20754) );
  AOI22_X1 U23717 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n20810), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n20768), .ZN(n20753) );
  OAI21_X1 U23718 ( .B1(n20754), .B2(n20775), .A(n20753), .ZN(P1_U3214) );
  AOI22_X1 U23719 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n20810), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n20769), .ZN(n20755) );
  OAI21_X1 U23720 ( .B1(n20756), .B2(n20771), .A(n20755), .ZN(P1_U3215) );
  INV_X1 U23721 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n20757) );
  OAI222_X1 U23722 ( .A1(n20771), .A2(n20759), .B1(n20757), .B2(n20823), .C1(
        n20756), .C2(n20775), .ZN(P1_U3216) );
  INV_X1 U23723 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20758) );
  OAI222_X1 U23724 ( .A1(n20775), .A2(n20759), .B1(n20758), .B2(n20823), .C1(
        n21030), .C2(n20771), .ZN(P1_U3217) );
  AOI22_X1 U23725 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n20810), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20768), .ZN(n20760) );
  OAI21_X1 U23726 ( .B1(n21030), .B2(n20775), .A(n20760), .ZN(P1_U3218) );
  INV_X1 U23727 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n21117) );
  OAI222_X1 U23728 ( .A1(n20775), .A2(n15052), .B1(n21117), .B2(n20823), .C1(
        n20762), .C2(n20771), .ZN(P1_U3219) );
  INV_X1 U23729 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n20761) );
  OAI222_X1 U23730 ( .A1(n20775), .A2(n20762), .B1(n20761), .B2(n20823), .C1(
        n14876), .C2(n20771), .ZN(P1_U3220) );
  INV_X1 U23731 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20764) );
  OAI222_X1 U23732 ( .A1(n20775), .A2(n14876), .B1(n20764), .B2(n20823), .C1(
        n20763), .C2(n20771), .ZN(P1_U3221) );
  AOI222_X1 U23733 ( .A1(n20769), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20810), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20768), .ZN(n20765) );
  INV_X1 U23734 ( .A(n20765), .ZN(P1_U3222) );
  AOI222_X1 U23735 ( .A1(n20769), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20810), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20768), .ZN(n20766) );
  INV_X1 U23736 ( .A(n20766), .ZN(P1_U3223) );
  AOI222_X1 U23737 ( .A1(n20769), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20810), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20768), .ZN(n20767) );
  INV_X1 U23738 ( .A(n20767), .ZN(P1_U3224) );
  AOI222_X1 U23739 ( .A1(n20769), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20810), .C1(P1_REIP_REG_30__SCAN_IN), 
        .C2(n20768), .ZN(n20770) );
  INV_X1 U23740 ( .A(n20770), .ZN(P1_U3225) );
  INV_X1 U23741 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20773) );
  OAI222_X1 U23742 ( .A1(n20775), .A2(n20774), .B1(n20773), .B2(n20823), .C1(
        n20772), .C2(n20771), .ZN(P1_U3226) );
  INV_X1 U23743 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20776) );
  AOI22_X1 U23744 ( .A1(n20823), .A2(n20777), .B1(n20776), .B2(n20810), .ZN(
        P1_U3458) );
  INV_X1 U23745 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20804) );
  INV_X1 U23746 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20778) );
  AOI22_X1 U23747 ( .A1(n20823), .A2(n20804), .B1(n20778), .B2(n20810), .ZN(
        P1_U3459) );
  INV_X1 U23748 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20779) );
  AOI22_X1 U23749 ( .A1(n20823), .A2(n20780), .B1(n20779), .B2(n20810), .ZN(
        P1_U3460) );
  INV_X1 U23750 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20809) );
  INV_X1 U23751 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20781) );
  AOI22_X1 U23752 ( .A1(n20823), .A2(n20809), .B1(n20781), .B2(n20810), .ZN(
        P1_U3461) );
  INV_X1 U23753 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20784) );
  INV_X1 U23754 ( .A(n20785), .ZN(n20782) );
  AOI21_X1 U23755 ( .B1(n20784), .B2(n20783), .A(n20782), .ZN(P1_U3464) );
  OAI21_X1 U23756 ( .B1(n20787), .B2(n20786), .A(n20785), .ZN(P1_U3465) );
  INV_X1 U23757 ( .A(n20788), .ZN(n20789) );
  OAI22_X1 U23758 ( .A1(n20791), .A2(n20790), .B1(n20794), .B2(n20789), .ZN(
        n20792) );
  MUX2_X1 U23759 ( .A(n20792), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n20799), .Z(P1_U3469) );
  OAI22_X1 U23760 ( .A1(n20796), .A2(n20795), .B1(n20794), .B2(n20793), .ZN(
        n20798) );
  AOI22_X1 U23761 ( .A1(n20799), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n20798), .B2(n20797), .ZN(n20800) );
  OAI21_X1 U23762 ( .B1(n20802), .B2(n20801), .A(n20800), .ZN(P1_U3472) );
  AOI21_X1 U23763 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20803) );
  AOI22_X1 U23764 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20803), .B2(n13981), .ZN(n20805) );
  AOI22_X1 U23765 ( .A1(n20806), .A2(n20805), .B1(n20804), .B2(n20808), .ZN(
        P1_U3481) );
  NOR2_X1 U23766 ( .A1(n20808), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20807) );
  AOI22_X1 U23767 ( .A1(n20809), .A2(n20808), .B1(n13493), .B2(n20807), .ZN(
        P1_U3482) );
  AOI22_X1 U23768 ( .A1(n20823), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20811), 
        .B2(n20810), .ZN(P1_U3483) );
  OAI21_X1 U23769 ( .B1(n20812), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20814) );
  OAI21_X1 U23770 ( .B1(n20815), .B2(n20814), .A(n20813), .ZN(n20822) );
  AOI211_X1 U23771 ( .C1(n20819), .C2(n20818), .A(n20817), .B(n20816), .ZN(
        n20821) );
  NAND2_X1 U23772 ( .A1(n20821), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20820) );
  OAI21_X1 U23773 ( .B1(n20822), .B2(n20821), .A(n20820), .ZN(P1_U3485) );
  MUX2_X1 U23774 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(P1_MEMORYFETCH_REG_SCAN_IN), 
        .S(n20823), .Z(P1_U3486) );
  AOI22_X1 U23775 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(keyinput245), .B1(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(keyinput201), .ZN(n20824) );
  OAI221_X1 U23776 ( .B1(P3_DATAWIDTH_REG_18__SCAN_IN), .B2(keyinput245), .C1(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(keyinput201), .A(n20824), 
        .ZN(n20831) );
  AOI22_X1 U23777 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(keyinput129), .B1(
        P1_INSTQUEUE_REG_4__6__SCAN_IN), .B2(keyinput179), .ZN(n20825) );
  OAI221_X1 U23778 ( .B1(P1_DATAO_REG_3__SCAN_IN), .B2(keyinput129), .C1(
        P1_INSTQUEUE_REG_4__6__SCAN_IN), .C2(keyinput179), .A(n20825), .ZN(
        n20830) );
  AOI22_X1 U23779 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(keyinput166), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(keyinput136), .ZN(n20826) );
  OAI221_X1 U23780 ( .B1(P3_EAX_REG_23__SCAN_IN), .B2(keyinput166), .C1(
        P2_REIP_REG_30__SCAN_IN), .C2(keyinput136), .A(n20826), .ZN(n20829) );
  AOI22_X1 U23781 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(keyinput207), 
        .B1(P2_ADDRESS_REG_3__SCAN_IN), .B2(keyinput148), .ZN(n20827) );
  OAI221_X1 U23782 ( .B1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B2(keyinput207), 
        .C1(P2_ADDRESS_REG_3__SCAN_IN), .C2(keyinput148), .A(n20827), .ZN(
        n20828) );
  NOR4_X1 U23783 ( .A1(n20831), .A2(n20830), .A3(n20829), .A4(n20828), .ZN(
        n20859) );
  AOI22_X1 U23784 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(keyinput255), .B1(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(keyinput228), .ZN(n20832) );
  OAI221_X1 U23785 ( .B1(P1_UWORD_REG_6__SCAN_IN), .B2(keyinput255), .C1(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(keyinput228), .A(n20832), .ZN(
        n20839) );
  AOI22_X1 U23786 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(keyinput145), .B1(
        P2_EBX_REG_9__SCAN_IN), .B2(keyinput190), .ZN(n20833) );
  OAI221_X1 U23787 ( .B1(P3_REIP_REG_8__SCAN_IN), .B2(keyinput145), .C1(
        P2_EBX_REG_9__SCAN_IN), .C2(keyinput190), .A(n20833), .ZN(n20838) );
  AOI22_X1 U23788 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(keyinput161), 
        .B1(P2_REIP_REG_29__SCAN_IN), .B2(keyinput226), .ZN(n20834) );
  OAI221_X1 U23789 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(keyinput161), 
        .C1(P2_REIP_REG_29__SCAN_IN), .C2(keyinput226), .A(n20834), .ZN(n20837) );
  AOI22_X1 U23790 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(keyinput167), .B1(
        P2_EBX_REG_29__SCAN_IN), .B2(keyinput206), .ZN(n20835) );
  OAI221_X1 U23791 ( .B1(P1_DATAWIDTH_REG_22__SCAN_IN), .B2(keyinput167), .C1(
        P2_EBX_REG_29__SCAN_IN), .C2(keyinput206), .A(n20835), .ZN(n20836) );
  NOR4_X1 U23792 ( .A1(n20839), .A2(n20838), .A3(n20837), .A4(n20836), .ZN(
        n20858) );
  AOI22_X1 U23793 ( .A1(P3_DATAO_REG_8__SCAN_IN), .A2(keyinput205), .B1(
        P3_DATAO_REG_16__SCAN_IN), .B2(keyinput253), .ZN(n20840) );
  OAI221_X1 U23794 ( .B1(P3_DATAO_REG_8__SCAN_IN), .B2(keyinput205), .C1(
        P3_DATAO_REG_16__SCAN_IN), .C2(keyinput253), .A(n20840), .ZN(n20847)
         );
  AOI22_X1 U23795 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(keyinput153), 
        .B1(P1_REIP_REG_22__SCAN_IN), .B2(keyinput195), .ZN(n20841) );
  OAI221_X1 U23796 ( .B1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B2(keyinput153), 
        .C1(P1_REIP_REG_22__SCAN_IN), .C2(keyinput195), .A(n20841), .ZN(n20846) );
  AOI22_X1 U23797 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(keyinput242), .B1(
        P2_INSTQUEUE_REG_7__4__SCAN_IN), .B2(keyinput224), .ZN(n20842) );
  OAI221_X1 U23798 ( .B1(P2_DATAO_REG_3__SCAN_IN), .B2(keyinput242), .C1(
        P2_INSTQUEUE_REG_7__4__SCAN_IN), .C2(keyinput224), .A(n20842), .ZN(
        n20845) );
  AOI22_X1 U23799 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(keyinput189), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(keyinput135), .ZN(n20843) );
  OAI221_X1 U23800 ( .B1(P1_LWORD_REG_5__SCAN_IN), .B2(keyinput189), .C1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .C2(keyinput135), .A(n20843), .ZN(
        n20844) );
  NOR4_X1 U23801 ( .A1(n20847), .A2(n20846), .A3(n20845), .A4(n20844), .ZN(
        n20857) );
  AOI22_X1 U23802 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(keyinput234), .B1(
        DATAI_9_), .B2(keyinput157), .ZN(n20848) );
  OAI221_X1 U23803 ( .B1(P3_REIP_REG_2__SCAN_IN), .B2(keyinput234), .C1(
        DATAI_9_), .C2(keyinput157), .A(n20848), .ZN(n20855) );
  AOI22_X1 U23804 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(keyinput141), .B1(
        P1_INSTQUEUE_REG_7__7__SCAN_IN), .B2(keyinput187), .ZN(n20849) );
  OAI221_X1 U23805 ( .B1(P3_DATAWIDTH_REG_19__SCAN_IN), .B2(keyinput141), .C1(
        P1_INSTQUEUE_REG_7__7__SCAN_IN), .C2(keyinput187), .A(n20849), .ZN(
        n20854) );
  AOI22_X1 U23806 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(keyinput169), .B1(
        P2_INSTQUEUE_REG_7__0__SCAN_IN), .B2(keyinput165), .ZN(n20850) );
  OAI221_X1 U23807 ( .B1(P3_DATAWIDTH_REG_26__SCAN_IN), .B2(keyinput169), .C1(
        P2_INSTQUEUE_REG_7__0__SCAN_IN), .C2(keyinput165), .A(n20850), .ZN(
        n20853) );
  AOI22_X1 U23808 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(keyinput159), 
        .B1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(keyinput139), .ZN(n20851) );
  OAI221_X1 U23809 ( .B1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B2(keyinput159), 
        .C1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .C2(keyinput139), .A(n20851), 
        .ZN(n20852) );
  NOR4_X1 U23810 ( .A1(n20855), .A2(n20854), .A3(n20853), .A4(n20852), .ZN(
        n20856) );
  NAND4_X1 U23811 ( .A1(n20859), .A2(n20858), .A3(n20857), .A4(n20856), .ZN(
        n21004) );
  AOI22_X1 U23812 ( .A1(P1_EAX_REG_20__SCAN_IN), .A2(keyinput223), .B1(
        P1_INSTQUEUE_REG_1__1__SCAN_IN), .B2(keyinput211), .ZN(n20860) );
  OAI221_X1 U23813 ( .B1(P1_EAX_REG_20__SCAN_IN), .B2(keyinput223), .C1(
        P1_INSTQUEUE_REG_1__1__SCAN_IN), .C2(keyinput211), .A(n20860), .ZN(
        n20867) );
  AOI22_X1 U23814 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(keyinput191), .B1(
        P1_EBX_REG_22__SCAN_IN), .B2(keyinput173), .ZN(n20861) );
  OAI221_X1 U23815 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(keyinput191), .C1(
        P1_EBX_REG_22__SCAN_IN), .C2(keyinput173), .A(n20861), .ZN(n20866) );
  AOI22_X1 U23816 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(keyinput186), 
        .B1(P2_EAX_REG_26__SCAN_IN), .B2(keyinput210), .ZN(n20862) );
  OAI221_X1 U23817 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(keyinput186), 
        .C1(P2_EAX_REG_26__SCAN_IN), .C2(keyinput210), .A(n20862), .ZN(n20865)
         );
  AOI22_X1 U23818 ( .A1(DATAI_26_), .A2(keyinput156), .B1(
        P2_INSTQUEUE_REG_0__3__SCAN_IN), .B2(keyinput181), .ZN(n20863) );
  OAI221_X1 U23819 ( .B1(DATAI_26_), .B2(keyinput156), .C1(
        P2_INSTQUEUE_REG_0__3__SCAN_IN), .C2(keyinput181), .A(n20863), .ZN(
        n20864) );
  NOR4_X1 U23820 ( .A1(n20867), .A2(n20866), .A3(n20865), .A4(n20864), .ZN(
        n20898) );
  AOI22_X1 U23821 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(keyinput185), .B1(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(keyinput128), .ZN(n20868) );
  OAI221_X1 U23822 ( .B1(P3_REIP_REG_13__SCAN_IN), .B2(keyinput185), .C1(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(keyinput128), .A(n20868), .ZN(
        n20875) );
  AOI22_X1 U23823 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(keyinput208), 
        .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(keyinput177), .ZN(n20869)
         );
  OAI221_X1 U23824 ( .B1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(keyinput208), 
        .C1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(keyinput177), .A(n20869), 
        .ZN(n20874) );
  AOI22_X1 U23825 ( .A1(P2_LWORD_REG_7__SCAN_IN), .A2(keyinput180), .B1(
        P2_INSTQUEUE_REG_14__2__SCAN_IN), .B2(keyinput196), .ZN(n20870) );
  OAI221_X1 U23826 ( .B1(P2_LWORD_REG_7__SCAN_IN), .B2(keyinput180), .C1(
        P2_INSTQUEUE_REG_14__2__SCAN_IN), .C2(keyinput196), .A(n20870), .ZN(
        n20873) );
  AOI22_X1 U23827 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(keyinput174), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(keyinput176), .ZN(n20871) );
  OAI221_X1 U23828 ( .B1(P1_UWORD_REG_12__SCAN_IN), .B2(keyinput174), .C1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(keyinput176), .A(n20871), .ZN(
        n20872) );
  NOR4_X1 U23829 ( .A1(n20875), .A2(n20874), .A3(n20873), .A4(n20872), .ZN(
        n20897) );
  AOI22_X1 U23830 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(keyinput137), .B1(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(keyinput138), .ZN(n20876) );
  OAI221_X1 U23831 ( .B1(P1_ADDRESS_REG_22__SCAN_IN), .B2(keyinput137), .C1(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(keyinput138), .A(n20876), .ZN(
        n20883) );
  AOI22_X1 U23832 ( .A1(P1_EAX_REG_25__SCAN_IN), .A2(keyinput251), .B1(
        P2_INSTQUEUE_REG_11__2__SCAN_IN), .B2(keyinput225), .ZN(n20877) );
  OAI221_X1 U23833 ( .B1(P1_EAX_REG_25__SCAN_IN), .B2(keyinput251), .C1(
        P2_INSTQUEUE_REG_11__2__SCAN_IN), .C2(keyinput225), .A(n20877), .ZN(
        n20882) );
  AOI22_X1 U23834 ( .A1(BUF1_REG_1__SCAN_IN), .A2(keyinput164), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(keyinput183), .ZN(n20878) );
  OAI221_X1 U23835 ( .B1(BUF1_REG_1__SCAN_IN), .B2(keyinput164), .C1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .C2(keyinput183), .A(n20878), .ZN(
        n20881) );
  AOI22_X1 U23836 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(keyinput220), .B1(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(keyinput144), .ZN(n20879) );
  OAI221_X1 U23837 ( .B1(P2_DATAWIDTH_REG_21__SCAN_IN), .B2(keyinput220), .C1(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(keyinput144), .A(n20879), 
        .ZN(n20880) );
  NOR4_X1 U23838 ( .A1(n20883), .A2(n20882), .A3(n20881), .A4(n20880), .ZN(
        n20896) );
  AOI22_X1 U23839 ( .A1(P1_DATAO_REG_31__SCAN_IN), .A2(keyinput175), .B1(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .B2(keyinput250), .ZN(n20884) );
  OAI221_X1 U23840 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(keyinput175), .C1(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .C2(keyinput250), .A(n20884), .ZN(
        n20894) );
  AOI22_X1 U23841 ( .A1(P3_DATAO_REG_23__SCAN_IN), .A2(keyinput130), .B1(
        BUF2_REG_28__SCAN_IN), .B2(keyinput142), .ZN(n20885) );
  OAI221_X1 U23842 ( .B1(P3_DATAO_REG_23__SCAN_IN), .B2(keyinput130), .C1(
        BUF2_REG_28__SCAN_IN), .C2(keyinput142), .A(n20885), .ZN(n20893) );
  INV_X1 U23843 ( .A(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n21125) );
  AOI22_X1 U23844 ( .A1(n21125), .A2(keyinput249), .B1(keyinput170), .B2(
        n20887), .ZN(n20886) );
  OAI221_X1 U23845 ( .B1(n21125), .B2(keyinput249), .C1(n20887), .C2(
        keyinput170), .A(n20886), .ZN(n20892) );
  AOI22_X1 U23846 ( .A1(n20890), .A2(keyinput162), .B1(n20889), .B2(
        keyinput184), .ZN(n20888) );
  OAI221_X1 U23847 ( .B1(n20890), .B2(keyinput162), .C1(n20889), .C2(
        keyinput184), .A(n20888), .ZN(n20891) );
  NOR4_X1 U23848 ( .A1(n20894), .A2(n20893), .A3(n20892), .A4(n20891), .ZN(
        n20895) );
  NAND4_X1 U23849 ( .A1(n20898), .A2(n20897), .A3(n20896), .A4(n20895), .ZN(
        n21003) );
  INV_X1 U23850 ( .A(P3_UWORD_REG_5__SCAN_IN), .ZN(n21092) );
  AOI22_X1 U23851 ( .A1(n21092), .A2(keyinput227), .B1(n20900), .B2(
        keyinput239), .ZN(n20899) );
  OAI221_X1 U23852 ( .B1(n21092), .B2(keyinput227), .C1(n20900), .C2(
        keyinput239), .A(n20899), .ZN(n20909) );
  INV_X1 U23853 ( .A(P2_UWORD_REG_12__SCAN_IN), .ZN(n21060) );
  AOI22_X1 U23854 ( .A1(n21038), .A2(keyinput171), .B1(n21060), .B2(
        keyinput197), .ZN(n20901) );
  OAI221_X1 U23855 ( .B1(n21038), .B2(keyinput171), .C1(n21060), .C2(
        keyinput197), .A(n20901), .ZN(n20908) );
  INV_X1 U23856 ( .A(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n21021) );
  AOI22_X1 U23857 ( .A1(n20903), .A2(keyinput151), .B1(n21021), .B2(
        keyinput194), .ZN(n20902) );
  OAI221_X1 U23858 ( .B1(n20903), .B2(keyinput151), .C1(n21021), .C2(
        keyinput194), .A(n20902), .ZN(n20907) );
  XOR2_X1 U23859 ( .A(n11312), .B(keyinput149), .Z(n20905) );
  XNOR2_X1 U23860 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B(keyinput254), .ZN(
        n20904) );
  NAND2_X1 U23861 ( .A1(n20905), .A2(n20904), .ZN(n20906) );
  NOR4_X1 U23862 ( .A1(n20909), .A2(n20908), .A3(n20907), .A4(n20906), .ZN(
        n20949) );
  INV_X1 U23863 ( .A(P3_DATAO_REG_0__SCAN_IN), .ZN(n21014) );
  INV_X1 U23864 ( .A(DATAI_29_), .ZN(n20911) );
  AOI22_X1 U23865 ( .A1(n21014), .A2(keyinput192), .B1(n20911), .B2(
        keyinput236), .ZN(n20910) );
  OAI221_X1 U23866 ( .B1(n21014), .B2(keyinput192), .C1(n20911), .C2(
        keyinput236), .A(n20910), .ZN(n20921) );
  INV_X1 U23867 ( .A(P3_UWORD_REG_0__SCAN_IN), .ZN(n21102) );
  AOI22_X1 U23868 ( .A1(n21102), .A2(keyinput204), .B1(n20913), .B2(
        keyinput182), .ZN(n20912) );
  OAI221_X1 U23869 ( .B1(n21102), .B2(keyinput204), .C1(n20913), .C2(
        keyinput182), .A(n20912), .ZN(n20920) );
  AOI22_X1 U23870 ( .A1(n21007), .A2(keyinput200), .B1(n20915), .B2(
        keyinput238), .ZN(n20914) );
  OAI221_X1 U23871 ( .B1(n21007), .B2(keyinput200), .C1(n20915), .C2(
        keyinput238), .A(n20914), .ZN(n20919) );
  INV_X1 U23872 ( .A(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n21096) );
  AOI22_X1 U23873 ( .A1(n20917), .A2(keyinput213), .B1(keyinput158), .B2(
        n21096), .ZN(n20916) );
  OAI221_X1 U23874 ( .B1(n20917), .B2(keyinput213), .C1(n21096), .C2(
        keyinput158), .A(n20916), .ZN(n20918) );
  NOR4_X1 U23875 ( .A1(n20921), .A2(n20920), .A3(n20919), .A4(n20918), .ZN(
        n20948) );
  INV_X1 U23876 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n21055) );
  AOI22_X1 U23877 ( .A1(n20926), .A2(keyinput143), .B1(keyinput237), .B2(
        n21055), .ZN(n20925) );
  OAI221_X1 U23878 ( .B1(n20926), .B2(keyinput143), .C1(n21055), .C2(
        keyinput237), .A(n20925), .ZN(n20931) );
  INV_X1 U23879 ( .A(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n21056) );
  AOI22_X1 U23880 ( .A1(n21053), .A2(keyinput241), .B1(n21056), .B2(
        keyinput230), .ZN(n20927) );
  OAI221_X1 U23881 ( .B1(n21053), .B2(keyinput241), .C1(n21056), .C2(
        keyinput230), .A(n20927), .ZN(n20930) );
  INV_X1 U23882 ( .A(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n21109) );
  AOI22_X1 U23883 ( .A1(n21109), .A2(keyinput160), .B1(keyinput163), .B2(
        n21031), .ZN(n20928) );
  OAI221_X1 U23884 ( .B1(n21109), .B2(keyinput160), .C1(n21031), .C2(
        keyinput163), .A(n20928), .ZN(n20929) );
  NOR4_X1 U23885 ( .A1(n20932), .A2(n20931), .A3(n20930), .A4(n20929), .ZN(
        n20947) );
  INV_X1 U23886 ( .A(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n20934) );
  AOI22_X1 U23887 ( .A1(n20935), .A2(keyinput247), .B1(keyinput221), .B2(
        n20934), .ZN(n20933) );
  OAI221_X1 U23888 ( .B1(n20935), .B2(keyinput247), .C1(n20934), .C2(
        keyinput221), .A(n20933), .ZN(n20945) );
  AOI22_X1 U23889 ( .A1(n20937), .A2(keyinput132), .B1(n21185), .B2(
        keyinput193), .ZN(n20936) );
  OAI221_X1 U23890 ( .B1(n20937), .B2(keyinput132), .C1(n21185), .C2(
        keyinput193), .A(n20936), .ZN(n20944) );
  INV_X1 U23891 ( .A(P1_LWORD_REG_1__SCAN_IN), .ZN(n20939) );
  AOI22_X1 U23892 ( .A1(n20940), .A2(keyinput133), .B1(n20939), .B2(
        keyinput222), .ZN(n20938) );
  OAI221_X1 U23893 ( .B1(n20940), .B2(keyinput133), .C1(n20939), .C2(
        keyinput222), .A(n20938), .ZN(n20943) );
  AOI22_X1 U23894 ( .A1(n11469), .A2(keyinput240), .B1(keyinput172), .B2(
        n21073), .ZN(n20941) );
  OAI221_X1 U23895 ( .B1(n11469), .B2(keyinput240), .C1(n21073), .C2(
        keyinput172), .A(n20941), .ZN(n20942) );
  NOR4_X1 U23896 ( .A1(n20945), .A2(n20944), .A3(n20943), .A4(n20942), .ZN(
        n20946) );
  NAND4_X1 U23897 ( .A1(n20949), .A2(n20948), .A3(n20947), .A4(n20946), .ZN(
        n21002) );
  INV_X1 U23898 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n21015) );
  AOI22_X1 U23899 ( .A1(n21015), .A2(keyinput252), .B1(keyinput198), .B2(
        n21006), .ZN(n20950) );
  OAI221_X1 U23900 ( .B1(n21015), .B2(keyinput252), .C1(n21006), .C2(
        keyinput198), .A(n20950), .ZN(n20961) );
  AOI22_X1 U23901 ( .A1(n20953), .A2(keyinput202), .B1(keyinput155), .B2(
        n20952), .ZN(n20951) );
  OAI221_X1 U23902 ( .B1(n20953), .B2(keyinput202), .C1(n20952), .C2(
        keyinput155), .A(n20951), .ZN(n20960) );
  AOI22_X1 U23903 ( .A1(n15040), .A2(keyinput244), .B1(n20955), .B2(
        keyinput248), .ZN(n20954) );
  OAI221_X1 U23904 ( .B1(n15040), .B2(keyinput244), .C1(n20955), .C2(
        keyinput248), .A(n20954), .ZN(n20959) );
  AOI22_X1 U23905 ( .A1(n21111), .A2(keyinput152), .B1(keyinput215), .B2(
        n20957), .ZN(n20956) );
  OAI221_X1 U23906 ( .B1(n21111), .B2(keyinput152), .C1(n20957), .C2(
        keyinput215), .A(n20956), .ZN(n20958) );
  NOR4_X1 U23907 ( .A1(n20961), .A2(n20960), .A3(n20959), .A4(n20958), .ZN(
        n21000) );
  INV_X1 U23908 ( .A(P3_DATAO_REG_26__SCAN_IN), .ZN(n21046) );
  XOR2_X1 U23909 ( .A(keyinput146), .B(n21046), .Z(n20966) );
  INV_X1 U23910 ( .A(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n20962) );
  XOR2_X1 U23911 ( .A(keyinput212), .B(n20962), .Z(n20965) );
  XNOR2_X1 U23912 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B(keyinput178), .ZN(
        n20964) );
  XNOR2_X1 U23913 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B(keyinput235), .ZN(
        n20963) );
  NAND4_X1 U23914 ( .A1(n20966), .A2(n20965), .A3(n20964), .A4(n20963), .ZN(
        n20972) );
  INV_X1 U23915 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n20968) );
  INV_X1 U23916 ( .A(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n21105) );
  AOI22_X1 U23917 ( .A1(n20968), .A2(keyinput147), .B1(n21105), .B2(
        keyinput232), .ZN(n20967) );
  OAI221_X1 U23918 ( .B1(n20968), .B2(keyinput147), .C1(n21105), .C2(
        keyinput232), .A(n20967), .ZN(n20971) );
  AOI22_X1 U23919 ( .A1(n21093), .A2(keyinput131), .B1(n21108), .B2(
        keyinput154), .ZN(n20969) );
  OAI221_X1 U23920 ( .B1(n21093), .B2(keyinput131), .C1(n21108), .C2(
        keyinput154), .A(n20969), .ZN(n20970) );
  NOR3_X1 U23921 ( .A1(n20972), .A2(n20971), .A3(n20970), .ZN(n20999) );
  INV_X1 U23922 ( .A(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n21082) );
  AOI22_X1 U23923 ( .A1(n21082), .A2(keyinput229), .B1(keyinput134), .B2(
        n20974), .ZN(n20973) );
  OAI221_X1 U23924 ( .B1(n21082), .B2(keyinput229), .C1(n20974), .C2(
        keyinput134), .A(n20973), .ZN(n20983) );
  AOI22_X1 U23925 ( .A1(n21078), .A2(keyinput243), .B1(n21095), .B2(
        keyinput140), .ZN(n20975) );
  OAI221_X1 U23926 ( .B1(n21078), .B2(keyinput243), .C1(n21095), .C2(
        keyinput140), .A(n20975), .ZN(n20982) );
  INV_X1 U23927 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n21087) );
  AOI22_X1 U23928 ( .A1(n20977), .A2(keyinput231), .B1(keyinput219), .B2(
        n21087), .ZN(n20976) );
  OAI221_X1 U23929 ( .B1(n20977), .B2(keyinput231), .C1(n21087), .C2(
        keyinput219), .A(n20976), .ZN(n20981) );
  AOI22_X1 U23930 ( .A1(n21188), .A2(keyinput233), .B1(keyinput218), .B2(
        n20979), .ZN(n20978) );
  OAI221_X1 U23931 ( .B1(n21188), .B2(keyinput233), .C1(n20979), .C2(
        keyinput218), .A(n20978), .ZN(n20980) );
  NOR4_X1 U23932 ( .A1(n20983), .A2(n20982), .A3(n20981), .A4(n20980), .ZN(
        n20998) );
  INV_X1 U23933 ( .A(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n20985) );
  AOI22_X1 U23934 ( .A1(n21103), .A2(keyinput214), .B1(n20985), .B2(
        keyinput246), .ZN(n20984) );
  OAI221_X1 U23935 ( .B1(n21103), .B2(keyinput214), .C1(n20985), .C2(
        keyinput246), .A(n20984), .ZN(n20996) );
  AOI22_X1 U23936 ( .A1(n21022), .A2(keyinput188), .B1(n21047), .B2(
        keyinput209), .ZN(n20986) );
  OAI221_X1 U23937 ( .B1(n21022), .B2(keyinput188), .C1(n21047), .C2(
        keyinput209), .A(n20986), .ZN(n20995) );
  AOI22_X1 U23938 ( .A1(n20989), .A2(keyinput217), .B1(keyinput150), .B2(
        n20988), .ZN(n20987) );
  OAI221_X1 U23939 ( .B1(n20989), .B2(keyinput217), .C1(n20988), .C2(
        keyinput150), .A(n20987), .ZN(n20994) );
  INV_X1 U23940 ( .A(P2_READREQUEST_REG_SCAN_IN), .ZN(n20992) );
  AOI22_X1 U23941 ( .A1(n20990), .A2(keyinput199), .B1(keyinput216), .B2(
        n20992), .ZN(n20991) );
  OAI221_X1 U23942 ( .B1(n20990), .B2(keyinput199), .C1(n20992), .C2(
        keyinput216), .A(n20991), .ZN(n20993) );
  NOR4_X1 U23943 ( .A1(n20996), .A2(n20995), .A3(n20994), .A4(n20993), .ZN(
        n20997) );
  NAND4_X1 U23944 ( .A1(n21000), .A2(n20999), .A3(n20998), .A4(n20997), .ZN(
        n21001) );
  NOR4_X1 U23945 ( .A1(n21004), .A2(n21003), .A3(n21002), .A4(n21001), .ZN(
        n21214) );
  AOI22_X1 U23946 ( .A1(n21007), .A2(keyinput72), .B1(keyinput70), .B2(n21006), 
        .ZN(n21005) );
  OAI221_X1 U23947 ( .B1(n21007), .B2(keyinput72), .C1(n21006), .C2(keyinput70), .A(n21005), .ZN(n21019) );
  AOI22_X1 U23948 ( .A1(n21010), .A2(keyinput58), .B1(keyinput25), .B2(n21009), 
        .ZN(n21008) );
  OAI221_X1 U23949 ( .B1(n21010), .B2(keyinput58), .C1(n21009), .C2(keyinput25), .A(n21008), .ZN(n21018) );
  INV_X1 U23950 ( .A(P3_DATAO_REG_16__SCAN_IN), .ZN(n21012) );
  AOI22_X1 U23951 ( .A1(n21012), .A2(keyinput125), .B1(n10721), .B2(keyinput96), .ZN(n21011) );
  OAI221_X1 U23952 ( .B1(n21012), .B2(keyinput125), .C1(n10721), .C2(
        keyinput96), .A(n21011), .ZN(n21017) );
  AOI22_X1 U23953 ( .A1(n21015), .A2(keyinput124), .B1(keyinput64), .B2(n21014), .ZN(n21013) );
  OAI221_X1 U23954 ( .B1(n21015), .B2(keyinput124), .C1(n21014), .C2(
        keyinput64), .A(n21013), .ZN(n21016) );
  NOR4_X1 U23955 ( .A1(n21019), .A2(n21018), .A3(n21017), .A4(n21016), .ZN(
        n21070) );
  AOI22_X1 U23956 ( .A1(n21022), .A2(keyinput60), .B1(n21021), .B2(keyinput66), 
        .ZN(n21020) );
  OAI221_X1 U23957 ( .B1(n21022), .B2(keyinput60), .C1(n21021), .C2(keyinput66), .A(n21020), .ZN(n21035) );
  INV_X1 U23958 ( .A(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n21024) );
  AOI22_X1 U23959 ( .A1(n21025), .A2(keyinput14), .B1(keyinput83), .B2(n21024), 
        .ZN(n21023) );
  OAI221_X1 U23960 ( .B1(n21025), .B2(keyinput14), .C1(n21024), .C2(keyinput83), .A(n21023), .ZN(n21034) );
  AOI22_X1 U23961 ( .A1(n21028), .A2(keyinput106), .B1(n21027), .B2(keyinput20), .ZN(n21026) );
  OAI221_X1 U23962 ( .B1(n21028), .B2(keyinput106), .C1(n21027), .C2(
        keyinput20), .A(n21026), .ZN(n21033) );
  AOI22_X1 U23963 ( .A1(n21031), .A2(keyinput35), .B1(n21030), .B2(keyinput67), 
        .ZN(n21029) );
  OAI221_X1 U23964 ( .B1(n21031), .B2(keyinput35), .C1(n21030), .C2(keyinput67), .A(n21029), .ZN(n21032) );
  NOR4_X1 U23965 ( .A1(n21035), .A2(n21034), .A3(n21033), .A4(n21032), .ZN(
        n21069) );
  AOI22_X1 U23966 ( .A1(n21038), .A2(keyinput43), .B1(n21037), .B2(keyinput92), 
        .ZN(n21036) );
  OAI221_X1 U23967 ( .B1(n21038), .B2(keyinput43), .C1(n21037), .C2(keyinput92), .A(n21036), .ZN(n21051) );
  AOI22_X1 U23968 ( .A1(n21041), .A2(keyinput31), .B1(keyinput114), .B2(n21040), .ZN(n21039) );
  OAI221_X1 U23969 ( .B1(n21041), .B2(keyinput31), .C1(n21040), .C2(
        keyinput114), .A(n21039), .ZN(n21050) );
  AOI22_X1 U23970 ( .A1(n21044), .A2(keyinput100), .B1(keyinput17), .B2(n21043), .ZN(n21042) );
  OAI221_X1 U23971 ( .B1(n21044), .B2(keyinput100), .C1(n21043), .C2(
        keyinput17), .A(n21042), .ZN(n21049) );
  AOI22_X1 U23972 ( .A1(n21047), .A2(keyinput81), .B1(keyinput18), .B2(n21046), 
        .ZN(n21045) );
  OAI221_X1 U23973 ( .B1(n21047), .B2(keyinput81), .C1(n21046), .C2(keyinput18), .A(n21045), .ZN(n21048) );
  NOR4_X1 U23974 ( .A1(n21051), .A2(n21050), .A3(n21049), .A4(n21048), .ZN(
        n21068) );
  AOI22_X1 U23975 ( .A1(n11933), .A2(keyinput49), .B1(keyinput113), .B2(n21053), .ZN(n21052) );
  OAI221_X1 U23976 ( .B1(n11933), .B2(keyinput49), .C1(n21053), .C2(
        keyinput113), .A(n21052), .ZN(n21066) );
  AOI22_X1 U23977 ( .A1(n21056), .A2(keyinput102), .B1(keyinput109), .B2(
        n21055), .ZN(n21054) );
  OAI221_X1 U23978 ( .B1(n21056), .B2(keyinput102), .C1(n21055), .C2(
        keyinput109), .A(n21054), .ZN(n21065) );
  INV_X1 U23979 ( .A(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n21059) );
  INV_X1 U23980 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n21058) );
  AOI22_X1 U23981 ( .A1(n21059), .A2(keyinput59), .B1(n21058), .B2(keyinput122), .ZN(n21057) );
  OAI221_X1 U23982 ( .B1(n21059), .B2(keyinput59), .C1(n21058), .C2(
        keyinput122), .A(n21057), .ZN(n21064) );
  XOR2_X1 U23983 ( .A(n21060), .B(keyinput69), .Z(n21062) );
  XNOR2_X1 U23984 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B(keyinput50), .ZN(
        n21061) );
  NAND2_X1 U23985 ( .A1(n21062), .A2(n21061), .ZN(n21063) );
  NOR4_X1 U23986 ( .A1(n21066), .A2(n21065), .A3(n21064), .A4(n21063), .ZN(
        n21067) );
  NAND4_X1 U23987 ( .A1(n21070), .A2(n21069), .A3(n21068), .A4(n21067), .ZN(
        n21213) );
  AOI22_X1 U23988 ( .A1(n11474), .A2(keyinput8), .B1(n21072), .B2(keyinput48), 
        .ZN(n21071) );
  OAI221_X1 U23989 ( .B1(n11474), .B2(keyinput8), .C1(n21072), .C2(keyinput48), 
        .A(n21071), .ZN(n21076) );
  XOR2_X1 U23990 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B(keyinput11), .Z(
        n21075) );
  XNOR2_X1 U23991 ( .A(n21073), .B(keyinput44), .ZN(n21074) );
  OR3_X1 U23992 ( .A1(n21076), .A2(n21075), .A3(n21074), .ZN(n21085) );
  AOI22_X1 U23993 ( .A1(n21079), .A2(keyinput38), .B1(keyinput115), .B2(n21078), .ZN(n21077) );
  OAI221_X1 U23994 ( .B1(n21079), .B2(keyinput38), .C1(n21078), .C2(
        keyinput115), .A(n21077), .ZN(n21084) );
  AOI22_X1 U23995 ( .A1(n21082), .A2(keyinput101), .B1(n21081), .B2(keyinput79), .ZN(n21080) );
  OAI221_X1 U23996 ( .B1(n21082), .B2(keyinput101), .C1(n21081), .C2(
        keyinput79), .A(n21080), .ZN(n21083) );
  NOR3_X1 U23997 ( .A1(n21085), .A2(n21084), .A3(n21083), .ZN(n21133) );
  AOI22_X1 U23998 ( .A1(n14410), .A2(keyinput45), .B1(n21087), .B2(keyinput91), 
        .ZN(n21086) );
  OAI221_X1 U23999 ( .B1(n14410), .B2(keyinput45), .C1(n21087), .C2(keyinput91), .A(n21086), .ZN(n21100) );
  INV_X1 U24000 ( .A(DATAI_26_), .ZN(n21090) );
  AOI22_X1 U24001 ( .A1(n21090), .A2(keyinput28), .B1(n21089), .B2(keyinput37), 
        .ZN(n21088) );
  OAI221_X1 U24002 ( .B1(n21090), .B2(keyinput28), .C1(n21089), .C2(keyinput37), .A(n21088), .ZN(n21099) );
  AOI22_X1 U24003 ( .A1(n21093), .A2(keyinput3), .B1(keyinput99), .B2(n21092), 
        .ZN(n21091) );
  OAI221_X1 U24004 ( .B1(n21093), .B2(keyinput3), .C1(n21092), .C2(keyinput99), 
        .A(n21091), .ZN(n21098) );
  AOI22_X1 U24005 ( .A1(n21096), .A2(keyinput30), .B1(n21095), .B2(keyinput12), 
        .ZN(n21094) );
  OAI221_X1 U24006 ( .B1(n21096), .B2(keyinput30), .C1(n21095), .C2(keyinput12), .A(n21094), .ZN(n21097) );
  NOR4_X1 U24007 ( .A1(n21100), .A2(n21099), .A3(n21098), .A4(n21097), .ZN(
        n21132) );
  AOI22_X1 U24008 ( .A1(n21103), .A2(keyinput86), .B1(keyinput76), .B2(n21102), 
        .ZN(n21101) );
  OAI221_X1 U24009 ( .B1(n21103), .B2(keyinput86), .C1(n21102), .C2(keyinput76), .A(n21101), .ZN(n21115) );
  INV_X1 U24010 ( .A(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n21106) );
  AOI22_X1 U24011 ( .A1(n21106), .A2(keyinput80), .B1(n21105), .B2(keyinput104), .ZN(n21104) );
  OAI221_X1 U24012 ( .B1(n21106), .B2(keyinput80), .C1(n21105), .C2(
        keyinput104), .A(n21104), .ZN(n21114) );
  AOI22_X1 U24013 ( .A1(n21109), .A2(keyinput32), .B1(keyinput26), .B2(n21108), 
        .ZN(n21107) );
  OAI221_X1 U24014 ( .B1(n21109), .B2(keyinput32), .C1(n21108), .C2(keyinput26), .A(n21107), .ZN(n21113) );
  AOI22_X1 U24015 ( .A1(n21111), .A2(keyinput24), .B1(n11939), .B2(keyinput53), 
        .ZN(n21110) );
  OAI221_X1 U24016 ( .B1(n21111), .B2(keyinput24), .C1(n11939), .C2(keyinput53), .A(n21110), .ZN(n21112) );
  NOR4_X1 U24017 ( .A1(n21115), .A2(n21114), .A3(n21113), .A4(n21112), .ZN(
        n21131) );
  AOI22_X1 U24018 ( .A1(n21118), .A2(keyinput78), .B1(keyinput9), .B2(n21117), 
        .ZN(n21116) );
  OAI221_X1 U24019 ( .B1(n21118), .B2(keyinput78), .C1(n21117), .C2(keyinput9), 
        .A(n21116), .ZN(n21129) );
  INV_X1 U24020 ( .A(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n21120) );
  AOI22_X1 U24021 ( .A1(n11312), .A2(keyinput21), .B1(keyinput51), .B2(n21120), 
        .ZN(n21119) );
  OAI221_X1 U24022 ( .B1(n11312), .B2(keyinput21), .C1(n21120), .C2(keyinput51), .A(n21119), .ZN(n21128) );
  AOI22_X1 U24023 ( .A1(n11037), .A2(keyinput16), .B1(keyinput1), .B2(n21122), 
        .ZN(n21121) );
  OAI221_X1 U24024 ( .B1(n11037), .B2(keyinput16), .C1(n21122), .C2(keyinput1), 
        .A(n21121), .ZN(n21127) );
  AOI22_X1 U24025 ( .A1(n21125), .A2(keyinput121), .B1(n21124), .B2(keyinput98), .ZN(n21123) );
  OAI221_X1 U24026 ( .B1(n21125), .B2(keyinput121), .C1(n21124), .C2(
        keyinput98), .A(n21123), .ZN(n21126) );
  NOR4_X1 U24027 ( .A1(n21129), .A2(n21128), .A3(n21127), .A4(n21126), .ZN(
        n21130) );
  NAND4_X1 U24028 ( .A1(n21133), .A2(n21132), .A3(n21131), .A4(n21130), .ZN(
        n21212) );
  AOI22_X1 U24029 ( .A1(P3_DATAO_REG_8__SCAN_IN), .A2(keyinput77), .B1(
        P3_REIP_REG_11__SCAN_IN), .B2(keyinput40), .ZN(n21134) );
  OAI221_X1 U24030 ( .B1(P3_DATAO_REG_8__SCAN_IN), .B2(keyinput77), .C1(
        P3_REIP_REG_11__SCAN_IN), .C2(keyinput40), .A(n21134), .ZN(n21141) );
  AOI22_X1 U24031 ( .A1(P1_EAX_REG_20__SCAN_IN), .A2(keyinput95), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(keyinput75), .ZN(n21135) );
  OAI221_X1 U24032 ( .B1(P1_EAX_REG_20__SCAN_IN), .B2(keyinput95), .C1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(keyinput75), .A(n21135), .ZN(
        n21140) );
  AOI22_X1 U24033 ( .A1(P2_ADDRESS_REG_28__SCAN_IN), .A2(keyinput120), .B1(
        P2_INSTQUEUE_REG_9__1__SCAN_IN), .B2(keyinput85), .ZN(n21136) );
  OAI221_X1 U24034 ( .B1(P2_ADDRESS_REG_28__SCAN_IN), .B2(keyinput120), .C1(
        P2_INSTQUEUE_REG_9__1__SCAN_IN), .C2(keyinput85), .A(n21136), .ZN(
        n21139) );
  AOI22_X1 U24035 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(keyinput110), 
        .B1(P2_ADDRESS_REG_15__SCAN_IN), .B2(keyinput119), .ZN(n21137) );
  OAI221_X1 U24036 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(keyinput110), 
        .C1(P2_ADDRESS_REG_15__SCAN_IN), .C2(keyinput119), .A(n21137), .ZN(
        n21138) );
  NOR4_X1 U24037 ( .A1(n21141), .A2(n21140), .A3(n21139), .A4(n21138), .ZN(
        n21210) );
  AOI22_X1 U24038 ( .A1(P2_UWORD_REG_1__SCAN_IN), .A2(keyinput19), .B1(
        DATAI_9_), .B2(keyinput29), .ZN(n21142) );
  OAI221_X1 U24039 ( .B1(P2_UWORD_REG_1__SCAN_IN), .B2(keyinput19), .C1(
        DATAI_9_), .C2(keyinput29), .A(n21142), .ZN(n21149) );
  AOI22_X1 U24040 ( .A1(P2_REIP_REG_28__SCAN_IN), .A2(keyinput112), .B1(
        P2_INSTQUEUE_REG_10__5__SCAN_IN), .B2(keyinput107), .ZN(n21143) );
  OAI221_X1 U24041 ( .B1(P2_REIP_REG_28__SCAN_IN), .B2(keyinput112), .C1(
        P2_INSTQUEUE_REG_10__5__SCAN_IN), .C2(keyinput107), .A(n21143), .ZN(
        n21148) );
  AOI22_X1 U24042 ( .A1(P3_ADDRESS_REG_10__SCAN_IN), .A2(keyinput87), .B1(
        P2_EAX_REG_26__SCAN_IN), .B2(keyinput82), .ZN(n21144) );
  OAI221_X1 U24043 ( .B1(P3_ADDRESS_REG_10__SCAN_IN), .B2(keyinput87), .C1(
        P2_EAX_REG_26__SCAN_IN), .C2(keyinput82), .A(n21144), .ZN(n21147) );
  AOI22_X1 U24044 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(keyinput89), .B1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(keyinput33), .ZN(n21145) );
  OAI221_X1 U24045 ( .B1(P3_DATAWIDTH_REG_30__SCAN_IN), .B2(keyinput89), .C1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C2(keyinput33), .A(n21145), .ZN(
        n21146) );
  NOR4_X1 U24046 ( .A1(n21149), .A2(n21148), .A3(n21147), .A4(n21146), .ZN(
        n21209) );
  OAI22_X1 U24047 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(keyinput127), .B1(
        keyinput61), .B2(P1_LWORD_REG_5__SCAN_IN), .ZN(n21150) );
  AOI221_X1 U24048 ( .B1(P1_UWORD_REG_6__SCAN_IN), .B2(keyinput127), .C1(
        P1_LWORD_REG_5__SCAN_IN), .C2(keyinput61), .A(n21150), .ZN(n21157) );
  OAI22_X1 U24049 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(keyinput56), 
        .B1(P2_LWORD_REG_7__SCAN_IN), .B2(keyinput52), .ZN(n21151) );
  AOI221_X1 U24050 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(keyinput56), 
        .C1(keyinput52), .C2(P2_LWORD_REG_7__SCAN_IN), .A(n21151), .ZN(n21156)
         );
  OAI22_X1 U24051 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(keyinput0), 
        .B1(keyinput27), .B2(P3_REIP_REG_6__SCAN_IN), .ZN(n21152) );
  AOI221_X1 U24052 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(keyinput0), 
        .C1(P3_REIP_REG_6__SCAN_IN), .C2(keyinput27), .A(n21152), .ZN(n21155)
         );
  OAI22_X1 U24053 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(keyinput126), 
        .B1(keyinput108), .B2(DATAI_29_), .ZN(n21153) );
  AOI221_X1 U24054 ( .B1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B2(keyinput126), 
        .C1(DATAI_29_), .C2(keyinput108), .A(n21153), .ZN(n21154) );
  NAND4_X1 U24055 ( .A1(n21157), .A2(n21156), .A3(n21155), .A4(n21154), .ZN(
        n21207) );
  OAI22_X1 U24056 ( .A1(BUF2_REG_31__SCAN_IN), .A2(keyinput6), .B1(
        P1_DATAWIDTH_REG_22__SCAN_IN), .B2(keyinput39), .ZN(n21158) );
  AOI221_X1 U24057 ( .B1(BUF2_REG_31__SCAN_IN), .B2(keyinput6), .C1(keyinput39), .C2(P1_DATAWIDTH_REG_22__SCAN_IN), .A(n21158), .ZN(n21165) );
  OAI22_X1 U24058 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(keyinput15), .B1(
        P3_DATAO_REG_23__SCAN_IN), .B2(keyinput2), .ZN(n21159) );
  AOI221_X1 U24059 ( .B1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B2(keyinput15), 
        .C1(keyinput2), .C2(P3_DATAO_REG_23__SCAN_IN), .A(n21159), .ZN(n21164)
         );
  OAI22_X1 U24060 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(keyinput116), 
        .B1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B2(keyinput118), .ZN(n21160) );
  AOI221_X1 U24061 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(keyinput116), 
        .C1(keyinput118), .C2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A(n21160), 
        .ZN(n21163) );
  OAI22_X1 U24062 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(keyinput23), 
        .B1(P3_DATAWIDTH_REG_26__SCAN_IN), .B2(keyinput41), .ZN(n21161) );
  AOI221_X1 U24063 ( .B1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(keyinput23), 
        .C1(keyinput41), .C2(P3_DATAWIDTH_REG_26__SCAN_IN), .A(n21161), .ZN(
        n21162) );
  NAND4_X1 U24064 ( .A1(n21165), .A2(n21164), .A3(n21163), .A4(n21162), .ZN(
        n21206) );
  AOI22_X1 U24065 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(keyinput5), .B1(
        P3_REIP_REG_13__SCAN_IN), .B2(keyinput57), .ZN(n21166) );
  OAI221_X1 U24066 ( .B1(P1_DATAWIDTH_REG_31__SCAN_IN), .B2(keyinput5), .C1(
        P3_REIP_REG_13__SCAN_IN), .C2(keyinput57), .A(n21166), .ZN(n21173) );
  AOI22_X1 U24067 ( .A1(P2_READREQUEST_REG_SCAN_IN), .A2(keyinput88), .B1(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(keyinput10), .ZN(n21167) );
  OAI221_X1 U24068 ( .B1(P2_READREQUEST_REG_SCAN_IN), .B2(keyinput88), .C1(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(keyinput10), .A(n21167), .ZN(
        n21172) );
  AOI22_X1 U24069 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(keyinput54), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(keyinput123), .ZN(n21168) );
  OAI221_X1 U24070 ( .B1(P1_DATAO_REG_5__SCAN_IN), .B2(keyinput54), .C1(
        P1_EAX_REG_25__SCAN_IN), .C2(keyinput123), .A(n21168), .ZN(n21171) );
  AOI22_X1 U24071 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(keyinput34), .B1(
        P3_INSTQUEUE_REG_10__4__SCAN_IN), .B2(keyinput111), .ZN(n21169) );
  OAI221_X1 U24072 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(keyinput34), .C1(
        P3_INSTQUEUE_REG_10__4__SCAN_IN), .C2(keyinput111), .A(n21169), .ZN(
        n21170) );
  NOR4_X1 U24073 ( .A1(n21173), .A2(n21172), .A3(n21171), .A4(n21170), .ZN(
        n21204) );
  AOI22_X1 U24074 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(keyinput94), .B1(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(keyinput42), .ZN(n21174) );
  OAI221_X1 U24075 ( .B1(P1_LWORD_REG_1__SCAN_IN), .B2(keyinput94), .C1(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .C2(keyinput42), .A(n21174), .ZN(
        n21181) );
  AOI22_X1 U24076 ( .A1(P1_DATAO_REG_31__SCAN_IN), .A2(keyinput47), .B1(
        P2_INSTQUEUE_REG_14__2__SCAN_IN), .B2(keyinput68), .ZN(n21175) );
  OAI221_X1 U24077 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(keyinput47), .C1(
        P2_INSTQUEUE_REG_14__2__SCAN_IN), .C2(keyinput68), .A(n21175), .ZN(
        n21180) );
  AOI22_X1 U24078 ( .A1(BUF1_REG_1__SCAN_IN), .A2(keyinput36), .B1(
        P2_EBX_REG_9__SCAN_IN), .B2(keyinput62), .ZN(n21176) );
  OAI221_X1 U24079 ( .B1(BUF1_REG_1__SCAN_IN), .B2(keyinput36), .C1(
        P2_EBX_REG_9__SCAN_IN), .C2(keyinput62), .A(n21176), .ZN(n21179) );
  AOI22_X1 U24080 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(keyinput13), .B1(
        P3_REIP_REG_24__SCAN_IN), .B2(keyinput63), .ZN(n21177) );
  OAI221_X1 U24081 ( .B1(P3_DATAWIDTH_REG_19__SCAN_IN), .B2(keyinput13), .C1(
        P3_REIP_REG_24__SCAN_IN), .C2(keyinput63), .A(n21177), .ZN(n21178) );
  NOR4_X1 U24082 ( .A1(n21181), .A2(n21180), .A3(n21179), .A4(n21178), .ZN(
        n21203) );
  AOI22_X1 U24083 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(keyinput4), 
        .B1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B2(keyinput84), .ZN(n21182) );
  OAI221_X1 U24084 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(keyinput4), 
        .C1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .C2(keyinput84), .A(n21182), 
        .ZN(n21192) );
  AOI22_X1 U24085 ( .A1(P2_EAX_REG_2__SCAN_IN), .A2(keyinput74), .B1(
        P2_STATE2_REG_3__SCAN_IN), .B2(keyinput71), .ZN(n21183) );
  OAI221_X1 U24086 ( .B1(P2_EAX_REG_2__SCAN_IN), .B2(keyinput74), .C1(
        P2_STATE2_REG_3__SCAN_IN), .C2(keyinput71), .A(n21183), .ZN(n21191) );
  AOI22_X1 U24087 ( .A1(n21186), .A2(keyinput73), .B1(n21185), .B2(keyinput65), 
        .ZN(n21184) );
  OAI221_X1 U24088 ( .B1(n21186), .B2(keyinput73), .C1(n21185), .C2(keyinput65), .A(n21184), .ZN(n21190) );
  AOI22_X1 U24089 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(keyinput22), .B1(
        n21188), .B2(keyinput105), .ZN(n21187) );
  OAI221_X1 U24090 ( .B1(P1_DATAWIDTH_REG_28__SCAN_IN), .B2(keyinput22), .C1(
        n21188), .C2(keyinput105), .A(n21187), .ZN(n21189) );
  NOR4_X1 U24091 ( .A1(n21192), .A2(n21191), .A3(n21190), .A4(n21189), .ZN(
        n21202) );
  AOI22_X1 U24092 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(keyinput117), .B1(
        P2_INSTQUEUE_REG_11__2__SCAN_IN), .B2(keyinput97), .ZN(n21193) );
  OAI221_X1 U24093 ( .B1(P3_DATAWIDTH_REG_18__SCAN_IN), .B2(keyinput117), .C1(
        P2_INSTQUEUE_REG_11__2__SCAN_IN), .C2(keyinput97), .A(n21193), .ZN(
        n21200) );
  AOI22_X1 U24094 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(keyinput103), 
        .B1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B2(keyinput93), .ZN(n21194) );
  OAI221_X1 U24095 ( .B1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(keyinput103), 
        .C1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .C2(keyinput93), .A(n21194), 
        .ZN(n21199) );
  AOI22_X1 U24096 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(keyinput90), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(keyinput55), .ZN(n21195) );
  OAI221_X1 U24097 ( .B1(P3_DATAWIDTH_REG_8__SCAN_IN), .B2(keyinput90), .C1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .C2(keyinput55), .A(n21195), .ZN(
        n21198) );
  AOI22_X1 U24098 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(keyinput46), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(keyinput7), .ZN(n21196) );
  OAI221_X1 U24099 ( .B1(P1_UWORD_REG_12__SCAN_IN), .B2(keyinput46), .C1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .C2(keyinput7), .A(n21196), .ZN(
        n21197) );
  NOR4_X1 U24100 ( .A1(n21200), .A2(n21199), .A3(n21198), .A4(n21197), .ZN(
        n21201) );
  NAND4_X1 U24101 ( .A1(n21204), .A2(n21203), .A3(n21202), .A4(n21201), .ZN(
        n21205) );
  NOR3_X1 U24102 ( .A1(n21207), .A2(n21206), .A3(n21205), .ZN(n21208) );
  NAND3_X1 U24103 ( .A1(n21210), .A2(n21209), .A3(n21208), .ZN(n21211) );
  NOR4_X1 U24104 ( .A1(n21214), .A2(n21213), .A3(n21212), .A4(n21211), .ZN(
        n21217) );
  AOI22_X1 U24105 ( .A1(n21215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(U215), .ZN(n21216) );
  XNOR2_X1 U24106 ( .A(n21217), .B(n21216), .ZN(U261) );
  AND2_X2 U15406 ( .A1(n12265), .A2(n13740), .ZN(n13045) );
  AND2_X1 U11711 ( .A1(n12273), .A2(n13739), .ZN(n12489) );
  XNOR2_X1 U11320 ( .A(n13170), .B(n12475), .ZN(n12515) );
  CLKBUF_X1 U11304 ( .A(n13045), .Z(n12983) );
  CLKBUF_X2 U11324 ( .A(n10548), .Z(n14539) );
  CLKBUF_X1 U11339 ( .A(n10672), .Z(n11190) );
  CLKBUF_X1 U11367 ( .A(n10438), .Z(n19860) );
  CLKBUF_X1 U11613 ( .A(n10407), .Z(n19160) );
  CLKBUF_X1 U11790 ( .A(n17447), .Z(n17455) );
endmodule

