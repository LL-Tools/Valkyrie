

module b21_C_gen_AntiSAT_k_128_2 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2, 
        keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7, 
        keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12, 
        keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17, 
        keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22, 
        keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27, 
        keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32, 
        keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37, 
        keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42, 
        keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47, 
        keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52, 
        keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57, 
        keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62, 
        keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3, 
        keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8, 
        keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13, 
        keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18, 
        keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23, 
        keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28, 
        keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33, 
        keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38, 
        keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43, 
        keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48, 
        keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53, 
        keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58, 
        keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63, 
        ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, 
        ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, 
        ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, 
        ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, 
        U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, 
        P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, 
        P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, 
        P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, 
        P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, 
        P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, 
        P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, 
        P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, 
        P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, 
        P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, 
        P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, 
        P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, 
        P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, 
        P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, 
        P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, 
        P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, 
        P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, 
        P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, 
        P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, 
        P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, 
        P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, 
        P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, 
        P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, 
        P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, 
        P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, 
        P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, 
        P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, 
        P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, 
        P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, 
        P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, 
        P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, 
        P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, 
        P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, 
        P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, 
        P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, 
        P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, 
        P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, 
        P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10130;

  INV_X1 U4815 ( .A(P1_STATE_REG_SCAN_IN), .ZN(n10130) );
  OAI21_X1 U4816 ( .B1(n7860), .B2(n4602), .A(n4601), .ZN(n7921) );
  NAND2_X1 U4817 ( .A1(n5201), .A2(n5200), .ZN(n8306) );
  INV_X1 U4819 ( .A(n5519), .ZN(n8252) );
  NAND4_X2 U4820 ( .A1(n4337), .A2(n5657), .A3(n5656), .A4(n5655), .ZN(n6259)
         );
  CLKBUF_X2 U4821 ( .A(n5075), .Z(n4315) );
  INV_X1 U4824 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U4825 ( .A(n8245), .ZN(n4583) );
  NAND2_X1 U4826 ( .A1(n7339), .A2(n4415), .ZN(n5024) );
  INV_X2 U4827 ( .A(n6117), .ZN(n5770) );
  NOR2_X1 U4828 ( .A1(n9262), .A2(n9261), .ZN(n9264) );
  NAND2_X1 U4829 ( .A1(n5110), .A2(n4916), .ZN(n4706) );
  OR2_X1 U4830 ( .A1(n8305), .A2(n5232), .ZN(n7500) );
  NAND2_X1 U4831 ( .A1(n7024), .A2(n8091), .ZN(n5510) );
  INV_X1 U4832 ( .A(n5677), .ZN(n6466) );
  NOR2_X1 U4833 ( .A1(n9230), .A2(n9228), .ZN(n9235) );
  XNOR2_X1 U4834 ( .A(n4911), .B(SI_5_), .ZN(n5074) );
  NAND2_X1 U4835 ( .A1(n4349), .A2(n5001), .ZN(n10003) );
  NAND2_X1 U4836 ( .A1(n4685), .A2(n4684), .ZN(n8348) );
  OAI22_X1 U4837 ( .A1(n7560), .A2(n5838), .B1(n7558), .B2(n7557), .ZN(n7692)
         );
  NAND2_X2 U4839 ( .A1(n5589), .A2(n5590), .ZN(n5675) );
  AOI21_X2 U4840 ( .B1(n8348), .B2(n5295), .A(n8347), .ZN(n8356) );
  OR2_X1 U4841 ( .A1(n6222), .A2(n9745), .ZN(n9054) );
  INV_X1 U4842 ( .A(n5675), .ZN(n6235) );
  NAND2_X1 U4843 ( .A1(n6662), .A2(n4968), .ZN(n4313) );
  NAND2_X2 U4844 ( .A1(n4887), .A2(n4886), .ZN(n4888) );
  NAND2_X2 U4845 ( .A1(n7659), .A2(n4686), .ZN(n4685) );
  NAND2_X2 U4846 ( .A1(n8336), .A2(n5163), .ZN(n7359) );
  NAND2_X2 U4847 ( .A1(n7660), .A2(n5271), .ZN(n7659) );
  XNOR2_X2 U4848 ( .A(n5273), .B(n5272), .ZN(n7660) );
  NAND2_X2 U4849 ( .A1(n7588), .A2(n5257), .ZN(n5273) );
  XNOR2_X2 U4850 ( .A(n6259), .B(n9936), .ZN(n7175) );
  INV_X4 U4851 ( .A(n6470), .ZN(n5636) );
  NAND2_X2 U4852 ( .A1(n8051), .A2(n8320), .ZN(n6470) );
  OR2_X2 U4853 ( .A1(n4854), .A2(n5093), .ZN(n4501) );
  NAND2_X1 U4855 ( .A1(n4522), .A2(n4520), .ZN(n8492) );
  INV_X4 U4856 ( .A(n6118), .ZN(n6179) );
  INV_X4 U4857 ( .A(n7167), .ZN(n6191) );
  XNOR2_X1 U4858 ( .A(n5024), .B(n10003), .ZN(n5012) );
  INV_X8 U4859 ( .A(n4968), .ZN(n6667) );
  INV_X2 U4860 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  AOI21_X1 U4861 ( .B1(n4343), .B2(n8292), .A(n8291), .ZN(n8297) );
  OAI21_X1 U4862 ( .B1(n6481), .B2(n6586), .A(n4367), .ZN(n6486) );
  OAI21_X1 U4863 ( .B1(n8492), .B2(n8490), .A(n4420), .ZN(n4419) );
  AOI21_X1 U4864 ( .B1(n6330), .B2(n9919), .A(n6329), .ZN(n8337) );
  AND2_X1 U4865 ( .A1(n4736), .A2(n4732), .ZN(n9012) );
  AND2_X1 U4866 ( .A1(n4614), .A2(n4613), .ZN(n9339) );
  NAND2_X1 U4867 ( .A1(n9011), .A2(n6122), .ZN(n8978) );
  OR2_X1 U4868 ( .A1(n8951), .A2(n8952), .ZN(n4736) );
  XNOR2_X1 U4869 ( .A(n4471), .B(n8066), .ZN(n8844) );
  NAND2_X1 U4870 ( .A1(n9030), .A2(n9033), .ZN(n6102) );
  NAND2_X1 U4871 ( .A1(n6100), .A2(n6099), .ZN(n9031) );
  NAND2_X1 U4872 ( .A1(n5549), .A2(n5548), .ZN(n8840) );
  NOR2_X1 U4873 ( .A1(n9264), .A2(n6316), .ZN(n9252) );
  NAND2_X1 U4874 ( .A1(n6315), .A2(n6528), .ZN(n9283) );
  NAND2_X1 U4875 ( .A1(n4606), .A2(n6572), .ZN(n9297) );
  NAND2_X1 U4876 ( .A1(n4421), .A2(n5272), .ZN(n5274) );
  NAND2_X1 U4877 ( .A1(n5394), .A2(n5393), .ZN(n8869) );
  AND2_X1 U4878 ( .A1(n9278), .A2(n9268), .ZN(n9269) );
  OAI21_X1 U4879 ( .B1(n4744), .B2(n4340), .A(n4475), .ZN(n5937) );
  OAI21_X1 U4880 ( .B1(n5385), .B2(n5384), .A(n5386), .ZN(n5407) );
  NAND2_X1 U4881 ( .A1(n4738), .A2(n4737), .ZN(n7520) );
  NAND2_X1 U4882 ( .A1(n7921), .A2(n7920), .ZN(n7919) );
  AND2_X1 U4883 ( .A1(n7308), .A2(n4739), .ZN(n4738) );
  INV_X1 U4884 ( .A(n9747), .ZN(n8048) );
  NAND2_X1 U4885 ( .A1(n5908), .A2(n5907), .ZN(n9407) );
  NAND2_X1 U4886 ( .A1(n5244), .A2(n5243), .ZN(n8177) );
  AND2_X1 U4887 ( .A1(n6391), .A2(n6540), .ZN(n9705) );
  NAND2_X1 U4888 ( .A1(n5887), .A2(n5886), .ZN(n9717) );
  NAND2_X1 U4889 ( .A1(n5863), .A2(n5862), .ZN(n9411) );
  NAND2_X1 U4890 ( .A1(n5842), .A2(n5841), .ZN(n9759) );
  NAND2_X1 U4891 ( .A1(n5172), .A2(n5171), .ZN(n7676) );
  NAND2_X1 U4892 ( .A1(n4473), .A2(n5133), .ZN(n8419) );
  NAND2_X1 U4893 ( .A1(n5533), .A2(n5512), .ZN(n8490) );
  INV_X2 U4894 ( .A(n10070), .ZN(n4316) );
  AND2_X1 U4895 ( .A1(n5761), .A2(n5760), .ZN(n9960) );
  NAND4_X1 U4896 ( .A1(n5641), .A2(n5640), .A3(n5639), .A4(n5638), .ZN(n6258)
         );
  NAND2_X2 U4897 ( .A1(n6299), .A2(n6238), .ZN(n7167) );
  INV_X1 U4898 ( .A(n5024), .ZN(n5309) );
  OR2_X2 U4899 ( .A1(n7163), .A2(n5644), .ZN(n6118) );
  NAND2_X1 U4900 ( .A1(n8252), .A2(n8815), .ZN(n8293) );
  NAND2_X1 U4901 ( .A1(n8320), .A2(n5590), .ZN(n5677) );
  OR2_X1 U4902 ( .A1(n7024), .A2(n8815), .ZN(n8285) );
  AOI21_X1 U4903 ( .B1(n4910), .B2(n4431), .A(n4348), .ZN(n4430) );
  NAND2_X2 U4904 ( .A1(n8936), .A2(n4866), .ZN(n5046) );
  XNOR2_X1 U4905 ( .A(n4877), .B(n4876), .ZN(n8091) );
  INV_X1 U4906 ( .A(n8939), .ZN(n4866) );
  NAND2_X1 U4907 ( .A1(n4883), .A2(n4882), .ZN(n8815) );
  OR2_X1 U4908 ( .A1(n9433), .A2(n5586), .ZN(n5588) );
  NAND2_X1 U4909 ( .A1(n4881), .A2(n4880), .ZN(n4883) );
  OR2_X1 U4910 ( .A1(n4973), .A2(n4969), .ZN(n4978) );
  AND2_X1 U4911 ( .A1(n4853), .A2(n4663), .ZN(n8939) );
  MUX2_X1 U4912 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5616), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5618) );
  MUX2_X1 U4913 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4970), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n4972) );
  NAND2_X2 U4914 ( .A1(n6667), .A2(n10130), .ZN(n9443) );
  AND2_X1 U4915 ( .A1(n4870), .A2(n4847), .ZN(n4546) );
  NAND4_X1 U4916 ( .A1(n4814), .A2(n4418), .A3(n4417), .A4(n4416), .ZN(n5055)
         );
  AND4_X1 U4917 ( .A1(n5572), .A2(n5571), .A3(n5570), .A4(n5569), .ZN(n5575)
         );
  NOR2_X1 U4918 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(n4341), .ZN(n4828) );
  AND2_X1 U4919 ( .A1(n4783), .A2(n6218), .ZN(n4781) );
  NOR2_X1 U4920 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5569) );
  NOR2_X1 U4921 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5570) );
  NOR2_X1 U4922 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5571) );
  INV_X1 U4923 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4783) );
  INV_X1 U4924 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5904) );
  NOR2_X1 U4925 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5619) );
  INV_X1 U4926 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4814) );
  INV_X1 U4927 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4416) );
  INV_X1 U4928 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4417) );
  INV_X1 U4929 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4418) );
  INV_X1 U4930 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5112) );
  NOR2_X1 U4931 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5576) );
  INV_X1 U4932 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5168) );
  INV_X1 U4933 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5166) );
  INV_X1 U4934 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5240) );
  INV_X1 U4935 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5237) );
  NOR2_X1 U4936 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n4842) );
  NOR3_X1 U4937 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .A3(
        P2_IR_REG_16__SCAN_IN), .ZN(n4841) );
  INV_X1 U4938 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5605) );
  AND2_X1 U4939 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n9656) );
  NOR2_X1 U4940 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5573) );
  XNOR2_X2 U4941 ( .A(n4647), .B(n5614), .ZN(n6323) );
  NAND2_X4 U4942 ( .A1(n8949), .A2(n5534), .ZN(n5006) );
  OR2_X2 U4943 ( .A1(n7681), .A2(n7367), .ZN(n7729) );
  NAND2_X2 U4944 ( .A1(n5186), .A2(n5185), .ZN(n7367) );
  INV_X4 U4945 ( .A(n4313), .ZN(n4317) );
  INV_X4 U4946 ( .A(n5044), .ZN(n4983) );
  INV_X1 U4947 ( .A(n5658), .ZN(n4318) );
  XNOR2_X2 U4948 ( .A(n5491), .B(n5490), .ZN(n7024) );
  INV_X1 U4949 ( .A(n5046), .ZN(n4319) );
  INV_X4 U4950 ( .A(n5046), .ZN(n5025) );
  INV_X1 U4951 ( .A(n5315), .ZN(n4320) );
  NAND2_X1 U4952 ( .A1(n8939), .A2(n4865), .ZN(n5315) );
  NAND2_X1 U4953 ( .A1(n8672), .A2(n8279), .ZN(n4499) );
  NAND2_X1 U4954 ( .A1(n5113), .A2(n4426), .ZN(n4427) );
  AND2_X1 U4955 ( .A1(n4870), .A2(n4372), .ZN(n4426) );
  OR2_X1 U4956 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n4873) );
  NAND2_X1 U4957 ( .A1(n6216), .A2(n9222), .ZN(n6299) );
  NOR2_X1 U4958 ( .A1(n5535), .A2(n10027), .ZN(n5533) );
  NAND2_X1 U4959 ( .A1(n5006), .A2(n4968), .ZN(n5044) );
  AOI21_X1 U4960 ( .B1(n8199), .B2(n8198), .A(n4565), .ZN(n4564) );
  INV_X1 U4961 ( .A(n8275), .ZN(n4565) );
  AOI21_X1 U4962 ( .B1(n8199), .B2(n8197), .A(n4569), .ZN(n4568) );
  INV_X1 U4963 ( .A(n8747), .ZN(n4569) );
  INV_X1 U4964 ( .A(n4708), .ZN(n4707) );
  OAI21_X1 U4965 ( .B1(n6444), .B2(n6442), .A(n6439), .ZN(n4708) );
  NOR2_X1 U4966 ( .A1(n4577), .A2(n8376), .ZN(n4576) );
  NOR2_X1 U4967 ( .A1(n4579), .A2(n4578), .ZN(n4577) );
  NOR2_X1 U4968 ( .A1(n4581), .A2(n4580), .ZN(n4579) );
  INV_X1 U4969 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5596) );
  NOR2_X1 U4970 ( .A1(n4952), .A2(n4528), .ZN(n4527) );
  INV_X1 U4971 ( .A(n4951), .ZN(n4528) );
  AOI21_X1 U4972 ( .B1(n4514), .B2(n4924), .A(n4512), .ZN(n4511) );
  INV_X1 U4973 ( .A(n5146), .ZN(n4512) );
  INV_X1 U4974 ( .A(SI_10_), .ZN(n9579) );
  OAI22_X1 U4975 ( .A1(n8425), .A2(n4679), .B1(n5359), .B2(n5360), .ZN(n4678)
         );
  AOI21_X1 U4976 ( .B1(n8619), .B2(n4805), .A(n4366), .ZN(n4804) );
  INV_X1 U4977 ( .A(n8375), .ZN(n4805) );
  OR2_X1 U4978 ( .A1(n8860), .A2(n8693), .ZN(n8217) );
  INV_X1 U4979 ( .A(n4468), .ZN(n4467) );
  OAI21_X1 U4980 ( .B1(n4338), .B2(n4469), .A(n8361), .ZN(n4468) );
  INV_X1 U4981 ( .A(n8269), .ZN(n4820) );
  OR2_X1 U4982 ( .A1(n8306), .A2(n8510), .ZN(n4819) );
  OAI22_X1 U4983 ( .A1(n7403), .A2(n6117), .B1(n7160), .B2(n6118), .ZN(n5712)
         );
  XNOR2_X1 U4984 ( .A(n5588), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5590) );
  OR2_X1 U4985 ( .A1(n9341), .A2(n9063), .ZN(n9166) );
  INV_X1 U4986 ( .A(n4771), .ZN(n4770) );
  AND2_X1 U4987 ( .A1(n9379), .A2(n8972), .ZN(n6491) );
  NAND2_X1 U4988 ( .A1(n9660), .A2(n9915), .ZN(n6377) );
  OR2_X1 U4989 ( .A1(n9660), .A2(n9915), .ZN(n6557) );
  OR2_X1 U4990 ( .A1(n6216), .A2(n4743), .ZN(n6300) );
  NAND2_X1 U4991 ( .A1(n6295), .A2(n6294), .ZN(n6446) );
  NAND2_X1 U4992 ( .A1(n5460), .A2(n5459), .ZN(n5545) );
  NAND2_X1 U4993 ( .A1(n5409), .A2(n5408), .ZN(n5422) );
  NAND2_X1 U4994 ( .A1(n5407), .A2(n5406), .ZN(n5409) );
  INV_X1 U4995 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6218) );
  NAND2_X1 U4996 ( .A1(n5366), .A2(n5365), .ZN(n5385) );
  OR2_X1 U4997 ( .A1(n5363), .A2(n5362), .ZN(n5366) );
  INV_X1 U4998 ( .A(SI_17_), .ZN(n4964) );
  AND2_X1 U4999 ( .A1(n5884), .A2(n5596), .ZN(n5973) );
  AND2_X1 U5000 ( .A1(n4963), .A2(n4962), .ZN(n4982) );
  INV_X1 U5001 ( .A(n5273), .ZN(n4421) );
  XNOR2_X1 U5002 ( .A(n5309), .B(n4425), .ZN(n7700) );
  NAND2_X1 U5003 ( .A1(n8447), .A2(n5105), .ZN(n8473) );
  INV_X1 U5004 ( .A(n5525), .ZN(n5558) );
  NOR2_X1 U5005 ( .A1(n8565), .A2(n8566), .ZN(n8577) );
  OR2_X1 U5006 ( .A1(n5523), .A2(n5522), .ZN(n8379) );
  NAND2_X1 U5007 ( .A1(n4655), .A2(n8230), .ZN(n4654) );
  NAND2_X1 U5008 ( .A1(n8066), .A2(n4656), .ZN(n4655) );
  OR2_X1 U5009 ( .A1(n8378), .A2(n8649), .ZN(n8375) );
  AOI21_X1 U5010 ( .B1(n4462), .B2(n4464), .A(n4365), .ZN(n4461) );
  AOI21_X1 U5011 ( .B1(n4823), .B2(n8371), .A(n4359), .ZN(n4822) );
  NAND2_X1 U5012 ( .A1(n8364), .A2(n8363), .ZN(n8729) );
  NAND2_X1 U5013 ( .A1(n4807), .A2(n4472), .ZN(n7534) );
  AOI21_X1 U5014 ( .B1(n4808), .B2(n8260), .A(n4388), .ZN(n4807) );
  NAND2_X1 U5015 ( .A1(n7413), .A2(n4808), .ZN(n4472) );
  NAND2_X1 U5016 ( .A1(n4812), .A2(n4811), .ZN(n4810) );
  INV_X1 U5017 ( .A(n7413), .ZN(n4812) );
  NAND2_X1 U5018 ( .A1(n5497), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4973) );
  INV_X1 U5019 ( .A(n4427), .ZN(n4878) );
  NAND2_X1 U5020 ( .A1(n4883), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4879) );
  NAND2_X1 U5021 ( .A1(n4427), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4881) );
  OR2_X1 U5022 ( .A1(n5280), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n5282) );
  NAND2_X1 U5023 ( .A1(n5113), .A2(n4870), .ZN(n5487) );
  NAND2_X1 U5024 ( .A1(n5648), .A2(n5650), .ZN(n5651) );
  NAND2_X1 U5025 ( .A1(n8038), .A2(n8041), .ZN(n4745) );
  AND2_X1 U5026 ( .A1(n4474), .A2(n4380), .ZN(n9011) );
  NAND2_X1 U5027 ( .A1(n4342), .A2(n4333), .ZN(n4731) );
  OR2_X1 U5028 ( .A1(n6143), .A2(n9059), .ZN(n6162) );
  NAND2_X1 U5029 ( .A1(n4741), .A2(n4740), .ZN(n5627) );
  AOI21_X1 U5030 ( .B1(n4742), .B2(n5586), .A(n5586), .ZN(n4740) );
  AOI21_X1 U5031 ( .B1(P1_IR_REG_19__SCAN_IN), .B2(P1_IR_REG_31__SCAN_IN), .A(
        P1_IR_REG_20__SCAN_IN), .ZN(n4742) );
  NAND2_X1 U5032 ( .A1(n4438), .A2(n4398), .ZN(n4704) );
  INV_X1 U5033 ( .A(n6486), .ZN(n4438) );
  OR2_X1 U5034 ( .A1(n5674), .A2(n5653), .ZN(n5656) );
  AND2_X1 U5035 ( .A1(n6583), .A2(n6524), .ZN(n9169) );
  NAND2_X1 U5036 ( .A1(n9200), .A2(n9191), .ZN(n9186) );
  INV_X1 U5037 ( .A(n4785), .ZN(n9199) );
  OAI21_X1 U5038 ( .B1(n9213), .B2(n4787), .A(n4786), .ZN(n4785) );
  AND2_X1 U5039 ( .A1(n9357), .A2(n9233), .ZN(n4787) );
  NAND2_X1 U5040 ( .A1(n9019), .A2(n6349), .ZN(n4786) );
  INV_X1 U5041 ( .A(n4780), .ZN(n4774) );
  INV_X1 U5042 ( .A(n6282), .ZN(n4778) );
  OAI22_X1 U5043 ( .A1(n6277), .A2(n4789), .B1(n8991), .B2(n9747), .ZN(n7975)
         );
  NOR2_X1 U5044 ( .A1(n8048), .A2(n9073), .ZN(n4789) );
  AOI21_X1 U5045 ( .B1(n4755), .B2(n4753), .A(n4363), .ZN(n4752) );
  INV_X1 U5046 ( .A(n4758), .ZN(n4753) );
  OR2_X1 U5047 ( .A1(n6478), .A2(n6639), .ZN(n9659) );
  AND2_X1 U5048 ( .A1(n4790), .A2(n4616), .ZN(n4615) );
  INV_X1 U5049 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4616) );
  XNOR2_X1 U5050 ( .A(n4445), .B(n4982), .ZN(n7037) );
  NAND2_X1 U5051 ( .A1(n4446), .A2(n4958), .ZN(n4445) );
  NAND2_X1 U5052 ( .A1(n4531), .A2(n4524), .ZN(n4446) );
  INV_X1 U5053 ( .A(n4529), .ZN(n4524) );
  AOI21_X1 U5054 ( .B1(n5517), .B2(n8474), .A(n4335), .ZN(n4420) );
  NAND2_X1 U5055 ( .A1(n8084), .A2(n8083), .ZN(n9676) );
  INV_X1 U5056 ( .A(n9222), .ZN(n9272) );
  NAND2_X1 U5057 ( .A1(n6411), .A2(n6532), .ZN(n4435) );
  NAND2_X1 U5058 ( .A1(n4566), .A2(n4562), .ZN(n8204) );
  OAI21_X1 U5059 ( .B1(n4564), .B2(n4563), .A(n8245), .ZN(n4562) );
  NAND2_X1 U5060 ( .A1(n8275), .A2(n8366), .ZN(n4567) );
  NAND2_X1 U5061 ( .A1(n4432), .A2(n6418), .ZN(n6419) );
  NAND2_X1 U5062 ( .A1(n6417), .A2(n4433), .ZN(n4432) );
  OAI21_X1 U5063 ( .B1(n8217), .B2(n8245), .A(n8225), .ZN(n4586) );
  INV_X1 U5064 ( .A(n9013), .ZN(n4735) );
  NAND2_X1 U5065 ( .A1(n4710), .A2(n4709), .ZN(n6477) );
  NAND2_X1 U5066 ( .A1(n6442), .A2(n4711), .ZN(n4709) );
  AND2_X1 U5067 ( .A1(n6440), .A2(n6439), .ZN(n6476) );
  INV_X1 U5068 ( .A(n6281), .ZN(n4454) );
  OAI21_X1 U5069 ( .B1(n6667), .B2(n4905), .A(n4904), .ZN(n4907) );
  INV_X1 U5070 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4884) );
  NOR2_X1 U5071 ( .A1(n4673), .A2(n4672), .ZN(n4671) );
  INV_X1 U5072 ( .A(n4395), .ZN(n4672) );
  NAND2_X1 U5073 ( .A1(n4515), .A2(n8031), .ZN(n4673) );
  INV_X1 U5074 ( .A(n8425), .ZN(n4515) );
  NAND2_X1 U5075 ( .A1(n4575), .A2(n4573), .ZN(n8241) );
  AOI21_X1 U5076 ( .B1(n4576), .B2(n4578), .A(n4574), .ZN(n4573) );
  INV_X1 U5077 ( .A(n8238), .ZN(n4574) );
  NOR2_X1 U5078 ( .A1(n8627), .A2(n4658), .ZN(n4657) );
  INV_X1 U5079 ( .A(n8220), .ZN(n4658) );
  NAND2_X1 U5080 ( .A1(n4490), .A2(n8061), .ZN(n4489) );
  INV_X1 U5081 ( .A(n4492), .ZN(n4490) );
  NAND2_X1 U5082 ( .A1(n8740), .A2(n4492), .ZN(n8706) );
  NOR2_X1 U5083 ( .A1(n8892), .A2(n8886), .ZN(n4552) );
  OR2_X1 U5084 ( .A1(n8886), .A2(n8428), .ZN(n8366) );
  INV_X1 U5085 ( .A(n8099), .ZN(n4496) );
  AND2_X1 U5086 ( .A1(n8191), .A2(n8099), .ZN(n8189) );
  INV_X1 U5087 ( .A(n4819), .ZN(n4817) );
  NAND2_X1 U5088 ( .A1(n7724), .A2(n4339), .ZN(n4818) );
  INV_X1 U5089 ( .A(n4652), .ZN(n4651) );
  OAI21_X1 U5090 ( .B1(n8263), .B2(n4653), .A(n8145), .ZN(n4652) );
  INV_X1 U5091 ( .A(n8160), .ZN(n4653) );
  INV_X1 U5092 ( .A(n7329), .ZN(n7327) );
  INV_X1 U5093 ( .A(n7088), .ZN(n4794) );
  OR2_X1 U5094 ( .A1(n4498), .A2(n4350), .ZN(n8784) );
  NOR2_X1 U5095 ( .A1(n7416), .A2(n8419), .ZN(n7541) );
  AND2_X1 U5096 ( .A1(n4871), .A2(n4691), .ZN(n4690) );
  NOR2_X1 U5097 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4691) );
  INV_X1 U5098 ( .A(n4476), .ZN(n4475) );
  OAI21_X1 U5099 ( .B1(n4326), .B2(n4340), .A(n7834), .ZN(n4476) );
  AND2_X1 U5100 ( .A1(n4726), .A2(n4479), .ZN(n4478) );
  OR2_X1 U5101 ( .A1(n4480), .A2(n8989), .ZN(n4479) );
  INV_X1 U5102 ( .A(n9001), .ZN(n4480) );
  NAND2_X1 U5103 ( .A1(n7990), .A2(n7992), .ZN(n5945) );
  NAND2_X1 U5104 ( .A1(n9793), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6713) );
  AND2_X1 U5105 ( .A1(n6525), .A2(n6526), .ZN(n4599) );
  OR2_X1 U5106 ( .A1(n9363), .A2(n9038), .ZN(n6577) );
  OR2_X1 U5107 ( .A1(n9372), .A2(n9035), .ZN(n6416) );
  AND2_X1 U5108 ( .A1(n7980), .A2(n6400), .ZN(n6569) );
  NAND2_X1 U5109 ( .A1(n6275), .A2(n4450), .ZN(n4449) );
  INV_X1 U5110 ( .A(n6273), .ZN(n4450) );
  AND2_X1 U5111 ( .A1(n4752), .A2(n4369), .ZN(n4748) );
  NOR2_X1 U5112 ( .A1(n6258), .A2(n7011), .ZN(n7173) );
  NOR2_X1 U5113 ( .A1(n9246), .A2(n9363), .ZN(n9237) );
  INV_X1 U5114 ( .A(n6603), .ZN(n4608) );
  INV_X1 U5115 ( .A(n7274), .ZN(n6266) );
  OR2_X1 U5116 ( .A1(n6334), .A2(n6333), .ZN(n7150) );
  AND2_X1 U5117 ( .A1(n4378), .A2(n5580), .ZN(n4790) );
  INV_X1 U5118 ( .A(n5583), .ZN(n4791) );
  NAND2_X1 U5119 ( .A1(n5547), .A2(n5546), .ZN(n6290) );
  AOI21_X1 U5120 ( .B1(n4719), .B2(n4721), .A(n4718), .ZN(n4717) );
  INV_X1 U5121 ( .A(n5440), .ZN(n4718) );
  INV_X1 U5122 ( .A(n5423), .ZN(n4721) );
  AND2_X1 U5123 ( .A1(n5408), .A2(n5392), .ZN(n5406) );
  AOI21_X1 U5124 ( .B1(n4695), .B2(n4697), .A(n4693), .ZN(n4692) );
  AND2_X1 U5125 ( .A1(n5354), .A2(n5329), .ZN(n5352) );
  AND2_X1 U5126 ( .A1(n5948), .A2(n5597), .ZN(n5972) );
  NAND2_X1 U5127 ( .A1(n4523), .A2(n4525), .ZN(n4712) );
  AOI21_X1 U5128 ( .B1(n4529), .B2(n4958), .A(n4526), .ZN(n4525) );
  INV_X1 U5129 ( .A(n4982), .ZN(n4526) );
  NOR2_X1 U5130 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5948) );
  NAND2_X1 U5131 ( .A1(n4722), .A2(n4527), .ZN(n4531) );
  NAND2_X1 U5132 ( .A1(n5212), .A2(n5211), .ZN(n4722) );
  NAND2_X1 U5133 ( .A1(n4511), .A2(n4513), .ZN(n4510) );
  AND2_X1 U5134 ( .A1(n4932), .A2(n4931), .ZN(n5164) );
  NAND2_X1 U5135 ( .A1(n4506), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4505) );
  INV_X1 U5136 ( .A(n5642), .ZN(n4506) );
  INV_X1 U5137 ( .A(n8518), .ZN(n7239) );
  INV_X1 U5138 ( .A(n5516), .ZN(n4519) );
  NAND2_X1 U5139 ( .A1(n5342), .A2(n5343), .ZN(n4679) );
  NAND2_X1 U5140 ( .A1(n4424), .A2(n5052), .ZN(n5053) );
  INV_X1 U5141 ( .A(n7700), .ZN(n4424) );
  NAND2_X1 U5142 ( .A1(n5210), .A2(n5209), .ZN(n7498) );
  INV_X1 U5143 ( .A(n7363), .ZN(n5210) );
  INV_X1 U5144 ( .A(n4682), .ZN(n4521) );
  OR2_X1 U5145 ( .A1(n8434), .A2(n8435), .ZN(n4682) );
  NOR2_X1 U5146 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4541) );
  XNOR2_X1 U5147 ( .A(n6848), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n6837) );
  NOR2_X1 U5148 ( .A1(n6870), .A2(n6869), .ZN(n6868) );
  OR2_X1 U5149 ( .A1(n6868), .A2(n4535), .ZN(n4534) );
  AND2_X1 U5150 ( .A1(n6858), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4535) );
  AND2_X1 U5151 ( .A1(n4534), .A2(n4533), .ZN(n6897) );
  INV_X1 U5152 ( .A(n6850), .ZN(n4533) );
  NOR2_X1 U5153 ( .A1(n8577), .A2(n4399), .ZN(n8590) );
  INV_X1 U5154 ( .A(n4804), .ZN(n4798) );
  NAND2_X1 U5155 ( .A1(n8376), .A2(n4802), .ZN(n4801) );
  NAND2_X1 U5156 ( .A1(n4804), .A2(n8066), .ZN(n4802) );
  NAND2_X1 U5157 ( .A1(n8629), .A2(n8229), .ZN(n8620) );
  NAND2_X1 U5158 ( .A1(n4499), .A2(n4360), .ZN(n8648) );
  INV_X1 U5159 ( .A(n4463), .ZN(n4462) );
  OAI21_X1 U5160 ( .B1(n8671), .B2(n4464), .A(n8645), .ZN(n4463) );
  INV_X1 U5161 ( .A(n8374), .ZN(n4464) );
  NAND2_X1 U5162 ( .A1(n8664), .A2(n8671), .ZN(n8663) );
  NAND2_X1 U5163 ( .A1(n4821), .A2(n4330), .ZN(n8678) );
  NOR2_X1 U5164 ( .A1(n8716), .A2(n8869), .ZN(n8701) );
  OR2_X1 U5165 ( .A1(n8874), .A2(n8742), .ZN(n4824) );
  AND2_X1 U5166 ( .A1(n8707), .A2(n4824), .ZN(n4823) );
  OAI21_X1 U5167 ( .B1(n8056), .B2(n4493), .A(n4494), .ZN(n8769) );
  AOI21_X1 U5168 ( .B1(n8057), .B2(n4350), .A(n4495), .ZN(n4494) );
  NAND2_X1 U5169 ( .A1(n8057), .A2(n8191), .ZN(n4493) );
  INV_X1 U5170 ( .A(n8198), .ZN(n4495) );
  AOI21_X1 U5171 ( .B1(n4467), .B2(n4469), .A(n4389), .ZN(n4466) );
  NOR2_X2 U5172 ( .A1(n8896), .A2(n8810), .ZN(n8779) );
  NAND2_X1 U5173 ( .A1(n8359), .A2(n4338), .ZN(n8799) );
  INV_X1 U5174 ( .A(n8189), .ZN(n8274) );
  INV_X1 U5175 ( .A(n7893), .ZN(n7894) );
  AND2_X1 U5176 ( .A1(n8174), .A2(n8173), .ZN(n8270) );
  NAND2_X1 U5177 ( .A1(n4327), .A2(n7598), .ZN(n7724) );
  AND2_X1 U5178 ( .A1(n8143), .A2(n8160), .ZN(n8263) );
  NAND2_X1 U5179 ( .A1(n7536), .A2(n8263), .ZN(n7594) );
  NOR2_X1 U5180 ( .A1(n8261), .A2(n4809), .ZN(n4808) );
  INV_X1 U5181 ( .A(n4813), .ZN(n4809) );
  OR2_X1 U5182 ( .A1(n7626), .A2(n8515), .ZN(n4813) );
  NAND2_X1 U5183 ( .A1(n4347), .A2(n7323), .ZN(n7413) );
  NAND2_X1 U5184 ( .A1(n7094), .A2(n8259), .ZN(n7326) );
  NAND2_X1 U5185 ( .A1(n7045), .A2(n8257), .ZN(n7089) );
  NAND2_X1 U5186 ( .A1(n7702), .A2(n7468), .ZN(n7092) );
  AND2_X1 U5187 ( .A1(n8285), .A2(n8089), .ZN(n8803) );
  NAND2_X1 U5188 ( .A1(n7039), .A2(n10003), .ZN(n4806) );
  INV_X1 U5189 ( .A(n7059), .ZN(n7049) );
  NAND2_X1 U5190 ( .A1(n7337), .A2(n7336), .ZN(n7342) );
  OR2_X1 U5191 ( .A1(n10064), .A2(n8815), .ZN(n7023) );
  AND2_X1 U5192 ( .A1(n6831), .A2(n5534), .ZN(n8790) );
  INV_X1 U5193 ( .A(n8803), .ZN(n8793) );
  OR2_X1 U5194 ( .A1(n10029), .A2(n5504), .ZN(n7073) );
  OR2_X1 U5195 ( .A1(n5510), .A2(n5519), .ZN(n10064) );
  INV_X1 U5196 ( .A(n10062), .ZN(n9677) );
  AND2_X1 U5197 ( .A1(n4826), .A2(n4871), .ZN(n4500) );
  AND2_X1 U5198 ( .A1(n4828), .A2(n4827), .ZN(n4826) );
  INV_X1 U5199 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4827) );
  AND2_X1 U5200 ( .A1(n4828), .A2(n4847), .ZN(n4589) );
  INV_X1 U5201 ( .A(n4974), .ZN(n4976) );
  AND2_X1 U5202 ( .A1(n4871), .A2(n4850), .ZN(n4689) );
  NAND2_X1 U5203 ( .A1(n5492), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5509) );
  INV_X1 U5204 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5508) );
  INV_X1 U5205 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n4880) );
  INV_X1 U5206 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n4872) );
  OAI22_X1 U5207 ( .A1(n7143), .A2(n6117), .B1(n9941), .B2(n6118), .ZN(n5634)
         );
  OR2_X1 U5208 ( .A1(n6055), .A2(n8971), .ZN(n6074) );
  NAND2_X1 U5209 ( .A1(n4390), .A2(n4745), .ZN(n8986) );
  NOR2_X1 U5210 ( .A1(n5647), .A2(n4355), .ZN(n6814) );
  NAND2_X1 U5211 ( .A1(n5646), .A2(n5645), .ZN(n5647) );
  NAND2_X1 U5212 ( .A1(n4725), .A2(n4723), .ZN(n9021) );
  AND2_X1 U5213 ( .A1(n4724), .A2(n8962), .ZN(n4723) );
  NAND2_X1 U5214 ( .A1(n4481), .A2(n4478), .ZN(n4725) );
  NAND2_X1 U5215 ( .A1(n4726), .A2(n4728), .ZN(n4724) );
  INV_X1 U5216 ( .A(n6098), .ZN(n6099) );
  OR2_X1 U5217 ( .A1(n5827), .A2(n7561), .ZN(n5845) );
  AND2_X1 U5218 ( .A1(n4481), .A2(n4479), .ZN(n8999) );
  OR2_X1 U5219 ( .A1(n9671), .A2(n9149), .ZN(n6633) );
  AND3_X1 U5220 ( .A1(n6011), .A2(n6010), .A3(n6009), .ZN(n6280) );
  AND4_X1 U5221 ( .A1(n5873), .A2(n5872), .A3(n5871), .A4(n5870), .ZN(n9729)
         );
  INV_X1 U5222 ( .A(n5674), .ZN(n6021) );
  NAND2_X1 U5223 ( .A1(n4402), .A2(n6713), .ZN(n9790) );
  OR2_X1 U5224 ( .A1(n9793), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4402) );
  NAND2_X1 U5225 ( .A1(n4401), .A2(n4400), .ZN(n6712) );
  NOR2_X1 U5226 ( .A1(n6724), .A2(n9786), .ZN(n4400) );
  INV_X1 U5227 ( .A(n9790), .ZN(n4401) );
  NAND2_X1 U5228 ( .A1(n9813), .A2(n9812), .ZN(n9817) );
  NAND2_X1 U5229 ( .A1(n6794), .A2(n4628), .ZN(n4627) );
  INV_X1 U5230 ( .A(n6753), .ZN(n4628) );
  INV_X1 U5231 ( .A(n4627), .ZN(n4626) );
  OR2_X1 U5232 ( .A1(n9862), .A2(n9861), .ZN(n4623) );
  NOR2_X1 U5233 ( .A1(n7738), .A2(n7739), .ZN(n9099) );
  OR2_X1 U5234 ( .A1(n9104), .A2(n9103), .ZN(n4618) );
  OR2_X1 U5235 ( .A1(n9110), .A2(n9109), .ZN(n4408) );
  INV_X1 U5236 ( .A(n6241), .ZN(n6727) );
  NOR2_X2 U5237 ( .A1(n9160), .A2(n6443), .ZN(n9154) );
  AND2_X1 U5238 ( .A1(n9336), .A2(n9180), .ZN(n6288) );
  AND2_X1 U5239 ( .A1(n9167), .A2(n9166), .ZN(n9170) );
  INV_X1 U5240 ( .A(n4599), .ZN(n4598) );
  INV_X1 U5241 ( .A(n6521), .ZN(n4595) );
  NAND2_X1 U5242 ( .A1(n9214), .A2(n4593), .ZN(n4592) );
  NOR2_X1 U5243 ( .A1(n6521), .A2(n4597), .ZN(n4593) );
  NAND2_X1 U5244 ( .A1(n9237), .A2(n9019), .ZN(n9219) );
  NAND2_X1 U5245 ( .A1(n4788), .A2(n4361), .ZN(n9213) );
  NAND2_X1 U5246 ( .A1(n9229), .A2(n6287), .ZN(n4788) );
  OAI21_X1 U5247 ( .B1(n9283), .B2(n6491), .A(n6490), .ZN(n9262) );
  AOI21_X1 U5248 ( .B1(n4773), .B2(n4777), .A(n4332), .ZN(n4771) );
  OR2_X1 U5249 ( .A1(n6492), .A2(n6491), .ZN(n9284) );
  NAND2_X1 U5250 ( .A1(n9305), .A2(n6281), .ZN(n6283) );
  NAND2_X1 U5251 ( .A1(n8017), .A2(n6279), .ZN(n9305) );
  NOR2_X1 U5252 ( .A1(n4637), .A2(n4638), .ZN(n4636) );
  NAND2_X1 U5253 ( .A1(n7858), .A2(n7929), .ZN(n4637) );
  AND2_X1 U5254 ( .A1(n6272), .A2(n4758), .ZN(n4756) );
  INV_X1 U5255 ( .A(n7610), .ZN(n4757) );
  AND2_X1 U5256 ( .A1(n9910), .A2(n6374), .ZN(n7442) );
  NAND2_X1 U5257 ( .A1(n7374), .A2(n7386), .ZN(n7373) );
  AND2_X1 U5258 ( .A1(n6548), .A2(n6366), .ZN(n7274) );
  INV_X1 U5259 ( .A(n7210), .ZN(n6264) );
  AND2_X1 U5260 ( .A1(n7272), .A2(n6361), .ZN(n7210) );
  NAND2_X1 U5261 ( .A1(n7141), .A2(n7144), .ZN(n7140) );
  NAND2_X1 U5262 ( .A1(n6555), .A2(n6599), .ZN(n7145) );
  AND4_X1 U5263 ( .A1(n5706), .A2(n5705), .A3(n5704), .A4(n5703), .ZN(n7403)
         );
  AND2_X1 U5264 ( .A1(n7170), .A2(n6260), .ZN(n7004) );
  XNOR2_X1 U5265 ( .A(n5692), .B(n6891), .ZN(n7006) );
  AND2_X1 U5266 ( .A1(n6217), .A2(n7549), .ZN(n7163) );
  AND2_X1 U5267 ( .A1(n6258), .A2(n7235), .ZN(n7171) );
  NAND2_X1 U5268 ( .A1(n6321), .A2(n6320), .ZN(n9919) );
  INV_X1 U5269 ( .A(n9914), .ZN(n9709) );
  NAND2_X1 U5270 ( .A1(n6453), .A2(n6452), .ZN(n9744) );
  AND2_X1 U5271 ( .A1(n5926), .A2(n5925), .ZN(n9747) );
  AND2_X1 U5272 ( .A1(n7157), .A2(n7549), .ZN(n9395) );
  AND2_X2 U5273 ( .A1(n7157), .A2(n4743), .ZN(n9745) );
  OR2_X1 U5274 ( .A1(n6198), .A2(n8015), .ZN(n9430) );
  XNOR2_X1 U5275 ( .A(n6463), .B(n6462), .ZN(n8933) );
  XNOR2_X1 U5276 ( .A(n6290), .B(n6289), .ZN(n8942) );
  XNOR2_X1 U5277 ( .A(n5545), .B(n5544), .ZN(n6158) );
  XNOR2_X1 U5278 ( .A(n5606), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6214) );
  NAND2_X1 U5279 ( .A1(n5610), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5606) );
  AND2_X1 U5280 ( .A1(n4346), .A2(n4781), .ZN(n4590) );
  XNOR2_X1 U5281 ( .A(n6219), .B(n6218), .ZN(n6660) );
  NAND2_X1 U5282 ( .A1(n4324), .A2(n4346), .ZN(n4782) );
  AND2_X1 U5283 ( .A1(n5906), .A2(n5922), .ZN(n7743) );
  NAND2_X1 U5284 ( .A1(n4706), .A2(n4918), .ZN(n5129) );
  XNOR2_X1 U5285 ( .A(n5058), .B(n5059), .ZN(n5707) );
  NAND2_X1 U5286 ( .A1(n5431), .A2(n5430), .ZN(n8860) );
  NOR2_X1 U5287 ( .A1(n8445), .A2(n4423), .ZN(n4422) );
  INV_X1 U5288 ( .A(n5072), .ZN(n4423) );
  NAND2_X1 U5289 ( .A1(n7698), .A2(n5072), .ZN(n8446) );
  NAND2_X1 U5290 ( .A1(n5263), .A2(n5262), .ZN(n8910) );
  NAND2_X1 U5291 ( .A1(n4830), .A2(n8290), .ZN(n8291) );
  NAND2_X1 U5292 ( .A1(n8289), .A2(n8288), .ZN(n8290) );
  INV_X1 U5293 ( .A(n8788), .ZN(n8808) );
  NAND2_X1 U5294 ( .A1(n5532), .A2(n5531), .ZN(n8632) );
  NAND2_X1 U5295 ( .A1(n5472), .A2(n5471), .ZN(n8649) );
  NAND2_X1 U5296 ( .A1(n5455), .A2(n5454), .ZN(n8673) );
  INV_X1 U5297 ( .A(n8815), .ZN(n8657) );
  XNOR2_X1 U5298 ( .A(n8604), .B(n9676), .ZN(n9673) );
  NOR2_X1 U5299 ( .A1(n8609), .A2(n4558), .ZN(n4557) );
  INV_X1 U5300 ( .A(n4559), .ZN(n4558) );
  NAND2_X1 U5301 ( .A1(n5285), .A2(n5284), .ZN(n8901) );
  OR2_X1 U5302 ( .A1(n5006), .A2(n4547), .ZN(n5022) );
  NAND2_X1 U5303 ( .A1(n6017), .A2(n6016), .ZN(n9384) );
  NAND2_X1 U5304 ( .A1(n9056), .A2(n4746), .ZN(n6257) );
  AND2_X1 U5305 ( .A1(n6648), .A2(n4383), .ZN(n4746) );
  NAND2_X1 U5306 ( .A1(n6124), .A2(n6123), .ZN(n9351) );
  NAND2_X1 U5307 ( .A1(n7932), .A2(n5685), .ZN(n6124) );
  NAND2_X1 U5308 ( .A1(n5952), .A2(n5951), .ZN(n9401) );
  AND4_X1 U5309 ( .A1(n5962), .A2(n5961), .A3(n5960), .A4(n5959), .ZN(n9005)
         );
  INV_X1 U5310 ( .A(n9254), .ZN(n9038) );
  NAND2_X1 U5311 ( .A1(n6150), .A2(n6149), .ZN(n9208) );
  INV_X1 U5312 ( .A(n6280), .ZN(n9299) );
  NOR2_X1 U5313 ( .A1(n7487), .A2(n7486), .ZN(n7738) );
  NAND2_X1 U5314 ( .A1(n4412), .A2(n4410), .ZN(n4409) );
  OR2_X1 U5315 ( .A1(n9141), .A2(n9843), .ZN(n4412) );
  INV_X1 U5316 ( .A(n4411), .ZN(n4410) );
  OAI21_X1 U5317 ( .B1(n9143), .B2(n9142), .A(n9114), .ZN(n4411) );
  AND2_X1 U5318 ( .A1(n6728), .A2(n6727), .ZN(n9895) );
  NOR2_X1 U5319 ( .A1(n9899), .A2(n9146), .ZN(n4632) );
  INV_X1 U5320 ( .A(n9744), .ZN(n9155) );
  XNOR2_X1 U5321 ( .A(n9154), .B(n9155), .ZN(n9742) );
  OR2_X1 U5322 ( .A1(n9659), .A2(n7152), .ZN(n9925) );
  NAND2_X1 U5323 ( .A1(n5630), .A2(n5633), .ZN(n9222) );
  NAND2_X1 U5324 ( .A1(n4584), .A2(n4582), .ZN(n8127) );
  NAND2_X1 U5325 ( .A1(n8106), .A2(n8245), .ZN(n4584) );
  INV_X1 U5326 ( .A(n6569), .ZN(n4441) );
  NAND2_X1 U5327 ( .A1(n4442), .A2(n4440), .ZN(n6403) );
  NAND2_X1 U5328 ( .A1(n6544), .A2(n6483), .ZN(n4442) );
  NAND2_X1 U5329 ( .A1(n4441), .A2(n6478), .ZN(n4440) );
  AND2_X1 U5330 ( .A1(n6416), .A2(n6490), .ZN(n4433) );
  NAND2_X1 U5331 ( .A1(n4436), .A2(n4434), .ZN(n6417) );
  NAND2_X1 U5332 ( .A1(n4437), .A2(n6483), .ZN(n4436) );
  NAND2_X1 U5333 ( .A1(n4435), .A2(n6478), .ZN(n4434) );
  NOR2_X1 U5334 ( .A1(n6426), .A2(n4443), .ZN(n6429) );
  NAND2_X1 U5335 ( .A1(n6428), .A2(n4444), .ZN(n4443) );
  NAND2_X1 U5336 ( .A1(n6427), .A2(n6478), .ZN(n4444) );
  INV_X1 U5337 ( .A(n4586), .ZN(n4585) );
  NAND2_X1 U5338 ( .A1(n8279), .A2(n8215), .ZN(n4587) );
  INV_X1 U5339 ( .A(n8231), .ZN(n4581) );
  INV_X1 U5340 ( .A(n8235), .ZN(n4578) );
  AND2_X1 U5341 ( .A1(n8371), .A2(n8095), .ZN(n4492) );
  INV_X1 U5342 ( .A(n8141), .ZN(n4661) );
  INV_X1 U5343 ( .A(n8109), .ZN(n4660) );
  INV_X1 U5344 ( .A(n8259), .ZN(n4486) );
  INV_X1 U5345 ( .A(n8148), .ZN(n4485) );
  INV_X1 U5346 ( .A(n5882), .ZN(n4477) );
  NOR2_X1 U5347 ( .A1(n9430), .A2(n6208), .ZN(n6333) );
  NOR2_X1 U5348 ( .A1(n5441), .A2(n4720), .ZN(n4719) );
  INV_X1 U5349 ( .A(n5425), .ZN(n4720) );
  INV_X1 U5350 ( .A(n5352), .ZN(n4693) );
  NOR2_X1 U5351 ( .A1(n5325), .A2(n4699), .ZN(n4698) );
  INV_X1 U5352 ( .A(n5302), .ZN(n4699) );
  INV_X1 U5353 ( .A(n4924), .ZN(n4513) );
  NAND2_X1 U5354 ( .A1(n8002), .A2(n4537), .ZN(n8536) );
  NAND2_X1 U5355 ( .A1(n7879), .A2(n4538), .ZN(n4537) );
  INV_X1 U5356 ( .A(n8229), .ZN(n4656) );
  NOR2_X1 U5357 ( .A1(n8840), .A2(n8378), .ZN(n4561) );
  INV_X1 U5358 ( .A(n8360), .ZN(n4469) );
  NOR2_X1 U5359 ( .A1(n7729), .A2(n4555), .ZN(n7899) );
  NAND2_X1 U5360 ( .A1(n7845), .A2(n4556), .ZN(n4555) );
  NOR2_X1 U5361 ( .A1(n7504), .A2(n8306), .ZN(n4556) );
  OR2_X1 U5362 ( .A1(n5152), .A2(n5151), .ZN(n5173) );
  OAI21_X1 U5363 ( .B1(n7094), .B2(n4487), .A(n4484), .ZN(n7329) );
  INV_X1 U5364 ( .A(n4659), .ZN(n4487) );
  AOI21_X1 U5365 ( .B1(n4659), .B2(n4486), .A(n4485), .ZN(n4484) );
  NOR2_X1 U5366 ( .A1(n4661), .A2(n4660), .ZN(n4659) );
  NAND2_X1 U5367 ( .A1(n7061), .A2(n8122), .ZN(n7461) );
  INV_X1 U5368 ( .A(n8823), .ZN(n7052) );
  INV_X1 U5369 ( .A(n6768), .ZN(n6831) );
  NAND2_X1 U5370 ( .A1(n4499), .A2(n8217), .ZN(n8646) );
  AND2_X1 U5371 ( .A1(n7425), .A2(n10044), .ZN(n7426) );
  NAND2_X1 U5372 ( .A1(n5506), .A2(n5505), .ZN(n7335) );
  INV_X1 U5373 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n4844) );
  OR2_X1 U5374 ( .A1(n5131), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5147) );
  INV_X1 U5375 ( .A(n8952), .ZN(n4733) );
  NAND2_X1 U5376 ( .A1(n4352), .A2(n6586), .ZN(n4439) );
  AND2_X1 U5377 ( .A1(n4596), .A2(n4375), .ZN(n4594) );
  NAND2_X1 U5378 ( .A1(n4599), .A2(n4597), .ZN(n4596) );
  INV_X1 U5379 ( .A(n6621), .ZN(n4597) );
  AND2_X1 U5380 ( .A1(n9251), .A2(n9265), .ZN(n6489) );
  NAND2_X1 U5381 ( .A1(n4646), .A2(n9314), .ZN(n4645) );
  NOR2_X1 U5382 ( .A1(n9394), .A2(n9401), .ZN(n4646) );
  OR2_X1 U5383 ( .A1(n9401), .A2(n9005), .ZN(n6400) );
  OR2_X1 U5384 ( .A1(n9407), .A2(n8042), .ZN(n6392) );
  NAND2_X1 U5385 ( .A1(n9752), .A2(n4639), .ZN(n4638) );
  INV_X1 U5386 ( .A(n7163), .ZN(n6238) );
  NAND2_X1 U5387 ( .A1(n4603), .A2(n6387), .ZN(n9707) );
  NAND2_X1 U5388 ( .A1(n7860), .A2(n6388), .ZN(n4603) );
  INV_X1 U5389 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5582) );
  AND2_X1 U5390 ( .A1(n5546), .A2(n5464), .ZN(n5544) );
  AND2_X1 U5391 ( .A1(n5459), .A2(n5445), .ZN(n5457) );
  INV_X1 U5392 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5579) );
  INV_X1 U5393 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5578) );
  INV_X1 U5394 ( .A(n5884), .ZN(n4784) );
  AOI21_X1 U5395 ( .B1(n5298), .B2(n4698), .A(n4696), .ZN(n4695) );
  INV_X1 U5396 ( .A(n5324), .ZN(n4696) );
  INV_X1 U5397 ( .A(n4698), .ZN(n4697) );
  NAND2_X1 U5398 ( .A1(n4530), .A2(n4954), .ZN(n4529) );
  INV_X1 U5399 ( .A(n5258), .ZN(n4530) );
  AND2_X1 U5400 ( .A1(n4951), .A2(n4950), .ZN(n5211) );
  NAND2_X1 U5401 ( .A1(n4933), .A2(n4714), .ZN(n4713) );
  NOR2_X1 U5402 ( .A1(n4938), .A2(n4715), .ZN(n4714) );
  INV_X1 U5403 ( .A(n4932), .ZN(n4715) );
  NAND2_X1 U5404 ( .A1(n4923), .A2(n4918), .ZN(n4514) );
  OR2_X1 U5405 ( .A1(n5758), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5781) );
  INV_X1 U5406 ( .A(n4908), .ZN(n4431) );
  NAND2_X1 U5407 ( .A1(n6667), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n4898) );
  NAND2_X1 U5408 ( .A1(n9656), .A2(n4885), .ZN(n4886) );
  INV_X1 U5409 ( .A(SI_9_), .ZN(n9520) );
  INV_X1 U5410 ( .A(SI_14_), .ZN(n9600) );
  INV_X1 U5411 ( .A(SI_13_), .ZN(n9562) );
  INV_X1 U5412 ( .A(SI_21_), .ZN(n9559) );
  XNOR2_X1 U5413 ( .A(n8177), .B(n5550), .ZN(n5254) );
  OR2_X1 U5414 ( .A1(n5344), .A2(n9564), .ZN(n5374) );
  XNOR2_X1 U5415 ( .A(n8879), .B(n5550), .ZN(n5358) );
  NAND2_X1 U5416 ( .A1(n5277), .A2(n5276), .ZN(n4688) );
  AND2_X1 U5417 ( .A1(n5274), .A2(n4687), .ZN(n4686) );
  OR2_X1 U5418 ( .A1(n5216), .A2(n7803), .ZN(n5246) );
  INV_X1 U5419 ( .A(n4678), .ZN(n4677) );
  NAND2_X1 U5420 ( .A1(n4671), .A2(n4675), .ZN(n4507) );
  NAND2_X1 U5421 ( .A1(n4862), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5311) );
  INV_X1 U5422 ( .A(n5288), .ZN(n4862) );
  INV_X1 U5423 ( .A(n5309), .ZN(n5097) );
  INV_X1 U5424 ( .A(n8649), .ZN(n8497) );
  OAI21_X1 U5425 ( .B1(n4322), .B2(n4321), .A(n8252), .ZN(n4570) );
  NAND2_X1 U5426 ( .A1(n4323), .A2(n8252), .ZN(n4571) );
  NOR2_X1 U5427 ( .A1(n6943), .A2(n4536), .ZN(n6870) );
  AND2_X1 U5428 ( .A1(n6857), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4536) );
  NOR2_X1 U5429 ( .A1(n6928), .A2(n4386), .ZN(n6931) );
  NOR2_X1 U5430 ( .A1(n6931), .A2(n6930), .ZN(n6953) );
  NOR2_X1 U5431 ( .A1(n6953), .A2(n4543), .ZN(n6957) );
  AND2_X1 U5432 ( .A1(n6954), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4543) );
  NOR2_X1 U5433 ( .A1(n6957), .A2(n6956), .ZN(n7121) );
  NOR2_X1 U5434 ( .A1(n7287), .A2(n4545), .ZN(n7290) );
  AND2_X1 U5435 ( .A1(n7293), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4545) );
  NOR2_X1 U5436 ( .A1(n7290), .A2(n7289), .ZN(n7648) );
  NOR2_X1 U5437 ( .A1(n7648), .A2(n4544), .ZN(n7650) );
  AND2_X1 U5438 ( .A1(n7649), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4544) );
  NOR2_X1 U5439 ( .A1(n7650), .A2(n7651), .ZN(n7798) );
  NAND2_X1 U5440 ( .A1(n7873), .A2(n4539), .ZN(n7875) );
  OR2_X1 U5441 ( .A1(n7874), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4539) );
  NAND2_X1 U5442 ( .A1(n7875), .A2(n7876), .ZN(n8002) );
  XNOR2_X1 U5443 ( .A(n8536), .B(n8537), .ZN(n8004) );
  NAND2_X1 U5444 ( .A1(n8563), .A2(n8564), .ZN(n8565) );
  AOI21_X1 U5445 ( .B1(n8590), .B2(n8591), .A(n4532), .ZN(n8592) );
  NOR2_X1 U5446 ( .A1(n8583), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n4532) );
  AND2_X1 U5447 ( .A1(n4560), .A2(n4561), .ZN(n4559) );
  AND2_X1 U5448 ( .A1(n5524), .A2(n8379), .ZN(n8616) );
  OR2_X1 U5449 ( .A1(n8860), .A2(n8681), .ZN(n8666) );
  OAI21_X1 U5450 ( .B1(n8740), .B2(n4491), .A(n4488), .ZN(n8695) );
  INV_X1 U5451 ( .A(n8061), .ZN(n4491) );
  AND2_X1 U5452 ( .A1(n8064), .A2(n4489), .ZN(n4488) );
  AND2_X1 U5453 ( .A1(n5439), .A2(n5438), .ZN(n8693) );
  NOR2_X1 U5454 ( .A1(n8874), .A2(n4550), .ZN(n4548) );
  NAND2_X1 U5455 ( .A1(n8779), .A2(n4552), .ZN(n8752) );
  AND2_X1 U5456 ( .A1(n8366), .A2(n8365), .ZN(n8751) );
  NAND2_X1 U5457 ( .A1(n8769), .A2(n8770), .ZN(n8768) );
  NAND2_X1 U5458 ( .A1(n8779), .A2(n8767), .ZN(n8762) );
  AND2_X1 U5459 ( .A1(n8275), .A2(n8747), .ZN(n8770) );
  OR2_X1 U5460 ( .A1(n8809), .A2(n8901), .ZN(n8810) );
  OR2_X1 U5461 ( .A1(n5286), .A2(n9604), .ZN(n5288) );
  INV_X1 U5462 ( .A(n8506), .ZN(n8807) );
  OR2_X1 U5463 ( .A1(n5264), .A2(n7661), .ZN(n5266) );
  NAND2_X1 U5464 ( .A1(n4861), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5286) );
  INV_X1 U5465 ( .A(n5266), .ZN(n4861) );
  NAND2_X1 U5466 ( .A1(n7949), .A2(n7948), .ZN(n8056) );
  OAI21_X1 U5467 ( .B1(n7906), .B2(n7905), .A(n7904), .ZN(n7907) );
  AND2_X1 U5468 ( .A1(n7899), .A2(n7903), .ZN(n7940) );
  OAI211_X1 U5469 ( .C1(n4815), .C2(n4339), .A(n4470), .B(n7770), .ZN(n7893)
         );
  NOR2_X1 U5470 ( .A1(n7729), .A2(n4554), .ZN(n7776) );
  INV_X1 U5471 ( .A(n4556), .ZN(n4554) );
  NAND2_X1 U5472 ( .A1(n4818), .A2(n4816), .ZN(n7771) );
  NAND2_X1 U5473 ( .A1(n4818), .A2(n4819), .ZN(n7752) );
  AOI21_X1 U5474 ( .B1(n4651), .B2(n4653), .A(n4650), .ZN(n4649) );
  INV_X1 U5475 ( .A(n8152), .ZN(n4650) );
  AND2_X1 U5476 ( .A1(n7541), .A2(n10055), .ZN(n7602) );
  INV_X1 U5477 ( .A(n4793), .ZN(n4792) );
  NOR2_X1 U5478 ( .A1(n7471), .A2(n7704), .ZN(n7425) );
  INV_X1 U5479 ( .A(n8517), .ZN(n7090) );
  NAND2_X1 U5480 ( .A1(n7461), .A2(n8254), .ZN(n7460) );
  OR2_X1 U5481 ( .A1(n7469), .A2(n7468), .ZN(n7471) );
  AND2_X1 U5482 ( .A1(n8113), .A2(n8120), .ZN(n4837) );
  NAND2_X1 U5483 ( .A1(n4837), .A2(n7049), .ZN(n7061) );
  OR2_X1 U5484 ( .A1(n8812), .A2(n8657), .ZN(n7760) );
  NOR2_X1 U5485 ( .A1(n10003), .A2(n7553), .ZN(n7063) );
  NAND2_X1 U5486 ( .A1(n7550), .A2(n7553), .ZN(n7048) );
  NAND2_X1 U5487 ( .A1(n5006), .A2(n4668), .ZN(n4667) );
  NAND2_X1 U5488 ( .A1(n8784), .A2(n8057), .ZN(n8785) );
  AND2_X1 U5489 ( .A1(n8359), .A2(n8358), .ZN(n8800) );
  AND2_X1 U5490 ( .A1(n7023), .A2(n7335), .ZN(n7071) );
  AND2_X1 U5491 ( .A1(n7075), .A2(n7022), .ZN(n7337) );
  OR2_X1 U5492 ( .A1(n5510), .A2(n5536), .ZN(n10062) );
  INV_X1 U5493 ( .A(n10064), .ZN(n9683) );
  XNOR2_X1 U5494 ( .A(n5509), .B(n5508), .ZN(n6765) );
  INV_X1 U5495 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5490) );
  OR3_X1 U5496 ( .A1(n5198), .A2(P2_IR_REG_10__SCAN_IN), .A3(
        P2_IR_REG_11__SCAN_IN), .ZN(n5213) );
  NAND2_X1 U5497 ( .A1(n5775), .A2(n5776), .ZN(n7184) );
  NAND2_X1 U5498 ( .A1(n6102), .A2(n9031), .ZN(n4730) );
  INV_X1 U5499 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6018) );
  AOI21_X1 U5500 ( .B1(n4351), .B2(n9042), .A(n4727), .ZN(n4726) );
  AND2_X1 U5501 ( .A1(n4729), .A2(n9043), .ZN(n4727) );
  NOR2_X1 U5502 ( .A1(n9043), .A2(n9042), .ZN(n4728) );
  NAND2_X1 U5503 ( .A1(n7692), .A2(n7691), .ZN(n4744) );
  NAND2_X1 U5504 ( .A1(n5954), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5981) );
  INV_X1 U5505 ( .A(n7522), .ZN(n4739) );
  NAND2_X1 U5506 ( .A1(n7307), .A2(n7310), .ZN(n4737) );
  INV_X1 U5507 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5888) );
  OR2_X1 U5508 ( .A1(n5889), .A2(n5888), .ZN(n5911) );
  NAND2_X1 U5509 ( .A1(n6001), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6019) );
  INV_X1 U5510 ( .A(n6003), .ZN(n6001) );
  INV_X1 U5511 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5927) );
  OR2_X1 U5512 ( .A1(n5928), .A2(n5927), .ZN(n5956) );
  NAND2_X1 U5513 ( .A1(n5947), .A2(n5946), .ZN(n8039) );
  AND2_X1 U5514 ( .A1(n6062), .A2(n6061), .ZN(n9035) );
  NAND2_X1 U5515 ( .A1(n9817), .A2(n6714), .ZN(n6717) );
  AND2_X1 U5516 ( .A1(n6717), .A2(n6716), .ZN(n6738) );
  NAND2_X1 U5517 ( .A1(n6786), .A2(n4404), .ZN(n6778) );
  OR2_X1 U5518 ( .A1(n6754), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n4404) );
  NAND2_X1 U5519 ( .A1(n6778), .A2(n6779), .ZN(n6777) );
  OR2_X1 U5520 ( .A1(n5781), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5801) );
  NAND2_X1 U5521 ( .A1(n6777), .A2(n4403), .ZN(n6744) );
  OR2_X1 U5522 ( .A1(n6746), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n4403) );
  NOR2_X1 U5523 ( .A1(n6744), .A2(n6743), .ZN(n6967) );
  NAND2_X1 U5524 ( .A1(n4623), .A2(n4622), .ZN(n4621) );
  NAND2_X1 U5525 ( .A1(n9866), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4622) );
  NAND2_X1 U5526 ( .A1(n9869), .A2(n4406), .ZN(n9086) );
  OR2_X1 U5527 ( .A1(n9879), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n4406) );
  NOR2_X1 U5528 ( .A1(n9873), .A2(n4619), .ZN(n9093) );
  AND2_X1 U5529 ( .A1(n9879), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4619) );
  NAND2_X1 U5530 ( .A1(n9086), .A2(n9087), .ZN(n9085) );
  NOR2_X1 U5531 ( .A1(n7484), .A2(n4394), .ZN(n7737) );
  AND2_X1 U5532 ( .A1(n4408), .A2(n4407), .ZN(n9120) );
  NAND2_X1 U5533 ( .A1(n9124), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n4407) );
  NOR2_X1 U5534 ( .A1(n9120), .A2(n9119), .ZN(n9137) );
  AND2_X1 U5535 ( .A1(n4618), .A2(n4617), .ZN(n9127) );
  NAND2_X1 U5536 ( .A1(n9124), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4617) );
  NOR2_X1 U5537 ( .A1(n9127), .A2(n9126), .ZN(n9132) );
  AND2_X1 U5538 ( .A1(n6230), .A2(n6182), .ZN(n9163) );
  NAND2_X1 U5539 ( .A1(n4766), .A2(n9063), .ZN(n4765) );
  NAND2_X1 U5540 ( .A1(n4768), .A2(n4767), .ZN(n4458) );
  NOR2_X1 U5541 ( .A1(n9169), .A2(n4763), .ZN(n4762) );
  INV_X1 U5542 ( .A(n4765), .ZN(n4763) );
  AND2_X1 U5543 ( .A1(n6430), .A2(n9205), .ZN(n6621) );
  OR2_X1 U5544 ( .A1(n6513), .A2(n6512), .ZN(n9192) );
  AND2_X1 U5545 ( .A1(n6525), .A2(n6430), .ZN(n9206) );
  NOR2_X1 U5546 ( .A1(n4453), .A2(n4452), .ZN(n9245) );
  NAND2_X1 U5547 ( .A1(n4353), .A2(n4769), .ZN(n4452) );
  NOR2_X1 U5548 ( .A1(n8017), .A2(n4364), .ZN(n4453) );
  AND2_X1 U5549 ( .A1(n6409), .A2(n6528), .ZN(n9296) );
  NAND2_X1 U5550 ( .A1(n6313), .A2(n4331), .ZN(n9316) );
  NOR2_X1 U5551 ( .A1(n7976), .A2(n4644), .ZN(n9307) );
  INV_X1 U5552 ( .A(n4646), .ZN(n4644) );
  NOR2_X1 U5553 ( .A1(n7976), .A2(n9401), .ZN(n8019) );
  AOI21_X1 U5554 ( .B1(n4325), .B2(n4451), .A(n4362), .ZN(n4448) );
  INV_X1 U5555 ( .A(n6275), .ZN(n4451) );
  NAND2_X1 U5556 ( .A1(n6540), .A2(n6387), .ZN(n4602) );
  NAND2_X1 U5557 ( .A1(n4600), .A2(n6540), .ZN(n4601) );
  NOR3_X1 U5558 ( .A1(n9721), .A2(n9411), .A3(n4638), .ZN(n9701) );
  NOR3_X1 U5559 ( .A1(n9721), .A2(n9411), .A3(n9759), .ZN(n9699) );
  AOI21_X1 U5560 ( .B1(n4748), .B2(n4754), .A(n4329), .ZN(n4749) );
  NOR2_X1 U5561 ( .A1(n9721), .A2(n9759), .ZN(n9722) );
  NAND2_X1 U5562 ( .A1(n4759), .A2(n7315), .ZN(n4758) );
  NAND2_X1 U5563 ( .A1(n6557), .A2(n6377), .ZN(n7610) );
  AND4_X1 U5564 ( .A1(n5791), .A2(n5790), .A3(n5789), .A4(n5788), .ZN(n9917)
         );
  NAND2_X1 U5565 ( .A1(n6267), .A2(n6266), .ZN(n7271) );
  AND4_X1 U5566 ( .A1(n5742), .A2(n5741), .A3(n5740), .A4(n5739), .ZN(n7388)
         );
  NAND2_X1 U5567 ( .A1(n6602), .A2(n6599), .ZN(n7401) );
  OR2_X1 U5568 ( .A1(n6659), .A2(n6727), .ZN(n9914) );
  NAND2_X1 U5569 ( .A1(n4317), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5686) );
  NAND2_X1 U5570 ( .A1(n5685), .A2(n5684), .ZN(n5687) );
  NAND2_X1 U5571 ( .A1(n7171), .A2(n7175), .ZN(n7170) );
  OR2_X1 U5572 ( .A1(n6299), .A2(n6238), .ZN(n7168) );
  NAND2_X1 U5573 ( .A1(n6297), .A2(n6296), .ZN(n6443) );
  NAND2_X1 U5574 ( .A1(n6142), .A2(n6141), .ZN(n9346) );
  NOR2_X1 U5575 ( .A1(n7150), .A2(n6335), .ZN(n6339) );
  NAND2_X1 U5576 ( .A1(n5581), .A2(n4790), .ZN(n5615) );
  NAND2_X1 U5577 ( .A1(n5604), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5607) );
  NAND2_X1 U5578 ( .A1(n5607), .A2(n5605), .ZN(n5610) );
  XNOR2_X1 U5579 ( .A(n5442), .B(n5441), .ZN(n7932) );
  AND2_X1 U5580 ( .A1(n5972), .A2(n5598), .ZN(n5599) );
  NOR2_X1 U5581 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5598) );
  NAND2_X1 U5582 ( .A1(n4700), .A2(n5302), .ZN(n5326) );
  NAND2_X1 U5583 ( .A1(n4712), .A2(n4963), .ZN(n5279) );
  NAND2_X1 U5584 ( .A1(n4531), .A2(n4954), .ZN(n5259) );
  XNOR2_X1 U5585 ( .A(n5236), .B(n5235), .ZN(n6818) );
  NAND2_X1 U5586 ( .A1(n4722), .A2(n4951), .ZN(n5236) );
  AND3_X1 U5587 ( .A1(n5575), .A2(n4783), .A3(n5574), .ZN(n5884) );
  XNOR2_X1 U5588 ( .A(n5182), .B(n5181), .ZN(n6706) );
  INV_X1 U5589 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5803) );
  NAND2_X1 U5590 ( .A1(n4909), .A2(n4908), .ZN(n5073) );
  XNOR2_X1 U5591 ( .A(n4895), .B(n4894), .ZN(n5017) );
  OR2_X1 U5592 ( .A1(n7361), .A2(n5179), .ZN(n5180) );
  AOI21_X1 U5593 ( .B1(n4520), .B2(n4683), .A(n4519), .ZN(n4518) );
  NAND2_X1 U5594 ( .A1(n6691), .A2(n4983), .ZN(n4473) );
  INV_X1 U5595 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9564) );
  XNOR2_X1 U5596 ( .A(n5358), .B(n4516), .ZN(n8425) );
  INV_X1 U5597 ( .A(n5359), .ZN(n4516) );
  AOI21_X1 U5598 ( .B1(n8032), .B2(n8031), .A(n4676), .ZN(n8426) );
  INV_X1 U5599 ( .A(n4679), .ZN(n4676) );
  NAND2_X1 U5600 ( .A1(n4987), .A2(n4986), .ZN(n8905) );
  AND2_X1 U5601 ( .A1(n7884), .A2(n4688), .ZN(n4684) );
  AND2_X1 U5602 ( .A1(n4685), .A2(n4688), .ZN(n7885) );
  NAND2_X1 U5603 ( .A1(n5411), .A2(n5410), .ZN(n8864) );
  NAND2_X1 U5604 ( .A1(n5068), .A2(n7247), .ZN(n7698) );
  AND4_X1 U5605 ( .A1(n5048), .A2(n4662), .A3(n5049), .A4(n5050), .ZN(n7702)
         );
  NAND2_X1 U5606 ( .A1(n5025), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4662) );
  INV_X1 U5607 ( .A(n8464), .ZN(n8495) );
  INV_X1 U5608 ( .A(n8465), .ZN(n8496) );
  XNOR2_X1 U5609 ( .A(n5342), .B(n5341), .ZN(n8031) );
  AND2_X1 U5610 ( .A1(n4674), .A2(n4395), .ZN(n8032) );
  OR2_X1 U5611 ( .A1(n8356), .A2(n4675), .ZN(n4674) );
  NAND2_X1 U5612 ( .A1(n5331), .A2(n5330), .ZN(n8886) );
  AND2_X1 U5613 ( .A1(n7516), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8479) );
  OR2_X1 U5614 ( .A1(n8490), .A2(n5514), .ZN(n8415) );
  AND2_X1 U5615 ( .A1(n8477), .A2(n8788), .ZN(n8464) );
  INV_X1 U5616 ( .A(n8468), .ZN(n5035) );
  NAND2_X1 U5617 ( .A1(n4981), .A2(n4980), .ZN(n8896) );
  INV_X1 U5618 ( .A(n7507), .ZN(n8500) );
  NAND2_X1 U5619 ( .A1(n4522), .A2(n4682), .ZN(n8489) );
  OAI21_X1 U5620 ( .B1(n5520), .B2(n7341), .A(n10025), .ZN(n8461) );
  NAND2_X1 U5621 ( .A1(n8090), .A2(n8089), .ZN(n8292) );
  NAND2_X1 U5622 ( .A1(n6833), .A2(n10033), .ZN(n10027) );
  INV_X1 U5623 ( .A(n7024), .ZN(n5511) );
  INV_X1 U5624 ( .A(n7702), .ZN(n8519) );
  INV_X2 U5625 ( .A(P2_U3966), .ZN(n8521) );
  AND2_X1 U5626 ( .A1(n4542), .A2(n4540), .ZN(n6848) );
  NAND2_X1 U5627 ( .A1(n4368), .A2(P2_IR_REG_1__SCAN_IN), .ZN(n4542) );
  NOR2_X1 U5628 ( .A1(n5000), .A2(n4541), .ZN(n4540) );
  INV_X1 U5629 ( .A(n4534), .ZN(n6851) );
  AND2_X1 U5630 ( .A1(n6842), .A2(n5534), .ZN(n8596) );
  INV_X1 U5631 ( .A(n9997), .ZN(n9992) );
  NAND2_X1 U5632 ( .A1(n8619), .A2(n8377), .ZN(n4803) );
  NAND2_X1 U5633 ( .A1(n4801), .A2(n4800), .ZN(n4799) );
  AOI21_X1 U5634 ( .B1(n8389), .B2(n8793), .A(n8388), .ZN(n8838) );
  NAND2_X1 U5635 ( .A1(n8387), .A2(n8386), .ZN(n8388) );
  NAND2_X1 U5636 ( .A1(n8626), .A2(n8375), .ZN(n4471) );
  AND2_X1 U5637 ( .A1(n8624), .A2(n8623), .ZN(n8843) );
  AOI22_X1 U5638 ( .A1(n8649), .A2(n8788), .B1(n8622), .B2(n8790), .ZN(n8623)
         );
  NAND2_X1 U5639 ( .A1(n8621), .A2(n8793), .ZN(n8624) );
  AND2_X1 U5640 ( .A1(n8648), .A2(n8220), .ZN(n8631) );
  OAI21_X1 U5641 ( .B1(n8664), .B2(n4464), .A(n4462), .ZN(n8644) );
  NAND2_X1 U5642 ( .A1(n8663), .A2(n8374), .ZN(n8642) );
  NAND2_X1 U5643 ( .A1(n5447), .A2(n5446), .ZN(n8851) );
  NAND2_X1 U5644 ( .A1(n4821), .A2(n4822), .ZN(n8680) );
  NAND2_X1 U5645 ( .A1(n4825), .A2(n4823), .ZN(n8700) );
  OR2_X1 U5646 ( .A1(n8715), .A2(n8371), .ZN(n4825) );
  NAND2_X1 U5647 ( .A1(n8740), .A2(n8095), .ZN(n8722) );
  NAND2_X1 U5648 ( .A1(n8799), .A2(n8360), .ZN(n8777) );
  AND2_X1 U5649 ( .A1(n7938), .A2(n7937), .ZN(n7939) );
  NAND2_X1 U5650 ( .A1(n7724), .A2(n7723), .ZN(n7750) );
  NAND2_X1 U5651 ( .A1(n7594), .A2(n8160), .ZN(n7679) );
  NAND2_X1 U5652 ( .A1(n4810), .A2(n4808), .ZN(n7530) );
  NAND2_X1 U5653 ( .A1(n4810), .A2(n4813), .ZN(n7324) );
  NAND2_X1 U5654 ( .A1(n7326), .A2(n8109), .ZN(n7419) );
  NAND2_X1 U5655 ( .A1(n7089), .A2(n7088), .ZN(n7424) );
  INV_X1 U5656 ( .A(n10018), .ZN(n8824) );
  NAND2_X1 U5657 ( .A1(n4806), .A2(n7041), .ZN(n7060) );
  INV_X1 U5658 ( .A(n10025), .ZN(n8827) );
  NOR2_X1 U5659 ( .A1(n7342), .A2(n8657), .ZN(n10011) );
  OR2_X1 U5660 ( .A1(n10027), .A2(n7023), .ZN(n10025) );
  NAND2_X1 U5661 ( .A1(n10009), .A2(n10004), .ZN(n10018) );
  INV_X2 U5662 ( .A(n10009), .ZN(n10022) );
  AOI211_X1 U5663 ( .C1(n9677), .C2(n9676), .A(n9675), .B(n9674), .ZN(n9693)
         );
  NAND2_X1 U5664 ( .A1(n7337), .A2(n7071), .ZN(n10070) );
  AND2_X1 U5665 ( .A1(n6765), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10033) );
  OR2_X1 U5666 ( .A1(n10027), .A2(n10026), .ZN(n10030) );
  NOR2_X1 U5667 ( .A1(n4976), .A2(n4975), .ZN(n4977) );
  NOR2_X1 U5668 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4975) );
  NAND2_X1 U5669 ( .A1(n5497), .A2(n5499), .ZN(n8030) );
  NAND2_X1 U5670 ( .A1(n5489), .A2(n4393), .ZN(n7936) );
  XNOR2_X1 U5671 ( .A(n5495), .B(n5494), .ZN(n7915) );
  INV_X1 U5672 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5494) );
  INV_X1 U5673 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4876) );
  INV_X1 U5674 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7511) );
  INV_X1 U5675 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7306) );
  OR2_X1 U5676 ( .A1(n4881), .A2(n4880), .ZN(n4882) );
  AND2_X1 U5677 ( .A1(n5283), .A2(n5282), .ZN(n8578) );
  INV_X1 U5678 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7000) );
  NOR2_X1 U5679 ( .A1(n4968), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8943) );
  INV_X1 U5680 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6708) );
  INV_X1 U5681 ( .A(n6848), .ZN(n6855) );
  NOR2_X1 U5682 ( .A1(n5625), .A2(n6658), .ZN(n9804) );
  NAND2_X1 U5683 ( .A1(n6158), .A2(n4318), .ZN(n4705) );
  NAND2_X1 U5684 ( .A1(n6087), .A2(n6086), .ZN(n9363) );
  OAI21_X1 U5685 ( .B1(n8999), .B2(n4728), .A(n4726), .ZN(n8963) );
  NAND2_X1 U5686 ( .A1(n6178), .A2(n6177), .ZN(n9336) );
  NAND2_X1 U5687 ( .A1(n5672), .A2(n5671), .ZN(n6881) );
  AOI21_X1 U5688 ( .B1(n9021), .B2(n6052), .A(n4344), .ZN(n8970) );
  NAND2_X1 U5689 ( .A1(n4744), .A2(n5858), .ZN(n7823) );
  NAND2_X1 U5690 ( .A1(n4745), .A2(n8039), .ZN(n8988) );
  NAND2_X1 U5691 ( .A1(n8986), .A2(n8989), .ZN(n9000) );
  INV_X1 U5692 ( .A(n9060), .ZN(n9048) );
  AND4_X1 U5693 ( .A1(n5723), .A2(n5722), .A3(n5721), .A4(n5720), .ZN(n7142)
         );
  INV_X1 U5694 ( .A(n6992), .ZN(n4482) );
  NAND2_X1 U5695 ( .A1(n5707), .A2(n5685), .ZN(n4483) );
  AND4_X1 U5696 ( .A1(n5833), .A2(n5832), .A3(n5831), .A4(n5830), .ZN(n9915)
         );
  NAND2_X1 U5697 ( .A1(n4737), .A2(n7308), .ZN(n7521) );
  NAND2_X1 U5698 ( .A1(n6032), .A2(n6031), .ZN(n9379) );
  NAND2_X1 U5699 ( .A1(n7821), .A2(n5882), .ZN(n7837) );
  NAND2_X1 U5700 ( .A1(n6073), .A2(n6072), .ZN(n9366) );
  AND4_X1 U5701 ( .A1(n5595), .A2(n5594), .A3(n5593), .A4(n5592), .ZN(n7143)
         );
  OR2_X1 U5702 ( .A1(n5675), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5594) );
  OR2_X1 U5703 ( .A1(n6242), .A2(n6727), .ZN(n9062) );
  NAND2_X1 U5704 ( .A1(n8999), .A2(n5996), .ZN(n9045) );
  NAND2_X1 U5705 ( .A1(n6000), .A2(n5999), .ZN(n9389) );
  AND2_X1 U5706 ( .A1(n6134), .A2(n6133), .ZN(n9061) );
  AOI21_X1 U5707 ( .B1(n8978), .B2(n8979), .A(n4384), .ZN(n9058) );
  NAND2_X1 U5708 ( .A1(n9058), .A2(n9057), .ZN(n9056) );
  AND2_X1 U5709 ( .A1(n6162), .A2(n6144), .ZN(n9189) );
  INV_X1 U5710 ( .A(n9066), .ZN(n9050) );
  AND2_X1 U5711 ( .A1(n7318), .A2(n9745), .ZN(n9052) );
  NAND2_X1 U5712 ( .A1(n5628), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5629) );
  OAI21_X1 U5713 ( .B1(n6640), .B2(n6639), .A(n6638), .ZN(n6641) );
  AND3_X1 U5714 ( .A1(n6473), .A2(n6472), .A3(n6471), .ZN(n9149) );
  INV_X1 U5715 ( .A(n9061), .ZN(n9217) );
  NAND2_X1 U5716 ( .A1(n6116), .A2(n6115), .ZN(n9233) );
  OR2_X1 U5717 ( .A1(n9224), .A2(n5675), .ZN(n6116) );
  NAND2_X1 U5718 ( .A1(n6093), .A2(n6092), .ZN(n9254) );
  INV_X1 U5719 ( .A(n9035), .ZN(n9285) );
  INV_X1 U5720 ( .A(n7142), .ZN(n9081) );
  OR2_X1 U5721 ( .A1(n5677), .A2(n5676), .ZN(n5679) );
  OR2_X1 U5722 ( .A1(n5675), .A2(n7180), .ZN(n5657) );
  OR2_X1 U5723 ( .A1(n5677), .A2(n5654), .ZN(n5655) );
  OR2_X1 U5724 ( .A1(n5677), .A2(n5635), .ZN(n5641) );
  OR2_X1 U5725 ( .A1(n5675), .A2(n5637), .ZN(n5638) );
  OR2_X1 U5726 ( .A1(n5674), .A2(n9786), .ZN(n5639) );
  INV_X1 U5727 ( .A(n6712), .ZN(n9789) );
  NOR2_X1 U5728 ( .A1(n9851), .A2(n9852), .ZN(n9850) );
  OR2_X1 U5729 ( .A1(n9850), .A2(n4627), .ZN(n6793) );
  NOR2_X1 U5730 ( .A1(n9850), .A2(n6753), .ZN(n6795) );
  AOI21_X1 U5731 ( .B1(n4626), .B2(n9852), .A(n4385), .ZN(n4625) );
  INV_X1 U5732 ( .A(n4623), .ZN(n9860) );
  AND2_X1 U5733 ( .A1(n4621), .A2(n4620), .ZN(n9873) );
  INV_X1 U5734 ( .A(n9874), .ZN(n4620) );
  INV_X1 U5735 ( .A(n4621), .ZN(n9875) );
  NAND2_X1 U5736 ( .A1(n9085), .A2(n4405), .ZN(n6973) );
  OR2_X1 U5737 ( .A1(n6983), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n4405) );
  NAND2_X1 U5738 ( .A1(n6973), .A2(n6972), .ZN(n7104) );
  XNOR2_X1 U5739 ( .A(n7737), .B(n7736), .ZN(n7487) );
  NOR2_X1 U5740 ( .A1(n9100), .A2(n9101), .ZN(n9104) );
  INV_X1 U5741 ( .A(n4618), .ZN(n9123) );
  INV_X1 U5742 ( .A(n9895), .ZN(n9872) );
  NOR2_X1 U5743 ( .A1(n9107), .A2(n9108), .ZN(n9110) );
  INV_X1 U5744 ( .A(n4408), .ZN(n9118) );
  INV_X1 U5745 ( .A(n9145), .ZN(n4631) );
  NAND2_X1 U5746 ( .A1(n6465), .A2(n6464), .ZN(n9671) );
  XNOR2_X1 U5747 ( .A(n6319), .B(n6298), .ZN(n6330) );
  XNOR2_X1 U5748 ( .A(n4764), .B(n6517), .ZN(n8346) );
  OAI21_X1 U5749 ( .B1(n4768), .B2(n4761), .A(n4760), .ZN(n4764) );
  AOI21_X1 U5750 ( .B1(n4762), .B2(n9179), .A(n6288), .ZN(n4760) );
  INV_X1 U5751 ( .A(n4762), .ZN(n4761) );
  NAND2_X1 U5752 ( .A1(n4456), .A2(n4455), .ZN(n9340) );
  NAND2_X1 U5753 ( .A1(n4457), .A2(n9169), .ZN(n4456) );
  NAND2_X1 U5754 ( .A1(n4458), .A2(n4762), .ZN(n4455) );
  NAND2_X1 U5755 ( .A1(n4458), .A2(n4765), .ZN(n4457) );
  AOI21_X1 U5756 ( .B1(n9171), .B2(n9709), .A(n4387), .ZN(n4613) );
  NAND2_X1 U5757 ( .A1(n9172), .A2(n9919), .ZN(n4614) );
  NAND2_X1 U5758 ( .A1(n4592), .A2(n4591), .ZN(n9178) );
  NAND2_X1 U5759 ( .A1(n4598), .A2(n4595), .ZN(n4591) );
  NAND2_X1 U5760 ( .A1(n6104), .A2(n6103), .ZN(n9357) );
  INV_X1 U5761 ( .A(n9366), .ZN(n9251) );
  OAI21_X1 U5762 ( .B1(n6283), .B2(n4772), .A(n4771), .ZN(n9259) );
  NAND2_X1 U5763 ( .A1(n6054), .A2(n6053), .ZN(n9372) );
  NAND2_X1 U5764 ( .A1(n4775), .A2(n4780), .ZN(n9277) );
  NAND2_X1 U5765 ( .A1(n6283), .A2(n4776), .ZN(n4775) );
  NAND2_X1 U5766 ( .A1(n6313), .A2(n6567), .ZN(n8023) );
  NAND2_X1 U5767 ( .A1(n9930), .A2(n4835), .ZN(n9924) );
  NAND2_X1 U5768 ( .A1(n4750), .A2(n4752), .ZN(n9720) );
  NAND2_X1 U5769 ( .A1(n4751), .A2(n4755), .ZN(n4750) );
  NAND2_X1 U5770 ( .A1(n4459), .A2(n5826), .ZN(n9660) );
  NAND2_X1 U5771 ( .A1(n5824), .A2(n4318), .ZN(n4459) );
  NAND2_X1 U5772 ( .A1(n7373), .A2(n6269), .ZN(n7439) );
  NAND2_X1 U5773 ( .A1(n7140), .A2(n6263), .ZN(n7205) );
  OAI211_X1 U5774 ( .C1(n5658), .C2(n6678), .A(n5624), .B(n5623), .ZN(n7400)
         );
  INV_X1 U5775 ( .A(n9925), .ZN(n9311) );
  INV_X1 U5776 ( .A(n9924), .ZN(n9739) );
  AND2_X1 U5777 ( .A1(n9930), .A2(n7158), .ZN(n9908) );
  NOR3_X1 U5778 ( .A1(n4641), .A2(n9743), .A3(n4640), .ZN(n9767) );
  AND2_X1 U5779 ( .A1(n9744), .A2(n9745), .ZN(n4640) );
  AND2_X1 U5780 ( .A1(n5625), .A2(n6220), .ZN(n9431) );
  NAND2_X1 U5781 ( .A1(n9431), .A2(n9430), .ZN(n9933) );
  XNOR2_X1 U5782 ( .A(n5585), .B(n5584), .ZN(n8320) );
  INV_X1 U5783 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5584) );
  NAND2_X1 U5784 ( .A1(n5617), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5585) );
  INV_X1 U5785 ( .A(n6214), .ZN(n8015) );
  XNOR2_X1 U5786 ( .A(n5612), .B(n5580), .ZN(n7892) );
  INV_X1 U5787 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7713) );
  INV_X1 U5788 ( .A(n6217), .ZN(n7579) );
  INV_X1 U5789 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7547) );
  NAND2_X1 U5790 ( .A1(n5630), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5602) );
  INV_X1 U5791 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7304) );
  AND2_X1 U5792 ( .A1(n5978), .A2(n5997), .ZN(n9138) );
  INV_X1 U5793 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7001) );
  INV_X1 U5794 ( .A(n7743), .ZN(n7736) );
  INV_X1 U5795 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6799) );
  INV_X1 U5796 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6771) );
  INV_X1 U5797 ( .A(n5707), .ZN(n6672) );
  XNOR2_X1 U5798 ( .A(n5660), .B(P1_IR_REG_1__SCAN_IN), .ZN(n9793) );
  OAI21_X1 U5799 ( .B1(n8838), .B2(n10022), .A(n4664), .ZN(P2_U3267) );
  AOI21_X1 U5800 ( .B1(n8836), .B2(n8829), .A(n4665), .ZN(n4664) );
  OAI21_X1 U5801 ( .B1(n8839), .B2(n8798), .A(n4666), .ZN(n4665) );
  INV_X1 U5802 ( .A(n8390), .ZN(n4666) );
  OAI21_X1 U5803 ( .B1(n8843), .B2(n10022), .A(n4502), .ZN(P2_U3268) );
  INV_X1 U5804 ( .A(n4503), .ZN(n4502) );
  OAI21_X1 U5805 ( .B1(n8844), .B2(n8798), .A(n4504), .ZN(n4503) );
  AOI21_X1 U5806 ( .B1(n8841), .B2(n8829), .A(n8625), .ZN(n4504) );
  OAI211_X1 U5807 ( .C1(n9144), .C2(n9272), .A(n4630), .B(n4629), .ZN(P1_U3260) );
  NOR2_X1 U5808 ( .A1(n4632), .A2(n4631), .ZN(n4630) );
  NAND2_X1 U5809 ( .A1(n4409), .A2(n9272), .ZN(n4629) );
  OAI21_X1 U5810 ( .B1(n9339), .B2(n9736), .A(n4610), .ZN(P1_U3263) );
  INV_X1 U5811 ( .A(n4611), .ZN(n4610) );
  OAI21_X1 U5812 ( .B1(n9340), .B2(n9325), .A(n4612), .ZN(n4611) );
  AOI21_X1 U5813 ( .B1(n9337), .B2(n9908), .A(n9173), .ZN(n4612) );
  NOR2_X1 U5814 ( .A1(n8246), .A2(n4583), .ZN(n4321) );
  AND2_X1 U5815 ( .A1(n4345), .A2(n4572), .ZN(n4322) );
  AND2_X1 U5816 ( .A1(n4345), .A2(n8242), .ZN(n4323) );
  MUX2_X1 U5817 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4852), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n4853) );
  AND4_X1 U5818 ( .A1(n5577), .A2(n5576), .A3(n5596), .A4(n5904), .ZN(n4324)
         );
  NOR2_X1 U5819 ( .A1(n8056), .A2(n8055), .ZN(n4498) );
  AOI21_X1 U5820 ( .B1(n4770), .B2(n9261), .A(n4779), .ZN(n4769) );
  AND2_X1 U5821 ( .A1(n6276), .A2(n4449), .ZN(n4325) );
  AND2_X1 U5822 ( .A1(n5881), .A2(n5858), .ZN(n4326) );
  AND2_X1 U5823 ( .A1(n7716), .A2(n7597), .ZN(n4327) );
  NAND2_X1 U5824 ( .A1(n4773), .A2(n9261), .ZN(n4328) );
  AND2_X1 U5825 ( .A1(n9759), .A2(n9075), .ZN(n4329) );
  AND2_X1 U5826 ( .A1(n4822), .A2(n8063), .ZN(n4330) );
  NAND2_X1 U5827 ( .A1(n5372), .A2(n5371), .ZN(n8874) );
  NOR2_X1 U5828 ( .A1(n6546), .A2(n4605), .ZN(n4331) );
  OR2_X1 U5829 ( .A1(n9351), .A2(n9061), .ZN(n6525) );
  INV_X1 U5830 ( .A(n8260), .ZN(n4811) );
  AND2_X1 U5831 ( .A1(n8148), .A2(n8141), .ZN(n8260) );
  AND2_X1 U5832 ( .A1(n9379), .A2(n9298), .ZN(n4332) );
  OR2_X1 U5833 ( .A1(n4735), .A2(n4734), .ZN(n4333) );
  NAND2_X1 U5834 ( .A1(n7968), .A2(n4681), .ZN(n4675) );
  INV_X1 U5835 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4850) );
  AND2_X1 U5836 ( .A1(n6270), .A2(n6269), .ZN(n4334) );
  NOR3_X1 U5837 ( .A1(n5515), .A2(n8440), .A3(n8415), .ZN(n4335) );
  INV_X1 U5838 ( .A(n9063), .ZN(n9194) );
  AND2_X1 U5839 ( .A1(n6169), .A2(n6168), .ZN(n9063) );
  AND2_X1 U5840 ( .A1(n8434), .A2(n8435), .ZN(n4683) );
  XNOR2_X1 U5841 ( .A(n4879), .B(P2_IR_REG_20__SCAN_IN), .ZN(n5519) );
  NOR2_X1 U5842 ( .A1(n4757), .A2(n4756), .ZN(n4755) );
  NAND2_X1 U5843 ( .A1(n5968), .A2(n5969), .ZN(n4336) );
  INV_X1 U5844 ( .A(n4317), .ZN(n5780) );
  INV_X1 U5845 ( .A(n7468), .ZN(n4425) );
  OR2_X1 U5846 ( .A1(n6470), .A2(n5652), .ZN(n4337) );
  AND2_X1 U5847 ( .A1(n5006), .A2(n6667), .ZN(n5075) );
  NAND2_X1 U5849 ( .A1(n5000), .A2(n4814), .ZN(n5019) );
  AND2_X1 U5850 ( .A1(n8801), .A2(n8358), .ZN(n4338) );
  AND2_X1 U5851 ( .A1(n9346), .A2(n8980), .ZN(n6521) );
  NAND3_X1 U5852 ( .A1(n4997), .A2(n4996), .A3(n4995), .ZN(n7025) );
  AND2_X1 U5853 ( .A1(n7723), .A2(n4820), .ZN(n4339) );
  OR2_X1 U5854 ( .A1(n7833), .A2(n4477), .ZN(n4340) );
  OR2_X1 U5855 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4341) );
  OR2_X1 U5856 ( .A1(n4735), .A2(n4733), .ZN(n4342) );
  XOR2_X1 U5857 ( .A(n8088), .B(n8815), .Z(n4343) );
  NOR2_X1 U5858 ( .A1(n6051), .A2(n9023), .ZN(n4344) );
  NAND2_X1 U5859 ( .A1(n8249), .A2(n8245), .ZN(n4345) );
  NAND2_X1 U5860 ( .A1(n5589), .A2(n8051), .ZN(n5674) );
  AND4_X1 U5861 ( .A1(n5600), .A2(n5597), .A3(n5579), .A4(n5578), .ZN(n4346)
         );
  OR2_X1 U5862 ( .A1(n7322), .A2(n7321), .ZN(n4347) );
  AND2_X1 U5863 ( .A1(n4911), .A2(SI_5_), .ZN(n4348) );
  AND2_X1 U5864 ( .A1(n4669), .A2(n4667), .ZN(n4349) );
  OR2_X1 U5865 ( .A1(n8801), .A2(n4496), .ZN(n4350) );
  OR2_X1 U5866 ( .A1(n4729), .A2(n9043), .ZN(n4351) );
  NOR2_X2 U5867 ( .A1(n5055), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n4871) );
  AND2_X1 U5868 ( .A1(n4849), .A2(n4500), .ZN(n4854) );
  AND2_X1 U5869 ( .A1(n6635), .A2(n6478), .ZN(n4352) );
  OR3_X1 U5870 ( .A1(n4328), .A2(n6279), .A3(n4454), .ZN(n4353) );
  INV_X1 U5871 ( .A(n6387), .ZN(n4604) );
  NAND2_X1 U5872 ( .A1(n5308), .A2(n5307), .ZN(n8892) );
  AND3_X1 U5873 ( .A1(n8241), .A2(n8243), .A3(n8240), .ZN(n4354) );
  INV_X1 U5874 ( .A(n9179), .ZN(n4767) );
  AND2_X1 U5875 ( .A1(n9166), .A2(n6523), .ZN(n9179) );
  NAND2_X1 U5876 ( .A1(n5980), .A2(n5979), .ZN(n9394) );
  AND3_X1 U5877 ( .A1(n6179), .A2(n6300), .A3(n6258), .ZN(n4355) );
  AND2_X1 U5878 ( .A1(n8213), .A2(n8214), .ZN(n8689) );
  AND3_X1 U5879 ( .A1(n6102), .A2(n9031), .A3(n6101), .ZN(n8951) );
  AND2_X1 U5880 ( .A1(n8142), .A2(n8150), .ZN(n8261) );
  NOR2_X1 U5881 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5000) );
  INV_X1 U5882 ( .A(n8372), .ZN(n8707) );
  AND2_X1 U5883 ( .A1(n8210), .A2(n8690), .ZN(n8372) );
  AND2_X1 U5884 ( .A1(n4825), .A2(n4824), .ZN(n4356) );
  INV_X1 U5885 ( .A(n8378), .ZN(n8845) );
  NAND2_X1 U5886 ( .A1(n5466), .A2(n5465), .ZN(n8378) );
  AND2_X1 U5887 ( .A1(n6264), .A2(n6263), .ZN(n4357) );
  AND2_X1 U5888 ( .A1(n8274), .A2(n7937), .ZN(n4358) );
  INV_X1 U5889 ( .A(n4777), .ZN(n4776) );
  OR2_X1 U5890 ( .A1(n6284), .A2(n4778), .ZN(n4777) );
  AND2_X1 U5891 ( .A1(n8869), .A2(n8505), .ZN(n4359) );
  INV_X1 U5892 ( .A(n4755), .ZN(n4754) );
  AND2_X1 U5893 ( .A1(n8065), .A2(n8217), .ZN(n4360) );
  OR2_X1 U5894 ( .A1(n8905), .A2(n8807), .ZN(n8191) );
  OR2_X1 U5895 ( .A1(n9242), .A2(n9038), .ZN(n4361) );
  INV_X1 U5896 ( .A(n8250), .ZN(n4563) );
  OR2_X1 U5897 ( .A1(n8840), .A2(n8234), .ZN(n8230) );
  INV_X1 U5898 ( .A(n8230), .ZN(n4580) );
  NOR2_X1 U5899 ( .A1(n9407), .A2(n9708), .ZN(n4362) );
  NOR2_X1 U5900 ( .A1(n9660), .A2(n9076), .ZN(n4363) );
  INV_X1 U5901 ( .A(n4681), .ZN(n4680) );
  NAND2_X1 U5902 ( .A1(n5296), .A2(n5297), .ZN(n4681) );
  OR2_X1 U5903 ( .A1(n4328), .A2(n4454), .ZN(n4364) );
  NOR2_X1 U5904 ( .A1(n8851), .A2(n8673), .ZN(n4365) );
  NOR2_X1 U5905 ( .A1(n8840), .A2(n8632), .ZN(n4366) );
  AND2_X1 U5906 ( .A1(n6484), .A2(n4439), .ZN(n4367) );
  INV_X1 U5907 ( .A(n4550), .ZN(n4549) );
  NAND2_X1 U5908 ( .A1(n4552), .A2(n4551), .ZN(n4550) );
  INV_X1 U5909 ( .A(n4773), .ZN(n4772) );
  NOR2_X1 U5910 ( .A1(n4774), .A2(n6285), .ZN(n4773) );
  AND2_X1 U5911 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4368) );
  NAND2_X1 U5912 ( .A1(n8706), .A2(n8061), .ZN(n8688) );
  INV_X1 U5913 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5603) );
  OR2_X1 U5914 ( .A1(n9759), .A2(n9075), .ZN(n4369) );
  XNOR2_X1 U5915 ( .A(n4891), .B(n4890), .ZN(n4998) );
  AND2_X1 U5916 ( .A1(n6667), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4370) );
  AND2_X1 U5917 ( .A1(n8094), .A2(n8096), .ZN(n8371) );
  AND2_X1 U5918 ( .A1(n4336), .A2(n9001), .ZN(n4371) );
  NOR2_X1 U5919 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(n4873), .ZN(n4372) );
  AND2_X1 U5920 ( .A1(n4527), .A2(n4958), .ZN(n4373) );
  NAND2_X1 U5921 ( .A1(n9407), .A2(n9708), .ZN(n4374) );
  NOR2_X1 U5922 ( .A1(n8491), .A2(n4521), .ZN(n4520) );
  AND2_X1 U5923 ( .A1(n9179), .A2(n4595), .ZN(n4375) );
  AND2_X1 U5924 ( .A1(n6429), .A2(n6513), .ZN(n4376) );
  AND2_X1 U5925 ( .A1(n8066), .A2(n4657), .ZN(n4377) );
  INV_X1 U5926 ( .A(n4816), .ZN(n4815) );
  NOR2_X1 U5927 ( .A1(n8270), .A2(n4817), .ZN(n4816) );
  AND2_X1 U5928 ( .A1(n4791), .A2(n5614), .ZN(n4378) );
  AND2_X1 U5929 ( .A1(n4944), .A2(n4937), .ZN(n4379) );
  OR2_X1 U5930 ( .A1(n4342), .A2(n4734), .ZN(n4380) );
  AND2_X1 U5931 ( .A1(n4510), .A2(n4928), .ZN(n4381) );
  NAND2_X1 U5932 ( .A1(n4730), .A2(n4734), .ZN(n4732) );
  INV_X1 U5933 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5597) );
  INV_X2 U5934 ( .A(n5658), .ZN(n5685) );
  XOR2_X1 U5935 ( .A(n8869), .B(n5550), .Z(n4382) );
  INV_X1 U5936 ( .A(n6101), .ZN(n4734) );
  AND2_X1 U5937 ( .A1(n7598), .A2(n7597), .ZN(n7717) );
  OR2_X1 U5938 ( .A1(n6157), .A2(n6156), .ZN(n4383) );
  AND2_X1 U5939 ( .A1(n6140), .A2(n6139), .ZN(n4384) );
  AND2_X1 U5940 ( .A1(n6754), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4385) );
  INV_X1 U5941 ( .A(n6567), .ZN(n4605) );
  AND2_X1 U5942 ( .A1(n6934), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4386) );
  OAI21_X1 U5943 ( .B1(n8729), .B2(n8367), .A(n8370), .ZN(n8715) );
  NAND2_X1 U5944 ( .A1(n6274), .A2(n6273), .ZN(n9698) );
  AND2_X1 U5945 ( .A1(n9194), .A2(n9710), .ZN(n4387) );
  NAND2_X1 U5946 ( .A1(n6283), .A2(n6282), .ZN(n9290) );
  INV_X1 U5947 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5580) );
  NAND2_X1 U5948 ( .A1(n7938), .A2(n4358), .ZN(n8359) );
  NAND2_X1 U5949 ( .A1(n8069), .A2(n8068), .ZN(n8835) );
  INV_X1 U5950 ( .A(n8835), .ZN(n4560) );
  NAND2_X1 U5951 ( .A1(n4705), .A2(n6159), .ZN(n9341) );
  INV_X1 U5952 ( .A(n9341), .ZN(n4766) );
  NAND2_X1 U5953 ( .A1(n9698), .A2(n6275), .ZN(n7916) );
  NAND2_X1 U5954 ( .A1(n5575), .A2(n5574), .ZN(n5860) );
  NOR3_X1 U5955 ( .A1(n7976), .A2(n9384), .A3(n4645), .ZN(n4642) );
  NAND2_X1 U5956 ( .A1(n8779), .A2(n4549), .ZN(n4553) );
  AND2_X1 U5957 ( .A1(n8419), .A2(n8514), .ZN(n4388) );
  NOR2_X1 U5958 ( .A1(n8896), .A2(n8771), .ZN(n4389) );
  INV_X1 U5959 ( .A(n4643), .ZN(n9308) );
  NOR2_X1 U5960 ( .A1(n7976), .A2(n4645), .ZN(n4643) );
  NAND2_X1 U5961 ( .A1(n4744), .A2(n4326), .ZN(n7821) );
  AND2_X1 U5962 ( .A1(n8039), .A2(n4336), .ZN(n4390) );
  AND2_X1 U5963 ( .A1(n5563), .A2(n5477), .ZN(n5517) );
  NOR2_X1 U5964 ( .A1(n8356), .A2(n4680), .ZN(n4391) );
  AND2_X1 U5965 ( .A1(n5278), .A2(n4963), .ZN(n4392) );
  XNOR2_X1 U5966 ( .A(n5627), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6217) );
  INV_X1 U5967 ( .A(n9904), .ZN(n4759) );
  NAND2_X1 U5968 ( .A1(n4849), .A2(n4871), .ZN(n4393) );
  NAND2_X1 U5969 ( .A1(n7714), .A2(n9272), .ZN(n6478) );
  NAND2_X1 U5970 ( .A1(n6993), .A2(n5715), .ZN(n7221) );
  INV_X1 U5971 ( .A(n8490), .ZN(n8474) );
  XNOR2_X1 U5972 ( .A(n5629), .B(P1_IR_REG_22__SCAN_IN), .ZN(n6216) );
  NAND2_X1 U5973 ( .A1(n7698), .A2(n4422), .ZN(n8447) );
  INV_X1 U5974 ( .A(n9759), .ZN(n4639) );
  AND2_X1 U5975 ( .A1(n7485), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4394) );
  NAND2_X1 U5976 ( .A1(n4747), .A2(n4749), .ZN(n7853) );
  NAND2_X1 U5977 ( .A1(n4795), .A2(n7091), .ZN(n7322) );
  NAND2_X1 U5978 ( .A1(n5357), .A2(n5356), .ZN(n8879) );
  INV_X1 U5979 ( .A(n8879), .ZN(n4551) );
  NAND2_X1 U5980 ( .A1(n5610), .A2(n5609), .ZN(n6196) );
  NAND2_X1 U5981 ( .A1(n5701), .A2(n5700), .ZN(n6991) );
  NAND2_X1 U5982 ( .A1(n7140), .A2(n4357), .ZN(n7204) );
  NAND2_X1 U5983 ( .A1(n5323), .A2(n5322), .ZN(n4395) );
  OR2_X1 U5984 ( .A1(n4782), .A2(n4784), .ZN(n4396) );
  AND2_X1 U5985 ( .A1(n5260), .A2(n5242), .ZN(n8003) );
  INV_X1 U5986 ( .A(n8003), .ZN(n7879) );
  OR2_X1 U5987 ( .A1(n7729), .A2(n8306), .ZN(n4397) );
  NAND2_X1 U5988 ( .A1(n4689), .A2(n4849), .ZN(n5497) );
  NAND2_X1 U5989 ( .A1(n5036), .A2(n5035), .ZN(n7244) );
  AND2_X1 U5990 ( .A1(n7549), .A2(n9222), .ZN(n7156) );
  INV_X1 U5991 ( .A(n7156), .ZN(n4743) );
  OR2_X1 U5992 ( .A1(n6659), .A2(n9222), .ZN(n4398) );
  NAND2_X1 U5993 ( .A1(n4972), .A2(n4971), .ZN(n5534) );
  AND2_X1 U5994 ( .A1(n6728), .A2(n6241), .ZN(n9886) );
  AND2_X1 U5995 ( .A1(n8578), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4399) );
  INV_X1 U5996 ( .A(n6857), .ZN(n4547) );
  XNOR2_X1 U5997 ( .A(n5602), .B(n5603), .ZN(n7549) );
  XNOR2_X1 U5998 ( .A(n5588), .B(n5587), .ZN(n8051) );
  INV_X1 U5999 ( .A(n4854), .ZN(n4663) );
  NOR2_X1 U6000 ( .A1(n5617), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n9433) );
  INV_X1 U6001 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n4538) );
  NOR2_X1 U6002 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n9655) );
  NOR2_X1 U6003 ( .A1(n6738), .A2(n6737), .ZN(n9829) );
  OAI21_X2 U6004 ( .B1(n8403), .B2(n8402), .A(n5405), .ZN(n4414) );
  OR2_X2 U6005 ( .A1(n8433), .A2(n4683), .ZN(n4522) );
  OAI21_X2 U6006 ( .B1(n8456), .B2(n8455), .A(n4413), .ZN(n8433) );
  NAND2_X1 U6007 ( .A1(n4414), .A2(n5421), .ZN(n4413) );
  XNOR2_X2 U6008 ( .A(n4414), .B(n5421), .ZN(n8456) );
  NAND3_X1 U6009 ( .A1(n8285), .A2(n5510), .A3(n8091), .ZN(n4415) );
  NAND2_X1 U6010 ( .A1(n4419), .A2(n5568), .ZN(n5543) );
  NAND2_X1 U6011 ( .A1(n7501), .A2(n5253), .ZN(n7588) );
  OAI21_X1 U6012 ( .B1(n5074), .B2(n4909), .A(n4430), .ZN(n5091) );
  NAND3_X1 U6013 ( .A1(n4429), .A2(n4428), .A3(n4912), .ZN(n4915) );
  NAND2_X1 U6014 ( .A1(n4430), .A2(n5074), .ZN(n4428) );
  NAND2_X1 U6015 ( .A1(n4909), .A2(n4430), .ZN(n4429) );
  NAND3_X1 U6016 ( .A1(n6408), .A2(n6528), .A3(n6407), .ZN(n4437) );
  NAND2_X1 U6017 ( .A1(n6274), .A2(n4325), .ZN(n4447) );
  NAND2_X1 U6018 ( .A1(n4447), .A2(n4448), .ZN(n6277) );
  NAND2_X1 U6019 ( .A1(n8664), .A2(n4462), .ZN(n4460) );
  NAND2_X1 U6020 ( .A1(n4460), .A2(n4461), .ZN(n8628) );
  NAND2_X1 U6021 ( .A1(n8359), .A2(n4467), .ZN(n4465) );
  NAND2_X1 U6022 ( .A1(n4465), .A2(n4466), .ZN(n8761) );
  NAND3_X1 U6023 ( .A1(n4327), .A2(n4816), .A3(n7598), .ZN(n4470) );
  XNOR2_X1 U6024 ( .A(n5129), .B(n5130), .ZN(n6691) );
  NAND3_X1 U6025 ( .A1(n6102), .A2(n4731), .A3(n9031), .ZN(n4474) );
  INV_X1 U6026 ( .A(n5937), .ZN(n5939) );
  NAND3_X1 U6027 ( .A1(n4745), .A2(n8039), .A3(n4371), .ZN(n4481) );
  NAND3_X1 U6028 ( .A1(n4482), .A2(n5701), .A3(n5700), .ZN(n6993) );
  NAND3_X1 U6029 ( .A1(n5710), .A2(n5711), .A3(n4483), .ZN(n7195) );
  INV_X1 U6030 ( .A(n4498), .ZN(n4497) );
  NAND2_X1 U6031 ( .A1(n4497), .A2(n8099), .ZN(n8802) );
  XNOR2_X2 U6032 ( .A(n4501), .B(n4851), .ZN(n4865) );
  INV_X1 U6033 ( .A(n7550), .ZN(n8522) );
  AND4_X2 U6034 ( .A1(n5010), .A2(n5009), .A3(n5008), .A4(n5007), .ZN(n7550)
         );
  NAND2_X1 U6035 ( .A1(n5005), .A2(n4505), .ZN(n4891) );
  NAND2_X1 U6036 ( .A1(n4968), .A2(n4889), .ZN(n5005) );
  INV_X2 U6037 ( .A(n4888), .ZN(n4968) );
  NAND3_X1 U6038 ( .A1(n4670), .A2(n4677), .A3(n4507), .ZN(n5382) );
  NAND2_X1 U6039 ( .A1(n4706), .A2(n4511), .ZN(n4509) );
  OAI21_X1 U6040 ( .B1(n4508), .B2(n4514), .A(n4924), .ZN(n5145) );
  INV_X1 U6041 ( .A(n4706), .ZN(n4508) );
  NAND2_X1 U6042 ( .A1(n4509), .A2(n4381), .ZN(n5165) );
  NAND2_X1 U6043 ( .A1(n8433), .A2(n4520), .ZN(n4517) );
  NAND2_X1 U6044 ( .A1(n4517), .A2(n4518), .ZN(n5518) );
  NAND2_X1 U6045 ( .A1(n4722), .A2(n4373), .ZN(n4523) );
  AND2_X2 U6046 ( .A1(n4546), .A2(n4848), .ZN(n4849) );
  INV_X2 U6047 ( .A(n5006), .ZN(n6766) );
  NAND2_X2 U6048 ( .A1(n4978), .A2(n4977), .ZN(n8949) );
  NAND2_X1 U6049 ( .A1(n4548), .A2(n8779), .ZN(n8716) );
  INV_X1 U6050 ( .A(n4553), .ZN(n8732) );
  AND2_X1 U6051 ( .A1(n8655), .A2(n4559), .ZN(n8610) );
  NAND2_X1 U6052 ( .A1(n8655), .A2(n4557), .ZN(n8604) );
  NAND2_X1 U6053 ( .A1(n8655), .A2(n4561), .ZN(n8614) );
  NAND2_X1 U6054 ( .A1(n8655), .A2(n8845), .ZN(n8635) );
  OAI21_X1 U6055 ( .B1(n4568), .B2(n4567), .A(n4583), .ZN(n4566) );
  OAI21_X1 U6056 ( .B1(n4354), .B2(n4571), .A(n4570), .ZN(n8247) );
  INV_X1 U6057 ( .A(n8244), .ZN(n4572) );
  NAND2_X1 U6058 ( .A1(n8232), .A2(n4576), .ZN(n4575) );
  NAND3_X1 U6059 ( .A1(n8105), .A2(n8108), .A3(n4583), .ZN(n4582) );
  OR2_X1 U6060 ( .A1(n8517), .A2(n10044), .ZN(n8108) );
  OR2_X1 U6061 ( .A1(n8518), .A2(n7087), .ZN(n8105) );
  OAI21_X1 U6062 ( .B1(n4588), .B2(n4587), .A(n4585), .ZN(n8218) );
  AOI21_X1 U6063 ( .B1(n8209), .B2(n8372), .A(n8216), .ZN(n4588) );
  NAND4_X1 U6064 ( .A1(n4589), .A2(n4848), .A3(n4870), .A4(n4871), .ZN(n4971)
         );
  NAND2_X1 U6065 ( .A1(n4971), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4852) );
  INV_X2 U6066 ( .A(n5315), .ZN(n5045) );
  NAND4_X1 U6067 ( .A1(n4590), .A2(n5574), .A3(n4324), .A4(n5575), .ZN(n5611)
         );
  OAI21_X1 U6068 ( .B1(n9214), .B2(n4598), .A(n4594), .ZN(n9167) );
  AOI21_X1 U6069 ( .B1(n9214), .B2(n6621), .A(n6318), .ZN(n9193) );
  OAI21_X1 U6070 ( .B1(n6388), .B2(n4604), .A(n9705), .ZN(n4600) );
  NAND2_X1 U6071 ( .A1(n9316), .A2(n6531), .ZN(n4606) );
  NAND3_X1 U6072 ( .A1(n6555), .A2(n6599), .A3(n6608), .ZN(n4609) );
  NAND3_X1 U6073 ( .A1(n4609), .A2(n6606), .A3(n4607), .ZN(n7385) );
  NAND2_X1 U6074 ( .A1(n6608), .A2(n4608), .ZN(n4607) );
  NAND2_X1 U6075 ( .A1(n7145), .A2(n6603), .ZN(n7208) );
  NAND2_X1 U6076 ( .A1(n5581), .A2(n4615), .ZN(n5617) );
  NOR2_X1 U6077 ( .A1(n8054), .A2(n6667), .ZN(n4668) );
  OR2_X2 U6078 ( .A1(n9728), .A2(n6383), .ZN(n7860) );
  NAND2_X1 U6079 ( .A1(n9851), .A2(n4626), .ZN(n4624) );
  NAND2_X1 U6080 ( .A1(n4624), .A2(n4625), .ZN(n6776) );
  INV_X1 U6081 ( .A(n4633), .ZN(n9808) );
  NAND2_X1 U6082 ( .A1(n4633), .A2(n9809), .ZN(n6726) );
  NAND2_X1 U6083 ( .A1(n9794), .A2(n4634), .ZN(n4633) );
  NAND2_X1 U6084 ( .A1(n9793), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4634) );
  INV_X1 U6085 ( .A(n9721), .ZN(n4635) );
  NAND2_X1 U6086 ( .A1(n4635), .A2(n4636), .ZN(n7960) );
  NOR2_X1 U6087 ( .A1(n9742), .A2(n9973), .ZN(n4641) );
  NOR2_X2 U6088 ( .A1(n9219), .A2(n9351), .ZN(n9200) );
  INV_X1 U6089 ( .A(n4642), .ZN(n9291) );
  OAI21_X2 U6090 ( .B1(n5604), .B2(n5583), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4647) );
  INV_X1 U6091 ( .A(n6891), .ZN(n9329) );
  NOR2_X1 U6092 ( .A1(n7395), .A2(n7400), .ZN(n7154) );
  NAND3_X1 U6093 ( .A1(n7011), .A2(n6891), .A3(n9936), .ZN(n7395) );
  AND3_X2 U6094 ( .A1(n5687), .A2(n5686), .A3(n5688), .ZN(n6891) );
  NAND2_X1 U6095 ( .A1(n7536), .A2(n4651), .ZN(n4648) );
  NAND2_X1 U6096 ( .A1(n4648), .A2(n4649), .ZN(n7725) );
  AOI21_X1 U6097 ( .B1(n8648), .B2(n4377), .A(n4654), .ZN(n8383) );
  NAND2_X1 U6098 ( .A1(n8648), .A2(n4657), .ZN(n8629) );
  OR2_X2 U6099 ( .A1(n7625), .A2(n7624), .ZN(n8412) );
  NAND2_X1 U6100 ( .A1(n8473), .A2(n5109), .ZN(n7625) );
  NAND2_X1 U6101 ( .A1(n5006), .A2(n4370), .ZN(n4669) );
  NAND2_X1 U6102 ( .A1(n8356), .A2(n4671), .ZN(n4670) );
  NAND2_X1 U6103 ( .A1(n7659), .A2(n5274), .ZN(n7810) );
  INV_X1 U6104 ( .A(n4685), .ZN(n7809) );
  INV_X1 U6105 ( .A(n7811), .ZN(n4687) );
  NAND2_X1 U6106 ( .A1(n4849), .A2(n4690), .ZN(n4974) );
  NAND2_X1 U6107 ( .A1(n5300), .A2(n5299), .ZN(n4700) );
  OAI21_X1 U6108 ( .B1(n5300), .B2(n4697), .A(n4695), .ZN(n5353) );
  NAND2_X1 U6109 ( .A1(n4694), .A2(n4692), .ZN(n5355) );
  NAND2_X1 U6110 ( .A1(n5300), .A2(n4695), .ZN(n4694) );
  NAND2_X1 U6111 ( .A1(n4701), .A2(n6647), .ZN(P1_U3240) );
  NAND2_X1 U6112 ( .A1(n4702), .A2(n6642), .ZN(n4701) );
  NAND3_X1 U6113 ( .A1(n4703), .A2(n6593), .A3(n6639), .ZN(n4702) );
  NAND3_X1 U6114 ( .A1(n6485), .A2(n4704), .A3(n6633), .ZN(n4703) );
  NAND2_X1 U6115 ( .A1(n9341), .A2(n9063), .ZN(n6523) );
  NAND2_X1 U6116 ( .A1(n6440), .A2(n4707), .ZN(n4710) );
  NAND2_X1 U6117 ( .A1(n8342), .A2(n9071), .ZN(n4711) );
  NAND2_X1 U6118 ( .A1(n4712), .A2(n4392), .ZN(n4967) );
  NAND2_X1 U6119 ( .A1(n4713), .A2(n4937), .ZN(n5197) );
  NAND2_X1 U6120 ( .A1(n4713), .A2(n4379), .ZN(n4946) );
  NAND2_X1 U6121 ( .A1(n4933), .A2(n4932), .ZN(n5182) );
  NAND2_X1 U6122 ( .A1(n5422), .A2(n4719), .ZN(n4716) );
  OAI21_X1 U6123 ( .B1(n5422), .B2(n4721), .A(n5425), .ZN(n5442) );
  NAND2_X1 U6124 ( .A1(n4716), .A2(n4717), .ZN(n5458) );
  MUX2_X1 U6125 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n4968), .Z(n4895) );
  MUX2_X1 U6126 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n4968), .Z(n4999) );
  INV_X1 U6127 ( .A(n5996), .ZN(n4729) );
  INV_X1 U6128 ( .A(n4736), .ZN(n8953) );
  INV_X1 U6129 ( .A(n7520), .ZN(n5820) );
  NAND2_X1 U6130 ( .A1(n5601), .A2(n4742), .ZN(n4741) );
  NAND2_X1 U6131 ( .A1(n5601), .A2(n5600), .ZN(n5630) );
  AND2_X2 U6132 ( .A1(n6300), .A2(n6179), .ZN(n6193) );
  INV_X1 U6133 ( .A(n6216), .ZN(n7714) );
  NAND2_X1 U6134 ( .A1(n9056), .A2(n4383), .ZN(n6650) );
  INV_X1 U6135 ( .A(n9902), .ZN(n4751) );
  NAND2_X1 U6136 ( .A1(n4748), .A2(n9902), .ZN(n4747) );
  OAI21_X1 U6137 ( .B1(n9902), .B2(n6272), .A(n4758), .ZN(n7608) );
  INV_X1 U6138 ( .A(n9174), .ZN(n4768) );
  AND2_X1 U6139 ( .A1(n9372), .A2(n9285), .ZN(n4779) );
  OR2_X1 U6140 ( .A1(n9384), .A2(n9319), .ZN(n4780) );
  NAND2_X1 U6141 ( .A1(n7975), .A2(n7982), .ZN(n8017) );
  NAND2_X1 U6142 ( .A1(n7373), .A2(n4334), .ZN(n7437) );
  NAND2_X1 U6143 ( .A1(n5581), .A2(n5580), .ZN(n5604) );
  OAI21_X1 U6144 ( .B1(n7045), .B2(n4794), .A(n4792), .ZN(n4795) );
  OAI21_X1 U6145 ( .B1(n4794), .B2(n8257), .A(n8256), .ZN(n4793) );
  OAI211_X1 U6146 ( .C1(n8626), .C2(n4803), .A(n4799), .B(n4796), .ZN(n8839)
         );
  NAND2_X1 U6147 ( .A1(n8626), .A2(n4797), .ZN(n4796) );
  NOR2_X1 U6148 ( .A1(n4798), .A2(n8377), .ZN(n4797) );
  NAND2_X1 U6149 ( .A1(n4804), .A2(n8377), .ZN(n4800) );
  NAND3_X1 U6150 ( .A1(n4806), .A2(n7041), .A3(n7059), .ZN(n7043) );
  INV_X1 U6151 ( .A(n7534), .ZN(n7532) );
  NAND2_X1 U6152 ( .A1(n8715), .A2(n4823), .ZN(n4821) );
  INV_X1 U6153 ( .A(n5670), .ZN(n5671) );
  NAND2_X1 U6154 ( .A1(n6812), .A2(n5651), .ZN(n5670) );
  OAI21_X2 U6155 ( .B1(n9252), .B2(n6489), .A(n6421), .ZN(n9230) );
  NAND2_X1 U6156 ( .A1(n6214), .A2(n5613), .ZN(n5625) );
  INV_X1 U6157 ( .A(n5631), .ZN(n5601) );
  NAND2_X1 U6158 ( .A1(n4903), .A2(n4902), .ZN(n5058) );
  INV_X2 U6159 ( .A(n6662), .ZN(n5708) );
  NAND2_X1 U6160 ( .A1(n6662), .A2(n6667), .ZN(n5658) );
  INV_X1 U6161 ( .A(n6097), .ZN(n6100) );
  NAND2_X1 U6162 ( .A1(n7026), .A2(n7025), .ZN(n8120) );
  OR2_X1 U6163 ( .A1(n8729), .A2(n8751), .ZN(n8885) );
  OAI21_X1 U6164 ( .B1(n8346), .B2(n9945), .A(n6332), .ZN(n6340) );
  NAND2_X1 U6165 ( .A1(n8076), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n4996) );
  OR2_X1 U6166 ( .A1(n5006), .A2(n6855), .ZN(n5001) );
  AOI21_X1 U6167 ( .B1(n8718), .B2(n5525), .A(n5379), .ZN(n8427) );
  NAND2_X1 U6168 ( .A1(n5525), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n4995) );
  INV_X1 U6169 ( .A(n8320), .ZN(n5589) );
  NAND2_X1 U6170 ( .A1(n5673), .A2(n6881), .ZN(n6889) );
  NOR2_X1 U6171 ( .A1(n8879), .A2(n8749), .ZN(n4829) );
  AND2_X2 U6172 ( .A1(n6339), .A2(n7151), .ZN(n9980) );
  NAND3_X1 U6173 ( .A1(n8247), .A2(n8285), .A3(n5510), .ZN(n4830) );
  INV_X1 U6174 ( .A(n6517), .ZN(n6298) );
  AND3_X1 U6175 ( .A1(n5564), .A2(n5563), .A3(n8474), .ZN(n4831) );
  AND2_X1 U6176 ( .A1(n9179), .A2(n6429), .ZN(n4832) );
  AND2_X1 U6177 ( .A1(n6649), .A2(n6648), .ZN(n4833) );
  AND2_X1 U6178 ( .A1(n6649), .A2(n6223), .ZN(n4834) );
  INV_X1 U6179 ( .A(n7549), .ZN(n6639) );
  INV_X1 U6180 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7661) );
  INV_X1 U6181 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n4905) );
  INV_X1 U6182 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5151) );
  INV_X1 U6183 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8437) );
  AND2_X1 U6184 ( .A1(n7157), .A2(n6639), .ZN(n4835) );
  OR2_X1 U6185 ( .A1(n4888), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8318) );
  INV_X1 U6186 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n4899) );
  NAND2_X1 U6187 ( .A1(n8123), .A2(n8122), .ZN(n7059) );
  INV_X2 U6188 ( .A(n10078), .ZN(n10080) );
  INV_X1 U6189 ( .A(n5799), .ZN(n5794) );
  AND2_X1 U6190 ( .A1(n5542), .A2(n5541), .ZN(n4836) );
  NAND2_X2 U6191 ( .A1(n7342), .A2(n10025), .ZN(n10009) );
  AND2_X1 U6192 ( .A1(n6443), .A2(n6478), .ZN(n6444) );
  INV_X1 U6193 ( .A(n7498), .ZN(n5225) );
  AND2_X1 U6194 ( .A1(n5649), .A2(n7167), .ZN(n5650) );
  OR4_X1 U6195 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6204) );
  INV_X1 U6196 ( .A(n8645), .ZN(n8065) );
  INV_X1 U6197 ( .A(n7442), .ZN(n6270) );
  INV_X1 U6198 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4885) );
  OR2_X1 U6199 ( .A1(n5404), .A2(n4382), .ZN(n5405) );
  INV_X1 U6200 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9541) );
  OR2_X1 U6201 ( .A1(n5432), .A2(n8437), .ZN(n5449) );
  NAND2_X1 U6202 ( .A1(n7242), .A2(n8823), .ZN(n8122) );
  INV_X1 U6203 ( .A(n5956), .ZN(n5954) );
  NAND2_X1 U6204 ( .A1(n5682), .A2(n7235), .ZN(n5646) );
  INV_X1 U6205 ( .A(n6035), .ZN(n6033) );
  AOI22_X1 U6206 ( .A1(n9180), .A2(n9710), .B1(n9148), .B2(n9070), .ZN(n6328)
         );
  INV_X1 U6207 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8971) );
  INV_X1 U6208 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5808) );
  INV_X1 U6209 ( .A(SI_27_), .ZN(n9518) );
  INV_X1 U6210 ( .A(SI_20_), .ZN(n9529) );
  INV_X1 U6211 ( .A(SI_16_), .ZN(n9577) );
  NAND2_X1 U6212 ( .A1(n6667), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n4904) );
  NAND2_X1 U6213 ( .A1(n5215), .A2(n5214), .ZN(n7504) );
  OR2_X1 U6214 ( .A1(n8299), .A2(n5194), .ZN(n5195) );
  OR2_X1 U6215 ( .A1(n5374), .A2(n9541), .ZN(n5396) );
  OR2_X1 U6216 ( .A1(n5311), .A2(n5310), .ZN(n5333) );
  OR2_X1 U6217 ( .A1(n5173), .A2(n9586), .ZN(n5188) );
  INV_X1 U6218 ( .A(n8091), .ZN(n8286) );
  NAND2_X1 U6219 ( .A1(n7894), .A2(n7905), .ZN(n7896) );
  INV_X1 U6220 ( .A(n8263), .ZN(n7531) );
  NAND2_X1 U6221 ( .A1(n8632), .A2(n8788), .ZN(n8387) );
  INV_X1 U6222 ( .A(n10032), .ZN(n5505) );
  INV_X1 U6223 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n4851) );
  NOR2_X1 U6224 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n4874) );
  INV_X1 U6225 ( .A(n7824), .ZN(n5881) );
  OR2_X1 U6226 ( .A1(n6181), .A2(n6180), .ZN(n6230) );
  OR2_X1 U6227 ( .A1(n6074), .A2(n9034), .ZN(n6109) );
  NAND2_X1 U6228 ( .A1(n6033), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6055) );
  INV_X1 U6229 ( .A(n6328), .ZN(n6329) );
  OR2_X1 U6230 ( .A1(n9363), .A2(n9254), .ZN(n6287) );
  OR2_X1 U6231 ( .A1(n5809), .A2(n5808), .ZN(n5827) );
  INV_X1 U6232 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6209) );
  OR2_X1 U6233 ( .A1(n9903), .A2(n9904), .ZN(n9905) );
  NOR2_X1 U6234 ( .A1(n6196), .A2(n7892), .ZN(n5613) );
  INV_X1 U6235 ( .A(SI_29_), .ZN(n6448) );
  INV_X1 U6236 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5600) );
  AND2_X1 U6237 ( .A1(n5540), .A2(n5539), .ZN(n5541) );
  NAND2_X1 U6238 ( .A1(n5054), .A2(n7245), .ZN(n7247) );
  INV_X1 U6239 ( .A(n5381), .ZN(n5373) );
  INV_X1 U6240 ( .A(n8293), .ZN(n5536) );
  INV_X1 U6241 ( .A(n8479), .ZN(n8494) );
  NAND2_X1 U6242 ( .A1(n5448), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5523) );
  AND2_X1 U6243 ( .A1(n5396), .A2(n5375), .ZN(n8718) );
  INV_X1 U6244 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9586) );
  INV_X1 U6245 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7803) );
  INV_X1 U6246 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9604) );
  INV_X1 U6247 ( .A(n9991), .ZN(n9996) );
  INV_X1 U6248 ( .A(n8512), .ZN(n8329) );
  INV_X1 U6249 ( .A(n8790), .ZN(n8806) );
  INV_X1 U6250 ( .A(n8451), .ZN(n10044) );
  NAND2_X1 U6251 ( .A1(n5937), .A2(n5921), .ZN(n7989) );
  OR2_X1 U6252 ( .A1(n5981), .A2(n9003), .ZN(n6003) );
  OR2_X1 U6253 ( .A1(n6019), .A2(n6018), .ZN(n6035) );
  INV_X1 U6254 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7561) );
  INV_X1 U6255 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9003) );
  INV_X1 U6256 ( .A(n9233), .ZN(n6349) );
  AND2_X1 U6257 ( .A1(n8337), .A2(n6331), .ZN(n6332) );
  AND2_X1 U6258 ( .A1(n6322), .A2(n6727), .ZN(n9710) );
  INV_X1 U6259 ( .A(n9395), .ZN(n9973) );
  INV_X1 U6260 ( .A(n9919), .ZN(n9732) );
  INV_X1 U6261 ( .A(n9745), .ZN(n9972) );
  NAND2_X1 U6262 ( .A1(n6451), .A2(n6450), .ZN(n6455) );
  AND2_X1 U6263 ( .A1(n4928), .A2(n4927), .ZN(n5146) );
  OAI21_X1 U6264 ( .B1(n6667), .B2(n4899), .A(n4898), .ZN(n4901) );
  OR3_X1 U6265 ( .A1(n7915), .A2(n7936), .A3(n8030), .ZN(n6833) );
  XNOR2_X1 U6266 ( .A(n8306), .B(n5550), .ZN(n5228) );
  NAND2_X1 U6267 ( .A1(n5144), .A2(n8410), .ZN(n8416) );
  AND2_X1 U6268 ( .A1(n8477), .A2(n8790), .ZN(n8465) );
  AND2_X1 U6269 ( .A1(n5533), .A2(n5536), .ZN(n8477) );
  OR2_X1 U6270 ( .A1(n8656), .A2(n5558), .ZN(n5455) );
  INV_X1 U6271 ( .A(n8076), .ZN(n5528) );
  AND2_X1 U6272 ( .A1(n6836), .A2(n6835), .ZN(n9991) );
  INV_X1 U6273 ( .A(n8376), .ZN(n8377) );
  INV_X1 U6274 ( .A(n8371), .ZN(n8723) );
  AND2_X1 U6275 ( .A1(n6831), .A2(n6830), .ZN(n8788) );
  AND2_X1 U6276 ( .A1(n8166), .A2(n8165), .ZN(n8269) );
  AND2_X1 U6277 ( .A1(n10009), .A2(n7340), .ZN(n7767) );
  AND2_X1 U6278 ( .A1(n10011), .A2(n9683), .ZN(n8829) );
  NOR2_X1 U6279 ( .A1(n7073), .A2(n7072), .ZN(n7074) );
  AND2_X1 U6280 ( .A1(n7021), .A2(n7020), .ZN(n7075) );
  AND2_X1 U6281 ( .A1(n7760), .A2(n9685), .ZN(n8914) );
  INV_X1 U6282 ( .A(n8914), .ZN(n10068) );
  AND2_X1 U6283 ( .A1(n5501), .A2(n5500), .ZN(n10026) );
  NAND2_X1 U6284 ( .A1(n5493), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5495) );
  AND2_X1 U6285 ( .A1(n5183), .A2(n5170), .ZN(n7649) );
  OAI22_X1 U6286 ( .A1(n6889), .A2(n6890), .B1(n5696), .B2(n5695), .ZN(n6823)
         );
  AND2_X1 U6287 ( .A1(n6247), .A2(n6229), .ZN(n7318) );
  INV_X1 U6288 ( .A(n9062), .ZN(n9024) );
  NAND2_X1 U6289 ( .A1(n6248), .A2(n6247), .ZN(n9066) );
  INV_X1 U6290 ( .A(n6641), .ZN(n6642) );
  AND2_X1 U6291 ( .A1(n6188), .A2(n6187), .ZN(n6651) );
  INV_X1 U6292 ( .A(n6703), .ZN(n9866) );
  INV_X1 U6293 ( .A(n9899), .ZN(n9880) );
  INV_X1 U6294 ( .A(n9886), .ZN(n9114) );
  AND2_X1 U6295 ( .A1(n6719), .A2(n6718), .ZN(n9894) );
  AOI21_X1 U6296 ( .B1(n9185), .B2(n6511), .A(n6513), .ZN(n9174) );
  AND2_X1 U6297 ( .A1(n6570), .A2(n9315), .ZN(n8022) );
  AND2_X1 U6298 ( .A1(n6392), .A2(n6563), .ZN(n7920) );
  INV_X1 U6299 ( .A(n9922), .ZN(n9735) );
  AND2_X1 U6300 ( .A1(n6211), .A2(n9432), .ZN(n7377) );
  AND2_X1 U6301 ( .A1(n9922), .A2(n9659), .ZN(n9945) );
  INV_X1 U6302 ( .A(n7377), .ZN(n7151) );
  AND2_X1 U6303 ( .A1(n5728), .A2(n5758), .ZN(n9849) );
  OAI21_X1 U6304 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10086), .ZN(n10117) );
  INV_X1 U6305 ( .A(n8602), .ZN(n9994) );
  INV_X1 U6306 ( .A(n7025), .ZN(n7556) );
  OR2_X1 U6307 ( .A1(n4992), .A2(n4991), .ZN(n8506) );
  INV_X1 U6308 ( .A(n8596), .ZN(n9995) );
  NAND2_X1 U6309 ( .A1(n6842), .A2(n6841), .ZN(n9997) );
  INV_X1 U6310 ( .A(n8829), .ZN(n10019) );
  NAND2_X1 U6311 ( .A1(n10009), .A2(n10014), .ZN(n8798) );
  NAND2_X1 U6312 ( .A1(n7075), .A2(n7074), .ZN(n10078) );
  INV_X1 U6313 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10031) );
  INV_X1 U6314 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8948) );
  INV_X1 U6315 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8401) );
  INV_X1 U6316 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6811) );
  NAND2_X1 U6317 ( .A1(n6224), .A2(n6223), .ZN(n6256) );
  INV_X1 U6318 ( .A(n9357), .ZN(n9019) );
  INV_X1 U6319 ( .A(n6651), .ZN(n9180) );
  NAND2_X1 U6320 ( .A1(n6081), .A2(n6080), .ZN(n9265) );
  INV_X1 U6321 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9842) );
  OR2_X1 U6322 ( .A1(P1_U3083), .A2(n9804), .ZN(n9899) );
  NAND2_X1 U6323 ( .A1(n9930), .A2(n7169), .ZN(n9325) );
  NAND2_X1 U6324 ( .A1(n6336), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6337) );
  AND2_X2 U6325 ( .A1(n6339), .A2(n7377), .ZN(n9990) );
  AND2_X1 U6326 ( .A1(n9757), .A2(n9756), .ZN(n9771) );
  AND2_X1 U6327 ( .A1(n9764), .A2(n9763), .ZN(n9773) );
  AND3_X1 U6328 ( .A1(n9952), .A2(n9951), .A3(n9950), .ZN(n9984) );
  INV_X1 U6329 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8014) );
  INV_X1 U6330 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7102) );
  INV_X1 U6331 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6709) );
  AND2_X1 U6332 ( .A1(n6663), .A2(n10033), .ZN(P2_U3966) );
  AND2_X2 U6333 ( .A1(n9804), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  NOR2_X1 U6334 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n4840) );
  NOR2_X1 U6335 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n4839) );
  NOR2_X1 U6336 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n4838) );
  NAND4_X1 U6337 ( .A1(n4841), .A2(n4840), .A3(n4839), .A4(n4838), .ZN(n5486)
         );
  INV_X1 U6338 ( .A(n5486), .ZN(n4848) );
  NOR2_X1 U6339 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n4847) );
  NOR2_X1 U6340 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n4843) );
  NAND4_X1 U6341 ( .A1(n4843), .A2(n4842), .A3(n5166), .A4(n5237), .ZN(n4846)
         );
  NAND4_X1 U6342 ( .A1(n4844), .A2(n5240), .A3(n5168), .A4(n5112), .ZN(n4845)
         );
  NOR2_X2 U6343 ( .A1(n4846), .A2(n4845), .ZN(n4870) );
  AND2_X4 U6344 ( .A1(n4865), .A2(n4866), .ZN(n8076) );
  INV_X1 U6345 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n4869) );
  NAND3_X1 U6346 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n5098) );
  INV_X1 U6347 ( .A(n5098), .ZN(n4855) );
  NAND2_X1 U6348 ( .A1(n4855), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5118) );
  INV_X1 U6349 ( .A(n5118), .ZN(n4856) );
  NAND2_X1 U6350 ( .A1(n4856), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5134) );
  INV_X1 U6351 ( .A(n5134), .ZN(n4857) );
  NAND2_X1 U6352 ( .A1(n4857), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5152) );
  INV_X1 U6353 ( .A(n5188), .ZN(n4858) );
  NAND2_X1 U6354 ( .A1(n4858), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5202) );
  INV_X1 U6355 ( .A(n5202), .ZN(n4859) );
  NAND2_X1 U6356 ( .A1(n4859), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5216) );
  INV_X1 U6357 ( .A(n5246), .ZN(n4860) );
  NAND2_X1 U6358 ( .A1(n4860), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5264) );
  INV_X1 U6359 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n4863) );
  NAND2_X1 U6360 ( .A1(n5288), .A2(n4863), .ZN(n4864) );
  NAND2_X1 U6361 ( .A1(n5311), .A2(n4864), .ZN(n8794) );
  INV_X2 U6362 ( .A(n4865), .ZN(n8936) );
  AND2_X4 U6363 ( .A1(n8939), .A2(n8936), .ZN(n5525) );
  OR2_X1 U6364 ( .A1(n8794), .A2(n5558), .ZN(n4868) );
  AOI22_X1 U6365 ( .A1(n5045), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n5025), .B2(
        P2_REG2_REG_18__SCAN_IN), .ZN(n4867) );
  OAI211_X1 U6366 ( .C1(n5528), .C2(n4869), .A(n4868), .B(n4867), .ZN(n8771)
         );
  AND2_X2 U6367 ( .A1(n4871), .A2(n4872), .ZN(n5113) );
  NAND2_X1 U6368 ( .A1(n4878), .A2(n4874), .ZN(n4875) );
  OAI21_X2 U6369 ( .B1(n4875), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5491) );
  NAND2_X1 U6370 ( .A1(n4875), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4877) );
  OR2_X4 U6371 ( .A1(n5510), .A2(n8293), .ZN(n8090) );
  NAND2_X1 U6372 ( .A1(n8771), .A2(n8090), .ZN(n5293) );
  INV_X1 U6373 ( .A(n5293), .ZN(n5297) );
  NAND2_X1 U6374 ( .A1(n9655), .A2(n4884), .ZN(n4887) );
  NAND2_X1 U6375 ( .A1(n4888), .A2(SI_0_), .ZN(n5642) );
  AND2_X1 U6376 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4889) );
  INV_X1 U6377 ( .A(SI_1_), .ZN(n4890) );
  NAND2_X1 U6378 ( .A1(n4998), .A2(n4999), .ZN(n4893) );
  NAND2_X1 U6379 ( .A1(n4891), .A2(SI_1_), .ZN(n4892) );
  NAND2_X1 U6380 ( .A1(n4893), .A2(n4892), .ZN(n5016) );
  INV_X1 U6381 ( .A(SI_2_), .ZN(n4894) );
  NAND2_X1 U6382 ( .A1(n5016), .A2(n5017), .ZN(n4897) );
  NAND2_X1 U6383 ( .A1(n4895), .A2(SI_2_), .ZN(n4896) );
  NAND2_X1 U6384 ( .A1(n4897), .A2(n4896), .ZN(n5038) );
  INV_X1 U6385 ( .A(SI_3_), .ZN(n4900) );
  XNOR2_X1 U6386 ( .A(n4901), .B(n4900), .ZN(n5039) );
  NAND2_X1 U6387 ( .A1(n5038), .A2(n5039), .ZN(n4903) );
  NAND2_X1 U6388 ( .A1(n4901), .A2(SI_3_), .ZN(n4902) );
  XNOR2_X1 U6389 ( .A(n4907), .B(SI_4_), .ZN(n5059) );
  INV_X1 U6390 ( .A(n5059), .ZN(n4906) );
  NAND2_X1 U6391 ( .A1(n5058), .A2(n4906), .ZN(n4909) );
  NAND2_X1 U6392 ( .A1(n4907), .A2(SI_4_), .ZN(n4908) );
  MUX2_X1 U6393 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n4888), .Z(n4911) );
  INV_X1 U6394 ( .A(n5074), .ZN(n4910) );
  MUX2_X1 U6395 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6667), .Z(n4913) );
  XNOR2_X1 U6396 ( .A(n4913), .B(SI_6_), .ZN(n5092) );
  INV_X1 U6397 ( .A(n5092), .ZN(n4912) );
  NAND2_X1 U6398 ( .A1(n4913), .A2(SI_6_), .ZN(n4914) );
  NAND2_X1 U6399 ( .A1(n4915), .A2(n4914), .ZN(n5110) );
  MUX2_X1 U6400 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6667), .Z(n4917) );
  XNOR2_X1 U6401 ( .A(n4917), .B(SI_7_), .ZN(n5111) );
  INV_X1 U6402 ( .A(n5111), .ZN(n4916) );
  NAND2_X1 U6403 ( .A1(n4917), .A2(SI_7_), .ZN(n4918) );
  INV_X1 U6404 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6694) );
  INV_X1 U6405 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6692) );
  MUX2_X1 U6406 ( .A(n6694), .B(n6692), .S(n6667), .Z(n4920) );
  INV_X1 U6407 ( .A(SI_8_), .ZN(n4919) );
  NAND2_X1 U6408 ( .A1(n4920), .A2(n4919), .ZN(n4924) );
  INV_X1 U6409 ( .A(n4920), .ZN(n4921) );
  NAND2_X1 U6410 ( .A1(n4921), .A2(SI_8_), .ZN(n4922) );
  NAND2_X1 U6411 ( .A1(n4924), .A2(n4922), .ZN(n5130) );
  INV_X1 U6412 ( .A(n5130), .ZN(n4923) );
  INV_X1 U6413 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6705) );
  INV_X1 U6414 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6702) );
  MUX2_X1 U6415 ( .A(n6705), .B(n6702), .S(n6667), .Z(n4925) );
  NAND2_X1 U6416 ( .A1(n4925), .A2(n9520), .ZN(n4928) );
  INV_X1 U6417 ( .A(n4925), .ZN(n4926) );
  NAND2_X1 U6418 ( .A1(n4926), .A2(SI_9_), .ZN(n4927) );
  MUX2_X1 U6419 ( .A(n6708), .B(n6709), .S(n6667), .Z(n4929) );
  NAND2_X1 U6420 ( .A1(n4929), .A2(n9579), .ZN(n4932) );
  INV_X1 U6421 ( .A(n4929), .ZN(n4930) );
  NAND2_X1 U6422 ( .A1(n4930), .A2(SI_10_), .ZN(n4931) );
  NAND2_X1 U6423 ( .A1(n5165), .A2(n5164), .ZN(n4933) );
  INV_X1 U6424 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n4934) );
  MUX2_X1 U6425 ( .A(n4934), .B(n6771), .S(n6667), .Z(n4935) );
  XNOR2_X1 U6426 ( .A(n4935), .B(SI_11_), .ZN(n5181) );
  INV_X1 U6427 ( .A(n5181), .ZN(n4938) );
  INV_X1 U6428 ( .A(n4935), .ZN(n4936) );
  NAND2_X1 U6429 ( .A1(n4936), .A2(SI_11_), .ZN(n4937) );
  INV_X1 U6430 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n4939) );
  MUX2_X1 U6431 ( .A(n4939), .B(n6799), .S(n6667), .Z(n4941) );
  INV_X1 U6432 ( .A(SI_12_), .ZN(n4940) );
  NAND2_X1 U6433 ( .A1(n4941), .A2(n4940), .ZN(n4945) );
  INV_X1 U6434 ( .A(n4941), .ZN(n4942) );
  NAND2_X1 U6435 ( .A1(n4942), .A2(SI_12_), .ZN(n4943) );
  NAND2_X1 U6436 ( .A1(n4945), .A2(n4943), .ZN(n5196) );
  INV_X1 U6437 ( .A(n5196), .ZN(n4944) );
  NAND2_X1 U6438 ( .A1(n4946), .A2(n4945), .ZN(n5212) );
  INV_X1 U6439 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n4947) );
  MUX2_X1 U6440 ( .A(n6811), .B(n4947), .S(n6667), .Z(n4948) );
  NAND2_X1 U6441 ( .A1(n4948), .A2(n9562), .ZN(n4951) );
  INV_X1 U6442 ( .A(n4948), .ZN(n4949) );
  NAND2_X1 U6443 ( .A1(n4949), .A2(SI_13_), .ZN(n4950) );
  MUX2_X1 U6444 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6667), .Z(n4953) );
  XNOR2_X1 U6445 ( .A(n4953), .B(n9600), .ZN(n5235) );
  INV_X1 U6446 ( .A(n5235), .ZN(n4952) );
  NAND2_X1 U6447 ( .A1(n4953), .A2(SI_14_), .ZN(n4954) );
  MUX2_X1 U6448 ( .A(n7000), .B(n7001), .S(n6667), .Z(n4955) );
  NAND2_X1 U6449 ( .A1(n4955), .A2(n9521), .ZN(n4958) );
  INV_X1 U6450 ( .A(n4955), .ZN(n4956) );
  NAND2_X1 U6451 ( .A1(n4956), .A2(SI_15_), .ZN(n4957) );
  NAND2_X1 U6452 ( .A1(n4958), .A2(n4957), .ZN(n5258) );
  INV_X1 U6453 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n4959) );
  MUX2_X1 U6454 ( .A(n4959), .B(n7102), .S(n6667), .Z(n4960) );
  NAND2_X1 U6455 ( .A1(n4960), .A2(n9577), .ZN(n4963) );
  INV_X1 U6456 ( .A(n4960), .ZN(n4961) );
  NAND2_X1 U6457 ( .A1(n4961), .A2(SI_16_), .ZN(n4962) );
  MUX2_X1 U6458 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n6667), .Z(n4965) );
  XNOR2_X1 U6459 ( .A(n4965), .B(n4964), .ZN(n5278) );
  NAND2_X1 U6460 ( .A1(n4965), .A2(SI_17_), .ZN(n4966) );
  NAND2_X1 U6461 ( .A1(n4967), .A2(n4966), .ZN(n5300) );
  MUX2_X1 U6462 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6667), .Z(n5301) );
  XNOR2_X1 U6463 ( .A(n5301), .B(SI_18_), .ZN(n5298) );
  XNOR2_X1 U6464 ( .A(n5300), .B(n5298), .ZN(n7252) );
  INV_X1 U6465 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4969) );
  NAND2_X1 U6466 ( .A1(n4974), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4970) );
  NAND2_X1 U6467 ( .A1(n7252), .A2(n4983), .ZN(n4981) );
  OR2_X1 U6468 ( .A1(n5487), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5280) );
  NAND2_X1 U6469 ( .A1(n5282), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4979) );
  XNOR2_X1 U6470 ( .A(n4979), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8583) );
  AOI22_X1 U6471 ( .A1(n4315), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6766), .B2(
        n8583), .ZN(n4980) );
  NAND2_X1 U6472 ( .A1(n8252), .A2(n8286), .ZN(n7339) );
  XNOR2_X1 U6473 ( .A(n8896), .B(n5309), .ZN(n5294) );
  INV_X1 U6474 ( .A(n5294), .ZN(n5296) );
  NAND2_X1 U6475 ( .A1(n7037), .A2(n4983), .ZN(n4987) );
  NAND2_X1 U6476 ( .A1(n5487), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4984) );
  MUX2_X1 U6477 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4984), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n4985) );
  AND2_X1 U6478 ( .A1(n4985), .A2(n5280), .ZN(n8553) );
  AOI22_X1 U6479 ( .A1(n4315), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6766), .B2(
        n8553), .ZN(n4986) );
  INV_X2 U6480 ( .A(n5309), .ZN(n5550) );
  XNOR2_X1 U6481 ( .A(n8905), .B(n5550), .ZN(n5275) );
  INV_X1 U6482 ( .A(n5275), .ZN(n5277) );
  INV_X1 U6483 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8544) );
  NAND2_X1 U6484 ( .A1(n5266), .A2(n8544), .ZN(n4988) );
  NAND2_X1 U6485 ( .A1(n5286), .A2(n4988), .ZN(n7944) );
  INV_X1 U6486 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n4989) );
  OAI22_X1 U6487 ( .A1(n7944), .A2(n5558), .B1(n5528), .B2(n4989), .ZN(n4992)
         );
  INV_X1 U6488 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n4990) );
  INV_X1 U6489 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7945) );
  OAI22_X1 U6490 ( .A1(n5315), .A2(n4990), .B1(n5046), .B2(n7945), .ZN(n4991)
         );
  NAND2_X1 U6491 ( .A1(n8090), .A2(n8506), .ZN(n5276) );
  NAND2_X1 U6492 ( .A1(n4319), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4994) );
  NAND2_X1 U6493 ( .A1(n4320), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4993) );
  AND2_X1 U6494 ( .A1(n4994), .A2(n4993), .ZN(n4997) );
  NAND2_X1 U6495 ( .A1(n8090), .A2(n7025), .ZN(n5013) );
  XNOR2_X1 U6496 ( .A(n4998), .B(n4999), .ZN(n8054) );
  XNOR2_X1 U6497 ( .A(n5013), .B(n5012), .ZN(n7513) );
  INV_X1 U6498 ( .A(SI_0_), .ZN(n5003) );
  INV_X1 U6499 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5002) );
  OAI21_X1 U6500 ( .B1(n6667), .B2(n5003), .A(n5002), .ZN(n5004) );
  AND2_X1 U6501 ( .A1(n5005), .A2(n5004), .ZN(n8950) );
  MUX2_X1 U6502 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8950), .S(n5006), .Z(n7553) );
  OR2_X1 U6503 ( .A1(n5024), .A2(n7553), .ZN(n5011) );
  NAND2_X1 U6504 ( .A1(n4319), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5008) );
  NAND2_X1 U6505 ( .A1(n4320), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5007) );
  NAND2_X1 U6506 ( .A1(n5525), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5010) );
  NAND2_X1 U6507 ( .A1(n8076), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5009) );
  AND2_X1 U6508 ( .A1(n8522), .A2(n7553), .ZN(n7040) );
  NAND2_X1 U6509 ( .A1(n7040), .A2(n8090), .ZN(n7551) );
  AND2_X1 U6510 ( .A1(n5011), .A2(n7551), .ZN(n7514) );
  NAND2_X1 U6511 ( .A1(n7513), .A2(n7514), .ZN(n7512) );
  INV_X1 U6512 ( .A(n5012), .ZN(n5014) );
  NAND2_X1 U6513 ( .A1(n5014), .A2(n5013), .ZN(n5015) );
  NAND2_X1 U6514 ( .A1(n7512), .A2(n5015), .ZN(n8467) );
  INV_X1 U6515 ( .A(n8467), .ZN(n5036) );
  XNOR2_X1 U6516 ( .A(n5017), .B(n5016), .ZN(n6669) );
  NAND2_X1 U6517 ( .A1(n4314), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5023) );
  INV_X1 U6518 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5093) );
  NOR2_X1 U6519 ( .A1(n5000), .A2(n5093), .ZN(n5018) );
  MUX2_X1 U6520 ( .A(n5093), .B(n5018), .S(P2_IR_REG_2__SCAN_IN), .Z(n5021) );
  INV_X1 U6521 ( .A(n5019), .ZN(n5020) );
  NOR2_X1 U6522 ( .A1(n5021), .A2(n5020), .ZN(n6857) );
  OAI211_X2 U6523 ( .C1(n5044), .C2(n6669), .A(n5023), .B(n5022), .ZN(n8823)
         );
  XNOR2_X1 U6524 ( .A(n5024), .B(n8823), .ZN(n5031) );
  NAND2_X1 U6525 ( .A1(n5025), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5027) );
  NAND2_X1 U6526 ( .A1(n4320), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5026) );
  AND2_X1 U6527 ( .A1(n5027), .A2(n5026), .ZN(n5030) );
  NAND2_X1 U6528 ( .A1(n8076), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5029) );
  NAND2_X1 U6529 ( .A1(n5525), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5028) );
  AND3_X2 U6530 ( .A1(n5030), .A2(n5029), .A3(n5028), .ZN(n7242) );
  INV_X1 U6531 ( .A(n7242), .ZN(n8520) );
  AND2_X1 U6532 ( .A1(n8090), .A2(n8520), .ZN(n5032) );
  NAND2_X1 U6533 ( .A1(n5031), .A2(n5032), .ZN(n5037) );
  INV_X1 U6534 ( .A(n5031), .ZN(n7243) );
  INV_X1 U6535 ( .A(n5032), .ZN(n5033) );
  NAND2_X1 U6536 ( .A1(n7243), .A2(n5033), .ZN(n5034) );
  NAND2_X1 U6537 ( .A1(n5037), .A2(n5034), .ZN(n8468) );
  NAND2_X1 U6538 ( .A1(n7244), .A2(n5037), .ZN(n5054) );
  XNOR2_X1 U6539 ( .A(n5038), .B(n5039), .ZN(n6678) );
  NAND2_X1 U6540 ( .A1(n4315), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5043) );
  NAND2_X1 U6541 ( .A1(n5019), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5040) );
  MUX2_X1 U6542 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5040), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5041) );
  AND2_X1 U6543 ( .A1(n5041), .A2(n5055), .ZN(n6858) );
  NAND2_X1 U6544 ( .A1(n6766), .A2(n6858), .ZN(n5042) );
  OAI211_X1 U6545 ( .C1(n5044), .C2(n6678), .A(n5043), .B(n5042), .ZN(n7468)
         );
  NAND2_X1 U6546 ( .A1(n5045), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5050) );
  INV_X1 U6547 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5047) );
  NAND2_X1 U6548 ( .A1(n5525), .A2(n5047), .ZN(n5049) );
  NAND2_X1 U6549 ( .A1(n8076), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5048) );
  AND2_X1 U6550 ( .A1(n8090), .A2(n8519), .ZN(n5051) );
  NAND2_X1 U6551 ( .A1(n7700), .A2(n5051), .ZN(n5067) );
  INV_X1 U6552 ( .A(n5051), .ZN(n5052) );
  AND2_X1 U6553 ( .A1(n5067), .A2(n5053), .ZN(n7245) );
  NAND2_X1 U6554 ( .A1(n5055), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5057) );
  INV_X1 U6555 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5056) );
  XNOR2_X1 U6556 ( .A(n5057), .B(n5056), .ZN(n6905) );
  NAND2_X1 U6557 ( .A1(n5707), .A2(n4983), .ZN(n5061) );
  NAND2_X1 U6558 ( .A1(n4315), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5060) );
  OAI211_X1 U6559 ( .C1(n5006), .C2(n6905), .A(n5061), .B(n5060), .ZN(n7704)
         );
  XNOR2_X1 U6560 ( .A(n5097), .B(n7704), .ZN(n5069) );
  NAND2_X1 U6561 ( .A1(n5045), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5066) );
  NAND2_X1 U6562 ( .A1(n5025), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5065) );
  INV_X1 U6563 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5062) );
  XNOR2_X1 U6564 ( .A(n5062), .B(P2_REG3_REG_3__SCAN_IN), .ZN(n7492) );
  NAND2_X1 U6565 ( .A1(n5525), .A2(n7492), .ZN(n5064) );
  NAND2_X1 U6566 ( .A1(n8076), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5063) );
  NAND4_X1 U6567 ( .A1(n5066), .A2(n5065), .A3(n5064), .A4(n5063), .ZN(n8518)
         );
  NAND2_X1 U6568 ( .A1(n8090), .A2(n8518), .ZN(n5070) );
  XNOR2_X1 U6569 ( .A(n5069), .B(n5070), .ZN(n7699) );
  AND2_X1 U6570 ( .A1(n7699), .A2(n5067), .ZN(n5068) );
  INV_X1 U6571 ( .A(n5069), .ZN(n5071) );
  NAND2_X1 U6572 ( .A1(n5071), .A2(n5070), .ZN(n5072) );
  XNOR2_X1 U6573 ( .A(n5073), .B(n5074), .ZN(n6673) );
  NAND2_X1 U6574 ( .A1(n6673), .A2(n4983), .ZN(n5079) );
  NOR2_X1 U6576 ( .A1(n4871), .A2(n5093), .ZN(n5076) );
  MUX2_X1 U6577 ( .A(n5093), .B(n5076), .S(P2_IR_REG_5__SCAN_IN), .Z(n5077) );
  OR2_X1 U6578 ( .A1(n5077), .A2(n5113), .ZN(n6912) );
  INV_X1 U6579 ( .A(n6912), .ZN(n6919) );
  AOI22_X1 U6580 ( .A1(n8067), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6766), .B2(
        n6919), .ZN(n5078) );
  NAND2_X1 U6581 ( .A1(n5079), .A2(n5078), .ZN(n8451) );
  XNOR2_X1 U6582 ( .A(n5097), .B(n8451), .ZN(n8482) );
  NAND2_X1 U6583 ( .A1(n5045), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5086) );
  NAND2_X1 U6584 ( .A1(n5025), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5085) );
  INV_X1 U6585 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5081) );
  NAND2_X1 U6586 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5080) );
  NAND2_X1 U6587 ( .A1(n5081), .A2(n5080), .ZN(n5082) );
  AND2_X1 U6588 ( .A1(n5098), .A2(n5082), .ZN(n8450) );
  NAND2_X1 U6589 ( .A1(n5525), .A2(n8450), .ZN(n5084) );
  NAND2_X1 U6590 ( .A1(n8076), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5083) );
  NAND4_X1 U6591 ( .A1(n5086), .A2(n5085), .A3(n5084), .A4(n5083), .ZN(n8517)
         );
  AND2_X1 U6592 ( .A1(n8090), .A2(n8517), .ZN(n5087) );
  NAND2_X1 U6593 ( .A1(n8482), .A2(n5087), .ZN(n5104) );
  INV_X1 U6594 ( .A(n8482), .ZN(n5089) );
  INV_X1 U6595 ( .A(n5087), .ZN(n5088) );
  NAND2_X1 U6596 ( .A1(n5089), .A2(n5088), .ZN(n5090) );
  NAND2_X1 U6597 ( .A1(n5104), .A2(n5090), .ZN(n8445) );
  XNOR2_X1 U6598 ( .A(n5091), .B(n5092), .ZN(n6683) );
  NAND2_X1 U6599 ( .A1(n6683), .A2(n4983), .ZN(n5096) );
  OR2_X1 U6600 ( .A1(n5113), .A2(n5093), .ZN(n5094) );
  XNOR2_X1 U6601 ( .A(n5094), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6934) );
  AOI22_X1 U6602 ( .A1(n8067), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6766), .B2(
        n6934), .ZN(n5095) );
  NAND2_X1 U6603 ( .A1(n5096), .A2(n5095), .ZN(n8480) );
  XNOR2_X1 U6604 ( .A(n5097), .B(n8480), .ZN(n5108) );
  NAND2_X1 U6605 ( .A1(n5045), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5103) );
  NAND2_X1 U6606 ( .A1(n5025), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5102) );
  INV_X1 U6607 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9558) );
  NAND2_X1 U6608 ( .A1(n5098), .A2(n9558), .ZN(n5099) );
  AND2_X1 U6609 ( .A1(n5118), .A2(n5099), .ZN(n8478) );
  NAND2_X1 U6610 ( .A1(n5525), .A2(n8478), .ZN(n5101) );
  NAND2_X1 U6611 ( .A1(n8076), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5100) );
  NAND4_X1 U6612 ( .A1(n5103), .A2(n5102), .A3(n5101), .A4(n5100), .ZN(n8516)
         );
  NAND2_X1 U6613 ( .A1(n8090), .A2(n8516), .ZN(n5106) );
  XNOR2_X1 U6614 ( .A(n5108), .B(n5106), .ZN(n8481) );
  AND2_X1 U6615 ( .A1(n8481), .A2(n5104), .ZN(n5105) );
  INV_X1 U6616 ( .A(n5106), .ZN(n5107) );
  OR2_X1 U6617 ( .A1(n5108), .A2(n5107), .ZN(n5109) );
  XNOR2_X1 U6618 ( .A(n5110), .B(n5111), .ZN(n6687) );
  NAND2_X1 U6619 ( .A1(n6687), .A2(n4983), .ZN(n5116) );
  NAND2_X1 U6620 ( .A1(n5113), .A2(n5112), .ZN(n5131) );
  NAND2_X1 U6621 ( .A1(n5131), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5114) );
  XNOR2_X1 U6622 ( .A(n5114), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6954) );
  AOI22_X1 U6623 ( .A1(n8067), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6766), .B2(
        n6954), .ZN(n5115) );
  NAND2_X1 U6624 ( .A1(n5116), .A2(n5115), .ZN(n7626) );
  XNOR2_X1 U6625 ( .A(n7626), .B(n5550), .ZN(n5124) );
  NAND2_X1 U6626 ( .A1(n5045), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5123) );
  NAND2_X1 U6627 ( .A1(n5025), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5122) );
  INV_X1 U6628 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5117) );
  NAND2_X1 U6629 ( .A1(n5118), .A2(n5117), .ZN(n5119) );
  AND2_X1 U6630 ( .A1(n5134), .A2(n5119), .ZN(n7627) );
  NAND2_X1 U6631 ( .A1(n5525), .A2(n7627), .ZN(n5121) );
  NAND2_X1 U6632 ( .A1(n8076), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5120) );
  NAND4_X1 U6633 ( .A1(n5123), .A2(n5122), .A3(n5121), .A4(n5120), .ZN(n8515)
         );
  AND2_X1 U6634 ( .A1(n8090), .A2(n8515), .ZN(n5125) );
  NAND2_X1 U6635 ( .A1(n5124), .A2(n5125), .ZN(n5128) );
  INV_X1 U6636 ( .A(n5124), .ZN(n8414) );
  INV_X1 U6637 ( .A(n5125), .ZN(n5126) );
  NAND2_X1 U6638 ( .A1(n8414), .A2(n5126), .ZN(n5127) );
  NAND2_X1 U6639 ( .A1(n5128), .A2(n5127), .ZN(n7624) );
  NAND2_X1 U6640 ( .A1(n8412), .A2(n5128), .ZN(n5144) );
  NAND2_X1 U6641 ( .A1(n5147), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5132) );
  XNOR2_X1 U6642 ( .A(n5132), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7122) );
  AOI22_X1 U6643 ( .A1(n8072), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6766), .B2(
        n7122), .ZN(n5133) );
  XNOR2_X1 U6644 ( .A(n8419), .B(n5550), .ZN(n8321) );
  NAND2_X1 U6645 ( .A1(n5045), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5139) );
  NAND2_X1 U6646 ( .A1(n5025), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5138) );
  INV_X1 U6647 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9573) );
  NAND2_X1 U6648 ( .A1(n5134), .A2(n9573), .ZN(n5135) );
  AND2_X1 U6649 ( .A1(n5152), .A2(n5135), .ZN(n8420) );
  NAND2_X1 U6650 ( .A1(n5525), .A2(n8420), .ZN(n5137) );
  NAND2_X1 U6651 ( .A1(n8076), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5136) );
  NAND4_X1 U6652 ( .A1(n5139), .A2(n5138), .A3(n5137), .A4(n5136), .ZN(n8514)
         );
  AND2_X1 U6653 ( .A1(n8090), .A2(n8514), .ZN(n5140) );
  NAND2_X1 U6654 ( .A1(n8321), .A2(n5140), .ZN(n5158) );
  INV_X1 U6655 ( .A(n8321), .ZN(n5142) );
  INV_X1 U6656 ( .A(n5140), .ZN(n5141) );
  NAND2_X1 U6657 ( .A1(n5142), .A2(n5141), .ZN(n5143) );
  AND2_X1 U6658 ( .A1(n5158), .A2(n5143), .ZN(n8410) );
  XNOR2_X1 U6659 ( .A(n5145), .B(n5146), .ZN(n6701) );
  NAND2_X1 U6660 ( .A1(n6701), .A2(n4983), .ZN(n5150) );
  NOR2_X1 U6661 ( .A1(n5147), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5167) );
  OR2_X1 U6662 ( .A1(n5167), .A2(n5093), .ZN(n5148) );
  XNOR2_X1 U6663 ( .A(n5148), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7293) );
  AOI22_X1 U6664 ( .A1(n8072), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7293), .B2(
        n6766), .ZN(n5149) );
  NAND2_X1 U6665 ( .A1(n5150), .A2(n5149), .ZN(n8333) );
  XNOR2_X1 U6666 ( .A(n8333), .B(n5550), .ZN(n5160) );
  NAND2_X1 U6667 ( .A1(n5045), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5157) );
  NAND2_X1 U6668 ( .A1(n5025), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5156) );
  NAND2_X1 U6669 ( .A1(n5152), .A2(n5151), .ZN(n5153) );
  AND2_X1 U6670 ( .A1(n5173), .A2(n5153), .ZN(n7540) );
  NAND2_X1 U6671 ( .A1(n5525), .A2(n7540), .ZN(n5155) );
  NAND2_X1 U6672 ( .A1(n8076), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5154) );
  NAND4_X1 U6673 ( .A1(n5157), .A2(n5156), .A3(n5155), .A4(n5154), .ZN(n8513)
         );
  NAND2_X1 U6674 ( .A1(n8090), .A2(n8513), .ZN(n5161) );
  XNOR2_X1 U6675 ( .A(n5160), .B(n5161), .ZN(n8323) );
  AND2_X1 U6676 ( .A1(n8323), .A2(n5158), .ZN(n5159) );
  NAND2_X1 U6677 ( .A1(n8416), .A2(n5159), .ZN(n8336) );
  INV_X1 U6678 ( .A(n5160), .ZN(n5162) );
  NAND2_X1 U6679 ( .A1(n5162), .A2(n5161), .ZN(n5163) );
  XNOR2_X1 U6680 ( .A(n5165), .B(n5164), .ZN(n5824) );
  NAND2_X1 U6681 ( .A1(n5824), .A2(n4983), .ZN(n5172) );
  NAND2_X1 U6682 ( .A1(n5167), .A2(n5166), .ZN(n5198) );
  NAND2_X1 U6683 ( .A1(n5198), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5169) );
  NAND2_X1 U6684 ( .A1(n5169), .A2(n5168), .ZN(n5183) );
  OR2_X1 U6685 ( .A1(n5169), .A2(n5168), .ZN(n5170) );
  AOI22_X1 U6686 ( .A1(n7649), .A2(n6766), .B1(n8067), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n5171) );
  XNOR2_X1 U6687 ( .A(n7676), .B(n5550), .ZN(n7361) );
  NAND2_X1 U6688 ( .A1(n5045), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5178) );
  NAND2_X1 U6689 ( .A1(n5025), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5177) );
  NAND2_X1 U6690 ( .A1(n5173), .A2(n9586), .ZN(n5174) );
  AND2_X1 U6691 ( .A1(n5188), .A2(n5174), .ZN(n7567) );
  NAND2_X1 U6692 ( .A1(n5525), .A2(n7567), .ZN(n5176) );
  NAND2_X1 U6693 ( .A1(n8076), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5175) );
  NAND4_X1 U6694 ( .A1(n5178), .A2(n5177), .A3(n5176), .A4(n5175), .ZN(n8512)
         );
  AND2_X1 U6695 ( .A1(n8090), .A2(n8512), .ZN(n5179) );
  NAND2_X1 U6696 ( .A1(n7361), .A2(n5179), .ZN(n5230) );
  NAND2_X1 U6697 ( .A1(n5230), .A2(n5180), .ZN(n7573) );
  NAND2_X1 U6698 ( .A1(n6706), .A2(n4983), .ZN(n5186) );
  NAND2_X1 U6699 ( .A1(n5183), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5184) );
  XNOR2_X1 U6700 ( .A(n5184), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7799) );
  AOI22_X1 U6701 ( .A1(n7799), .A2(n6766), .B1(n8072), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n5185) );
  XNOR2_X1 U6702 ( .A(n7367), .B(n5550), .ZN(n8299) );
  NAND2_X1 U6703 ( .A1(n5045), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5193) );
  NAND2_X1 U6704 ( .A1(n5025), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5192) );
  INV_X1 U6705 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5187) );
  NAND2_X1 U6706 ( .A1(n5188), .A2(n5187), .ZN(n5189) );
  AND2_X1 U6707 ( .A1(n5202), .A2(n5189), .ZN(n7368) );
  NAND2_X1 U6708 ( .A1(n5525), .A2(n7368), .ZN(n5191) );
  NAND2_X1 U6709 ( .A1(n8076), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5190) );
  NAND4_X1 U6710 ( .A1(n5193), .A2(n5192), .A3(n5191), .A4(n5190), .ZN(n8511)
         );
  AND2_X1 U6711 ( .A1(n8090), .A2(n8511), .ZN(n5194) );
  NAND2_X1 U6712 ( .A1(n8299), .A2(n5194), .ZN(n5229) );
  NAND2_X1 U6713 ( .A1(n5229), .A2(n5195), .ZN(n7360) );
  OR2_X1 U6714 ( .A1(n7573), .A2(n7360), .ZN(n7363) );
  XNOR2_X1 U6715 ( .A(n5197), .B(n5196), .ZN(n5859) );
  NAND2_X1 U6716 ( .A1(n5859), .A2(n4983), .ZN(n5201) );
  NAND2_X1 U6717 ( .A1(n5213), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5199) );
  XNOR2_X1 U6718 ( .A(n5199), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8527) );
  AOI22_X1 U6719 ( .A1(n8527), .A2(n6766), .B1(n8067), .B2(
        P1_DATAO_REG_12__SCAN_IN), .ZN(n5200) );
  INV_X1 U6720 ( .A(n5228), .ZN(n5208) );
  NAND2_X1 U6721 ( .A1(n5045), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5207) );
  NAND2_X1 U6722 ( .A1(n5025), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5206) );
  INV_X1 U6723 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9596) );
  NAND2_X1 U6724 ( .A1(n5202), .A2(n9596), .ZN(n5203) );
  AND2_X1 U6725 ( .A1(n5216), .A2(n5203), .ZN(n8307) );
  NAND2_X1 U6726 ( .A1(n5525), .A2(n8307), .ZN(n5205) );
  NAND2_X1 U6727 ( .A1(n8076), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5204) );
  NAND4_X1 U6728 ( .A1(n5207), .A2(n5206), .A3(n5205), .A4(n5204), .ZN(n8510)
         );
  NAND2_X1 U6729 ( .A1(n8090), .A2(n8510), .ZN(n5227) );
  NAND2_X1 U6730 ( .A1(n5208), .A2(n5227), .ZN(n5209) );
  INV_X1 U6731 ( .A(n5209), .ZN(n5232) );
  XNOR2_X1 U6732 ( .A(n5212), .B(n5211), .ZN(n5883) );
  NAND2_X1 U6733 ( .A1(n5883), .A2(n4983), .ZN(n5215) );
  OAI21_X1 U6734 ( .B1(n5213), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5238) );
  XNOR2_X1 U6735 ( .A(n5238), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7874) );
  AOI22_X1 U6736 ( .A1(n7874), .A2(n6766), .B1(n8067), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n5214) );
  XNOR2_X1 U6737 ( .A(n7504), .B(n5550), .ZN(n7580) );
  NAND2_X1 U6738 ( .A1(n5045), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5221) );
  NAND2_X1 U6739 ( .A1(n5025), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5220) );
  NAND2_X1 U6740 ( .A1(n5216), .A2(n7803), .ZN(n5217) );
  AND2_X1 U6741 ( .A1(n5246), .A2(n5217), .ZN(n7763) );
  NAND2_X1 U6742 ( .A1(n5525), .A2(n7763), .ZN(n5219) );
  NAND2_X1 U6743 ( .A1(n8076), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5218) );
  NAND4_X1 U6744 ( .A1(n5221), .A2(n5220), .A3(n5219), .A4(n5218), .ZN(n8509)
         );
  AND2_X1 U6745 ( .A1(n8090), .A2(n8509), .ZN(n5222) );
  NAND2_X1 U6746 ( .A1(n7580), .A2(n5222), .ZN(n5252) );
  OR2_X1 U6747 ( .A1(n7580), .A2(n5222), .ZN(n5223) );
  NAND2_X1 U6748 ( .A1(n5252), .A2(n5223), .ZN(n7503) );
  INV_X1 U6749 ( .A(n7503), .ZN(n5224) );
  NAND2_X1 U6750 ( .A1(n5225), .A2(n5224), .ZN(n5226) );
  NOR2_X1 U6751 ( .A1(n7359), .A2(n5226), .ZN(n5234) );
  XNOR2_X1 U6752 ( .A(n5228), .B(n5227), .ZN(n8315) );
  AND2_X1 U6753 ( .A1(n8315), .A2(n5229), .ZN(n5231) );
  OR2_X1 U6754 ( .A1(n7360), .A2(n5230), .ZN(n7364) );
  AND2_X1 U6755 ( .A1(n5231), .A2(n7364), .ZN(n8305) );
  NOR2_X1 U6756 ( .A1(n7503), .A2(n7500), .ZN(n5233) );
  NOR2_X1 U6757 ( .A1(n5234), .A2(n5233), .ZN(n7501) );
  NAND2_X1 U6758 ( .A1(n6818), .A2(n4983), .ZN(n5244) );
  NAND2_X1 U6759 ( .A1(n5238), .A2(n5237), .ZN(n5239) );
  NAND2_X1 U6760 ( .A1(n5239), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5241) );
  NAND2_X1 U6761 ( .A1(n5241), .A2(n5240), .ZN(n5260) );
  OR2_X1 U6762 ( .A1(n5241), .A2(n5240), .ZN(n5242) );
  AOI22_X1 U6763 ( .A1(n8003), .A2(n6766), .B1(n8067), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5243) );
  NAND2_X1 U6764 ( .A1(n5045), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5251) );
  NAND2_X1 U6765 ( .A1(n5025), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5250) );
  INV_X1 U6766 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5245) );
  NAND2_X1 U6767 ( .A1(n5246), .A2(n5245), .ZN(n5247) );
  AND2_X1 U6768 ( .A1(n5264), .A2(n5247), .ZN(n7777) );
  NAND2_X1 U6769 ( .A1(n5525), .A2(n7777), .ZN(n5249) );
  NAND2_X1 U6770 ( .A1(n8076), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5248) );
  NAND4_X1 U6771 ( .A1(n5251), .A2(n5250), .A3(n5249), .A4(n5248), .ZN(n8508)
         );
  NAND2_X1 U6772 ( .A1(n8090), .A2(n8508), .ZN(n5255) );
  XNOR2_X1 U6773 ( .A(n5254), .B(n5255), .ZN(n7592) );
  AND2_X1 U6774 ( .A1(n7592), .A2(n5252), .ZN(n5253) );
  INV_X1 U6775 ( .A(n5254), .ZN(n5256) );
  NAND2_X1 U6776 ( .A1(n5256), .A2(n5255), .ZN(n5257) );
  XNOR2_X1 U6777 ( .A(n5259), .B(n5258), .ZN(n6999) );
  NAND2_X1 U6778 ( .A1(n6999), .A2(n4983), .ZN(n5263) );
  NAND2_X1 U6779 ( .A1(n5260), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5261) );
  XNOR2_X1 U6780 ( .A(n5261), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8547) );
  AOI22_X1 U6781 ( .A1(n8547), .A2(n6766), .B1(n8072), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5262) );
  XNOR2_X1 U6782 ( .A(n8910), .B(n5550), .ZN(n5272) );
  NAND2_X1 U6783 ( .A1(n5045), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5270) );
  NAND2_X1 U6784 ( .A1(n5025), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5269) );
  NAND2_X1 U6785 ( .A1(n5264), .A2(n7661), .ZN(n5265) );
  AND2_X1 U6786 ( .A1(n5266), .A2(n5265), .ZN(n7901) );
  NAND2_X1 U6787 ( .A1(n5525), .A2(n7901), .ZN(n5268) );
  NAND2_X1 U6788 ( .A1(n8076), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5267) );
  NAND4_X1 U6789 ( .A1(n5270), .A2(n5269), .A3(n5268), .A4(n5267), .ZN(n8507)
         );
  AND2_X1 U6790 ( .A1(n8507), .A2(n8090), .ZN(n5271) );
  XOR2_X1 U6791 ( .A(n5276), .B(n5275), .Z(n7811) );
  XNOR2_X1 U6792 ( .A(n5279), .B(n5278), .ZN(n7136) );
  NAND2_X1 U6793 ( .A1(n7136), .A2(n4983), .ZN(n5285) );
  NAND2_X1 U6794 ( .A1(n5280), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5281) );
  MUX2_X1 U6795 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5281), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n5283) );
  AOI22_X1 U6796 ( .A1(n8072), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6766), .B2(
        n8578), .ZN(n5284) );
  XNOR2_X1 U6797 ( .A(n8901), .B(n5309), .ZN(n8350) );
  NAND2_X1 U6798 ( .A1(n5286), .A2(n9604), .ZN(n5287) );
  NAND2_X1 U6799 ( .A1(n5288), .A2(n5287), .ZN(n8816) );
  AOI22_X1 U6800 ( .A1(n5045), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n5025), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n5290) );
  NAND2_X1 U6801 ( .A1(n8076), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5289) );
  OAI211_X1 U6802 ( .C1(n8816), .C2(n5558), .A(n5290), .B(n5289), .ZN(n8789)
         );
  NAND2_X1 U6803 ( .A1(n8789), .A2(n8090), .ZN(n5291) );
  NOR2_X1 U6804 ( .A1(n8350), .A2(n5291), .ZN(n5292) );
  AOI21_X1 U6805 ( .B1(n8350), .B2(n5291), .A(n5292), .ZN(n7884) );
  INV_X1 U6806 ( .A(n5292), .ZN(n5295) );
  XNOR2_X1 U6807 ( .A(n5294), .B(n5293), .ZN(n8347) );
  INV_X1 U6808 ( .A(n5298), .ZN(n5299) );
  NAND2_X1 U6809 ( .A1(n5301), .A2(SI_18_), .ZN(n5302) );
  MUX2_X1 U6810 ( .A(n7306), .B(n7304), .S(n6667), .Z(n5304) );
  INV_X1 U6811 ( .A(SI_19_), .ZN(n5303) );
  NAND2_X1 U6812 ( .A1(n5304), .A2(n5303), .ZN(n5324) );
  INV_X1 U6813 ( .A(n5304), .ZN(n5305) );
  NAND2_X1 U6814 ( .A1(n5305), .A2(SI_19_), .ZN(n5306) );
  NAND2_X1 U6815 ( .A1(n5324), .A2(n5306), .ZN(n5325) );
  XNOR2_X1 U6816 ( .A(n5326), .B(n5325), .ZN(n7303) );
  NAND2_X1 U6817 ( .A1(n7303), .A2(n4983), .ZN(n5308) );
  AOI22_X1 U6818 ( .A1(n8657), .A2(n6766), .B1(n4315), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n5307) );
  XNOR2_X1 U6819 ( .A(n8892), .B(n5309), .ZN(n5323) );
  INV_X1 U6820 ( .A(n5323), .ZN(n5321) );
  INV_X1 U6821 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5310) );
  NAND2_X1 U6822 ( .A1(n5311), .A2(n5310), .ZN(n5312) );
  AND2_X1 U6823 ( .A1(n5333), .A2(n5312), .ZN(n8765) );
  NAND2_X1 U6824 ( .A1(n8765), .A2(n5525), .ZN(n5319) );
  INV_X1 U6825 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n5316) );
  NAND2_X1 U6826 ( .A1(n4319), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5314) );
  NAND2_X1 U6827 ( .A1(n8076), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5313) );
  OAI211_X1 U6828 ( .C1(n5316), .C2(n5315), .A(n5314), .B(n5313), .ZN(n5317)
         );
  INV_X1 U6829 ( .A(n5317), .ZN(n5318) );
  NAND2_X1 U6830 ( .A1(n5319), .A2(n5318), .ZN(n8791) );
  NAND2_X1 U6831 ( .A1(n8791), .A2(n8090), .ZN(n5322) );
  INV_X1 U6832 ( .A(n5322), .ZN(n5320) );
  NAND2_X1 U6833 ( .A1(n5321), .A2(n5320), .ZN(n7968) );
  MUX2_X1 U6834 ( .A(n7511), .B(n7547), .S(n6667), .Z(n5327) );
  NAND2_X1 U6835 ( .A1(n5327), .A2(n9529), .ZN(n5354) );
  INV_X1 U6836 ( .A(n5327), .ZN(n5328) );
  NAND2_X1 U6837 ( .A1(n5328), .A2(SI_20_), .ZN(n5329) );
  XNOR2_X1 U6838 ( .A(n5353), .B(n5352), .ZN(n7510) );
  NAND2_X1 U6839 ( .A1(n7510), .A2(n4983), .ZN(n5331) );
  NAND2_X1 U6840 ( .A1(n8072), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5330) );
  XNOR2_X1 U6841 ( .A(n8886), .B(n5550), .ZN(n5342) );
  INV_X1 U6842 ( .A(n5333), .ZN(n5332) );
  NAND2_X1 U6843 ( .A1(n5332), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5344) );
  INV_X1 U6844 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8033) );
  NAND2_X1 U6845 ( .A1(n5333), .A2(n8033), .ZN(n5334) );
  NAND2_X1 U6846 ( .A1(n5344), .A2(n5334), .ZN(n8754) );
  OR2_X1 U6847 ( .A1(n8754), .A2(n5558), .ZN(n5340) );
  INV_X1 U6848 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n5337) );
  NAND2_X1 U6849 ( .A1(n5025), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5336) );
  NAND2_X1 U6850 ( .A1(n5045), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5335) );
  OAI211_X1 U6851 ( .C1(n5337), .C2(n5528), .A(n5336), .B(n5335), .ZN(n5338)
         );
  INV_X1 U6852 ( .A(n5338), .ZN(n5339) );
  NAND2_X1 U6853 ( .A1(n5340), .A2(n5339), .ZN(n8772) );
  NAND2_X1 U6854 ( .A1(n8772), .A2(n8090), .ZN(n5341) );
  INV_X1 U6855 ( .A(n5341), .ZN(n5343) );
  NAND2_X1 U6856 ( .A1(n5344), .A2(n9564), .ZN(n5345) );
  NAND2_X1 U6857 ( .A1(n5374), .A2(n5345), .ZN(n8733) );
  OR2_X1 U6858 ( .A1(n8733), .A2(n5558), .ZN(n5351) );
  INV_X1 U6859 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n5348) );
  NAND2_X1 U6860 ( .A1(n5025), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5347) );
  NAND2_X1 U6861 ( .A1(n5045), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5346) );
  OAI211_X1 U6862 ( .C1(n5348), .C2(n5528), .A(n5347), .B(n5346), .ZN(n5349)
         );
  INV_X1 U6863 ( .A(n5349), .ZN(n5350) );
  NAND2_X1 U6864 ( .A1(n5351), .A2(n5350), .ZN(n8749) );
  NAND2_X1 U6865 ( .A1(n8749), .A2(n8090), .ZN(n5359) );
  NAND2_X1 U6866 ( .A1(n5355), .A2(n5354), .ZN(n5363) );
  MUX2_X1 U6867 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n6667), .Z(n5364) );
  XNOR2_X1 U6868 ( .A(n5364), .B(n9559), .ZN(n5361) );
  XNOR2_X1 U6869 ( .A(n5363), .B(n5361), .ZN(n7577) );
  NAND2_X1 U6870 ( .A1(n7577), .A2(n4983), .ZN(n5357) );
  NAND2_X1 U6871 ( .A1(n8067), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5356) );
  INV_X1 U6872 ( .A(n5358), .ZN(n5360) );
  INV_X1 U6873 ( .A(n5361), .ZN(n5362) );
  NAND2_X1 U6874 ( .A1(n5364), .A2(SI_21_), .ZN(n5365) );
  MUX2_X1 U6875 ( .A(n8401), .B(n7713), .S(n6667), .Z(n5368) );
  INV_X1 U6876 ( .A(SI_22_), .ZN(n5367) );
  NAND2_X1 U6877 ( .A1(n5368), .A2(n5367), .ZN(n5386) );
  INV_X1 U6878 ( .A(n5368), .ZN(n5369) );
  NAND2_X1 U6879 ( .A1(n5369), .A2(SI_22_), .ZN(n5370) );
  NAND2_X1 U6880 ( .A1(n5386), .A2(n5370), .ZN(n5384) );
  XNOR2_X1 U6881 ( .A(n5385), .B(n5384), .ZN(n7712) );
  NAND2_X1 U6882 ( .A1(n7712), .A2(n4983), .ZN(n5372) );
  NAND2_X1 U6883 ( .A1(n4315), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5371) );
  XNOR2_X1 U6884 ( .A(n8874), .B(n5550), .ZN(n5381) );
  XNOR2_X1 U6885 ( .A(n5382), .B(n5373), .ZN(n8395) );
  NAND2_X1 U6886 ( .A1(n5374), .A2(n9541), .ZN(n5375) );
  INV_X1 U6887 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n5378) );
  NAND2_X1 U6888 ( .A1(n5025), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5377) );
  NAND2_X1 U6889 ( .A1(n5045), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5376) );
  OAI211_X1 U6890 ( .C1(n5378), .C2(n5528), .A(n5377), .B(n5376), .ZN(n5379)
         );
  INV_X1 U6891 ( .A(n8090), .ZN(n5514) );
  OR2_X1 U6892 ( .A1(n8427), .A2(n5514), .ZN(n5380) );
  NAND2_X1 U6893 ( .A1(n8395), .A2(n5380), .ZN(n8399) );
  OR2_X1 U6894 ( .A1(n5382), .A2(n5381), .ZN(n5383) );
  NAND2_X2 U6895 ( .A1(n8399), .A2(n5383), .ZN(n5404) );
  INV_X1 U6896 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5388) );
  INV_X1 U6897 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5387) );
  MUX2_X1 U6898 ( .A(n5388), .B(n5387), .S(n6667), .Z(n5390) );
  INV_X1 U6899 ( .A(SI_23_), .ZN(n5389) );
  NAND2_X1 U6900 ( .A1(n5390), .A2(n5389), .ZN(n5408) );
  INV_X1 U6901 ( .A(n5390), .ZN(n5391) );
  NAND2_X1 U6902 ( .A1(n5391), .A2(SI_23_), .ZN(n5392) );
  XNOR2_X1 U6903 ( .A(n5407), .B(n5406), .ZN(n7816) );
  NAND2_X1 U6904 ( .A1(n7816), .A2(n4983), .ZN(n5394) );
  NAND2_X1 U6905 ( .A1(n4315), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5393) );
  XNOR2_X2 U6906 ( .A(n5404), .B(n4382), .ZN(n8403) );
  INV_X1 U6907 ( .A(n5396), .ZN(n5395) );
  NAND2_X1 U6908 ( .A1(n5395), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5413) );
  INV_X1 U6909 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9561) );
  NAND2_X1 U6910 ( .A1(n5396), .A2(n9561), .ZN(n5397) );
  NAND2_X1 U6911 ( .A1(n5413), .A2(n5397), .ZN(n8702) );
  OR2_X1 U6912 ( .A1(n8702), .A2(n5558), .ZN(n5403) );
  INV_X1 U6913 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n5400) );
  NAND2_X1 U6914 ( .A1(n5025), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5399) );
  NAND2_X1 U6915 ( .A1(n5045), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5398) );
  OAI211_X1 U6916 ( .C1(n5528), .C2(n5400), .A(n5399), .B(n5398), .ZN(n5401)
         );
  INV_X1 U6917 ( .A(n5401), .ZN(n5402) );
  NAND2_X1 U6918 ( .A1(n5403), .A2(n5402), .ZN(n8505) );
  NAND2_X1 U6919 ( .A1(n8505), .A2(n8090), .ZN(n8402) );
  MUX2_X1 U6920 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n6667), .Z(n5424) );
  INV_X1 U6921 ( .A(SI_24_), .ZN(n9598) );
  XNOR2_X1 U6922 ( .A(n5424), .B(n9598), .ZN(n5423) );
  XNOR2_X1 U6923 ( .A(n5422), .B(n5423), .ZN(n7890) );
  NAND2_X1 U6924 ( .A1(n7890), .A2(n4983), .ZN(n5411) );
  NAND2_X1 U6925 ( .A1(n8072), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5410) );
  XNOR2_X1 U6926 ( .A(n8864), .B(n5550), .ZN(n5421) );
  INV_X1 U6927 ( .A(n5413), .ZN(n5412) );
  NAND2_X1 U6928 ( .A1(n5412), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5432) );
  INV_X1 U6929 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9565) );
  NAND2_X1 U6930 ( .A1(n5413), .A2(n9565), .ZN(n5414) );
  NAND2_X1 U6931 ( .A1(n5432), .A2(n5414), .ZN(n8684) );
  OR2_X1 U6932 ( .A1(n8684), .A2(n5558), .ZN(n5420) );
  INV_X1 U6933 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n5417) );
  NAND2_X1 U6934 ( .A1(n5025), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5416) );
  NAND2_X1 U6935 ( .A1(n5045), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5415) );
  OAI211_X1 U6936 ( .C1(n5528), .C2(n5417), .A(n5416), .B(n5415), .ZN(n5418)
         );
  INV_X1 U6937 ( .A(n5418), .ZN(n5419) );
  NAND2_X1 U6938 ( .A1(n5420), .A2(n5419), .ZN(n8710) );
  NAND2_X1 U6939 ( .A1(n8710), .A2(n8090), .ZN(n8455) );
  NAND2_X1 U6940 ( .A1(n5424), .A2(SI_24_), .ZN(n5425) );
  INV_X1 U6941 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7934) );
  INV_X1 U6942 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7933) );
  MUX2_X1 U6943 ( .A(n7934), .B(n7933), .S(n6667), .Z(n5427) );
  INV_X1 U6944 ( .A(SI_25_), .ZN(n5426) );
  NAND2_X1 U6945 ( .A1(n5427), .A2(n5426), .ZN(n5440) );
  INV_X1 U6946 ( .A(n5427), .ZN(n5428) );
  NAND2_X1 U6947 ( .A1(n5428), .A2(SI_25_), .ZN(n5429) );
  NAND2_X1 U6948 ( .A1(n5440), .A2(n5429), .ZN(n5441) );
  NAND2_X1 U6949 ( .A1(n7932), .A2(n4983), .ZN(n5431) );
  NAND2_X1 U6950 ( .A1(n8072), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5430) );
  XNOR2_X1 U6951 ( .A(n8860), .B(n5550), .ZN(n8434) );
  NAND2_X1 U6952 ( .A1(n5432), .A2(n8437), .ZN(n5433) );
  AND2_X1 U6953 ( .A1(n5449), .A2(n5433), .ZN(n8668) );
  NAND2_X1 U6954 ( .A1(n8668), .A2(n5525), .ZN(n5439) );
  INV_X1 U6955 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U6956 ( .A1(n5045), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5435) );
  NAND2_X1 U6957 ( .A1(n4319), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5434) );
  OAI211_X1 U6958 ( .C1(n5436), .C2(n5528), .A(n5435), .B(n5434), .ZN(n5437)
         );
  INV_X1 U6959 ( .A(n5437), .ZN(n5438) );
  NOR2_X1 U6960 ( .A1(n8693), .A2(n5514), .ZN(n8435) );
  INV_X1 U6961 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8029) );
  MUX2_X1 U6962 ( .A(n8029), .B(n8014), .S(n6667), .Z(n5443) );
  NAND2_X1 U6963 ( .A1(n5443), .A2(n9601), .ZN(n5459) );
  INV_X1 U6964 ( .A(n5443), .ZN(n5444) );
  NAND2_X1 U6965 ( .A1(n5444), .A2(SI_26_), .ZN(n5445) );
  XNOR2_X1 U6966 ( .A(n5458), .B(n5457), .ZN(n8013) );
  NAND2_X1 U6967 ( .A1(n8013), .A2(n4983), .ZN(n5447) );
  NAND2_X1 U6968 ( .A1(n4315), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5446) );
  XNOR2_X1 U6969 ( .A(n8851), .B(n5550), .ZN(n5513) );
  INV_X1 U6970 ( .A(n5449), .ZN(n5448) );
  INV_X1 U6971 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9539) );
  NAND2_X1 U6972 ( .A1(n5449), .A2(n9539), .ZN(n5450) );
  NAND2_X1 U6973 ( .A1(n5523), .A2(n5450), .ZN(n8656) );
  INV_X1 U6974 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8919) );
  NAND2_X1 U6975 ( .A1(n5045), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5452) );
  NAND2_X1 U6976 ( .A1(n5025), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5451) );
  OAI211_X1 U6977 ( .C1(n8919), .C2(n5528), .A(n5452), .B(n5451), .ZN(n5453)
         );
  INV_X1 U6978 ( .A(n5453), .ZN(n5454) );
  AND2_X1 U6979 ( .A1(n8673), .A2(n8090), .ZN(n5456) );
  NAND2_X1 U6980 ( .A1(n5513), .A2(n5456), .ZN(n5516) );
  OAI21_X1 U6981 ( .B1(n5513), .B2(n5456), .A(n5516), .ZN(n8491) );
  NAND2_X1 U6982 ( .A1(n5458), .A2(n5457), .ZN(n5460) );
  INV_X1 U6983 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5461) );
  MUX2_X1 U6984 ( .A(n8948), .B(n5461), .S(n6667), .Z(n5462) );
  NAND2_X1 U6985 ( .A1(n5462), .A2(n9518), .ZN(n5546) );
  INV_X1 U6986 ( .A(n5462), .ZN(n5463) );
  NAND2_X1 U6987 ( .A1(n5463), .A2(SI_27_), .ZN(n5464) );
  NAND2_X1 U6988 ( .A1(n6158), .A2(n4983), .ZN(n5466) );
  NAND2_X1 U6989 ( .A1(n4315), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5465) );
  XNOR2_X1 U6990 ( .A(n8378), .B(n5550), .ZN(n5473) );
  XNOR2_X1 U6991 ( .A(n5523), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8636) );
  NAND2_X1 U6992 ( .A1(n8636), .A2(n5525), .ZN(n5472) );
  INV_X1 U6993 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n5469) );
  NAND2_X1 U6994 ( .A1(n5045), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5468) );
  NAND2_X1 U6995 ( .A1(n5025), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5467) );
  OAI211_X1 U6996 ( .C1(n5469), .C2(n5528), .A(n5468), .B(n5467), .ZN(n5470)
         );
  INV_X1 U6997 ( .A(n5470), .ZN(n5471) );
  AND2_X1 U6998 ( .A1(n8649), .A2(n8090), .ZN(n5474) );
  NAND2_X1 U6999 ( .A1(n5473), .A2(n5474), .ZN(n5563) );
  INV_X1 U7000 ( .A(n5473), .ZN(n5476) );
  INV_X1 U7001 ( .A(n5474), .ZN(n5475) );
  NAND2_X1 U7002 ( .A1(n5476), .A2(n5475), .ZN(n5477) );
  NOR4_X1 U7003 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n5481) );
  NOR4_X1 U7004 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n5480) );
  NOR4_X1 U7005 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5479) );
  NOR4_X1 U7006 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5478) );
  NAND4_X1 U7007 ( .A1(n5481), .A2(n5480), .A3(n5479), .A4(n5478), .ZN(n5503)
         );
  NOR2_X1 U7008 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n5485) );
  NOR4_X1 U7009 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n5484) );
  NOR4_X1 U7010 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5483) );
  NOR4_X1 U7011 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n5482) );
  NAND4_X1 U7012 ( .A1(n5485), .A2(n5484), .A3(n5483), .A4(n5482), .ZN(n5502)
         );
  OAI21_X1 U7013 ( .B1(n5487), .B2(n5486), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5488) );
  MUX2_X1 U7014 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5488), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n5489) );
  NAND2_X1 U7015 ( .A1(n5491), .A2(n5490), .ZN(n5492) );
  NAND2_X1 U7016 ( .A1(n5509), .A2(n5508), .ZN(n5493) );
  INV_X1 U7017 ( .A(P2_B_REG_SCAN_IN), .ZN(n8384) );
  XOR2_X1 U7018 ( .A(n7915), .B(n8384), .Z(n5496) );
  NAND2_X1 U7019 ( .A1(n7936), .A2(n5496), .ZN(n5501) );
  NAND2_X1 U7020 ( .A1(n4393), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5498) );
  MUX2_X1 U7021 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5498), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5499) );
  INV_X1 U7022 ( .A(n8030), .ZN(n5500) );
  OAI21_X1 U7023 ( .B1(n5503), .B2(n5502), .A(n10026), .ZN(n7021) );
  AND2_X1 U7024 ( .A1(n7915), .A2(n8030), .ZN(n10029) );
  INV_X1 U7025 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10028) );
  AND2_X1 U7026 ( .A1(n10026), .A2(n10028), .ZN(n5504) );
  NAND2_X1 U7027 ( .A1(n10026), .A2(n10031), .ZN(n5506) );
  AND2_X1 U7028 ( .A1(n7936), .A2(n8030), .ZN(n10032) );
  NOR2_X1 U7029 ( .A1(n7073), .A2(n7335), .ZN(n5507) );
  NAND2_X1 U7030 ( .A1(n7021), .A2(n5507), .ZN(n5535) );
  NAND2_X1 U7031 ( .A1(n5511), .A2(n8286), .ZN(n6768) );
  AND2_X1 U7032 ( .A1(n10062), .A2(n6768), .ZN(n5512) );
  INV_X1 U7033 ( .A(n5513), .ZN(n5515) );
  INV_X1 U7034 ( .A(n8673), .ZN(n8440) );
  NAND2_X1 U7035 ( .A1(n5518), .A2(n5517), .ZN(n5568) );
  INV_X1 U7036 ( .A(n5533), .ZN(n5520) );
  OR2_X1 U7037 ( .A1(n5510), .A2(n8252), .ZN(n7341) );
  INV_X1 U7038 ( .A(n8461), .ZN(n7507) );
  NAND2_X1 U7039 ( .A1(n8378), .A2(n8500), .ZN(n5542) );
  INV_X1 U7040 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9533) );
  INV_X1 U7041 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5521) );
  OAI21_X1 U7042 ( .B1(n5523), .B2(n9533), .A(n5521), .ZN(n5524) );
  NAND2_X1 U7043 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n5522) );
  NAND2_X1 U7044 ( .A1(n8616), .A2(n5525), .ZN(n5532) );
  INV_X1 U7045 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n5529) );
  NAND2_X1 U7046 ( .A1(n5045), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5527) );
  NAND2_X1 U7047 ( .A1(n5025), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5526) );
  OAI211_X1 U7048 ( .C1(n5529), .C2(n5528), .A(n5527), .B(n5526), .ZN(n5530)
         );
  INV_X1 U7049 ( .A(n5530), .ZN(n5531) );
  INV_X1 U7050 ( .A(n5534), .ZN(n6830) );
  AOI22_X1 U7051 ( .A1(n8632), .A2(n8465), .B1(n8464), .B2(n8673), .ZN(n5540)
         );
  NAND2_X1 U7052 ( .A1(n5535), .A2(n7023), .ZN(n5538) );
  OR2_X1 U7053 ( .A1(n6768), .A2(n5536), .ZN(n7070) );
  AND3_X1 U7054 ( .A1(n6833), .A2(n6765), .A3(n7070), .ZN(n5537) );
  NAND2_X1 U7055 ( .A1(n5538), .A2(n5537), .ZN(n7516) );
  AOI22_X1 U7056 ( .A1(n8636), .A2(n8479), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n5539) );
  NAND2_X1 U7057 ( .A1(n5543), .A2(n4836), .ZN(P2_U3216) );
  NAND2_X1 U7058 ( .A1(n5545), .A2(n5544), .ZN(n5547) );
  MUX2_X1 U7059 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n6667), .Z(n6291) );
  INV_X1 U7060 ( .A(SI_28_), .ZN(n6292) );
  XNOR2_X1 U7061 ( .A(n6291), .B(n6292), .ZN(n6289) );
  NAND2_X1 U7062 ( .A1(n8942), .A2(n4983), .ZN(n5549) );
  NAND2_X1 U7063 ( .A1(n8072), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5548) );
  NAND2_X1 U7064 ( .A1(n8632), .A2(n8090), .ZN(n5551) );
  XNOR2_X1 U7065 ( .A(n5551), .B(n5550), .ZN(n5552) );
  XNOR2_X1 U7066 ( .A(n8840), .B(n5552), .ZN(n5564) );
  INV_X1 U7067 ( .A(n5564), .ZN(n5553) );
  NAND2_X1 U7068 ( .A1(n5553), .A2(n8474), .ZN(n5567) );
  NAND2_X1 U7069 ( .A1(n5045), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5556) );
  NAND2_X1 U7070 ( .A1(n4319), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5555) );
  NAND2_X1 U7071 ( .A1(n8076), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5554) );
  AND3_X1 U7072 ( .A1(n5556), .A2(n5555), .A3(n5554), .ZN(n5557) );
  OAI21_X1 U7073 ( .B1(n8379), .B2(n5558), .A(n5557), .ZN(n8622) );
  AOI22_X1 U7074 ( .A1(n8649), .A2(n8464), .B1(n8622), .B2(n8465), .ZN(n5560)
         );
  AOI22_X1 U7075 ( .A1(n8616), .A2(n8479), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n5559) );
  NAND2_X1 U7076 ( .A1(n5560), .A2(n5559), .ZN(n5562) );
  NOR3_X1 U7077 ( .A1(n5564), .A2(n5563), .A3(n8490), .ZN(n5561) );
  AOI211_X1 U7078 ( .C1(n8840), .C2(n8461), .A(n5562), .B(n5561), .ZN(n5566)
         );
  NAND2_X1 U7079 ( .A1(n5568), .A2(n4831), .ZN(n5565) );
  OAI211_X1 U7080 ( .C1(n5568), .C2(n5567), .A(n5566), .B(n5565), .ZN(P2_U3222) );
  NOR2_X1 U7081 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5572) );
  NAND2_X1 U7082 ( .A1(n5619), .A2(n5573), .ZN(n5724) );
  INV_X1 U7083 ( .A(n5724), .ZN(n5574) );
  NOR2_X1 U7084 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5577) );
  INV_X1 U7085 ( .A(n5611), .ZN(n5581) );
  NAND2_X1 U7086 ( .A1(n5605), .A2(n5582), .ZN(n5583) );
  INV_X1 U7087 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5614) );
  INV_X1 U7088 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5586) );
  INV_X1 U7089 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U7090 ( .A1(n6021), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5595) );
  INV_X1 U7091 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6723) );
  OR2_X1 U7092 ( .A1(n5677), .A2(n6723), .ZN(n5593) );
  INV_X1 U7093 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5591) );
  OR2_X1 U7094 ( .A1(n6470), .A2(n5591), .ZN(n5592) );
  NAND2_X1 U7095 ( .A1(n5973), .A2(n5599), .ZN(n5631) );
  INV_X1 U7096 ( .A(n5607), .ZN(n5608) );
  NAND2_X1 U7097 ( .A1(n5608), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U7098 ( .A1(n5611), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5612) );
  AND2_X2 U7099 ( .A1(n7163), .A2(n5625), .ZN(n5682) );
  NAND2_X1 U7100 ( .A1(n5615), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5616) );
  NAND2_X1 U7101 ( .A1(n5618), .A2(n5617), .ZN(n6241) );
  NAND2_X2 U7102 ( .A1(n6323), .A2(n6241), .ZN(n6662) );
  NAND2_X1 U7103 ( .A1(n4317), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5624) );
  OR2_X1 U7104 ( .A1(n5619), .A2(n5586), .ZN(n5683) );
  INV_X1 U7105 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5620) );
  NAND2_X1 U7106 ( .A1(n5683), .A2(n5620), .ZN(n5621) );
  NAND2_X1 U7107 ( .A1(n5621), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5622) );
  XNOR2_X1 U7108 ( .A(n5622), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6748) );
  NAND2_X1 U7109 ( .A1(n5708), .A2(n6748), .ZN(n5623) );
  INV_X1 U7110 ( .A(n7400), .ZN(n9941) );
  INV_X1 U7111 ( .A(n5625), .ZN(n5644) );
  INV_X1 U7112 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5626) );
  NAND2_X1 U7113 ( .A1(n5627), .A2(n5626), .ZN(n5628) );
  NAND2_X1 U7114 ( .A1(n5631), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5632) );
  MUX2_X1 U7115 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5632), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n5633) );
  XNOR2_X1 U7116 ( .A(n5634), .B(n6191), .ZN(n5697) );
  INV_X2 U7117 ( .A(n6193), .ZN(n6173) );
  OAI22_X1 U7118 ( .A1(n7143), .A2(n6173), .B1(n9941), .B2(n6117), .ZN(n5698)
         );
  XNOR2_X1 U7119 ( .A(n5697), .B(n5698), .ZN(n6822) );
  INV_X1 U7120 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5635) );
  NAND2_X1 U7121 ( .A1(n5636), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5640) );
  INV_X1 U7122 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9786) );
  INV_X1 U7123 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n5637) );
  NAND2_X1 U7124 ( .A1(n6258), .A2(n5682), .ZN(n5648) );
  XNOR2_X1 U7125 ( .A(n5642), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n6664) );
  MUX2_X1 U7126 ( .A(P1_IR_REG_0__SCAN_IN), .B(n6664), .S(n6662), .Z(n7235) );
  NOR2_X1 U7127 ( .A1(n5625), .A2(n9786), .ZN(n5643) );
  AOI21_X1 U7128 ( .B1(n6179), .B2(n7235), .A(n5643), .ZN(n5649) );
  NAND2_X1 U7129 ( .A1(n5648), .A2(n5649), .ZN(n6813) );
  NAND2_X1 U7130 ( .A1(n5644), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n5645) );
  NAND2_X1 U7131 ( .A1(n6813), .A2(n6814), .ZN(n6812) );
  INV_X1 U7132 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5652) );
  INV_X1 U7133 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7180) );
  INV_X1 U7134 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n5653) );
  INV_X1 U7135 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5654) );
  NAND2_X1 U7136 ( .A1(n6259), .A2(n5682), .ZN(n5665) );
  NAND2_X1 U7137 ( .A1(n4317), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5663) );
  INV_X1 U7138 ( .A(n8054), .ZN(n5659) );
  NAND2_X1 U7139 ( .A1(n4318), .A2(n5659), .ZN(n5662) );
  NAND2_X1 U7140 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5660) );
  NAND2_X1 U7141 ( .A1(n5708), .A2(n9793), .ZN(n5661) );
  AND3_X4 U7142 ( .A1(n5663), .A2(n5662), .A3(n5661), .ZN(n9936) );
  INV_X1 U7143 ( .A(n9936), .ZN(n6304) );
  NAND2_X1 U7144 ( .A1(n6304), .A2(n6179), .ZN(n5664) );
  NAND2_X1 U7145 ( .A1(n5665), .A2(n5664), .ZN(n5666) );
  XNOR2_X1 U7146 ( .A(n5666), .B(n6191), .ZN(n5669) );
  NAND2_X1 U7147 ( .A1(n5670), .A2(n5669), .ZN(n6880) );
  NAND2_X1 U7148 ( .A1(n6193), .A2(n6259), .ZN(n5668) );
  NAND2_X1 U7149 ( .A1(n6304), .A2(n5682), .ZN(n5667) );
  NAND2_X1 U7150 ( .A1(n5668), .A2(n5667), .ZN(n6882) );
  NAND2_X1 U7151 ( .A1(n6880), .A2(n6882), .ZN(n5673) );
  INV_X1 U7152 ( .A(n5669), .ZN(n5672) );
  INV_X1 U7153 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6711) );
  OR2_X1 U7154 ( .A1(n5674), .A2(n6711), .ZN(n5681) );
  INV_X1 U7155 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9327) );
  OR2_X1 U7156 ( .A1(n5675), .A2(n9327), .ZN(n5680) );
  INV_X1 U7157 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5676) );
  NAND2_X1 U7158 ( .A1(n5636), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5678) );
  NAND4_X1 U7159 ( .A1(n5681), .A2(n5680), .A3(n5679), .A4(n5678), .ZN(n5692)
         );
  NAND2_X1 U7160 ( .A1(n5692), .A2(n5682), .ZN(n5690) );
  XNOR2_X1 U7161 ( .A(n5683), .B(P1_IR_REG_2__SCAN_IN), .ZN(n9811) );
  NAND2_X1 U7162 ( .A1(n5708), .A2(n9811), .ZN(n5688) );
  INV_X1 U7163 ( .A(n6669), .ZN(n5684) );
  NAND2_X1 U7164 ( .A1(n9329), .A2(n6179), .ZN(n5689) );
  NAND2_X1 U7165 ( .A1(n5690), .A2(n5689), .ZN(n5691) );
  XNOR2_X1 U7166 ( .A(n5691), .B(n7167), .ZN(n5695) );
  NAND2_X1 U7167 ( .A1(n6193), .A2(n5692), .ZN(n5694) );
  NAND2_X1 U7168 ( .A1(n9329), .A2(n5682), .ZN(n5693) );
  NAND2_X1 U7169 ( .A1(n5694), .A2(n5693), .ZN(n5696) );
  XNOR2_X1 U7170 ( .A(n5695), .B(n5696), .ZN(n6890) );
  NAND2_X1 U7171 ( .A1(n6822), .A2(n6823), .ZN(n5701) );
  INV_X1 U7172 ( .A(n5697), .ZN(n5699) );
  OR2_X1 U7173 ( .A1(n5699), .A2(n5698), .ZN(n5700) );
  NAND2_X1 U7174 ( .A1(n5636), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5706) );
  INV_X1 U7175 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5702) );
  OR2_X1 U7176 ( .A1(n5677), .A2(n5702), .ZN(n5705) );
  XNOR2_X1 U7177 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n7159) );
  OR2_X1 U7178 ( .A1(n5675), .A2(n7159), .ZN(n5704) );
  INV_X1 U7179 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6739) );
  OR2_X1 U7180 ( .A1(n5674), .A2(n6739), .ZN(n5703) );
  NAND2_X1 U7181 ( .A1(n4317), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5711) );
  NAND2_X1 U7182 ( .A1(n5724), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5709) );
  XNOR2_X1 U7183 ( .A(n5709), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9830) );
  NAND2_X1 U7184 ( .A1(n5708), .A2(n9830), .ZN(n5710) );
  INV_X1 U7185 ( .A(n7195), .ZN(n7160) );
  XNOR2_X1 U7186 ( .A(n5712), .B(n7167), .ZN(n5714) );
  OAI22_X1 U7187 ( .A1(n7403), .A2(n6173), .B1(n7160), .B2(n6117), .ZN(n5713)
         );
  XNOR2_X1 U7188 ( .A(n5714), .B(n5713), .ZN(n6992) );
  NAND2_X1 U7189 ( .A1(n5714), .A2(n5713), .ZN(n5715) );
  NAND2_X1 U7190 ( .A1(n6021), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5723) );
  INV_X1 U7191 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7213) );
  OR2_X1 U7192 ( .A1(n5677), .A2(n7213), .ZN(n5722) );
  NAND3_X1 U7193 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5736) );
  INV_X1 U7194 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5717) );
  NAND2_X1 U7195 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5716) );
  NAND2_X1 U7196 ( .A1(n5717), .A2(n5716), .ZN(n5718) );
  NAND2_X1 U7197 ( .A1(n5736), .A2(n5718), .ZN(n7225) );
  OR2_X1 U7198 ( .A1(n5675), .A2(n7225), .ZN(n5721) );
  INV_X1 U7199 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5719) );
  OR2_X1 U7200 ( .A1(n6470), .A2(n5719), .ZN(n5720) );
  OR2_X1 U7201 ( .A1(n7142), .A2(n6173), .ZN(n5732) );
  INV_X1 U7202 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6675) );
  NAND2_X1 U7203 ( .A1(n5685), .A2(n6673), .ZN(n5730) );
  NOR2_X1 U7204 ( .A1(n5724), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5727) );
  OR2_X1 U7205 ( .A1(n5727), .A2(n5586), .ZN(n5725) );
  MUX2_X1 U7206 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5725), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5728) );
  INV_X1 U7207 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5726) );
  NAND2_X1 U7208 ( .A1(n5727), .A2(n5726), .ZN(n5758) );
  NAND2_X1 U7209 ( .A1(n5708), .A2(n9849), .ZN(n5729) );
  OAI211_X1 U7210 ( .C1(n5780), .C2(n6675), .A(n5730), .B(n5729), .ZN(n7227)
         );
  NAND2_X1 U7211 ( .A1(n7227), .A2(n5770), .ZN(n5731) );
  NAND2_X1 U7212 ( .A1(n5732), .A2(n5731), .ZN(n5750) );
  INV_X1 U7213 ( .A(n5750), .ZN(n7224) );
  INV_X1 U7214 ( .A(n7227), .ZN(n7216) );
  OAI22_X1 U7215 ( .A1(n7142), .A2(n6117), .B1(n7216), .B2(n6118), .ZN(n5733)
         );
  XNOR2_X1 U7216 ( .A(n5733), .B(n6191), .ZN(n7222) );
  NAND2_X1 U7217 ( .A1(n6021), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5742) );
  INV_X1 U7218 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n5734) );
  OR2_X1 U7219 ( .A1(n5677), .A2(n5734), .ZN(n5741) );
  INV_X1 U7220 ( .A(n5736), .ZN(n5735) );
  NAND2_X1 U7221 ( .A1(n5735), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5764) );
  INV_X1 U7222 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6789) );
  NAND2_X1 U7223 ( .A1(n5736), .A2(n6789), .ZN(n5737) );
  NAND2_X1 U7224 ( .A1(n5764), .A2(n5737), .ZN(n7282) );
  OR2_X1 U7225 ( .A1(n5675), .A2(n7282), .ZN(n5740) );
  INV_X1 U7226 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5738) );
  OR2_X1 U7227 ( .A1(n6470), .A2(n5738), .ZN(n5739) );
  NAND2_X1 U7228 ( .A1(n5758), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5743) );
  XNOR2_X1 U7229 ( .A(n5743), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6754) );
  AOI22_X1 U7230 ( .A1(n4317), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5708), .B2(
        n6754), .ZN(n5745) );
  NAND2_X1 U7231 ( .A1(n6683), .A2(n5685), .ZN(n5744) );
  NAND2_X1 U7232 ( .A1(n5745), .A2(n5744), .ZN(n7281) );
  INV_X1 U7233 ( .A(n7281), .ZN(n9954) );
  OAI22_X1 U7234 ( .A1(n7388), .A2(n6117), .B1(n9954), .B2(n6118), .ZN(n5746)
         );
  XNOR2_X1 U7235 ( .A(n5746), .B(n6191), .ZN(n7259) );
  OR2_X1 U7236 ( .A1(n7388), .A2(n6173), .ZN(n5748) );
  NAND2_X1 U7237 ( .A1(n7281), .A2(n5770), .ZN(n5747) );
  NAND2_X1 U7238 ( .A1(n5748), .A2(n5747), .ZN(n5752) );
  INV_X1 U7239 ( .A(n5752), .ZN(n7258) );
  AOI22_X1 U7240 ( .A1(n7224), .A2(n7222), .B1(n7259), .B2(n7258), .ZN(n5749)
         );
  NAND2_X1 U7241 ( .A1(n7221), .A2(n5749), .ZN(n5757) );
  INV_X1 U7242 ( .A(n7259), .ZN(n5755) );
  INV_X1 U7243 ( .A(n7222), .ZN(n7257) );
  NAND2_X1 U7244 ( .A1(n7257), .A2(n5750), .ZN(n5751) );
  NAND2_X1 U7245 ( .A1(n5751), .A2(n7258), .ZN(n5754) );
  INV_X1 U7246 ( .A(n5751), .ZN(n5753) );
  AOI22_X1 U7247 ( .A1(n5755), .A2(n5754), .B1(n5753), .B2(n5752), .ZN(n5756)
         );
  NAND2_X1 U7248 ( .A1(n5757), .A2(n5756), .ZN(n7186) );
  NAND2_X1 U7249 ( .A1(n6687), .A2(n5685), .ZN(n5761) );
  NAND2_X1 U7250 ( .A1(n5781), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5759) );
  XNOR2_X1 U7251 ( .A(n5759), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6746) );
  AOI22_X1 U7252 ( .A1(n4317), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5708), .B2(
        n6746), .ZN(n5760) );
  NAND2_X1 U7253 ( .A1(n5636), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5769) );
  NAND2_X1 U7254 ( .A1(n6466), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5768) );
  INV_X1 U7255 ( .A(n5764), .ZN(n5762) );
  NAND2_X1 U7256 ( .A1(n5762), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5786) );
  INV_X1 U7257 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5763) );
  NAND2_X1 U7258 ( .A1(n5764), .A2(n5763), .ZN(n5765) );
  NAND2_X1 U7259 ( .A1(n5786), .A2(n5765), .ZN(n7380) );
  OR2_X1 U7260 ( .A1(n5675), .A2(n7380), .ZN(n5767) );
  INV_X1 U7261 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6735) );
  OR2_X1 U7262 ( .A1(n6468), .A2(n6735), .ZN(n5766) );
  NAND4_X1 U7263 ( .A1(n5769), .A2(n5768), .A3(n5767), .A4(n5766), .ZN(n9079)
         );
  NAND2_X1 U7264 ( .A1(n9079), .A2(n5770), .ZN(n5771) );
  OAI21_X1 U7265 ( .B1(n9960), .B2(n6118), .A(n5771), .ZN(n5772) );
  XNOR2_X1 U7266 ( .A(n5772), .B(n6191), .ZN(n5775) );
  OR2_X1 U7267 ( .A1(n9960), .A2(n6117), .ZN(n5774) );
  NAND2_X1 U7268 ( .A1(n6193), .A2(n9079), .ZN(n5773) );
  AND2_X1 U7269 ( .A1(n5774), .A2(n5773), .ZN(n5776) );
  NAND2_X1 U7270 ( .A1(n7186), .A2(n7184), .ZN(n5779) );
  INV_X1 U7271 ( .A(n5775), .ZN(n5778) );
  INV_X1 U7272 ( .A(n5776), .ZN(n5777) );
  NAND2_X1 U7273 ( .A1(n5778), .A2(n5777), .ZN(n7185) );
  NAND2_X1 U7274 ( .A1(n5779), .A2(n7185), .ZN(n5800) );
  INV_X1 U7275 ( .A(n5800), .ZN(n5795) );
  NAND2_X1 U7276 ( .A1(n6691), .A2(n5685), .ZN(n5784) );
  NAND2_X1 U7277 ( .A1(n5801), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5782) );
  XNOR2_X1 U7278 ( .A(n5782), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6968) );
  AOI22_X1 U7279 ( .A1(n4317), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5708), .B2(
        n6968), .ZN(n5783) );
  NAND2_X1 U7280 ( .A1(n5784), .A2(n5783), .ZN(n7450) );
  NAND2_X1 U7281 ( .A1(n7450), .A2(n5770), .ZN(n5793) );
  NAND2_X1 U7282 ( .A1(n5636), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5791) );
  INV_X1 U7283 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6758) );
  OR2_X1 U7284 ( .A1(n5677), .A2(n6758), .ZN(n5790) );
  INV_X1 U7285 ( .A(n5786), .ZN(n5785) );
  NAND2_X1 U7286 ( .A1(n5785), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5809) );
  INV_X1 U7287 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6734) );
  NAND2_X1 U7288 ( .A1(n5786), .A2(n6734), .ZN(n5787) );
  NAND2_X1 U7289 ( .A1(n5809), .A2(n5787), .ZN(n7311) );
  OR2_X1 U7290 ( .A1(n5675), .A2(n7311), .ZN(n5789) );
  INV_X1 U7291 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6742) );
  OR2_X1 U7292 ( .A1(n6468), .A2(n6742), .ZN(n5788) );
  OR2_X1 U7293 ( .A1(n9917), .A2(n6173), .ZN(n5792) );
  NAND2_X1 U7294 ( .A1(n5793), .A2(n5792), .ZN(n5799) );
  NAND2_X1 U7295 ( .A1(n5795), .A2(n5794), .ZN(n7307) );
  NAND2_X1 U7296 ( .A1(n7450), .A2(n6179), .ZN(n5797) );
  OR2_X1 U7297 ( .A1(n9917), .A2(n6117), .ZN(n5796) );
  NAND2_X1 U7298 ( .A1(n5797), .A2(n5796), .ZN(n5798) );
  XNOR2_X1 U7299 ( .A(n5798), .B(n7167), .ZN(n7310) );
  NAND2_X1 U7300 ( .A1(n5800), .A2(n5799), .ZN(n7308) );
  NAND2_X1 U7301 ( .A1(n6701), .A2(n5685), .ZN(n5807) );
  NOR2_X1 U7302 ( .A1(n5801), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5804) );
  OR2_X1 U7303 ( .A1(n5804), .A2(n5586), .ZN(n5802) );
  MUX2_X1 U7304 ( .A(n5802), .B(P1_IR_REG_31__SCAN_IN), .S(n5803), .Z(n5805)
         );
  NAND2_X1 U7305 ( .A1(n5804), .A2(n5803), .ZN(n5839) );
  NAND2_X1 U7306 ( .A1(n5805), .A2(n5839), .ZN(n6703) );
  AOI22_X1 U7307 ( .A1(n4317), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5708), .B2(
        n9866), .ZN(n5806) );
  NAND2_X1 U7308 ( .A1(n5807), .A2(n5806), .ZN(n9904) );
  NAND2_X1 U7309 ( .A1(n9904), .A2(n6179), .ZN(n5817) );
  NAND2_X1 U7310 ( .A1(n6466), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5815) );
  NAND2_X1 U7311 ( .A1(n5636), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5814) );
  NAND2_X1 U7312 ( .A1(n5809), .A2(n5808), .ZN(n5810) );
  NAND2_X1 U7313 ( .A1(n5827), .A2(n5810), .ZN(n9926) );
  OR2_X1 U7314 ( .A1(n5675), .A2(n9926), .ZN(n5813) );
  INV_X1 U7315 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5811) );
  OR2_X1 U7316 ( .A1(n6468), .A2(n5811), .ZN(n5812) );
  NAND4_X1 U7317 ( .A1(n5815), .A2(n5814), .A3(n5813), .A4(n5812), .ZN(n9077)
         );
  NAND2_X1 U7318 ( .A1(n9077), .A2(n5770), .ZN(n5816) );
  NAND2_X1 U7319 ( .A1(n5817), .A2(n5816), .ZN(n5818) );
  XNOR2_X1 U7320 ( .A(n5818), .B(n6191), .ZN(n5822) );
  AND2_X1 U7321 ( .A1(n6193), .A2(n9077), .ZN(n5819) );
  AOI21_X1 U7322 ( .B1(n9904), .B2(n5770), .A(n5819), .ZN(n5821) );
  XNOR2_X1 U7323 ( .A(n5822), .B(n5821), .ZN(n7522) );
  NAND2_X1 U7324 ( .A1(n5822), .A2(n5821), .ZN(n5823) );
  NAND2_X1 U7325 ( .A1(n7520), .A2(n5823), .ZN(n7560) );
  NAND2_X1 U7326 ( .A1(n5839), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5825) );
  XNOR2_X1 U7327 ( .A(n5825), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9879) );
  AOI22_X1 U7328 ( .A1(n4317), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5708), .B2(
        n9879), .ZN(n5826) );
  NAND2_X1 U7329 ( .A1(n9660), .A2(n6179), .ZN(n5835) );
  NAND2_X1 U7330 ( .A1(n5636), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5833) );
  INV_X1 U7331 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7617) );
  OR2_X1 U7332 ( .A1(n5677), .A2(n7617), .ZN(n5832) );
  NAND2_X1 U7333 ( .A1(n5827), .A2(n7561), .ZN(n5828) );
  NAND2_X1 U7334 ( .A1(n5845), .A2(n5828), .ZN(n7616) );
  OR2_X1 U7335 ( .A1(n5675), .A2(n7616), .ZN(n5831) );
  INV_X1 U7336 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n5829) );
  OR2_X1 U7337 ( .A1(n6468), .A2(n5829), .ZN(n5830) );
  OR2_X1 U7338 ( .A1(n9915), .A2(n6117), .ZN(n5834) );
  NAND2_X1 U7339 ( .A1(n5835), .A2(n5834), .ZN(n5836) );
  XNOR2_X1 U7340 ( .A(n5836), .B(n6191), .ZN(n7558) );
  NOR2_X1 U7341 ( .A1(n9915), .A2(n6173), .ZN(n5837) );
  AOI21_X1 U7342 ( .B1(n9660), .B2(n5770), .A(n5837), .ZN(n7557) );
  AND2_X1 U7343 ( .A1(n7558), .A2(n7557), .ZN(n5838) );
  NAND2_X1 U7344 ( .A1(n6706), .A2(n5685), .ZN(n5842) );
  OAI21_X1 U7345 ( .B1(n5839), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5840) );
  XNOR2_X1 U7346 ( .A(n5840), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6983) );
  AOI22_X1 U7347 ( .A1(n4317), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5708), .B2(
        n6983), .ZN(n5841) );
  NAND2_X1 U7348 ( .A1(n9759), .A2(n6179), .ZN(n5852) );
  NAND2_X1 U7349 ( .A1(n6021), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5850) );
  NAND2_X1 U7350 ( .A1(n5636), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5849) );
  INV_X1 U7351 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9726) );
  OR2_X1 U7352 ( .A1(n5677), .A2(n9726), .ZN(n5848) );
  INV_X1 U7353 ( .A(n5845), .ZN(n5843) );
  NAND2_X1 U7354 ( .A1(n5843), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5867) );
  INV_X1 U7355 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5844) );
  NAND2_X1 U7356 ( .A1(n5845), .A2(n5844), .ZN(n5846) );
  NAND2_X1 U7357 ( .A1(n5867), .A2(n5846), .ZN(n9725) );
  OR2_X1 U7358 ( .A1(n5675), .A2(n9725), .ZN(n5847) );
  NAND4_X1 U7359 ( .A1(n5850), .A2(n5849), .A3(n5848), .A4(n5847), .ZN(n9075)
         );
  NAND2_X1 U7360 ( .A1(n9075), .A2(n5770), .ZN(n5851) );
  NAND2_X1 U7361 ( .A1(n5852), .A2(n5851), .ZN(n5853) );
  XNOR2_X1 U7362 ( .A(n5853), .B(n7167), .ZN(n5857) );
  AND2_X1 U7363 ( .A1(n6193), .A2(n9075), .ZN(n5854) );
  AOI21_X1 U7364 ( .B1(n9759), .B2(n5770), .A(n5854), .ZN(n5855) );
  XNOR2_X1 U7365 ( .A(n5857), .B(n5855), .ZN(n7691) );
  INV_X1 U7366 ( .A(n5855), .ZN(n5856) );
  NAND2_X1 U7367 ( .A1(n5857), .A2(n5856), .ZN(n5858) );
  NAND2_X1 U7368 ( .A1(n5859), .A2(n5685), .ZN(n5863) );
  NAND2_X1 U7369 ( .A1(n5860), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5861) );
  XNOR2_X1 U7370 ( .A(n5861), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7111) );
  AOI22_X1 U7371 ( .A1(n4317), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5708), .B2(
        n7111), .ZN(n5862) );
  NAND2_X1 U7372 ( .A1(n9411), .A2(n6179), .ZN(n5875) );
  NAND2_X1 U7373 ( .A1(n6466), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5873) );
  INV_X1 U7374 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n5864) );
  OR2_X1 U7375 ( .A1(n6470), .A2(n5864), .ZN(n5872) );
  INV_X1 U7376 ( .A(n5867), .ZN(n5865) );
  NAND2_X1 U7377 ( .A1(n5865), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5889) );
  INV_X1 U7378 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5866) );
  NAND2_X1 U7379 ( .A1(n5867), .A2(n5866), .ZN(n5868) );
  NAND2_X1 U7380 ( .A1(n5889), .A2(n5868), .ZN(n7855) );
  OR2_X1 U7381 ( .A1(n5675), .A2(n7855), .ZN(n5871) );
  INV_X1 U7382 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n5869) );
  OR2_X1 U7383 ( .A1(n6468), .A2(n5869), .ZN(n5870) );
  OR2_X1 U7384 ( .A1(n9729), .A2(n6117), .ZN(n5874) );
  NAND2_X1 U7385 ( .A1(n5875), .A2(n5874), .ZN(n5876) );
  XNOR2_X1 U7386 ( .A(n5876), .B(n6191), .ZN(n5879) );
  NOR2_X1 U7387 ( .A1(n9729), .A2(n6173), .ZN(n5877) );
  AOI21_X1 U7388 ( .B1(n9411), .B2(n5770), .A(n5877), .ZN(n5878) );
  NAND2_X1 U7389 ( .A1(n5879), .A2(n5878), .ZN(n5882) );
  OR2_X1 U7390 ( .A1(n5879), .A2(n5878), .ZN(n5880) );
  NAND2_X1 U7391 ( .A1(n5882), .A2(n5880), .ZN(n7824) );
  NAND2_X1 U7392 ( .A1(n5883), .A2(n5685), .ZN(n5887) );
  OR2_X1 U7393 ( .A1(n5884), .A2(n5586), .ZN(n5885) );
  XNOR2_X1 U7394 ( .A(n5885), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7485) );
  AOI22_X1 U7395 ( .A1(n4317), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5708), .B2(
        n7485), .ZN(n5886) );
  NAND2_X1 U7396 ( .A1(n9717), .A2(n6179), .ZN(n5896) );
  NAND2_X1 U7397 ( .A1(n5636), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U7398 ( .A1(n6021), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5893) );
  INV_X1 U7399 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9704) );
  OR2_X1 U7400 ( .A1(n5677), .A2(n9704), .ZN(n5892) );
  NAND2_X1 U7401 ( .A1(n5889), .A2(n5888), .ZN(n5890) );
  NAND2_X1 U7402 ( .A1(n5911), .A2(n5890), .ZN(n9703) );
  OR2_X1 U7403 ( .A1(n5675), .A2(n9703), .ZN(n5891) );
  NAND4_X1 U7404 ( .A1(n5894), .A2(n5893), .A3(n5892), .A4(n5891), .ZN(n9074)
         );
  NAND2_X1 U7405 ( .A1(n9074), .A2(n5770), .ZN(n5895) );
  NAND2_X1 U7406 ( .A1(n5896), .A2(n5895), .ZN(n5897) );
  XNOR2_X1 U7407 ( .A(n5897), .B(n6191), .ZN(n5899) );
  AND2_X1 U7408 ( .A1(n6193), .A2(n9074), .ZN(n5898) );
  AOI21_X1 U7409 ( .B1(n9717), .B2(n5770), .A(n5898), .ZN(n5900) );
  AND2_X1 U7410 ( .A1(n5899), .A2(n5900), .ZN(n7833) );
  INV_X1 U7411 ( .A(n5899), .ZN(n5902) );
  INV_X1 U7412 ( .A(n5900), .ZN(n5901) );
  NAND2_X1 U7413 ( .A1(n5902), .A2(n5901), .ZN(n7834) );
  NAND2_X1 U7414 ( .A1(n6818), .A2(n5685), .ZN(n5908) );
  OR2_X1 U7415 ( .A1(n5973), .A2(n5586), .ZN(n5905) );
  INV_X1 U7416 ( .A(n5905), .ZN(n5903) );
  NAND2_X1 U7417 ( .A1(n5903), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5906) );
  NAND2_X1 U7418 ( .A1(n5905), .A2(n5904), .ZN(n5922) );
  AOI22_X1 U7419 ( .A1(n4317), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5708), .B2(
        n7743), .ZN(n5907) );
  NAND2_X1 U7420 ( .A1(n9407), .A2(n6179), .ZN(n5919) );
  NAND2_X1 U7421 ( .A1(n6466), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5917) );
  NAND2_X1 U7422 ( .A1(n5636), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5916) );
  INV_X1 U7423 ( .A(n5911), .ZN(n5909) );
  NAND2_X1 U7424 ( .A1(n5909), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5928) );
  INV_X1 U7425 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5910) );
  NAND2_X1 U7426 ( .A1(n5911), .A2(n5910), .ZN(n5912) );
  NAND2_X1 U7427 ( .A1(n5928), .A2(n5912), .ZN(n7995) );
  OR2_X1 U7428 ( .A1(n5675), .A2(n7995), .ZN(n5915) );
  INV_X1 U7429 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n5913) );
  OR2_X1 U7430 ( .A1(n6468), .A2(n5913), .ZN(n5914) );
  NAND4_X1 U7431 ( .A1(n5917), .A2(n5916), .A3(n5915), .A4(n5914), .ZN(n9708)
         );
  NAND2_X1 U7432 ( .A1(n9708), .A2(n5770), .ZN(n5918) );
  NAND2_X1 U7433 ( .A1(n5919), .A2(n5918), .ZN(n5920) );
  XNOR2_X1 U7434 ( .A(n5920), .B(n6191), .ZN(n5938) );
  INV_X1 U7435 ( .A(n5938), .ZN(n5921) );
  NAND2_X1 U7436 ( .A1(n6999), .A2(n5685), .ZN(n5926) );
  NAND2_X1 U7437 ( .A1(n5922), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5924) );
  INV_X1 U7438 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5923) );
  XNOR2_X1 U7439 ( .A(n5924), .B(n5923), .ZN(n9106) );
  INV_X1 U7440 ( .A(n9106), .ZN(n7746) );
  AOI22_X1 U7441 ( .A1(n4317), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5708), .B2(
        n7746), .ZN(n5925) );
  NAND2_X1 U7442 ( .A1(n6466), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5934) );
  NAND2_X1 U7443 ( .A1(n5636), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5933) );
  NAND2_X1 U7444 ( .A1(n5928), .A2(n5927), .ZN(n5929) );
  NAND2_X1 U7445 ( .A1(n5956), .A2(n5929), .ZN(n8046) );
  OR2_X1 U7446 ( .A1(n5675), .A2(n8046), .ZN(n5932) );
  INV_X1 U7447 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n5930) );
  OR2_X1 U7448 ( .A1(n6468), .A2(n5930), .ZN(n5931) );
  NAND4_X1 U7449 ( .A1(n5934), .A2(n5933), .A3(n5932), .A4(n5931), .ZN(n9073)
         );
  INV_X1 U7450 ( .A(n9073), .ZN(n8991) );
  OAI22_X1 U7451 ( .A1(n9747), .A2(n6118), .B1(n8991), .B2(n6117), .ZN(n5935)
         );
  XNOR2_X1 U7452 ( .A(n5935), .B(n7167), .ZN(n5946) );
  INV_X1 U7453 ( .A(n5946), .ZN(n5936) );
  AND2_X1 U7454 ( .A1(n7989), .A2(n5936), .ZN(n5942) );
  NAND2_X1 U7455 ( .A1(n5939), .A2(n5938), .ZN(n7990) );
  NAND2_X1 U7456 ( .A1(n9407), .A2(n5770), .ZN(n5941) );
  NAND2_X1 U7457 ( .A1(n6193), .A2(n9708), .ZN(n5940) );
  NAND2_X1 U7458 ( .A1(n5941), .A2(n5940), .ZN(n7992) );
  NAND2_X1 U7459 ( .A1(n5942), .A2(n5945), .ZN(n8038) );
  OR2_X1 U7460 ( .A1(n9747), .A2(n6117), .ZN(n5944) );
  NAND2_X1 U7461 ( .A1(n6193), .A2(n9073), .ZN(n5943) );
  NAND2_X1 U7462 ( .A1(n5944), .A2(n5943), .ZN(n8041) );
  NAND2_X1 U7463 ( .A1(n5945), .A2(n7989), .ZN(n5947) );
  NAND2_X1 U7464 ( .A1(n7037), .A2(n4318), .ZN(n5952) );
  NAND2_X1 U7465 ( .A1(n5973), .A2(n5948), .ZN(n5949) );
  NAND2_X1 U7466 ( .A1(n5949), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5950) );
  XNOR2_X1 U7467 ( .A(n5950), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9124) );
  AOI22_X1 U7468 ( .A1(n4317), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5708), .B2(
        n9124), .ZN(n5951) );
  NAND2_X1 U7469 ( .A1(n9401), .A2(n6179), .ZN(n5964) );
  NAND2_X1 U7470 ( .A1(n6466), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5962) );
  INV_X1 U7471 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n5953) );
  OR2_X1 U7472 ( .A1(n6470), .A2(n5953), .ZN(n5961) );
  INV_X1 U7473 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5955) );
  NAND2_X1 U7474 ( .A1(n5956), .A2(n5955), .ZN(n5957) );
  NAND2_X1 U7475 ( .A1(n5981), .A2(n5957), .ZN(n8995) );
  OR2_X1 U7476 ( .A1(n5675), .A2(n8995), .ZN(n5960) );
  INV_X1 U7477 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n5958) );
  OR2_X1 U7478 ( .A1(n6468), .A2(n5958), .ZN(n5959) );
  OR2_X1 U7479 ( .A1(n9005), .A2(n6117), .ZN(n5963) );
  NAND2_X1 U7480 ( .A1(n5964), .A2(n5963), .ZN(n5965) );
  XNOR2_X1 U7481 ( .A(n5965), .B(n7167), .ZN(n5968) );
  NAND2_X1 U7482 ( .A1(n9401), .A2(n5682), .ZN(n5967) );
  OR2_X1 U7483 ( .A1(n9005), .A2(n6173), .ZN(n5966) );
  NAND2_X1 U7484 ( .A1(n5967), .A2(n5966), .ZN(n5969) );
  INV_X1 U7485 ( .A(n5968), .ZN(n5971) );
  INV_X1 U7486 ( .A(n5969), .ZN(n5970) );
  NAND2_X1 U7487 ( .A1(n5971), .A2(n5970), .ZN(n8989) );
  NAND2_X1 U7488 ( .A1(n7136), .A2(n4318), .ZN(n5980) );
  NAND2_X1 U7489 ( .A1(n5973), .A2(n5972), .ZN(n5974) );
  NAND2_X1 U7490 ( .A1(n5974), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5977) );
  INV_X1 U7491 ( .A(n5977), .ZN(n5975) );
  NAND2_X1 U7492 ( .A1(n5975), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n5978) );
  INV_X1 U7493 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5976) );
  NAND2_X1 U7494 ( .A1(n5977), .A2(n5976), .ZN(n5997) );
  AOI22_X1 U7495 ( .A1(n4317), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5708), .B2(
        n9138), .ZN(n5979) );
  NAND2_X1 U7496 ( .A1(n9394), .A2(n6179), .ZN(n5990) );
  NAND2_X1 U7497 ( .A1(n5981), .A2(n9003), .ZN(n5982) );
  AND2_X1 U7498 ( .A1(n6003), .A2(n5982), .ZN(n9007) );
  NAND2_X1 U7499 ( .A1(n9007), .A2(n6235), .ZN(n5988) );
  NAND2_X1 U7500 ( .A1(n5636), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5987) );
  INV_X1 U7501 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n5983) );
  OR2_X1 U7502 ( .A1(n5677), .A2(n5983), .ZN(n5986) );
  INV_X1 U7503 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n5984) );
  OR2_X1 U7504 ( .A1(n6468), .A2(n5984), .ZN(n5985) );
  NAND4_X1 U7505 ( .A1(n5988), .A2(n5987), .A3(n5986), .A4(n5985), .ZN(n9320)
         );
  NAND2_X1 U7506 ( .A1(n9320), .A2(n5770), .ZN(n5989) );
  NAND2_X1 U7507 ( .A1(n5990), .A2(n5989), .ZN(n5991) );
  XNOR2_X1 U7508 ( .A(n5991), .B(n7167), .ZN(n5993) );
  AND2_X1 U7509 ( .A1(n6193), .A2(n9320), .ZN(n5992) );
  AOI21_X1 U7510 ( .B1(n9394), .B2(n5770), .A(n5992), .ZN(n5994) );
  XNOR2_X1 U7511 ( .A(n5993), .B(n5994), .ZN(n9001) );
  INV_X1 U7512 ( .A(n5993), .ZN(n5995) );
  NAND2_X1 U7513 ( .A1(n5995), .A2(n5994), .ZN(n5996) );
  NAND2_X1 U7514 ( .A1(n7252), .A2(n5685), .ZN(n6000) );
  NAND2_X1 U7515 ( .A1(n5997), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5998) );
  XNOR2_X1 U7516 ( .A(n5998), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9885) );
  AOI22_X1 U7517 ( .A1(n4317), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5708), .B2(
        n9885), .ZN(n5999) );
  NAND2_X1 U7518 ( .A1(n9389), .A2(n6179), .ZN(n6013) );
  INV_X1 U7519 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6002) );
  NAND2_X1 U7520 ( .A1(n6003), .A2(n6002), .ZN(n6004) );
  NAND2_X1 U7521 ( .A1(n6019), .A2(n6004), .ZN(n9310) );
  OR2_X1 U7522 ( .A1(n9310), .A2(n5675), .ZN(n6011) );
  INV_X1 U7523 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n6005) );
  OR2_X1 U7524 ( .A1(n5677), .A2(n6005), .ZN(n6008) );
  INV_X1 U7525 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n6006) );
  OR2_X1 U7526 ( .A1(n6470), .A2(n6006), .ZN(n6007) );
  AND2_X1 U7527 ( .A1(n6008), .A2(n6007), .ZN(n6010) );
  INV_X1 U7528 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9136) );
  OR2_X1 U7529 ( .A1(n6468), .A2(n9136), .ZN(n6009) );
  NAND2_X1 U7530 ( .A1(n9299), .A2(n5770), .ZN(n6012) );
  NAND2_X1 U7531 ( .A1(n6013), .A2(n6012), .ZN(n6014) );
  XNOR2_X1 U7532 ( .A(n6014), .B(n6191), .ZN(n9043) );
  NOR2_X1 U7533 ( .A1(n6280), .A2(n6173), .ZN(n6015) );
  AOI21_X1 U7534 ( .B1(n9389), .B2(n5770), .A(n6015), .ZN(n9042) );
  NAND2_X1 U7535 ( .A1(n7303), .A2(n4318), .ZN(n6017) );
  AOI22_X1 U7536 ( .A1(n4317), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n5708), .B2(
        n9272), .ZN(n6016) );
  NAND2_X1 U7537 ( .A1(n9384), .A2(n6179), .ZN(n6025) );
  NAND2_X1 U7538 ( .A1(n6019), .A2(n6018), .ZN(n6020) );
  NAND2_X1 U7539 ( .A1(n6035), .A2(n6020), .ZN(n9292) );
  AOI22_X1 U7540 ( .A1(n6021), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n6466), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U7541 ( .A1(n5636), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6022) );
  OAI211_X1 U7542 ( .C1(n9292), .C2(n5675), .A(n6023), .B(n6022), .ZN(n9319)
         );
  NAND2_X1 U7543 ( .A1(n9319), .A2(n5682), .ZN(n6024) );
  NAND2_X1 U7544 ( .A1(n6025), .A2(n6024), .ZN(n6026) );
  XNOR2_X1 U7545 ( .A(n6026), .B(n7167), .ZN(n6028) );
  AND2_X1 U7546 ( .A1(n9319), .A2(n6193), .ZN(n6027) );
  AOI21_X1 U7547 ( .B1(n9384), .B2(n5770), .A(n6027), .ZN(n6029) );
  XNOR2_X1 U7548 ( .A(n6028), .B(n6029), .ZN(n8962) );
  INV_X1 U7549 ( .A(n6028), .ZN(n6030) );
  NAND2_X1 U7550 ( .A1(n6030), .A2(n6029), .ZN(n9020) );
  NAND2_X1 U7551 ( .A1(n7510), .A2(n4318), .ZN(n6032) );
  NAND2_X1 U7552 ( .A1(n4317), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U7553 ( .A1(n9379), .A2(n6179), .ZN(n6044) );
  INV_X1 U7554 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U7555 ( .A1(n6035), .A2(n6034), .ZN(n6036) );
  NAND2_X1 U7556 ( .A1(n6055), .A2(n6036), .ZN(n9279) );
  OR2_X1 U7557 ( .A1(n9279), .A2(n5675), .ZN(n6042) );
  INV_X1 U7558 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n6039) );
  NAND2_X1 U7559 ( .A1(n6466), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6038) );
  NAND2_X1 U7560 ( .A1(n5636), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6037) );
  OAI211_X1 U7561 ( .C1(n6468), .C2(n6039), .A(n6038), .B(n6037), .ZN(n6040)
         );
  INV_X1 U7562 ( .A(n6040), .ZN(n6041) );
  NAND2_X1 U7563 ( .A1(n6042), .A2(n6041), .ZN(n9298) );
  NAND2_X1 U7564 ( .A1(n9298), .A2(n5682), .ZN(n6043) );
  NAND2_X1 U7565 ( .A1(n6044), .A2(n6043), .ZN(n6045) );
  XNOR2_X1 U7566 ( .A(n6045), .B(n7167), .ZN(n6050) );
  INV_X1 U7567 ( .A(n6050), .ZN(n6047) );
  AND2_X1 U7568 ( .A1(n9298), .A2(n6193), .ZN(n6046) );
  AOI21_X1 U7569 ( .B1(n9379), .B2(n5682), .A(n6046), .ZN(n6049) );
  NAND2_X1 U7570 ( .A1(n6047), .A2(n6049), .ZN(n6048) );
  AND2_X1 U7571 ( .A1(n9020), .A2(n6048), .ZN(n6052) );
  INV_X1 U7572 ( .A(n6048), .ZN(n6051) );
  XNOR2_X1 U7573 ( .A(n6050), .B(n6049), .ZN(n9023) );
  NAND2_X1 U7574 ( .A1(n7577), .A2(n5685), .ZN(n6054) );
  NAND2_X1 U7575 ( .A1(n4317), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U7576 ( .A1(n9372), .A2(n6179), .ZN(n6064) );
  NAND2_X1 U7577 ( .A1(n6055), .A2(n8971), .ZN(n6056) );
  NAND2_X1 U7578 ( .A1(n6074), .A2(n6056), .ZN(n9271) );
  OR2_X1 U7579 ( .A1(n9271), .A2(n5675), .ZN(n6062) );
  INV_X1 U7580 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n6059) );
  NAND2_X1 U7581 ( .A1(n6466), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6058) );
  NAND2_X1 U7582 ( .A1(n5636), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6057) );
  OAI211_X1 U7583 ( .C1(n6059), .C2(n6468), .A(n6058), .B(n6057), .ZN(n6060)
         );
  INV_X1 U7584 ( .A(n6060), .ZN(n6061) );
  NAND2_X1 U7585 ( .A1(n9285), .A2(n5770), .ZN(n6063) );
  NAND2_X1 U7586 ( .A1(n6064), .A2(n6063), .ZN(n6065) );
  XNOR2_X1 U7587 ( .A(n6065), .B(n7167), .ZN(n6067) );
  NOR2_X1 U7588 ( .A1(n9035), .A2(n6173), .ZN(n6066) );
  AOI21_X1 U7589 ( .B1(n9372), .B2(n5682), .A(n6066), .ZN(n6068) );
  XNOR2_X1 U7590 ( .A(n6067), .B(n6068), .ZN(n8969) );
  NAND2_X1 U7591 ( .A1(n8970), .A2(n8969), .ZN(n6071) );
  INV_X1 U7592 ( .A(n6067), .ZN(n6069) );
  NAND2_X1 U7593 ( .A1(n6069), .A2(n6068), .ZN(n6070) );
  NAND2_X1 U7594 ( .A1(n6071), .A2(n6070), .ZN(n6097) );
  NAND2_X1 U7595 ( .A1(n7712), .A2(n5685), .ZN(n6073) );
  NAND2_X1 U7596 ( .A1(n4317), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6072) );
  INV_X1 U7597 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9034) );
  NAND2_X1 U7598 ( .A1(n6074), .A2(n9034), .ZN(n6075) );
  AND2_X1 U7599 ( .A1(n6109), .A2(n6075), .ZN(n9249) );
  NAND2_X1 U7600 ( .A1(n9249), .A2(n6235), .ZN(n6081) );
  INV_X1 U7601 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n6078) );
  NAND2_X1 U7602 ( .A1(n5636), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6077) );
  NAND2_X1 U7603 ( .A1(n6466), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6076) );
  OAI211_X1 U7604 ( .C1(n6078), .C2(n6468), .A(n6077), .B(n6076), .ZN(n6079)
         );
  INV_X1 U7605 ( .A(n6079), .ZN(n6080) );
  AND2_X1 U7606 ( .A1(n9265), .A2(n6193), .ZN(n6082) );
  AOI21_X1 U7607 ( .B1(n9366), .B2(n5682), .A(n6082), .ZN(n6098) );
  NAND2_X1 U7608 ( .A1(n6097), .A2(n6098), .ZN(n9030) );
  NAND2_X1 U7609 ( .A1(n9366), .A2(n6179), .ZN(n6084) );
  NAND2_X1 U7610 ( .A1(n9265), .A2(n5770), .ZN(n6083) );
  NAND2_X1 U7611 ( .A1(n6084), .A2(n6083), .ZN(n6085) );
  XNOR2_X1 U7612 ( .A(n6085), .B(n7167), .ZN(n9033) );
  NAND2_X1 U7613 ( .A1(n7816), .A2(n5685), .ZN(n6087) );
  NAND2_X1 U7614 ( .A1(n4317), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7615 ( .A1(n9363), .A2(n6179), .ZN(n6095) );
  XNOR2_X1 U7616 ( .A(n6109), .B(P1_REG3_REG_23__SCAN_IN), .ZN(n9239) );
  NAND2_X1 U7617 ( .A1(n9239), .A2(n6235), .ZN(n6093) );
  INV_X1 U7618 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n6090) );
  NAND2_X1 U7619 ( .A1(n6466), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6089) );
  NAND2_X1 U7620 ( .A1(n5636), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6088) );
  OAI211_X1 U7621 ( .C1(n6468), .C2(n6090), .A(n6089), .B(n6088), .ZN(n6091)
         );
  INV_X1 U7622 ( .A(n6091), .ZN(n6092) );
  NAND2_X1 U7623 ( .A1(n9254), .A2(n5770), .ZN(n6094) );
  NAND2_X1 U7624 ( .A1(n6095), .A2(n6094), .ZN(n6096) );
  XNOR2_X1 U7625 ( .A(n6096), .B(n6191), .ZN(n6101) );
  AOI22_X1 U7626 ( .A1(n9363), .A2(n5682), .B1(n6193), .B2(n9254), .ZN(n8952)
         );
  NAND2_X1 U7627 ( .A1(n7890), .A2(n4318), .ZN(n6104) );
  NAND2_X1 U7628 ( .A1(n4317), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6103) );
  INV_X1 U7629 ( .A(n6109), .ZN(n6106) );
  AND2_X1 U7630 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(P1_REG3_REG_23__SCAN_IN), 
        .ZN(n6105) );
  NAND2_X1 U7631 ( .A1(n6106), .A2(n6105), .ZN(n6127) );
  INV_X1 U7632 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6108) );
  INV_X1 U7633 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6107) );
  OAI21_X1 U7634 ( .B1(n6109), .B2(n6108), .A(n6107), .ZN(n6110) );
  NAND2_X1 U7635 ( .A1(n6127), .A2(n6110), .ZN(n9224) );
  INV_X1 U7636 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n6113) );
  NAND2_X1 U7637 ( .A1(n6466), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6112) );
  NAND2_X1 U7638 ( .A1(n5636), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6111) );
  OAI211_X1 U7639 ( .C1(n6468), .C2(n6113), .A(n6112), .B(n6111), .ZN(n6114)
         );
  INV_X1 U7640 ( .A(n6114), .ZN(n6115) );
  OAI22_X1 U7641 ( .A1(n9019), .A2(n6117), .B1(n6349), .B2(n6173), .ZN(n6120)
         );
  OAI22_X1 U7642 ( .A1(n9019), .A2(n6118), .B1(n6349), .B2(n6117), .ZN(n6119)
         );
  XNOR2_X1 U7643 ( .A(n6119), .B(n7167), .ZN(n6121) );
  XOR2_X1 U7644 ( .A(n6120), .B(n6121), .Z(n9013) );
  OR2_X1 U7645 ( .A1(n6121), .A2(n6120), .ZN(n6122) );
  NAND2_X1 U7646 ( .A1(n4317), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6123) );
  NAND2_X1 U7647 ( .A1(n9351), .A2(n6179), .ZN(n6136) );
  INV_X1 U7648 ( .A(n6127), .ZN(n6125) );
  NAND2_X1 U7649 ( .A1(n6125), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6143) );
  INV_X1 U7650 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6126) );
  NAND2_X1 U7651 ( .A1(n6127), .A2(n6126), .ZN(n6128) );
  NAND2_X1 U7652 ( .A1(n6143), .A2(n6128), .ZN(n9201) );
  OR2_X1 U7653 ( .A1(n9201), .A2(n5675), .ZN(n6134) );
  INV_X1 U7654 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n6131) );
  NAND2_X1 U7655 ( .A1(n6466), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6130) );
  NAND2_X1 U7656 ( .A1(n5636), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6129) );
  OAI211_X1 U7657 ( .C1(n6468), .C2(n6131), .A(n6130), .B(n6129), .ZN(n6132)
         );
  INV_X1 U7658 ( .A(n6132), .ZN(n6133) );
  NAND2_X1 U7659 ( .A1(n9217), .A2(n5682), .ZN(n6135) );
  NAND2_X1 U7660 ( .A1(n6136), .A2(n6135), .ZN(n6137) );
  XNOR2_X1 U7661 ( .A(n6137), .B(n7167), .ZN(n6138) );
  AOI22_X1 U7662 ( .A1(n9351), .A2(n5682), .B1(n6193), .B2(n9217), .ZN(n6139)
         );
  XNOR2_X1 U7663 ( .A(n6138), .B(n6139), .ZN(n8979) );
  INV_X1 U7664 ( .A(n6138), .ZN(n6140) );
  NAND2_X1 U7665 ( .A1(n8013), .A2(n5685), .ZN(n6142) );
  NAND2_X1 U7666 ( .A1(n4317), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6141) );
  NAND2_X1 U7667 ( .A1(n9346), .A2(n6179), .ZN(n6152) );
  INV_X1 U7668 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9059) );
  NAND2_X1 U7669 ( .A1(n6143), .A2(n9059), .ZN(n6144) );
  NAND2_X1 U7670 ( .A1(n9189), .A2(n6235), .ZN(n6150) );
  INV_X1 U7671 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U7672 ( .A1(n5636), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6146) );
  NAND2_X1 U7673 ( .A1(n6466), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6145) );
  OAI211_X1 U7674 ( .C1(n6147), .C2(n6468), .A(n6146), .B(n6145), .ZN(n6148)
         );
  INV_X1 U7675 ( .A(n6148), .ZN(n6149) );
  NAND2_X1 U7676 ( .A1(n9208), .A2(n5770), .ZN(n6151) );
  NAND2_X1 U7677 ( .A1(n6152), .A2(n6151), .ZN(n6153) );
  XNOR2_X1 U7678 ( .A(n6153), .B(n7167), .ZN(n6155) );
  AND2_X1 U7679 ( .A1(n9208), .A2(n6193), .ZN(n6154) );
  AOI21_X1 U7680 ( .B1(n9346), .B2(n5682), .A(n6154), .ZN(n6156) );
  XNOR2_X1 U7681 ( .A(n6155), .B(n6156), .ZN(n9057) );
  INV_X1 U7682 ( .A(n6155), .ZN(n6157) );
  NAND2_X1 U7683 ( .A1(n4317), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6159) );
  NAND2_X1 U7684 ( .A1(n9341), .A2(n6179), .ZN(n6171) );
  INV_X1 U7685 ( .A(n6162), .ZN(n6160) );
  NAND2_X1 U7686 ( .A1(n6160), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n6181) );
  INV_X1 U7687 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6161) );
  NAND2_X1 U7688 ( .A1(n6162), .A2(n6161), .ZN(n6163) );
  NAND2_X1 U7689 ( .A1(n6181), .A2(n6163), .ZN(n6652) );
  OR2_X1 U7690 ( .A1(n6652), .A2(n5675), .ZN(n6169) );
  INV_X1 U7691 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n6166) );
  NAND2_X1 U7692 ( .A1(n6466), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6165) );
  NAND2_X1 U7693 ( .A1(n5636), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6164) );
  OAI211_X1 U7694 ( .C1(n6468), .C2(n6166), .A(n6165), .B(n6164), .ZN(n6167)
         );
  INV_X1 U7695 ( .A(n6167), .ZN(n6168) );
  NAND2_X1 U7696 ( .A1(n9194), .A2(n5770), .ZN(n6170) );
  NAND2_X1 U7697 ( .A1(n6171), .A2(n6170), .ZN(n6172) );
  XNOR2_X1 U7698 ( .A(n6172), .B(n6191), .ZN(n6226) );
  INV_X1 U7699 ( .A(n6226), .ZN(n6176) );
  NOR2_X1 U7700 ( .A1(n9063), .A2(n6173), .ZN(n6174) );
  AOI21_X1 U7701 ( .B1(n9341), .B2(n5770), .A(n6174), .ZN(n6225) );
  INV_X1 U7702 ( .A(n6225), .ZN(n6175) );
  NAND2_X1 U7703 ( .A1(n6176), .A2(n6175), .ZN(n6648) );
  NAND2_X1 U7704 ( .A1(n8942), .A2(n4318), .ZN(n6178) );
  NAND2_X1 U7705 ( .A1(n4317), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6177) );
  NAND2_X1 U7706 ( .A1(n9336), .A2(n6179), .ZN(n6190) );
  INV_X1 U7707 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6180) );
  NAND2_X1 U7708 ( .A1(n6181), .A2(n6180), .ZN(n6182) );
  NAND2_X1 U7709 ( .A1(n9163), .A2(n6235), .ZN(n6188) );
  INV_X1 U7710 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6185) );
  NAND2_X1 U7711 ( .A1(n6466), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6184) );
  NAND2_X1 U7712 ( .A1(n5636), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6183) );
  OAI211_X1 U7713 ( .C1(n6185), .C2(n6468), .A(n6184), .B(n6183), .ZN(n6186)
         );
  INV_X1 U7714 ( .A(n6186), .ZN(n6187) );
  NAND2_X1 U7715 ( .A1(n9180), .A2(n5770), .ZN(n6189) );
  NAND2_X1 U7716 ( .A1(n6190), .A2(n6189), .ZN(n6192) );
  XNOR2_X1 U7717 ( .A(n6192), .B(n6191), .ZN(n6195) );
  AOI22_X1 U7718 ( .A1(n9336), .A2(n5770), .B1(n6193), .B2(n9180), .ZN(n6194)
         );
  XNOR2_X1 U7719 ( .A(n6195), .B(n6194), .ZN(n6251) );
  INV_X1 U7720 ( .A(n6251), .ZN(n6224) );
  NAND3_X1 U7721 ( .A1(n6196), .A2(P1_B_REG_SCAN_IN), .A3(n7892), .ZN(n6197)
         );
  OAI21_X1 U7722 ( .B1(P1_B_REG_SCAN_IN), .B2(n7892), .A(n6197), .ZN(n6198) );
  NOR4_X1 U7723 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6207) );
  NOR4_X1 U7724 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6206) );
  NOR4_X1 U7725 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6202) );
  NOR4_X1 U7726 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6201) );
  NOR4_X1 U7727 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6200) );
  NOR4_X1 U7728 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6199) );
  NAND4_X1 U7729 ( .A1(n6202), .A2(n6201), .A3(n6200), .A4(n6199), .ZN(n6203)
         );
  NOR4_X1 U7730 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n6204), .A4(n6203), .ZN(n6205) );
  AND3_X1 U7731 ( .A1(n6207), .A2(n6206), .A3(n6205), .ZN(n6208) );
  INV_X1 U7732 ( .A(n6333), .ZN(n6212) );
  INV_X1 U7733 ( .A(n9430), .ZN(n6210) );
  NAND2_X1 U7734 ( .A1(n6210), .A2(n6209), .ZN(n6211) );
  NAND2_X1 U7735 ( .A1(n8015), .A2(n7892), .ZN(n9432) );
  NAND2_X1 U7736 ( .A1(n6212), .A2(n7377), .ZN(n6215) );
  INV_X1 U7737 ( .A(n6196), .ZN(n6213) );
  OAI22_X1 U7738 ( .A1(n9430), .A2(P1_D_REG_1__SCAN_IN), .B1(n6214), .B2(n6213), .ZN(n7149) );
  OR2_X1 U7739 ( .A1(n6215), .A2(n7149), .ZN(n6237) );
  INV_X1 U7740 ( .A(n6237), .ZN(n6244) );
  NAND2_X1 U7741 ( .A1(n6216), .A2(n6217), .ZN(n6659) );
  NAND2_X1 U7742 ( .A1(n4396), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6219) );
  AND2_X1 U7743 ( .A1(n6660), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6220) );
  AND2_X1 U7744 ( .A1(n6659), .A2(n9431), .ZN(n6221) );
  NAND2_X1 U7745 ( .A1(n6244), .A2(n6221), .ZN(n6222) );
  AND2_X1 U7746 ( .A1(n7714), .A2(n7579), .ZN(n7157) );
  INV_X1 U7747 ( .A(n9054), .ZN(n6223) );
  NAND2_X1 U7748 ( .A1(n6226), .A2(n6225), .ZN(n6649) );
  AND2_X1 U7749 ( .A1(n6251), .A2(n4834), .ZN(n6227) );
  NAND2_X1 U7750 ( .A1(n6257), .A2(n6227), .ZN(n6255) );
  AND2_X1 U7751 ( .A1(n6237), .A2(n9431), .ZN(n6228) );
  NAND2_X1 U7752 ( .A1(n4835), .A2(n6228), .ZN(n6247) );
  OR2_X1 U7753 ( .A1(n6659), .A2(n7156), .ZN(n6243) );
  NAND2_X1 U7754 ( .A1(n6243), .A2(n9431), .ZN(n6334) );
  INV_X1 U7755 ( .A(n6334), .ZN(n6229) );
  INV_X1 U7756 ( .A(n6230), .ZN(n8339) );
  INV_X1 U7757 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6233) );
  NAND2_X1 U7758 ( .A1(n6466), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6232) );
  NAND2_X1 U7759 ( .A1(n5636), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6231) );
  OAI211_X1 U7760 ( .C1(n6468), .C2(n6233), .A(n6232), .B(n6231), .ZN(n6234)
         );
  AOI21_X1 U7761 ( .B1(n8339), .B2(n6235), .A(n6234), .ZN(n9071) );
  INV_X1 U7762 ( .A(n9431), .ZN(n6236) );
  NOR2_X1 U7763 ( .A1(n6237), .A2(n6236), .ZN(n6240) );
  INV_X1 U7764 ( .A(n7168), .ZN(n6239) );
  NAND2_X1 U7765 ( .A1(n6240), .A2(n6239), .ZN(n6242) );
  OR2_X1 U7766 ( .A1(n6242), .A2(n6241), .ZN(n9060) );
  NAND2_X1 U7767 ( .A1(n9194), .A2(n9048), .ZN(n6250) );
  AND3_X1 U7768 ( .A1(n6243), .A2(n5625), .A3(n6660), .ZN(n6245) );
  OR2_X1 U7769 ( .A1(n9745), .A2(n6244), .ZN(n6815) );
  NAND2_X1 U7770 ( .A1(n6245), .A2(n6815), .ZN(n6246) );
  NAND2_X1 U7771 ( .A1(n6246), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6248) );
  AOI22_X1 U7772 ( .A1(n9163), .A2(n9066), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n6249) );
  OAI211_X1 U7773 ( .C1(n9071), .C2(n9062), .A(n6250), .B(n6249), .ZN(n6253)
         );
  NOR3_X1 U7774 ( .A1(n6251), .A2(n9054), .A3(n6649), .ZN(n6252) );
  AOI211_X1 U7775 ( .C1(n9052), .C2(n9336), .A(n6253), .B(n6252), .ZN(n6254)
         );
  OAI211_X1 U7776 ( .C1(n6257), .C2(n6256), .A(n6255), .B(n6254), .ZN(P1_U3218) );
  INV_X1 U7777 ( .A(n9363), .ZN(n9242) );
  NAND2_X1 U7778 ( .A1(n6259), .A2(n6304), .ZN(n6260) );
  NAND2_X1 U7779 ( .A1(n7004), .A2(n7006), .ZN(n7003) );
  INV_X1 U7780 ( .A(n5692), .ZN(n7404) );
  NAND2_X1 U7781 ( .A1(n7404), .A2(n6891), .ZN(n6261) );
  NAND2_X1 U7782 ( .A1(n7003), .A2(n6261), .ZN(n7394) );
  INV_X1 U7783 ( .A(n7143), .ZN(n9083) );
  NAND2_X1 U7784 ( .A1(n9083), .A2(n9941), .ZN(n6602) );
  NAND2_X1 U7785 ( .A1(n7143), .A2(n7400), .ZN(n6599) );
  NAND2_X1 U7786 ( .A1(n7394), .A2(n7401), .ZN(n7393) );
  NAND2_X1 U7787 ( .A1(n7143), .A2(n9941), .ZN(n6262) );
  NAND2_X1 U7788 ( .A1(n7393), .A2(n6262), .ZN(n7141) );
  NAND2_X1 U7789 ( .A1(n7403), .A2(n7195), .ZN(n7207) );
  INV_X1 U7790 ( .A(n7403), .ZN(n9082) );
  NAND2_X1 U7791 ( .A1(n9082), .A2(n7160), .ZN(n6603) );
  NAND2_X1 U7792 ( .A1(n7207), .A2(n6603), .ZN(n7144) );
  NAND2_X1 U7793 ( .A1(n7403), .A2(n7160), .ZN(n6263) );
  NAND2_X1 U7794 ( .A1(n7142), .A2(n7227), .ZN(n7272) );
  NAND2_X1 U7795 ( .A1(n9081), .A2(n7216), .ZN(n6361) );
  NAND2_X1 U7796 ( .A1(n9081), .A2(n7227), .ZN(n6265) );
  NAND2_X1 U7797 ( .A1(n7204), .A2(n6265), .ZN(n7269) );
  INV_X1 U7798 ( .A(n7269), .ZN(n6267) );
  NAND2_X1 U7799 ( .A1(n7388), .A2(n7281), .ZN(n6548) );
  INV_X1 U7800 ( .A(n7388), .ZN(n9080) );
  NAND2_X1 U7801 ( .A1(n9080), .A2(n9954), .ZN(n6366) );
  NAND2_X1 U7802 ( .A1(n7388), .A2(n9954), .ZN(n6268) );
  NAND2_X1 U7803 ( .A1(n7271), .A2(n6268), .ZN(n7374) );
  NAND2_X1 U7804 ( .A1(n9960), .A2(n9079), .ZN(n6605) );
  INV_X1 U7805 ( .A(n9079), .ZN(n7262) );
  INV_X1 U7806 ( .A(n9960), .ZN(n7382) );
  NAND2_X1 U7807 ( .A1(n7262), .A2(n7382), .ZN(n7440) );
  NAND2_X1 U7808 ( .A1(n6605), .A2(n7440), .ZN(n7386) );
  NAND2_X1 U7809 ( .A1(n9960), .A2(n7262), .ZN(n6269) );
  OR2_X1 U7810 ( .A1(n7450), .A2(n9917), .ZN(n9910) );
  NAND2_X1 U7811 ( .A1(n7450), .A2(n9917), .ZN(n6374) );
  INV_X1 U7812 ( .A(n9917), .ZN(n9078) );
  NAND2_X1 U7813 ( .A1(n7450), .A2(n9078), .ZN(n6271) );
  NAND2_X1 U7814 ( .A1(n7437), .A2(n6271), .ZN(n9902) );
  AND2_X1 U7815 ( .A1(n9904), .A2(n9077), .ZN(n6272) );
  INV_X1 U7816 ( .A(n9915), .ZN(n9076) );
  OR2_X1 U7817 ( .A1(n9411), .A2(n9729), .ZN(n6385) );
  NAND2_X1 U7818 ( .A1(n9411), .A2(n9729), .ZN(n6387) );
  NAND2_X1 U7819 ( .A1(n6385), .A2(n6387), .ZN(n7861) );
  NAND2_X1 U7820 ( .A1(n7853), .A2(n7861), .ZN(n6274) );
  INV_X1 U7821 ( .A(n9729), .ZN(n9711) );
  NAND2_X1 U7822 ( .A1(n9411), .A2(n9711), .ZN(n6273) );
  OR2_X1 U7823 ( .A1(n9717), .A2(n9074), .ZN(n6275) );
  NAND2_X1 U7824 ( .A1(n9717), .A2(n9074), .ZN(n7917) );
  AND2_X1 U7825 ( .A1(n4374), .A2(n7917), .ZN(n6276) );
  NAND2_X1 U7826 ( .A1(n9401), .A2(n9005), .ZN(n6567) );
  NAND2_X1 U7827 ( .A1(n6400), .A2(n6567), .ZN(n7982) );
  INV_X1 U7828 ( .A(n9005), .ZN(n9072) );
  NAND2_X1 U7829 ( .A1(n9401), .A2(n9072), .ZN(n8016) );
  NAND2_X1 U7830 ( .A1(n9394), .A2(n9320), .ZN(n6278) );
  AND2_X1 U7831 ( .A1(n8016), .A2(n6278), .ZN(n6279) );
  OR2_X1 U7832 ( .A1(n9389), .A2(n6280), .ZN(n6406) );
  NAND2_X1 U7833 ( .A1(n9389), .A2(n6280), .ZN(n6572) );
  NAND2_X1 U7834 ( .A1(n6406), .A2(n6572), .ZN(n9317) );
  OR2_X1 U7835 ( .A1(n9394), .A2(n9320), .ZN(n9304) );
  AND2_X1 U7836 ( .A1(n9317), .A2(n9304), .ZN(n6281) );
  NAND2_X1 U7837 ( .A1(n9389), .A2(n9299), .ZN(n6282) );
  AND2_X1 U7838 ( .A1(n9384), .A2(n9319), .ZN(n6284) );
  NOR2_X1 U7839 ( .A1(n9379), .A2(n9298), .ZN(n6285) );
  NAND2_X1 U7840 ( .A1(n9372), .A2(n9035), .ZN(n6418) );
  NAND2_X1 U7841 ( .A1(n6416), .A2(n6418), .ZN(n9261) );
  NAND2_X1 U7842 ( .A1(n9366), .A2(n9265), .ZN(n6286) );
  INV_X1 U7843 ( .A(n9265), .ZN(n6317) );
  AOI22_X1 U7844 ( .A1(n9245), .A2(n6286), .B1(n6317), .B2(n9251), .ZN(n9229)
         );
  NAND2_X1 U7845 ( .A1(n9351), .A2(n9061), .ZN(n6430) );
  OAI22_X1 U7846 ( .A1(n9199), .A2(n9206), .B1(n9217), .B2(n9351), .ZN(n9185)
         );
  NAND2_X1 U7847 ( .A1(n9346), .A2(n9208), .ZN(n6511) );
  NOR2_X1 U7848 ( .A1(n9346), .A2(n9208), .ZN(n6513) );
  OR2_X1 U7849 ( .A1(n9336), .A2(n6651), .ZN(n6583) );
  NAND2_X1 U7850 ( .A1(n9336), .A2(n6651), .ZN(n6524) );
  NAND2_X1 U7851 ( .A1(n6290), .A2(n6289), .ZN(n6295) );
  INV_X1 U7852 ( .A(n6291), .ZN(n6293) );
  NAND2_X1 U7853 ( .A1(n6293), .A2(n6292), .ZN(n6294) );
  MUX2_X1 U7854 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n6667), .Z(n6447) );
  XNOR2_X1 U7855 ( .A(n6447), .B(n6448), .ZN(n6445) );
  XNOR2_X1 U7856 ( .A(n6446), .B(n6445), .ZN(n8317) );
  NAND2_X1 U7857 ( .A1(n8317), .A2(n4318), .ZN(n6297) );
  NAND2_X1 U7858 ( .A1(n4317), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6296) );
  OR2_X1 U7859 ( .A1(n6443), .A2(n9071), .ZN(n6584) );
  NAND2_X1 U7860 ( .A1(n6443), .A2(n9071), .ZN(n6627) );
  NAND2_X1 U7861 ( .A1(n6584), .A2(n6627), .ZN(n6517) );
  OR2_X1 U7862 ( .A1(n6299), .A2(n7163), .ZN(n6302) );
  OR2_X1 U7863 ( .A1(n6300), .A2(n7579), .ZN(n6301) );
  AND2_X1 U7864 ( .A1(n6302), .A2(n6301), .ZN(n9922) );
  INV_X1 U7865 ( .A(n7175), .ZN(n6303) );
  INV_X1 U7866 ( .A(n7235), .ZN(n7011) );
  NAND2_X1 U7867 ( .A1(n6303), .A2(n7173), .ZN(n6306) );
  INV_X1 U7868 ( .A(n6259), .ZN(n7005) );
  NAND2_X1 U7869 ( .A1(n7005), .A2(n6304), .ZN(n6305) );
  NAND2_X1 U7870 ( .A1(n6306), .A2(n6305), .ZN(n7007) );
  INV_X1 U7871 ( .A(n7006), .ZN(n6493) );
  NAND2_X1 U7872 ( .A1(n7007), .A2(n6493), .ZN(n6308) );
  NAND2_X1 U7873 ( .A1(n7404), .A2(n9329), .ZN(n6307) );
  NAND2_X1 U7874 ( .A1(n6308), .A2(n6307), .ZN(n7402) );
  NAND2_X1 U7875 ( .A1(n7402), .A2(n6602), .ZN(n6555) );
  AND2_X1 U7876 ( .A1(n7272), .A2(n7207), .ZN(n6360) );
  AND2_X1 U7877 ( .A1(n6360), .A2(n6548), .ZN(n6608) );
  INV_X1 U7878 ( .A(n6361), .ZN(n6309) );
  NAND2_X1 U7879 ( .A1(n6548), .A2(n6309), .ZN(n6310) );
  AND2_X1 U7880 ( .A1(n6310), .A2(n6366), .ZN(n6606) );
  OR2_X2 U7881 ( .A1(n7385), .A2(n7386), .ZN(n7441) );
  AND2_X1 U7882 ( .A1(n6374), .A2(n7440), .ZN(n6541) );
  NAND2_X1 U7883 ( .A1(n7441), .A2(n6541), .ZN(n9911) );
  INV_X1 U7884 ( .A(n9077), .ZN(n7315) );
  OR2_X1 U7885 ( .A1(n9904), .A2(n7315), .ZN(n9901) );
  AND2_X1 U7886 ( .A1(n9901), .A2(n9910), .ZN(n6556) );
  NAND2_X1 U7887 ( .A1(n9911), .A2(n6556), .ZN(n7609) );
  INV_X1 U7888 ( .A(n6557), .ZN(n6311) );
  NAND2_X1 U7889 ( .A1(n9904), .A2(n7315), .ZN(n9900) );
  NAND2_X1 U7890 ( .A1(n6377), .A2(n9900), .ZN(n6368) );
  NAND2_X1 U7891 ( .A1(n6368), .A2(n6557), .ZN(n6538) );
  OAI21_X2 U7892 ( .B1(n7609), .B2(n6311), .A(n6538), .ZN(n9728) );
  INV_X1 U7893 ( .A(n9075), .ZN(n7826) );
  AND2_X1 U7894 ( .A1(n9759), .A2(n7826), .ZN(n6383) );
  OR2_X1 U7895 ( .A1(n9759), .A2(n7826), .ZN(n7859) );
  AND2_X1 U7896 ( .A1(n6385), .A2(n7859), .ZN(n6388) );
  INV_X1 U7897 ( .A(n9074), .ZN(n6312) );
  OR2_X1 U7898 ( .A1(n9717), .A2(n6312), .ZN(n6391) );
  NAND2_X1 U7899 ( .A1(n9717), .A2(n6312), .ZN(n6540) );
  INV_X1 U7900 ( .A(n6540), .ZN(n6558) );
  INV_X1 U7901 ( .A(n9708), .ZN(n8042) );
  NAND2_X1 U7902 ( .A1(n9407), .A2(n8042), .ZN(n6563) );
  NAND2_X1 U7903 ( .A1(n7919), .A2(n6392), .ZN(n7956) );
  NAND2_X1 U7904 ( .A1(n8048), .A2(n8991), .ZN(n6564) );
  NAND2_X1 U7905 ( .A1(n7956), .A2(n6564), .ZN(n7981) );
  OR2_X1 U7906 ( .A1(n8048), .A2(n8991), .ZN(n7980) );
  NAND2_X1 U7907 ( .A1(n7981), .A2(n6569), .ZN(n6313) );
  INV_X1 U7908 ( .A(n9320), .ZN(n6314) );
  AND2_X1 U7909 ( .A1(n9394), .A2(n6314), .ZN(n6546) );
  OR2_X1 U7910 ( .A1(n9394), .A2(n6314), .ZN(n9315) );
  AND2_X1 U7911 ( .A1(n6406), .A2(n9315), .ZN(n6531) );
  INV_X1 U7912 ( .A(n9319), .ZN(n9046) );
  OR2_X1 U7913 ( .A1(n9384), .A2(n9046), .ZN(n6409) );
  NAND2_X1 U7914 ( .A1(n9384), .A2(n9046), .ZN(n6528) );
  NAND2_X1 U7915 ( .A1(n9297), .A2(n9296), .ZN(n6315) );
  INV_X1 U7916 ( .A(n9298), .ZN(n8972) );
  OR2_X1 U7917 ( .A1(n9379), .A2(n8972), .ZN(n6490) );
  INV_X1 U7918 ( .A(n6418), .ZN(n6316) );
  NAND2_X1 U7919 ( .A1(n9366), .A2(n6317), .ZN(n6421) );
  NAND2_X1 U7920 ( .A1(n9363), .A2(n9038), .ZN(n6616) );
  NAND2_X1 U7921 ( .A1(n6577), .A2(n6616), .ZN(n9228) );
  INV_X1 U7922 ( .A(n6577), .ZN(n6351) );
  NOR2_X1 U7923 ( .A1(n9235), .A2(n6351), .ZN(n9216) );
  XNOR2_X1 U7924 ( .A(n9357), .B(n9233), .ZN(n9215) );
  NAND2_X1 U7925 ( .A1(n9216), .A2(n9215), .ZN(n9214) );
  NAND2_X1 U7926 ( .A1(n9357), .A2(n6349), .ZN(n9205) );
  INV_X1 U7927 ( .A(n6525), .ZN(n6318) );
  INV_X1 U7928 ( .A(n9208), .ZN(n8980) );
  OR2_X1 U7929 ( .A1(n9346), .A2(n8980), .ZN(n6526) );
  NAND3_X1 U7930 ( .A1(n9167), .A2(n9169), .A3(n9166), .ZN(n9168) );
  NAND2_X1 U7931 ( .A1(n9168), .A2(n6524), .ZN(n6319) );
  NAND2_X1 U7932 ( .A1(n6216), .A2(n9272), .ZN(n6321) );
  NAND2_X1 U7933 ( .A1(n6217), .A2(n6639), .ZN(n6320) );
  INV_X1 U7934 ( .A(n6659), .ZN(n6322) );
  INV_X1 U7935 ( .A(n6323), .ZN(n6643) );
  AND2_X1 U7936 ( .A1(n6643), .A2(P1_B_REG_SCAN_IN), .ZN(n6324) );
  NOR2_X1 U7937 ( .A1(n9914), .A2(n6324), .ZN(n9148) );
  INV_X1 U7938 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n6327) );
  NAND2_X1 U7939 ( .A1(n6466), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6326) );
  NAND2_X1 U7940 ( .A1(n5636), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6325) );
  OAI211_X1 U7941 ( .C1(n6468), .C2(n6327), .A(n6326), .B(n6325), .ZN(n9070)
         );
  INV_X1 U7942 ( .A(n9346), .ZN(n9191) );
  NAND2_X1 U7943 ( .A1(n7154), .A2(n7160), .ZN(n7214) );
  OR2_X1 U7944 ( .A1(n7214), .A2(n7227), .ZN(n7280) );
  NOR2_X2 U7945 ( .A1(n7280), .A2(n7281), .ZN(n7375) );
  AND2_X1 U7946 ( .A1(n7375), .A2(n9960), .ZN(n7448) );
  INV_X1 U7947 ( .A(n7450), .ZN(n7447) );
  NAND2_X1 U7948 ( .A1(n7448), .A2(n7447), .ZN(n9903) );
  OR2_X1 U7949 ( .A1(n9905), .A2(n9660), .ZN(n9721) );
  INV_X1 U7950 ( .A(n9411), .ZN(n7858) );
  INV_X1 U7951 ( .A(n9717), .ZN(n9752) );
  INV_X1 U7952 ( .A(n9407), .ZN(n7929) );
  OR2_X2 U7953 ( .A1(n7960), .A2(n8048), .ZN(n7976) );
  INV_X1 U7954 ( .A(n9394), .ZN(n9010) );
  INV_X1 U7955 ( .A(n9389), .ZN(n9314) );
  NOR2_X2 U7956 ( .A1(n9291), .A2(n9379), .ZN(n9278) );
  INV_X1 U7957 ( .A(n9372), .ZN(n9268) );
  NAND2_X1 U7958 ( .A1(n9269), .A2(n9251), .ZN(n9246) );
  NOR2_X2 U7959 ( .A1(n9341), .A2(n9186), .ZN(n9175) );
  INV_X1 U7960 ( .A(n9336), .ZN(n9165) );
  NAND2_X1 U7961 ( .A1(n9175), .A2(n9165), .ZN(n9160) );
  AOI21_X1 U7962 ( .B1(n6443), .B2(n9160), .A(n9154), .ZN(n8338) );
  AOI22_X1 U7963 ( .A1(n8338), .A2(n9395), .B1(n9745), .B2(n6443), .ZN(n6331)
         );
  OAI21_X1 U7964 ( .B1(n9659), .B2(n6217), .A(n7149), .ZN(n6335) );
  NAND2_X1 U7965 ( .A1(n6340), .A2(n9990), .ZN(n6338) );
  INV_X1 U7966 ( .A(n9990), .ZN(n6336) );
  NAND2_X1 U7967 ( .A1(n6338), .A2(n6337), .ZN(P1_U3552) );
  NAND2_X1 U7968 ( .A1(n6340), .A2(n9980), .ZN(n6343) );
  INV_X1 U7969 ( .A(n9980), .ZN(n6341) );
  NAND2_X1 U7970 ( .A1(n6341), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6342) );
  NAND2_X1 U7971 ( .A1(n6343), .A2(n6342), .ZN(P1_U3520) );
  NAND2_X1 U7972 ( .A1(n9346), .A2(n6525), .ZN(n6344) );
  NAND2_X1 U7973 ( .A1(n6523), .A2(n6344), .ZN(n6347) );
  NAND2_X1 U7974 ( .A1(n6430), .A2(n9208), .ZN(n6345) );
  NAND2_X1 U7975 ( .A1(n9166), .A2(n6345), .ZN(n6346) );
  MUX2_X1 U7976 ( .A(n6347), .B(n6346), .S(n6478), .Z(n6348) );
  INV_X1 U7977 ( .A(n6348), .ZN(n6436) );
  NOR2_X1 U7978 ( .A1(n9357), .A2(n6349), .ZN(n6415) );
  OAI21_X1 U7979 ( .B1(n6415), .B2(n6616), .A(n6621), .ZN(n6350) );
  INV_X1 U7980 ( .A(n6478), .ZN(n6483) );
  NAND2_X1 U7981 ( .A1(n6350), .A2(n6483), .ZN(n6428) );
  NAND2_X1 U7982 ( .A1(n9205), .A2(n6351), .ZN(n6352) );
  NAND2_X1 U7983 ( .A1(n6525), .A2(n6352), .ZN(n6427) );
  NAND2_X1 U7984 ( .A1(n6415), .A2(n6478), .ZN(n6425) );
  NAND2_X1 U7985 ( .A1(n6416), .A2(n6491), .ZN(n6353) );
  AND2_X1 U7986 ( .A1(n6353), .A2(n6418), .ZN(n6354) );
  NAND2_X1 U7987 ( .A1(n6354), .A2(n6421), .ZN(n6533) );
  OR2_X1 U7988 ( .A1(n6533), .A2(n6416), .ZN(n6356) );
  INV_X1 U7989 ( .A(n6489), .ZN(n6355) );
  AND2_X1 U7990 ( .A1(n6356), .A2(n6355), .ZN(n6535) );
  INV_X1 U7991 ( .A(n6533), .ZN(n6412) );
  INV_X1 U7992 ( .A(n6546), .ZN(n6570) );
  AND2_X1 U7993 ( .A1(n6572), .A2(n6570), .ZN(n6357) );
  MUX2_X1 U7994 ( .A(n6357), .B(n6531), .S(n6478), .Z(n6405) );
  NAND2_X1 U7995 ( .A1(n6567), .A2(n6564), .ZN(n6544) );
  INV_X1 U7996 ( .A(n7207), .ZN(n6358) );
  OR2_X1 U7997 ( .A1(n7145), .A2(n6358), .ZN(n6359) );
  MUX2_X1 U7998 ( .A(n6359), .B(n7208), .S(n6478), .Z(n6365) );
  AND2_X1 U7999 ( .A1(n6603), .A2(n6361), .ZN(n6495) );
  MUX2_X1 U8000 ( .A(n6495), .B(n6360), .S(n6478), .Z(n6364) );
  MUX2_X1 U8001 ( .A(n6361), .B(n7272), .S(n6483), .Z(n6362) );
  NAND2_X1 U8002 ( .A1(n6362), .A2(n7274), .ZN(n6363) );
  AOI21_X1 U8003 ( .B1(n6365), .B2(n6364), .A(n6363), .ZN(n6373) );
  NAND2_X1 U8004 ( .A1(n6605), .A2(n6366), .ZN(n6499) );
  OAI21_X1 U8005 ( .B1(n6373), .B2(n6499), .A(n6541), .ZN(n6367) );
  NAND2_X1 U8006 ( .A1(n6367), .A2(n6556), .ZN(n6371) );
  INV_X1 U8007 ( .A(n6368), .ZN(n6370) );
  NAND2_X1 U8008 ( .A1(n6385), .A2(n6557), .ZN(n6369) );
  AOI21_X1 U8009 ( .B1(n6371), .B2(n6370), .A(n6369), .ZN(n6381) );
  NAND2_X1 U8010 ( .A1(n6548), .A2(n7440), .ZN(n6372) );
  OAI211_X1 U8011 ( .C1(n6373), .C2(n6372), .A(n6556), .B(n6605), .ZN(n6376)
         );
  NAND2_X1 U8012 ( .A1(n9900), .A2(n6374), .ZN(n6498) );
  NAND2_X1 U8013 ( .A1(n6498), .A2(n9901), .ZN(n6375) );
  NAND2_X1 U8014 ( .A1(n6376), .A2(n6375), .ZN(n6379) );
  INV_X1 U8015 ( .A(n6377), .ZN(n6378) );
  AOI21_X1 U8016 ( .B1(n6379), .B2(n6557), .A(n6378), .ZN(n6380) );
  MUX2_X1 U8017 ( .A(n6381), .B(n6380), .S(n6478), .Z(n6382) );
  XNOR2_X1 U8018 ( .A(n9759), .B(n9075), .ZN(n6502) );
  NAND3_X1 U8019 ( .A1(n6382), .A2(n6387), .A3(n6502), .ZN(n6399) );
  NAND2_X1 U8020 ( .A1(n6563), .A2(n6540), .ZN(n6393) );
  INV_X1 U8021 ( .A(n6383), .ZN(n6384) );
  NAND2_X1 U8022 ( .A1(n6387), .A2(n6384), .ZN(n6537) );
  NAND2_X1 U8023 ( .A1(n6537), .A2(n6385), .ZN(n6386) );
  NAND2_X1 U8024 ( .A1(n6386), .A2(n6483), .ZN(n6390) );
  OR2_X1 U8025 ( .A1(n6388), .A2(n4604), .ZN(n6559) );
  NAND4_X1 U8026 ( .A1(n6392), .A2(n6391), .A3(n6559), .A4(n6478), .ZN(n6389)
         );
  OAI21_X1 U8027 ( .B1(n6393), .B2(n6390), .A(n6389), .ZN(n6398) );
  NAND2_X1 U8028 ( .A1(n7980), .A2(n6564), .ZN(n7954) );
  NAND2_X1 U8029 ( .A1(n6392), .A2(n6391), .ZN(n6565) );
  NAND3_X1 U8030 ( .A1(n6565), .A2(n6483), .A3(n6563), .ZN(n6395) );
  NAND3_X1 U8031 ( .A1(n6393), .A2(n6392), .A3(n6478), .ZN(n6394) );
  NAND2_X1 U8032 ( .A1(n6395), .A2(n6394), .ZN(n6396) );
  OR2_X1 U8033 ( .A1(n7954), .A2(n6396), .ZN(n6397) );
  AOI21_X1 U8034 ( .B1(n6399), .B2(n6398), .A(n6397), .ZN(n6402) );
  MUX2_X1 U8035 ( .A(n6400), .B(n6567), .S(n6478), .Z(n6401) );
  OAI211_X1 U8036 ( .C1(n6403), .C2(n6402), .A(n8022), .B(n6401), .ZN(n6404)
         );
  NAND2_X1 U8037 ( .A1(n6405), .A2(n6404), .ZN(n6410) );
  NAND3_X1 U8038 ( .A1(n6410), .A2(n6406), .A3(n6409), .ZN(n6408) );
  INV_X1 U8039 ( .A(n6491), .ZN(n6407) );
  AND2_X1 U8040 ( .A1(n6490), .A2(n6409), .ZN(n6532) );
  NAND3_X1 U8041 ( .A1(n6410), .A2(n6572), .A3(n6528), .ZN(n6411) );
  NAND2_X1 U8042 ( .A1(n6412), .A2(n6417), .ZN(n6413) );
  NAND2_X1 U8043 ( .A1(n6535), .A2(n6413), .ZN(n6414) );
  NAND4_X1 U8044 ( .A1(n6414), .A2(n9205), .A3(n6616), .A4(n6478), .ZN(n6424)
         );
  INV_X1 U8045 ( .A(n9228), .ZN(n9231) );
  NOR2_X1 U8046 ( .A1(n6489), .A2(n6478), .ZN(n6420) );
  INV_X1 U8047 ( .A(n6415), .ZN(n6578) );
  NAND4_X1 U8048 ( .A1(n9231), .A2(n6420), .A3(n6578), .A4(n6419), .ZN(n6423)
         );
  INV_X1 U8049 ( .A(n6421), .ZN(n6488) );
  NAND4_X1 U8050 ( .A1(n6578), .A2(n6488), .A3(n6483), .A4(n6577), .ZN(n6422)
         );
  NAND4_X1 U8051 ( .A1(n6425), .A2(n6424), .A3(n6423), .A4(n6422), .ZN(n6426)
         );
  NOR2_X1 U8052 ( .A1(n6430), .A2(n9208), .ZN(n6431) );
  OR2_X1 U8053 ( .A1(n6431), .A2(n9346), .ZN(n6434) );
  AND2_X1 U8054 ( .A1(n6525), .A2(n8980), .ZN(n6432) );
  NOR2_X1 U8055 ( .A1(n6521), .A2(n6432), .ZN(n6433) );
  MUX2_X1 U8056 ( .A(n6434), .B(n6433), .S(n6483), .Z(n6435) );
  OAI22_X1 U8057 ( .A1(n6436), .A2(n4832), .B1(n4376), .B2(n6435), .ZN(n6438)
         );
  MUX2_X1 U8058 ( .A(n9166), .B(n6523), .S(n6478), .Z(n6437) );
  NAND3_X1 U8059 ( .A1(n6438), .A2(n9169), .A3(n6437), .ZN(n6440) );
  MUX2_X1 U8060 ( .A(n6524), .B(n6583), .S(n6478), .Z(n6439) );
  INV_X1 U8061 ( .A(n6443), .ZN(n8342) );
  NOR2_X1 U8062 ( .A1(n9071), .A2(n6483), .ZN(n6441) );
  AOI21_X1 U8063 ( .B1(n6443), .B2(n6483), .A(n6441), .ZN(n6442) );
  NAND2_X1 U8064 ( .A1(n6446), .A2(n6445), .ZN(n6451) );
  INV_X1 U8065 ( .A(n6447), .ZN(n6449) );
  NAND2_X1 U8066 ( .A1(n6449), .A2(n6448), .ZN(n6450) );
  MUX2_X1 U8067 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n6667), .Z(n6456) );
  INV_X1 U8068 ( .A(SI_30_), .ZN(n9595) );
  XNOR2_X1 U8069 ( .A(n6456), .B(n9595), .ZN(n6454) );
  XNOR2_X1 U8070 ( .A(n6455), .B(n6454), .ZN(n8071) );
  NAND2_X1 U8071 ( .A1(n8071), .A2(n5685), .ZN(n6453) );
  NAND2_X1 U8072 ( .A1(n4317), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n6452) );
  INV_X1 U8073 ( .A(n9070), .ZN(n6479) );
  NOR2_X1 U8074 ( .A1(n9744), .A2(n6479), .ZN(n6487) );
  NAND2_X1 U8075 ( .A1(n6455), .A2(n6454), .ZN(n6459) );
  INV_X1 U8076 ( .A(n6456), .ZN(n6457) );
  NAND2_X1 U8077 ( .A1(n6457), .A2(n9595), .ZN(n6458) );
  NAND2_X1 U8078 ( .A1(n6459), .A2(n6458), .ZN(n6463) );
  MUX2_X1 U8079 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n6667), .Z(n6461) );
  INV_X1 U8080 ( .A(SI_31_), .ZN(n6460) );
  XNOR2_X1 U8081 ( .A(n6461), .B(n6460), .ZN(n6462) );
  NAND2_X1 U8082 ( .A1(n8933), .A2(n4318), .ZN(n6465) );
  NAND2_X1 U8083 ( .A1(n4317), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n6464) );
  NAND2_X1 U8084 ( .A1(n6487), .A2(n9671), .ZN(n6474) );
  NAND2_X1 U8085 ( .A1(n6466), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6473) );
  INV_X1 U8086 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6467) );
  OR2_X1 U8087 ( .A1(n6468), .A2(n6467), .ZN(n6472) );
  INV_X1 U8088 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6469) );
  OR2_X1 U8089 ( .A1(n6470), .A2(n6469), .ZN(n6471) );
  NAND2_X1 U8090 ( .A1(n9671), .A2(n9149), .ZN(n6635) );
  AND2_X1 U8091 ( .A1(n6474), .A2(n6635), .ZN(n6482) );
  NOR2_X1 U8092 ( .A1(n9071), .A2(n6478), .ZN(n6475) );
  AOI22_X1 U8093 ( .A1(n6477), .A2(n6482), .B1(n6476), .B2(n6475), .ZN(n6481)
         );
  NAND2_X1 U8094 ( .A1(n9744), .A2(n6479), .ZN(n6632) );
  NAND2_X1 U8095 ( .A1(n9744), .A2(n9149), .ZN(n6480) );
  NAND2_X1 U8096 ( .A1(n6632), .A2(n6480), .ZN(n6586) );
  INV_X1 U8097 ( .A(n6482), .ZN(n6588) );
  NAND2_X1 U8098 ( .A1(n6588), .A2(n6483), .ZN(n6484) );
  OAI21_X1 U8099 ( .B1(n6216), .B2(n7579), .A(n6486), .ZN(n6485) );
  INV_X1 U8100 ( .A(n6487), .ZN(n6630) );
  AND2_X1 U8101 ( .A1(n6630), .A2(n6632), .ZN(n6519) );
  NOR2_X1 U8102 ( .A1(n6489), .A2(n6488), .ZN(n9253) );
  INV_X1 U8103 ( .A(n6490), .ZN(n6492) );
  INV_X1 U8104 ( .A(n9317), .ZN(n6508) );
  AND2_X1 U8105 ( .A1(n6258), .A2(n7011), .ZN(n6594) );
  NOR2_X1 U8106 ( .A1(n7173), .A2(n6594), .ZN(n6804) );
  INV_X1 U8107 ( .A(n7401), .ZN(n6494) );
  AND3_X1 U8108 ( .A1(n6804), .A2(n6494), .A3(n6493), .ZN(n6497) );
  INV_X1 U8109 ( .A(n6495), .ZN(n6549) );
  NOR2_X1 U8110 ( .A1(n7175), .A2(n6549), .ZN(n6496) );
  AND4_X1 U8111 ( .A1(n6497), .A2(n6608), .A3(n6496), .A4(n7440), .ZN(n6501)
         );
  INV_X1 U8112 ( .A(n6498), .ZN(n6500) );
  INV_X1 U8113 ( .A(n6499), .ZN(n6551) );
  NAND4_X1 U8114 ( .A1(n6501), .A2(n6556), .A3(n6500), .A4(n6551), .ZN(n6503)
         );
  INV_X1 U8115 ( .A(n6502), .ZN(n9727) );
  NOR4_X1 U8116 ( .A1(n7861), .A2(n6503), .A3(n9727), .A4(n7610), .ZN(n6504)
         );
  NAND3_X1 U8117 ( .A1(n7920), .A2(n9705), .A3(n6504), .ZN(n6505) );
  OR2_X1 U8118 ( .A1(n7954), .A2(n6505), .ZN(n6506) );
  NOR2_X1 U8119 ( .A1(n7982), .A2(n6506), .ZN(n6507) );
  NAND4_X1 U8120 ( .A1(n9296), .A2(n8022), .A3(n6508), .A4(n6507), .ZN(n6509)
         );
  NOR3_X1 U8121 ( .A1(n9261), .A2(n9284), .A3(n6509), .ZN(n6510) );
  AND4_X1 U8122 ( .A1(n9206), .A2(n9231), .A3(n9253), .A4(n6510), .ZN(n6514)
         );
  INV_X1 U8123 ( .A(n6511), .ZN(n6512) );
  AND4_X1 U8124 ( .A1(n9179), .A2(n6514), .A3(n9215), .A4(n9192), .ZN(n6515)
         );
  NAND2_X1 U8125 ( .A1(n9169), .A2(n6515), .ZN(n6516) );
  NOR2_X1 U8126 ( .A1(n6517), .A2(n6516), .ZN(n6518) );
  NAND4_X1 U8127 ( .A1(n6633), .A2(n6635), .A3(n6519), .A4(n6518), .ZN(n6520)
         );
  NAND2_X1 U8128 ( .A1(n6520), .A2(n7579), .ZN(n6592) );
  NAND2_X1 U8129 ( .A1(n9166), .A2(n6521), .ZN(n6522) );
  NAND3_X1 U8130 ( .A1(n6524), .A2(n6523), .A3(n6522), .ZN(n6626) );
  AND2_X1 U8131 ( .A1(n6526), .A2(n6525), .ZN(n6527) );
  NAND2_X1 U8132 ( .A1(n9166), .A2(n6527), .ZN(n6624) );
  INV_X1 U8133 ( .A(n6528), .ZN(n6529) );
  OR2_X1 U8134 ( .A1(n6533), .A2(n6529), .ZN(n6615) );
  INV_X1 U8135 ( .A(n6572), .ZN(n6530) );
  OR2_X1 U8136 ( .A1(n6531), .A2(n6530), .ZN(n6536) );
  OR2_X1 U8137 ( .A1(n6533), .A2(n6532), .ZN(n6534) );
  OAI211_X1 U8138 ( .C1(n6615), .C2(n6536), .A(n6535), .B(n6534), .ZN(n6618)
         );
  INV_X1 U8139 ( .A(n6537), .ZN(n6539) );
  NAND3_X1 U8140 ( .A1(n6540), .A2(n6539), .A3(n6538), .ZN(n6562) );
  INV_X1 U8141 ( .A(n6562), .ZN(n6542) );
  NAND3_X1 U8142 ( .A1(n6542), .A2(n6541), .A3(n6563), .ZN(n6543) );
  OR2_X1 U8143 ( .A1(n6544), .A2(n6543), .ZN(n6545) );
  NOR2_X1 U8144 ( .A1(n6546), .A2(n6545), .ZN(n6547) );
  NAND2_X1 U8145 ( .A1(n6572), .A2(n6547), .ZN(n6612) );
  NAND3_X1 U8146 ( .A1(n6606), .A2(n6603), .A3(n6605), .ZN(n6554) );
  NAND2_X1 U8147 ( .A1(n6608), .A2(n6599), .ZN(n6552) );
  NAND3_X1 U8148 ( .A1(n6549), .A2(n6548), .A3(n7272), .ZN(n6550) );
  NAND3_X1 U8149 ( .A1(n6552), .A2(n6551), .A3(n6550), .ZN(n6553) );
  OAI21_X1 U8150 ( .B1(n6555), .B2(n6554), .A(n6553), .ZN(n6573) );
  AND2_X1 U8151 ( .A1(n6557), .A2(n6556), .ZN(n6561) );
  OR2_X1 U8152 ( .A1(n6559), .A2(n6558), .ZN(n6560) );
  OAI21_X1 U8153 ( .B1(n6562), .B2(n6561), .A(n6560), .ZN(n6566) );
  OAI211_X1 U8154 ( .C1(n6566), .C2(n6565), .A(n6564), .B(n6563), .ZN(n6568)
         );
  AOI21_X1 U8155 ( .B1(n6569), .B2(n6568), .A(n4605), .ZN(n6571) );
  NAND3_X1 U8156 ( .A1(n6572), .A2(n6571), .A3(n6570), .ZN(n6610) );
  OAI21_X1 U8157 ( .B1(n6612), .B2(n6573), .A(n6610), .ZN(n6574) );
  INV_X1 U8158 ( .A(n6574), .ZN(n6575) );
  NOR2_X1 U8159 ( .A1(n6615), .A2(n6575), .ZN(n6576) );
  OAI21_X1 U8160 ( .B1(n6618), .B2(n6576), .A(n6616), .ZN(n6579) );
  AND2_X1 U8161 ( .A1(n6578), .A2(n6577), .ZN(n6619) );
  NAND2_X1 U8162 ( .A1(n6579), .A2(n6619), .ZN(n6580) );
  AND2_X1 U8163 ( .A1(n6580), .A2(n6621), .ZN(n6581) );
  NOR2_X1 U8164 ( .A1(n6624), .A2(n6581), .ZN(n6582) );
  NOR2_X1 U8165 ( .A1(n6626), .A2(n6582), .ZN(n6585) );
  NAND2_X1 U8166 ( .A1(n6584), .A2(n6583), .ZN(n6628) );
  OAI21_X1 U8167 ( .B1(n6585), .B2(n6628), .A(n6627), .ZN(n6587) );
  NOR2_X1 U8168 ( .A1(n6587), .A2(n6586), .ZN(n6589) );
  OAI211_X1 U8169 ( .C1(n6589), .C2(n6588), .A(n6217), .B(n6633), .ZN(n6590)
         );
  NAND2_X1 U8170 ( .A1(n6590), .A2(n6592), .ZN(n6591) );
  MUX2_X1 U8171 ( .A(n6592), .B(n6591), .S(n9222), .Z(n6593) );
  AOI21_X1 U8172 ( .B1(n6259), .B2(n9936), .A(n7579), .ZN(n6596) );
  INV_X1 U8173 ( .A(n6594), .ZN(n6595) );
  AND2_X1 U8174 ( .A1(n6596), .A2(n6595), .ZN(n6597) );
  OR2_X1 U8175 ( .A1(n7007), .A2(n6597), .ZN(n6598) );
  AOI21_X1 U8176 ( .B1(n6598), .B2(n9329), .A(n7404), .ZN(n6601) );
  NOR2_X1 U8177 ( .A1(n6598), .A2(n9329), .ZN(n6600) );
  OAI21_X1 U8178 ( .B1(n6601), .B2(n6600), .A(n6599), .ZN(n6604) );
  NAND3_X1 U8179 ( .A1(n6604), .A2(n6603), .A3(n6602), .ZN(n6609) );
  NAND2_X1 U8180 ( .A1(n6606), .A2(n6605), .ZN(n6607) );
  AOI21_X1 U8181 ( .B1(n6609), .B2(n6608), .A(n6607), .ZN(n6611) );
  OAI21_X1 U8182 ( .B1(n6612), .B2(n6611), .A(n6610), .ZN(n6613) );
  INV_X1 U8183 ( .A(n6613), .ZN(n6614) );
  NOR2_X1 U8184 ( .A1(n6615), .A2(n6614), .ZN(n6617) );
  OAI21_X1 U8185 ( .B1(n6618), .B2(n6617), .A(n6616), .ZN(n6620) );
  NAND2_X1 U8186 ( .A1(n6620), .A2(n6619), .ZN(n6622) );
  AND2_X1 U8187 ( .A1(n6622), .A2(n6621), .ZN(n6623) );
  NOR2_X1 U8188 ( .A1(n6624), .A2(n6623), .ZN(n6625) );
  NOR2_X1 U8189 ( .A1(n6626), .A2(n6625), .ZN(n6629) );
  OAI21_X1 U8190 ( .B1(n6629), .B2(n6628), .A(n6627), .ZN(n6631) );
  NAND2_X1 U8191 ( .A1(n6631), .A2(n6630), .ZN(n6634) );
  NAND3_X1 U8192 ( .A1(n6634), .A2(n6633), .A3(n6632), .ZN(n6636) );
  NAND2_X1 U8193 ( .A1(n6636), .A2(n6635), .ZN(n6637) );
  OR2_X1 U8194 ( .A1(n6637), .A2(n9222), .ZN(n6640) );
  OR2_X1 U8195 ( .A1(n6660), .A2(n10130), .ZN(n7818) );
  AOI21_X1 U8196 ( .B1(n6637), .B2(n7156), .A(n7818), .ZN(n6638) );
  NAND3_X1 U8197 ( .A1(n9431), .A2(n6727), .A3(n6643), .ZN(n6644) );
  NOR2_X1 U8198 ( .A1(n7168), .A2(n6644), .ZN(n6646) );
  OAI21_X1 U8199 ( .B1(n6216), .B2(n7818), .A(P1_B_REG_SCAN_IN), .ZN(n6645) );
  OR2_X1 U8200 ( .A1(n6646), .A2(n6645), .ZN(n6647) );
  XNOR2_X1 U8201 ( .A(n6650), .B(n4833), .ZN(n6657) );
  NOR2_X1 U8202 ( .A1(n6651), .A2(n9062), .ZN(n6655) );
  INV_X1 U8203 ( .A(n6652), .ZN(n9176) );
  AOI22_X1 U8204 ( .A1(n9176), .A2(n9066), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n6653) );
  OAI21_X1 U8205 ( .B1(n8980), .B2(n9060), .A(n6653), .ZN(n6654) );
  AOI211_X1 U8206 ( .C1(n9341), .C2(n9052), .A(n6655), .B(n6654), .ZN(n6656)
         );
  OAI21_X1 U8207 ( .B1(n6657), .B2(n9054), .A(n6656), .ZN(P1_U3212) );
  INV_X1 U8208 ( .A(n6660), .ZN(n6658) );
  NAND2_X1 U8209 ( .A1(n6659), .A2(n5625), .ZN(n6661) );
  NAND2_X1 U8210 ( .A1(n6661), .A2(n6660), .ZN(n6719) );
  NAND2_X1 U8211 ( .A1(n6719), .A2(n6662), .ZN(n9783) );
  NAND2_X1 U8212 ( .A1(n9783), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U8213 ( .A(n6833), .ZN(n6663) );
  XNOR2_X1 U8214 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U8215 ( .A(n6664), .ZN(n6665) );
  NAND2_X1 U8216 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_STATE_REG_SCAN_IN), .ZN(
        n9777) );
  OAI21_X1 U8217 ( .B1(n6665), .B2(P1_STATE_REG_SCAN_IN), .A(n9777), .ZN(
        P1_U3353) );
  INV_X1 U8218 ( .A(n8943), .ZN(n8947) );
  INV_X1 U8219 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6666) );
  OR2_X2 U8220 ( .A1(n6667), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8946) );
  OAI222_X1 U8221 ( .A1(n8947), .A2(n6666), .B1(n8946), .B2(n6669), .C1(
        P2_U3152), .C2(n4547), .ZN(P2_U3356) );
  INV_X1 U8222 ( .A(n8318), .ZN(n9441) );
  AOI22_X1 U8223 ( .A1(n9441), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n9811), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6668) );
  OAI21_X1 U8224 ( .B1(n6669), .B2(n9443), .A(n6668), .ZN(P1_U3351) );
  AOI22_X1 U8225 ( .A1(n6748), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n9441), .ZN(n6670) );
  OAI21_X1 U8226 ( .B1(n6678), .B2(n9443), .A(n6670), .ZN(P1_U3350) );
  OAI222_X1 U8227 ( .A1(n8947), .A2(n4905), .B1(n8946), .B2(n6672), .C1(
        P2_U3152), .C2(n6905), .ZN(P2_U3354) );
  INV_X1 U8228 ( .A(n9830), .ZN(n6751) );
  INV_X1 U8229 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6671) );
  OAI222_X1 U8230 ( .A1(n6751), .A2(P1_U3084), .B1(n9443), .B2(n6672), .C1(
        n6671), .C2(n8318), .ZN(P1_U3349) );
  INV_X1 U8231 ( .A(n6673), .ZN(n6676) );
  INV_X1 U8232 ( .A(n9849), .ZN(n6674) );
  OAI222_X1 U8233 ( .A1(n8318), .A2(n6675), .B1(n9443), .B2(n6676), .C1(n6674), 
        .C2(P1_U3084), .ZN(P1_U3348) );
  INV_X1 U8234 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6677) );
  OAI222_X1 U8235 ( .A1(n8947), .A2(n6677), .B1(n8946), .B2(n6676), .C1(
        P2_U3152), .C2(n6912), .ZN(P2_U3353) );
  INV_X1 U8236 ( .A(n6858), .ZN(n6879) );
  OAI222_X1 U8237 ( .A1(n8947), .A2(n4899), .B1(n8946), .B2(n6678), .C1(
        P2_U3152), .C2(n6879), .ZN(P2_U3355) );
  INV_X1 U8238 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6679) );
  OAI222_X1 U8239 ( .A1(n8947), .A2(n6679), .B1(n8946), .B2(n8054), .C1(
        P2_U3152), .C2(n6855), .ZN(P2_U3357) );
  INV_X1 U8240 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6682) );
  INV_X1 U8241 ( .A(n7149), .ZN(n6680) );
  NAND2_X1 U8242 ( .A1(n6680), .A2(n9431), .ZN(n6681) );
  OAI21_X1 U8243 ( .B1(n9431), .B2(n6682), .A(n6681), .ZN(P1_U3441) );
  INV_X1 U8244 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6684) );
  INV_X1 U8245 ( .A(n6683), .ZN(n6686) );
  INV_X1 U8246 ( .A(n6934), .ZN(n6927) );
  OAI222_X1 U8247 ( .A1(n8947), .A2(n6684), .B1(n8946), .B2(n6686), .C1(
        P2_U3152), .C2(n6927), .ZN(P2_U3352) );
  INV_X1 U8248 ( .A(n6754), .ZN(n6790) );
  INV_X1 U8249 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6685) );
  OAI222_X1 U8250 ( .A1(n6790), .A2(n10130), .B1(n9443), .B2(n6686), .C1(n6685), .C2(n8318), .ZN(P1_U3347) );
  INV_X1 U8251 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6688) );
  INV_X1 U8252 ( .A(n6687), .ZN(n6689) );
  INV_X1 U8253 ( .A(n6746), .ZN(n6780) );
  OAI222_X1 U8254 ( .A1(n8318), .A2(n6688), .B1(n9443), .B2(n6689), .C1(n6780), 
        .C2(n10130), .ZN(P1_U3346) );
  INV_X1 U8255 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6690) );
  INV_X1 U8256 ( .A(n6954), .ZN(n6961) );
  OAI222_X1 U8257 ( .A1(n8947), .A2(n6690), .B1(n8946), .B2(n6689), .C1(
        P2_U3152), .C2(n6961), .ZN(P2_U3351) );
  INV_X1 U8258 ( .A(n6968), .ZN(n6977) );
  INV_X1 U8259 ( .A(n6691), .ZN(n6693) );
  OAI222_X1 U8260 ( .A1(n6977), .A2(P1_U3084), .B1(n9443), .B2(n6693), .C1(
        n6692), .C2(n8318), .ZN(P1_U3345) );
  INV_X1 U8261 ( .A(n7122), .ZN(n7128) );
  OAI222_X1 U8262 ( .A1(n8947), .A2(n6694), .B1(n8946), .B2(n6693), .C1(
        P2_U3152), .C2(n7128), .ZN(P2_U3350) );
  INV_X1 U8263 ( .A(P1_U4006), .ZN(n9084) );
  NAND2_X1 U8264 ( .A1(n9084), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n6695) );
  OAI21_X1 U8265 ( .B1(n9149), .B2(n9084), .A(n6695), .ZN(P1_U3586) );
  INV_X1 U8266 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6700) );
  NAND2_X1 U8267 ( .A1(n5045), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6698) );
  NAND2_X1 U8268 ( .A1(n5025), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6697) );
  NAND2_X1 U8269 ( .A1(n8076), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6696) );
  NAND3_X1 U8270 ( .A1(n6698), .A2(n6697), .A3(n6696), .ZN(n8605) );
  NAND2_X1 U8271 ( .A1(n8605), .A2(P2_U3966), .ZN(n6699) );
  OAI21_X1 U8272 ( .B1(n6700), .B2(P2_U3966), .A(n6699), .ZN(P2_U3583) );
  INV_X1 U8273 ( .A(n6701), .ZN(n6704) );
  OAI222_X1 U8274 ( .A1(n10130), .A2(n6703), .B1(n9443), .B2(n6704), .C1(n6702), .C2(n8318), .ZN(P1_U3344) );
  INV_X1 U8275 ( .A(n7293), .ZN(n7135) );
  OAI222_X1 U8276 ( .A1(n8947), .A2(n6705), .B1(n8946), .B2(n6704), .C1(n7135), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U8277 ( .A(n6706), .ZN(n6772) );
  AOI22_X1 U8278 ( .A1(n7799), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n8943), .ZN(n6707) );
  OAI21_X1 U8279 ( .B1(n6772), .B2(n8946), .A(n6707), .ZN(P2_U3347) );
  INV_X1 U8280 ( .A(n5824), .ZN(n6710) );
  INV_X1 U8281 ( .A(n7649), .ZN(n7302) );
  OAI222_X1 U8282 ( .A1(n8947), .A2(n6708), .B1(n8946), .B2(n6710), .C1(n7302), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U8283 ( .A(n9879), .ZN(n6966) );
  OAI222_X1 U8284 ( .A1(P1_U3084), .A2(n6966), .B1(n9443), .B2(n6710), .C1(
        n6709), .C2(n8318), .ZN(P1_U3343) );
  INV_X1 U8285 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6733) );
  NOR2_X1 U8286 ( .A1(n6323), .A2(P1_U3084), .ZN(n9440) );
  NAND2_X1 U8287 ( .A1(n6719), .A2(n9440), .ZN(n9142) );
  INV_X1 U8288 ( .A(n9142), .ZN(n6728) );
  AND2_X1 U8289 ( .A1(n10130), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6824) );
  XNOR2_X1 U8290 ( .A(n9811), .B(n6711), .ZN(n9812) );
  INV_X1 U8291 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6724) );
  NAND2_X1 U8292 ( .A1(n6713), .A2(n6712), .ZN(n9813) );
  NAND2_X1 U8293 ( .A1(n9811), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6714) );
  INV_X1 U8294 ( .A(n6717), .ZN(n6721) );
  INV_X1 U8295 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6715) );
  XNOR2_X1 U8296 ( .A(n6748), .B(n6715), .ZN(n6716) );
  INV_X1 U8297 ( .A(n6716), .ZN(n6720) );
  NOR2_X1 U8298 ( .A1(n6241), .A2(n10130), .ZN(n9776) );
  AND2_X1 U8299 ( .A1(n9776), .A2(n6323), .ZN(n6718) );
  INV_X1 U8300 ( .A(n9894), .ZN(n9843) );
  AOI211_X1 U8301 ( .C1(n6721), .C2(n6720), .A(n6738), .B(n9843), .ZN(n6722)
         );
  AOI211_X1 U8302 ( .C1(n9886), .C2(n6748), .A(n6824), .B(n6722), .ZN(n6732)
         );
  MUX2_X1 U8303 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6723), .S(n6748), .Z(n6730)
         );
  XNOR2_X1 U8304 ( .A(n9811), .B(n5676), .ZN(n9809) );
  NOR2_X1 U8305 ( .A1(n6724), .A2(n5635), .ZN(n9796) );
  XNOR2_X1 U8306 ( .A(n9793), .B(n5654), .ZN(n9795) );
  NAND2_X1 U8307 ( .A1(n9796), .A2(n9795), .ZN(n9794) );
  NAND2_X1 U8308 ( .A1(n9811), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6725) );
  NAND2_X1 U8309 ( .A1(n6726), .A2(n6725), .ZN(n6729) );
  NAND2_X1 U8310 ( .A1(n6729), .A2(n6730), .ZN(n6750) );
  OAI211_X1 U8311 ( .C1(n6730), .C2(n6729), .A(n9895), .B(n6750), .ZN(n6731)
         );
  OAI211_X1 U8312 ( .C1(n6733), .C2(n9899), .A(n6732), .B(n6731), .ZN(P1_U3244) );
  INV_X1 U8313 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6764) );
  NOR2_X1 U8314 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6734), .ZN(n7312) );
  MUX2_X1 U8315 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n6735), .S(n6746), .Z(n6779)
         );
  NAND2_X1 U8316 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n9849), .ZN(n6736) );
  OAI21_X1 U8317 ( .B1(n9849), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6736), .ZN(
        n9845) );
  AND2_X1 U8318 ( .A1(n6748), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6737) );
  MUX2_X1 U8319 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6739), .S(n9830), .Z(n6740)
         );
  NAND2_X1 U8320 ( .A1(n9829), .A2(n6740), .ZN(n9834) );
  OAI21_X1 U8321 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n9830), .A(n9834), .ZN(
        n9846) );
  NOR2_X1 U8322 ( .A1(n9845), .A2(n9846), .ZN(n9844) );
  AOI21_X1 U8323 ( .B1(n9849), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9844), .ZN(
        n6787) );
  NOR2_X1 U8324 ( .A1(n6754), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6741) );
  AOI21_X1 U8325 ( .B1(n6754), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6741), .ZN(
        n6788) );
  NAND2_X1 U8326 ( .A1(n6787), .A2(n6788), .ZN(n6786) );
  MUX2_X1 U8327 ( .A(n6742), .B(P1_REG1_REG_8__SCAN_IN), .S(n6968), .Z(n6743)
         );
  AOI211_X1 U8328 ( .C1(n6744), .C2(n6743), .A(n6967), .B(n9843), .ZN(n6745)
         );
  AOI211_X1 U8329 ( .C1(n9886), .C2(n6968), .A(n7312), .B(n6745), .ZN(n6763)
         );
  INV_X1 U8330 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6747) );
  OR2_X1 U8331 ( .A1(n6746), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6757) );
  MUX2_X1 U8332 ( .A(n6747), .B(P1_REG2_REG_7__SCAN_IN), .S(n6746), .Z(n6775)
         );
  NOR2_X1 U8333 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n9849), .ZN(n6753) );
  NAND2_X1 U8334 ( .A1(n6748), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6749) );
  NAND2_X1 U8335 ( .A1(n6750), .A2(n6749), .ZN(n9826) );
  AOI22_X1 U8336 ( .A1(n9830), .A2(n5702), .B1(P1_REG2_REG_4__SCAN_IN), .B2(
        n6751), .ZN(n9825) );
  NOR2_X1 U8337 ( .A1(n9826), .A2(n9825), .ZN(n9828) );
  AOI21_X1 U8338 ( .B1(n6751), .B2(n5702), .A(n9828), .ZN(n9851) );
  MUX2_X1 U8339 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n7213), .S(n9849), .Z(n6752)
         );
  INV_X1 U8340 ( .A(n6752), .ZN(n9852) );
  MUX2_X1 U8341 ( .A(n5734), .B(P1_REG2_REG_6__SCAN_IN), .S(n6754), .Z(n6755)
         );
  INV_X1 U8342 ( .A(n6755), .ZN(n6794) );
  NOR2_X1 U8343 ( .A1(n6775), .A2(n6776), .ZN(n6774) );
  INV_X1 U8344 ( .A(n6774), .ZN(n6756) );
  AND2_X1 U8345 ( .A1(n6757), .A2(n6756), .ZN(n6980) );
  MUX2_X1 U8346 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n6758), .S(n6968), .Z(n6761)
         );
  NOR2_X1 U8347 ( .A1(n6977), .A2(n6758), .ZN(n6978) );
  INV_X1 U8348 ( .A(n6978), .ZN(n6759) );
  OAI211_X1 U8349 ( .C1(n6968), .C2(P1_REG2_REG_8__SCAN_IN), .A(n6759), .B(
        n6980), .ZN(n6760) );
  OAI211_X1 U8350 ( .C1(n6980), .C2(n6761), .A(n9895), .B(n6760), .ZN(n6762)
         );
  OAI211_X1 U8351 ( .C1(n6764), .C2(n9899), .A(n6763), .B(n6762), .ZN(P1_U3249) );
  OR2_X1 U8352 ( .A1(n6765), .A2(P2_U3152), .ZN(n8296) );
  NAND2_X1 U8353 ( .A1(n10027), .A2(n8296), .ZN(n6767) );
  NAND2_X1 U8354 ( .A1(n6767), .A2(n6766), .ZN(n6770) );
  OR2_X1 U8355 ( .A1(n10027), .A2(n6768), .ZN(n6769) );
  AND2_X1 U8356 ( .A1(n6770), .A2(n6769), .ZN(n8602) );
  NOR2_X1 U8357 ( .A1(n9994), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8358 ( .A(n6983), .ZN(n9089) );
  OAI222_X1 U8359 ( .A1(n10130), .A2(n9089), .B1(n9443), .B2(n6772), .C1(n6771), .C2(n8318), .ZN(P1_U3342) );
  INV_X1 U8360 ( .A(n5859), .ZN(n6800) );
  AOI22_X1 U8361 ( .A1(n8527), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n8943), .ZN(n6773) );
  OAI21_X1 U8362 ( .B1(n6800), .B2(n8946), .A(n6773), .ZN(P2_U3346) );
  AOI21_X1 U8363 ( .B1(n6776), .B2(n6775), .A(n6774), .ZN(n6785) );
  OAI21_X1 U8364 ( .B1(n6779), .B2(n6778), .A(n6777), .ZN(n6782) );
  AND2_X1 U8365 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7189) );
  NOR2_X1 U8366 ( .A1(n9114), .A2(n6780), .ZN(n6781) );
  AOI211_X1 U8367 ( .C1(n9894), .C2(n6782), .A(n7189), .B(n6781), .ZN(n6784)
         );
  NAND2_X1 U8368 ( .A1(n9880), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n6783) );
  OAI211_X1 U8369 ( .C1(n6785), .C2(n9872), .A(n6784), .B(n6783), .ZN(P1_U3248) );
  INV_X1 U8370 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6798) );
  OAI21_X1 U8371 ( .B1(n6788), .B2(n6787), .A(n6786), .ZN(n6792) );
  NOR2_X1 U8372 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6789), .ZN(n7264) );
  NOR2_X1 U8373 ( .A1(n9114), .A2(n6790), .ZN(n6791) );
  AOI211_X1 U8374 ( .C1(n9894), .C2(n6792), .A(n7264), .B(n6791), .ZN(n6797)
         );
  OAI211_X1 U8375 ( .C1(n6795), .C2(n6794), .A(n9895), .B(n6793), .ZN(n6796)
         );
  OAI211_X1 U8376 ( .C1(n6798), .C2(n9899), .A(n6797), .B(n6796), .ZN(P1_U3247) );
  INV_X1 U8377 ( .A(n7111), .ZN(n6975) );
  OAI222_X1 U8378 ( .A1(n6975), .A2(n10130), .B1(n9443), .B2(n6800), .C1(n6799), .C2(n8318), .ZN(P1_U3341) );
  INV_X1 U8379 ( .A(n5883), .ZN(n6810) );
  AOI22_X1 U8380 ( .A1(n7485), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9441), .ZN(n6801) );
  OAI21_X1 U8381 ( .B1(n6810), .B2(n9443), .A(n6801), .ZN(P1_U3340) );
  INV_X1 U8382 ( .A(n7157), .ZN(n6802) );
  NAND2_X1 U8383 ( .A1(n6802), .A2(n7168), .ZN(n6803) );
  OR2_X1 U8384 ( .A1(n6804), .A2(n6803), .ZN(n6806) );
  NAND2_X1 U8385 ( .A1(n6259), .A2(n9709), .ZN(n6805) );
  NAND2_X1 U8386 ( .A1(n6806), .A2(n6805), .ZN(n7236) );
  AOI21_X1 U8387 ( .B1(n7235), .B2(n7157), .A(n7236), .ZN(n6809) );
  NAND2_X1 U8388 ( .A1(n6336), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6807) );
  OAI21_X1 U8389 ( .B1(n6809), .B2(n6336), .A(n6807), .ZN(P1_U3523) );
  NAND2_X1 U8390 ( .A1(n6341), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6808) );
  OAI21_X1 U8391 ( .B1(n6809), .B2(n6341), .A(n6808), .ZN(P1_U3454) );
  INV_X1 U8392 ( .A(n7874), .ZN(n7869) );
  OAI222_X1 U8393 ( .A1(n8947), .A2(n6811), .B1(n8946), .B2(n6810), .C1(n7869), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  OAI21_X1 U8394 ( .B1(n6814), .B2(n6813), .A(n6812), .ZN(n9800) );
  AOI22_X1 U8395 ( .A1(n9800), .A2(n6223), .B1(n9052), .B2(n7235), .ZN(n6817)
         );
  NAND2_X1 U8396 ( .A1(n7318), .A2(n6815), .ZN(n6894) );
  AOI22_X1 U8397 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n6894), .B1(n9024), .B2(
        n6259), .ZN(n6816) );
  NAND2_X1 U8398 ( .A1(n6817), .A2(n6816), .ZN(P1_U3230) );
  INV_X1 U8399 ( .A(n6818), .ZN(n6820) );
  INV_X1 U8400 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6819) );
  OAI222_X1 U8401 ( .A1(P1_U3084), .A2(n7736), .B1(n9443), .B2(n6820), .C1(
        n6819), .C2(n8318), .ZN(P1_U3339) );
  INV_X1 U8402 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6821) );
  OAI222_X1 U8403 ( .A1(n8947), .A2(n6821), .B1(n8946), .B2(n6820), .C1(n7879), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  XOR2_X1 U8404 ( .A(n6823), .B(n6822), .Z(n6829) );
  AOI21_X1 U8405 ( .B1(n9024), .B2(n9082), .A(n6824), .ZN(n6825) );
  OAI21_X1 U8406 ( .B1(n7404), .B2(n9060), .A(n6825), .ZN(n6827) );
  NOR2_X1 U8407 ( .A1(n9050), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6826) );
  AOI211_X1 U8408 ( .C1(n9052), .C2(n7400), .A(n6827), .B(n6826), .ZN(n6828)
         );
  OAI21_X1 U8409 ( .B1(n6829), .B2(n9054), .A(n6828), .ZN(P1_U3216) );
  NAND2_X1 U8410 ( .A1(n6830), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8945) );
  OR2_X1 U8411 ( .A1(n10027), .A2(n6831), .ZN(n6832) );
  OAI211_X1 U8412 ( .C1(n6833), .C2(n8945), .A(n6832), .B(n8296), .ZN(n6836)
         );
  NAND2_X1 U8413 ( .A1(n6836), .A2(n5006), .ZN(n6834) );
  NAND2_X1 U8414 ( .A1(n6834), .A2(n8521), .ZN(n6842) );
  INV_X1 U8415 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10085) );
  INV_X1 U8416 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9567) );
  OAI22_X1 U8417 ( .A1(n8602), .A2(n10085), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9567), .ZN(n6840) );
  NAND2_X1 U8418 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n6838) );
  NOR2_X1 U8419 ( .A1(n6837), .A2(n6838), .ZN(n6847) );
  AND2_X1 U8420 ( .A1(n5006), .A2(n8949), .ZN(n6835) );
  AOI211_X1 U8421 ( .C1(n6838), .C2(n6837), .A(n6847), .B(n9996), .ZN(n6839)
         );
  AOI211_X1 U8422 ( .C1(n8596), .C2(n6848), .A(n6840), .B(n6839), .ZN(n6846)
         );
  AND2_X1 U8423 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(
        n6844) );
  INV_X1 U8424 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6856) );
  MUX2_X1 U8425 ( .A(n6856), .B(P2_REG2_REG_1__SCAN_IN), .S(n6855), .Z(n6843)
         );
  NOR2_X1 U8426 ( .A1(n5534), .A2(n8949), .ZN(n6841) );
  NAND3_X1 U8427 ( .A1(n6843), .A2(P2_REG2_REG_0__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n6854) );
  OAI211_X1 U8428 ( .C1(n6844), .C2(n6843), .A(n9992), .B(n6854), .ZN(n6845)
         );
  NAND2_X1 U8429 ( .A1(n6846), .A2(n6845), .ZN(P2_U3246) );
  NAND2_X1 U8430 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n7705) );
  INV_X1 U8431 ( .A(n7705), .ZN(n6853) );
  AOI21_X1 U8432 ( .B1(P2_REG1_REG_1__SCAN_IN), .B2(n6848), .A(n6847), .ZN(
        n6945) );
  XNOR2_X1 U8433 ( .A(n6857), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n6944) );
  NOR2_X1 U8434 ( .A1(n6945), .A2(n6944), .ZN(n6943) );
  XNOR2_X1 U8435 ( .A(n6858), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n6869) );
  INV_X1 U8436 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6849) );
  MUX2_X1 U8437 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6849), .S(n6905), .Z(n6850)
         );
  AOI211_X1 U8438 ( .C1(n6851), .C2(n6850), .A(n6897), .B(n9996), .ZN(n6852)
         );
  AOI211_X1 U8439 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n9994), .A(n6853), .B(
        n6852), .ZN(n6867) );
  INV_X1 U8440 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n8831) );
  MUX2_X1 U8441 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n8831), .S(n6857), .Z(n6950)
         );
  OAI21_X1 U8442 ( .B1(n6856), .B2(n6855), .A(n6854), .ZN(n6949) );
  NAND2_X1 U8443 ( .A1(n6950), .A2(n6949), .ZN(n6948) );
  NAND2_X1 U8444 ( .A1(n6857), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6874) );
  INV_X1 U8445 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7472) );
  MUX2_X1 U8446 ( .A(n7472), .B(P2_REG2_REG_3__SCAN_IN), .S(n6858), .Z(n6873)
         );
  AOI21_X1 U8447 ( .B1(n6948), .B2(n6874), .A(n6873), .ZN(n6861) );
  NOR2_X1 U8448 ( .A1(n6879), .A2(n7472), .ZN(n6862) );
  INV_X1 U8449 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6859) );
  MUX2_X1 U8450 ( .A(n6859), .B(P2_REG2_REG_4__SCAN_IN), .S(n6905), .Z(n6860)
         );
  OAI21_X1 U8451 ( .B1(n6861), .B2(n6862), .A(n6860), .ZN(n6904) );
  INV_X1 U8452 ( .A(n6861), .ZN(n6876) );
  INV_X1 U8453 ( .A(n6862), .ZN(n6864) );
  MUX2_X1 U8454 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6859), .S(n6905), .Z(n6863)
         );
  NAND3_X1 U8455 ( .A1(n6876), .A2(n6864), .A3(n6863), .ZN(n6865) );
  NAND3_X1 U8456 ( .A1(n9992), .A2(n6904), .A3(n6865), .ZN(n6866) );
  OAI211_X1 U8457 ( .C1(n9995), .C2(n6905), .A(n6867), .B(n6866), .ZN(P2_U3249) );
  NOR2_X1 U8458 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5047), .ZN(n6872) );
  AOI211_X1 U8459 ( .C1(n6870), .C2(n6869), .A(n6868), .B(n9996), .ZN(n6871)
         );
  AOI211_X1 U8460 ( .C1(P2_ADDR_REG_3__SCAN_IN), .C2(n9994), .A(n6872), .B(
        n6871), .ZN(n6878) );
  NAND3_X1 U8461 ( .A1(n6948), .A2(n6874), .A3(n6873), .ZN(n6875) );
  NAND3_X1 U8462 ( .A1(n9992), .A2(n6876), .A3(n6875), .ZN(n6877) );
  OAI211_X1 U8463 ( .C1(n9995), .C2(n6879), .A(n6878), .B(n6877), .ZN(P2_U3248) );
  NAND2_X1 U8464 ( .A1(n6881), .A2(n6880), .ZN(n6883) );
  XOR2_X1 U8465 ( .A(n6883), .B(n6882), .Z(n6888) );
  INV_X1 U8466 ( .A(n6258), .ZN(n6884) );
  OAI22_X1 U8467 ( .A1(n6884), .A2(n9060), .B1(n9062), .B2(n7404), .ZN(n6886)
         );
  INV_X1 U8468 ( .A(n9052), .ZN(n9069) );
  NOR2_X1 U8469 ( .A1(n9069), .A2(n9936), .ZN(n6885) );
  AOI211_X1 U8470 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n6894), .A(n6886), .B(
        n6885), .ZN(n6887) );
  OAI21_X1 U8471 ( .B1(n6888), .B2(n9054), .A(n6887), .ZN(P1_U3220) );
  XOR2_X1 U8472 ( .A(n6890), .B(n6889), .Z(n6896) );
  OAI22_X1 U8473 ( .A1(n7005), .A2(n9060), .B1(n9062), .B2(n7143), .ZN(n6893)
         );
  NOR2_X1 U8474 ( .A1(n9069), .A2(n6891), .ZN(n6892) );
  AOI211_X1 U8475 ( .C1(P1_REG3_REG_2__SCAN_IN), .C2(n6894), .A(n6893), .B(
        n6892), .ZN(n6895) );
  OAI21_X1 U8476 ( .B1(n6896), .B2(n9054), .A(n6895), .ZN(P1_U3235) );
  AND2_X1 U8477 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6903) );
  INV_X1 U8478 ( .A(n6905), .ZN(n6898) );
  AOI21_X1 U8479 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(n6898), .A(n6897), .ZN(
        n6901) );
  NAND2_X1 U8480 ( .A1(n6919), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6899) );
  OAI21_X1 U8481 ( .B1(n6919), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6899), .ZN(
        n6900) );
  NOR2_X1 U8482 ( .A1(n6901), .A2(n6900), .ZN(n6913) );
  AOI211_X1 U8483 ( .C1(n6901), .C2(n6900), .A(n6913), .B(n9996), .ZN(n6902)
         );
  AOI211_X1 U8484 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n9994), .A(n6903), .B(
        n6902), .ZN(n6911) );
  OAI21_X1 U8485 ( .B1(n6859), .B2(n6905), .A(n6904), .ZN(n6909) );
  INV_X1 U8486 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6906) );
  MUX2_X1 U8487 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n6906), .S(n6912), .Z(n6907)
         );
  INV_X1 U8488 ( .A(n6907), .ZN(n6908) );
  NAND2_X1 U8489 ( .A1(n6908), .A2(n6909), .ZN(n6920) );
  OAI211_X1 U8490 ( .C1(n6909), .C2(n6908), .A(n9992), .B(n6920), .ZN(n6910)
         );
  OAI211_X1 U8491 ( .C1(n9995), .C2(n6912), .A(n6911), .B(n6910), .ZN(P2_U3250) );
  NOR2_X1 U8492 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9558), .ZN(n6918) );
  AOI21_X1 U8493 ( .B1(n6919), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6913), .ZN(
        n6916) );
  NAND2_X1 U8494 ( .A1(n6934), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6914) );
  OAI21_X1 U8495 ( .B1(n6934), .B2(P2_REG1_REG_6__SCAN_IN), .A(n6914), .ZN(
        n6915) );
  NOR2_X1 U8496 ( .A1(n6916), .A2(n6915), .ZN(n6928) );
  AOI211_X1 U8497 ( .C1(n6916), .C2(n6915), .A(n6928), .B(n9996), .ZN(n6917)
         );
  AOI211_X1 U8498 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n9994), .A(n6918), .B(
        n6917), .ZN(n6926) );
  NAND2_X1 U8499 ( .A1(n6919), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6921) );
  NAND2_X1 U8500 ( .A1(n6921), .A2(n6920), .ZN(n6924) );
  INV_X1 U8501 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6922) );
  MUX2_X1 U8502 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6922), .S(n6934), .Z(n6923)
         );
  NAND2_X1 U8503 ( .A1(n6923), .A2(n6924), .ZN(n6935) );
  OAI211_X1 U8504 ( .C1(n6924), .C2(n6923), .A(n9992), .B(n6935), .ZN(n6925)
         );
  OAI211_X1 U8505 ( .C1(n9995), .C2(n6927), .A(n6926), .B(n6925), .ZN(P2_U3251) );
  NOR2_X1 U8506 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5117), .ZN(n6933) );
  INV_X1 U8507 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6929) );
  MUX2_X1 U8508 ( .A(n6929), .B(P2_REG1_REG_7__SCAN_IN), .S(n6954), .Z(n6930)
         );
  AOI211_X1 U8509 ( .C1(n6931), .C2(n6930), .A(n6953), .B(n9996), .ZN(n6932)
         );
  AOI211_X1 U8510 ( .C1(P2_ADDR_REG_7__SCAN_IN), .C2(n9994), .A(n6933), .B(
        n6932), .ZN(n6941) );
  NAND2_X1 U8511 ( .A1(n6934), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6936) );
  NAND2_X1 U8512 ( .A1(n6936), .A2(n6935), .ZN(n6939) );
  INV_X1 U8513 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6937) );
  MUX2_X1 U8514 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n6937), .S(n6954), .Z(n6938)
         );
  NAND2_X1 U8515 ( .A1(n6938), .A2(n6939), .ZN(n6960) );
  OAI211_X1 U8516 ( .C1(n6939), .C2(n6938), .A(n9992), .B(n6960), .ZN(n6940)
         );
  OAI211_X1 U8517 ( .C1(n9995), .C2(n6961), .A(n6941), .B(n6940), .ZN(P2_U3252) );
  INV_X1 U8518 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6942) );
  NOR2_X1 U8519 ( .A1(n6942), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6947) );
  AOI211_X1 U8520 ( .C1(n6945), .C2(n6944), .A(n6943), .B(n9996), .ZN(n6946)
         );
  AOI211_X1 U8521 ( .C1(P2_ADDR_REG_2__SCAN_IN), .C2(n9994), .A(n6947), .B(
        n6946), .ZN(n6952) );
  OAI211_X1 U8522 ( .C1(n6950), .C2(n6949), .A(n9992), .B(n6948), .ZN(n6951)
         );
  OAI211_X1 U8523 ( .C1(n9995), .C2(n4547), .A(n6952), .B(n6951), .ZN(P2_U3247) );
  NOR2_X1 U8524 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9573), .ZN(n6959) );
  INV_X1 U8525 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6955) );
  MUX2_X1 U8526 ( .A(n6955), .B(P2_REG1_REG_8__SCAN_IN), .S(n7122), .Z(n6956)
         );
  AOI211_X1 U8527 ( .C1(n6957), .C2(n6956), .A(n7121), .B(n9996), .ZN(n6958)
         );
  AOI211_X1 U8528 ( .C1(P2_ADDR_REG_8__SCAN_IN), .C2(n9994), .A(n6959), .B(
        n6958), .ZN(n6965) );
  OAI21_X1 U8529 ( .B1(n6961), .B2(n6937), .A(n6960), .ZN(n6963) );
  INV_X1 U8530 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7338) );
  MUX2_X1 U8531 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n7338), .S(n7122), .Z(n6962)
         );
  NAND2_X1 U8532 ( .A1(n6962), .A2(n6963), .ZN(n7127) );
  OAI211_X1 U8533 ( .C1(n6963), .C2(n6962), .A(n9992), .B(n7127), .ZN(n6964)
         );
  OAI211_X1 U8534 ( .C1(n9995), .C2(n7128), .A(n6965), .B(n6964), .ZN(P2_U3253) );
  INV_X1 U8535 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9765) );
  AOI22_X1 U8536 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n6983), .B1(n9089), .B2(
        n9765), .ZN(n9087) );
  AOI22_X1 U8537 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n9879), .B1(n6966), .B2(
        n5829), .ZN(n9871) );
  AOI21_X1 U8538 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n6968), .A(n6967), .ZN(
        n9859) );
  NOR2_X1 U8539 ( .A1(n9866), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6969) );
  AOI21_X1 U8540 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9866), .A(n6969), .ZN(
        n9858) );
  NAND2_X1 U8541 ( .A1(n9859), .A2(n9858), .ZN(n9857) );
  OAI21_X1 U8542 ( .B1(n9866), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9857), .ZN(
        n9870) );
  NAND2_X1 U8543 ( .A1(n9871), .A2(n9870), .ZN(n9869) );
  OR2_X1 U8544 ( .A1(n7111), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6971) );
  NAND2_X1 U8545 ( .A1(n7111), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6970) );
  AND2_X1 U8546 ( .A1(n6971), .A2(n6970), .ZN(n6972) );
  OAI21_X1 U8547 ( .B1(n6973), .B2(n6972), .A(n7104), .ZN(n6989) );
  NAND2_X1 U8548 ( .A1(n9880), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6974) );
  NAND2_X1 U8549 ( .A1(n10130), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7825) );
  OAI211_X1 U8550 ( .C1(n9114), .C2(n6975), .A(n6974), .B(n7825), .ZN(n6988)
         );
  NOR2_X1 U8551 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n6983), .ZN(n6976) );
  AOI21_X1 U8552 ( .B1(n6983), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6976), .ZN(
        n9094) );
  NAND2_X1 U8553 ( .A1(n6977), .A2(n6758), .ZN(n6979) );
  AOI21_X1 U8554 ( .B1(n6980), .B2(n6979), .A(n6978), .ZN(n9862) );
  NAND2_X1 U8555 ( .A1(n9866), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6981) );
  OAI21_X1 U8556 ( .B1(n9866), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6981), .ZN(
        n9861) );
  NAND2_X1 U8557 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n9879), .ZN(n6982) );
  OAI21_X1 U8558 ( .B1(n9879), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6982), .ZN(
        n9874) );
  NAND2_X1 U8559 ( .A1(n9094), .A2(n9093), .ZN(n9092) );
  OAI21_X1 U8560 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n6983), .A(n9092), .ZN(
        n6986) );
  NAND2_X1 U8561 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7111), .ZN(n6984) );
  OAI21_X1 U8562 ( .B1(n7111), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6984), .ZN(
        n6985) );
  NOR2_X1 U8563 ( .A1(n6985), .A2(n6986), .ZN(n7110) );
  AOI211_X1 U8564 ( .C1(n6986), .C2(n6985), .A(n7110), .B(n9872), .ZN(n6987)
         );
  AOI211_X1 U8565 ( .C1(n9894), .C2(n6989), .A(n6988), .B(n6987), .ZN(n6990)
         );
  INV_X1 U8566 ( .A(n6990), .ZN(P1_U3253) );
  AOI21_X1 U8567 ( .B1(n6991), .B2(n6992), .A(n9054), .ZN(n6994) );
  NAND2_X1 U8568 ( .A1(n6994), .A2(n6993), .ZN(n6998) );
  AND2_X1 U8569 ( .A1(n10130), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9835) );
  AOI21_X1 U8570 ( .B1(n9048), .B2(n9083), .A(n9835), .ZN(n6995) );
  OAI21_X1 U8571 ( .B1(n7142), .B2(n9062), .A(n6995), .ZN(n6996) );
  AOI21_X1 U8572 ( .B1(n9052), .B2(n7195), .A(n6996), .ZN(n6997) );
  OAI211_X1 U8573 ( .C1(n9050), .C2(n7159), .A(n6998), .B(n6997), .ZN(P1_U3228) );
  INV_X1 U8574 ( .A(n6999), .ZN(n7002) );
  INV_X1 U8575 ( .A(n8547), .ZN(n8537) );
  OAI222_X1 U8576 ( .A1(n8947), .A2(n7000), .B1(n8946), .B2(n7002), .C1(
        P2_U3152), .C2(n8537), .ZN(P2_U3343) );
  OAI222_X1 U8577 ( .A1(n9106), .A2(P1_U3084), .B1(n9443), .B2(n7002), .C1(
        n7001), .C2(n8318), .ZN(P1_U3338) );
  OAI21_X1 U8578 ( .B1(n7004), .B2(n7006), .A(n7003), .ZN(n9330) );
  INV_X1 U8579 ( .A(n9330), .ZN(n7015) );
  INV_X1 U8580 ( .A(n9710), .ZN(n9916) );
  OAI22_X1 U8581 ( .A1(n7005), .A2(n9916), .B1(n7143), .B2(n9914), .ZN(n7010)
         );
  XNOR2_X1 U8582 ( .A(n7007), .B(n7006), .ZN(n7008) );
  NOR2_X1 U8583 ( .A1(n7008), .A2(n9732), .ZN(n7009) );
  AOI211_X1 U8584 ( .C1(n9735), .C2(n9330), .A(n7010), .B(n7009), .ZN(n9326)
         );
  NAND2_X1 U8585 ( .A1(n9936), .A2(n7011), .ZN(n7012) );
  NAND2_X1 U8586 ( .A1(n9329), .A2(n7012), .ZN(n7013) );
  AND2_X1 U8587 ( .A1(n7013), .A2(n7395), .ZN(n9331) );
  AOI22_X1 U8588 ( .A1(n9331), .A2(n9395), .B1(n9745), .B2(n9329), .ZN(n7014)
         );
  OAI211_X1 U8589 ( .C1(n7015), .C2(n9659), .A(n9326), .B(n7014), .ZN(n7017)
         );
  NAND2_X1 U8590 ( .A1(n7017), .A2(n9990), .ZN(n7016) );
  OAI21_X1 U8591 ( .B1(n9990), .B2(n6711), .A(n7016), .ZN(P1_U3525) );
  INV_X1 U8592 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7019) );
  NAND2_X1 U8593 ( .A1(n7017), .A2(n9980), .ZN(n7018) );
  OAI21_X1 U8594 ( .B1(n9980), .B2(n7019), .A(n7018), .ZN(P1_U3460) );
  INV_X1 U8595 ( .A(n10027), .ZN(n7020) );
  AND2_X1 U8596 ( .A1(n7073), .A2(n7070), .ZN(n7022) );
  INV_X1 U8597 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7033) );
  XNOR2_X1 U8598 ( .A(n7339), .B(n7024), .ZN(n8812) );
  NAND3_X1 U8599 ( .A1(n8252), .A2(n8657), .A3(n7024), .ZN(n9685) );
  NAND2_X1 U8600 ( .A1(n7556), .A2(n10003), .ZN(n7047) );
  INV_X1 U8601 ( .A(n10003), .ZN(n7026) );
  NAND2_X1 U8602 ( .A1(n7047), .A2(n8120), .ZN(n7027) );
  INV_X1 U8603 ( .A(n7040), .ZN(n7028) );
  NAND2_X1 U8604 ( .A1(n7027), .A2(n7028), .ZN(n7039) );
  OAI21_X1 U8605 ( .B1(n7027), .B2(n7028), .A(n7039), .ZN(n10005) );
  INV_X1 U8606 ( .A(n10005), .ZN(n7031) );
  NAND2_X1 U8607 ( .A1(n5519), .A2(n8286), .ZN(n8089) );
  XNOR2_X1 U8608 ( .A(n7027), .B(n7048), .ZN(n7029) );
  OAI22_X1 U8609 ( .A1(n7550), .A2(n8808), .B1(n8806), .B2(n7242), .ZN(n7517)
         );
  AOI21_X1 U8610 ( .B1(n8793), .B2(n7029), .A(n7517), .ZN(n10007) );
  AOI211_X1 U8611 ( .C1(n7553), .C2(n10003), .A(n7063), .B(n10064), .ZN(n10010) );
  AOI21_X1 U8612 ( .B1(n9677), .B2(n10003), .A(n10010), .ZN(n7030) );
  OAI211_X1 U8613 ( .C1(n8914), .C2(n7031), .A(n10007), .B(n7030), .ZN(n7076)
         );
  NAND2_X1 U8614 ( .A1(n4316), .A2(n7076), .ZN(n7032) );
  OAI21_X1 U8615 ( .B1(n4316), .B2(n7033), .A(n7032), .ZN(P2_U3454) );
  INV_X1 U8616 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7036) );
  INV_X1 U8617 ( .A(n7553), .ZN(n10017) );
  NAND2_X1 U8618 ( .A1(n8522), .A2(n10017), .ZN(n8119) );
  NAND2_X1 U8619 ( .A1(n7048), .A2(n8119), .ZN(n10013) );
  NAND2_X1 U8620 ( .A1(n10068), .A2(n10013), .ZN(n7034) );
  AOI22_X1 U8621 ( .A1(n10013), .A2(n8793), .B1(n8790), .B2(n7025), .ZN(n10016) );
  OAI211_X1 U8622 ( .C1(n10017), .C2(n5510), .A(n7034), .B(n10016), .ZN(n7084)
         );
  NAND2_X1 U8623 ( .A1(n4316), .A2(n7084), .ZN(n7035) );
  OAI21_X1 U8624 ( .B1(n4316), .B2(n7036), .A(n7035), .ZN(P2_U3451) );
  INV_X1 U8625 ( .A(n7037), .ZN(n7101) );
  AOI22_X1 U8626 ( .A1(n8553), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n8943), .ZN(n7038) );
  OAI21_X1 U8627 ( .B1(n7101), .B2(n8946), .A(n7038), .ZN(P2_U3342) );
  INV_X1 U8628 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n7058) );
  NAND2_X1 U8629 ( .A1(n7040), .A2(n7025), .ZN(n7041) );
  NAND2_X1 U8630 ( .A1(n8520), .A2(n7052), .ZN(n8123) );
  NAND2_X1 U8631 ( .A1(n7242), .A2(n7052), .ZN(n7042) );
  NAND2_X1 U8632 ( .A1(n7043), .A2(n7042), .ZN(n7458) );
  NAND2_X1 U8633 ( .A1(n8519), .A2(n4425), .ZN(n8128) );
  NAND2_X1 U8634 ( .A1(n7092), .A2(n8128), .ZN(n7457) );
  NAND2_X1 U8635 ( .A1(n7458), .A2(n7457), .ZN(n7456) );
  NAND2_X1 U8636 ( .A1(n7702), .A2(n4425), .ZN(n7044) );
  NAND2_X1 U8637 ( .A1(n7456), .A2(n7044), .ZN(n7045) );
  INV_X1 U8638 ( .A(n7704), .ZN(n7087) );
  NAND2_X1 U8639 ( .A1(n8518), .A2(n7087), .ZN(n8129) );
  NAND2_X1 U8640 ( .A1(n8105), .A2(n8129), .ZN(n8257) );
  OAI21_X1 U8641 ( .B1(n7045), .B2(n8257), .A(n7089), .ZN(n7046) );
  INV_X1 U8642 ( .A(n7046), .ZN(n7497) );
  NAND2_X1 U8643 ( .A1(n7047), .A2(n7048), .ZN(n8113) );
  INV_X1 U8644 ( .A(n7457), .ZN(n8254) );
  NAND2_X1 U8645 ( .A1(n7460), .A2(n7092), .ZN(n7050) );
  XNOR2_X1 U8646 ( .A(n7050), .B(n8257), .ZN(n7051) );
  OAI222_X1 U8647 ( .A1(n8806), .A2(n7090), .B1(n8808), .B2(n7702), .C1(n7051), 
        .C2(n8803), .ZN(n7494) );
  INV_X1 U8648 ( .A(n7494), .ZN(n7056) );
  NAND2_X1 U8649 ( .A1(n7063), .A2(n7052), .ZN(n7469) );
  AND2_X1 U8650 ( .A1(n7471), .A2(n7704), .ZN(n7053) );
  NOR2_X1 U8651 ( .A1(n7425), .A2(n7053), .ZN(n7491) );
  NOR2_X1 U8652 ( .A1(n10062), .A2(n7087), .ZN(n7054) );
  AOI21_X1 U8653 ( .B1(n7491), .B2(n9683), .A(n7054), .ZN(n7055) );
  OAI211_X1 U8654 ( .C1(n8914), .C2(n7497), .A(n7056), .B(n7055), .ZN(n7079)
         );
  NAND2_X1 U8655 ( .A1(n7079), .A2(n4316), .ZN(n7057) );
  OAI21_X1 U8656 ( .B1(n4316), .B2(n7058), .A(n7057), .ZN(P2_U3463) );
  INV_X1 U8657 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n7069) );
  XNOR2_X1 U8658 ( .A(n7060), .B(n7049), .ZN(n8826) );
  INV_X1 U8659 ( .A(n8826), .ZN(n7067) );
  OAI21_X1 U8660 ( .B1(n4837), .B2(n7049), .A(n7061), .ZN(n7062) );
  AOI222_X1 U8661 ( .A1(n8793), .A2(n7062), .B1(n7025), .B2(n8788), .C1(n8519), 
        .C2(n8790), .ZN(n8830) );
  INV_X1 U8662 ( .A(n7063), .ZN(n7065) );
  INV_X1 U8663 ( .A(n7469), .ZN(n7064) );
  AOI21_X1 U8664 ( .B1(n8823), .B2(n7065), .A(n7064), .ZN(n8828) );
  AOI22_X1 U8665 ( .A1(n8828), .A2(n9683), .B1(n9677), .B2(n8823), .ZN(n7066)
         );
  OAI211_X1 U8666 ( .C1(n8914), .C2(n7067), .A(n8830), .B(n7066), .ZN(n7081)
         );
  NAND2_X1 U8667 ( .A1(n7081), .A2(n4316), .ZN(n7068) );
  OAI21_X1 U8668 ( .B1(n4316), .B2(n7069), .A(n7068), .ZN(P2_U3457) );
  NAND2_X1 U8669 ( .A1(n7071), .A2(n7070), .ZN(n7072) );
  INV_X1 U8670 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7078) );
  NAND2_X1 U8671 ( .A1(n10080), .A2(n7076), .ZN(n7077) );
  OAI21_X1 U8672 ( .B1(n10080), .B2(n7078), .A(n7077), .ZN(P2_U3521) );
  NAND2_X1 U8673 ( .A1(n7079), .A2(n10080), .ZN(n7080) );
  OAI21_X1 U8674 ( .B1(n10080), .B2(n6849), .A(n7080), .ZN(P2_U3524) );
  INV_X1 U8675 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7083) );
  NAND2_X1 U8676 ( .A1(n7081), .A2(n10080), .ZN(n7082) );
  OAI21_X1 U8677 ( .B1(n10080), .B2(n7083), .A(n7082), .ZN(P2_U3522) );
  INV_X1 U8678 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7086) );
  NAND2_X1 U8679 ( .A1(n10080), .A2(n7084), .ZN(n7085) );
  OAI21_X1 U8680 ( .B1(n10080), .B2(n7086), .A(n7085), .ZN(P2_U3520) );
  NAND2_X1 U8681 ( .A1(n7239), .A2(n7087), .ZN(n7088) );
  NAND2_X1 U8682 ( .A1(n10044), .A2(n8517), .ZN(n8131) );
  NAND2_X1 U8683 ( .A1(n8108), .A2(n8131), .ZN(n8256) );
  NAND2_X1 U8684 ( .A1(n7090), .A2(n10044), .ZN(n7091) );
  XNOR2_X1 U8685 ( .A(n8480), .B(n8516), .ZN(n8259) );
  XOR2_X1 U8686 ( .A(n7322), .B(n8259), .Z(n7639) );
  INV_X1 U8687 ( .A(n8480), .ZN(n8118) );
  AND2_X1 U8688 ( .A1(n8105), .A2(n7092), .ZN(n8107) );
  NAND2_X1 U8689 ( .A1(n7460), .A2(n8107), .ZN(n7430) );
  AND2_X1 U8690 ( .A1(n8131), .A2(n8129), .ZN(n8106) );
  NAND2_X1 U8691 ( .A1(n7430), .A2(n8106), .ZN(n7093) );
  NAND2_X1 U8692 ( .A1(n7093), .A2(n8108), .ZN(n7094) );
  OAI21_X1 U8693 ( .B1(n8259), .B2(n7094), .A(n7326), .ZN(n7097) );
  NAND2_X1 U8694 ( .A1(n8788), .A2(n8517), .ZN(n7096) );
  NAND2_X1 U8695 ( .A1(n8790), .A2(n8515), .ZN(n7095) );
  NAND2_X1 U8696 ( .A1(n7096), .A2(n7095), .ZN(n8476) );
  AOI21_X1 U8697 ( .B1(n7097), .B2(n8793), .A(n8476), .ZN(n7632) );
  NAND2_X1 U8698 ( .A1(n7426), .A2(n8118), .ZN(n7414) );
  OAI211_X1 U8699 ( .C1(n7426), .C2(n8118), .A(n9683), .B(n7414), .ZN(n7633)
         );
  OAI211_X1 U8700 ( .C1(n8118), .C2(n10062), .A(n7632), .B(n7633), .ZN(n7098)
         );
  AOI21_X1 U8701 ( .B1(n7639), .B2(n10068), .A(n7098), .ZN(n7120) );
  INV_X1 U8702 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7099) );
  OR2_X1 U8703 ( .A1(n10080), .A2(n7099), .ZN(n7100) );
  OAI21_X1 U8704 ( .B1(n7120), .B2(n10078), .A(n7100), .ZN(P2_U3526) );
  INV_X1 U8705 ( .A(n9124), .ZN(n9113) );
  OAI222_X1 U8706 ( .A1(n8318), .A2(n7102), .B1(n9443), .B2(n7101), .C1(
        P1_U3084), .C2(n9113), .ZN(P1_U3337) );
  INV_X1 U8707 ( .A(n7485), .ZN(n7109) );
  NAND2_X1 U8708 ( .A1(n10130), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7838) );
  INV_X1 U8709 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9758) );
  NOR2_X1 U8710 ( .A1(n7109), .A2(n9758), .ZN(n7103) );
  AOI21_X1 U8711 ( .B1(n9758), .B2(n7109), .A(n7103), .ZN(n7106) );
  OAI21_X1 U8712 ( .B1(n7111), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7104), .ZN(
        n7105) );
  NAND2_X1 U8713 ( .A1(n7106), .A2(n7105), .ZN(n7478) );
  OAI21_X1 U8714 ( .B1(n7106), .B2(n7105), .A(n7478), .ZN(n7107) );
  NAND2_X1 U8715 ( .A1(n9894), .A2(n7107), .ZN(n7108) );
  OAI211_X1 U8716 ( .C1(n9114), .C2(n7109), .A(n7838), .B(n7108), .ZN(n7116)
         );
  AOI21_X1 U8717 ( .B1(n7111), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7110), .ZN(
        n7114) );
  NOR2_X1 U8718 ( .A1(n7485), .A2(n9704), .ZN(n7112) );
  AOI21_X1 U8719 ( .B1(n7485), .B2(n9704), .A(n7112), .ZN(n7113) );
  NOR2_X1 U8720 ( .A1(n7114), .A2(n7113), .ZN(n7484) );
  AOI211_X1 U8721 ( .C1(n7114), .C2(n7113), .A(n7484), .B(n9872), .ZN(n7115)
         );
  AOI211_X1 U8722 ( .C1(P1_ADDR_REG_13__SCAN_IN), .C2(n9880), .A(n7116), .B(
        n7115), .ZN(n7117) );
  INV_X1 U8723 ( .A(n7117), .ZN(P1_U3254) );
  INV_X1 U8724 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n7118) );
  OR2_X1 U8725 ( .A1(n4316), .A2(n7118), .ZN(n7119) );
  OAI21_X1 U8726 ( .B1(n7120), .B2(n10070), .A(n7119), .ZN(P2_U3469) );
  NOR2_X1 U8727 ( .A1(n5151), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8326) );
  AOI21_X1 U8728 ( .B1(n7122), .B2(P2_REG1_REG_8__SCAN_IN), .A(n7121), .ZN(
        n7125) );
  INV_X1 U8729 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7123) );
  MUX2_X1 U8730 ( .A(n7123), .B(P2_REG1_REG_9__SCAN_IN), .S(n7293), .Z(n7124)
         );
  NOR2_X1 U8731 ( .A1(n7125), .A2(n7124), .ZN(n7287) );
  AOI211_X1 U8732 ( .C1(n7125), .C2(n7124), .A(n7287), .B(n9996), .ZN(n7126)
         );
  AOI211_X1 U8733 ( .C1(P2_ADDR_REG_9__SCAN_IN), .C2(n9994), .A(n8326), .B(
        n7126), .ZN(n7134) );
  OAI21_X1 U8734 ( .B1(n7128), .B2(n7338), .A(n7127), .ZN(n7132) );
  INV_X1 U8735 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7129) );
  MUX2_X1 U8736 ( .A(n7129), .B(P2_REG2_REG_9__SCAN_IN), .S(n7293), .Z(n7130)
         );
  INV_X1 U8737 ( .A(n7130), .ZN(n7131) );
  NAND2_X1 U8738 ( .A1(n7131), .A2(n7132), .ZN(n7294) );
  OAI211_X1 U8739 ( .C1(n7132), .C2(n7131), .A(n9992), .B(n7294), .ZN(n7133)
         );
  OAI211_X1 U8740 ( .C1(n9995), .C2(n7135), .A(n7134), .B(n7133), .ZN(P2_U3254) );
  INV_X1 U8741 ( .A(n7136), .ZN(n7139) );
  AOI22_X1 U8742 ( .A1(n9138), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9441), .ZN(n7137) );
  OAI21_X1 U8743 ( .B1(n7139), .B2(n9443), .A(n7137), .ZN(P1_U3336) );
  AOI22_X1 U8744 ( .A1(n8578), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n8943), .ZN(n7138) );
  OAI21_X1 U8745 ( .B1(n7139), .B2(n8946), .A(n7138), .ZN(P2_U3341) );
  OAI21_X1 U8746 ( .B1(n7141), .B2(n7144), .A(n7140), .ZN(n7194) );
  OAI22_X1 U8747 ( .A1(n7143), .A2(n9916), .B1(n7142), .B2(n9914), .ZN(n7148)
         );
  XNOR2_X1 U8748 ( .A(n7145), .B(n7144), .ZN(n7146) );
  NOR2_X1 U8749 ( .A1(n7146), .A2(n9732), .ZN(n7147) );
  AOI211_X1 U8750 ( .C1(n9735), .C2(n7194), .A(n7148), .B(n7147), .ZN(n7198)
         );
  NOR2_X1 U8751 ( .A1(n7150), .A2(n7149), .ZN(n7379) );
  NAND2_X1 U8752 ( .A1(n7379), .A2(n7151), .ZN(n7153) );
  NAND2_X1 U8753 ( .A1(n7579), .A2(n9431), .ZN(n7152) );
  NAND2_X2 U8754 ( .A1(n7153), .A2(n9925), .ZN(n9930) );
  INV_X2 U8755 ( .A(n9930), .ZN(n9736) );
  INV_X1 U8756 ( .A(n7154), .ZN(n7396) );
  INV_X1 U8757 ( .A(n7214), .ZN(n7155) );
  AOI21_X1 U8758 ( .B1(n7195), .B2(n7396), .A(n7155), .ZN(n7196) );
  AND2_X1 U8759 ( .A1(n7157), .A2(n7156), .ZN(n7158) );
  OAI22_X1 U8760 ( .A1(n9930), .A2(n5702), .B1(n7159), .B2(n9925), .ZN(n7162)
         );
  NOR2_X1 U8761 ( .A1(n9924), .A2(n7160), .ZN(n7161) );
  AOI211_X1 U8762 ( .C1(n7196), .C2(n9908), .A(n7162), .B(n7161), .ZN(n7166)
         );
  AND2_X1 U8763 ( .A1(n7163), .A2(n9272), .ZN(n7164) );
  AND2_X1 U8764 ( .A1(n9930), .A2(n7164), .ZN(n9909) );
  NAND2_X1 U8765 ( .A1(n7194), .A2(n9909), .ZN(n7165) );
  OAI211_X1 U8766 ( .C1(n7198), .C2(n9736), .A(n7166), .B(n7165), .ZN(P1_U3287) );
  AND2_X1 U8767 ( .A1(n7168), .A2(n7167), .ZN(n7169) );
  OAI21_X1 U8768 ( .B1(n7175), .B2(n7171), .A(n7170), .ZN(n9934) );
  OAI22_X1 U8769 ( .A1(n9924), .A2(n9936), .B1(n9930), .B2(n5654), .ZN(n7172)
         );
  INV_X1 U8770 ( .A(n7172), .ZN(n7183) );
  INV_X1 U8771 ( .A(n7173), .ZN(n7174) );
  XNOR2_X1 U8772 ( .A(n7175), .B(n7174), .ZN(n7176) );
  NAND2_X1 U8773 ( .A1(n7176), .A2(n9919), .ZN(n7178) );
  AOI22_X1 U8774 ( .A1(n9709), .A2(n5692), .B1(n6258), .B2(n9710), .ZN(n7177)
         );
  NAND2_X1 U8775 ( .A1(n7178), .A2(n7177), .ZN(n9937) );
  XNOR2_X1 U8776 ( .A(n9936), .B(n7235), .ZN(n7179) );
  NAND2_X1 U8777 ( .A1(n7179), .A2(n9395), .ZN(n9935) );
  OAI22_X1 U8778 ( .A1(n9935), .A2(n9272), .B1(n9925), .B2(n7180), .ZN(n7181)
         );
  OAI21_X1 U8779 ( .B1(n9937), .B2(n7181), .A(n9930), .ZN(n7182) );
  OAI211_X1 U8780 ( .C1(n9325), .C2(n9934), .A(n7183), .B(n7182), .ZN(P1_U3290) );
  NAND2_X1 U8781 ( .A1(n7185), .A2(n7184), .ZN(n7187) );
  XOR2_X1 U8782 ( .A(n7187), .B(n7186), .Z(n7193) );
  NOR2_X1 U8783 ( .A1(n9062), .A2(n9917), .ZN(n7188) );
  AOI211_X1 U8784 ( .C1(n9048), .C2(n9080), .A(n7189), .B(n7188), .ZN(n7190)
         );
  OAI21_X1 U8785 ( .B1(n9050), .B2(n7380), .A(n7190), .ZN(n7191) );
  AOI21_X1 U8786 ( .B1(n9052), .B2(n7382), .A(n7191), .ZN(n7192) );
  OAI21_X1 U8787 ( .B1(n7193), .B2(n9054), .A(n7192), .ZN(P1_U3211) );
  INV_X1 U8788 ( .A(n7194), .ZN(n7199) );
  AOI22_X1 U8789 ( .A1(n7196), .A2(n9395), .B1(n9745), .B2(n7195), .ZN(n7197)
         );
  OAI211_X1 U8790 ( .C1(n7199), .C2(n9659), .A(n7198), .B(n7197), .ZN(n7201)
         );
  NAND2_X1 U8791 ( .A1(n7201), .A2(n9990), .ZN(n7200) );
  OAI21_X1 U8792 ( .B1(n9990), .B2(n6739), .A(n7200), .ZN(P1_U3527) );
  INV_X1 U8793 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7203) );
  NAND2_X1 U8794 ( .A1(n7201), .A2(n9980), .ZN(n7202) );
  OAI21_X1 U8795 ( .B1(n9980), .B2(n7203), .A(n7202), .ZN(P1_U3466) );
  NAND2_X1 U8796 ( .A1(n7205), .A2(n7210), .ZN(n7206) );
  NAND2_X1 U8797 ( .A1(n7204), .A2(n7206), .ZN(n9946) );
  NAND2_X1 U8798 ( .A1(n7208), .A2(n7207), .ZN(n7209) );
  NAND2_X1 U8799 ( .A1(n7209), .A2(n7210), .ZN(n7273) );
  OAI21_X1 U8800 ( .B1(n7210), .B2(n7209), .A(n7273), .ZN(n7212) );
  OAI22_X1 U8801 ( .A1(n7403), .A2(n9916), .B1(n7388), .B2(n9914), .ZN(n7211)
         );
  AOI21_X1 U8802 ( .B1(n7212), .B2(n9919), .A(n7211), .ZN(n9952) );
  MUX2_X1 U8803 ( .A(n7213), .B(n9952), .S(n9930), .Z(n7220) );
  NOR2_X1 U8804 ( .A1(n9736), .A2(n9272), .ZN(n9238) );
  AOI21_X1 U8805 ( .B1(n7214), .B2(n7227), .A(n9973), .ZN(n7215) );
  NAND2_X1 U8806 ( .A1(n7215), .A2(n7280), .ZN(n9949) );
  INV_X1 U8807 ( .A(n9949), .ZN(n7218) );
  OAI22_X1 U8808 ( .A1(n9924), .A2(n7216), .B1(n7225), .B2(n9925), .ZN(n7217)
         );
  AOI21_X1 U8809 ( .B1(n9238), .B2(n7218), .A(n7217), .ZN(n7219) );
  OAI211_X1 U8810 ( .C1(n9325), .C2(n9946), .A(n7220), .B(n7219), .ZN(P1_U3286) );
  XNOR2_X1 U8811 ( .A(n7221), .B(n7222), .ZN(n7223) );
  NAND2_X1 U8812 ( .A1(n7223), .A2(n7224), .ZN(n7256) );
  OAI21_X1 U8813 ( .B1(n7224), .B2(n7223), .A(n7256), .ZN(n7233) );
  INV_X1 U8814 ( .A(n7225), .ZN(n7226) );
  NAND2_X1 U8815 ( .A1(n9066), .A2(n7226), .ZN(n7231) );
  AND2_X1 U8816 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9848) );
  AOI21_X1 U8817 ( .B1(n9048), .B2(n9082), .A(n9848), .ZN(n7230) );
  AND2_X1 U8818 ( .A1(n9745), .A2(n7227), .ZN(n9947) );
  NAND2_X1 U8819 ( .A1(n7318), .A2(n9947), .ZN(n7229) );
  NAND2_X1 U8820 ( .A1(n9024), .A2(n9080), .ZN(n7228) );
  NAND4_X1 U8821 ( .A1(n7231), .A2(n7230), .A3(n7229), .A4(n7228), .ZN(n7232)
         );
  AOI21_X1 U8822 ( .B1(n7233), .B2(n6223), .A(n7232), .ZN(n7234) );
  INV_X1 U8823 ( .A(n7234), .ZN(P1_U3225) );
  OAI21_X1 U8824 ( .B1(n9739), .B2(n9908), .A(n7235), .ZN(n7238) );
  AOI22_X1 U8825 ( .A1(n7236), .A2(n9930), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n9311), .ZN(n7237) );
  OAI211_X1 U8826 ( .C1(n5635), .C2(n9930), .A(n7238), .B(n7237), .ZN(P1_U3291) );
  MUX2_X1 U8827 ( .A(P2_U3152), .B(n8479), .S(n5047), .Z(n7241) );
  OAI22_X1 U8828 ( .A1(n8496), .A2(n7239), .B1(n4425), .B2(n7507), .ZN(n7240)
         );
  AOI211_X1 U8829 ( .C1(n8464), .C2(n8520), .A(n7241), .B(n7240), .ZN(n7251)
         );
  NOR3_X1 U8830 ( .A1(n8415), .A2(n7243), .A3(n7242), .ZN(n7249) );
  INV_X1 U8831 ( .A(n7245), .ZN(n7246) );
  AOI21_X1 U8832 ( .B1(n7244), .B2(n7246), .A(n8490), .ZN(n7248) );
  OAI21_X1 U8833 ( .B1(n7249), .B2(n7248), .A(n7247), .ZN(n7250) );
  NAND2_X1 U8834 ( .A1(n7251), .A2(n7250), .ZN(P2_U3220) );
  INV_X1 U8835 ( .A(n9885), .ZN(n9135) );
  INV_X1 U8836 ( .A(n7252), .ZN(n7254) );
  INV_X1 U8837 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7253) );
  OAI222_X1 U8838 ( .A1(n9135), .A2(n10130), .B1(n9443), .B2(n7254), .C1(n7253), .C2(n8318), .ZN(P1_U3335) );
  INV_X1 U8839 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7255) );
  INV_X1 U8840 ( .A(n8583), .ZN(n8589) );
  OAI222_X1 U8841 ( .A1(n8947), .A2(n7255), .B1(n8946), .B2(n7254), .C1(
        P2_U3152), .C2(n8589), .ZN(P2_U3340) );
  OAI21_X1 U8842 ( .B1(n7257), .B2(n7221), .A(n7256), .ZN(n7261) );
  XNOR2_X1 U8843 ( .A(n7259), .B(n7258), .ZN(n7260) );
  XNOR2_X1 U8844 ( .A(n7261), .B(n7260), .ZN(n7268) );
  NOR2_X1 U8845 ( .A1(n9062), .A2(n7262), .ZN(n7263) );
  AOI211_X1 U8846 ( .C1(n9048), .C2(n9081), .A(n7264), .B(n7263), .ZN(n7265)
         );
  OAI21_X1 U8847 ( .B1(n9050), .B2(n7282), .A(n7265), .ZN(n7266) );
  AOI21_X1 U8848 ( .B1(n9052), .B2(n7281), .A(n7266), .ZN(n7267) );
  OAI21_X1 U8849 ( .B1(n7268), .B2(n9054), .A(n7267), .ZN(P1_U3237) );
  NAND2_X1 U8850 ( .A1(n7269), .A2(n7274), .ZN(n7270) );
  NAND2_X1 U8851 ( .A1(n7271), .A2(n7270), .ZN(n9958) );
  INV_X1 U8852 ( .A(n9958), .ZN(n7286) );
  INV_X1 U8853 ( .A(n9909), .ZN(n7410) );
  NAND2_X1 U8854 ( .A1(n7273), .A2(n7272), .ZN(n7275) );
  XNOR2_X1 U8855 ( .A(n7275), .B(n6266), .ZN(n7278) );
  NAND2_X1 U8856 ( .A1(n9958), .A2(n9735), .ZN(n7277) );
  AOI22_X1 U8857 ( .A1(n9081), .A2(n9710), .B1(n9709), .B2(n9079), .ZN(n7276)
         );
  OAI211_X1 U8858 ( .C1(n9732), .C2(n7278), .A(n7277), .B(n7276), .ZN(n9956)
         );
  MUX2_X1 U8859 ( .A(n9956), .B(P1_REG2_REG_6__SCAN_IN), .S(n9736), .Z(n7279)
         );
  INV_X1 U8860 ( .A(n7279), .ZN(n7285) );
  AOI21_X1 U8861 ( .B1(n7281), .B2(n7280), .A(n7375), .ZN(n9953) );
  OAI22_X1 U8862 ( .A1(n9924), .A2(n9954), .B1(n7282), .B2(n9925), .ZN(n7283)
         );
  AOI21_X1 U8863 ( .B1(n9953), .B2(n9908), .A(n7283), .ZN(n7284) );
  OAI211_X1 U8864 ( .C1(n7286), .C2(n7410), .A(n7285), .B(n7284), .ZN(P1_U3285) );
  NOR2_X1 U8865 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9586), .ZN(n7292) );
  INV_X1 U8866 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7288) );
  MUX2_X1 U8867 ( .A(n7288), .B(P2_REG1_REG_10__SCAN_IN), .S(n7649), .Z(n7289)
         );
  AOI211_X1 U8868 ( .C1(n7290), .C2(n7289), .A(n7648), .B(n9996), .ZN(n7291)
         );
  AOI211_X1 U8869 ( .C1(P2_ADDR_REG_10__SCAN_IN), .C2(n9994), .A(n7292), .B(
        n7291), .ZN(n7301) );
  NAND2_X1 U8870 ( .A1(n7293), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7295) );
  NAND2_X1 U8871 ( .A1(n7295), .A2(n7294), .ZN(n7299) );
  INV_X1 U8872 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7296) );
  MUX2_X1 U8873 ( .A(n7296), .B(P2_REG2_REG_10__SCAN_IN), .S(n7649), .Z(n7297)
         );
  INV_X1 U8874 ( .A(n7297), .ZN(n7298) );
  NAND2_X1 U8875 ( .A1(n7298), .A2(n7299), .ZN(n7641) );
  OAI211_X1 U8876 ( .C1(n7299), .C2(n7298), .A(n9992), .B(n7641), .ZN(n7300)
         );
  OAI211_X1 U8877 ( .C1(n9995), .C2(n7302), .A(n7301), .B(n7300), .ZN(P2_U3255) );
  INV_X1 U8878 ( .A(n7303), .ZN(n7305) );
  OAI222_X1 U8879 ( .A1(n10130), .A2(n9222), .B1(n9443), .B2(n7305), .C1(n7304), .C2(n8318), .ZN(P1_U3334) );
  OAI222_X1 U8880 ( .A1(n8947), .A2(n7306), .B1(n8946), .B2(n7305), .C1(n8815), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  NAND2_X1 U8881 ( .A1(n7307), .A2(n7308), .ZN(n7309) );
  XOR2_X1 U8882 ( .A(n7310), .B(n7309), .Z(n7320) );
  NAND2_X1 U8883 ( .A1(n7450), .A2(n9745), .ZN(n9965) );
  INV_X1 U8884 ( .A(n9965), .ZN(n7317) );
  INV_X1 U8885 ( .A(n7311), .ZN(n7449) );
  NAND2_X1 U8886 ( .A1(n9066), .A2(n7449), .ZN(n7314) );
  AOI21_X1 U8887 ( .B1(n9048), .B2(n9079), .A(n7312), .ZN(n7313) );
  OAI211_X1 U8888 ( .C1(n7315), .C2(n9062), .A(n7314), .B(n7313), .ZN(n7316)
         );
  AOI21_X1 U8889 ( .B1(n7318), .B2(n7317), .A(n7316), .ZN(n7319) );
  OAI21_X1 U8890 ( .B1(n7320), .B2(n9054), .A(n7319), .ZN(P1_U3219) );
  NOR2_X1 U8891 ( .A1(n8480), .A2(n8516), .ZN(n7321) );
  NAND2_X1 U8892 ( .A1(n8480), .A2(n8516), .ZN(n7323) );
  INV_X1 U8893 ( .A(n8515), .ZN(n8413) );
  OR2_X1 U8894 ( .A1(n7626), .A2(n8413), .ZN(n8148) );
  NAND2_X1 U8895 ( .A1(n7626), .A2(n8413), .ZN(n8141) );
  INV_X1 U8896 ( .A(n8514), .ZN(n8330) );
  OR2_X1 U8897 ( .A1(n8419), .A2(n8330), .ZN(n8142) );
  NAND2_X1 U8898 ( .A1(n8419), .A2(n8330), .ZN(n8150) );
  NAND2_X1 U8899 ( .A1(n7324), .A2(n8261), .ZN(n7325) );
  AND2_X1 U8900 ( .A1(n7530), .A2(n7325), .ZN(n7350) );
  INV_X1 U8901 ( .A(n7760), .ZN(n7459) );
  INV_X1 U8902 ( .A(n8516), .ZN(n8137) );
  NAND2_X1 U8903 ( .A1(n8480), .A2(n8137), .ZN(n8109) );
  INV_X1 U8904 ( .A(n8261), .ZN(n7328) );
  NAND2_X1 U8905 ( .A1(n7327), .A2(n8261), .ZN(n7535) );
  NAND2_X1 U8906 ( .A1(n7329), .A2(n7328), .ZN(n7330) );
  NAND2_X1 U8907 ( .A1(n7535), .A2(n7330), .ZN(n7331) );
  NAND2_X1 U8908 ( .A1(n7331), .A2(n8793), .ZN(n7333) );
  AOI22_X1 U8909 ( .A1(n8788), .A2(n8515), .B1(n8790), .B2(n8513), .ZN(n7332)
         );
  NAND2_X1 U8910 ( .A1(n7333), .A2(n7332), .ZN(n7334) );
  AOI21_X1 U8911 ( .B1(n7350), .B2(n7459), .A(n7334), .ZN(n7353) );
  INV_X1 U8912 ( .A(n7335), .ZN(n7336) );
  MUX2_X1 U8913 ( .A(n7338), .B(n7353), .S(n10009), .Z(n7349) );
  OR2_X1 U8914 ( .A1(n7339), .A2(n8815), .ZN(n7412) );
  INV_X1 U8915 ( .A(n7412), .ZN(n7340) );
  INV_X1 U8916 ( .A(n8419), .ZN(n7346) );
  INV_X1 U8917 ( .A(n7341), .ZN(n10004) );
  OR2_X1 U8918 ( .A1(n7414), .A2(n7626), .ZN(n7416) );
  AND2_X1 U8919 ( .A1(n7416), .A2(n8419), .ZN(n7343) );
  NOR2_X1 U8920 ( .A1(n7541), .A2(n7343), .ZN(n7351) );
  NAND2_X1 U8921 ( .A1(n8829), .A2(n7351), .ZN(n7345) );
  NAND2_X1 U8922 ( .A1(n8827), .A2(n8420), .ZN(n7344) );
  OAI211_X1 U8923 ( .C1(n7346), .C2(n10018), .A(n7345), .B(n7344), .ZN(n7347)
         );
  AOI21_X1 U8924 ( .B1(n7350), .B2(n7767), .A(n7347), .ZN(n7348) );
  NAND2_X1 U8925 ( .A1(n7349), .A2(n7348), .ZN(P2_U3288) );
  INV_X1 U8926 ( .A(n7350), .ZN(n7354) );
  AOI22_X1 U8927 ( .A1(n7351), .A2(n9683), .B1(n9677), .B2(n8419), .ZN(n7352)
         );
  OAI211_X1 U8928 ( .C1(n7354), .C2(n9685), .A(n7353), .B(n7352), .ZN(n7356)
         );
  NAND2_X1 U8929 ( .A1(n7356), .A2(n10080), .ZN(n7355) );
  OAI21_X1 U8930 ( .B1(n10080), .B2(n6955), .A(n7355), .ZN(P2_U3528) );
  INV_X1 U8931 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7358) );
  NAND2_X1 U8932 ( .A1(n7356), .A2(n4316), .ZN(n7357) );
  OAI21_X1 U8933 ( .B1(n4316), .B2(n7358), .A(n7357), .ZN(P2_U3475) );
  OR2_X1 U8934 ( .A1(n7359), .A2(n7573), .ZN(n7571) );
  AOI21_X1 U8935 ( .B1(n7571), .B2(n7360), .A(n8490), .ZN(n7366) );
  INV_X1 U8936 ( .A(n7361), .ZN(n7362) );
  NOR3_X1 U8937 ( .A1(n8415), .A2(n7362), .A3(n8329), .ZN(n7365) );
  OR2_X1 U8938 ( .A1(n7359), .A2(n7363), .ZN(n8304) );
  AND2_X1 U8939 ( .A1(n8304), .A2(n7364), .ZN(n8298) );
  OAI21_X1 U8940 ( .B1(n7366), .B2(n7365), .A(n8298), .ZN(n7372) );
  INV_X1 U8941 ( .A(n7368), .ZN(n7683) );
  OAI22_X1 U8942 ( .A1(n8494), .A2(n7683), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5187), .ZN(n7370) );
  INV_X1 U8943 ( .A(n8510), .ZN(n7756) );
  OAI22_X1 U8944 ( .A1(n8329), .A2(n8495), .B1(n8496), .B2(n7756), .ZN(n7369)
         );
  AOI211_X1 U8945 ( .C1(n7367), .C2(n8461), .A(n7370), .B(n7369), .ZN(n7371)
         );
  NAND2_X1 U8946 ( .A1(n7372), .A2(n7371), .ZN(P2_U3238) );
  INV_X1 U8947 ( .A(n9325), .ZN(n7391) );
  OAI21_X1 U8948 ( .B1(n7374), .B2(n7386), .A(n7373), .ZN(n9963) );
  OAI21_X1 U8949 ( .B1(n7375), .B2(n9960), .A(n9395), .ZN(n7376) );
  OR2_X1 U8950 ( .A1(n7376), .A2(n7448), .ZN(n9959) );
  NOR2_X1 U8951 ( .A1(n7377), .A2(n9272), .ZN(n7378) );
  AND2_X1 U8952 ( .A1(n7379), .A2(n7378), .ZN(n7987) );
  INV_X1 U8953 ( .A(n7987), .ZN(n7620) );
  INV_X1 U8954 ( .A(n7380), .ZN(n7381) );
  AOI22_X1 U8955 ( .A1(n9739), .A2(n7382), .B1(n7381), .B2(n9311), .ZN(n7383)
         );
  OAI21_X1 U8956 ( .B1(n9959), .B2(n7620), .A(n7383), .ZN(n7390) );
  INV_X1 U8957 ( .A(n7441), .ZN(n7384) );
  AOI21_X1 U8958 ( .B1(n7386), .B2(n7385), .A(n7384), .ZN(n7387) );
  OAI222_X1 U8959 ( .A1(n9916), .A2(n7388), .B1(n9914), .B2(n9917), .C1(n9732), 
        .C2(n7387), .ZN(n9961) );
  MUX2_X1 U8960 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n9961), .S(n9930), .Z(n7389)
         );
  AOI211_X1 U8961 ( .C1(n7391), .C2(n9963), .A(n7390), .B(n7389), .ZN(n7392)
         );
  INV_X1 U8962 ( .A(n7392), .ZN(P1_U3284) );
  OAI21_X1 U8963 ( .B1(n7394), .B2(n7401), .A(n7393), .ZN(n9944) );
  INV_X1 U8964 ( .A(n9944), .ZN(n7411) );
  OAI22_X1 U8965 ( .A1(n9930), .A2(n6723), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9925), .ZN(n7399) );
  INV_X1 U8966 ( .A(n9238), .ZN(n7965) );
  INV_X1 U8967 ( .A(n7395), .ZN(n7397) );
  OAI211_X1 U8968 ( .C1(n9941), .C2(n7397), .A(n7396), .B(n9395), .ZN(n9940)
         );
  NOR2_X1 U8969 ( .A1(n7965), .A2(n9940), .ZN(n7398) );
  AOI211_X1 U8970 ( .C1(n9739), .C2(n7400), .A(n7399), .B(n7398), .ZN(n7409)
         );
  XNOR2_X1 U8971 ( .A(n7402), .B(n7401), .ZN(n7407) );
  OAI22_X1 U8972 ( .A1(n7404), .A2(n9916), .B1(n7403), .B2(n9914), .ZN(n7405)
         );
  AOI21_X1 U8973 ( .B1(n9944), .B2(n9735), .A(n7405), .ZN(n7406) );
  OAI21_X1 U8974 ( .B1(n9732), .B2(n7407), .A(n7406), .ZN(n9942) );
  NAND2_X1 U8975 ( .A1(n9942), .A2(n9930), .ZN(n7408) );
  OAI211_X1 U8976 ( .C1(n7411), .C2(n7410), .A(n7409), .B(n7408), .ZN(P1_U3288) );
  NAND2_X1 U8977 ( .A1(n7760), .A2(n7412), .ZN(n10014) );
  INV_X1 U8978 ( .A(n8798), .ZN(n8825) );
  XNOR2_X1 U8979 ( .A(n7413), .B(n8260), .ZN(n10052) );
  INV_X1 U8980 ( .A(n7626), .ZN(n10048) );
  NAND2_X1 U8981 ( .A1(n7414), .A2(n7626), .ZN(n7415) );
  NAND2_X1 U8982 ( .A1(n7416), .A2(n7415), .ZN(n10049) );
  INV_X1 U8983 ( .A(n10049), .ZN(n7417) );
  AOI22_X1 U8984 ( .A1(n8829), .A2(n7417), .B1(n7627), .B2(n8827), .ZN(n7418)
         );
  OAI21_X1 U8985 ( .B1(n10048), .B2(n10018), .A(n7418), .ZN(n7422) );
  XOR2_X1 U8986 ( .A(n8260), .B(n7419), .Z(n7420) );
  OAI222_X1 U8987 ( .A1(n8808), .A2(n8137), .B1(n8806), .B2(n8330), .C1(n7420), 
        .C2(n8803), .ZN(n10050) );
  MUX2_X1 U8988 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10050), .S(n10009), .Z(n7421) );
  AOI211_X1 U8989 ( .C1(n8825), .C2(n10052), .A(n7422), .B(n7421), .ZN(n7423)
         );
  INV_X1 U8990 ( .A(n7423), .ZN(P2_U3289) );
  XNOR2_X1 U8991 ( .A(n7424), .B(n8256), .ZN(n10046) );
  OAI21_X1 U8992 ( .B1(n7425), .B2(n10044), .A(n9683), .ZN(n7427) );
  NOR2_X1 U8993 ( .A1(n7427), .A2(n7426), .ZN(n10041) );
  AOI22_X1 U8994 ( .A1(n10011), .A2(n10041), .B1(n8450), .B2(n8827), .ZN(n7428) );
  OAI21_X1 U8995 ( .B1(n10044), .B2(n10018), .A(n7428), .ZN(n7429) );
  AOI21_X1 U8996 ( .B1(n8825), .B2(n10046), .A(n7429), .ZN(n7436) );
  NAND2_X1 U8997 ( .A1(n7430), .A2(n8129), .ZN(n7431) );
  XNOR2_X1 U8998 ( .A(n7431), .B(n8256), .ZN(n7434) );
  NAND2_X1 U8999 ( .A1(n8788), .A2(n8518), .ZN(n7433) );
  NAND2_X1 U9000 ( .A1(n8790), .A2(n8516), .ZN(n7432) );
  NAND2_X1 U9001 ( .A1(n7433), .A2(n7432), .ZN(n8449) );
  AOI21_X1 U9002 ( .B1(n7434), .B2(n8793), .A(n8449), .ZN(n10043) );
  MUX2_X1 U9003 ( .A(n6906), .B(n10043), .S(n10009), .Z(n7435) );
  NAND2_X1 U9004 ( .A1(n7436), .A2(n7435), .ZN(P2_U3291) );
  INV_X1 U9005 ( .A(n7437), .ZN(n7438) );
  AOI21_X1 U9006 ( .B1(n7442), .B2(n7439), .A(n7438), .ZN(n9970) );
  INV_X1 U9007 ( .A(n9970), .ZN(n7455) );
  NAND2_X1 U9008 ( .A1(n7441), .A2(n7440), .ZN(n7443) );
  XNOR2_X1 U9009 ( .A(n7443), .B(n7442), .ZN(n7444) );
  NAND2_X1 U9010 ( .A1(n7444), .A2(n9919), .ZN(n7446) );
  AOI22_X1 U9011 ( .A1(n9709), .A2(n9077), .B1(n9079), .B2(n9710), .ZN(n7445)
         );
  NAND2_X1 U9012 ( .A1(n7446), .A2(n7445), .ZN(n9968) );
  OAI21_X1 U9013 ( .B1(n7448), .B2(n7447), .A(n9903), .ZN(n9966) );
  INV_X1 U9014 ( .A(n9908), .ZN(n9159) );
  AOI22_X1 U9015 ( .A1(n9736), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7449), .B2(
        n9311), .ZN(n7452) );
  NAND2_X1 U9016 ( .A1(n9739), .A2(n7450), .ZN(n7451) );
  OAI211_X1 U9017 ( .C1(n9966), .C2(n9159), .A(n7452), .B(n7451), .ZN(n7453)
         );
  AOI21_X1 U9018 ( .B1(n9968), .B2(n9930), .A(n7453), .ZN(n7454) );
  OAI21_X1 U9019 ( .B1(n7455), .B2(n9325), .A(n7454), .ZN(P1_U3283) );
  OAI21_X1 U9020 ( .B1(n7458), .B2(n7457), .A(n7456), .ZN(n10037) );
  NAND2_X1 U9021 ( .A1(n10037), .A2(n7459), .ZN(n7467) );
  OAI21_X1 U9022 ( .B1(n8254), .B2(n7461), .A(n7460), .ZN(n7465) );
  NAND2_X1 U9023 ( .A1(n8788), .A2(n8520), .ZN(n7463) );
  NAND2_X1 U9024 ( .A1(n8790), .A2(n8518), .ZN(n7462) );
  NAND2_X1 U9025 ( .A1(n7463), .A2(n7462), .ZN(n7464) );
  AOI21_X1 U9026 ( .B1(n7465), .B2(n8793), .A(n7464), .ZN(n7466) );
  AND2_X1 U9027 ( .A1(n7467), .A2(n7466), .ZN(n10039) );
  AOI22_X1 U9028 ( .A1(n8824), .A2(n7468), .B1(n7767), .B2(n10037), .ZN(n7475)
         );
  NAND2_X1 U9029 ( .A1(n7469), .A2(n7468), .ZN(n7470) );
  AND3_X1 U9030 ( .A1(n7471), .A2(n9683), .A3(n7470), .ZN(n10034) );
  OAI22_X1 U9031 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(n10025), .B1(n7472), .B2(
        n10009), .ZN(n7473) );
  AOI21_X1 U9032 ( .B1(n10011), .B2(n10034), .A(n7473), .ZN(n7474) );
  OAI211_X1 U9033 ( .C1(n10022), .C2(n10039), .A(n7475), .B(n7474), .ZN(
        P2_U3293) );
  NAND2_X1 U9034 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3084), .ZN(n7483) );
  OR2_X1 U9035 ( .A1(n7743), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7477) );
  NAND2_X1 U9036 ( .A1(n7743), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7476) );
  AND2_X1 U9037 ( .A1(n7477), .A2(n7476), .ZN(n7480) );
  OAI21_X1 U9038 ( .B1(n7485), .B2(P1_REG1_REG_13__SCAN_IN), .A(n7478), .ZN(
        n7479) );
  NAND2_X1 U9039 ( .A1(n7480), .A2(n7479), .ZN(n7742) );
  OAI21_X1 U9040 ( .B1(n7480), .B2(n7479), .A(n7742), .ZN(n7481) );
  NAND2_X1 U9041 ( .A1(n9894), .A2(n7481), .ZN(n7482) );
  OAI211_X1 U9042 ( .C1(n9114), .C2(n7736), .A(n7483), .B(n7482), .ZN(n7489)
         );
  INV_X1 U9043 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7486) );
  AOI211_X1 U9044 ( .C1(n7487), .C2(n7486), .A(n7738), .B(n9872), .ZN(n7488)
         );
  AOI211_X1 U9045 ( .C1(P1_ADDR_REG_14__SCAN_IN), .C2(n9880), .A(n7489), .B(
        n7488), .ZN(n7490) );
  INV_X1 U9046 ( .A(n7490), .ZN(P1_U3255) );
  AOI22_X1 U9047 ( .A1(n8829), .A2(n7491), .B1(n8824), .B2(n7704), .ZN(n7496)
         );
  INV_X1 U9048 ( .A(n7492), .ZN(n7707) );
  OAI22_X1 U9049 ( .A1(n10009), .A2(n6859), .B1(n7707), .B2(n10025), .ZN(n7493) );
  AOI21_X1 U9050 ( .B1(n10009), .B2(n7494), .A(n7493), .ZN(n7495) );
  OAI211_X1 U9051 ( .C1(n7497), .C2(n8798), .A(n7496), .B(n7495), .ZN(P2_U3292) );
  OR2_X1 U9052 ( .A1(n7359), .A2(n7498), .ZN(n7499) );
  AND2_X1 U9053 ( .A1(n7500), .A2(n7499), .ZN(n7502) );
  INV_X1 U9054 ( .A(n7501), .ZN(n7583) );
  AOI211_X1 U9055 ( .C1(n7503), .C2(n7502), .A(n8490), .B(n7583), .ZN(n7509)
         );
  INV_X1 U9056 ( .A(n7504), .ZN(n9686) );
  AOI22_X1 U9057 ( .A1(n8464), .A2(n8510), .B1(n8465), .B2(n8508), .ZN(n7506)
         );
  AOI22_X1 U9058 ( .A1(n8479), .A2(n7763), .B1(P2_U3152), .B2(
        P2_REG3_REG_13__SCAN_IN), .ZN(n7505) );
  OAI211_X1 U9059 ( .C1(n9686), .C2(n7507), .A(n7506), .B(n7505), .ZN(n7508)
         );
  OR2_X1 U9060 ( .A1(n7509), .A2(n7508), .ZN(P2_U3236) );
  INV_X1 U9061 ( .A(n7510), .ZN(n7548) );
  OAI222_X1 U9062 ( .A1(n8946), .A2(n7548), .B1(P2_U3152), .B2(n8252), .C1(
        n7511), .C2(n8947), .ZN(P2_U3338) );
  OAI21_X1 U9063 ( .B1(n7514), .B2(n7513), .A(n7512), .ZN(n7515) );
  AOI22_X1 U9064 ( .A1(n10003), .A2(n8500), .B1(n8474), .B2(n7515), .ZN(n7519)
         );
  OR2_X1 U9065 ( .A1(n7516), .A2(P2_U3152), .ZN(n8466) );
  AOI22_X1 U9066 ( .A1(n8477), .A2(n7517), .B1(n8466), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n7518) );
  NAND2_X1 U9067 ( .A1(n7519), .A2(n7518), .ZN(P2_U3224) );
  AOI21_X1 U9068 ( .B1(n7522), .B2(n7521), .A(n5820), .ZN(n7528) );
  INV_X1 U9069 ( .A(n9926), .ZN(n7523) );
  NAND2_X1 U9070 ( .A1(n9066), .A2(n7523), .ZN(n7525) );
  AND2_X1 U9071 ( .A1(n10130), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9864) );
  AOI21_X1 U9072 ( .B1(n9048), .B2(n9078), .A(n9864), .ZN(n7524) );
  OAI211_X1 U9073 ( .C1(n9915), .C2(n9062), .A(n7525), .B(n7524), .ZN(n7526)
         );
  AOI21_X1 U9074 ( .B1(n9052), .B2(n9904), .A(n7526), .ZN(n7527) );
  OAI21_X1 U9075 ( .B1(n7528), .B2(n9054), .A(n7527), .ZN(P1_U3229) );
  INV_X1 U9076 ( .A(n8513), .ZN(n7529) );
  OR2_X1 U9077 ( .A1(n8333), .A2(n7529), .ZN(n8143) );
  NAND2_X1 U9078 ( .A1(n8333), .A2(n7529), .ZN(n8160) );
  NAND2_X1 U9079 ( .A1(n7532), .A2(n7531), .ZN(n7598) );
  INV_X1 U9080 ( .A(n7598), .ZN(n7533) );
  AOI21_X1 U9081 ( .B1(n8263), .B2(n7534), .A(n7533), .ZN(n10054) );
  INV_X1 U9082 ( .A(n7767), .ZN(n8821) );
  NAND2_X1 U9083 ( .A1(n7535), .A2(n8150), .ZN(n7536) );
  OAI21_X1 U9084 ( .B1(n8263), .B2(n7536), .A(n7594), .ZN(n7538) );
  OAI22_X1 U9085 ( .A1(n8330), .A2(n8808), .B1(n8806), .B2(n8329), .ZN(n7537)
         );
  AOI21_X1 U9086 ( .B1(n7538), .B2(n8793), .A(n7537), .ZN(n7539) );
  OAI21_X1 U9087 ( .B1(n10054), .B2(n7760), .A(n7539), .ZN(n10057) );
  NAND2_X1 U9088 ( .A1(n10057), .A2(n10009), .ZN(n7546) );
  INV_X1 U9089 ( .A(n7540), .ZN(n8328) );
  OAI22_X1 U9090 ( .A1(n10009), .A2(n7129), .B1(n8328), .B2(n10025), .ZN(n7544) );
  INV_X1 U9091 ( .A(n8333), .ZN(n10055) );
  NOR2_X1 U9092 ( .A1(n7541), .A2(n10055), .ZN(n7542) );
  OR2_X1 U9093 ( .A1(n7602), .A2(n7542), .ZN(n10056) );
  NOR2_X1 U9094 ( .A1(n10019), .A2(n10056), .ZN(n7543) );
  AOI211_X1 U9095 ( .C1(n8824), .C2(n8333), .A(n7544), .B(n7543), .ZN(n7545)
         );
  OAI211_X1 U9096 ( .C1(n10054), .C2(n8821), .A(n7546), .B(n7545), .ZN(
        P2_U3287) );
  OAI222_X1 U9097 ( .A1(n7549), .A2(P1_U3084), .B1(n9443), .B2(n7548), .C1(
        n7547), .C2(n8318), .ZN(P1_U3333) );
  OAI22_X1 U9098 ( .A1(n8415), .A2(n7550), .B1(n10017), .B2(n8490), .ZN(n7552)
         );
  NAND2_X1 U9099 ( .A1(n7552), .A2(n7551), .ZN(n7555) );
  INV_X1 U9100 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10024) );
  AOI22_X1 U9101 ( .A1(n8500), .A2(n7553), .B1(n8466), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n7554) );
  OAI211_X1 U9102 ( .C1(n8496), .C2(n7556), .A(n7555), .B(n7554), .ZN(P2_U3234) );
  XNOR2_X1 U9103 ( .A(n7558), .B(n7557), .ZN(n7559) );
  XNOR2_X1 U9104 ( .A(n7560), .B(n7559), .ZN(n7566) );
  NOR2_X1 U9105 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7561), .ZN(n9877) );
  NOR2_X1 U9106 ( .A1(n9062), .A2(n7826), .ZN(n7562) );
  AOI211_X1 U9107 ( .C1(n9048), .C2(n9077), .A(n9877), .B(n7562), .ZN(n7563)
         );
  OAI21_X1 U9108 ( .B1(n9050), .B2(n7616), .A(n7563), .ZN(n7564) );
  AOI21_X1 U9109 ( .B1(n9052), .B2(n9660), .A(n7564), .ZN(n7565) );
  OAI21_X1 U9110 ( .B1(n7566), .B2(n9054), .A(n7565), .ZN(P1_U3215) );
  INV_X1 U9111 ( .A(n7567), .ZN(n7599) );
  NAND2_X1 U9112 ( .A1(n8788), .A2(n8513), .ZN(n7569) );
  NAND2_X1 U9113 ( .A1(n8790), .A2(n8511), .ZN(n7568) );
  NAND2_X1 U9114 ( .A1(n7569), .A2(n7568), .ZN(n7595) );
  AOI22_X1 U9115 ( .A1(n8477), .A2(n7595), .B1(P2_REG3_REG_10__SCAN_IN), .B2(
        P2_U3152), .ZN(n7570) );
  OAI21_X1 U9116 ( .B1(n7599), .B2(n8494), .A(n7570), .ZN(n7575) );
  INV_X1 U9117 ( .A(n7571), .ZN(n7572) );
  AOI211_X1 U9118 ( .C1(n7573), .C2(n7359), .A(n8490), .B(n7572), .ZN(n7574)
         );
  AOI211_X1 U9119 ( .C1(n7676), .C2(n8500), .A(n7575), .B(n7574), .ZN(n7576)
         );
  INV_X1 U9120 ( .A(n7576), .ZN(P2_U3219) );
  INV_X1 U9121 ( .A(n7577), .ZN(n7690) );
  INV_X1 U9122 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7578) );
  OAI222_X1 U9123 ( .A1(n7579), .A2(n10130), .B1(n9443), .B2(n7690), .C1(n7578), .C2(n8318), .ZN(P1_U3332) );
  INV_X1 U9124 ( .A(n7580), .ZN(n7581) );
  INV_X1 U9125 ( .A(n8509), .ZN(n7751) );
  NOR3_X1 U9126 ( .A1(n7581), .A2(n7751), .A3(n8415), .ZN(n7582) );
  AOI21_X1 U9127 ( .B1(n7583), .B2(n8474), .A(n7582), .ZN(n7593) );
  INV_X1 U9128 ( .A(n8477), .ZN(n7587) );
  NAND2_X1 U9129 ( .A1(n8790), .A2(n8507), .ZN(n7585) );
  NAND2_X1 U9130 ( .A1(n8788), .A2(n8509), .ZN(n7584) );
  AND2_X1 U9131 ( .A1(n7585), .A2(n7584), .ZN(n7774) );
  NAND2_X1 U9132 ( .A1(n8479), .A2(n7777), .ZN(n7586) );
  NAND2_X1 U9133 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7878) );
  OAI211_X1 U9134 ( .C1(n7587), .C2(n7774), .A(n7586), .B(n7878), .ZN(n7590)
         );
  NOR2_X1 U9135 ( .A1(n7588), .A2(n8490), .ZN(n7589) );
  AOI211_X1 U9136 ( .C1(n8177), .C2(n8461), .A(n7590), .B(n7589), .ZN(n7591)
         );
  OAI21_X1 U9137 ( .B1(n7593), .B2(n7592), .A(n7591), .ZN(P2_U3217) );
  OR2_X1 U9138 ( .A1(n7676), .A2(n8329), .ZN(n8145) );
  NAND2_X1 U9139 ( .A1(n7676), .A2(n8329), .ZN(n8152) );
  NAND2_X1 U9140 ( .A1(n8145), .A2(n8152), .ZN(n8265) );
  XOR2_X1 U9141 ( .A(n7679), .B(n8265), .Z(n7596) );
  AOI21_X1 U9142 ( .B1(n7596), .B2(n8793), .A(n7595), .ZN(n7670) );
  OR2_X1 U9143 ( .A1(n8333), .A2(n8513), .ZN(n7597) );
  NAND2_X1 U9144 ( .A1(n7717), .A2(n8265), .ZN(n7677) );
  OAI21_X1 U9145 ( .B1(n7717), .B2(n8265), .A(n7677), .ZN(n7671) );
  OAI22_X1 U9146 ( .A1(n10009), .A2(n7296), .B1(n7599), .B2(n10025), .ZN(n7600) );
  AOI21_X1 U9147 ( .B1(n8824), .B2(n7676), .A(n7600), .ZN(n7605) );
  INV_X1 U9148 ( .A(n7676), .ZN(n7601) );
  NAND2_X1 U9149 ( .A1(n7602), .A2(n7601), .ZN(n7681) );
  OR2_X1 U9150 ( .A1(n7602), .A2(n7601), .ZN(n7603) );
  AND2_X1 U9151 ( .A1(n7681), .A2(n7603), .ZN(n7668) );
  NAND2_X1 U9152 ( .A1(n8829), .A2(n7668), .ZN(n7604) );
  OAI211_X1 U9153 ( .C1(n7671), .C2(n8798), .A(n7605), .B(n7604), .ZN(n7606)
         );
  INV_X1 U9154 ( .A(n7606), .ZN(n7607) );
  OAI21_X1 U9155 ( .B1(n10022), .B2(n7670), .A(n7607), .ZN(P2_U3286) );
  XNOR2_X1 U9156 ( .A(n7608), .B(n7610), .ZN(n9664) );
  NAND2_X1 U9157 ( .A1(n7609), .A2(n9900), .ZN(n7611) );
  XNOR2_X1 U9158 ( .A(n7611), .B(n7610), .ZN(n7613) );
  AOI22_X1 U9159 ( .A1(n9709), .A2(n9075), .B1(n9077), .B2(n9710), .ZN(n7612)
         );
  OAI21_X1 U9160 ( .B1(n7613), .B2(n9732), .A(n7612), .ZN(n7614) );
  AOI21_X1 U9161 ( .B1(n9664), .B2(n9735), .A(n7614), .ZN(n9666) );
  AOI21_X1 U9162 ( .B1(n9905), .B2(n9660), .A(n9973), .ZN(n7615) );
  NAND2_X1 U9163 ( .A1(n7615), .A2(n9721), .ZN(n9661) );
  OAI22_X1 U9164 ( .A1(n9930), .A2(n7617), .B1(n7616), .B2(n9925), .ZN(n7618)
         );
  AOI21_X1 U9165 ( .B1(n9739), .B2(n9660), .A(n7618), .ZN(n7619) );
  OAI21_X1 U9166 ( .B1(n9661), .B2(n7620), .A(n7619), .ZN(n7621) );
  AOI21_X1 U9167 ( .B1(n9664), .B2(n9909), .A(n7621), .ZN(n7622) );
  OAI21_X1 U9168 ( .B1(n9666), .B2(n9736), .A(n7622), .ZN(P1_U3281) );
  INV_X1 U9169 ( .A(n8412), .ZN(n7623) );
  AOI211_X1 U9170 ( .C1(n7625), .C2(n7624), .A(n8490), .B(n7623), .ZN(n7631)
         );
  AOI22_X1 U9171 ( .A1(n8465), .A2(n8514), .B1(n7626), .B2(n8500), .ZN(n7629)
         );
  AOI22_X1 U9172 ( .A1(n8479), .A2(n7627), .B1(P2_U3152), .B2(
        P2_REG3_REG_7__SCAN_IN), .ZN(n7628) );
  OAI211_X1 U9173 ( .C1(n8495), .C2(n8137), .A(n7629), .B(n7628), .ZN(n7630)
         );
  OR2_X1 U9174 ( .A1(n7631), .A2(n7630), .ZN(P2_U3215) );
  NOR2_X1 U9175 ( .A1(n7632), .A2(n10022), .ZN(n7638) );
  INV_X1 U9176 ( .A(n7633), .ZN(n7634) );
  AOI22_X1 U9177 ( .A1(n10011), .A2(n7634), .B1(n8478), .B2(n8827), .ZN(n7636)
         );
  NAND2_X1 U9178 ( .A1(n8824), .A2(n8480), .ZN(n7635) );
  OAI211_X1 U9179 ( .C1(n6922), .C2(n10009), .A(n7636), .B(n7635), .ZN(n7637)
         );
  AOI211_X1 U9180 ( .C1(n7639), .C2(n8825), .A(n7638), .B(n7637), .ZN(n7640)
         );
  INV_X1 U9181 ( .A(n7640), .ZN(P2_U3290) );
  NAND2_X1 U9182 ( .A1(n7649), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7642) );
  NAND2_X1 U9183 ( .A1(n7642), .A2(n7641), .ZN(n7646) );
  INV_X1 U9184 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7643) );
  MUX2_X1 U9185 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n7643), .S(n7799), .Z(n7644)
         );
  INV_X1 U9186 ( .A(n7644), .ZN(n7645) );
  NOR2_X1 U9187 ( .A1(n7646), .A2(n7645), .ZN(n7793) );
  AOI21_X1 U9188 ( .B1(n7646), .B2(n7645), .A(n7793), .ZN(n7658) );
  INV_X1 U9189 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7655) );
  INV_X1 U9190 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7647) );
  MUX2_X1 U9191 ( .A(n7647), .B(P2_REG1_REG_11__SCAN_IN), .S(n7799), .Z(n7651)
         );
  AOI21_X1 U9192 ( .B1(n7651), .B2(n7650), .A(n7798), .ZN(n7652) );
  NAND2_X1 U9193 ( .A1(n9991), .A2(n7652), .ZN(n7654) );
  OR2_X1 U9194 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5187), .ZN(n7653) );
  OAI211_X1 U9195 ( .C1(n8602), .C2(n7655), .A(n7654), .B(n7653), .ZN(n7656)
         );
  AOI21_X1 U9196 ( .B1(n7799), .B2(n8596), .A(n7656), .ZN(n7657) );
  OAI21_X1 U9197 ( .B1(n7658), .B2(n9997), .A(n7657), .ZN(P2_U3256) );
  INV_X1 U9198 ( .A(n7659), .ZN(n7667) );
  INV_X1 U9199 ( .A(n8415), .ZN(n8484) );
  AOI22_X1 U9200 ( .A1(n7660), .A2(n8474), .B1(n8484), .B2(n8507), .ZN(n7666)
         );
  INV_X1 U9201 ( .A(n7901), .ZN(n7662) );
  OAI22_X1 U9202 ( .A1(n8494), .A2(n7662), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7661), .ZN(n7664) );
  INV_X1 U9203 ( .A(n8508), .ZN(n8176) );
  OAI22_X1 U9204 ( .A1(n8176), .A2(n8495), .B1(n8496), .B2(n8807), .ZN(n7663)
         );
  AOI211_X1 U9205 ( .C1(n8910), .C2(n8461), .A(n7664), .B(n7663), .ZN(n7665)
         );
  OAI21_X1 U9206 ( .B1(n7667), .B2(n7666), .A(n7665), .ZN(P2_U3243) );
  AOI22_X1 U9207 ( .A1(n7668), .A2(n9683), .B1(n9677), .B2(n7676), .ZN(n7669)
         );
  OAI211_X1 U9208 ( .C1(n7671), .C2(n8914), .A(n7670), .B(n7669), .ZN(n7673)
         );
  NAND2_X1 U9209 ( .A1(n7673), .A2(n10080), .ZN(n7672) );
  OAI21_X1 U9210 ( .B1(n10080), .B2(n7288), .A(n7672), .ZN(P2_U3530) );
  INV_X1 U9211 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n7675) );
  NAND2_X1 U9212 ( .A1(n7673), .A2(n4316), .ZN(n7674) );
  OAI21_X1 U9213 ( .B1(n4316), .B2(n7675), .A(n7674), .ZN(P2_U3481) );
  INV_X1 U9214 ( .A(n8511), .ZN(n8300) );
  OR2_X1 U9215 ( .A1(n7367), .A2(n8300), .ZN(n8163) );
  NAND2_X1 U9216 ( .A1(n7367), .A2(n8300), .ZN(n8161) );
  NAND2_X1 U9217 ( .A1(n8163), .A2(n8161), .ZN(n8267) );
  NAND2_X1 U9218 ( .A1(n7676), .A2(n8512), .ZN(n7720) );
  NAND2_X1 U9219 ( .A1(n7677), .A2(n7720), .ZN(n7678) );
  XOR2_X1 U9220 ( .A(n8267), .B(n7678), .Z(n10069) );
  INV_X1 U9221 ( .A(n10069), .ZN(n7688) );
  XNOR2_X1 U9222 ( .A(n7725), .B(n8267), .ZN(n7680) );
  OAI222_X1 U9223 ( .A1(n8806), .A2(n7756), .B1(n8808), .B2(n8329), .C1(n7680), 
        .C2(n8803), .ZN(n10067) );
  INV_X1 U9224 ( .A(n7681), .ZN(n7682) );
  INV_X1 U9225 ( .A(n7367), .ZN(n10063) );
  OAI21_X1 U9226 ( .B1(n7682), .B2(n10063), .A(n7729), .ZN(n10065) );
  OAI22_X1 U9227 ( .A1(n10009), .A2(n7643), .B1(n7683), .B2(n10025), .ZN(n7684) );
  AOI21_X1 U9228 ( .B1(n8824), .B2(n7367), .A(n7684), .ZN(n7685) );
  OAI21_X1 U9229 ( .B1(n10019), .B2(n10065), .A(n7685), .ZN(n7686) );
  AOI21_X1 U9230 ( .B1(n10067), .B2(n10009), .A(n7686), .ZN(n7687) );
  OAI21_X1 U9231 ( .B1(n7688), .B2(n8798), .A(n7687), .ZN(P2_U3285) );
  INV_X1 U9232 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7689) );
  OAI222_X1 U9233 ( .A1(n8946), .A2(n7690), .B1(P2_U3152), .B2(n8091), .C1(
        n7689), .C2(n8947), .ZN(P2_U3337) );
  XNOR2_X1 U9234 ( .A(n7692), .B(n7691), .ZN(n7697) );
  AND2_X1 U9235 ( .A1(n10130), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9091) );
  NOR2_X1 U9236 ( .A1(n9062), .A2(n9729), .ZN(n7693) );
  AOI211_X1 U9237 ( .C1(n9048), .C2(n9076), .A(n9091), .B(n7693), .ZN(n7694)
         );
  OAI21_X1 U9238 ( .B1(n9050), .B2(n9725), .A(n7694), .ZN(n7695) );
  AOI21_X1 U9239 ( .B1(n9052), .B2(n9759), .A(n7695), .ZN(n7696) );
  OAI21_X1 U9240 ( .B1(n7697), .B2(n9054), .A(n7696), .ZN(P1_U3234) );
  OAI21_X1 U9241 ( .B1(n7699), .B2(n7247), .A(n7698), .ZN(n7710) );
  INV_X1 U9242 ( .A(n7699), .ZN(n7701) );
  NAND3_X1 U9243 ( .A1(n8484), .A2(n7701), .A3(n7700), .ZN(n7703) );
  AOI21_X1 U9244 ( .B1(n7703), .B2(n8495), .A(n7702), .ZN(n7709) );
  AOI22_X1 U9245 ( .A1(n8465), .A2(n8517), .B1(n7704), .B2(n8500), .ZN(n7706)
         );
  OAI211_X1 U9246 ( .C1(n7707), .C2(n8494), .A(n7706), .B(n7705), .ZN(n7708)
         );
  AOI211_X1 U9247 ( .C1(n8474), .C2(n7710), .A(n7709), .B(n7708), .ZN(n7711)
         );
  INV_X1 U9248 ( .A(n7711), .ZN(P2_U3232) );
  INV_X1 U9249 ( .A(n7712), .ZN(n8400) );
  OAI222_X1 U9250 ( .A1(P1_U3084), .A2(n7714), .B1(n9443), .B2(n8400), .C1(
        n7713), .C2(n8318), .ZN(P1_U3331) );
  INV_X1 U9251 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7732) );
  OR2_X1 U9252 ( .A1(n8306), .A2(n7756), .ZN(n8166) );
  NAND2_X1 U9253 ( .A1(n8306), .A2(n7756), .ZN(n8165) );
  NAND2_X1 U9254 ( .A1(n7367), .A2(n8511), .ZN(n7719) );
  INV_X1 U9255 ( .A(n7719), .ZN(n7715) );
  OR2_X1 U9256 ( .A1(n7715), .A2(n8267), .ZN(n7718) );
  AND2_X1 U9257 ( .A1(n8265), .A2(n7718), .ZN(n7716) );
  INV_X1 U9258 ( .A(n7718), .ZN(n7722) );
  AND2_X1 U9259 ( .A1(n7720), .A2(n7719), .ZN(n7721) );
  OR2_X1 U9260 ( .A1(n7722), .A2(n7721), .ZN(n7723) );
  XOR2_X1 U9261 ( .A(n8269), .B(n7750), .Z(n7790) );
  NAND2_X1 U9262 ( .A1(n7725), .A2(n8163), .ZN(n7726) );
  NAND2_X1 U9263 ( .A1(n7726), .A2(n8161), .ZN(n7754) );
  XNOR2_X1 U9264 ( .A(n7754), .B(n8269), .ZN(n7727) );
  AOI222_X1 U9265 ( .A1(n8793), .A2(n7727), .B1(n8509), .B2(n8790), .C1(n8511), 
        .C2(n8788), .ZN(n7785) );
  INV_X1 U9266 ( .A(n4397), .ZN(n7728) );
  AOI21_X1 U9267 ( .B1(n8306), .B2(n7729), .A(n7728), .ZN(n7788) );
  AOI22_X1 U9268 ( .A1(n7788), .A2(n9683), .B1(n9677), .B2(n8306), .ZN(n7730)
         );
  OAI211_X1 U9269 ( .C1(n7790), .C2(n8914), .A(n7785), .B(n7730), .ZN(n7733)
         );
  NAND2_X1 U9270 ( .A1(n7733), .A2(n10080), .ZN(n7731) );
  OAI21_X1 U9271 ( .B1(n10080), .B2(n7732), .A(n7731), .ZN(P2_U3532) );
  INV_X1 U9272 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7735) );
  NAND2_X1 U9273 ( .A1(n7733), .A2(n4316), .ZN(n7734) );
  OAI21_X1 U9274 ( .B1(n4316), .B2(n7735), .A(n7734), .ZN(P2_U3487) );
  INV_X1 U9275 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7749) );
  NOR2_X1 U9276 ( .A1(n7737), .A2(n7736), .ZN(n7739) );
  XNOR2_X1 U9277 ( .A(n9099), .B(n9106), .ZN(n7740) );
  INV_X1 U9278 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7962) );
  NOR2_X1 U9279 ( .A1(n7962), .A2(n7740), .ZN(n9100) );
  AOI211_X1 U9280 ( .C1(n7740), .C2(n7962), .A(n9100), .B(n9872), .ZN(n7741)
         );
  INV_X1 U9281 ( .A(n7741), .ZN(n7748) );
  AND2_X1 U9282 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8044) );
  OAI21_X1 U9283 ( .B1(n7743), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7742), .ZN(
        n9105) );
  XNOR2_X1 U9284 ( .A(n9106), .B(n9105), .ZN(n7744) );
  NOR2_X1 U9285 ( .A1(n5930), .A2(n7744), .ZN(n9107) );
  AOI211_X1 U9286 ( .C1(n7744), .C2(n5930), .A(n9107), .B(n9843), .ZN(n7745)
         );
  AOI211_X1 U9287 ( .C1(n9886), .C2(n7746), .A(n8044), .B(n7745), .ZN(n7747)
         );
  OAI211_X1 U9288 ( .C1(n9899), .C2(n7749), .A(n7748), .B(n7747), .ZN(P1_U3256) );
  OR2_X1 U9289 ( .A1(n7504), .A2(n7751), .ZN(n8174) );
  NAND2_X1 U9290 ( .A1(n7504), .A2(n7751), .ZN(n8173) );
  NAND2_X1 U9291 ( .A1(n7752), .A2(n8270), .ZN(n7753) );
  NAND2_X1 U9292 ( .A1(n7771), .A2(n7753), .ZN(n7761) );
  NAND2_X1 U9293 ( .A1(n7754), .A2(n8166), .ZN(n7755) );
  NAND2_X1 U9294 ( .A1(n7755), .A2(n8165), .ZN(n7772) );
  XNOR2_X1 U9295 ( .A(n7772), .B(n8270), .ZN(n7758) );
  OAI22_X1 U9296 ( .A1(n7756), .A2(n8808), .B1(n8806), .B2(n8176), .ZN(n7757)
         );
  AOI21_X1 U9297 ( .B1(n7758), .B2(n8793), .A(n7757), .ZN(n7759) );
  OAI21_X1 U9298 ( .B1(n7761), .B2(n7760), .A(n7759), .ZN(n9688) );
  INV_X1 U9299 ( .A(n9688), .ZN(n7769) );
  INV_X1 U9300 ( .A(n7761), .ZN(n9690) );
  AND2_X1 U9301 ( .A1(n4397), .A2(n7504), .ZN(n7762) );
  OR2_X1 U9302 ( .A1(n7762), .A2(n7776), .ZN(n9687) );
  AOI22_X1 U9303 ( .A1(n10022), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7763), .B2(
        n8827), .ZN(n7765) );
  NAND2_X1 U9304 ( .A1(n8824), .A2(n7504), .ZN(n7764) );
  OAI211_X1 U9305 ( .C1(n9687), .C2(n10019), .A(n7765), .B(n7764), .ZN(n7766)
         );
  AOI21_X1 U9306 ( .B1(n9690), .B2(n7767), .A(n7766), .ZN(n7768) );
  OAI21_X1 U9307 ( .B1(n7769), .B2(n10022), .A(n7768), .ZN(P2_U3283) );
  NAND2_X1 U9308 ( .A1(n7504), .A2(n8509), .ZN(n7770) );
  XNOR2_X1 U9309 ( .A(n8177), .B(n8508), .ZN(n8271) );
  XNOR2_X1 U9310 ( .A(n7893), .B(n8271), .ZN(n7849) );
  INV_X1 U9311 ( .A(n7849), .ZN(n7782) );
  NAND2_X1 U9312 ( .A1(n7772), .A2(n8270), .ZN(n7773) );
  NAND2_X1 U9313 ( .A1(n7773), .A2(n8173), .ZN(n7906) );
  INV_X1 U9314 ( .A(n8271), .ZN(n7905) );
  XNOR2_X1 U9315 ( .A(n7906), .B(n7905), .ZN(n7775) );
  OAI21_X1 U9316 ( .B1(n7775), .B2(n8803), .A(n7774), .ZN(n7848) );
  INV_X1 U9317 ( .A(n8177), .ZN(n7845) );
  INV_X1 U9318 ( .A(n7899), .ZN(n7900) );
  OAI21_X1 U9319 ( .B1(n7845), .B2(n7776), .A(n7900), .ZN(n7846) );
  AOI22_X1 U9320 ( .A1(n10022), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7777), .B2(
        n8827), .ZN(n7779) );
  NAND2_X1 U9321 ( .A1(n8177), .A2(n8824), .ZN(n7778) );
  OAI211_X1 U9322 ( .C1(n7846), .C2(n10019), .A(n7779), .B(n7778), .ZN(n7780)
         );
  AOI21_X1 U9323 ( .B1(n7848), .B2(n10009), .A(n7780), .ZN(n7781) );
  OAI21_X1 U9324 ( .B1(n7782), .B2(n8798), .A(n7781), .ZN(P2_U3282) );
  INV_X1 U9325 ( .A(n8306), .ZN(n7784) );
  AOI22_X1 U9326 ( .A1(n10022), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n8307), .B2(
        n8827), .ZN(n7783) );
  OAI21_X1 U9327 ( .B1(n7784), .B2(n10018), .A(n7783), .ZN(n7787) );
  NOR2_X1 U9328 ( .A1(n7785), .A2(n10022), .ZN(n7786) );
  AOI211_X1 U9329 ( .C1(n7788), .C2(n8829), .A(n7787), .B(n7786), .ZN(n7789)
         );
  OAI21_X1 U9330 ( .B1(n8798), .B2(n7790), .A(n7789), .ZN(P2_U3284) );
  NAND2_X1 U9331 ( .A1(n8527), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7795) );
  INV_X1 U9332 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7791) );
  MUX2_X1 U9333 ( .A(n7791), .B(P2_REG2_REG_12__SCAN_IN), .S(n8527), .Z(n7792)
         );
  INV_X1 U9334 ( .A(n7792), .ZN(n8524) );
  NOR2_X1 U9335 ( .A1(n7799), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7794) );
  NOR2_X1 U9336 ( .A1(n7794), .A2(n7793), .ZN(n8525) );
  NAND2_X1 U9337 ( .A1(n8524), .A2(n8525), .ZN(n8523) );
  NAND2_X1 U9338 ( .A1(n7795), .A2(n8523), .ZN(n7797) );
  INV_X1 U9339 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7868) );
  AOI22_X1 U9340 ( .A1(n7874), .A2(n7868), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n7869), .ZN(n7796) );
  NOR2_X1 U9341 ( .A1(n7797), .A2(n7796), .ZN(n7867) );
  AOI21_X1 U9342 ( .B1(n7797), .B2(n7796), .A(n7867), .ZN(n7808) );
  INV_X1 U9343 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9691) );
  AOI22_X1 U9344 ( .A1(n7874), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n9691), .B2(
        n7869), .ZN(n7801) );
  AOI21_X1 U9345 ( .B1(n7799), .B2(P2_REG1_REG_11__SCAN_IN), .A(n7798), .ZN(
        n8530) );
  MUX2_X1 U9346 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7732), .S(n8527), .Z(n8529)
         );
  NAND2_X1 U9347 ( .A1(n8530), .A2(n8529), .ZN(n8528) );
  OAI21_X1 U9348 ( .B1(n8527), .B2(P2_REG1_REG_12__SCAN_IN), .A(n8528), .ZN(
        n7800) );
  NAND2_X1 U9349 ( .A1(n7801), .A2(n7800), .ZN(n7873) );
  OAI21_X1 U9350 ( .B1(n7801), .B2(n7800), .A(n7873), .ZN(n7802) );
  NAND2_X1 U9351 ( .A1(n7802), .A2(n9991), .ZN(n7807) );
  INV_X1 U9352 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7804) );
  OAI22_X1 U9353 ( .A1(n8602), .A2(n7804), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7803), .ZN(n7805) );
  AOI21_X1 U9354 ( .B1(n8596), .B2(n7874), .A(n7805), .ZN(n7806) );
  OAI211_X1 U9355 ( .C1(n7808), .C2(n9997), .A(n7807), .B(n7806), .ZN(P2_U3258) );
  AOI21_X1 U9356 ( .B1(n7811), .B2(n7810), .A(n7809), .ZN(n7815) );
  INV_X1 U9357 ( .A(n8789), .ZN(n8349) );
  INV_X1 U9358 ( .A(n8507), .ZN(n8184) );
  OAI22_X1 U9359 ( .A1(n8349), .A2(n8806), .B1(n8808), .B2(n8184), .ZN(n7950)
         );
  AOI22_X1 U9360 ( .A1(n8477), .A2(n7950), .B1(P2_REG3_REG_16__SCAN_IN), .B2(
        P2_U3152), .ZN(n7812) );
  OAI21_X1 U9361 ( .B1(n7944), .B2(n8494), .A(n7812), .ZN(n7813) );
  AOI21_X1 U9362 ( .B1(n8905), .B2(n8500), .A(n7813), .ZN(n7814) );
  OAI21_X1 U9363 ( .B1(n7815), .B2(n8490), .A(n7814), .ZN(P2_U3228) );
  INV_X1 U9364 ( .A(n7816), .ZN(n7820) );
  NAND2_X1 U9365 ( .A1(n9441), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7817) );
  OAI211_X1 U9366 ( .C1(n7820), .C2(n9443), .A(n7818), .B(n7817), .ZN(P1_U3330) );
  NAND2_X1 U9367 ( .A1(n8943), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7819) );
  OAI211_X1 U9368 ( .C1(n7820), .C2(n8946), .A(n8296), .B(n7819), .ZN(P2_U3335) );
  INV_X1 U9369 ( .A(n7821), .ZN(n7822) );
  AOI21_X1 U9370 ( .B1(n7824), .B2(n7823), .A(n7822), .ZN(n7832) );
  INV_X1 U9371 ( .A(n7825), .ZN(n7828) );
  NOR2_X1 U9372 ( .A1(n9060), .A2(n7826), .ZN(n7827) );
  AOI211_X1 U9373 ( .C1(n9024), .C2(n9074), .A(n7828), .B(n7827), .ZN(n7829)
         );
  OAI21_X1 U9374 ( .B1(n9050), .B2(n7855), .A(n7829), .ZN(n7830) );
  AOI21_X1 U9375 ( .B1(n9411), .B2(n9052), .A(n7830), .ZN(n7831) );
  OAI21_X1 U9376 ( .B1(n7832), .B2(n9054), .A(n7831), .ZN(P1_U3222) );
  INV_X1 U9377 ( .A(n7833), .ZN(n7835) );
  NAND2_X1 U9378 ( .A1(n7835), .A2(n7834), .ZN(n7836) );
  XNOR2_X1 U9379 ( .A(n7837), .B(n7836), .ZN(n7844) );
  INV_X1 U9380 ( .A(n7838), .ZN(n7840) );
  NOR2_X1 U9381 ( .A1(n9060), .A2(n9729), .ZN(n7839) );
  AOI211_X1 U9382 ( .C1(n9024), .C2(n9708), .A(n7840), .B(n7839), .ZN(n7841)
         );
  OAI21_X1 U9383 ( .B1(n9050), .B2(n9703), .A(n7841), .ZN(n7842) );
  AOI21_X1 U9384 ( .B1(n9717), .B2(n9052), .A(n7842), .ZN(n7843) );
  OAI21_X1 U9385 ( .B1(n7844), .B2(n9054), .A(n7843), .ZN(P1_U3232) );
  OAI22_X1 U9386 ( .A1(n7846), .A2(n10064), .B1(n7845), .B2(n10062), .ZN(n7847) );
  AOI211_X1 U9387 ( .C1(n7849), .C2(n10068), .A(n7848), .B(n7847), .ZN(n7852)
         );
  NAND2_X1 U9388 ( .A1(n10078), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7850) );
  OAI21_X1 U9389 ( .B1(n7852), .B2(n10078), .A(n7850), .ZN(P2_U3534) );
  NAND2_X1 U9390 ( .A1(n10070), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n7851) );
  OAI21_X1 U9391 ( .B1(n7852), .B2(n10070), .A(n7851), .ZN(P2_U3493) );
  XNOR2_X1 U9392 ( .A(n7853), .B(n7861), .ZN(n9414) );
  INV_X1 U9393 ( .A(n9722), .ZN(n7854) );
  AOI211_X1 U9394 ( .C1(n9411), .C2(n7854), .A(n9973), .B(n9699), .ZN(n9410)
         );
  INV_X1 U9395 ( .A(n7855), .ZN(n7856) );
  AOI22_X1 U9396 ( .A1(n9736), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7856), .B2(
        n9311), .ZN(n7857) );
  OAI21_X1 U9397 ( .B1(n7858), .B2(n9924), .A(n7857), .ZN(n7865) );
  NAND2_X1 U9398 ( .A1(n7860), .A2(n7859), .ZN(n7862) );
  XNOR2_X1 U9399 ( .A(n7862), .B(n7861), .ZN(n7863) );
  AOI222_X1 U9400 ( .A1(n9919), .A2(n7863), .B1(n9074), .B2(n9709), .C1(n9075), 
        .C2(n9710), .ZN(n9413) );
  NOR2_X1 U9401 ( .A1(n9413), .A2(n9736), .ZN(n7864) );
  AOI211_X1 U9402 ( .C1(n9410), .C2(n7987), .A(n7865), .B(n7864), .ZN(n7866)
         );
  OAI21_X1 U9403 ( .B1(n9325), .B2(n9414), .A(n7866), .ZN(P1_U3279) );
  AOI21_X1 U9404 ( .B1(n7869), .B2(n7868), .A(n7867), .ZN(n7872) );
  INV_X1 U9405 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7870) );
  AOI22_X1 U9406 ( .A1(n8003), .A2(n7870), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n7879), .ZN(n7871) );
  NOR2_X1 U9407 ( .A1(n7872), .A2(n7871), .ZN(n7999) );
  AOI21_X1 U9408 ( .B1(n7872), .B2(n7871), .A(n7999), .ZN(n7883) );
  AOI22_X1 U9409 ( .A1(n8003), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n4538), .B2(
        n7879), .ZN(n7876) );
  OAI21_X1 U9410 ( .B1(n7876), .B2(n7875), .A(n8002), .ZN(n7881) );
  NAND2_X1 U9411 ( .A1(n9994), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n7877) );
  OAI211_X1 U9412 ( .C1(n9995), .C2(n7879), .A(n7878), .B(n7877), .ZN(n7880)
         );
  AOI21_X1 U9413 ( .B1(n7881), .B2(n9991), .A(n7880), .ZN(n7882) );
  OAI21_X1 U9414 ( .B1(n7883), .B2(n9997), .A(n7882), .ZN(P2_U3259) );
  OAI211_X1 U9415 ( .C1(n7885), .C2(n7884), .A(n8348), .B(n8474), .ZN(n7889)
         );
  OAI22_X1 U9416 ( .A1(n8494), .A2(n8816), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9604), .ZN(n7887) );
  INV_X1 U9417 ( .A(n8771), .ZN(n8805) );
  OAI22_X1 U9418 ( .A1(n8805), .A2(n8496), .B1(n8495), .B2(n8807), .ZN(n7886)
         );
  AOI211_X1 U9419 ( .C1(n8901), .C2(n8461), .A(n7887), .B(n7886), .ZN(n7888)
         );
  NAND2_X1 U9420 ( .A1(n7889), .A2(n7888), .ZN(P2_U3230) );
  INV_X1 U9421 ( .A(n7890), .ZN(n7913) );
  INV_X1 U9422 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7891) );
  OAI222_X1 U9423 ( .A1(n7892), .A2(P1_U3084), .B1(n9443), .B2(n7913), .C1(
        n7891), .C2(n8318), .ZN(P1_U3329) );
  OR2_X1 U9424 ( .A1(n8177), .A2(n8508), .ZN(n7895) );
  NAND2_X1 U9425 ( .A1(n7896), .A2(n7895), .ZN(n7897) );
  XNOR2_X1 U9426 ( .A(n8910), .B(n8184), .ZN(n8273) );
  NAND2_X1 U9427 ( .A1(n7897), .A2(n8273), .ZN(n7938) );
  OAI21_X1 U9428 ( .B1(n7897), .B2(n8273), .A(n7938), .ZN(n7898) );
  INV_X1 U9429 ( .A(n7898), .ZN(n8915) );
  INV_X1 U9430 ( .A(n8910), .ZN(n7903) );
  AOI21_X1 U9431 ( .B1(n8910), .B2(n7900), .A(n7940), .ZN(n8911) );
  AOI22_X1 U9432 ( .A1(n10022), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n7901), .B2(
        n8827), .ZN(n7902) );
  OAI21_X1 U9433 ( .B1(n7903), .B2(n10018), .A(n7902), .ZN(n7911) );
  OR2_X1 U9434 ( .A1(n8177), .A2(n8176), .ZN(n7904) );
  INV_X1 U9435 ( .A(n8273), .ZN(n8181) );
  NAND2_X1 U9436 ( .A1(n7907), .A2(n8181), .ZN(n7949) );
  OAI211_X1 U9437 ( .C1(n7907), .C2(n8181), .A(n7949), .B(n8793), .ZN(n7909)
         );
  AOI22_X1 U9438 ( .A1(n8788), .A2(n8508), .B1(n8790), .B2(n8506), .ZN(n7908)
         );
  AND2_X1 U9439 ( .A1(n7909), .A2(n7908), .ZN(n8913) );
  NOR2_X1 U9440 ( .A1(n8913), .A2(n10022), .ZN(n7910) );
  AOI211_X1 U9441 ( .C1(n8911), .C2(n8829), .A(n7911), .B(n7910), .ZN(n7912)
         );
  OAI21_X1 U9442 ( .B1(n8915), .B2(n8798), .A(n7912), .ZN(P2_U3281) );
  INV_X1 U9443 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7914) );
  OAI222_X1 U9444 ( .A1(P2_U3152), .A2(n7915), .B1(n8947), .B2(n7914), .C1(
        n8946), .C2(n7913), .ZN(P2_U3334) );
  NAND2_X1 U9445 ( .A1(n7916), .A2(n7917), .ZN(n7918) );
  XOR2_X1 U9446 ( .A(n7920), .B(n7918), .Z(n9409) );
  OAI211_X1 U9447 ( .C1(n7921), .C2(n7920), .A(n7919), .B(n9919), .ZN(n7923)
         );
  AOI22_X1 U9448 ( .A1(n9709), .A2(n9073), .B1(n9074), .B2(n9710), .ZN(n7922)
         );
  NAND2_X1 U9449 ( .A1(n7923), .A2(n7922), .ZN(n9406) );
  INV_X1 U9450 ( .A(n9701), .ZN(n7925) );
  INV_X1 U9451 ( .A(n7960), .ZN(n7924) );
  AOI211_X1 U9452 ( .C1(n9407), .C2(n7925), .A(n9973), .B(n7924), .ZN(n9405)
         );
  NAND2_X1 U9453 ( .A1(n9405), .A2(n7987), .ZN(n7928) );
  INV_X1 U9454 ( .A(n7995), .ZN(n7926) );
  AOI22_X1 U9455 ( .A1(n9736), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7926), .B2(
        n9311), .ZN(n7927) );
  OAI211_X1 U9456 ( .C1(n7929), .C2(n9924), .A(n7928), .B(n7927), .ZN(n7930)
         );
  AOI21_X1 U9457 ( .B1(n9930), .B2(n9406), .A(n7930), .ZN(n7931) );
  OAI21_X1 U9458 ( .B1(n9409), .B2(n9325), .A(n7931), .ZN(P1_U3277) );
  INV_X1 U9459 ( .A(n7932), .ZN(n7935) );
  OAI222_X1 U9460 ( .A1(P1_U3084), .A2(n6196), .B1(n9443), .B2(n7935), .C1(
        n7933), .C2(n8318), .ZN(P1_U3328) );
  OAI222_X1 U9461 ( .A1(n7936), .A2(P2_U3152), .B1(n8946), .B2(n7935), .C1(
        n7934), .C2(n8947), .ZN(P2_U3333) );
  OR2_X1 U9462 ( .A1(n8910), .A2(n8507), .ZN(n7937) );
  NAND2_X1 U9463 ( .A1(n8905), .A2(n8807), .ZN(n8099) );
  OAI21_X1 U9464 ( .B1(n7939), .B2(n8274), .A(n8359), .ZN(n8909) );
  INV_X1 U9465 ( .A(n7940), .ZN(n7942) );
  INV_X1 U9466 ( .A(n8905), .ZN(n7943) );
  NAND2_X1 U9467 ( .A1(n7940), .A2(n7943), .ZN(n8809) );
  INV_X1 U9468 ( .A(n8809), .ZN(n7941) );
  AOI21_X1 U9469 ( .B1(n8905), .B2(n7942), .A(n7941), .ZN(n8906) );
  NOR2_X1 U9470 ( .A1(n7943), .A2(n10018), .ZN(n7947) );
  OAI22_X1 U9471 ( .A1(n10009), .A2(n7945), .B1(n7944), .B2(n10025), .ZN(n7946) );
  AOI211_X1 U9472 ( .C1(n8906), .C2(n8829), .A(n7947), .B(n7946), .ZN(n7953)
         );
  OR2_X1 U9473 ( .A1(n8910), .A2(n8184), .ZN(n7948) );
  XNOR2_X1 U9474 ( .A(n8056), .B(n8274), .ZN(n7951) );
  AOI21_X1 U9475 ( .B1(n7951), .B2(n8793), .A(n7950), .ZN(n8908) );
  OR2_X1 U9476 ( .A1(n8908), .A2(n10022), .ZN(n7952) );
  OAI211_X1 U9477 ( .C1(n8909), .C2(n8798), .A(n7953), .B(n7952), .ZN(P2_U3280) );
  XNOR2_X1 U9478 ( .A(n6277), .B(n7954), .ZN(n9749) );
  INV_X1 U9479 ( .A(n7954), .ZN(n7955) );
  XNOR2_X1 U9480 ( .A(n7956), .B(n7955), .ZN(n7958) );
  AOI22_X1 U9481 ( .A1(n9072), .A2(n9709), .B1(n9710), .B2(n9708), .ZN(n7957)
         );
  OAI21_X1 U9482 ( .B1(n7958), .B2(n9732), .A(n7957), .ZN(n7959) );
  AOI21_X1 U9483 ( .B1(n9749), .B2(n9735), .A(n7959), .ZN(n9751) );
  AOI21_X1 U9484 ( .B1(n7960), .B2(n8048), .A(n9973), .ZN(n7961) );
  NAND2_X1 U9485 ( .A1(n7961), .A2(n7976), .ZN(n9746) );
  OAI22_X1 U9486 ( .A1(n9930), .A2(n7962), .B1(n8046), .B2(n9925), .ZN(n7963)
         );
  AOI21_X1 U9487 ( .B1(n8048), .B2(n9739), .A(n7963), .ZN(n7964) );
  OAI21_X1 U9488 ( .B1(n9746), .B2(n7965), .A(n7964), .ZN(n7966) );
  AOI21_X1 U9489 ( .B1(n9749), .B2(n9909), .A(n7966), .ZN(n7967) );
  OAI21_X1 U9490 ( .B1(n9751), .B2(n9736), .A(n7967), .ZN(P1_U3276) );
  NAND2_X1 U9491 ( .A1(n4395), .A2(n7968), .ZN(n7969) );
  XNOR2_X1 U9492 ( .A(n4391), .B(n7969), .ZN(n7974) );
  INV_X1 U9493 ( .A(n8765), .ZN(n7971) );
  AOI22_X1 U9494 ( .A1(n8464), .A2(n8771), .B1(n8465), .B2(n8772), .ZN(n7970)
         );
  NAND2_X1 U9495 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8600) );
  OAI211_X1 U9496 ( .C1(n8494), .C2(n7971), .A(n7970), .B(n8600), .ZN(n7972)
         );
  AOI21_X1 U9497 ( .B1(n8892), .B2(n8500), .A(n7972), .ZN(n7973) );
  OAI21_X1 U9498 ( .B1(n7974), .B2(n8490), .A(n7973), .ZN(P2_U3221) );
  XNOR2_X1 U9499 ( .A(n7975), .B(n7982), .ZN(n9404) );
  AOI211_X1 U9500 ( .C1(n9401), .C2(n7976), .A(n9973), .B(n8019), .ZN(n9400)
         );
  INV_X1 U9501 ( .A(n9401), .ZN(n7979) );
  INV_X1 U9502 ( .A(n8995), .ZN(n7977) );
  AOI22_X1 U9503 ( .A1(n9736), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n7977), .B2(
        n9311), .ZN(n7978) );
  OAI21_X1 U9504 ( .B1(n7979), .B2(n9924), .A(n7978), .ZN(n7986) );
  NAND2_X1 U9505 ( .A1(n7981), .A2(n7980), .ZN(n7983) );
  XNOR2_X1 U9506 ( .A(n7983), .B(n7982), .ZN(n7984) );
  AOI222_X1 U9507 ( .A1(n9919), .A2(n7984), .B1(n9320), .B2(n9709), .C1(n9073), 
        .C2(n9710), .ZN(n9403) );
  NOR2_X1 U9508 ( .A1(n9403), .A2(n9736), .ZN(n7985) );
  AOI211_X1 U9509 ( .C1(n9400), .C2(n7987), .A(n7986), .B(n7985), .ZN(n7988)
         );
  OAI21_X1 U9510 ( .B1(n9325), .B2(n9404), .A(n7988), .ZN(P1_U3275) );
  NAND2_X1 U9511 ( .A1(n7990), .A2(n7989), .ZN(n7991) );
  XOR2_X1 U9512 ( .A(n7992), .B(n7991), .Z(n7998) );
  AOI22_X1 U9513 ( .A1(n9048), .A2(n9074), .B1(P1_REG3_REG_14__SCAN_IN), .B2(
        P1_U3084), .ZN(n7994) );
  NAND2_X1 U9514 ( .A1(n9024), .A2(n9073), .ZN(n7993) );
  OAI211_X1 U9515 ( .C1(n9050), .C2(n7995), .A(n7994), .B(n7993), .ZN(n7996)
         );
  AOI21_X1 U9516 ( .B1(n9407), .B2(n9052), .A(n7996), .ZN(n7997) );
  OAI21_X1 U9517 ( .B1(n7998), .B2(n9054), .A(n7997), .ZN(P1_U3213) );
  NOR2_X1 U9518 ( .A1(n8003), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8000) );
  NOR2_X1 U9519 ( .A1(n8000), .A2(n7999), .ZN(n8546) );
  XNOR2_X1 U9520 ( .A(n8546), .B(n8547), .ZN(n8001) );
  NOR2_X1 U9521 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n8001), .ZN(n8548) );
  AOI21_X1 U9522 ( .B1(n8001), .B2(P2_REG2_REG_15__SCAN_IN), .A(n8548), .ZN(
        n8012) );
  INV_X1 U9523 ( .A(n8004), .ZN(n8007) );
  INV_X1 U9524 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8005) );
  NOR2_X1 U9525 ( .A1(n8005), .A2(n8004), .ZN(n8538) );
  INV_X1 U9526 ( .A(n8538), .ZN(n8006) );
  OAI211_X1 U9527 ( .C1(n8007), .C2(P2_REG1_REG_15__SCAN_IN), .A(n9991), .B(
        n8006), .ZN(n8011) );
  NOR2_X1 U9528 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7661), .ZN(n8009) );
  NOR2_X1 U9529 ( .A1(n9995), .A2(n8537), .ZN(n8008) );
  AOI211_X1 U9530 ( .C1(P2_ADDR_REG_15__SCAN_IN), .C2(n9994), .A(n8009), .B(
        n8008), .ZN(n8010) );
  OAI211_X1 U9531 ( .C1(n8012), .C2(n9997), .A(n8011), .B(n8010), .ZN(P2_U3260) );
  INV_X1 U9532 ( .A(n8013), .ZN(n8028) );
  OAI222_X1 U9533 ( .A1(n8015), .A2(n10130), .B1(n9443), .B2(n8028), .C1(n8014), .C2(n8318), .ZN(P1_U3327) );
  NAND2_X1 U9534 ( .A1(n8017), .A2(n8016), .ZN(n8018) );
  XOR2_X1 U9535 ( .A(n8022), .B(n8018), .Z(n9399) );
  INV_X1 U9536 ( .A(n8019), .ZN(n8020) );
  AOI21_X1 U9537 ( .B1(n9394), .B2(n8020), .A(n9307), .ZN(n9396) );
  AOI22_X1 U9538 ( .A1(n9736), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9007), .B2(
        n9311), .ZN(n8021) );
  OAI21_X1 U9539 ( .B1(n9010), .B2(n9924), .A(n8021), .ZN(n8026) );
  XNOR2_X1 U9540 ( .A(n8023), .B(n8022), .ZN(n8024) );
  AOI222_X1 U9541 ( .A1(n9919), .A2(n8024), .B1(n9299), .B2(n9709), .C1(n9072), 
        .C2(n9710), .ZN(n9398) );
  NOR2_X1 U9542 ( .A1(n9398), .A2(n9736), .ZN(n8025) );
  AOI211_X1 U9543 ( .C1(n9396), .C2(n9908), .A(n8026), .B(n8025), .ZN(n8027)
         );
  OAI21_X1 U9544 ( .B1(n9399), .B2(n9325), .A(n8027), .ZN(P1_U3274) );
  OAI222_X1 U9545 ( .A1(P2_U3152), .A2(n8030), .B1(n8947), .B2(n8029), .C1(
        n8946), .C2(n8028), .ZN(P2_U3332) );
  XNOR2_X1 U9546 ( .A(n8032), .B(n8031), .ZN(n8037) );
  OAI22_X1 U9547 ( .A1(n8494), .A2(n8754), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8033), .ZN(n8035) );
  INV_X1 U9548 ( .A(n8791), .ZN(n8058) );
  INV_X1 U9549 ( .A(n8749), .ZN(n8059) );
  OAI22_X1 U9550 ( .A1(n8058), .A2(n8495), .B1(n8496), .B2(n8059), .ZN(n8034)
         );
  AOI211_X1 U9551 ( .C1(n8886), .C2(n8461), .A(n8035), .B(n8034), .ZN(n8036)
         );
  OAI21_X1 U9552 ( .B1(n8037), .B2(n8490), .A(n8036), .ZN(P2_U3235) );
  NAND2_X1 U9553 ( .A1(n8039), .A2(n8038), .ZN(n8040) );
  XOR2_X1 U9554 ( .A(n8041), .B(n8040), .Z(n8050) );
  NOR2_X1 U9555 ( .A1(n9060), .A2(n8042), .ZN(n8043) );
  AOI211_X1 U9556 ( .C1(n9024), .C2(n9072), .A(n8044), .B(n8043), .ZN(n8045)
         );
  OAI21_X1 U9557 ( .B1(n9050), .B2(n8046), .A(n8045), .ZN(n8047) );
  AOI21_X1 U9558 ( .B1(n8048), .B2(n9052), .A(n8047), .ZN(n8049) );
  OAI21_X1 U9559 ( .B1(n8050), .B2(n9054), .A(n8049), .ZN(P1_U3239) );
  INV_X1 U9560 ( .A(n8071), .ZN(n8938) );
  INV_X1 U9561 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8052) );
  OAI222_X1 U9562 ( .A1(n9443), .A2(n8938), .B1(n8051), .B2(n10130), .C1(n8052), .C2(n8318), .ZN(P1_U3323) );
  AOI22_X1 U9563 ( .A1(n9441), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        P1_STATE_REG_SCAN_IN), .B2(n9793), .ZN(n8053) );
  OAI21_X1 U9564 ( .B1(n8054), .B2(n9443), .A(n8053), .ZN(P1_U3352) );
  INV_X1 U9565 ( .A(n8191), .ZN(n8055) );
  OR2_X1 U9566 ( .A1(n8901), .A2(n8349), .ZN(n8783) );
  NAND2_X1 U9567 ( .A1(n8901), .A2(n8349), .ZN(n8098) );
  NAND2_X1 U9568 ( .A1(n8783), .A2(n8098), .ZN(n8801) );
  OR2_X1 U9569 ( .A1(n8896), .A2(n8805), .ZN(n8197) );
  NAND2_X1 U9570 ( .A1(n8896), .A2(n8805), .ZN(n8198) );
  NAND2_X1 U9571 ( .A1(n8197), .A2(n8198), .ZN(n8251) );
  INV_X1 U9572 ( .A(n8783), .ZN(n8101) );
  NOR2_X1 U9573 ( .A1(n8251), .A2(n8101), .ZN(n8057) );
  OR2_X1 U9574 ( .A1(n8892), .A2(n8058), .ZN(n8275) );
  NAND2_X1 U9575 ( .A1(n8892), .A2(n8058), .ZN(n8747) );
  INV_X1 U9576 ( .A(n8772), .ZN(n8428) );
  NAND2_X1 U9577 ( .A1(n8886), .A2(n8428), .ZN(n8365) );
  AND2_X1 U9578 ( .A1(n8365), .A2(n8747), .ZN(n8250) );
  NAND2_X1 U9579 ( .A1(n8768), .A2(n8250), .ZN(n8736) );
  OR2_X1 U9580 ( .A1(n8879), .A2(n8059), .ZN(n8093) );
  NAND2_X1 U9581 ( .A1(n8879), .A2(n8059), .ZN(n8095) );
  NAND2_X1 U9582 ( .A1(n8093), .A2(n8095), .ZN(n8737) );
  INV_X1 U9583 ( .A(n8366), .ZN(n8738) );
  NOR2_X1 U9584 ( .A1(n8737), .A2(n8738), .ZN(n8060) );
  NAND2_X1 U9585 ( .A1(n8736), .A2(n8060), .ZN(n8740) );
  OR2_X1 U9586 ( .A1(n8874), .A2(n8427), .ZN(n8094) );
  NAND2_X1 U9587 ( .A1(n8874), .A2(n8427), .ZN(n8096) );
  INV_X1 U9588 ( .A(n8505), .ZN(n8692) );
  OR2_X1 U9589 ( .A1(n8869), .A2(n8692), .ZN(n8210) );
  NAND2_X1 U9590 ( .A1(n8869), .A2(n8692), .ZN(n8690) );
  INV_X1 U9591 ( .A(n8094), .ZN(n8708) );
  NOR2_X1 U9592 ( .A1(n8707), .A2(n8708), .ZN(n8061) );
  INV_X1 U9593 ( .A(n8710), .ZN(n8439) );
  OR2_X1 U9594 ( .A1(n8864), .A2(n8439), .ZN(n8213) );
  NAND2_X1 U9595 ( .A1(n8864), .A2(n8439), .ZN(n8214) );
  INV_X1 U9596 ( .A(n8689), .ZN(n8063) );
  INV_X1 U9597 ( .A(n8690), .ZN(n8062) );
  NOR2_X1 U9598 ( .A1(n8063), .A2(n8062), .ZN(n8064) );
  NAND2_X1 U9599 ( .A1(n8695), .A2(n8213), .ZN(n8672) );
  NAND2_X1 U9600 ( .A1(n8860), .A2(n8693), .ZN(n8219) );
  NAND2_X1 U9601 ( .A1(n8217), .A2(n8219), .ZN(n8671) );
  INV_X1 U9602 ( .A(n8671), .ZN(n8279) );
  OR2_X1 U9603 ( .A1(n8851), .A2(n8440), .ZN(n8225) );
  NAND2_X1 U9604 ( .A1(n8851), .A2(n8440), .ZN(n8220) );
  NAND2_X1 U9605 ( .A1(n8225), .A2(n8220), .ZN(n8645) );
  XNOR2_X1 U9606 ( .A(n8378), .B(n8497), .ZN(n8627) );
  INV_X1 U9607 ( .A(n8627), .ZN(n8630) );
  OR2_X1 U9608 ( .A1(n8378), .A2(n8497), .ZN(n8229) );
  INV_X1 U9609 ( .A(n8632), .ZN(n8234) );
  NAND2_X1 U9610 ( .A1(n8840), .A2(n8234), .ZN(n8227) );
  NAND2_X1 U9611 ( .A1(n8230), .A2(n8227), .ZN(n8619) );
  INV_X1 U9612 ( .A(n8619), .ZN(n8066) );
  NAND2_X1 U9613 ( .A1(n8317), .A2(n4983), .ZN(n8069) );
  NAND2_X1 U9614 ( .A1(n8067), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8068) );
  INV_X1 U9615 ( .A(n8622), .ZN(n8070) );
  OR2_X1 U9616 ( .A1(n8835), .A2(n8070), .ZN(n8236) );
  NAND2_X1 U9617 ( .A1(n8835), .A2(n8070), .ZN(n8237) );
  NAND2_X1 U9618 ( .A1(n8236), .A2(n8237), .ZN(n8376) );
  NAND2_X1 U9619 ( .A1(n8383), .A2(n8377), .ZN(n8382) );
  NOR2_X1 U9620 ( .A1(n8605), .A2(n8091), .ZN(n8080) );
  NAND2_X1 U9621 ( .A1(n8071), .A2(n4983), .ZN(n8074) );
  NAND2_X1 U9622 ( .A1(n8072), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8073) );
  NAND2_X1 U9623 ( .A1(n8074), .A2(n8073), .ZN(n8609) );
  INV_X1 U9624 ( .A(n8237), .ZN(n8075) );
  AOI21_X1 U9625 ( .B1(n8080), .B2(n8609), .A(n8075), .ZN(n8082) );
  NAND2_X1 U9626 ( .A1(n5045), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8079) );
  NAND2_X1 U9627 ( .A1(n5025), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8078) );
  NAND2_X1 U9628 ( .A1(n8076), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8077) );
  NAND3_X1 U9629 ( .A1(n8079), .A2(n8078), .A3(n8077), .ZN(n8503) );
  INV_X1 U9630 ( .A(n8503), .ZN(n8085) );
  NOR2_X1 U9631 ( .A1(n8609), .A2(n8085), .ZN(n8239) );
  INV_X1 U9632 ( .A(n8080), .ZN(n8081) );
  AOI22_X1 U9633 ( .A1(n8382), .A2(n8082), .B1(n8239), .B2(n8081), .ZN(n8087)
         );
  NAND2_X1 U9634 ( .A1(n8933), .A2(n4983), .ZN(n8084) );
  NAND2_X1 U9635 ( .A1(n4315), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8083) );
  INV_X1 U9636 ( .A(n8605), .ZN(n8086) );
  OR2_X1 U9637 ( .A1(n9676), .A2(n8086), .ZN(n8246) );
  NAND2_X1 U9638 ( .A1(n8609), .A2(n8085), .ZN(n8240) );
  NAND2_X1 U9639 ( .A1(n8246), .A2(n8240), .ZN(n8248) );
  NAND2_X1 U9640 ( .A1(n9676), .A2(n8086), .ZN(n8244) );
  OAI21_X1 U9641 ( .B1(n8087), .B2(n8248), .A(n8244), .ZN(n8088) );
  NOR2_X1 U9642 ( .A1(n8091), .A2(n8815), .ZN(n8092) );
  NAND2_X1 U9643 ( .A1(n7024), .A2(n8092), .ZN(n8245) );
  NAND2_X1 U9644 ( .A1(n8094), .A2(n8093), .ZN(n8203) );
  OR2_X1 U9645 ( .A1(n8203), .A2(n8095), .ZN(n8097) );
  NAND2_X1 U9646 ( .A1(n8097), .A2(n8096), .ZN(n8205) );
  INV_X1 U9647 ( .A(n8205), .ZN(n8202) );
  INV_X1 U9648 ( .A(n8203), .ZN(n8200) );
  OAI211_X1 U9649 ( .C1(n8801), .C2(n8099), .A(n8198), .B(n8098), .ZN(n8100)
         );
  MUX2_X1 U9650 ( .A(n8101), .B(n8100), .S(n4583), .Z(n8102) );
  INV_X1 U9651 ( .A(n8102), .ZN(n8196) );
  INV_X1 U9652 ( .A(n8801), .ZN(n8193) );
  AND2_X1 U9653 ( .A1(n8145), .A2(n8143), .ZN(n8103) );
  MUX2_X1 U9654 ( .A(n8160), .B(n8103), .S(n4583), .Z(n8104) );
  AND2_X1 U9655 ( .A1(n8104), .A2(n8152), .ZN(n8155) );
  INV_X1 U9656 ( .A(n8155), .ZN(n8159) );
  INV_X1 U9657 ( .A(n8107), .ZN(n8111) );
  NAND2_X1 U9658 ( .A1(n8109), .A2(n8108), .ZN(n8110) );
  AOI21_X1 U9659 ( .B1(n8127), .B2(n8111), .A(n8110), .ZN(n8117) );
  AND2_X1 U9660 ( .A1(n8119), .A2(n8286), .ZN(n8112) );
  OAI211_X1 U9661 ( .C1(n8113), .C2(n8112), .A(n8123), .B(n8120), .ZN(n8114)
         );
  NAND3_X1 U9662 ( .A1(n8114), .A2(n8122), .A3(n8245), .ZN(n8115) );
  NAND3_X1 U9663 ( .A1(n8127), .A2(n8254), .A3(n8115), .ZN(n8116) );
  OAI21_X1 U9664 ( .B1(n8117), .B2(n4583), .A(n8116), .ZN(n8126) );
  NAND2_X1 U9665 ( .A1(n8118), .A2(n8516), .ZN(n8130) );
  NAND2_X1 U9666 ( .A1(n8120), .A2(n8119), .ZN(n8121) );
  NAND3_X1 U9667 ( .A1(n8122), .A2(n7047), .A3(n8121), .ZN(n8124) );
  NAND3_X1 U9668 ( .A1(n8124), .A2(n4583), .A3(n8123), .ZN(n8125) );
  NAND3_X1 U9669 ( .A1(n8126), .A2(n8130), .A3(n8125), .ZN(n8136) );
  INV_X1 U9670 ( .A(n8127), .ZN(n8133) );
  AND2_X1 U9671 ( .A1(n8129), .A2(n8128), .ZN(n8132) );
  OAI211_X1 U9672 ( .C1(n8133), .C2(n8132), .A(n8131), .B(n8130), .ZN(n8134)
         );
  NAND2_X1 U9673 ( .A1(n8134), .A2(n4583), .ZN(n8135) );
  NAND2_X1 U9674 ( .A1(n8136), .A2(n8135), .ZN(n8140) );
  NAND3_X1 U9675 ( .A1(n8480), .A2(n8137), .A3(n4583), .ZN(n8138) );
  AND2_X1 U9676 ( .A1(n8260), .A2(n8138), .ZN(n8139) );
  NAND2_X1 U9677 ( .A1(n8140), .A2(n8139), .ZN(n8149) );
  NAND3_X1 U9678 ( .A1(n8149), .A2(n8261), .A3(n8141), .ZN(n8144) );
  NAND3_X1 U9679 ( .A1(n8144), .A2(n8143), .A3(n8142), .ZN(n8147) );
  NAND2_X1 U9680 ( .A1(n8163), .A2(n8145), .ZN(n8146) );
  AOI21_X1 U9681 ( .B1(n8155), .B2(n8147), .A(n8146), .ZN(n8157) );
  NAND3_X1 U9682 ( .A1(n8149), .A2(n8261), .A3(n8148), .ZN(n8151) );
  NAND2_X1 U9683 ( .A1(n8151), .A2(n8150), .ZN(n8154) );
  NAND2_X1 U9684 ( .A1(n8161), .A2(n8152), .ZN(n8153) );
  AOI21_X1 U9685 ( .B1(n8155), .B2(n8154), .A(n8153), .ZN(n8156) );
  MUX2_X1 U9686 ( .A(n8157), .B(n8156), .S(n4583), .Z(n8158) );
  OAI211_X1 U9687 ( .C1(n8160), .C2(n8159), .A(n8158), .B(n8269), .ZN(n8172)
         );
  NAND2_X1 U9688 ( .A1(n8165), .A2(n8161), .ZN(n8162) );
  NAND2_X1 U9689 ( .A1(n8162), .A2(n8166), .ZN(n8169) );
  INV_X1 U9690 ( .A(n8163), .ZN(n8164) );
  NAND2_X1 U9691 ( .A1(n8165), .A2(n8164), .ZN(n8167) );
  AND2_X1 U9692 ( .A1(n8167), .A2(n8166), .ZN(n8168) );
  MUX2_X1 U9693 ( .A(n8169), .B(n8168), .S(n4583), .Z(n8171) );
  INV_X1 U9694 ( .A(n8270), .ZN(n8170) );
  AOI21_X1 U9695 ( .B1(n8172), .B2(n8171), .A(n8170), .ZN(n8183) );
  MUX2_X1 U9696 ( .A(n8174), .B(n8173), .S(n8245), .Z(n8175) );
  NAND2_X1 U9697 ( .A1(n8271), .A2(n8175), .ZN(n8182) );
  NAND2_X1 U9698 ( .A1(n8508), .A2(n8245), .ZN(n8179) );
  NAND2_X1 U9699 ( .A1(n8176), .A2(n4583), .ZN(n8178) );
  MUX2_X1 U9700 ( .A(n8179), .B(n8178), .S(n8177), .Z(n8180) );
  OAI211_X1 U9701 ( .C1(n8183), .C2(n8182), .A(n8181), .B(n8180), .ZN(n8188)
         );
  OR2_X1 U9702 ( .A1(n8910), .A2(n8245), .ZN(n8186) );
  NAND2_X1 U9703 ( .A1(n8910), .A2(n8245), .ZN(n8185) );
  MUX2_X1 U9704 ( .A(n8186), .B(n8185), .S(n8184), .Z(n8187) );
  NAND3_X1 U9705 ( .A1(n8189), .A2(n8188), .A3(n8187), .ZN(n8190) );
  OAI21_X1 U9706 ( .B1(n4583), .B2(n8191), .A(n8190), .ZN(n8192) );
  NAND2_X1 U9707 ( .A1(n8193), .A2(n8192), .ZN(n8194) );
  AND2_X1 U9708 ( .A1(n8194), .A2(n8197), .ZN(n8195) );
  NAND2_X1 U9709 ( .A1(n8196), .A2(n8195), .ZN(n8199) );
  NAND3_X1 U9710 ( .A1(n8200), .A2(n8366), .A3(n8204), .ZN(n8201) );
  NAND2_X1 U9711 ( .A1(n8202), .A2(n8201), .ZN(n8208) );
  AOI21_X1 U9712 ( .B1(n8365), .B2(n8204), .A(n8203), .ZN(n8206) );
  NOR2_X1 U9713 ( .A1(n8206), .A2(n8205), .ZN(n8207) );
  MUX2_X1 U9714 ( .A(n8208), .B(n8207), .S(n4583), .Z(n8209) );
  NAND2_X1 U9715 ( .A1(n8689), .A2(n8210), .ZN(n8212) );
  NAND2_X1 U9716 ( .A1(n8214), .A2(n8690), .ZN(n8211) );
  MUX2_X1 U9717 ( .A(n8212), .B(n8211), .S(n8245), .Z(n8216) );
  MUX2_X1 U9718 ( .A(n8214), .B(n8213), .S(n8245), .Z(n8215) );
  NAND2_X1 U9719 ( .A1(n8218), .A2(n8220), .ZN(n8223) );
  NAND2_X1 U9720 ( .A1(n8220), .A2(n8219), .ZN(n8221) );
  NAND2_X1 U9721 ( .A1(n8221), .A2(n8245), .ZN(n8222) );
  NAND2_X1 U9722 ( .A1(n8223), .A2(n8222), .ZN(n8224) );
  OAI211_X1 U9723 ( .C1(n4583), .C2(n8225), .A(n8224), .B(n8630), .ZN(n8232)
         );
  NAND2_X1 U9724 ( .A1(n8378), .A2(n8497), .ZN(n8226) );
  AND2_X1 U9725 ( .A1(n8227), .A2(n8226), .ZN(n8228) );
  MUX2_X1 U9726 ( .A(n8229), .B(n8228), .S(n8245), .Z(n8231) );
  INV_X1 U9727 ( .A(n8840), .ZN(n8618) );
  MUX2_X1 U9728 ( .A(n8632), .B(n8840), .S(n4583), .Z(n8233) );
  OAI21_X1 U9729 ( .B1(n8618), .B2(n8234), .A(n8233), .ZN(n8235) );
  MUX2_X1 U9730 ( .A(n8237), .B(n8236), .S(n8245), .Z(n8238) );
  INV_X1 U9731 ( .A(n8239), .ZN(n8243) );
  NAND2_X1 U9732 ( .A1(n8248), .A2(n4583), .ZN(n8242) );
  NAND2_X1 U9733 ( .A1(n8244), .A2(n8243), .ZN(n8249) );
  INV_X1 U9734 ( .A(n8247), .ZN(n8289) );
  INV_X1 U9735 ( .A(n8248), .ZN(n8283) );
  INV_X1 U9736 ( .A(n8249), .ZN(n8282) );
  INV_X1 U9737 ( .A(n8251), .ZN(n8786) );
  NOR2_X1 U9738 ( .A1(n10013), .A2(n8252), .ZN(n8255) );
  INV_X1 U9739 ( .A(n7027), .ZN(n8253) );
  NAND4_X1 U9740 ( .A1(n8255), .A2(n8254), .A3(n8253), .A4(n7049), .ZN(n8258)
         );
  NOR3_X1 U9741 ( .A1(n8258), .A2(n8257), .A3(n8256), .ZN(n8262) );
  NAND4_X1 U9742 ( .A1(n8262), .A2(n8261), .A3(n8260), .A4(n8259), .ZN(n8264)
         );
  OR3_X1 U9743 ( .A1(n8265), .A2(n8264), .A3(n7531), .ZN(n8266) );
  NOR2_X1 U9744 ( .A1(n8267), .A2(n8266), .ZN(n8268) );
  NAND4_X1 U9745 ( .A1(n8271), .A2(n8270), .A3(n8269), .A4(n8268), .ZN(n8272)
         );
  NOR4_X1 U9746 ( .A1(n8801), .A2(n8274), .A3(n8273), .A4(n8272), .ZN(n8276)
         );
  NAND4_X1 U9747 ( .A1(n8366), .A2(n8786), .A3(n8276), .A4(n8275), .ZN(n8277)
         );
  NOR4_X1 U9748 ( .A1(n8723), .A2(n4563), .A3(n8737), .A4(n8277), .ZN(n8278)
         );
  NAND4_X1 U9749 ( .A1(n8279), .A2(n8689), .A3(n8372), .A4(n8278), .ZN(n8280)
         );
  NOR4_X1 U9750 ( .A1(n8619), .A2(n8627), .A3(n8645), .A4(n8280), .ZN(n8281)
         );
  NAND4_X1 U9751 ( .A1(n8283), .A2(n8282), .A3(n8377), .A4(n8281), .ZN(n8284)
         );
  XNOR2_X1 U9752 ( .A(n8284), .B(n8815), .ZN(n8287) );
  OAI22_X1 U9753 ( .A1(n8287), .A2(n8286), .B1(n5519), .B2(n8285), .ZN(n8288)
         );
  NOR4_X1 U9754 ( .A1(n10027), .A2(n8808), .A3(n8949), .A4(n8293), .ZN(n8295)
         );
  OAI21_X1 U9755 ( .B1(n8296), .B2(n5511), .A(P2_B_REG_SCAN_IN), .ZN(n8294) );
  OAI22_X1 U9756 ( .A1(n8297), .A2(n8296), .B1(n8295), .B2(n8294), .ZN(
        P2_U3244) );
  INV_X1 U9757 ( .A(n8298), .ZN(n8303) );
  INV_X1 U9758 ( .A(n8299), .ZN(n8301) );
  NOR3_X1 U9759 ( .A1(n8301), .A2(n8415), .A3(n8300), .ZN(n8302) );
  AOI21_X1 U9760 ( .B1(n8303), .B2(n8474), .A(n8302), .ZN(n8316) );
  AND2_X1 U9761 ( .A1(n8305), .A2(n8304), .ZN(n8313) );
  AOI22_X1 U9762 ( .A1(n8464), .A2(n8511), .B1(n8465), .B2(n8509), .ZN(n8311)
         );
  NOR2_X1 U9763 ( .A1(n9596), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8526) );
  INV_X1 U9764 ( .A(n8526), .ZN(n8310) );
  NAND2_X1 U9765 ( .A1(n8500), .A2(n8306), .ZN(n8309) );
  NAND2_X1 U9766 ( .A1(n8479), .A2(n8307), .ZN(n8308) );
  NAND4_X1 U9767 ( .A1(n8311), .A2(n8310), .A3(n8309), .A4(n8308), .ZN(n8312)
         );
  AOI21_X1 U9768 ( .B1(n8313), .B2(n8474), .A(n8312), .ZN(n8314) );
  OAI21_X1 U9769 ( .B1(n8316), .B2(n8315), .A(n8314), .ZN(P2_U3226) );
  INV_X1 U9770 ( .A(n8317), .ZN(n8941) );
  INV_X1 U9771 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8319) );
  OAI222_X1 U9772 ( .A1(n9443), .A2(n8941), .B1(n8320), .B2(P1_U3084), .C1(
        n8319), .C2(n8318), .ZN(P1_U3324) );
  NAND3_X1 U9773 ( .A1(n8484), .A2(n8321), .A3(n8514), .ZN(n8322) );
  OAI21_X1 U9774 ( .B1(n8416), .B2(n8490), .A(n8322), .ZN(n8325) );
  INV_X1 U9775 ( .A(n8323), .ZN(n8324) );
  NAND2_X1 U9776 ( .A1(n8325), .A2(n8324), .ZN(n8335) );
  INV_X1 U9777 ( .A(n8326), .ZN(n8327) );
  OAI21_X1 U9778 ( .B1(n8494), .B2(n8328), .A(n8327), .ZN(n8332) );
  OAI22_X1 U9779 ( .A1(n8330), .A2(n8495), .B1(n8496), .B2(n8329), .ZN(n8331)
         );
  AOI211_X1 U9780 ( .C1(n8333), .C2(n8500), .A(n8332), .B(n8331), .ZN(n8334)
         );
  OAI211_X1 U9781 ( .C1(n8490), .C2(n8336), .A(n8335), .B(n8334), .ZN(P2_U3233) );
  INV_X1 U9782 ( .A(n8337), .ZN(n8344) );
  NAND2_X1 U9783 ( .A1(n8338), .A2(n9908), .ZN(n8341) );
  AOI22_X1 U9784 ( .A1(n8339), .A2(n9311), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9736), .ZN(n8340) );
  OAI211_X1 U9785 ( .C1(n8342), .C2(n9924), .A(n8341), .B(n8340), .ZN(n8343)
         );
  AOI21_X1 U9786 ( .B1(n8344), .B2(n9930), .A(n8343), .ZN(n8345) );
  OAI21_X1 U9787 ( .B1(n8346), .B2(n9325), .A(n8345), .ZN(P1_U3355) );
  AOI21_X1 U9788 ( .B1(n8348), .B2(n8347), .A(n8490), .ZN(n8352) );
  NOR3_X1 U9789 ( .A1(n8350), .A2(n8349), .A3(n8415), .ZN(n8351) );
  NOR2_X1 U9790 ( .A1(n8352), .A2(n8351), .ZN(n8357) );
  AOI22_X1 U9791 ( .A1(n8464), .A2(n8789), .B1(n8465), .B2(n8791), .ZN(n8353)
         );
  NAND2_X1 U9792 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8580) );
  OAI211_X1 U9793 ( .C1(n8494), .C2(n8794), .A(n8353), .B(n8580), .ZN(n8354)
         );
  AOI21_X1 U9794 ( .B1(n8896), .B2(n8500), .A(n8354), .ZN(n8355) );
  OAI21_X1 U9795 ( .B1(n8357), .B2(n8356), .A(n8355), .ZN(P2_U3240) );
  NAND2_X1 U9796 ( .A1(n8905), .A2(n8506), .ZN(n8358) );
  OR2_X1 U9797 ( .A1(n8901), .A2(n8789), .ZN(n8360) );
  NAND2_X1 U9798 ( .A1(n8896), .A2(n8771), .ZN(n8361) );
  NAND2_X1 U9799 ( .A1(n8892), .A2(n8791), .ZN(n8362) );
  NAND2_X1 U9800 ( .A1(n8761), .A2(n8362), .ZN(n8364) );
  OR2_X1 U9801 ( .A1(n8892), .A2(n8791), .ZN(n8363) );
  OR2_X1 U9802 ( .A1(n8751), .A2(n4829), .ZN(n8367) );
  NAND2_X1 U9803 ( .A1(n8886), .A2(n8772), .ZN(n8730) );
  NAND2_X1 U9804 ( .A1(n8879), .A2(n8749), .ZN(n8368) );
  AND2_X1 U9805 ( .A1(n8730), .A2(n8368), .ZN(n8369) );
  OR2_X1 U9806 ( .A1(n4829), .A2(n8369), .ZN(n8370) );
  INV_X1 U9807 ( .A(n8427), .ZN(n8742) );
  OR2_X1 U9808 ( .A1(n8864), .A2(n8710), .ZN(n8373) );
  NAND2_X1 U9809 ( .A1(n8678), .A2(n8373), .ZN(n8664) );
  INV_X1 U9810 ( .A(n8693), .ZN(n8504) );
  OR2_X1 U9811 ( .A1(n8860), .A2(n8504), .ZN(n8374) );
  NAND2_X1 U9812 ( .A1(n8628), .A2(n8627), .ZN(n8626) );
  INV_X1 U9813 ( .A(n8864), .ZN(n8687) );
  INV_X1 U9814 ( .A(n8874), .ZN(n8720) );
  INV_X1 U9815 ( .A(n8892), .ZN(n8767) );
  NAND2_X1 U9816 ( .A1(n8687), .A2(n8701), .ZN(n8681) );
  NOR2_X4 U9817 ( .A1(n8851), .A2(n8666), .ZN(n8655) );
  AOI21_X1 U9818 ( .B1(n8835), .B2(n8614), .A(n8610), .ZN(n8836) );
  INV_X1 U9819 ( .A(n8379), .ZN(n8380) );
  AOI22_X1 U9820 ( .A1(n10022), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8380), .B2(
        n8827), .ZN(n8381) );
  OAI21_X1 U9821 ( .B1(n4560), .B2(n10018), .A(n8381), .ZN(n8390) );
  OAI21_X1 U9822 ( .B1(n8377), .B2(n8383), .A(n8382), .ZN(n8389) );
  OR2_X1 U9823 ( .A1(n8949), .A2(n8384), .ZN(n8385) );
  AND2_X1 U9824 ( .A1(n8790), .A2(n8385), .ZN(n8606) );
  NAND2_X1 U9825 ( .A1(n8606), .A2(n8503), .ZN(n8386) );
  INV_X1 U9826 ( .A(n8718), .ZN(n8394) );
  NAND2_X1 U9827 ( .A1(n8505), .A2(n8790), .ZN(n8392) );
  NAND2_X1 U9828 ( .A1(n8749), .A2(n8788), .ZN(n8391) );
  NAND2_X1 U9829 ( .A1(n8392), .A2(n8391), .ZN(n8724) );
  AOI22_X1 U9830 ( .A1(n8477), .A2(n8724), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3152), .ZN(n8393) );
  OAI21_X1 U9831 ( .B1(n8394), .B2(n8494), .A(n8393), .ZN(n8397) );
  NOR3_X1 U9832 ( .A1(n8395), .A2(n8427), .A3(n8415), .ZN(n8396) );
  AOI211_X1 U9833 ( .C1(n8874), .C2(n8500), .A(n8397), .B(n8396), .ZN(n8398)
         );
  OAI21_X1 U9834 ( .B1(n8399), .B2(n8490), .A(n8398), .ZN(P2_U3237) );
  OAI222_X1 U9835 ( .A1(n8947), .A2(n8401), .B1(n8946), .B2(n8400), .C1(n7024), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  NAND2_X1 U9836 ( .A1(n8474), .A2(n8402), .ZN(n8405) );
  NAND2_X1 U9837 ( .A1(n8484), .A2(n8505), .ZN(n8404) );
  MUX2_X1 U9838 ( .A(n8405), .B(n8404), .S(n8403), .Z(n8409) );
  OAI22_X1 U9839 ( .A1(n8494), .A2(n8702), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9561), .ZN(n8407) );
  OAI22_X1 U9840 ( .A1(n8439), .A2(n8496), .B1(n8495), .B2(n8427), .ZN(n8406)
         );
  AOI211_X1 U9841 ( .C1(n8869), .C2(n8461), .A(n8407), .B(n8406), .ZN(n8408)
         );
  NAND2_X1 U9842 ( .A1(n8409), .A2(n8408), .ZN(P2_U3218) );
  INV_X1 U9843 ( .A(n8410), .ZN(n8411) );
  AOI21_X1 U9844 ( .B1(n8412), .B2(n8411), .A(n8490), .ZN(n8418) );
  NOR3_X1 U9845 ( .A1(n8415), .A2(n8414), .A3(n8413), .ZN(n8417) );
  OAI21_X1 U9846 ( .B1(n8418), .B2(n8417), .A(n8416), .ZN(n8424) );
  AOI22_X1 U9847 ( .A1(n8465), .A2(n8513), .B1(n8419), .B2(n8500), .ZN(n8423)
         );
  AOI22_X1 U9848 ( .A1(n8479), .A2(n8420), .B1(P2_REG3_REG_8__SCAN_IN), .B2(
        P2_U3152), .ZN(n8422) );
  NAND2_X1 U9849 ( .A1(n8464), .A2(n8515), .ZN(n8421) );
  NAND4_X1 U9850 ( .A1(n8424), .A2(n8423), .A3(n8422), .A4(n8421), .ZN(
        P2_U3223) );
  XNOR2_X1 U9851 ( .A(n8426), .B(n8425), .ZN(n8432) );
  OAI22_X1 U9852 ( .A1(n8494), .A2(n8733), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9564), .ZN(n8430) );
  OAI22_X1 U9853 ( .A1(n8428), .A2(n8495), .B1(n8496), .B2(n8427), .ZN(n8429)
         );
  AOI211_X1 U9854 ( .C1(n8879), .C2(n8461), .A(n8430), .B(n8429), .ZN(n8431)
         );
  OAI21_X1 U9855 ( .B1(n8432), .B2(n8490), .A(n8431), .ZN(P2_U3225) );
  XOR2_X1 U9856 ( .A(n8435), .B(n8434), .Z(n8436) );
  XNOR2_X1 U9857 ( .A(n8433), .B(n8436), .ZN(n8444) );
  INV_X1 U9858 ( .A(n8668), .ZN(n8438) );
  OAI22_X1 U9859 ( .A1(n8494), .A2(n8438), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8437), .ZN(n8442) );
  OAI22_X1 U9860 ( .A1(n8440), .A2(n8496), .B1(n8495), .B2(n8439), .ZN(n8441)
         );
  AOI211_X1 U9861 ( .C1(n8860), .C2(n8461), .A(n8442), .B(n8441), .ZN(n8443)
         );
  OAI21_X1 U9862 ( .B1(n8444), .B2(n8490), .A(n8443), .ZN(P2_U3227) );
  AOI21_X1 U9863 ( .B1(n8446), .B2(n8445), .A(n8490), .ZN(n8448) );
  NAND2_X1 U9864 ( .A1(n8448), .A2(n8447), .ZN(n8454) );
  AOI22_X1 U9865 ( .A1(n8477), .A2(n8449), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n8453) );
  AOI22_X1 U9866 ( .A1(n8500), .A2(n8451), .B1(n8479), .B2(n8450), .ZN(n8452)
         );
  NAND3_X1 U9867 ( .A1(n8454), .A2(n8453), .A3(n8452), .ZN(P2_U3229) );
  NAND2_X1 U9868 ( .A1(n8474), .A2(n8455), .ZN(n8458) );
  NAND2_X1 U9869 ( .A1(n8484), .A2(n8710), .ZN(n8457) );
  MUX2_X1 U9870 ( .A(n8458), .B(n8457), .S(n8456), .Z(n8463) );
  OAI22_X1 U9871 ( .A1(n8494), .A2(n8684), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9565), .ZN(n8460) );
  OAI22_X1 U9872 ( .A1(n8692), .A2(n8495), .B1(n8496), .B2(n8693), .ZN(n8459)
         );
  AOI211_X1 U9873 ( .C1(n8864), .C2(n8461), .A(n8460), .B(n8459), .ZN(n8462)
         );
  NAND2_X1 U9874 ( .A1(n8463), .A2(n8462), .ZN(P2_U3231) );
  AOI22_X1 U9875 ( .A1(n8465), .A2(n8519), .B1(n8464), .B2(n7025), .ZN(n8472)
         );
  AOI22_X1 U9876 ( .A1(n8500), .A2(n8823), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n8466), .ZN(n8471) );
  AOI21_X1 U9877 ( .B1(n8467), .B2(n8468), .A(n8490), .ZN(n8469) );
  NAND2_X1 U9878 ( .A1(n8469), .A2(n7244), .ZN(n8470) );
  NAND3_X1 U9879 ( .A1(n8472), .A2(n8471), .A3(n8470), .ZN(P2_U3239) );
  OAI21_X1 U9880 ( .B1(n8481), .B2(n8447), .A(n8473), .ZN(n8475) );
  NAND2_X1 U9881 ( .A1(n8475), .A2(n8474), .ZN(n8488) );
  AOI22_X1 U9882 ( .A1(n8477), .A2(n8476), .B1(P2_REG3_REG_6__SCAN_IN), .B2(
        P2_U3152), .ZN(n8487) );
  AOI22_X1 U9883 ( .A1(n8500), .A2(n8480), .B1(n8479), .B2(n8478), .ZN(n8486)
         );
  INV_X1 U9884 ( .A(n8481), .ZN(n8483) );
  NAND4_X1 U9885 ( .A1(n8484), .A2(n8483), .A3(n8482), .A4(n8517), .ZN(n8485)
         );
  NAND4_X1 U9886 ( .A1(n8488), .A2(n8487), .A3(n8486), .A4(n8485), .ZN(
        P2_U3241) );
  AOI21_X1 U9887 ( .B1(n8489), .B2(n8491), .A(n8490), .ZN(n8493) );
  NAND2_X1 U9888 ( .A1(n8493), .A2(n8492), .ZN(n8502) );
  OAI22_X1 U9889 ( .A1(n8494), .A2(n8656), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9539), .ZN(n8499) );
  OAI22_X1 U9890 ( .A1(n8497), .A2(n8496), .B1(n8693), .B2(n8495), .ZN(n8498)
         );
  AOI211_X1 U9891 ( .C1(n8851), .C2(n8500), .A(n8499), .B(n8498), .ZN(n8501)
         );
  NAND2_X1 U9892 ( .A1(n8502), .A2(n8501), .ZN(P2_U3242) );
  MUX2_X1 U9893 ( .A(n8503), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8521), .Z(
        P2_U3582) );
  MUX2_X1 U9894 ( .A(n8622), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8521), .Z(
        P2_U3581) );
  MUX2_X1 U9895 ( .A(n8632), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8521), .Z(
        P2_U3580) );
  MUX2_X1 U9896 ( .A(n8649), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8521), .Z(
        P2_U3579) );
  MUX2_X1 U9897 ( .A(n8673), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8521), .Z(
        P2_U3578) );
  MUX2_X1 U9898 ( .A(n8504), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8521), .Z(
        P2_U3577) );
  MUX2_X1 U9899 ( .A(n8710), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8521), .Z(
        P2_U3576) );
  MUX2_X1 U9900 ( .A(n8505), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8521), .Z(
        P2_U3575) );
  MUX2_X1 U9901 ( .A(n8742), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8521), .Z(
        P2_U3574) );
  MUX2_X1 U9902 ( .A(n8749), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8521), .Z(
        P2_U3573) );
  MUX2_X1 U9903 ( .A(n8772), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8521), .Z(
        P2_U3572) );
  MUX2_X1 U9904 ( .A(n8791), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8521), .Z(
        P2_U3571) );
  MUX2_X1 U9905 ( .A(n8771), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8521), .Z(
        P2_U3570) );
  MUX2_X1 U9906 ( .A(n8789), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8521), .Z(
        P2_U3569) );
  MUX2_X1 U9907 ( .A(n8506), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8521), .Z(
        P2_U3568) );
  MUX2_X1 U9908 ( .A(n8507), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8521), .Z(
        P2_U3567) );
  MUX2_X1 U9909 ( .A(n8508), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8521), .Z(
        P2_U3566) );
  MUX2_X1 U9910 ( .A(n8509), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8521), .Z(
        P2_U3565) );
  MUX2_X1 U9911 ( .A(n8510), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8521), .Z(
        P2_U3564) );
  MUX2_X1 U9912 ( .A(n8511), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8521), .Z(
        P2_U3563) );
  MUX2_X1 U9913 ( .A(n8512), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8521), .Z(
        P2_U3562) );
  MUX2_X1 U9914 ( .A(n8513), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8521), .Z(
        P2_U3561) );
  MUX2_X1 U9915 ( .A(n8514), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8521), .Z(
        P2_U3560) );
  MUX2_X1 U9916 ( .A(n8515), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8521), .Z(
        P2_U3559) );
  MUX2_X1 U9917 ( .A(n8516), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8521), .Z(
        P2_U3558) );
  MUX2_X1 U9918 ( .A(n8517), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8521), .Z(
        P2_U3557) );
  MUX2_X1 U9919 ( .A(n8518), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8521), .Z(
        P2_U3556) );
  MUX2_X1 U9920 ( .A(n8519), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8521), .Z(
        P2_U3555) );
  MUX2_X1 U9921 ( .A(n8520), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8521), .Z(
        P2_U3554) );
  MUX2_X1 U9922 ( .A(n7025), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8521), .Z(
        P2_U3553) );
  MUX2_X1 U9923 ( .A(n8522), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8521), .Z(
        P2_U3552) );
  OAI211_X1 U9924 ( .C1(n8525), .C2(n8524), .A(n9992), .B(n8523), .ZN(n8535)
         );
  AOI21_X1 U9925 ( .B1(n9994), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n8526), .ZN(
        n8534) );
  NAND2_X1 U9926 ( .A1(n8596), .A2(n8527), .ZN(n8533) );
  OAI21_X1 U9927 ( .B1(n8530), .B2(n8529), .A(n8528), .ZN(n8531) );
  NAND2_X1 U9928 ( .A1(n9991), .A2(n8531), .ZN(n8532) );
  NAND4_X1 U9929 ( .A1(n8535), .A2(n8534), .A3(n8533), .A4(n8532), .ZN(
        P2_U3257) );
  NOR2_X1 U9930 ( .A1(n8537), .A2(n8536), .ZN(n8539) );
  NOR2_X1 U9931 ( .A1(n8539), .A2(n8538), .ZN(n8542) );
  OR2_X1 U9932 ( .A1(n8553), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8564) );
  NAND2_X1 U9933 ( .A1(n8553), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8540) );
  AND2_X1 U9934 ( .A1(n8564), .A2(n8540), .ZN(n8541) );
  NAND2_X1 U9935 ( .A1(n8541), .A2(n8542), .ZN(n8563) );
  OAI21_X1 U9936 ( .B1(n8542), .B2(n8541), .A(n8563), .ZN(n8543) );
  NAND2_X1 U9937 ( .A1(n8543), .A2(n9991), .ZN(n8557) );
  NOR2_X1 U9938 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8544), .ZN(n8545) );
  AOI21_X1 U9939 ( .B1(n9994), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8545), .ZN(
        n8556) );
  NOR2_X1 U9940 ( .A1(n8547), .A2(n8546), .ZN(n8549) );
  NOR2_X1 U9941 ( .A1(n8549), .A2(n8548), .ZN(n8552) );
  OR2_X1 U9942 ( .A1(n8553), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8550) );
  NAND2_X1 U9943 ( .A1(n8553), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8559) );
  AND2_X1 U9944 ( .A1(n8550), .A2(n8559), .ZN(n8551) );
  NAND2_X1 U9945 ( .A1(n8551), .A2(n8552), .ZN(n8558) );
  OAI211_X1 U9946 ( .C1(n8552), .C2(n8551), .A(n9992), .B(n8558), .ZN(n8555)
         );
  NAND2_X1 U9947 ( .A1(n8596), .A2(n8553), .ZN(n8554) );
  NAND4_X1 U9948 ( .A1(n8557), .A2(n8556), .A3(n8555), .A4(n8554), .ZN(
        P2_U3261) );
  NAND2_X1 U9949 ( .A1(n8559), .A2(n8558), .ZN(n8561) );
  INV_X1 U9950 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8817) );
  XNOR2_X1 U9951 ( .A(n8578), .B(n8817), .ZN(n8560) );
  NAND2_X1 U9952 ( .A1(n8560), .A2(n8561), .ZN(n8572) );
  OAI211_X1 U9953 ( .C1(n8561), .C2(n8560), .A(n9992), .B(n8572), .ZN(n8571)
         );
  NOR2_X1 U9954 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9604), .ZN(n8562) );
  AOI21_X1 U9955 ( .B1(n9994), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8562), .ZN(
        n8570) );
  NAND2_X1 U9956 ( .A1(n8596), .A2(n8578), .ZN(n8569) );
  XNOR2_X1 U9957 ( .A(n8578), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8566) );
  AOI21_X1 U9958 ( .B1(n8566), .B2(n8565), .A(n8577), .ZN(n8567) );
  NAND2_X1 U9959 ( .A1(n9991), .A2(n8567), .ZN(n8568) );
  NAND4_X1 U9960 ( .A1(n8571), .A2(n8570), .A3(n8569), .A4(n8568), .ZN(
        P2_U3262) );
  INV_X1 U9961 ( .A(n8572), .ZN(n8573) );
  AOI21_X1 U9962 ( .B1(n8578), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8573), .ZN(
        n8575) );
  AND2_X1 U9963 ( .A1(n8575), .A2(n8589), .ZN(n8587) );
  INV_X1 U9964 ( .A(n8587), .ZN(n8574) );
  OAI21_X1 U9965 ( .B1(n8575), .B2(n8589), .A(n8574), .ZN(n8576) );
  NOR2_X1 U9966 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8576), .ZN(n8586) );
  AOI21_X1 U9967 ( .B1(n8576), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8586), .ZN(
        n8585) );
  XOR2_X1 U9968 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8583), .Z(n8591) );
  XOR2_X1 U9969 ( .A(n8590), .B(n8591), .Z(n8581) );
  NAND2_X1 U9970 ( .A1(n9994), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n8579) );
  OAI211_X1 U9971 ( .C1(n9996), .C2(n8581), .A(n8580), .B(n8579), .ZN(n8582)
         );
  AOI21_X1 U9972 ( .B1(n8583), .B2(n8596), .A(n8582), .ZN(n8584) );
  OAI21_X1 U9973 ( .B1(n8585), .B2(n9997), .A(n8584), .ZN(P2_U3263) );
  INV_X1 U9974 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8603) );
  NOR2_X1 U9975 ( .A1(n8587), .A2(n8586), .ZN(n8588) );
  XOR2_X1 U9976 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8588), .Z(n8594) );
  XNOR2_X1 U9977 ( .A(n8592), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8597) );
  INV_X1 U9978 ( .A(n8597), .ZN(n8593) );
  AOI22_X1 U9979 ( .A1(n8594), .A2(n9992), .B1(n8593), .B2(n9991), .ZN(n8599)
         );
  NOR2_X1 U9980 ( .A1(n8594), .A2(n9997), .ZN(n8595) );
  AOI211_X1 U9981 ( .C1(n9991), .C2(n8597), .A(n8596), .B(n8595), .ZN(n8598)
         );
  MUX2_X1 U9982 ( .A(n8599), .B(n8598), .S(n8657), .Z(n8601) );
  OAI211_X1 U9983 ( .C1(n8603), .C2(n8602), .A(n8601), .B(n8600), .ZN(P2_U3264) );
  INV_X1 U9984 ( .A(n8609), .ZN(n9680) );
  AND2_X1 U9985 ( .A1(n8606), .A2(n8605), .ZN(n9675) );
  INV_X1 U9986 ( .A(n9675), .ZN(n9679) );
  NOR2_X1 U9987 ( .A1(n10022), .A2(n9679), .ZN(n8611) );
  AOI21_X1 U9988 ( .B1(n10022), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8611), .ZN(
        n8608) );
  NAND2_X1 U9989 ( .A1(n9676), .A2(n8824), .ZN(n8607) );
  OAI211_X1 U9990 ( .C1(n9673), .C2(n10019), .A(n8608), .B(n8607), .ZN(
        P2_U3265) );
  XNOR2_X1 U9991 ( .A(n8610), .B(n8609), .ZN(n9682) );
  NAND2_X1 U9992 ( .A1(n9682), .A2(n8829), .ZN(n8613) );
  AOI21_X1 U9993 ( .B1(n10022), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8611), .ZN(
        n8612) );
  OAI211_X1 U9994 ( .C1(n9680), .C2(n10018), .A(n8613), .B(n8612), .ZN(
        P2_U3266) );
  INV_X1 U9995 ( .A(n8614), .ZN(n8615) );
  AOI21_X1 U9996 ( .B1(n8840), .B2(n8635), .A(n8615), .ZN(n8841) );
  AOI22_X1 U9997 ( .A1(n8616), .A2(n8827), .B1(n10022), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n8617) );
  OAI21_X1 U9998 ( .B1(n8618), .B2(n10018), .A(n8617), .ZN(n8625) );
  XNOR2_X1 U9999 ( .A(n8620), .B(n8619), .ZN(n8621) );
  OAI21_X1 U10000 ( .B1(n8628), .B2(n8627), .A(n8626), .ZN(n8849) );
  INV_X1 U10001 ( .A(n8849), .ZN(n8641) );
  OAI211_X1 U10002 ( .C1(n8631), .C2(n8630), .A(n8629), .B(n8793), .ZN(n8634)
         );
  AOI22_X1 U10003 ( .A1(n8632), .A2(n8790), .B1(n8788), .B2(n8673), .ZN(n8633)
         );
  NAND2_X1 U10004 ( .A1(n8634), .A2(n8633), .ZN(n8848) );
  OAI21_X1 U10005 ( .B1(n8845), .B2(n8655), .A(n8635), .ZN(n8846) );
  NOR2_X1 U10006 ( .A1(n8846), .A2(n10019), .ZN(n8639) );
  AOI22_X1 U10007 ( .A1(P2_REG2_REG_27__SCAN_IN), .A2(n10022), .B1(n8636), 
        .B2(n8827), .ZN(n8637) );
  OAI21_X1 U10008 ( .B1(n8845), .B2(n10018), .A(n8637), .ZN(n8638) );
  AOI211_X1 U10009 ( .C1(n8848), .C2(n10009), .A(n8639), .B(n8638), .ZN(n8640)
         );
  OAI21_X1 U10010 ( .B1(n8641), .B2(n8798), .A(n8640), .ZN(P2_U3269) );
  OR2_X1 U10011 ( .A1(n8642), .A2(n8645), .ZN(n8643) );
  NAND2_X1 U10012 ( .A1(n8644), .A2(n8643), .ZN(n8856) );
  INV_X1 U10013 ( .A(n8856), .ZN(n8662) );
  AOI22_X1 U10014 ( .A1(n8851), .A2(n8824), .B1(n10022), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8661) );
  NAND2_X1 U10015 ( .A1(n8646), .A2(n8645), .ZN(n8647) );
  NAND2_X1 U10016 ( .A1(n8648), .A2(n8647), .ZN(n8652) );
  NAND2_X1 U10017 ( .A1(n8649), .A2(n8790), .ZN(n8650) );
  OAI21_X1 U10018 ( .B1(n8693), .B2(n8808), .A(n8650), .ZN(n8651) );
  AOI21_X1 U10019 ( .B1(n8652), .B2(n8793), .A(n8651), .ZN(n8854) );
  INV_X1 U10020 ( .A(n8854), .ZN(n8659) );
  NAND2_X1 U10021 ( .A1(n8851), .A2(n8666), .ZN(n8653) );
  NAND2_X1 U10022 ( .A1(n8653), .A2(n9683), .ZN(n8654) );
  OR2_X1 U10023 ( .A1(n8655), .A2(n8654), .ZN(n8852) );
  OAI22_X1 U10024 ( .A1(n8852), .A2(n8657), .B1(n10025), .B2(n8656), .ZN(n8658) );
  OAI21_X1 U10025 ( .B1(n8659), .B2(n8658), .A(n10009), .ZN(n8660) );
  OAI211_X1 U10026 ( .C1(n8662), .C2(n8798), .A(n8661), .B(n8660), .ZN(
        P2_U3270) );
  OAI21_X1 U10027 ( .B1(n8664), .B2(n8671), .A(n8663), .ZN(n8665) );
  INV_X1 U10028 ( .A(n8665), .ZN(n8863) );
  INV_X1 U10029 ( .A(n8666), .ZN(n8667) );
  AOI211_X1 U10030 ( .C1(n8860), .C2(n8681), .A(n10064), .B(n8667), .ZN(n8859)
         );
  INV_X1 U10031 ( .A(n8860), .ZN(n8670) );
  AOI22_X1 U10032 ( .A1(n10022), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8668), 
        .B2(n8827), .ZN(n8669) );
  OAI21_X1 U10033 ( .B1(n8670), .B2(n10018), .A(n8669), .ZN(n8676) );
  XNOR2_X1 U10034 ( .A(n8672), .B(n8671), .ZN(n8674) );
  AOI222_X1 U10035 ( .A1(n8793), .A2(n8674), .B1(n8673), .B2(n8790), .C1(n8710), .C2(n8788), .ZN(n8862) );
  NOR2_X1 U10036 ( .A1(n8862), .A2(n10022), .ZN(n8675) );
  AOI211_X1 U10037 ( .C1(n8859), .C2(n10011), .A(n8676), .B(n8675), .ZN(n8677)
         );
  OAI21_X1 U10038 ( .B1(n8863), .B2(n8798), .A(n8677), .ZN(P2_U3271) );
  INV_X1 U10039 ( .A(n8678), .ZN(n8679) );
  AOI21_X1 U10040 ( .B1(n8689), .B2(n8680), .A(n8679), .ZN(n8868) );
  INV_X1 U10041 ( .A(n8701), .ZN(n8683) );
  INV_X1 U10042 ( .A(n8681), .ZN(n8682) );
  AOI21_X1 U10043 ( .B1(n8864), .B2(n8683), .A(n8682), .ZN(n8865) );
  INV_X1 U10044 ( .A(n8684), .ZN(n8685) );
  AOI22_X1 U10045 ( .A1(n10022), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8685), 
        .B2(n8827), .ZN(n8686) );
  OAI21_X1 U10046 ( .B1(n8687), .B2(n10018), .A(n8686), .ZN(n8698) );
  AOI21_X1 U10047 ( .B1(n8688), .B2(n8690), .A(n8689), .ZN(n8691) );
  NOR2_X1 U10048 ( .A1(n8691), .A2(n8803), .ZN(n8696) );
  OAI22_X1 U10049 ( .A1(n8693), .A2(n8806), .B1(n8692), .B2(n8808), .ZN(n8694)
         );
  AOI21_X1 U10050 ( .B1(n8696), .B2(n8695), .A(n8694), .ZN(n8867) );
  NOR2_X1 U10051 ( .A1(n8867), .A2(n10022), .ZN(n8697) );
  AOI211_X1 U10052 ( .C1(n8865), .C2(n8829), .A(n8698), .B(n8697), .ZN(n8699)
         );
  OAI21_X1 U10053 ( .B1(n8868), .B2(n8798), .A(n8699), .ZN(P2_U3272) );
  OAI21_X1 U10054 ( .B1(n4356), .B2(n8707), .A(n8700), .ZN(n8873) );
  AOI21_X1 U10055 ( .B1(n8869), .B2(n8716), .A(n8701), .ZN(n8870) );
  INV_X1 U10056 ( .A(n8869), .ZN(n8705) );
  INV_X1 U10057 ( .A(n8702), .ZN(n8703) );
  AOI22_X1 U10058 ( .A1(n10022), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8703), 
        .B2(n8827), .ZN(n8704) );
  OAI21_X1 U10059 ( .B1(n8705), .B2(n10018), .A(n8704), .ZN(n8713) );
  INV_X1 U10060 ( .A(n8706), .ZN(n8721) );
  OAI21_X1 U10061 ( .B1(n8721), .B2(n8708), .A(n8707), .ZN(n8709) );
  NAND2_X1 U10062 ( .A1(n8709), .A2(n8688), .ZN(n8711) );
  AOI222_X1 U10063 ( .A1(n8793), .A2(n8711), .B1(n8742), .B2(n8788), .C1(n8710), .C2(n8790), .ZN(n8872) );
  NOR2_X1 U10064 ( .A1(n8872), .A2(n10022), .ZN(n8712) );
  AOI211_X1 U10065 ( .C1(n8870), .C2(n8829), .A(n8713), .B(n8712), .ZN(n8714)
         );
  OAI21_X1 U10066 ( .B1(n8798), .B2(n8873), .A(n8714), .ZN(P2_U3273) );
  XNOR2_X1 U10067 ( .A(n8715), .B(n8723), .ZN(n8878) );
  INV_X1 U10068 ( .A(n8716), .ZN(n8717) );
  AOI21_X1 U10069 ( .B1(n8874), .B2(n4553), .A(n8717), .ZN(n8875) );
  AOI22_X1 U10070 ( .A1(n10022), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8718), 
        .B2(n8827), .ZN(n8719) );
  OAI21_X1 U10071 ( .B1(n8720), .B2(n10018), .A(n8719), .ZN(n8727) );
  AOI211_X1 U10072 ( .C1(n8723), .C2(n8722), .A(n8803), .B(n8721), .ZN(n8725)
         );
  NOR2_X1 U10073 ( .A1(n8725), .A2(n8724), .ZN(n8877) );
  NOR2_X1 U10074 ( .A1(n8877), .A2(n10022), .ZN(n8726) );
  AOI211_X1 U10075 ( .C1(n8875), .C2(n8829), .A(n8727), .B(n8726), .ZN(n8728)
         );
  OAI21_X1 U10076 ( .B1(n8798), .B2(n8878), .A(n8728), .ZN(P2_U3274) );
  NAND2_X1 U10077 ( .A1(n8885), .A2(n8730), .ZN(n8731) );
  XNOR2_X1 U10078 ( .A(n8731), .B(n8737), .ZN(n8883) );
  AOI21_X1 U10079 ( .B1(n8879), .B2(n8752), .A(n8732), .ZN(n8880) );
  INV_X1 U10080 ( .A(n8733), .ZN(n8734) );
  AOI22_X1 U10081 ( .A1(n10022), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8734), 
        .B2(n8827), .ZN(n8735) );
  OAI21_X1 U10082 ( .B1(n4551), .B2(n10018), .A(n8735), .ZN(n8745) );
  INV_X1 U10083 ( .A(n8736), .ZN(n8739) );
  OAI21_X1 U10084 ( .B1(n8739), .B2(n8738), .A(n8737), .ZN(n8741) );
  NAND2_X1 U10085 ( .A1(n8741), .A2(n8740), .ZN(n8743) );
  AOI222_X1 U10086 ( .A1(n8793), .A2(n8743), .B1(n8742), .B2(n8790), .C1(n8772), .C2(n8788), .ZN(n8882) );
  NOR2_X1 U10087 ( .A1(n8882), .A2(n10022), .ZN(n8744) );
  AOI211_X1 U10088 ( .C1(n8880), .C2(n8829), .A(n8745), .B(n8744), .ZN(n8746)
         );
  OAI21_X1 U10089 ( .B1(n8798), .B2(n8883), .A(n8746), .ZN(P2_U3275) );
  NAND2_X1 U10090 ( .A1(n8768), .A2(n8747), .ZN(n8748) );
  XNOR2_X1 U10091 ( .A(n8748), .B(n8751), .ZN(n8750) );
  AOI222_X1 U10092 ( .A1(n8793), .A2(n8750), .B1(n8749), .B2(n8790), .C1(n8791), .C2(n8788), .ZN(n8889) );
  NAND2_X1 U10093 ( .A1(n8729), .A2(n8751), .ZN(n8884) );
  NAND3_X1 U10094 ( .A1(n8885), .A2(n8884), .A3(n8825), .ZN(n8760) );
  INV_X1 U10095 ( .A(n8752), .ZN(n8753) );
  AOI21_X1 U10096 ( .B1(n8886), .B2(n8762), .A(n8753), .ZN(n8887) );
  INV_X1 U10097 ( .A(n8886), .ZN(n8757) );
  INV_X1 U10098 ( .A(n8754), .ZN(n8755) );
  AOI22_X1 U10099 ( .A1(n10022), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8755), 
        .B2(n8827), .ZN(n8756) );
  OAI21_X1 U10100 ( .B1(n8757), .B2(n10018), .A(n8756), .ZN(n8758) );
  AOI21_X1 U10101 ( .B1(n8887), .B2(n8829), .A(n8758), .ZN(n8759) );
  OAI211_X1 U10102 ( .C1(n10022), .C2(n8889), .A(n8760), .B(n8759), .ZN(
        P2_U3276) );
  XNOR2_X1 U10103 ( .A(n8761), .B(n8770), .ZN(n8895) );
  INV_X1 U10104 ( .A(n8779), .ZN(n8764) );
  INV_X1 U10105 ( .A(n8762), .ZN(n8763) );
  AOI211_X1 U10106 ( .C1(n8892), .C2(n8764), .A(n10064), .B(n8763), .ZN(n8891)
         );
  AOI22_X1 U10107 ( .A1(n10022), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8765), 
        .B2(n8827), .ZN(n8766) );
  OAI21_X1 U10108 ( .B1(n8767), .B2(n10018), .A(n8766), .ZN(n8775) );
  OAI21_X1 U10109 ( .B1(n8770), .B2(n8769), .A(n8768), .ZN(n8773) );
  AOI222_X1 U10110 ( .A1(n8793), .A2(n8773), .B1(n8772), .B2(n8790), .C1(n8771), .C2(n8788), .ZN(n8894) );
  NOR2_X1 U10111 ( .A1(n8894), .A2(n10022), .ZN(n8774) );
  AOI211_X1 U10112 ( .C1(n8891), .C2(n10011), .A(n8775), .B(n8774), .ZN(n8776)
         );
  OAI21_X1 U10113 ( .B1(n8798), .B2(n8895), .A(n8776), .ZN(P2_U3277) );
  XNOR2_X1 U10114 ( .A(n8777), .B(n8786), .ZN(n8900) );
  AND2_X1 U10115 ( .A1(n8896), .A2(n8810), .ZN(n8778) );
  NOR2_X1 U10116 ( .A1(n8779), .A2(n8778), .ZN(n8897) );
  INV_X1 U10117 ( .A(n8896), .ZN(n8781) );
  INV_X1 U10118 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8780) );
  OAI22_X1 U10119 ( .A1(n8781), .A2(n10018), .B1(n8780), .B2(n10009), .ZN(
        n8782) );
  AOI21_X1 U10120 ( .B1(n8897), .B2(n8829), .A(n8782), .ZN(n8797) );
  AND2_X1 U10121 ( .A1(n8784), .A2(n8783), .ZN(n8787) );
  OAI21_X1 U10122 ( .B1(n8787), .B2(n8786), .A(n8785), .ZN(n8792) );
  AOI222_X1 U10123 ( .A1(n8793), .A2(n8792), .B1(n8791), .B2(n8790), .C1(n8789), .C2(n8788), .ZN(n8899) );
  OAI21_X1 U10124 ( .B1(n8794), .B2(n10025), .A(n8899), .ZN(n8795) );
  NAND2_X1 U10125 ( .A1(n8795), .A2(n10009), .ZN(n8796) );
  OAI211_X1 U10126 ( .C1(n8900), .C2(n8798), .A(n8797), .B(n8796), .ZN(
        P2_U3278) );
  OAI21_X1 U10127 ( .B1(n8800), .B2(n8801), .A(n8799), .ZN(n8902) );
  INV_X1 U10128 ( .A(n8902), .ZN(n8822) );
  XNOR2_X1 U10129 ( .A(n8802), .B(n8801), .ZN(n8804) );
  OAI222_X1 U10130 ( .A1(n8808), .A2(n8807), .B1(n8806), .B2(n8805), .C1(n8804), .C2(n8803), .ZN(n8814) );
  AOI21_X1 U10131 ( .B1(n8809), .B2(n8901), .A(n10064), .ZN(n8811) );
  AOI21_X1 U10132 ( .B1(n8811), .B2(n8810), .A(n8814), .ZN(n8903) );
  OAI21_X1 U10133 ( .B1(n8822), .B2(n8812), .A(n8903), .ZN(n8813) );
  OAI211_X1 U10134 ( .C1(n8815), .C2(n8814), .A(n8813), .B(n10009), .ZN(n8820)
         );
  OAI22_X1 U10135 ( .A1(n10009), .A2(n8817), .B1(n8816), .B2(n10025), .ZN(
        n8818) );
  AOI21_X1 U10136 ( .B1(n8901), .B2(n8824), .A(n8818), .ZN(n8819) );
  OAI211_X1 U10137 ( .C1(n8822), .C2(n8821), .A(n8820), .B(n8819), .ZN(
        P2_U3279) );
  AOI22_X1 U10138 ( .A1(n8826), .A2(n8825), .B1(n8824), .B2(n8823), .ZN(n8834)
         );
  AOI22_X1 U10139 ( .A1(n8829), .A2(n8828), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n8827), .ZN(n8833) );
  MUX2_X1 U10140 ( .A(n8831), .B(n8830), .S(n10009), .Z(n8832) );
  NAND3_X1 U10141 ( .A1(n8834), .A2(n8833), .A3(n8832), .ZN(P2_U3294) );
  AOI22_X1 U10142 ( .A1(n8836), .A2(n9683), .B1(n9677), .B2(n8835), .ZN(n8837)
         );
  OAI211_X1 U10143 ( .C1(n8839), .C2(n8914), .A(n8838), .B(n8837), .ZN(n8916)
         );
  MUX2_X1 U10144 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8916), .S(n10080), .Z(
        P2_U3549) );
  AOI22_X1 U10145 ( .A1(n8841), .A2(n9683), .B1(n9677), .B2(n8840), .ZN(n8842)
         );
  OAI211_X1 U10146 ( .C1(n8844), .C2(n8914), .A(n8843), .B(n8842), .ZN(n8917)
         );
  MUX2_X1 U10147 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8917), .S(n10080), .Z(
        P2_U3548) );
  OAI22_X1 U10148 ( .A1(n8846), .A2(n10064), .B1(n8845), .B2(n10062), .ZN(
        n8847) );
  AOI211_X1 U10149 ( .C1(n8849), .C2(n10068), .A(n8848), .B(n8847), .ZN(n8850)
         );
  INV_X1 U10150 ( .A(n8850), .ZN(n8918) );
  MUX2_X1 U10151 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8918), .S(n10080), .Z(
        P2_U3547) );
  NAND2_X1 U10152 ( .A1(n8851), .A2(n9677), .ZN(n8853) );
  NAND3_X1 U10153 ( .A1(n8854), .A2(n8853), .A3(n8852), .ZN(n8855) );
  AOI21_X1 U10154 ( .B1(n8856), .B2(n10068), .A(n8855), .ZN(n8920) );
  INV_X1 U10155 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8857) );
  MUX2_X1 U10156 ( .A(n8920), .B(n8857), .S(n10078), .Z(n8858) );
  INV_X1 U10157 ( .A(n8858), .ZN(P2_U3546) );
  AOI21_X1 U10158 ( .B1(n9677), .B2(n8860), .A(n8859), .ZN(n8861) );
  OAI211_X1 U10159 ( .C1(n8863), .C2(n8914), .A(n8862), .B(n8861), .ZN(n8922)
         );
  MUX2_X1 U10160 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8922), .S(n10080), .Z(
        P2_U3545) );
  AOI22_X1 U10161 ( .A1(n8865), .A2(n9683), .B1(n9677), .B2(n8864), .ZN(n8866)
         );
  OAI211_X1 U10162 ( .C1(n8868), .C2(n8914), .A(n8867), .B(n8866), .ZN(n8923)
         );
  MUX2_X1 U10163 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8923), .S(n10080), .Z(
        P2_U3544) );
  AOI22_X1 U10164 ( .A1(n8870), .A2(n9683), .B1(n9677), .B2(n8869), .ZN(n8871)
         );
  OAI211_X1 U10165 ( .C1(n8873), .C2(n8914), .A(n8872), .B(n8871), .ZN(n8924)
         );
  MUX2_X1 U10166 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8924), .S(n10080), .Z(
        P2_U3543) );
  AOI22_X1 U10167 ( .A1(n8875), .A2(n9683), .B1(n9677), .B2(n8874), .ZN(n8876)
         );
  OAI211_X1 U10168 ( .C1(n8878), .C2(n8914), .A(n8877), .B(n8876), .ZN(n8925)
         );
  MUX2_X1 U10169 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8925), .S(n10080), .Z(
        P2_U3542) );
  AOI22_X1 U10170 ( .A1(n8880), .A2(n9683), .B1(n9677), .B2(n8879), .ZN(n8881)
         );
  OAI211_X1 U10171 ( .C1(n8883), .C2(n8914), .A(n8882), .B(n8881), .ZN(n8926)
         );
  MUX2_X1 U10172 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8926), .S(n10080), .Z(
        P2_U3541) );
  NAND3_X1 U10173 ( .A1(n8885), .A2(n10068), .A3(n8884), .ZN(n8890) );
  AOI22_X1 U10174 ( .A1(n8887), .A2(n9683), .B1(n9677), .B2(n8886), .ZN(n8888)
         );
  NAND3_X1 U10175 ( .A1(n8890), .A2(n8889), .A3(n8888), .ZN(n8927) );
  MUX2_X1 U10176 ( .A(n8927), .B(P2_REG1_REG_20__SCAN_IN), .S(n10078), .Z(
        P2_U3540) );
  AOI21_X1 U10177 ( .B1(n9677), .B2(n8892), .A(n8891), .ZN(n8893) );
  OAI211_X1 U10178 ( .C1(n8895), .C2(n8914), .A(n8894), .B(n8893), .ZN(n8928)
         );
  MUX2_X1 U10179 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8928), .S(n10080), .Z(
        P2_U3539) );
  AOI22_X1 U10180 ( .A1(n8897), .A2(n9683), .B1(n9677), .B2(n8896), .ZN(n8898)
         );
  OAI211_X1 U10181 ( .C1(n8900), .C2(n8914), .A(n8899), .B(n8898), .ZN(n8929)
         );
  MUX2_X1 U10182 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8929), .S(n10080), .Z(
        P2_U3538) );
  AOI22_X1 U10183 ( .A1(n8902), .A2(n10068), .B1(n9677), .B2(n8901), .ZN(n8904) );
  NAND2_X1 U10184 ( .A1(n8904), .A2(n8903), .ZN(n8930) );
  MUX2_X1 U10185 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8930), .S(n10080), .Z(
        P2_U3537) );
  AOI22_X1 U10186 ( .A1(n8906), .A2(n9683), .B1(n9677), .B2(n8905), .ZN(n8907)
         );
  OAI211_X1 U10187 ( .C1(n8909), .C2(n8914), .A(n8908), .B(n8907), .ZN(n8931)
         );
  MUX2_X1 U10188 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8931), .S(n10080), .Z(
        P2_U3536) );
  AOI22_X1 U10189 ( .A1(n8911), .A2(n9683), .B1(n9677), .B2(n8910), .ZN(n8912)
         );
  OAI211_X1 U10190 ( .C1(n8915), .C2(n8914), .A(n8913), .B(n8912), .ZN(n8932)
         );
  MUX2_X1 U10191 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8932), .S(n10080), .Z(
        P2_U3535) );
  MUX2_X1 U10192 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8916), .S(n4316), .Z(
        P2_U3517) );
  MUX2_X1 U10193 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8917), .S(n4316), .Z(
        P2_U3516) );
  MUX2_X1 U10194 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8918), .S(n4316), .Z(
        P2_U3515) );
  MUX2_X1 U10195 ( .A(n8920), .B(n8919), .S(n10070), .Z(n8921) );
  INV_X1 U10196 ( .A(n8921), .ZN(P2_U3514) );
  MUX2_X1 U10197 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8922), .S(n4316), .Z(
        P2_U3513) );
  MUX2_X1 U10198 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8923), .S(n4316), .Z(
        P2_U3512) );
  MUX2_X1 U10199 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8924), .S(n4316), .Z(
        P2_U3511) );
  MUX2_X1 U10200 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8925), .S(n4316), .Z(
        P2_U3510) );
  MUX2_X1 U10201 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8926), .S(n4316), .Z(
        P2_U3509) );
  MUX2_X1 U10202 ( .A(n8927), .B(P2_REG0_REG_20__SCAN_IN), .S(n10070), .Z(
        P2_U3508) );
  MUX2_X1 U10203 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8928), .S(n4316), .Z(
        P2_U3507) );
  MUX2_X1 U10204 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8929), .S(n4316), .Z(
        P2_U3505) );
  MUX2_X1 U10205 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8930), .S(n4316), .Z(
        P2_U3502) );
  MUX2_X1 U10206 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8931), .S(n4316), .Z(
        P2_U3499) );
  MUX2_X1 U10207 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8932), .S(n4316), .Z(
        P2_U3496) );
  INV_X1 U10208 ( .A(n8933), .ZN(n9437) );
  NOR4_X1 U10209 ( .A1(n4663), .A2(P2_IR_REG_30__SCAN_IN), .A3(n5093), .A4(
        P2_U3152), .ZN(n8934) );
  AOI21_X1 U10210 ( .B1(n8943), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8934), .ZN(
        n8935) );
  OAI21_X1 U10211 ( .B1(n9437), .B2(n8946), .A(n8935), .ZN(P2_U3327) );
  AOI22_X1 U10212 ( .A1(n8936), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8943), .ZN(n8937) );
  OAI21_X1 U10213 ( .B1(n8938), .B2(n8946), .A(n8937), .ZN(P2_U3328) );
  AOI22_X1 U10214 ( .A1(n8939), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n8943), .ZN(n8940) );
  OAI21_X1 U10215 ( .B1(n8941), .B2(n8946), .A(n8940), .ZN(P2_U3329) );
  INV_X1 U10216 ( .A(n8942), .ZN(n9439) );
  NAND2_X1 U10217 ( .A1(n8943), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8944) );
  OAI211_X1 U10218 ( .C1(n9439), .C2(n8946), .A(n8945), .B(n8944), .ZN(
        P2_U3330) );
  INV_X1 U10219 ( .A(n6158), .ZN(n9444) );
  OAI222_X1 U10220 ( .A1(n8946), .A2(n9444), .B1(P2_U3152), .B2(n8949), .C1(
        n8948), .C2(n8947), .ZN(P2_U3331) );
  MUX2_X1 U10221 ( .A(n8950), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U10222 ( .A(n8951), .ZN(n8955) );
  AOI21_X1 U10223 ( .B1(n8953), .B2(n4732), .A(n8952), .ZN(n8954) );
  AOI21_X1 U10224 ( .B1(n9012), .B2(n8955), .A(n8954), .ZN(n8961) );
  INV_X1 U10225 ( .A(n9239), .ZN(n8958) );
  NAND2_X1 U10226 ( .A1(n9233), .A2(n9024), .ZN(n8957) );
  AOI22_X1 U10227 ( .A1(n9265), .A2(n9048), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8956) );
  OAI211_X1 U10228 ( .C1(n9050), .C2(n8958), .A(n8957), .B(n8956), .ZN(n8959)
         );
  AOI21_X1 U10229 ( .B1(n9363), .B2(n9052), .A(n8959), .ZN(n8960) );
  OAI21_X1 U10230 ( .B1(n8961), .B2(n9054), .A(n8960), .ZN(P1_U3214) );
  XOR2_X1 U10231 ( .A(n8963), .B(n8962), .Z(n8968) );
  NAND2_X1 U10232 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9145) );
  OAI21_X1 U10233 ( .B1(n8972), .B2(n9062), .A(n9145), .ZN(n8964) );
  AOI21_X1 U10234 ( .B1(n9048), .B2(n9299), .A(n8964), .ZN(n8965) );
  OAI21_X1 U10235 ( .B1(n9050), .B2(n9292), .A(n8965), .ZN(n8966) );
  AOI21_X1 U10236 ( .B1(n9384), .B2(n9052), .A(n8966), .ZN(n8967) );
  OAI21_X1 U10237 ( .B1(n8968), .B2(n9054), .A(n8967), .ZN(P1_U3217) );
  XOR2_X1 U10238 ( .A(n8970), .B(n8969), .Z(n8977) );
  OAI22_X1 U10239 ( .A1(n8972), .A2(n9060), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8971), .ZN(n8973) );
  AOI21_X1 U10240 ( .B1(n9024), .B2(n9265), .A(n8973), .ZN(n8974) );
  OAI21_X1 U10241 ( .B1(n9050), .B2(n9271), .A(n8974), .ZN(n8975) );
  AOI21_X1 U10242 ( .B1(n9372), .B2(n9052), .A(n8975), .ZN(n8976) );
  OAI21_X1 U10243 ( .B1(n8977), .B2(n9054), .A(n8976), .ZN(P1_U3221) );
  XOR2_X1 U10244 ( .A(n8979), .B(n8978), .Z(n8985) );
  NOR2_X1 U10245 ( .A1(n8980), .A2(n9062), .ZN(n8983) );
  AOI22_X1 U10246 ( .A1(n9233), .A2(n9048), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8981) );
  OAI21_X1 U10247 ( .B1(n9050), .B2(n9201), .A(n8981), .ZN(n8982) );
  AOI211_X1 U10248 ( .C1(n9351), .C2(n9052), .A(n8983), .B(n8982), .ZN(n8984)
         );
  OAI21_X1 U10249 ( .B1(n8985), .B2(n9054), .A(n8984), .ZN(P1_U3223) );
  INV_X1 U10250 ( .A(n8986), .ZN(n8990) );
  NAND2_X1 U10251 ( .A1(n4336), .A2(n8989), .ZN(n8987) );
  AOI22_X1 U10252 ( .A1(n8990), .A2(n8989), .B1(n8988), .B2(n8987), .ZN(n8998)
         );
  NAND2_X1 U10253 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9111) );
  INV_X1 U10254 ( .A(n9111), .ZN(n8993) );
  NOR2_X1 U10255 ( .A1(n9060), .A2(n8991), .ZN(n8992) );
  AOI211_X1 U10256 ( .C1(n9024), .C2(n9320), .A(n8993), .B(n8992), .ZN(n8994)
         );
  OAI21_X1 U10257 ( .B1(n9050), .B2(n8995), .A(n8994), .ZN(n8996) );
  AOI21_X1 U10258 ( .B1(n9401), .B2(n9052), .A(n8996), .ZN(n8997) );
  OAI21_X1 U10259 ( .B1(n8998), .B2(n9054), .A(n8997), .ZN(P1_U3224) );
  OAI21_X1 U10260 ( .B1(n9001), .B2(n9000), .A(n8999), .ZN(n9002) );
  NAND2_X1 U10261 ( .A1(n9002), .A2(n6223), .ZN(n9009) );
  NOR2_X1 U10262 ( .A1(n9003), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9122) );
  AOI21_X1 U10263 ( .B1(n9024), .B2(n9299), .A(n9122), .ZN(n9004) );
  OAI21_X1 U10264 ( .B1(n9005), .B2(n9060), .A(n9004), .ZN(n9006) );
  AOI21_X1 U10265 ( .B1(n9007), .B2(n9066), .A(n9006), .ZN(n9008) );
  OAI211_X1 U10266 ( .C1(n9010), .C2(n9069), .A(n9009), .B(n9008), .ZN(
        P1_U3226) );
  OAI21_X1 U10267 ( .B1(n9013), .B2(n9012), .A(n9011), .ZN(n9014) );
  NAND2_X1 U10268 ( .A1(n9014), .A2(n6223), .ZN(n9018) );
  AOI22_X1 U10269 ( .A1(n9217), .A2(n9024), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        n10130), .ZN(n9015) );
  OAI21_X1 U10270 ( .B1(n9050), .B2(n9224), .A(n9015), .ZN(n9016) );
  AOI21_X1 U10271 ( .B1(n9048), .B2(n9254), .A(n9016), .ZN(n9017) );
  OAI211_X1 U10272 ( .C1(n9019), .C2(n9069), .A(n9018), .B(n9017), .ZN(
        P1_U3227) );
  NAND2_X1 U10273 ( .A1(n9021), .A2(n9020), .ZN(n9022) );
  XOR2_X1 U10274 ( .A(n9023), .B(n9022), .Z(n9029) );
  AOI22_X1 U10275 ( .A1(n9285), .A2(n9024), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        n10130), .ZN(n9026) );
  NAND2_X1 U10276 ( .A1(n9048), .A2(n9319), .ZN(n9025) );
  OAI211_X1 U10277 ( .C1(n9050), .C2(n9279), .A(n9026), .B(n9025), .ZN(n9027)
         );
  AOI21_X1 U10278 ( .B1(n9379), .B2(n9052), .A(n9027), .ZN(n9028) );
  OAI21_X1 U10279 ( .B1(n9029), .B2(n9054), .A(n9028), .ZN(P1_U3231) );
  NAND2_X1 U10280 ( .A1(n9031), .A2(n9030), .ZN(n9032) );
  XOR2_X1 U10281 ( .A(n9033), .B(n9032), .Z(n9041) );
  OAI22_X1 U10282 ( .A1(n9035), .A2(n9060), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9034), .ZN(n9036) );
  AOI21_X1 U10283 ( .B1(n9249), .B2(n9066), .A(n9036), .ZN(n9037) );
  OAI21_X1 U10284 ( .B1(n9038), .B2(n9062), .A(n9037), .ZN(n9039) );
  AOI21_X1 U10285 ( .B1(n9366), .B2(n9052), .A(n9039), .ZN(n9040) );
  OAI21_X1 U10286 ( .B1(n9041), .B2(n9054), .A(n9040), .ZN(P1_U3233) );
  XNOR2_X1 U10287 ( .A(n9043), .B(n9042), .ZN(n9044) );
  XNOR2_X1 U10288 ( .A(n9045), .B(n9044), .ZN(n9055) );
  NAND2_X1 U10289 ( .A1(n10130), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9883) );
  OAI21_X1 U10290 ( .B1(n9046), .B2(n9062), .A(n9883), .ZN(n9047) );
  AOI21_X1 U10291 ( .B1(n9048), .B2(n9320), .A(n9047), .ZN(n9049) );
  OAI21_X1 U10292 ( .B1(n9050), .B2(n9310), .A(n9049), .ZN(n9051) );
  AOI21_X1 U10293 ( .B1(n9389), .B2(n9052), .A(n9051), .ZN(n9053) );
  OAI21_X1 U10294 ( .B1(n9055), .B2(n9054), .A(n9053), .ZN(P1_U3236) );
  OAI211_X1 U10295 ( .C1(n9058), .C2(n9057), .A(n9056), .B(n6223), .ZN(n9068)
         );
  OAI22_X1 U10296 ( .A1(n9061), .A2(n9060), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9059), .ZN(n9065) );
  NOR2_X1 U10297 ( .A1(n9063), .A2(n9062), .ZN(n9064) );
  AOI211_X1 U10298 ( .C1(n9189), .C2(n9066), .A(n9065), .B(n9064), .ZN(n9067)
         );
  OAI211_X1 U10299 ( .C1(n9191), .C2(n9069), .A(n9068), .B(n9067), .ZN(
        P1_U3238) );
  MUX2_X1 U10300 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9070), .S(P1_U4006), .Z(
        P1_U3585) );
  INV_X1 U10301 ( .A(n9071), .ZN(n9171) );
  MUX2_X1 U10302 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9171), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10303 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9180), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10304 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9194), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10305 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9208), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10306 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9217), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10307 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9233), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10308 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9254), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10309 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9265), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10310 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9285), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10311 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9298), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10312 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9319), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10313 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9299), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10314 ( .A(n9320), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9084), .Z(
        P1_U3572) );
  MUX2_X1 U10315 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9072), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10316 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9073), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10317 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9708), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10318 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9074), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10319 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9711), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10320 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9075), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10321 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9076), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10322 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9077), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10323 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9078), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10324 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9079), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10325 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9080), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10326 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9081), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10327 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9082), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10328 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9083), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10329 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n5692), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10330 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6259), .S(P1_U4006), .Z(
        P1_U3556) );
  MUX2_X1 U10331 ( .A(n6258), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9084), .Z(
        P1_U3555) );
  OAI21_X1 U10332 ( .B1(n9087), .B2(n9086), .A(n9085), .ZN(n9088) );
  NAND2_X1 U10333 ( .A1(n9088), .A2(n9894), .ZN(n9098) );
  NOR2_X1 U10334 ( .A1(n9114), .A2(n9089), .ZN(n9090) );
  AOI211_X1 U10335 ( .C1(n9880), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n9091), .B(
        n9090), .ZN(n9097) );
  OAI21_X1 U10336 ( .B1(n9094), .B2(n9093), .A(n9092), .ZN(n9095) );
  NAND2_X1 U10337 ( .A1(n9095), .A2(n9895), .ZN(n9096) );
  NAND3_X1 U10338 ( .A1(n9098), .A2(n9097), .A3(n9096), .ZN(P1_U3252) );
  NOR2_X1 U10339 ( .A1(n9099), .A2(n9106), .ZN(n9101) );
  NAND2_X1 U10340 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9124), .ZN(n9102) );
  OAI21_X1 U10341 ( .B1(n9124), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9102), .ZN(
        n9103) );
  AOI211_X1 U10342 ( .C1(n9104), .C2(n9103), .A(n9123), .B(n9872), .ZN(n9117)
         );
  NOR2_X1 U10343 ( .A1(n9106), .A2(n9105), .ZN(n9108) );
  XNOR2_X1 U10344 ( .A(n9124), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9109) );
  AOI211_X1 U10345 ( .C1(n9110), .C2(n9109), .A(n9118), .B(n9843), .ZN(n9116)
         );
  NAND2_X1 U10346 ( .A1(n9880), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9112) );
  OAI211_X1 U10347 ( .C1(n9114), .C2(n9113), .A(n9112), .B(n9111), .ZN(n9115)
         );
  OR3_X1 U10348 ( .A1(n9117), .A2(n9116), .A3(n9115), .ZN(P1_U3257) );
  INV_X1 U10349 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9131) );
  XNOR2_X1 U10350 ( .A(n9138), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9119) );
  AOI211_X1 U10351 ( .C1(n9120), .C2(n9119), .A(n9137), .B(n9843), .ZN(n9121)
         );
  AOI211_X1 U10352 ( .C1(n9886), .C2(n9138), .A(n9122), .B(n9121), .ZN(n9130)
         );
  NAND2_X1 U10353 ( .A1(n9138), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9125) );
  OAI21_X1 U10354 ( .B1(n9138), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9125), .ZN(
        n9126) );
  AOI211_X1 U10355 ( .C1(n9127), .C2(n9126), .A(n9132), .B(n9872), .ZN(n9128)
         );
  INV_X1 U10356 ( .A(n9128), .ZN(n9129) );
  OAI211_X1 U10357 ( .C1(n9131), .C2(n9899), .A(n9130), .B(n9129), .ZN(
        P1_U3258) );
  INV_X1 U10358 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9146) );
  AOI21_X1 U10359 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n9138), .A(n9132), .ZN(
        n9889) );
  NAND2_X1 U10360 ( .A1(n9885), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9133) );
  OAI21_X1 U10361 ( .B1(n9885), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9133), .ZN(
        n9888) );
  NOR2_X1 U10362 ( .A1(n9889), .A2(n9888), .ZN(n9887) );
  AOI21_X1 U10363 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n9885), .A(n9887), .ZN(
        n9134) );
  XNOR2_X1 U10364 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9134), .ZN(n9143) );
  AOI22_X1 U10365 ( .A1(n9885), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n9136), .B2(
        n9135), .ZN(n9892) );
  AOI21_X1 U10366 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n9138), .A(n9137), .ZN(
        n9891) );
  NAND2_X1 U10367 ( .A1(n9892), .A2(n9891), .ZN(n9890) );
  OAI21_X1 U10368 ( .B1(n9885), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9890), .ZN(
        n9140) );
  INV_X1 U10369 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9139) );
  XOR2_X1 U10370 ( .A(n9140), .B(n9139), .Z(n9141) );
  AOI22_X1 U10371 ( .A1(n9143), .A2(n9895), .B1(n9894), .B2(n9141), .ZN(n9144)
         );
  NAND2_X1 U10372 ( .A1(n9155), .A2(n9154), .ZN(n9147) );
  XNOR2_X2 U10373 ( .A(n9147), .B(n9671), .ZN(n9669) );
  INV_X1 U10374 ( .A(n9148), .ZN(n9150) );
  NOR2_X1 U10375 ( .A1(n9150), .A2(n9149), .ZN(n9743) );
  INV_X1 U10376 ( .A(n9743), .ZN(n9151) );
  NOR2_X1 U10377 ( .A1(n9736), .A2(n9151), .ZN(n9157) );
  AOI21_X1 U10378 ( .B1(n9736), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9157), .ZN(
        n9153) );
  NAND2_X1 U10379 ( .A1(n9671), .A2(n9739), .ZN(n9152) );
  OAI211_X1 U10380 ( .C1(n9669), .C2(n9159), .A(n9153), .B(n9152), .ZN(
        P1_U3261) );
  NOR2_X1 U10381 ( .A1(n9155), .A2(n9924), .ZN(n9156) );
  AOI211_X1 U10382 ( .C1(n9736), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9157), .B(
        n9156), .ZN(n9158) );
  OAI21_X1 U10383 ( .B1(n9159), .B2(n9742), .A(n9158), .ZN(P1_U3262) );
  INV_X1 U10384 ( .A(n9175), .ZN(n9162) );
  INV_X1 U10385 ( .A(n9160), .ZN(n9161) );
  AOI21_X1 U10386 ( .B1(n9336), .B2(n9162), .A(n9161), .ZN(n9337) );
  AOI22_X1 U10387 ( .A1(n9163), .A2(n9311), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9736), .ZN(n9164) );
  OAI21_X1 U10388 ( .B1(n9165), .B2(n9924), .A(n9164), .ZN(n9173) );
  OAI21_X1 U10389 ( .B1(n9170), .B2(n9169), .A(n9168), .ZN(n9172) );
  XOR2_X1 U10390 ( .A(n9179), .B(n9174), .Z(n9345) );
  AOI21_X1 U10391 ( .B1(n9341), .B2(n9186), .A(n9175), .ZN(n9342) );
  AOI22_X1 U10392 ( .A1(n9176), .A2(n9311), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9736), .ZN(n9177) );
  OAI21_X1 U10393 ( .B1(n4766), .B2(n9924), .A(n9177), .ZN(n9183) );
  XOR2_X1 U10394 ( .A(n9179), .B(n9178), .Z(n9181) );
  AOI222_X1 U10395 ( .A1(n9919), .A2(n9181), .B1(n9208), .B2(n9710), .C1(n9180), .C2(n9709), .ZN(n9344) );
  NOR2_X1 U10396 ( .A1(n9344), .A2(n9736), .ZN(n9182) );
  AOI211_X1 U10397 ( .C1(n9908), .C2(n9342), .A(n9183), .B(n9182), .ZN(n9184)
         );
  OAI21_X1 U10398 ( .B1(n9345), .B2(n9325), .A(n9184), .ZN(P1_U3264) );
  XNOR2_X1 U10399 ( .A(n9185), .B(n9192), .ZN(n9350) );
  INV_X1 U10400 ( .A(n9200), .ZN(n9188) );
  INV_X1 U10401 ( .A(n9186), .ZN(n9187) );
  AOI21_X1 U10402 ( .B1(n9346), .B2(n9188), .A(n9187), .ZN(n9347) );
  AOI22_X1 U10403 ( .A1(n9189), .A2(n9311), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9736), .ZN(n9190) );
  OAI21_X1 U10404 ( .B1(n9191), .B2(n9924), .A(n9190), .ZN(n9197) );
  XNOR2_X1 U10405 ( .A(n9193), .B(n9192), .ZN(n9195) );
  AOI222_X1 U10406 ( .A1(n9919), .A2(n9195), .B1(n9217), .B2(n9710), .C1(n9194), .C2(n9709), .ZN(n9349) );
  NOR2_X1 U10407 ( .A1(n9349), .A2(n9736), .ZN(n9196) );
  AOI211_X1 U10408 ( .C1(n9347), .C2(n9908), .A(n9197), .B(n9196), .ZN(n9198)
         );
  OAI21_X1 U10409 ( .B1(n9350), .B2(n9325), .A(n9198), .ZN(P1_U3265) );
  XOR2_X1 U10410 ( .A(n9206), .B(n9199), .Z(n9355) );
  AOI21_X1 U10411 ( .B1(n9351), .B2(n9219), .A(n9200), .ZN(n9352) );
  INV_X1 U10412 ( .A(n9351), .ZN(n9204) );
  INV_X1 U10413 ( .A(n9201), .ZN(n9202) );
  AOI22_X1 U10414 ( .A1(n9202), .A2(n9311), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9736), .ZN(n9203) );
  OAI21_X1 U10415 ( .B1(n9204), .B2(n9924), .A(n9203), .ZN(n9211) );
  NAND2_X1 U10416 ( .A1(n9214), .A2(n9205), .ZN(n9207) );
  XNOR2_X1 U10417 ( .A(n9207), .B(n9206), .ZN(n9209) );
  AOI222_X1 U10418 ( .A1(n9919), .A2(n9209), .B1(n9233), .B2(n9710), .C1(n9208), .C2(n9709), .ZN(n9354) );
  NOR2_X1 U10419 ( .A1(n9354), .A2(n9736), .ZN(n9210) );
  AOI211_X1 U10420 ( .C1(n9352), .C2(n9908), .A(n9211), .B(n9210), .ZN(n9212)
         );
  OAI21_X1 U10421 ( .B1(n9355), .B2(n9325), .A(n9212), .ZN(P1_U3266) );
  XOR2_X1 U10422 ( .A(n9215), .B(n9213), .Z(n9360) );
  AOI22_X1 U10423 ( .A1(n9357), .A2(n9739), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9736), .ZN(n9227) );
  OAI21_X1 U10424 ( .B1(n9216), .B2(n9215), .A(n9214), .ZN(n9218) );
  AOI222_X1 U10425 ( .A1(n9919), .A2(n9218), .B1(n9217), .B2(n9709), .C1(n9254), .C2(n9710), .ZN(n9359) );
  INV_X1 U10426 ( .A(n9237), .ZN(n9221) );
  INV_X1 U10427 ( .A(n9219), .ZN(n9220) );
  AOI211_X1 U10428 ( .C1(n9357), .C2(n9221), .A(n9973), .B(n9220), .ZN(n9356)
         );
  NAND2_X1 U10429 ( .A1(n9356), .A2(n9222), .ZN(n9223) );
  OAI211_X1 U10430 ( .C1(n9925), .C2(n9224), .A(n9359), .B(n9223), .ZN(n9225)
         );
  NAND2_X1 U10431 ( .A1(n9225), .A2(n9930), .ZN(n9226) );
  OAI211_X1 U10432 ( .C1(n9360), .C2(n9325), .A(n9227), .B(n9226), .ZN(
        P1_U3267) );
  XNOR2_X1 U10433 ( .A(n9229), .B(n9228), .ZN(n9365) );
  INV_X1 U10434 ( .A(n9230), .ZN(n9232) );
  OAI21_X1 U10435 ( .B1(n9232), .B2(n9231), .A(n9919), .ZN(n9236) );
  AOI22_X1 U10436 ( .A1(n9233), .A2(n9709), .B1(n9710), .B2(n9265), .ZN(n9234)
         );
  OAI21_X1 U10437 ( .B1(n9236), .B2(n9235), .A(n9234), .ZN(n9361) );
  AOI211_X1 U10438 ( .C1(n9363), .C2(n9246), .A(n9973), .B(n9237), .ZN(n9362)
         );
  NAND2_X1 U10439 ( .A1(n9362), .A2(n9238), .ZN(n9241) );
  AOI22_X1 U10440 ( .A1(P1_REG2_REG_23__SCAN_IN), .A2(n9736), .B1(n9239), .B2(
        n9311), .ZN(n9240) );
  OAI211_X1 U10441 ( .C1(n9242), .C2(n9924), .A(n9241), .B(n9240), .ZN(n9243)
         );
  AOI21_X1 U10442 ( .B1(n9361), .B2(n9930), .A(n9243), .ZN(n9244) );
  OAI21_X1 U10443 ( .B1(n9365), .B2(n9325), .A(n9244), .ZN(P1_U3268) );
  XNOR2_X1 U10444 ( .A(n9245), .B(n9253), .ZN(n9370) );
  INV_X1 U10445 ( .A(n9269), .ZN(n9248) );
  INV_X1 U10446 ( .A(n9246), .ZN(n9247) );
  AOI21_X1 U10447 ( .B1(n9366), .B2(n9248), .A(n9247), .ZN(n9367) );
  AOI22_X1 U10448 ( .A1(n9736), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9249), .B2(
        n9311), .ZN(n9250) );
  OAI21_X1 U10449 ( .B1(n9251), .B2(n9924), .A(n9250), .ZN(n9257) );
  XOR2_X1 U10450 ( .A(n9253), .B(n9252), .Z(n9255) );
  AOI222_X1 U10451 ( .A1(n9919), .A2(n9255), .B1(n9254), .B2(n9709), .C1(n9285), .C2(n9710), .ZN(n9369) );
  NOR2_X1 U10452 ( .A1(n9369), .A2(n9736), .ZN(n9256) );
  AOI211_X1 U10453 ( .C1(n9367), .C2(n9908), .A(n9257), .B(n9256), .ZN(n9258)
         );
  OAI21_X1 U10454 ( .B1(n9325), .B2(n9370), .A(n9258), .ZN(P1_U3269) );
  INV_X1 U10455 ( .A(n9261), .ZN(n9260) );
  XNOR2_X1 U10456 ( .A(n9259), .B(n9260), .ZN(n9371) );
  INV_X1 U10457 ( .A(n9371), .ZN(n9276) );
  AOI22_X1 U10458 ( .A1(n9372), .A2(n9739), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9736), .ZN(n9275) );
  AND2_X1 U10459 ( .A1(n9262), .A2(n9261), .ZN(n9263) );
  OAI21_X1 U10460 ( .B1(n9264), .B2(n9263), .A(n9919), .ZN(n9267) );
  AOI22_X1 U10461 ( .A1(n9265), .A2(n9709), .B1(n9710), .B2(n9298), .ZN(n9266)
         );
  NAND2_X1 U10462 ( .A1(n9267), .A2(n9266), .ZN(n9376) );
  OAI21_X1 U10463 ( .B1(n9278), .B2(n9268), .A(n9395), .ZN(n9270) );
  OR2_X1 U10464 ( .A1(n9270), .A2(n9269), .ZN(n9374) );
  OAI22_X1 U10465 ( .A1(n9374), .A2(n9272), .B1(n9925), .B2(n9271), .ZN(n9273)
         );
  OAI21_X1 U10466 ( .B1(n9376), .B2(n9273), .A(n9930), .ZN(n9274) );
  OAI211_X1 U10467 ( .C1(n9276), .C2(n9325), .A(n9275), .B(n9274), .ZN(
        P1_U3270) );
  XOR2_X1 U10468 ( .A(n9277), .B(n9284), .Z(n9383) );
  AOI21_X1 U10469 ( .B1(n9379), .B2(n9291), .A(n9278), .ZN(n9380) );
  INV_X1 U10470 ( .A(n9379), .ZN(n9282) );
  INV_X1 U10471 ( .A(n9279), .ZN(n9280) );
  AOI22_X1 U10472 ( .A1(n9736), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9280), .B2(
        n9311), .ZN(n9281) );
  OAI21_X1 U10473 ( .B1(n9282), .B2(n9924), .A(n9281), .ZN(n9288) );
  XOR2_X1 U10474 ( .A(n9284), .B(n9283), .Z(n9286) );
  AOI222_X1 U10475 ( .A1(n9919), .A2(n9286), .B1(n9319), .B2(n9710), .C1(n9285), .C2(n9709), .ZN(n9382) );
  NOR2_X1 U10476 ( .A1(n9382), .A2(n9736), .ZN(n9287) );
  AOI211_X1 U10477 ( .C1(n9380), .C2(n9908), .A(n9288), .B(n9287), .ZN(n9289)
         );
  OAI21_X1 U10478 ( .B1(n9383), .B2(n9325), .A(n9289), .ZN(P1_U3271) );
  XOR2_X1 U10479 ( .A(n9290), .B(n9296), .Z(n9388) );
  AOI21_X1 U10480 ( .B1(n9384), .B2(n9308), .A(n4642), .ZN(n9385) );
  INV_X1 U10481 ( .A(n9384), .ZN(n9295) );
  INV_X1 U10482 ( .A(n9292), .ZN(n9293) );
  AOI22_X1 U10483 ( .A1(n9736), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9293), .B2(
        n9311), .ZN(n9294) );
  OAI21_X1 U10484 ( .B1(n9295), .B2(n9924), .A(n9294), .ZN(n9302) );
  XNOR2_X1 U10485 ( .A(n9297), .B(n9296), .ZN(n9300) );
  AOI222_X1 U10486 ( .A1(n9919), .A2(n9300), .B1(n9299), .B2(n9710), .C1(n9298), .C2(n9709), .ZN(n9387) );
  NOR2_X1 U10487 ( .A1(n9387), .A2(n9736), .ZN(n9301) );
  AOI211_X1 U10488 ( .C1(n9385), .C2(n9908), .A(n9302), .B(n9301), .ZN(n9303)
         );
  OAI21_X1 U10489 ( .B1(n9388), .B2(n9325), .A(n9303), .ZN(P1_U3272) );
  AND2_X1 U10490 ( .A1(n9305), .A2(n9304), .ZN(n9306) );
  XNOR2_X1 U10491 ( .A(n9306), .B(n9317), .ZN(n9393) );
  INV_X1 U10492 ( .A(n9307), .ZN(n9309) );
  AOI21_X1 U10493 ( .B1(n9389), .B2(n9309), .A(n4643), .ZN(n9390) );
  INV_X1 U10494 ( .A(n9310), .ZN(n9312) );
  AOI22_X1 U10495 ( .A1(n9736), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9312), .B2(
        n9311), .ZN(n9313) );
  OAI21_X1 U10496 ( .B1(n9314), .B2(n9924), .A(n9313), .ZN(n9323) );
  NAND2_X1 U10497 ( .A1(n9316), .A2(n9315), .ZN(n9318) );
  XNOR2_X1 U10498 ( .A(n9318), .B(n9317), .ZN(n9321) );
  AOI222_X1 U10499 ( .A1(n9919), .A2(n9321), .B1(n9320), .B2(n9710), .C1(n9319), .C2(n9709), .ZN(n9392) );
  NOR2_X1 U10500 ( .A1(n9392), .A2(n9736), .ZN(n9322) );
  AOI211_X1 U10501 ( .C1(n9390), .C2(n9908), .A(n9323), .B(n9322), .ZN(n9324)
         );
  OAI21_X1 U10502 ( .B1(n9325), .B2(n9393), .A(n9324), .ZN(P1_U3273) );
  OR2_X1 U10503 ( .A1(n9326), .A2(n9736), .ZN(n9335) );
  OAI22_X1 U10504 ( .A1(n9930), .A2(n5676), .B1(n9327), .B2(n9925), .ZN(n9328)
         );
  AOI21_X1 U10505 ( .B1(n9739), .B2(n9329), .A(n9328), .ZN(n9334) );
  NAND2_X1 U10506 ( .A1(n9330), .A2(n9909), .ZN(n9333) );
  NAND2_X1 U10507 ( .A1(n9908), .A2(n9331), .ZN(n9332) );
  NAND4_X1 U10508 ( .A1(n9335), .A2(n9334), .A3(n9333), .A4(n9332), .ZN(
        P1_U3289) );
  AOI22_X1 U10509 ( .A1(n9337), .A2(n9395), .B1(n9745), .B2(n9336), .ZN(n9338)
         );
  OAI211_X1 U10510 ( .C1(n9340), .C2(n9945), .A(n9339), .B(n9338), .ZN(n9415)
         );
  MUX2_X1 U10511 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9415), .S(n9990), .Z(
        P1_U3551) );
  AOI22_X1 U10512 ( .A1(n9342), .A2(n9395), .B1(n9745), .B2(n9341), .ZN(n9343)
         );
  OAI211_X1 U10513 ( .C1(n9345), .C2(n9945), .A(n9344), .B(n9343), .ZN(n9416)
         );
  MUX2_X1 U10514 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9416), .S(n9990), .Z(
        P1_U3550) );
  AOI22_X1 U10515 ( .A1(n9347), .A2(n9395), .B1(n9745), .B2(n9346), .ZN(n9348)
         );
  OAI211_X1 U10516 ( .C1(n9350), .C2(n9945), .A(n9349), .B(n9348), .ZN(n9417)
         );
  MUX2_X1 U10517 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9417), .S(n9990), .Z(
        P1_U3549) );
  AOI22_X1 U10518 ( .A1(n9352), .A2(n9395), .B1(n9745), .B2(n9351), .ZN(n9353)
         );
  OAI211_X1 U10519 ( .C1(n9355), .C2(n9945), .A(n9354), .B(n9353), .ZN(n9418)
         );
  MUX2_X1 U10520 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9418), .S(n9990), .Z(
        P1_U3548) );
  AOI21_X1 U10521 ( .B1(n9745), .B2(n9357), .A(n9356), .ZN(n9358) );
  OAI211_X1 U10522 ( .C1(n9360), .C2(n9945), .A(n9359), .B(n9358), .ZN(n9419)
         );
  MUX2_X1 U10523 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9419), .S(n9990), .Z(
        P1_U3547) );
  AOI211_X1 U10524 ( .C1(n9745), .C2(n9363), .A(n9362), .B(n9361), .ZN(n9364)
         );
  OAI21_X1 U10525 ( .B1(n9365), .B2(n9945), .A(n9364), .ZN(n9420) );
  MUX2_X1 U10526 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9420), .S(n9990), .Z(
        P1_U3546) );
  AOI22_X1 U10527 ( .A1(n9367), .A2(n9395), .B1(n9745), .B2(n9366), .ZN(n9368)
         );
  OAI211_X1 U10528 ( .C1(n9370), .C2(n9945), .A(n9369), .B(n9368), .ZN(n9421)
         );
  MUX2_X1 U10529 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9421), .S(n9990), .Z(
        P1_U3545) );
  INV_X1 U10530 ( .A(n9945), .ZN(n9969) );
  NAND2_X1 U10531 ( .A1(n9371), .A2(n9969), .ZN(n9378) );
  NAND2_X1 U10532 ( .A1(n9372), .A2(n9745), .ZN(n9373) );
  NAND2_X1 U10533 ( .A1(n9374), .A2(n9373), .ZN(n9375) );
  NOR2_X1 U10534 ( .A1(n9376), .A2(n9375), .ZN(n9377) );
  NAND2_X1 U10535 ( .A1(n9378), .A2(n9377), .ZN(n9422) );
  MUX2_X1 U10536 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9422), .S(n9990), .Z(
        P1_U3544) );
  AOI22_X1 U10537 ( .A1(n9380), .A2(n9395), .B1(n9745), .B2(n9379), .ZN(n9381)
         );
  OAI211_X1 U10538 ( .C1(n9383), .C2(n9945), .A(n9382), .B(n9381), .ZN(n9423)
         );
  MUX2_X1 U10539 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9423), .S(n9990), .Z(
        P1_U3543) );
  AOI22_X1 U10540 ( .A1(n9385), .A2(n9395), .B1(n9745), .B2(n9384), .ZN(n9386)
         );
  OAI211_X1 U10541 ( .C1(n9388), .C2(n9945), .A(n9387), .B(n9386), .ZN(n9424)
         );
  MUX2_X1 U10542 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9424), .S(n9990), .Z(
        P1_U3542) );
  AOI22_X1 U10543 ( .A1(n9390), .A2(n9395), .B1(n9745), .B2(n9389), .ZN(n9391)
         );
  OAI211_X1 U10544 ( .C1(n9393), .C2(n9945), .A(n9392), .B(n9391), .ZN(n9425)
         );
  MUX2_X1 U10545 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9425), .S(n9990), .Z(
        P1_U3541) );
  AOI22_X1 U10546 ( .A1(n9396), .A2(n9395), .B1(n9745), .B2(n9394), .ZN(n9397)
         );
  OAI211_X1 U10547 ( .C1(n9399), .C2(n9945), .A(n9398), .B(n9397), .ZN(n9426)
         );
  MUX2_X1 U10548 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9426), .S(n9990), .Z(
        P1_U3540) );
  AOI21_X1 U10549 ( .B1(n9745), .B2(n9401), .A(n9400), .ZN(n9402) );
  OAI211_X1 U10550 ( .C1(n9404), .C2(n9945), .A(n9403), .B(n9402), .ZN(n9427)
         );
  MUX2_X1 U10551 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9427), .S(n9990), .Z(
        P1_U3539) );
  AOI211_X1 U10552 ( .C1(n9745), .C2(n9407), .A(n9406), .B(n9405), .ZN(n9408)
         );
  OAI21_X1 U10553 ( .B1(n9409), .B2(n9945), .A(n9408), .ZN(n9428) );
  MUX2_X1 U10554 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9428), .S(n9990), .Z(
        P1_U3537) );
  AOI21_X1 U10555 ( .B1(n9745), .B2(n9411), .A(n9410), .ZN(n9412) );
  OAI211_X1 U10556 ( .C1(n9414), .C2(n9945), .A(n9413), .B(n9412), .ZN(n9429)
         );
  MUX2_X1 U10557 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9429), .S(n9990), .Z(
        P1_U3535) );
  MUX2_X1 U10558 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9415), .S(n9980), .Z(
        P1_U3519) );
  MUX2_X1 U10559 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9416), .S(n9980), .Z(
        P1_U3518) );
  MUX2_X1 U10560 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9417), .S(n9980), .Z(
        P1_U3517) );
  MUX2_X1 U10561 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9418), .S(n9980), .Z(
        P1_U3516) );
  MUX2_X1 U10562 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9419), .S(n9980), .Z(
        P1_U3515) );
  MUX2_X1 U10563 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9420), .S(n9980), .Z(
        P1_U3514) );
  MUX2_X1 U10564 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9421), .S(n9980), .Z(
        P1_U3513) );
  MUX2_X1 U10565 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9422), .S(n9980), .Z(
        P1_U3512) );
  MUX2_X1 U10566 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9423), .S(n9980), .Z(
        P1_U3511) );
  MUX2_X1 U10567 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9424), .S(n9980), .Z(
        P1_U3510) );
  MUX2_X1 U10568 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9425), .S(n9980), .Z(
        P1_U3508) );
  MUX2_X1 U10569 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9426), .S(n9980), .Z(
        P1_U3505) );
  MUX2_X1 U10570 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9427), .S(n9980), .Z(
        P1_U3502) );
  MUX2_X1 U10571 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9428), .S(n9980), .Z(
        P1_U3496) );
  MUX2_X1 U10572 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n9429), .S(n9980), .Z(
        P1_U3490) );
  MUX2_X1 U10573 ( .A(n9432), .B(P1_D_REG_0__SCAN_IN), .S(n9933), .Z(P1_U3440)
         );
  INV_X1 U10574 ( .A(n9433), .ZN(n9434) );
  NOR4_X1 U10575 ( .A1(n9434), .A2(P1_IR_REG_30__SCAN_IN), .A3(n10130), .A4(
        n5586), .ZN(n9435) );
  AOI21_X1 U10576 ( .B1(n9441), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9435), .ZN(
        n9436) );
  OAI21_X1 U10577 ( .B1(n9437), .B2(n9443), .A(n9436), .ZN(P1_U3322) );
  AOI21_X1 U10578 ( .B1(n9441), .B2(P2_DATAO_REG_28__SCAN_IN), .A(n9776), .ZN(
        n9438) );
  OAI21_X1 U10579 ( .B1(n9439), .B2(n9443), .A(n9438), .ZN(P1_U3325) );
  AOI21_X1 U10580 ( .B1(n9441), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n9440), .ZN(
        n9442) );
  OAI21_X1 U10581 ( .B1(n9444), .B2(n9443), .A(n9442), .ZN(P1_U3326) );
  INV_X1 U10582 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10118) );
  NOR2_X1 U10583 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9445) );
  AOI21_X1 U10584 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9445), .ZN(n10088) );
  NOR2_X1 U10585 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9446) );
  AOI21_X1 U10586 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9446), .ZN(n10091) );
  NOR2_X1 U10587 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9447) );
  AOI21_X1 U10588 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9447), .ZN(n10094) );
  NOR2_X1 U10589 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9448) );
  AOI21_X1 U10590 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9448), .ZN(n10097) );
  NOR2_X1 U10591 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9449) );
  AOI21_X1 U10592 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9449), .ZN(n10100) );
  INV_X1 U10593 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9856) );
  NOR2_X1 U10594 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9455) );
  XOR2_X1 U10595 ( .A(n9842), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n10128) );
  NAND2_X1 U10596 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9453) );
  XOR2_X1 U10597 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10126) );
  NAND2_X1 U10598 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9451) );
  INV_X1 U10599 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9824) );
  XNOR2_X1 U10600 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n9824), .ZN(n10114) );
  AOI21_X1 U10601 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10081) );
  NAND3_X1 U10602 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10083) );
  OAI21_X1 U10603 ( .B1(n10081), .B2(n10085), .A(n10083), .ZN(n10113) );
  NAND2_X1 U10604 ( .A1(n10114), .A2(n10113), .ZN(n9450) );
  NAND2_X1 U10605 ( .A1(n9451), .A2(n9450), .ZN(n10125) );
  NAND2_X1 U10606 ( .A1(n10126), .A2(n10125), .ZN(n9452) );
  NAND2_X1 U10607 ( .A1(n9453), .A2(n9452), .ZN(n10127) );
  NOR2_X1 U10608 ( .A1(n10128), .A2(n10127), .ZN(n9454) );
  NOR2_X1 U10609 ( .A1(n9455), .A2(n9454), .ZN(n10123) );
  NAND2_X1 U10610 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10123), .ZN(n9456) );
  NOR2_X1 U10611 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10123), .ZN(n10122) );
  AOI21_X1 U10612 ( .B1(n9856), .B2(n9456), .A(n10122), .ZN(n9457) );
  NAND2_X1 U10613 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n9457), .ZN(n9459) );
  XOR2_X1 U10614 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n9457), .Z(n10121) );
  NAND2_X1 U10615 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10121), .ZN(n9458) );
  NAND2_X1 U10616 ( .A1(n9459), .A2(n9458), .ZN(n9460) );
  NAND2_X1 U10617 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9460), .ZN(n9462) );
  XOR2_X1 U10618 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9460), .Z(n10120) );
  NAND2_X1 U10619 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10120), .ZN(n9461) );
  NAND2_X1 U10620 ( .A1(n9462), .A2(n9461), .ZN(n9463) );
  NAND2_X1 U10621 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9463), .ZN(n9465) );
  XOR2_X1 U10622 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n9463), .Z(n10115) );
  NAND2_X1 U10623 ( .A1(n10115), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n9464) );
  NAND2_X1 U10624 ( .A1(n9465), .A2(n9464), .ZN(n9466) );
  AND2_X1 U10625 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9466), .ZN(n9467) );
  XNOR2_X1 U10626 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n9466), .ZN(n10112) );
  INV_X1 U10627 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10111) );
  NOR2_X1 U10628 ( .A1(n10112), .A2(n10111), .ZN(n10110) );
  NOR2_X1 U10629 ( .A1(n9467), .A2(n10110), .ZN(n10109) );
  NAND2_X1 U10630 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9468) );
  OAI21_X1 U10631 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9468), .ZN(n10108) );
  NOR2_X1 U10632 ( .A1(n10109), .A2(n10108), .ZN(n10107) );
  AOI21_X1 U10633 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10107), .ZN(n10106) );
  NAND2_X1 U10634 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9469) );
  OAI21_X1 U10635 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9469), .ZN(n10105) );
  NOR2_X1 U10636 ( .A1(n10106), .A2(n10105), .ZN(n10104) );
  AOI21_X1 U10637 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10104), .ZN(n10103) );
  NOR2_X1 U10638 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9470) );
  AOI21_X1 U10639 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9470), .ZN(n10102) );
  NAND2_X1 U10640 ( .A1(n10103), .A2(n10102), .ZN(n10101) );
  OAI21_X1 U10641 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10101), .ZN(n10099) );
  NAND2_X1 U10642 ( .A1(n10100), .A2(n10099), .ZN(n10098) );
  OAI21_X1 U10643 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10098), .ZN(n10096) );
  NAND2_X1 U10644 ( .A1(n10097), .A2(n10096), .ZN(n10095) );
  OAI21_X1 U10645 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10095), .ZN(n10093) );
  NAND2_X1 U10646 ( .A1(n10094), .A2(n10093), .ZN(n10092) );
  OAI21_X1 U10647 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10092), .ZN(n10090) );
  NAND2_X1 U10648 ( .A1(n10091), .A2(n10090), .ZN(n10089) );
  OAI21_X1 U10649 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10089), .ZN(n10087) );
  NAND2_X1 U10650 ( .A1(n10088), .A2(n10087), .ZN(n10086) );
  NOR2_X1 U10651 ( .A1(n10118), .A2(n10117), .ZN(n9471) );
  NAND2_X1 U10652 ( .A1(n10118), .A2(n10117), .ZN(n10116) );
  OAI21_X1 U10653 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n9471), .A(n10116), .ZN(
        n9654) );
  INV_X1 U10654 ( .A(SI_11_), .ZN(n9652) );
  AOI22_X1 U10655 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_f54), .B1(SI_21_), .B2(keyinput_f11), .ZN(n9472) );
  OAI221_X1 U10656 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_f54), .C1(
        SI_21_), .C2(keyinput_f11), .A(n9472), .ZN(n9479) );
  AOI22_X1 U10657 ( .A1(P2_STATE_REG_SCAN_IN), .A2(keyinput_f34), .B1(SI_17_), 
        .B2(keyinput_f15), .ZN(n9473) );
  OAI221_X1 U10658 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_f34), .C1(SI_17_), 
        .C2(keyinput_f15), .A(n9473), .ZN(n9478) );
  AOI22_X1 U10659 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput_f53), .B1(
        P2_REG3_REG_20__SCAN_IN), .B2(keyinput_f55), .ZN(n9474) );
  OAI221_X1 U10660 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_f53), .C1(
        P2_REG3_REG_20__SCAN_IN), .C2(keyinput_f55), .A(n9474), .ZN(n9477) );
  AOI22_X1 U10661 ( .A1(SI_1_), .A2(keyinput_f31), .B1(SI_8_), .B2(
        keyinput_f24), .ZN(n9475) );
  OAI221_X1 U10662 ( .B1(SI_1_), .B2(keyinput_f31), .C1(SI_8_), .C2(
        keyinput_f24), .A(n9475), .ZN(n9476) );
  NOR4_X1 U10663 ( .A1(n9479), .A2(n9478), .A3(n9477), .A4(n9476), .ZN(n9506)
         );
  XOR2_X1 U10664 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput_f37), .Z(n9486) );
  AOI22_X1 U10665 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(keyinput_f52), .B1(SI_23_), .B2(keyinput_f9), .ZN(n9480) );
  OAI221_X1 U10666 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput_f52), .C1(
        SI_23_), .C2(keyinput_f9), .A(n9480), .ZN(n9485) );
  AOI22_X1 U10667 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput_f41), .B1(
        P2_REG3_REG_21__SCAN_IN), .B2(keyinput_f45), .ZN(n9481) );
  OAI221_X1 U10668 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_f41), .C1(
        P2_REG3_REG_21__SCAN_IN), .C2(keyinput_f45), .A(n9481), .ZN(n9484) );
  AOI22_X1 U10669 ( .A1(SI_4_), .A2(keyinput_f28), .B1(SI_6_), .B2(
        keyinput_f26), .ZN(n9482) );
  OAI221_X1 U10670 ( .B1(SI_4_), .B2(keyinput_f28), .C1(SI_6_), .C2(
        keyinput_f26), .A(n9482), .ZN(n9483) );
  NOR4_X1 U10671 ( .A1(n9486), .A2(n9485), .A3(n9484), .A4(n9483), .ZN(n9505)
         );
  AOI22_X1 U10672 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput_f47), .B1(
        SI_19_), .B2(keyinput_f13), .ZN(n9487) );
  OAI221_X1 U10673 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_f47), .C1(
        SI_19_), .C2(keyinput_f13), .A(n9487), .ZN(n9494) );
  AOI22_X1 U10674 ( .A1(SI_28_), .A2(keyinput_f4), .B1(SI_12_), .B2(
        keyinput_f20), .ZN(n9488) );
  OAI221_X1 U10675 ( .B1(SI_28_), .B2(keyinput_f4), .C1(SI_12_), .C2(
        keyinput_f20), .A(n9488), .ZN(n9493) );
  AOI22_X1 U10676 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput_f51), .B1(
        SI_25_), .B2(keyinput_f7), .ZN(n9489) );
  OAI221_X1 U10677 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .C1(
        SI_25_), .C2(keyinput_f7), .A(n9489), .ZN(n9492) );
  AOI22_X1 U10678 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput_f50), .B1(
        SI_24_), .B2(keyinput_f8), .ZN(n9490) );
  OAI221_X1 U10679 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput_f50), .C1(
        SI_24_), .C2(keyinput_f8), .A(n9490), .ZN(n9491) );
  NOR4_X1 U10680 ( .A1(n9494), .A2(n9493), .A3(n9492), .A4(n9491), .ZN(n9504)
         );
  AOI22_X1 U10681 ( .A1(SI_31_), .A2(keyinput_f1), .B1(SI_22_), .B2(
        keyinput_f10), .ZN(n9495) );
  OAI221_X1 U10682 ( .B1(SI_31_), .B2(keyinput_f1), .C1(SI_22_), .C2(
        keyinput_f10), .A(n9495), .ZN(n9502) );
  AOI22_X1 U10683 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_f59), .B1(SI_10_), .B2(keyinput_f22), .ZN(n9496) );
  OAI221_X1 U10684 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_f59), .C1(
        SI_10_), .C2(keyinput_f22), .A(n9496), .ZN(n9501) );
  AOI22_X1 U10685 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_f49), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .ZN(n9497) );
  OAI221_X1 U10686 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_f49), .C1(
        P2_REG3_REG_18__SCAN_IN), .C2(keyinput_f60), .A(n9497), .ZN(n9500) );
  AOI22_X1 U10687 ( .A1(SI_29_), .A2(keyinput_f3), .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .ZN(n9498) );
  OAI221_X1 U10688 ( .B1(SI_29_), .B2(keyinput_f3), .C1(
        P2_REG3_REG_12__SCAN_IN), .C2(keyinput_f46), .A(n9498), .ZN(n9499) );
  NOR4_X1 U10689 ( .A1(n9502), .A2(n9501), .A3(n9500), .A4(n9499), .ZN(n9503)
         );
  NAND4_X1 U10690 ( .A1(n9506), .A2(n9505), .A3(n9504), .A4(n9503), .ZN(n9555)
         );
  INV_X1 U10691 ( .A(SI_18_), .ZN(n9603) );
  AOI22_X1 U10692 ( .A1(n5117), .A2(keyinput_f35), .B1(n9603), .B2(
        keyinput_f14), .ZN(n9507) );
  OAI221_X1 U10693 ( .B1(n5117), .B2(keyinput_f35), .C1(n9603), .C2(
        keyinput_f14), .A(n9507), .ZN(n9515) );
  INV_X1 U10694 ( .A(SI_5_), .ZN(n9574) );
  AOI22_X1 U10695 ( .A1(n9561), .A2(keyinput_f38), .B1(n9574), .B2(
        keyinput_f27), .ZN(n9508) );
  OAI221_X1 U10696 ( .B1(n9561), .B2(keyinput_f38), .C1(n9574), .C2(
        keyinput_f27), .A(n9508), .ZN(n9514) );
  XNOR2_X1 U10697 ( .A(SI_13_), .B(keyinput_f19), .ZN(n9512) );
  XNOR2_X1 U10698 ( .A(SI_0_), .B(keyinput_f32), .ZN(n9511) );
  XNOR2_X1 U10699 ( .A(SI_3_), .B(keyinput_f29), .ZN(n9510) );
  XNOR2_X1 U10700 ( .A(keyinput_f44), .B(P2_REG3_REG_1__SCAN_IN), .ZN(n9509)
         );
  NAND4_X1 U10701 ( .A1(n9512), .A2(n9511), .A3(n9510), .A4(n9509), .ZN(n9513)
         );
  NOR3_X1 U10702 ( .A1(n9515), .A2(n9514), .A3(n9513), .ZN(n9553) );
  AOI22_X1 U10703 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(keyinput_f48), .B1(n5047), .B2(keyinput_f40), .ZN(n9516) );
  OAI221_X1 U10704 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput_f48), .C1(
        n5047), .C2(keyinput_f40), .A(n9516), .ZN(n9527) );
  AOI22_X1 U10705 ( .A1(n7803), .A2(keyinput_f56), .B1(n9518), .B2(keyinput_f5), .ZN(n9517) );
  OAI221_X1 U10706 ( .B1(n7803), .B2(keyinput_f56), .C1(n9518), .C2(
        keyinput_f5), .A(n9517), .ZN(n9526) );
  INV_X1 U10707 ( .A(SI_15_), .ZN(n9521) );
  AOI22_X1 U10708 ( .A1(n9521), .A2(keyinput_f17), .B1(keyinput_f23), .B2(
        n9520), .ZN(n9519) );
  OAI221_X1 U10709 ( .B1(n9521), .B2(keyinput_f17), .C1(n9520), .C2(
        keyinput_f23), .A(n9519), .ZN(n9525) );
  XOR2_X1 U10710 ( .A(n5521), .B(keyinput_f42), .Z(n9523) );
  XNOR2_X1 U10711 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_f33), .ZN(n9522) );
  NAND2_X1 U10712 ( .A1(n9523), .A2(n9522), .ZN(n9524) );
  NOR4_X1 U10713 ( .A1(n9527), .A2(n9526), .A3(n9525), .A4(n9524), .ZN(n9552)
         );
  AOI22_X1 U10714 ( .A1(n5187), .A2(keyinput_f58), .B1(n9529), .B2(
        keyinput_f12), .ZN(n9528) );
  OAI221_X1 U10715 ( .B1(n5187), .B2(keyinput_f58), .C1(n9529), .C2(
        keyinput_f12), .A(n9528), .ZN(n9537) );
  AOI22_X1 U10716 ( .A1(n9573), .A2(keyinput_f43), .B1(n9577), .B2(
        keyinput_f16), .ZN(n9530) );
  OAI221_X1 U10717 ( .B1(n9573), .B2(keyinput_f43), .C1(n9577), .C2(
        keyinput_f16), .A(n9530), .ZN(n9536) );
  AOI22_X1 U10718 ( .A1(n9586), .A2(keyinput_f39), .B1(n7661), .B2(
        keyinput_f63), .ZN(n9531) );
  OAI221_X1 U10719 ( .B1(n9586), .B2(keyinput_f39), .C1(n7661), .C2(
        keyinput_f63), .A(n9531), .ZN(n9535) );
  AOI22_X1 U10720 ( .A1(n9533), .A2(keyinput_f36), .B1(keyinput_f61), .B2(
        n9558), .ZN(n9532) );
  OAI221_X1 U10721 ( .B1(n9533), .B2(keyinput_f36), .C1(n9558), .C2(
        keyinput_f61), .A(n9532), .ZN(n9534) );
  NOR4_X1 U10722 ( .A1(n9537), .A2(n9536), .A3(n9535), .A4(n9534), .ZN(n9551)
         );
  INV_X1 U10723 ( .A(P2_WR_REG_SCAN_IN), .ZN(n9774) );
  AOI22_X1 U10724 ( .A1(n9539), .A2(keyinput_f62), .B1(keyinput_f0), .B2(n9774), .ZN(n9538) );
  OAI221_X1 U10725 ( .B1(n9539), .B2(keyinput_f62), .C1(n9774), .C2(
        keyinput_f0), .A(n9538), .ZN(n9549) );
  INV_X1 U10726 ( .A(SI_26_), .ZN(n9601) );
  AOI22_X1 U10727 ( .A1(n9541), .A2(keyinput_f57), .B1(n9601), .B2(keyinput_f6), .ZN(n9540) );
  OAI221_X1 U10728 ( .B1(n9541), .B2(keyinput_f57), .C1(n9601), .C2(
        keyinput_f6), .A(n9540), .ZN(n9548) );
  INV_X1 U10729 ( .A(SI_7_), .ZN(n9543) );
  AOI22_X1 U10730 ( .A1(n9543), .A2(keyinput_f25), .B1(keyinput_f2), .B2(n9595), .ZN(n9542) );
  OAI221_X1 U10731 ( .B1(n9543), .B2(keyinput_f25), .C1(n9595), .C2(
        keyinput_f2), .A(n9542), .ZN(n9547) );
  XNOR2_X1 U10732 ( .A(SI_2_), .B(keyinput_f30), .ZN(n9545) );
  XNOR2_X1 U10733 ( .A(SI_14_), .B(keyinput_f18), .ZN(n9544) );
  NAND2_X1 U10734 ( .A1(n9545), .A2(n9544), .ZN(n9546) );
  NOR4_X1 U10735 ( .A1(n9549), .A2(n9548), .A3(n9547), .A4(n9546), .ZN(n9550)
         );
  NAND4_X1 U10736 ( .A1(n9553), .A2(n9552), .A3(n9551), .A4(n9550), .ZN(n9554)
         );
  OAI22_X1 U10737 ( .A1(keyinput_f21), .A2(n9652), .B1(n9555), .B2(n9554), 
        .ZN(n9556) );
  AOI21_X1 U10738 ( .B1(keyinput_f21), .B2(n9652), .A(n9556), .ZN(n9651) );
  AOI22_X1 U10739 ( .A1(n9559), .A2(keyinput_g11), .B1(keyinput_g61), .B2(
        n9558), .ZN(n9557) );
  OAI221_X1 U10740 ( .B1(n9559), .B2(keyinput_g11), .C1(n9558), .C2(
        keyinput_g61), .A(n9557), .ZN(n9571) );
  AOI22_X1 U10741 ( .A1(n9562), .A2(keyinput_g19), .B1(keyinput_g38), .B2(
        n9561), .ZN(n9560) );
  OAI221_X1 U10742 ( .B1(n9562), .B2(keyinput_g19), .C1(n9561), .C2(
        keyinput_g38), .A(n9560), .ZN(n9570) );
  AOI22_X1 U10743 ( .A1(n9565), .A2(keyinput_g51), .B1(keyinput_g45), .B2(
        n9564), .ZN(n9563) );
  OAI221_X1 U10744 ( .B1(n9565), .B2(keyinput_g51), .C1(n9564), .C2(
        keyinput_g45), .A(n9563), .ZN(n9569) );
  AOI22_X1 U10745 ( .A1(n9567), .A2(keyinput_g44), .B1(keyinput_g54), .B2(
        n10024), .ZN(n9566) );
  OAI221_X1 U10746 ( .B1(n9567), .B2(keyinput_g44), .C1(n10024), .C2(
        keyinput_g54), .A(n9566), .ZN(n9568) );
  NOR4_X1 U10747 ( .A1(n9571), .A2(n9570), .A3(n9569), .A4(n9568), .ZN(n9612)
         );
  AOI22_X1 U10748 ( .A1(n9574), .A2(keyinput_g27), .B1(keyinput_g43), .B2(
        n9573), .ZN(n9572) );
  OAI221_X1 U10749 ( .B1(n9574), .B2(keyinput_g27), .C1(n9573), .C2(
        keyinput_g43), .A(n9572), .ZN(n9583) );
  AOI22_X1 U10750 ( .A1(SI_22_), .A2(keyinput_g10), .B1(SI_23_), .B2(
        keyinput_g9), .ZN(n9575) );
  OAI221_X1 U10751 ( .B1(SI_22_), .B2(keyinput_g10), .C1(SI_23_), .C2(
        keyinput_g9), .A(n9575), .ZN(n9582) );
  AOI22_X1 U10752 ( .A1(n5117), .A2(keyinput_g35), .B1(n9577), .B2(
        keyinput_g16), .ZN(n9576) );
  OAI221_X1 U10753 ( .B1(n5117), .B2(keyinput_g35), .C1(n9577), .C2(
        keyinput_g16), .A(n9576), .ZN(n9581) );
  AOI22_X1 U10754 ( .A1(n7803), .A2(keyinput_g56), .B1(n9579), .B2(
        keyinput_g22), .ZN(n9578) );
  OAI221_X1 U10755 ( .B1(n7803), .B2(keyinput_g56), .C1(n9579), .C2(
        keyinput_g22), .A(n9578), .ZN(n9580) );
  NOR4_X1 U10756 ( .A1(n9583), .A2(n9582), .A3(n9581), .A4(n9580), .ZN(n9611)
         );
  AOI22_X1 U10757 ( .A1(n8437), .A2(keyinput_g47), .B1(keyinput_g53), .B2(
        n5151), .ZN(n9584) );
  OAI221_X1 U10758 ( .B1(n8437), .B2(keyinput_g47), .C1(n5151), .C2(
        keyinput_g53), .A(n9584), .ZN(n9593) );
  AOI22_X1 U10759 ( .A1(n9586), .A2(keyinput_g39), .B1(P2_U3152), .B2(
        keyinput_g34), .ZN(n9585) );
  OAI221_X1 U10760 ( .B1(n9586), .B2(keyinput_g39), .C1(P2_U3152), .C2(
        keyinput_g34), .A(n9585), .ZN(n9592) );
  XNOR2_X1 U10761 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_g33), .ZN(n9590) );
  XNOR2_X1 U10762 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_g60), .ZN(n9589)
         );
  XNOR2_X1 U10763 ( .A(SI_1_), .B(keyinput_g31), .ZN(n9588) );
  XNOR2_X1 U10764 ( .A(SI_31_), .B(keyinput_g1), .ZN(n9587) );
  NAND4_X1 U10765 ( .A1(n9590), .A2(n9589), .A3(n9588), .A4(n9587), .ZN(n9591)
         );
  NOR3_X1 U10766 ( .A1(n9593), .A2(n9592), .A3(n9591), .ZN(n9610) );
  AOI22_X1 U10767 ( .A1(n9596), .A2(keyinput_g46), .B1(keyinput_g2), .B2(n9595), .ZN(n9594) );
  OAI221_X1 U10768 ( .B1(n9596), .B2(keyinput_g46), .C1(n9595), .C2(
        keyinput_g2), .A(n9594), .ZN(n9608) );
  AOI22_X1 U10769 ( .A1(n5521), .A2(keyinput_g42), .B1(n9598), .B2(keyinput_g8), .ZN(n9597) );
  OAI221_X1 U10770 ( .B1(n5521), .B2(keyinput_g42), .C1(n9598), .C2(
        keyinput_g8), .A(n9597), .ZN(n9607) );
  AOI22_X1 U10771 ( .A1(n9601), .A2(keyinput_g6), .B1(keyinput_g18), .B2(n9600), .ZN(n9599) );
  OAI221_X1 U10772 ( .B1(n9601), .B2(keyinput_g6), .C1(n9600), .C2(
        keyinput_g18), .A(n9599), .ZN(n9606) );
  AOI22_X1 U10773 ( .A1(n9604), .A2(keyinput_g50), .B1(n9603), .B2(
        keyinput_g14), .ZN(n9602) );
  OAI221_X1 U10774 ( .B1(n9604), .B2(keyinput_g50), .C1(n9603), .C2(
        keyinput_g14), .A(n9602), .ZN(n9605) );
  NOR4_X1 U10775 ( .A1(n9608), .A2(n9607), .A3(n9606), .A4(n9605), .ZN(n9609)
         );
  NAND4_X1 U10776 ( .A1(n9612), .A2(n9611), .A3(n9610), .A4(n9609), .ZN(n9649)
         );
  AOI22_X1 U10777 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(keyinput_g48), .B1(
        P2_REG3_REG_20__SCAN_IN), .B2(keyinput_g55), .ZN(n9613) );
  OAI221_X1 U10778 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput_g48), .C1(
        P2_REG3_REG_20__SCAN_IN), .C2(keyinput_g55), .A(n9613), .ZN(n9620) );
  AOI22_X1 U10779 ( .A1(SI_0_), .A2(keyinput_g32), .B1(SI_2_), .B2(
        keyinput_g30), .ZN(n9614) );
  OAI221_X1 U10780 ( .B1(SI_0_), .B2(keyinput_g32), .C1(SI_2_), .C2(
        keyinput_g30), .A(n9614), .ZN(n9619) );
  AOI22_X1 U10781 ( .A1(SI_29_), .A2(keyinput_g3), .B1(SI_6_), .B2(
        keyinput_g26), .ZN(n9615) );
  OAI221_X1 U10782 ( .B1(SI_29_), .B2(keyinput_g3), .C1(SI_6_), .C2(
        keyinput_g26), .A(n9615), .ZN(n9618) );
  AOI22_X1 U10783 ( .A1(SI_4_), .A2(keyinput_g28), .B1(SI_27_), .B2(
        keyinput_g5), .ZN(n9616) );
  OAI221_X1 U10784 ( .B1(SI_4_), .B2(keyinput_g28), .C1(SI_27_), .C2(
        keyinput_g5), .A(n9616), .ZN(n9617) );
  NOR4_X1 U10785 ( .A1(n9620), .A2(n9619), .A3(n9618), .A4(n9617), .ZN(n9647)
         );
  XOR2_X1 U10786 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput_g37), .Z(n9627) );
  AOI22_X1 U10787 ( .A1(SI_7_), .A2(keyinput_g25), .B1(SI_20_), .B2(
        keyinput_g12), .ZN(n9621) );
  OAI221_X1 U10788 ( .B1(SI_7_), .B2(keyinput_g25), .C1(SI_20_), .C2(
        keyinput_g12), .A(n9621), .ZN(n9626) );
  AOI22_X1 U10789 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput_g41), .B1(
        P2_REG3_REG_26__SCAN_IN), .B2(keyinput_g62), .ZN(n9622) );
  OAI221_X1 U10790 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .C1(
        P2_REG3_REG_26__SCAN_IN), .C2(keyinput_g62), .A(n9622), .ZN(n9625) );
  AOI22_X1 U10791 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput_g36), .B1(SI_8_), .B2(keyinput_g24), .ZN(n9623) );
  OAI221_X1 U10792 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput_g36), .C1(
        SI_8_), .C2(keyinput_g24), .A(n9623), .ZN(n9624) );
  NOR4_X1 U10793 ( .A1(n9627), .A2(n9626), .A3(n9625), .A4(n9624), .ZN(n9646)
         );
  AOI22_X1 U10794 ( .A1(SI_12_), .A2(keyinput_g20), .B1(SI_17_), .B2(
        keyinput_g15), .ZN(n9628) );
  OAI221_X1 U10795 ( .B1(SI_12_), .B2(keyinput_g20), .C1(SI_17_), .C2(
        keyinput_g15), .A(n9628), .ZN(n9635) );
  AOI22_X1 U10796 ( .A1(SI_28_), .A2(keyinput_g4), .B1(SI_3_), .B2(
        keyinput_g29), .ZN(n9629) );
  OAI221_X1 U10797 ( .B1(SI_28_), .B2(keyinput_g4), .C1(SI_3_), .C2(
        keyinput_g29), .A(n9629), .ZN(n9634) );
  AOI22_X1 U10798 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_g59), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .ZN(n9630) );
  OAI221_X1 U10799 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .C1(
        P2_REG3_REG_15__SCAN_IN), .C2(keyinput_g63), .A(n9630), .ZN(n9633) );
  AOI22_X1 U10800 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(keyinput_g52), .B1(SI_19_), .B2(keyinput_g13), .ZN(n9631) );
  OAI221_X1 U10801 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput_g52), .C1(
        SI_19_), .C2(keyinput_g13), .A(n9631), .ZN(n9632) );
  NOR4_X1 U10802 ( .A1(n9635), .A2(n9634), .A3(n9633), .A4(n9632), .ZN(n9645)
         );
  AOI22_X1 U10803 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput_g57), .B1(
        SI_25_), .B2(keyinput_g7), .ZN(n9636) );
  OAI221_X1 U10804 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .C1(
        SI_25_), .C2(keyinput_g7), .A(n9636), .ZN(n9643) );
  AOI22_X1 U10805 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_g40), .B1(SI_15_), .B2(keyinput_g17), .ZN(n9637) );
  OAI221_X1 U10806 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_g40), .C1(
        SI_15_), .C2(keyinput_g17), .A(n9637), .ZN(n9642) );
  AOI22_X1 U10807 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_g0), .B1(SI_9_), .B2(
        keyinput_g23), .ZN(n9638) );
  OAI221_X1 U10808 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_g0), .C1(SI_9_), 
        .C2(keyinput_g23), .A(n9638), .ZN(n9641) );
  AOI22_X1 U10809 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_g49), .B1(
        P2_REG3_REG_11__SCAN_IN), .B2(keyinput_g58), .ZN(n9639) );
  OAI221_X1 U10810 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_g49), .C1(
        P2_REG3_REG_11__SCAN_IN), .C2(keyinput_g58), .A(n9639), .ZN(n9640) );
  NOR4_X1 U10811 ( .A1(n9643), .A2(n9642), .A3(n9641), .A4(n9640), .ZN(n9644)
         );
  NAND4_X1 U10812 ( .A1(n9647), .A2(n9646), .A3(n9645), .A4(n9644), .ZN(n9648)
         );
  OAI22_X1 U10813 ( .A1(keyinput_g21), .A2(n9652), .B1(n9649), .B2(n9648), 
        .ZN(n9650) );
  AOI211_X1 U10814 ( .C1(keyinput_g21), .C2(n9652), .A(n9651), .B(n9650), .ZN(
        n9653) );
  XNOR2_X1 U10815 ( .A(n9654), .B(n9653), .ZN(n9658) );
  NOR2_X1 U10816 ( .A1(n9655), .A2(n9656), .ZN(n9657) );
  XOR2_X1 U10817 ( .A(n9658), .B(n9657), .Z(ADD_1071_U4) );
  INV_X1 U10818 ( .A(n9659), .ZN(n9978) );
  INV_X1 U10819 ( .A(n9660), .ZN(n9662) );
  OAI21_X1 U10820 ( .B1(n9662), .B2(n9972), .A(n9661), .ZN(n9663) );
  AOI21_X1 U10821 ( .B1(n9664), .B2(n9978), .A(n9663), .ZN(n9665) );
  AND2_X1 U10822 ( .A1(n9666), .A2(n9665), .ZN(n9668) );
  INV_X1 U10823 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9667) );
  AOI22_X1 U10824 ( .A1(n9980), .A2(n9668), .B1(n9667), .B2(n6341), .ZN(
        P1_U3484) );
  AOI22_X1 U10825 ( .A1(n9990), .A2(n9668), .B1(n5829), .B2(n6336), .ZN(
        P1_U3533) );
  NOR2_X1 U10826 ( .A1(n9669), .A2(n9973), .ZN(n9670) );
  AOI211_X2 U10827 ( .C1(n9745), .C2(n9671), .A(n9743), .B(n9670), .ZN(n9672)
         );
  AOI22_X1 U10828 ( .A1(n9990), .A2(n9672), .B1(n6467), .B2(n6336), .ZN(
        P1_U3554) );
  AOI22_X1 U10829 ( .A1(n9980), .A2(n9672), .B1(n6469), .B2(n6341), .ZN(
        P1_U3522) );
  NOR2_X1 U10830 ( .A1(n9673), .A2(n10064), .ZN(n9674) );
  INV_X1 U10831 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9678) );
  AOI22_X1 U10832 ( .A1(n10080), .A2(n9693), .B1(n9678), .B2(n10078), .ZN(
        P2_U3551) );
  OAI21_X1 U10833 ( .B1(n9680), .B2(n10062), .A(n9679), .ZN(n9681) );
  AOI21_X1 U10834 ( .B1(n9683), .B2(n9682), .A(n9681), .ZN(n9695) );
  INV_X1 U10835 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9684) );
  AOI22_X1 U10836 ( .A1(n10080), .A2(n9695), .B1(n9684), .B2(n10078), .ZN(
        P2_U3550) );
  INV_X1 U10837 ( .A(n9685), .ZN(n10060) );
  OAI22_X1 U10838 ( .A1(n9687), .A2(n10064), .B1(n9686), .B2(n10062), .ZN(
        n9689) );
  AOI211_X1 U10839 ( .C1(n10060), .C2(n9690), .A(n9689), .B(n9688), .ZN(n9697)
         );
  AOI22_X1 U10840 ( .A1(n10080), .A2(n9697), .B1(n9691), .B2(n10078), .ZN(
        P2_U3533) );
  INV_X1 U10841 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9692) );
  AOI22_X1 U10842 ( .A1(n4316), .A2(n9693), .B1(n9692), .B2(n10070), .ZN(
        P2_U3519) );
  INV_X1 U10843 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9694) );
  AOI22_X1 U10844 ( .A1(n4316), .A2(n9695), .B1(n9694), .B2(n10070), .ZN(
        P2_U3518) );
  INV_X1 U10845 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9696) );
  AOI22_X1 U10846 ( .A1(n4316), .A2(n9697), .B1(n9696), .B2(n10070), .ZN(
        P2_U3490) );
  XNOR2_X1 U10847 ( .A(n9698), .B(n9705), .ZN(n9755) );
  NOR2_X1 U10848 ( .A1(n9699), .A2(n9752), .ZN(n9700) );
  OR2_X1 U10849 ( .A1(n9701), .A2(n9700), .ZN(n9753) );
  INV_X1 U10850 ( .A(n9753), .ZN(n9702) );
  AOI22_X1 U10851 ( .A1(n9755), .A2(n9909), .B1(n9908), .B2(n9702), .ZN(n9719)
         );
  OAI22_X1 U10852 ( .A1(n9930), .A2(n9704), .B1(n9703), .B2(n9925), .ZN(n9716)
         );
  INV_X1 U10853 ( .A(n9705), .ZN(n9706) );
  XNOR2_X1 U10854 ( .A(n9707), .B(n9706), .ZN(n9713) );
  AOI22_X1 U10855 ( .A1(n9711), .A2(n9710), .B1(n9709), .B2(n9708), .ZN(n9712)
         );
  OAI21_X1 U10856 ( .B1(n9713), .B2(n9732), .A(n9712), .ZN(n9714) );
  AOI21_X1 U10857 ( .B1(n9755), .B2(n9735), .A(n9714), .ZN(n9757) );
  NOR2_X1 U10858 ( .A1(n9757), .A2(n9736), .ZN(n9715) );
  AOI211_X1 U10859 ( .C1(n9739), .C2(n9717), .A(n9716), .B(n9715), .ZN(n9718)
         );
  NAND2_X1 U10860 ( .A1(n9719), .A2(n9718), .ZN(P1_U3278) );
  XNOR2_X1 U10861 ( .A(n9720), .B(n9727), .ZN(n9762) );
  AND2_X1 U10862 ( .A1(n9721), .A2(n9759), .ZN(n9723) );
  OR2_X1 U10863 ( .A1(n9723), .A2(n9722), .ZN(n9760) );
  INV_X1 U10864 ( .A(n9760), .ZN(n9724) );
  AOI22_X1 U10865 ( .A1(n9762), .A2(n9909), .B1(n9908), .B2(n9724), .ZN(n9741)
         );
  OAI22_X1 U10866 ( .A1(n9930), .A2(n9726), .B1(n9725), .B2(n9925), .ZN(n9738)
         );
  XNOR2_X1 U10867 ( .A(n9728), .B(n9727), .ZN(n9733) );
  OAI22_X1 U10868 ( .A1(n9915), .A2(n9916), .B1(n9729), .B2(n9914), .ZN(n9730)
         );
  INV_X1 U10869 ( .A(n9730), .ZN(n9731) );
  OAI21_X1 U10870 ( .B1(n9733), .B2(n9732), .A(n9731), .ZN(n9734) );
  AOI21_X1 U10871 ( .B1(n9762), .B2(n9735), .A(n9734), .ZN(n9764) );
  NOR2_X1 U10872 ( .A1(n9764), .A2(n9736), .ZN(n9737) );
  AOI211_X1 U10873 ( .C1(n9739), .C2(n9759), .A(n9738), .B(n9737), .ZN(n9740)
         );
  NAND2_X1 U10874 ( .A1(n9741), .A2(n9740), .ZN(P1_U3280) );
  AOI22_X1 U10875 ( .A1(n9990), .A2(n9767), .B1(n6327), .B2(n6336), .ZN(
        P1_U3553) );
  OAI21_X1 U10876 ( .B1(n9747), .B2(n9972), .A(n9746), .ZN(n9748) );
  AOI21_X1 U10877 ( .B1(n9749), .B2(n9978), .A(n9748), .ZN(n9750) );
  AND2_X1 U10878 ( .A1(n9751), .A2(n9750), .ZN(n9769) );
  AOI22_X1 U10879 ( .A1(n9990), .A2(n9769), .B1(n5930), .B2(n6336), .ZN(
        P1_U3538) );
  OAI22_X1 U10880 ( .A1(n9753), .A2(n9973), .B1(n9752), .B2(n9972), .ZN(n9754)
         );
  AOI21_X1 U10881 ( .B1(n9755), .B2(n9978), .A(n9754), .ZN(n9756) );
  AOI22_X1 U10882 ( .A1(n9990), .A2(n9771), .B1(n9758), .B2(n6336), .ZN(
        P1_U3536) );
  OAI22_X1 U10883 ( .A1(n9760), .A2(n9973), .B1(n4639), .B2(n9972), .ZN(n9761)
         );
  AOI21_X1 U10884 ( .B1(n9762), .B2(n9978), .A(n9761), .ZN(n9763) );
  AOI22_X1 U10885 ( .A1(n9990), .A2(n9773), .B1(n9765), .B2(n6336), .ZN(
        P1_U3534) );
  INV_X1 U10886 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9766) );
  AOI22_X1 U10887 ( .A1(n9980), .A2(n9767), .B1(n9766), .B2(n6341), .ZN(
        P1_U3521) );
  INV_X1 U10888 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9768) );
  AOI22_X1 U10889 ( .A1(n9980), .A2(n9769), .B1(n9768), .B2(n6341), .ZN(
        P1_U3499) );
  INV_X1 U10890 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9770) );
  AOI22_X1 U10891 ( .A1(n9980), .A2(n9771), .B1(n9770), .B2(n6341), .ZN(
        P1_U3493) );
  INV_X1 U10892 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9772) );
  AOI22_X1 U10893 ( .A1(n9980), .A2(n9773), .B1(n9772), .B2(n6341), .ZN(
        P1_U3487) );
  XOR2_X1 U10894 ( .A(n9774), .B(P1_WR_REG_SCAN_IN), .Z(U123) );
  INV_X1 U10895 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9784) );
  OR2_X1 U10896 ( .A1(n6323), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9775) );
  NAND2_X1 U10897 ( .A1(n9776), .A2(n9775), .ZN(n9778) );
  NAND2_X1 U10898 ( .A1(n9778), .A2(n9777), .ZN(n9805) );
  INV_X1 U10899 ( .A(n9796), .ZN(n9779) );
  NOR2_X1 U10900 ( .A1(n6241), .A2(n9779), .ZN(n9802) );
  INV_X1 U10901 ( .A(n9802), .ZN(n9781) );
  OAI21_X1 U10902 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(n9786), .A(n6323), .ZN(
        n9780) );
  NAND3_X1 U10903 ( .A1(n9805), .A2(n9781), .A3(n9780), .ZN(n9782) );
  OAI22_X1 U10904 ( .A1(n9899), .A2(n9784), .B1(n9783), .B2(n9782), .ZN(n9785)
         );
  INV_X1 U10905 ( .A(n9785), .ZN(n9788) );
  NAND3_X1 U10906 ( .A1(n9894), .A2(P1_IR_REG_0__SCAN_IN), .A3(n9786), .ZN(
        n9787) );
  OAI211_X1 U10907 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n5637), .A(n9788), .B(
        n9787), .ZN(P1_U3241) );
  NAND2_X1 U10908 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9791) );
  AOI211_X1 U10909 ( .C1(n9791), .C2(n9790), .A(n9789), .B(n9843), .ZN(n9792)
         );
  AOI21_X1 U10910 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n10130), .A(n9792), .ZN(
        n9799) );
  AOI22_X1 U10911 ( .A1(n9880), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(n9793), .B2(
        n9886), .ZN(n9798) );
  OAI211_X1 U10912 ( .C1(n9796), .C2(n9795), .A(n9895), .B(n9794), .ZN(n9797)
         );
  NAND3_X1 U10913 ( .A1(n9799), .A2(n9798), .A3(n9797), .ZN(P1_U3242) );
  NOR2_X1 U10914 ( .A1(n9800), .A2(n6241), .ZN(n9801) );
  MUX2_X1 U10915 ( .A(n9802), .B(n9801), .S(n6323), .Z(n9803) );
  INV_X1 U10916 ( .A(n9803), .ZN(n9807) );
  AND2_X1 U10917 ( .A1(n9805), .A2(n9804), .ZN(n9806) );
  NAND2_X1 U10918 ( .A1(n9807), .A2(n9806), .ZN(n9840) );
  XNOR2_X1 U10919 ( .A(n9809), .B(n9808), .ZN(n9810) );
  NAND2_X1 U10920 ( .A1(n9895), .A2(n9810), .ZN(n9821) );
  NAND2_X1 U10921 ( .A1(n9886), .A2(n9811), .ZN(n9820) );
  NAND2_X1 U10922 ( .A1(P1_U3084), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9819) );
  INV_X1 U10923 ( .A(n9812), .ZN(n9815) );
  INV_X1 U10924 ( .A(n9813), .ZN(n9814) );
  NAND2_X1 U10925 ( .A1(n9815), .A2(n9814), .ZN(n9816) );
  NAND3_X1 U10926 ( .A1(n9894), .A2(n9817), .A3(n9816), .ZN(n9818) );
  AND4_X1 U10927 ( .A1(n9821), .A2(n9820), .A3(n9819), .A4(n9818), .ZN(n9822)
         );
  AND2_X1 U10928 ( .A1(n9840), .A2(n9822), .ZN(n9823) );
  OAI21_X1 U10929 ( .B1(n9899), .B2(n9824), .A(n9823), .ZN(P1_U3243) );
  AND2_X1 U10930 ( .A1(n9826), .A2(n9825), .ZN(n9827) );
  OAI21_X1 U10931 ( .B1(n9828), .B2(n9827), .A(n9895), .ZN(n9839) );
  NAND2_X1 U10932 ( .A1(n9886), .A2(n9830), .ZN(n9838) );
  INV_X1 U10933 ( .A(n9829), .ZN(n9832) );
  MUX2_X1 U10934 ( .A(n6739), .B(P1_REG1_REG_4__SCAN_IN), .S(n9830), .Z(n9831)
         );
  NAND2_X1 U10935 ( .A1(n9832), .A2(n9831), .ZN(n9833) );
  NAND2_X1 U10936 ( .A1(n9834), .A2(n9833), .ZN(n9836) );
  AOI21_X1 U10937 ( .B1(n9894), .B2(n9836), .A(n9835), .ZN(n9837) );
  AND3_X1 U10938 ( .A1(n9839), .A2(n9838), .A3(n9837), .ZN(n9841) );
  OAI211_X1 U10939 ( .C1(n9842), .C2(n9899), .A(n9841), .B(n9840), .ZN(
        P1_U3245) );
  AOI211_X1 U10940 ( .C1(n9846), .C2(n9845), .A(n9844), .B(n9843), .ZN(n9847)
         );
  AOI211_X1 U10941 ( .C1(n9886), .C2(n9849), .A(n9848), .B(n9847), .ZN(n9855)
         );
  AOI21_X1 U10942 ( .B1(n9852), .B2(n9851), .A(n9850), .ZN(n9853) );
  OR2_X1 U10943 ( .A1(n9872), .A2(n9853), .ZN(n9854) );
  OAI211_X1 U10944 ( .C1(n9856), .C2(n9899), .A(n9855), .B(n9854), .ZN(
        P1_U3246) );
  OAI21_X1 U10945 ( .B1(n9859), .B2(n9858), .A(n9857), .ZN(n9865) );
  AOI211_X1 U10946 ( .C1(n9862), .C2(n9861), .A(n9860), .B(n9872), .ZN(n9863)
         );
  AOI211_X1 U10947 ( .C1(n9894), .C2(n9865), .A(n9864), .B(n9863), .ZN(n9868)
         );
  AOI22_X1 U10948 ( .A1(n9880), .A2(P1_ADDR_REG_9__SCAN_IN), .B1(n9866), .B2(
        n9886), .ZN(n9867) );
  NAND2_X1 U10949 ( .A1(n9868), .A2(n9867), .ZN(P1_U3250) );
  OAI21_X1 U10950 ( .B1(n9871), .B2(n9870), .A(n9869), .ZN(n9878) );
  AOI211_X1 U10951 ( .C1(n9875), .C2(n9874), .A(n9873), .B(n9872), .ZN(n9876)
         );
  AOI211_X1 U10952 ( .C1(n9878), .C2(n9894), .A(n9877), .B(n9876), .ZN(n9882)
         );
  AOI22_X1 U10953 ( .A1(n9880), .A2(P1_ADDR_REG_10__SCAN_IN), .B1(n9879), .B2(
        n9886), .ZN(n9881) );
  NAND2_X1 U10954 ( .A1(n9882), .A2(n9881), .ZN(P1_U3251) );
  INV_X1 U10955 ( .A(n9883), .ZN(n9884) );
  AOI21_X1 U10956 ( .B1(n9886), .B2(n9885), .A(n9884), .ZN(n9898) );
  AOI21_X1 U10957 ( .B1(n9889), .B2(n9888), .A(n9887), .ZN(n9896) );
  OAI21_X1 U10958 ( .B1(n9892), .B2(n9891), .A(n9890), .ZN(n9893) );
  AOI22_X1 U10959 ( .A1(n9896), .A2(n9895), .B1(n9894), .B2(n9893), .ZN(n9897)
         );
  OAI211_X1 U10960 ( .C1(n9899), .C2(n10118), .A(n9898), .B(n9897), .ZN(
        P1_U3259) );
  NAND2_X1 U10961 ( .A1(n9901), .A2(n9900), .ZN(n9912) );
  XNOR2_X1 U10962 ( .A(n9902), .B(n9912), .ZN(n9923) );
  INV_X1 U10963 ( .A(n9923), .ZN(n9977) );
  INV_X1 U10964 ( .A(n9903), .ZN(n9906) );
  OAI21_X1 U10965 ( .B1(n9906), .B2(n4759), .A(n9905), .ZN(n9974) );
  INV_X1 U10966 ( .A(n9974), .ZN(n9907) );
  AOI22_X1 U10967 ( .A1(n9977), .A2(n9909), .B1(n9908), .B2(n9907), .ZN(n9932)
         );
  NAND2_X1 U10968 ( .A1(n9911), .A2(n9910), .ZN(n9913) );
  XNOR2_X1 U10969 ( .A(n9913), .B(n9912), .ZN(n9920) );
  OAI22_X1 U10970 ( .A1(n9917), .A2(n9916), .B1(n9915), .B2(n9914), .ZN(n9918)
         );
  AOI21_X1 U10971 ( .B1(n9920), .B2(n9919), .A(n9918), .ZN(n9921) );
  OAI21_X1 U10972 ( .B1(n9923), .B2(n9922), .A(n9921), .ZN(n9975) );
  NOR2_X1 U10973 ( .A1(n9924), .A2(n4759), .ZN(n9929) );
  INV_X1 U10974 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9927) );
  OAI22_X1 U10975 ( .A1(n9930), .A2(n9927), .B1(n9926), .B2(n9925), .ZN(n9928)
         );
  AOI211_X1 U10976 ( .C1(n9975), .C2(n9930), .A(n9929), .B(n9928), .ZN(n9931)
         );
  NAND2_X1 U10977 ( .A1(n9932), .A2(n9931), .ZN(P1_U3282) );
  AND2_X1 U10978 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9933), .ZN(P1_U3292) );
  AND2_X1 U10979 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9933), .ZN(P1_U3293) );
  AND2_X1 U10980 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9933), .ZN(P1_U3294) );
  AND2_X1 U10981 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9933), .ZN(P1_U3295) );
  AND2_X1 U10982 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9933), .ZN(P1_U3296) );
  AND2_X1 U10983 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9933), .ZN(P1_U3297) );
  AND2_X1 U10984 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9933), .ZN(P1_U3298) );
  AND2_X1 U10985 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9933), .ZN(P1_U3299) );
  AND2_X1 U10986 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9933), .ZN(P1_U3300) );
  AND2_X1 U10987 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9933), .ZN(P1_U3301) );
  AND2_X1 U10988 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9933), .ZN(P1_U3302) );
  AND2_X1 U10989 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9933), .ZN(P1_U3303) );
  AND2_X1 U10990 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9933), .ZN(P1_U3304) );
  AND2_X1 U10991 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9933), .ZN(P1_U3305) );
  AND2_X1 U10992 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9933), .ZN(P1_U3306) );
  AND2_X1 U10993 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9933), .ZN(P1_U3307) );
  AND2_X1 U10994 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9933), .ZN(P1_U3308) );
  AND2_X1 U10995 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9933), .ZN(P1_U3309) );
  AND2_X1 U10996 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9933), .ZN(P1_U3310) );
  AND2_X1 U10997 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9933), .ZN(P1_U3311) );
  AND2_X1 U10998 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9933), .ZN(P1_U3312) );
  AND2_X1 U10999 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9933), .ZN(P1_U3313) );
  AND2_X1 U11000 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9933), .ZN(P1_U3314) );
  AND2_X1 U11001 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9933), .ZN(P1_U3315) );
  AND2_X1 U11002 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9933), .ZN(P1_U3316) );
  AND2_X1 U11003 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9933), .ZN(P1_U3317) );
  AND2_X1 U11004 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9933), .ZN(P1_U3318) );
  AND2_X1 U11005 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9933), .ZN(P1_U3319) );
  AND2_X1 U11006 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9933), .ZN(P1_U3320) );
  AND2_X1 U11007 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9933), .ZN(P1_U3321) );
  INV_X1 U11008 ( .A(n9934), .ZN(n9939) );
  OAI21_X1 U11009 ( .B1(n9936), .B2(n9972), .A(n9935), .ZN(n9938) );
  AOI211_X1 U11010 ( .C1(n9939), .C2(n9969), .A(n9938), .B(n9937), .ZN(n9981)
         );
  AOI22_X1 U11011 ( .A1(n9980), .A2(n9981), .B1(n5652), .B2(n6341), .ZN(
        P1_U3457) );
  OAI21_X1 U11012 ( .B1(n9941), .B2(n9972), .A(n9940), .ZN(n9943) );
  AOI211_X1 U11013 ( .C1(n9978), .C2(n9944), .A(n9943), .B(n9942), .ZN(n9982)
         );
  AOI22_X1 U11014 ( .A1(n9980), .A2(n9982), .B1(n5591), .B2(n6341), .ZN(
        P1_U3463) );
  OR2_X1 U11015 ( .A1(n9946), .A2(n9945), .ZN(n9951) );
  INV_X1 U11016 ( .A(n9947), .ZN(n9948) );
  AND2_X1 U11017 ( .A1(n9949), .A2(n9948), .ZN(n9950) );
  AOI22_X1 U11018 ( .A1(n9980), .A2(n9984), .B1(n5719), .B2(n6341), .ZN(
        P1_U3469) );
  INV_X1 U11019 ( .A(n9953), .ZN(n9955) );
  OAI22_X1 U11020 ( .A1(n9955), .A2(n9973), .B1(n9954), .B2(n9972), .ZN(n9957)
         );
  AOI211_X1 U11021 ( .C1(n9978), .C2(n9958), .A(n9957), .B(n9956), .ZN(n9986)
         );
  AOI22_X1 U11022 ( .A1(n9980), .A2(n9986), .B1(n5738), .B2(n6341), .ZN(
        P1_U3472) );
  OAI21_X1 U11023 ( .B1(n9960), .B2(n9972), .A(n9959), .ZN(n9962) );
  AOI211_X1 U11024 ( .C1(n9969), .C2(n9963), .A(n9962), .B(n9961), .ZN(n9987)
         );
  INV_X1 U11025 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9964) );
  AOI22_X1 U11026 ( .A1(n9980), .A2(n9987), .B1(n9964), .B2(n6341), .ZN(
        P1_U3475) );
  OAI21_X1 U11027 ( .B1(n9966), .B2(n9973), .A(n9965), .ZN(n9967) );
  AOI211_X1 U11028 ( .C1(n9970), .C2(n9969), .A(n9968), .B(n9967), .ZN(n9988)
         );
  INV_X1 U11029 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9971) );
  AOI22_X1 U11030 ( .A1(n9980), .A2(n9988), .B1(n9971), .B2(n6341), .ZN(
        P1_U3478) );
  OAI22_X1 U11031 ( .A1(n9974), .A2(n9973), .B1(n4759), .B2(n9972), .ZN(n9976)
         );
  AOI211_X1 U11032 ( .C1(n9978), .C2(n9977), .A(n9976), .B(n9975), .ZN(n9989)
         );
  INV_X1 U11033 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9979) );
  AOI22_X1 U11034 ( .A1(n9980), .A2(n9989), .B1(n9979), .B2(n6341), .ZN(
        P1_U3481) );
  AOI22_X1 U11035 ( .A1(n9990), .A2(n9981), .B1(n5653), .B2(n6336), .ZN(
        P1_U3524) );
  AOI22_X1 U11036 ( .A1(n9990), .A2(n9982), .B1(n6715), .B2(n6336), .ZN(
        P1_U3526) );
  INV_X1 U11037 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9983) );
  AOI22_X1 U11038 ( .A1(n9990), .A2(n9984), .B1(n9983), .B2(n6336), .ZN(
        P1_U3528) );
  INV_X1 U11039 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9985) );
  AOI22_X1 U11040 ( .A1(n9990), .A2(n9986), .B1(n9985), .B2(n6336), .ZN(
        P1_U3529) );
  AOI22_X1 U11041 ( .A1(n9990), .A2(n9987), .B1(n6735), .B2(n6336), .ZN(
        P1_U3530) );
  AOI22_X1 U11042 ( .A1(n9990), .A2(n9988), .B1(n6742), .B2(n6336), .ZN(
        P1_U3531) );
  AOI22_X1 U11043 ( .A1(n9990), .A2(n9989), .B1(n5811), .B2(n6336), .ZN(
        P1_U3532) );
  AOI22_X1 U11044 ( .A1(n9992), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9991), .ZN(n10002) );
  AOI22_X1 U11045 ( .A1(n9994), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10001) );
  OAI21_X1 U11046 ( .B1(P2_REG1_REG_0__SCAN_IN), .B2(n9996), .A(n9995), .ZN(
        n9999) );
  NOR2_X1 U11047 ( .A1(n9997), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9998) );
  OAI21_X1 U11048 ( .B1(n9999), .B2(n9998), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n10000) );
  OAI211_X1 U11049 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n10002), .A(n10001), .B(
        n10000), .ZN(P2_U3245) );
  AOI22_X1 U11050 ( .A1(n10005), .A2(n10014), .B1(n10004), .B2(n10003), .ZN(
        n10006) );
  OAI211_X1 U11051 ( .C1(n9567), .C2(n10025), .A(n10007), .B(n10006), .ZN(
        n10008) );
  AOI22_X1 U11052 ( .A1(n10011), .A2(n10010), .B1(n10009), .B2(n10008), .ZN(
        n10012) );
  OAI21_X1 U11053 ( .B1(n6856), .B2(n10009), .A(n10012), .ZN(P2_U3295) );
  NAND2_X1 U11054 ( .A1(n10014), .A2(n10013), .ZN(n10015) );
  AOI21_X1 U11055 ( .B1(n10016), .B2(n10015), .A(n10022), .ZN(n10021) );
  AOI21_X1 U11056 ( .B1(n10019), .B2(n10018), .A(n10017), .ZN(n10020) );
  AOI211_X1 U11057 ( .C1(n10022), .C2(P2_REG2_REG_0__SCAN_IN), .A(n10021), .B(
        n10020), .ZN(n10023) );
  OAI21_X1 U11058 ( .B1(n10025), .B2(n10024), .A(n10023), .ZN(P2_U3296) );
  AND2_X1 U11059 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10030), .ZN(P2_U3297) );
  AND2_X1 U11060 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10030), .ZN(P2_U3298) );
  AND2_X1 U11061 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10030), .ZN(P2_U3299) );
  AND2_X1 U11062 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10030), .ZN(P2_U3300) );
  AND2_X1 U11063 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10030), .ZN(P2_U3301) );
  AND2_X1 U11064 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10030), .ZN(P2_U3302) );
  AND2_X1 U11065 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10030), .ZN(P2_U3303) );
  AND2_X1 U11066 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10030), .ZN(P2_U3304) );
  AND2_X1 U11067 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10030), .ZN(P2_U3305) );
  AND2_X1 U11068 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10030), .ZN(P2_U3306) );
  AND2_X1 U11069 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10030), .ZN(P2_U3307) );
  AND2_X1 U11070 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10030), .ZN(P2_U3308) );
  AND2_X1 U11071 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10030), .ZN(P2_U3309) );
  AND2_X1 U11072 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10030), .ZN(P2_U3310) );
  AND2_X1 U11073 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10030), .ZN(P2_U3311) );
  AND2_X1 U11074 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10030), .ZN(P2_U3312) );
  AND2_X1 U11075 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10030), .ZN(P2_U3313) );
  AND2_X1 U11076 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10030), .ZN(P2_U3314) );
  AND2_X1 U11077 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10030), .ZN(P2_U3315) );
  AND2_X1 U11078 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10030), .ZN(P2_U3316) );
  AND2_X1 U11079 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10030), .ZN(P2_U3317) );
  AND2_X1 U11080 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10030), .ZN(P2_U3318) );
  AND2_X1 U11081 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10030), .ZN(P2_U3319) );
  AND2_X1 U11082 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10030), .ZN(P2_U3320) );
  AND2_X1 U11083 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10030), .ZN(P2_U3321) );
  AND2_X1 U11084 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10030), .ZN(P2_U3322) );
  AND2_X1 U11085 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10030), .ZN(P2_U3323) );
  AND2_X1 U11086 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10030), .ZN(P2_U3324) );
  AND2_X1 U11087 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10030), .ZN(P2_U3325) );
  AND2_X1 U11088 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10030), .ZN(P2_U3326) );
  AOI22_X1 U11089 ( .A1(n10033), .A2(n10029), .B1(n10028), .B2(n10030), .ZN(
        P2_U3437) );
  AOI22_X1 U11090 ( .A1(n10033), .A2(n10032), .B1(n10031), .B2(n10030), .ZN(
        P2_U3438) );
  INV_X1 U11091 ( .A(n10034), .ZN(n10035) );
  OAI21_X1 U11092 ( .B1(n4425), .B2(n10062), .A(n10035), .ZN(n10036) );
  AOI21_X1 U11093 ( .B1(n10037), .B2(n10060), .A(n10036), .ZN(n10038) );
  AND2_X1 U11094 ( .A1(n10039), .A2(n10038), .ZN(n10073) );
  INV_X1 U11095 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10040) );
  AOI22_X1 U11096 ( .A1(n4316), .A2(n10073), .B1(n10040), .B2(n10070), .ZN(
        P2_U3460) );
  INV_X1 U11097 ( .A(n10041), .ZN(n10042) );
  OAI211_X1 U11098 ( .C1(n10044), .C2(n10062), .A(n10043), .B(n10042), .ZN(
        n10045) );
  AOI21_X1 U11099 ( .B1(n10068), .B2(n10046), .A(n10045), .ZN(n10075) );
  INV_X1 U11100 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10047) );
  AOI22_X1 U11101 ( .A1(n4316), .A2(n10075), .B1(n10047), .B2(n10070), .ZN(
        P2_U3466) );
  OAI22_X1 U11102 ( .A1(n10049), .A2(n10064), .B1(n10048), .B2(n10062), .ZN(
        n10051) );
  AOI211_X1 U11103 ( .C1(n10052), .C2(n10068), .A(n10051), .B(n10050), .ZN(
        n10076) );
  INV_X1 U11104 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10053) );
  AOI22_X1 U11105 ( .A1(n4316), .A2(n10076), .B1(n10053), .B2(n10070), .ZN(
        P2_U3472) );
  INV_X1 U11106 ( .A(n10054), .ZN(n10059) );
  OAI22_X1 U11107 ( .A1(n10056), .A2(n10064), .B1(n10055), .B2(n10062), .ZN(
        n10058) );
  AOI211_X1 U11108 ( .C1(n10060), .C2(n10059), .A(n10058), .B(n10057), .ZN(
        n10077) );
  INV_X1 U11109 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10061) );
  AOI22_X1 U11110 ( .A1(n4316), .A2(n10077), .B1(n10061), .B2(n10070), .ZN(
        P2_U3478) );
  OAI22_X1 U11111 ( .A1(n10065), .A2(n10064), .B1(n10063), .B2(n10062), .ZN(
        n10066) );
  AOI211_X1 U11112 ( .C1(n10069), .C2(n10068), .A(n10067), .B(n10066), .ZN(
        n10079) );
  INV_X1 U11113 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10071) );
  AOI22_X1 U11114 ( .A1(n4316), .A2(n10079), .B1(n10071), .B2(n10070), .ZN(
        P2_U3484) );
  INV_X1 U11115 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10072) );
  AOI22_X1 U11116 ( .A1(n10080), .A2(n10073), .B1(n10072), .B2(n10078), .ZN(
        P2_U3523) );
  INV_X1 U11117 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10074) );
  AOI22_X1 U11118 ( .A1(n10080), .A2(n10075), .B1(n10074), .B2(n10078), .ZN(
        P2_U3525) );
  AOI22_X1 U11119 ( .A1(n10080), .A2(n10076), .B1(n6929), .B2(n10078), .ZN(
        P2_U3527) );
  AOI22_X1 U11120 ( .A1(n10080), .A2(n10077), .B1(n7123), .B2(n10078), .ZN(
        P2_U3529) );
  AOI22_X1 U11121 ( .A1(n10080), .A2(n10079), .B1(n7647), .B2(n10078), .ZN(
        P2_U3531) );
  INV_X1 U11122 ( .A(n10081), .ZN(n10082) );
  NAND2_X1 U11123 ( .A1(n10083), .A2(n10082), .ZN(n10084) );
  XOR2_X1 U11124 ( .A(n10085), .B(n10084), .Z(ADD_1071_U5) );
  XOR2_X1 U11125 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11126 ( .B1(n10088), .B2(n10087), .A(n10086), .ZN(ADD_1071_U56) );
  OAI21_X1 U11127 ( .B1(n10091), .B2(n10090), .A(n10089), .ZN(ADD_1071_U57) );
  OAI21_X1 U11128 ( .B1(n10094), .B2(n10093), .A(n10092), .ZN(ADD_1071_U58) );
  OAI21_X1 U11129 ( .B1(n10097), .B2(n10096), .A(n10095), .ZN(ADD_1071_U59) );
  OAI21_X1 U11130 ( .B1(n10100), .B2(n10099), .A(n10098), .ZN(ADD_1071_U60) );
  OAI21_X1 U11131 ( .B1(n10103), .B2(n10102), .A(n10101), .ZN(ADD_1071_U61) );
  AOI21_X1 U11132 ( .B1(n10106), .B2(n10105), .A(n10104), .ZN(ADD_1071_U62) );
  AOI21_X1 U11133 ( .B1(n10109), .B2(n10108), .A(n10107), .ZN(ADD_1071_U63) );
  AOI21_X1 U11134 ( .B1(n10112), .B2(n10111), .A(n10110), .ZN(ADD_1071_U47) );
  XOR2_X1 U11135 ( .A(n10114), .B(n10113), .Z(ADD_1071_U54) );
  XOR2_X1 U11136 ( .A(n10115), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1071_U48) );
  OAI21_X1 U11137 ( .B1(n10118), .B2(n10117), .A(n10116), .ZN(n10119) );
  XNOR2_X1 U11138 ( .A(n10119), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XOR2_X1 U11139 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10120), .Z(ADD_1071_U49) );
  XOR2_X1 U11140 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10121), .Z(ADD_1071_U50) );
  AOI21_X1 U11141 ( .B1(n10123), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n10122), .ZN(
        n10124) );
  XOR2_X1 U11142 ( .A(n10124), .B(P1_ADDR_REG_5__SCAN_IN), .Z(ADD_1071_U51) );
  XOR2_X1 U11143 ( .A(n10126), .B(n10125), .Z(ADD_1071_U53) );
  XNOR2_X1 U11144 ( .A(n10128), .B(n10127), .ZN(ADD_1071_U52) );
  INV_X1 U4818 ( .A(n5682), .ZN(n6117) );
  CLKBUF_X1 U4822 ( .A(n4314), .Z(n8067) );
  CLKBUF_X1 U4823 ( .A(n8067), .Z(n8072) );
  CLKBUF_X1 U4838 ( .A(n5075), .Z(n4314) );
  CLKBUF_X1 U4854 ( .A(n5674), .Z(n6468) );
endmodule

