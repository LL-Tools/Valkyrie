

module b22_C_AntiSAT_k_256_2 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, SUB_1596_U4, SUB_1596_U62, 
        SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, 
        SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, 
        SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, 
        SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, 
        P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, 
        P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, 
        P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, 
        P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, 
        P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, 
        P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, 
        P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, 
        P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, 
        P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, 
        P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, 
        P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, 
        P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, 
        P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, 
        P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, 
        P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, 
        P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, 
        P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, 
        P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, 
        P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, 
        P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, 
        P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, 
        P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, 
        P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, 
        P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, 
        P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, 
        P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, 
        P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, 
        P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, 
        P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, 
        P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, 
        P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, 
        P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, 
        P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, 
        P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, 
        P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, 
        P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, 
        P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, 
        P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, 
        P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, 
        P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, 
        P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, 
        P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, 
        P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, 
        P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, 
        P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, 
        P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, 
        P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, 
        P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, 
        P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, 
        P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, 
        P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, 
        P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, 
        P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, 
        P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, 
        P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, 
        P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, 
        P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, 
        P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, 
        P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, 
        P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, 
        P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, 
        P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, 
        P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, 
        P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, 
        P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, 
        P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, 
        P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, 
        P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, 
        P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, 
        P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, 
        P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, 
        P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, 
        P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, 
        P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, 
        P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, 
        P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, 
        P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, 
        P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, 
        P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, 
        P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, 
        P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, 
        P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, 
        P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, 
        P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, 
        P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, 
        P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, 
        P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, 
        P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, 
        P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, 
        P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, 
        P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127,
         keyinput128, keyinput129, keyinput130, keyinput131, keyinput132,
         keyinput133, keyinput134, keyinput135, keyinput136, keyinput137,
         keyinput138, keyinput139, keyinput140, keyinput141, keyinput142,
         keyinput143, keyinput144, keyinput145, keyinput146, keyinput147,
         keyinput148, keyinput149, keyinput150, keyinput151, keyinput152,
         keyinput153, keyinput154, keyinput155, keyinput156, keyinput157,
         keyinput158, keyinput159, keyinput160, keyinput161, keyinput162,
         keyinput163, keyinput164, keyinput165, keyinput166, keyinput167,
         keyinput168, keyinput169, keyinput170, keyinput171, keyinput172,
         keyinput173, keyinput174, keyinput175, keyinput176, keyinput177,
         keyinput178, keyinput179, keyinput180, keyinput181, keyinput182,
         keyinput183, keyinput184, keyinput185, keyinput186, keyinput187,
         keyinput188, keyinput189, keyinput190, keyinput191, keyinput192,
         keyinput193, keyinput194, keyinput195, keyinput196, keyinput197,
         keyinput198, keyinput199, keyinput200, keyinput201, keyinput202,
         keyinput203, keyinput204, keyinput205, keyinput206, keyinput207,
         keyinput208, keyinput209, keyinput210, keyinput211, keyinput212,
         keyinput213, keyinput214, keyinput215, keyinput216, keyinput217,
         keyinput218, keyinput219, keyinput220, keyinput221, keyinput222,
         keyinput223, keyinput224, keyinput225, keyinput226, keyinput227,
         keyinput228, keyinput229, keyinput230, keyinput231, keyinput232,
         keyinput233, keyinput234, keyinput235, keyinput236, keyinput237,
         keyinput238, keyinput239, keyinput240, keyinput241, keyinput242,
         keyinput243, keyinput244, keyinput245, keyinput246, keyinput247,
         keyinput248, keyinput249, keyinput250, keyinput251, keyinput252,
         keyinput253, keyinput254, keyinput255;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6687, n6688, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453;

  OR2_X1 U7353 ( .A1(n7468), .A2(n6715), .ZN(n7167) );
  INV_X4 U7354 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  OR2_X1 U7355 ( .A1(n13814), .A2(n13990), .ZN(n13794) );
  OAI21_X1 U7356 ( .B1(n11666), .B2(n11665), .A(n14075), .ZN(n11956) );
  CLKBUF_X1 U7357 ( .A(n7684), .Z(n8102) );
  CLKBUF_X3 U7358 ( .A(n9932), .Z(n12895) );
  INV_X2 U7359 ( .A(n10243), .ZN(n12120) );
  XNOR2_X1 U7360 ( .A(n15106), .B(n13274), .ZN(n13961) );
  INV_X1 U7361 ( .A(n9932), .ZN(n11155) );
  NAND2_X2 U7362 ( .A1(n10367), .A2(n10083), .ZN(n10243) );
  AND2_X1 U7363 ( .A1(n10367), .A2(n10084), .ZN(n10245) );
  BUF_X2 U7364 ( .A(n8541), .Z(n9079) );
  CLKBUF_X2 U7365 ( .A(n8437), .Z(n8661) );
  INV_X1 U7366 ( .A(n7700), .ZN(n7870) );
  INV_X1 U7368 ( .A(n7672), .ZN(n6993) );
  NAND2_X1 U7369 ( .A1(n8264), .A2(n6688), .ZN(n9973) );
  NAND4_X2 U7370 ( .A1(n9948), .A2(n9947), .A3(n9946), .A4(n9945), .ZN(n13274)
         );
  XNOR2_X2 U7371 ( .A(n8795), .B(n8794), .ZN(n8900) );
  AND2_X1 U7372 ( .A1(n10052), .A2(n7606), .ZN(n7694) );
  CLKBUF_X2 U7373 ( .A(n9907), .Z(n6610) );
  INV_X1 U7374 ( .A(n9794), .ZN(n9486) );
  INV_X1 U7376 ( .A(n12063), .ZN(n12112) );
  INV_X1 U7377 ( .A(n9082), .ZN(n9026) );
  OR2_X1 U7378 ( .A1(n12398), .A2(n9397), .ZN(n8245) );
  INV_X1 U7379 ( .A(n13000), .ZN(n13173) );
  AND2_X1 U7380 ( .A1(n9907), .A2(n9906), .ZN(n12971) );
  INV_X1 U7381 ( .A(n11374), .ZN(n12855) );
  INV_X2 U7382 ( .A(n10245), .ZN(n12063) );
  INV_X1 U7383 ( .A(n8295), .ZN(n8297) );
  INV_X1 U7384 ( .A(n10209), .ZN(n9255) );
  INV_X1 U7385 ( .A(n12422), .ZN(n12449) );
  INV_X1 U7386 ( .A(n7700), .ZN(n8045) );
  OR2_X1 U7387 ( .A1(n12274), .A2(n7249), .ZN(n7248) );
  INV_X1 U7388 ( .A(n7040), .ZN(n7039) );
  INV_X1 U7389 ( .A(n10442), .ZN(n7214) );
  INV_X2 U7390 ( .A(n9973), .ZN(n7946) );
  NAND2_X1 U7391 ( .A1(n8029), .A2(n8028), .ZN(n8040) );
  INV_X1 U7392 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8267) );
  INV_X1 U7394 ( .A(n10406), .ZN(n12845) );
  INV_X1 U7395 ( .A(n13404), .ZN(n9915) );
  XNOR2_X1 U7396 ( .A(n15113), .B(n13950), .ZN(n13190) );
  CLKBUF_X3 U7397 ( .A(n13404), .Z(n6611) );
  INV_X1 U7398 ( .A(n14249), .ZN(n10939) );
  OR2_X1 U7401 ( .A1(n11972), .A2(n14561), .ZN(n7601) );
  INV_X2 U7402 ( .A(n10252), .ZN(n12121) );
  XNOR2_X1 U7403 ( .A(n8323), .B(SI_5_), .ZN(n8447) );
  INV_X1 U7404 ( .A(n7674), .ZN(n8099) );
  OAI211_X1 U7405 ( .C1(n9525), .C2(n7674), .A(n6992), .B(n6990), .ZN(n10187)
         );
  XNOR2_X1 U7406 ( .A(n12794), .B(n12793), .ZN(n12872) );
  INV_X1 U7407 ( .A(n13394), .ZN(n13980) );
  NAND2_X1 U7410 ( .A1(n14077), .A2(n14076), .ZN(n14075) );
  INV_X1 U7411 ( .A(n10794), .ZN(n10746) );
  AND2_X1 U7412 ( .A1(n8384), .A2(n6791), .ZN(n8385) );
  XNOR2_X1 U7413 ( .A(n7555), .B(n8447), .ZN(n10259) );
  INV_X1 U7414 ( .A(n10565), .ZN(n15192) );
  AND2_X1 U7415 ( .A1(n11544), .A2(n11543), .ZN(n13064) );
  AND4_X1 U7416 ( .A1(n6621), .A2(n6620), .A3(n6619), .A4(n9493), .ZN(n6606)
         );
  XNOR2_X1 U7417 ( .A(n9619), .B(P2_IR_REG_21__SCAN_IN), .ZN(n9907) );
  INV_X1 U7418 ( .A(n12340), .ZN(n14735) );
  AND4_X1 U7419 ( .A1(n8404), .A2(n8403), .A3(n8402), .A4(n8401), .ZN(n6607)
         );
  INV_X1 U7420 ( .A(n8918), .ZN(n6612) );
  OR2_X2 U7421 ( .A1(n11380), .A2(n13197), .ZN(n7517) );
  OAI21_X2 U7422 ( .B1(n10231), .B2(n8914), .A(n6838), .ZN(n10829) );
  OAI21_X1 U7423 ( .B1(n8066), .B2(n8065), .A(n8067), .ZN(n8078) );
  NOR2_X2 U7424 ( .A1(n15444), .A2(n9347), .ZN(n9350) );
  NAND2_X1 U7425 ( .A1(n8264), .A2(n6688), .ZN(n6608) );
  OR2_X2 U7426 ( .A1(n10052), .A2(n8267), .ZN(n7630) );
  NAND2_X2 U7427 ( .A1(n9627), .A2(n13253), .ZN(n10878) );
  NAND2_X2 U7428 ( .A1(n6864), .A2(n6862), .ZN(n8310) );
  AOI211_X2 U7429 ( .C1(n8109), .C2(n8252), .A(n8256), .B(n8108), .ZN(n8111)
         );
  OR2_X2 U7430 ( .A1(n13183), .A2(n10170), .ZN(n10471) );
  XNOR2_X2 U7431 ( .A(n9360), .B(n9359), .ZN(n14877) );
  INV_X1 U7432 ( .A(n6607), .ZN(n6609) );
  XNOR2_X2 U7433 ( .A(n7967), .B(n11203), .ZN(n7966) );
  NAND2_X2 U7434 ( .A1(n7156), .A2(n7155), .ZN(n7967) );
  NAND2_X1 U7435 ( .A1(n8321), .A2(n8320), .ZN(n7555) );
  NAND2_X2 U7436 ( .A1(n7621), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7622) );
  AOI211_X2 U7437 ( .C1(n15329), .C2(n12350), .A(n12349), .B(n12348), .ZN(
        n12351) );
  OAI22_X2 U7438 ( .A1(n11150), .A2(n11149), .B1(n11148), .B2(n11147), .ZN(
        n11159) );
  OAI21_X2 U7439 ( .B1(n12164), .B2(n7383), .A(n7381), .ZN(n9390) );
  OAI21_X2 U7440 ( .B1(n12185), .B2(n12166), .A(n12165), .ZN(n12164) );
  XNOR2_X2 U7441 ( .A(n7696), .B(n7695), .ZN(n10062) );
  XNOR2_X1 U7442 ( .A(n8312), .B(SI_2_), .ZN(n8417) );
  NAND2_X2 U7443 ( .A1(n8482), .A2(n8481), .ZN(n14954) );
  XNOR2_X2 U7444 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n7656) );
  OAI21_X2 U7445 ( .B1(n8040), .B2(n8039), .A(n8041), .ZN(n8053) );
  AOI21_X2 U7446 ( .B1(n12461), .B2(n12399), .A(n6739), .ZN(n12432) );
  OAI22_X2 U7447 ( .A1(n11180), .A2(n11179), .B1(n13268), .B2(n15061), .ZN(
        n11379) );
  INV_X1 U7448 ( .A(n15063), .ZN(n11180) );
  NAND2_X2 U7449 ( .A1(n12391), .A2(n12390), .ZN(n12475) );
  OAI21_X2 U7450 ( .B1(n9356), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n14872), .ZN(
        n9360) );
  AND2_X2 U7451 ( .A1(n12969), .A2(n6610), .ZN(n13000) );
  NAND2_X1 U7452 ( .A1(n10198), .A2(n9906), .ZN(n13404) );
  NAND2_X1 U7453 ( .A1(n7305), .A2(n7304), .ZN(n12922) );
  XNOR2_X2 U7454 ( .A(n12591), .B(n12422), .ZN(n7040) );
  AOI21_X1 U7455 ( .B1(n14754), .B2(n12322), .A(n12323), .ZN(n12335) );
  AND2_X1 U7456 ( .A1(n6972), .A2(n6730), .ZN(n13788) );
  INV_X1 U7457 ( .A(n13357), .ZN(n6614) );
  NAND2_X1 U7458 ( .A1(n13917), .A2(n7586), .ZN(n13894) );
  NAND2_X1 U7459 ( .A1(n13390), .A2(n13182), .ZN(n13409) );
  NAND2_X1 U7460 ( .A1(n13919), .A2(n13918), .ZN(n13917) );
  NAND2_X1 U7461 ( .A1(n11449), .A2(n6849), .ZN(n11509) );
  OR2_X1 U7462 ( .A1(n13985), .A2(n13790), .ZN(n13182) );
  OR2_X1 U7463 ( .A1(n9000), .A2(n8999), .ZN(n6662) );
  NOR2_X1 U7464 ( .A1(n6645), .A2(n7229), .ZN(n7228) );
  INV_X1 U7465 ( .A(n12464), .ZN(n9397) );
  AOI21_X1 U7466 ( .B1(n8939), .B2(n6615), .A(n6786), .ZN(n6658) );
  AND2_X1 U7467 ( .A1(n14830), .A2(n11371), .ZN(n6983) );
  NAND2_X1 U7468 ( .A1(n8527), .A2(n8526), .ZN(n14964) );
  INV_X1 U7469 ( .A(n8941), .ZN(n6615) );
  XNOR2_X1 U7470 ( .A(n7579), .B(n8540), .ZN(n11151) );
  OAI21_X1 U7471 ( .B1(n8534), .B2(n8335), .A(n8537), .ZN(n7579) );
  INV_X4 U7472 ( .A(n12063), .ZN(n12073) );
  INV_X2 U7473 ( .A(n12063), .ZN(n12054) );
  AND2_X1 U7474 ( .A1(n8907), .A2(n8813), .ZN(n11138) );
  INV_X2 U7475 ( .A(n14251), .ZN(n11135) );
  INV_X1 U7476 ( .A(n14248), .ZN(n10961) );
  AND2_X1 U7477 ( .A1(n11952), .A2(n10448), .ZN(n9154) );
  INV_X1 U7478 ( .A(n9160), .ZN(n10214) );
  NOR2_X2 U7479 ( .A1(n11130), .A2(n14125), .ZN(n11129) );
  INV_X1 U7480 ( .A(n10255), .ZN(n10594) );
  INV_X1 U7481 ( .A(n12988), .ZN(n15100) );
  INV_X1 U7482 ( .A(n15360), .ZN(n7649) );
  INV_X1 U7484 ( .A(n10317), .ZN(n15093) );
  NAND2_X1 U7485 ( .A1(n8125), .A2(n8124), .ZN(n11952) );
  CLKBUF_X3 U7486 ( .A(n8436), .Z(n6617) );
  CLKBUF_X1 U7488 ( .A(n8112), .Z(n6687) );
  INV_X2 U7489 ( .A(n14671), .ZN(n8296) );
  NAND2_X4 U7490 ( .A1(n10878), .A2(n9794), .ZN(n13164) );
  INV_X1 U7491 ( .A(n9919), .ZN(n6613) );
  NAND2_X1 U7492 ( .A1(n9545), .A2(n9544), .ZN(n10135) );
  NAND2_X1 U7493 ( .A1(n9545), .A2(n11989), .ZN(n10407) );
  BUF_X1 U7494 ( .A(n9541), .Z(n11989) );
  INV_X1 U7495 ( .A(n7638), .ZN(n12340) );
  NAND2_X2 U7496 ( .A1(n9794), .A2(P1_U3086), .ZN(n12137) );
  INV_X8 U7497 ( .A(n9910), .ZN(n9794) );
  AND3_X2 U7498 ( .A1(n10052), .A2(n7605), .A3(n7604), .ZN(n6722) );
  NOR2_X1 U7499 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n8284) );
  NOR2_X1 U7500 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n8283) );
  NOR2_X1 U7501 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n8282) );
  NOR2_X1 U7502 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n6621) );
  INV_X4 U7504 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  AND3_X1 U7505 ( .A1(n13251), .A2(n7125), .A3(n13250), .ZN(n13258) );
  AOI21_X1 U7506 ( .B1(n13154), .B2(n13153), .A(n13152), .ZN(n13236) );
  NAND2_X1 U7507 ( .A1(n6670), .A2(n6669), .ZN(n9138) );
  OAI22_X1 U7508 ( .A1(n9047), .A2(n6668), .B1(n6671), .B2(n9048), .ZN(n9093)
         );
  NAND2_X1 U7509 ( .A1(n9035), .A2(n9036), .ZN(n9034) );
  OAI22_X1 U7510 ( .A1(n9031), .A2(n6672), .B1(n6673), .B2(n9032), .ZN(n9035)
         );
  AOI211_X1 U7511 ( .C1(n14716), .C2(n12002), .A(n12001), .B(n12000), .ZN(
        n12003) );
  NAND2_X1 U7512 ( .A1(n6648), .A2(n6646), .ZN(n7234) );
  OR2_X1 U7513 ( .A1(n14564), .A2(n14959), .ZN(n7109) );
  INV_X1 U7514 ( .A(n12408), .ZN(n7194) );
  AND2_X1 U7515 ( .A1(n14563), .A2(n6826), .ZN(n7107) );
  OAI21_X1 U7516 ( .B1(n12828), .B2(n7336), .A(n7334), .ZN(n12899) );
  OR2_X1 U7517 ( .A1(n14102), .A2(n14103), .ZN(n14188) );
  NAND2_X1 U7518 ( .A1(n12922), .A2(n12921), .ZN(n12828) );
  OR2_X1 U7519 ( .A1(n13993), .A2(n13941), .ZN(n13803) );
  NAND2_X1 U7520 ( .A1(n12426), .A2(n12435), .ZN(n7210) );
  OAI21_X1 U7521 ( .B1(n13802), .B2(n7538), .A(n7534), .ZN(n13399) );
  INV_X1 U7522 ( .A(n8245), .ZN(n7463) );
  NAND2_X1 U7523 ( .A1(n7216), .A2(n7217), .ZN(n12486) );
  OAI21_X2 U7524 ( .B1(n14199), .B2(n7438), .A(n7436), .ZN(n14176) );
  OAI21_X1 U7525 ( .B1(n12795), .B2(n7308), .A(n12810), .ZN(n7306) );
  OR2_X1 U7526 ( .A1(n14388), .A2(n7494), .ZN(n7493) );
  NAND2_X1 U7527 ( .A1(n6636), .A2(n6634), .ZN(n13982) );
  OR2_X1 U7528 ( .A1(n6661), .A2(n9002), .ZN(n9003) );
  NOR2_X1 U7529 ( .A1(n13414), .A2(n13413), .ZN(n13987) );
  NAND2_X1 U7530 ( .A1(n6637), .A2(n6635), .ZN(n6634) );
  AND2_X1 U7531 ( .A1(n9048), .A2(n6671), .ZN(n6668) );
  OR2_X1 U7532 ( .A1(n6988), .A2(n13391), .ZN(n6636) );
  AND2_X1 U7533 ( .A1(n13357), .A2(n6638), .ZN(n6635) );
  AND2_X1 U7534 ( .A1(n6663), .A2(n6662), .ZN(n6661) );
  NAND2_X1 U7535 ( .A1(n13411), .A2(n13390), .ZN(n6637) );
  AND2_X1 U7536 ( .A1(n7601), .A2(n11973), .ZN(n14559) );
  XNOR2_X1 U7537 ( .A(n12023), .B(n12021), .ZN(n14219) );
  AND2_X1 U7538 ( .A1(n7254), .A2(n14737), .ZN(n12309) );
  INV_X1 U7539 ( .A(n7536), .ZN(n7534) );
  NAND2_X1 U7540 ( .A1(n9025), .A2(n6650), .ZN(n6649) );
  NAND2_X1 U7541 ( .A1(n14461), .A2(n8699), .ZN(n14434) );
  NOR2_X1 U7542 ( .A1(n6789), .A2(n6647), .ZN(n6646) );
  AND2_X1 U7543 ( .A1(n9032), .A2(n6673), .ZN(n6672) );
  NAND2_X1 U7544 ( .A1(n11931), .A2(n11930), .ZN(n12013) );
  OR2_X1 U7545 ( .A1(n13369), .A2(n6976), .ZN(n6972) );
  AND2_X1 U7546 ( .A1(n9028), .A2(n7235), .ZN(n6789) );
  XNOR2_X1 U7547 ( .A(n7248), .B(n12317), .ZN(n12275) );
  INV_X1 U7548 ( .A(n9030), .ZN(n6673) );
  NAND2_X1 U7549 ( .A1(n7572), .A2(n7567), .ZN(n13369) );
  OR2_X1 U7550 ( .A1(n6718), .A2(n12368), .ZN(n12567) );
  NAND2_X1 U7551 ( .A1(n13874), .A2(n7568), .ZN(n7572) );
  NOR2_X1 U7552 ( .A1(n6650), .A2(n9025), .ZN(n6647) );
  OAI21_X1 U7553 ( .B1(n13888), .B2(n13872), .A(n13878), .ZN(n13874) );
  NAND2_X1 U7554 ( .A1(n6643), .A2(n6644), .ZN(n8969) );
  NAND2_X1 U7555 ( .A1(n7969), .A2(n7968), .ZN(n7980) );
  OR2_X1 U7556 ( .A1(n12288), .A2(n12287), .ZN(n12295) );
  NAND2_X1 U7557 ( .A1(n11451), .A2(n11450), .ZN(n11449) );
  NAND2_X1 U7558 ( .A1(n12831), .A2(n12830), .ZN(n13990) );
  NOR2_X1 U7559 ( .A1(n13889), .A2(n13893), .ZN(n13888) );
  OAI21_X1 U7560 ( .B1(n8951), .B2(n8950), .A(n8949), .ZN(n8956) );
  NAND2_X1 U7561 ( .A1(n13903), .A2(n13364), .ZN(n13889) );
  NAND2_X1 U7562 ( .A1(n11752), .A2(n7588), .ZN(n11754) );
  NAND2_X1 U7563 ( .A1(n9000), .A2(n8999), .ZN(n6664) );
  NAND2_X1 U7564 ( .A1(n12253), .A2(n12252), .ZN(n12286) );
  NAND2_X1 U7565 ( .A1(n13905), .A2(n13904), .ZN(n13903) );
  INV_X1 U7566 ( .A(n13391), .ZN(n6638) );
  NOR2_X1 U7567 ( .A1(n11649), .A2(n11648), .ZN(n14296) );
  NAND2_X1 U7568 ( .A1(n6660), .A2(n7236), .ZN(n8947) );
  NAND2_X1 U7569 ( .A1(n14806), .A2(n6861), .ZN(n11596) );
  NAND2_X1 U7570 ( .A1(n7928), .A2(n7927), .ZN(n7941) );
  OAI21_X1 U7571 ( .B1(n8940), .B2(n6659), .A(n6658), .ZN(n6660) );
  NAND3_X1 U7572 ( .A1(n7793), .A2(n7813), .A3(n7792), .ZN(n15417) );
  NAND2_X1 U7573 ( .A1(n8676), .A2(n8675), .ZN(n14609) );
  AOI21_X1 U7574 ( .B1(n14801), .B2(n14800), .A(n6982), .ZN(n11582) );
  NAND2_X1 U7575 ( .A1(n7911), .A2(n7910), .ZN(n7926) );
  NAND2_X1 U7576 ( .A1(n6633), .A2(n6794), .ZN(n14801) );
  AOI21_X1 U7577 ( .B1(n7228), .B2(n7231), .A(n7227), .ZN(n6644) );
  NAND2_X1 U7578 ( .A1(n6628), .A2(n6625), .ZN(n6633) );
  NAND2_X1 U7579 ( .A1(n6628), .A2(n6626), .ZN(n11561) );
  NAND2_X1 U7580 ( .A1(n6632), .A2(n6631), .ZN(n11406) );
  NAND2_X1 U7581 ( .A1(n6632), .A2(n6629), .ZN(n6628) );
  AND2_X1 U7582 ( .A1(n6918), .A2(n6916), .ZN(n7263) );
  NAND2_X1 U7583 ( .A1(n6677), .A2(n6867), .ZN(n8930) );
  AND2_X1 U7584 ( .A1(n6762), .A2(n8957), .ZN(n6645) );
  OR2_X1 U7585 ( .A1(n11054), .A2(n7247), .ZN(n7244) );
  OR2_X1 U7586 ( .A1(n11357), .A2(n11378), .ZN(n6632) );
  AND2_X1 U7587 ( .A1(n6626), .A2(n13197), .ZN(n6625) );
  NOR2_X1 U7588 ( .A1(n10659), .A2(n10660), .ZN(n11057) );
  NOR2_X1 U7589 ( .A1(n6630), .A2(n6983), .ZN(n6629) );
  AOI22_X1 U7590 ( .A1(n15052), .A2(n15062), .B1(n11178), .B2(n15061), .ZN(
        n11357) );
  OR2_X1 U7591 ( .A1(n14634), .A2(n14095), .ZN(n8960) );
  NAND2_X1 U7592 ( .A1(n7863), .A2(n7862), .ZN(n7879) );
  OAI22_X1 U7593 ( .A1(n11174), .A2(n11173), .B1(n7074), .B2(n13269), .ZN(
        n15052) );
  NOR2_X1 U7594 ( .A1(n7416), .A2(n7415), .ZN(n7414) );
  NAND2_X1 U7595 ( .A1(n6627), .A2(n13196), .ZN(n6626) );
  INV_X1 U7596 ( .A(n6631), .ZN(n6630) );
  AND2_X1 U7597 ( .A1(n15327), .A2(n10658), .ZN(n10659) );
  OR2_X1 U7598 ( .A1(n15064), .A2(n13040), .ZN(n11412) );
  NAND2_X1 U7599 ( .A1(n11741), .A2(n11740), .ZN(n14037) );
  NAND2_X1 U7600 ( .A1(n6622), .A2(n7528), .ZN(n11174) );
  XNOR2_X1 U7601 ( .A(n7861), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n7860) );
  INV_X1 U7602 ( .A(n6983), .ZN(n6627) );
  NAND2_X1 U7603 ( .A1(n7529), .A2(n10892), .ZN(n6622) );
  NOR2_X1 U7604 ( .A1(n6615), .A2(n8939), .ZN(n6659) );
  AOI21_X1 U7605 ( .B1(n10349), .B2(n10350), .A(n9167), .ZN(n15196) );
  OR2_X1 U7606 ( .A1(n15151), .A2(n13267), .ZN(n6631) );
  OAI21_X1 U7607 ( .B1(n10846), .B2(n7531), .A(n7530), .ZN(n7529) );
  NAND2_X1 U7608 ( .A1(n8585), .A2(n8584), .ZN(n14639) );
  NAND2_X1 U7609 ( .A1(n6842), .A2(n10656), .ZN(n10657) );
  NAND2_X1 U7610 ( .A1(n8546), .A2(n8545), .ZN(n14843) );
  NOR2_X1 U7611 ( .A1(n15446), .A2(n15445), .ZN(n15444) );
  NAND2_X1 U7612 ( .A1(n10990), .A2(n10989), .ZN(n15061) );
  AOI21_X1 U7613 ( .B1(n10522), .B2(n10521), .A(n10520), .ZN(n10698) );
  NOR2_X1 U7614 ( .A1(n8944), .A2(n8942), .ZN(n6786) );
  NAND2_X1 U7615 ( .A1(n10387), .A2(n10386), .ZN(n13947) );
  NOR2_X1 U7616 ( .A1(n14685), .A2(n9343), .ZN(n9344) );
  NAND2_X1 U7617 ( .A1(n13946), .A2(n10389), .ZN(n10522) );
  INV_X2 U7618 ( .A(n10738), .ZN(n12119) );
  OAI211_X1 U7619 ( .C1(n6641), .C2(n6640), .A(n13961), .B(n6623), .ZN(n13946)
         );
  CLKBUF_X1 U7620 ( .A(n10738), .Z(n12062) );
  NAND2_X1 U7621 ( .A1(n6641), .A2(n10327), .ZN(n10387) );
  XOR2_X1 U7622 ( .A(n10654), .B(n15279), .Z(n15278) );
  NAND2_X1 U7623 ( .A1(n10753), .A2(n10752), .ZN(n13022) );
  INV_X1 U7624 ( .A(n8921), .ZN(n6674) );
  NAND2_X2 U7625 ( .A1(n10405), .A2(n10404), .ZN(n13009) );
  OR2_X1 U7626 ( .A1(n13190), .A2(n10382), .ZN(n10508) );
  NAND2_X1 U7627 ( .A1(n10386), .A2(n13186), .ZN(n6623) );
  NAND2_X1 U7628 ( .A1(n10328), .A2(n10329), .ZN(n6641) );
  INV_X1 U7629 ( .A(n11138), .ZN(n9097) );
  NAND2_X1 U7630 ( .A1(n10653), .A2(n10652), .ZN(n10654) );
  INV_X1 U7631 ( .A(n8915), .ZN(n6653) );
  CLKBUF_X1 U7632 ( .A(n11374), .Z(n15065) );
  INV_X1 U7633 ( .A(n13186), .ZN(n10327) );
  AND2_X1 U7634 ( .A1(n7222), .A2(n7224), .ZN(n8918) );
  NAND2_X1 U7635 ( .A1(n10325), .A2(n10465), .ZN(n10326) );
  INV_X1 U7636 ( .A(n10386), .ZN(n6640) );
  NAND2_X1 U7637 ( .A1(n6667), .A2(n6666), .ZN(n8903) );
  NAND2_X1 U7638 ( .A1(n6909), .A2(n8446), .ZN(n14249) );
  AND4_X1 U7639 ( .A1(n7727), .A2(n7726), .A3(n7725), .A4(n7724), .ZN(n10858)
         );
  NOR2_X1 U7640 ( .A1(n10324), .A2(n9915), .ZN(n9916) );
  NAND2_X1 U7641 ( .A1(n8901), .A2(n9070), .ZN(n6667) );
  NAND2_X1 U7642 ( .A1(n10542), .A2(n10427), .ZN(n10458) );
  NAND2_X1 U7643 ( .A1(n10173), .A2(n13183), .ZN(n10325) );
  BUF_X4 U7644 ( .A(n8085), .Z(n7991) );
  AND2_X2 U7645 ( .A1(n9822), .A2(n8900), .ZN(n14712) );
  NAND2_X1 U7646 ( .A1(n7743), .A2(n7742), .ZN(n7745) );
  AND2_X1 U7647 ( .A1(n8900), .A2(n9089), .ZN(n10084) );
  OR2_X1 U7648 ( .A1(n8900), .A2(n11277), .ZN(n8901) );
  NAND4_X2 U7649 ( .A1(n8400), .A2(n8399), .A3(n8398), .A4(n8397), .ZN(n10246)
         );
  NAND2_X1 U7650 ( .A1(n10121), .A2(n10120), .ZN(n15106) );
  OAI211_X1 U7651 ( .C1(n9430), .C2(n9836), .A(n8433), .B(n8432), .ZN(n14939)
         );
  INV_X1 U7652 ( .A(n9993), .ZN(n12979) );
  NAND2_X1 U7653 ( .A1(n9936), .A2(n9935), .ZN(n12988) );
  OAI211_X1 U7654 ( .C1(n9057), .C2(n9920), .A(n7300), .B(n7299), .ZN(n10255)
         );
  INV_X1 U7655 ( .A(n10448), .ZN(n10504) );
  NAND2_X1 U7656 ( .A1(n8409), .A2(n6869), .ZN(n11130) );
  INV_X1 U7657 ( .A(n8112), .ZN(n9145) );
  INV_X1 U7658 ( .A(n13275), .ZN(n10324) );
  INV_X1 U7659 ( .A(n13275), .ZN(n6624) );
  OR2_X1 U7660 ( .A1(n9922), .A2(n9921), .ZN(n10317) );
  NAND4_X1 U7661 ( .A1(n9927), .A2(n9926), .A3(n9925), .A4(n9924), .ZN(n10319)
         );
  OR2_X1 U7662 ( .A1(n9070), .A2(n11277), .ZN(n6666) );
  AND2_X1 U7663 ( .A1(n12726), .A2(n7624), .ZN(n7666) );
  NAND4_X1 U7664 ( .A1(n9549), .A2(n9548), .A3(n9547), .A4(n9546), .ZN(n10172)
         );
  NAND4_X1 U7665 ( .A1(n10139), .A2(n10138), .A3(n10137), .A4(n10136), .ZN(
        n13950) );
  BUF_X2 U7666 ( .A(n7672), .Z(n7673) );
  AND2_X2 U7667 ( .A1(n8129), .A2(n8128), .ZN(n10448) );
  NAND4_X1 U7668 ( .A1(n9763), .A2(n9762), .A3(n9761), .A4(n9760), .ZN(n13275)
         );
  AND2_X1 U7669 ( .A1(n7089), .A2(n7088), .ZN(n9875) );
  OR2_X1 U7670 ( .A1(n13164), .A2(n9909), .ZN(n9914) );
  MUX2_X1 U7671 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8127), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n8129) );
  NAND2_X1 U7672 ( .A1(n8793), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8795) );
  XNOR2_X1 U7673 ( .A(n7945), .B(n8114), .ZN(n8112) );
  AND2_X1 U7674 ( .A1(n8297), .A2(n14671), .ZN(n8460) );
  CLKBUF_X1 U7675 ( .A(n10407), .Z(n13172) );
  NAND2_X1 U7676 ( .A1(n8294), .A2(n7512), .ZN(n14671) );
  XNOR2_X1 U7677 ( .A(n8792), .B(n8791), .ZN(n14334) );
  NAND2_X1 U7678 ( .A1(n7944), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7945) );
  OR2_X1 U7679 ( .A1(n10878), .A2(n6639), .ZN(n9912) );
  AND2_X2 U7680 ( .A1(n11939), .A2(n11989), .ZN(n10406) );
  NAND2_X1 U7681 ( .A1(n8660), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8792) );
  OAI21_X1 U7682 ( .B1(n9618), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9617) );
  NAND2_X1 U7683 ( .A1(n9618), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9619) );
  NAND2_X1 U7684 ( .A1(n7633), .A2(n7634), .ZN(n8264) );
  NAND2_X1 U7685 ( .A1(n9542), .A2(n9544), .ZN(n12775) );
  XNOR2_X1 U7686 ( .A(n8292), .B(n8291), .ZN(n8295) );
  INV_X1 U7687 ( .A(n9542), .ZN(n9545) );
  NAND2_X1 U7688 ( .A1(n7153), .A2(n7691), .ZN(n7709) );
  INV_X1 U7689 ( .A(n9089), .ZN(n11277) );
  MUX2_X1 U7690 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7632), .S(
        P3_IR_REG_28__SCAN_IN), .Z(n7634) );
  INV_X2 U7691 ( .A(n12719), .ZN(n11991) );
  NAND2_X1 U7692 ( .A1(n7512), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8292) );
  NAND2_X2 U7693 ( .A1(n9486), .A2(P1_U3086), .ZN(n14668) );
  NAND2_X1 U7694 ( .A1(n9623), .A2(n9622), .ZN(n13253) );
  XNOR2_X1 U7695 ( .A(n8799), .B(P1_IR_REG_22__SCAN_IN), .ZN(n8899) );
  XNOR2_X1 U7696 ( .A(n9537), .B(n9536), .ZN(n9542) );
  XNOR2_X1 U7697 ( .A(n8326), .B(SI_6_), .ZN(n8465) );
  INV_X1 U7698 ( .A(n9541), .ZN(n9544) );
  XNOR2_X1 U7699 ( .A(n8319), .B(SI_4_), .ZN(n8434) );
  XNOR2_X1 U7700 ( .A(n7637), .B(n7636), .ZN(n7638) );
  MUX2_X1 U7701 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9621), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n9623) );
  XNOR2_X1 U7702 ( .A(n9540), .B(n9539), .ZN(n9541) );
  NOR2_X1 U7703 ( .A1(n10107), .A2(n10108), .ZN(n10106) );
  XNOR2_X1 U7704 ( .A(n8308), .B(SI_1_), .ZN(n8392) );
  OAI21_X1 U7705 ( .B1(n8796), .B2(n7242), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n8798) );
  INV_X2 U7706 ( .A(n11849), .ZN(n6618) );
  NAND2_X1 U7707 ( .A1(n14069), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9537) );
  OAI21_X1 U7708 ( .B1(n8310), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n6839), .ZN(
        n8308) );
  NAND2_X1 U7709 ( .A1(n8573), .A2(n8572), .ZN(n8796) );
  OR2_X1 U7710 ( .A1(n9538), .A2(n6642), .ZN(n9540) );
  NAND2_X1 U7711 ( .A1(n9622), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9620) );
  AND2_X1 U7712 ( .A1(n9425), .A2(n7340), .ZN(n9783) );
  AND3_X1 U7713 ( .A1(n9425), .A2(n6695), .A3(n6986), .ZN(n9538) );
  CLKBUF_X1 U7714 ( .A(n9425), .Z(n6837) );
  OR2_X1 U7715 ( .A1(n9425), .A2(n6642), .ZN(n10191) );
  INV_X2 U7716 ( .A(n8310), .ZN(n9910) );
  NOR2_X1 U7717 ( .A1(n8864), .A2(n8280), .ZN(n8287) );
  NOR2_X1 U7718 ( .A1(n9286), .A2(n9285), .ZN(n9328) );
  AND2_X1 U7719 ( .A1(n9426), .A2(n6731), .ZN(n6695) );
  INV_X1 U7720 ( .A(n9911), .ZN(n6639) );
  AND2_X1 U7721 ( .A1(n7189), .A2(n7590), .ZN(n7188) );
  AND3_X1 U7722 ( .A1(n9409), .A2(n9408), .A3(n9407), .ZN(n9728) );
  AND2_X1 U7723 ( .A1(n7474), .A2(n8281), .ZN(n7471) );
  AND3_X1 U7724 ( .A1(n7610), .A2(n7609), .A3(n7914), .ZN(n8120) );
  AND2_X1 U7725 ( .A1(n7011), .A2(n7010), .ZN(n7189) );
  AND2_X1 U7726 ( .A1(n7342), .A2(n7341), .ZN(n7340) );
  AND2_X1 U7727 ( .A1(n7473), .A2(n7472), .ZN(n8419) );
  AND2_X1 U7728 ( .A1(n6875), .A2(n6874), .ZN(n7406) );
  AND2_X1 U7729 ( .A1(n9470), .A2(n9471), .ZN(n9494) );
  INV_X1 U7730 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n8858) );
  NOR2_X1 U7731 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n6874) );
  INV_X1 U7732 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n8281) );
  NOR2_X1 U7733 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n6875) );
  INV_X4 U7734 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7735 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n9493) );
  NOR2_X1 U7736 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n9407) );
  NOR2_X1 U7737 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n9408) );
  NOR2_X1 U7738 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n9409) );
  INV_X1 U7739 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n10190) );
  INV_X1 U7740 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6642) );
  NOR2_X1 U7741 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n6619) );
  NOR2_X1 U7742 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n6620) );
  NOR2_X1 U7743 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n7010) );
  NOR2_X1 U7744 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n7011) );
  NOR2_X1 U7745 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_8__SCAN_IN), .ZN(
        n7604) );
  NOR2_X1 U7746 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n7605) );
  INV_X1 U7747 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n7847) );
  INV_X1 U7748 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n7894) );
  INV_X1 U7749 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n7914) );
  NOR2_X1 U7750 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_18__SCAN_IN), .ZN(
        n7609) );
  NOR2_X1 U7751 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), .ZN(
        n7610) );
  INV_X1 U7752 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n13648) );
  INV_X1 U7753 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n13643) );
  INV_X1 U7754 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n13642) );
  NOR2_X1 U7755 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n9410) );
  NOR3_X1 U7756 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .A3(
        P2_IR_REG_24__SCAN_IN), .ZN(n9412) );
  INV_X1 U7757 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n9614) );
  INV_X1 U7758 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n13636) );
  INV_X4 U7759 ( .A(n13164), .ZN(n10117) );
  XNOR2_X2 U7760 ( .A(n6624), .B(n9993), .ZN(n13183) );
  OAI211_X1 U7761 ( .C1(n13983), .C2(n15117), .A(n13982), .B(n13981), .ZN(
        n14054) );
  AOI21_X1 U7762 ( .B1(n11738), .B2(n6736), .A(n7544), .ZN(n13905) );
  INV_X2 U7763 ( .A(n10878), .ZN(n12733) );
  XNOR2_X2 U7764 ( .A(n9620), .B(n13637), .ZN(n9627) );
  AND3_X2 U7765 ( .A1(n6606), .A2(n9494), .A3(n9728), .ZN(n9425) );
  NAND2_X1 U7766 ( .A1(n8969), .A2(n8968), .ZN(n8971) );
  NAND2_X1 U7767 ( .A1(n8956), .A2(n7228), .ZN(n6643) );
  NAND3_X1 U7768 ( .A1(n9023), .A2(n9022), .A3(n6649), .ZN(n6648) );
  INV_X1 U7769 ( .A(n9024), .ZN(n6650) );
  NAND2_X1 U7770 ( .A1(n6651), .A2(n8916), .ZN(n8917) );
  NAND3_X1 U7771 ( .A1(n6654), .A2(n8913), .A3(n6652), .ZN(n6651) );
  NAND2_X1 U7772 ( .A1(n8898), .A2(n6653), .ZN(n6652) );
  NAND2_X1 U7773 ( .A1(n6655), .A2(n9097), .ZN(n6654) );
  NAND3_X1 U7774 ( .A1(n6656), .A2(n8905), .A3(n8906), .ZN(n6655) );
  NAND2_X1 U7775 ( .A1(n6657), .A2(n9082), .ZN(n6656) );
  INV_X1 U7776 ( .A(n9096), .ZN(n6657) );
  NAND3_X1 U7777 ( .A1(n6665), .A2(n8998), .A3(n6664), .ZN(n6663) );
  NAND2_X1 U7778 ( .A1(n8990), .A2(n7585), .ZN(n6665) );
  NOR2_X1 U7779 ( .A1(n9125), .A2(n9120), .ZN(n6669) );
  INV_X1 U7780 ( .A(n9093), .ZN(n6670) );
  INV_X1 U7781 ( .A(n9046), .ZN(n6671) );
  NOR2_X1 U7782 ( .A1(n8924), .A2(n6674), .ZN(n6675) );
  NAND2_X1 U7783 ( .A1(n8922), .A2(n6675), .ZN(n6676) );
  NAND2_X1 U7784 ( .A1(n8922), .A2(n8921), .ZN(n6680) );
  NAND2_X1 U7785 ( .A1(n6676), .A2(n8923), .ZN(n6679) );
  NAND3_X1 U7786 ( .A1(n6679), .A2(n6790), .A3(n6678), .ZN(n6677) );
  NAND2_X1 U7787 ( .A1(n6680), .A2(n8924), .ZN(n6678) );
  NAND2_X1 U7789 ( .A1(n8419), .A2(n7471), .ZN(n8438) );
  AOI21_X2 U7790 ( .B1(n11852), .B2(n11854), .A(n11853), .ZN(n12175) );
  NAND2_X1 U7791 ( .A1(n9627), .A2(n13253), .ZN(n6681) );
  AND2_X1 U7792 ( .A1(n8297), .A2(n8296), .ZN(n6682) );
  AND2_X1 U7793 ( .A1(n8297), .A2(n8296), .ZN(n6683) );
  NAND2_X2 U7794 ( .A1(n9908), .A2(n13331), .ZN(n10171) );
  NOR3_X2 U7795 ( .A1(n14435), .A2(n14572), .A3(n7102), .ZN(n8854) );
  OAI22_X1 U7796 ( .A1(n10698), .A2(n13191), .B1(n15122), .B2(n13272), .ZN(
        n10846) );
  CLKBUF_X1 U7797 ( .A(n14253), .Z(n6684) );
  OAI211_X1 U7798 ( .C1(P1_IR_REG_31__SCAN_IN), .C2(P1_IR_REG_27__SCAN_IN), 
        .A(n7289), .B(n8389), .ZN(n14253) );
  AOI22_X2 U7799 ( .A1(n11177), .A2(n13194), .B1(n13027), .B2(n13269), .ZN(
        n15063) );
  AOI21_X2 U7800 ( .B1(n11596), .B2(n11595), .A(n6749), .ZN(n11597) );
  INV_X1 U7801 ( .A(n13000), .ZN(n6685) );
  XNOR2_X1 U7803 ( .A(n7637), .B(n7636), .ZN(n6688) );
  NOR2_X2 U7804 ( .A1(n11159), .A2(n11158), .ZN(n11301) );
  AOI21_X2 U7805 ( .B1(n7562), .B2(n7564), .A(n7561), .ZN(n13919) );
  OAI21_X2 U7806 ( .B1(n10845), .B2(n10844), .A(n10843), .ZN(n10893) );
  NAND2_X2 U7807 ( .A1(n10691), .A2(n10690), .ZN(n10845) );
  INV_X1 U7808 ( .A(n8102), .ZN(n6690) );
  NOR2_X2 U7809 ( .A1(n7625), .A2(n7624), .ZN(n7595) );
  OAI22_X2 U7810 ( .A1(n10893), .A2(n10892), .B1(n15137), .B2(n10922), .ZN(
        n11177) );
  AND2_X1 U7811 ( .A1(n7036), .A2(n12419), .ZN(n7035) );
  NAND2_X1 U7812 ( .A1(n7037), .A2(n7039), .ZN(n7036) );
  INV_X1 U7813 ( .A(n8820), .ZN(n7296) );
  OR2_X1 U7814 ( .A1(n12387), .A2(n12488), .ZN(n8230) );
  NAND2_X1 U7815 ( .A1(n6694), .A2(n6949), .ZN(n6946) );
  INV_X1 U7816 ( .A(n9057), .ZN(n8436) );
  OAI21_X1 U7817 ( .B1(n8596), .B2(n8350), .A(n8355), .ZN(n8619) );
  AOI21_X1 U7818 ( .B1(n8354), .B2(n8600), .A(n8353), .ZN(n8355) );
  OAI21_X1 U7819 ( .B1(n8349), .B2(n9661), .A(n8600), .ZN(n8350) );
  INV_X1 U7820 ( .A(n13801), .ZN(n6971) );
  NAND2_X1 U7821 ( .A1(n14877), .A2(n15036), .ZN(n14876) );
  OAI21_X1 U7822 ( .B1(n12982), .B2(n12981), .A(n12980), .ZN(n12984) );
  OR2_X1 U7823 ( .A1(n12985), .A2(n12987), .ZN(n7365) );
  NAND2_X1 U7824 ( .A1(n9013), .A2(n9015), .ZN(n7225) );
  AOI21_X1 U7825 ( .B1(n7049), .B2(n7047), .A(n6758), .ZN(n7046) );
  INV_X1 U7826 ( .A(n7050), .ZN(n7047) );
  INV_X1 U7827 ( .A(n8163), .ZN(n7445) );
  NOR2_X1 U7828 ( .A1(n7287), .A2(n8834), .ZN(n7286) );
  INV_X1 U7829 ( .A(n8832), .ZN(n7287) );
  INV_X1 U7830 ( .A(n8674), .ZN(n8684) );
  AOI21_X1 U7831 ( .B1(n7035), .B2(n7033), .A(n7032), .ZN(n7031) );
  INV_X1 U7832 ( .A(n8251), .ZN(n7032) );
  OR2_X1 U7833 ( .A1(n12426), .A2(n12402), .ZN(n8249) );
  INV_X1 U7834 ( .A(n8241), .ZN(n7009) );
  NOR2_X1 U7835 ( .A1(n12388), .A2(n7220), .ZN(n7219) );
  INV_X1 U7836 ( .A(n12385), .ZN(n7220) );
  INV_X1 U7837 ( .A(n7666), .ZN(n7700) );
  AND2_X1 U7838 ( .A1(n7174), .A2(n7744), .ZN(n7173) );
  INV_X1 U7839 ( .A(n7747), .ZN(n7174) );
  OAI21_X1 U7840 ( .B1(n7315), .B2(n7314), .A(n10757), .ZN(n7313) );
  INV_X1 U7841 ( .A(n7523), .ZN(n7522) );
  OAI21_X1 U7842 ( .B1(n7598), .B2(n7526), .A(n7524), .ZN(n7523) );
  NAND2_X1 U7843 ( .A1(n7527), .A2(n7525), .ZN(n7524) );
  INV_X1 U7844 ( .A(n13374), .ZN(n7525) );
  NAND2_X1 U7845 ( .A1(n13403), .A2(n13394), .ZN(n13381) );
  INV_X1 U7846 ( .A(n13354), .ZN(n13373) );
  INV_X1 U7847 ( .A(n7549), .ZN(n7548) );
  NAND2_X1 U7848 ( .A1(n13366), .A2(n13875), .ZN(n7571) );
  NOR2_X1 U7849 ( .A1(n13867), .A2(n7569), .ZN(n7568) );
  INV_X1 U7850 ( .A(n7583), .ZN(n7569) );
  NAND2_X1 U7851 ( .A1(n6857), .A2(n6856), .ZN(n10738) );
  INV_X1 U7852 ( .A(n14712), .ZN(n6856) );
  INV_X1 U7853 ( .A(n10243), .ZN(n6857) );
  NAND2_X1 U7854 ( .A1(n7491), .A2(n7496), .ZN(n14357) );
  XNOR2_X1 U7855 ( .A(n14585), .B(n8728), .ZN(n14406) );
  OR2_X1 U7856 ( .A1(n14620), .A2(n8987), .ZN(n8992) );
  OAI21_X1 U7857 ( .B1(n11193), .B2(n7296), .A(n8821), .ZN(n7295) );
  NAND2_X1 U7858 ( .A1(n6607), .A2(n11130), .ZN(n9096) );
  NAND2_X1 U7859 ( .A1(n14514), .A2(n8992), .ZN(n14494) );
  NAND2_X1 U7860 ( .A1(n7124), .A2(n9074), .ZN(n7114) );
  AOI21_X1 U7861 ( .B1(n8746), .B2(n7149), .A(n7148), .ZN(n7147) );
  INV_X1 U7862 ( .A(n8759), .ZN(n7148) );
  OAI21_X1 U7863 ( .B1(n8733), .B2(n8732), .A(n8731), .ZN(n8747) );
  XNOR2_X1 U7864 ( .A(n8730), .B(SI_24_), .ZN(n8733) );
  NAND2_X1 U7865 ( .A1(n8369), .A2(n6955), .ZN(n8656) );
  INV_X1 U7866 ( .A(n8642), .ZN(n6956) );
  AND2_X1 U7867 ( .A1(n8373), .A2(n8372), .ZN(n8655) );
  NAND2_X1 U7868 ( .A1(n8361), .A2(n8360), .ZN(n8632) );
  NAND2_X1 U7869 ( .A1(n8619), .A2(n8618), .ZN(n8361) );
  NAND2_X1 U7870 ( .A1(n6961), .A2(n6959), .ZN(n8568) );
  AOI21_X1 U7871 ( .B1(n6963), .B2(n6966), .A(n6960), .ZN(n6959) );
  INV_X1 U7872 ( .A(n8345), .ZN(n6960) );
  NAND2_X1 U7873 ( .A1(n8506), .A2(n8332), .ZN(n7151) );
  INV_X1 U7874 ( .A(n8505), .ZN(n8332) );
  XNOR2_X1 U7875 ( .A(n9291), .B(n15273), .ZN(n9323) );
  AOI22_X1 U7876 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n9296), .B1(n9295), .B2(
        n9345), .ZN(n9349) );
  AOI21_X1 U7877 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n9300), .A(n9299), .ZN(
        n9301) );
  NOR2_X1 U7878 ( .A1(n9353), .A2(n9352), .ZN(n9299) );
  AOI21_X1 U7879 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n9307), .A(n9306), .ZN(
        n9363) );
  NOR2_X1 U7880 ( .A1(n9357), .A2(n9358), .ZN(n9306) );
  NAND2_X1 U7881 ( .A1(n6608), .A2(n9794), .ZN(n7672) );
  OR2_X1 U7882 ( .A1(n12410), .A2(n12232), .ZN(n8252) );
  CLKBUF_X1 U7883 ( .A(n7595), .Z(n7684) );
  INV_X1 U7884 ( .A(n7624), .ZN(n7623) );
  INV_X1 U7885 ( .A(n8237), .ZN(n7470) );
  INV_X1 U7886 ( .A(n12386), .ZN(n12488) );
  AOI21_X1 U7887 ( .B1(n7451), .B2(n7449), .A(n6761), .ZN(n7448) );
  INV_X1 U7888 ( .A(n7454), .ZN(n7449) );
  AND2_X1 U7889 ( .A1(n12375), .A2(n12373), .ZN(n7221) );
  NAND2_X1 U7890 ( .A1(n11353), .A2(n8186), .ZN(n11527) );
  NAND2_X1 U7891 ( .A1(n8081), .A2(n8080), .ZN(n8090) );
  NAND2_X1 U7892 ( .A1(n8004), .A2(n8003), .ZN(n8017) );
  NAND2_X1 U7893 ( .A1(n7980), .A2(n7979), .ZN(n7187) );
  AND2_X1 U7894 ( .A1(n7780), .A2(n7767), .ZN(n7768) );
  NAND2_X1 U7895 ( .A1(n7745), .A2(n7173), .ZN(n7766) );
  NAND2_X1 U7896 ( .A1(n7732), .A2(n7731), .ZN(n7743) );
  OR2_X1 U7897 ( .A1(n13165), .A2(n13164), .ZN(n13167) );
  AND2_X1 U7898 ( .A1(n14010), .A2(n13875), .ZN(n6871) );
  XNOR2_X1 U7899 ( .A(n14010), .B(n13207), .ZN(n13867) );
  OR2_X1 U7900 ( .A1(n7079), .A2(n11751), .ZN(n7588) );
  OAI21_X1 U7901 ( .B1(n14083), .B2(n6752), .A(n6898), .ZN(n6897) );
  NAND2_X1 U7902 ( .A1(n14083), .A2(n12111), .ZN(n6898) );
  AND2_X1 U7903 ( .A1(n14083), .A2(n7429), .ZN(n7428) );
  OR2_X1 U7904 ( .A1(n14209), .A2(n7430), .ZN(n7429) );
  NAND2_X1 U7905 ( .A1(n11906), .A2(n11905), .ZN(n14852) );
  INV_X1 U7906 ( .A(n14848), .ZN(n11906) );
  INV_X1 U7907 ( .A(n8455), .ZN(n8803) );
  XNOR2_X1 U7908 ( .A(n14561), .B(n12129), .ZN(n11970) );
  NOR2_X1 U7909 ( .A1(n9094), .A2(n6936), .ZN(n6935) );
  INV_X1 U7910 ( .A(n8846), .ZN(n6936) );
  NAND2_X1 U7911 ( .A1(n14580), .A2(n8843), .ZN(n14382) );
  NAND2_X1 U7912 ( .A1(n14382), .A2(n14381), .ZN(n14380) );
  XNOR2_X1 U7913 ( .A(n14572), .B(n14086), .ZN(n14381) );
  INV_X1 U7914 ( .A(n14454), .ZN(n6969) );
  INV_X1 U7915 ( .A(n7488), .ZN(n7487) );
  OAI21_X1 U7916 ( .B1(n7489), .B2(n8566), .A(n8583), .ZN(n7488) );
  AND2_X1 U7917 ( .A1(n10092), .A2(n12005), .ZN(n14540) );
  XNOR2_X1 U7918 ( .A(n8710), .B(n8700), .ZN(n11941) );
  OR2_X1 U7919 ( .A1(n14691), .A2(n7264), .ZN(n6920) );
  NAND2_X1 U7920 ( .A1(n8780), .A2(n8779), .ZN(n12132) );
  OR2_X1 U7921 ( .A1(n12030), .A2(n12029), .ZN(n12031) );
  OAI21_X1 U7922 ( .B1(n14219), .B2(n7411), .A(n7409), .ZN(n6873) );
  OR2_X1 U7923 ( .A1(n14354), .A2(n14353), .ZN(n14569) );
  INV_X1 U7924 ( .A(n9361), .ZN(n9359) );
  NAND2_X1 U7925 ( .A1(n9372), .A2(n9373), .ZN(n14891) );
  INV_X1 U7926 ( .A(n6932), .ZN(n6929) );
  NAND2_X1 U7927 ( .A1(n14887), .A2(n6931), .ZN(n6930) );
  INV_X1 U7928 ( .A(n12985), .ZN(n7368) );
  INV_X1 U7929 ( .A(n13010), .ZN(n7349) );
  NOR2_X1 U7930 ( .A1(n8955), .A2(n7230), .ZN(n7229) );
  NOR2_X1 U7931 ( .A1(n8958), .A2(n8957), .ZN(n7231) );
  INV_X1 U7932 ( .A(n13049), .ZN(n7351) );
  NAND2_X1 U7933 ( .A1(n7016), .A2(n7015), .ZN(n7014) );
  NAND2_X1 U7934 ( .A1(n7020), .A2(n7017), .ZN(n7016) );
  INV_X1 U7935 ( .A(n8158), .ZN(n7015) );
  NAND2_X1 U7936 ( .A1(n7354), .A2(n13103), .ZN(n7353) );
  NAND2_X1 U7937 ( .A1(n7061), .A2(n7059), .ZN(n7058) );
  NAND2_X1 U7938 ( .A1(n6802), .A2(n6708), .ZN(n7061) );
  NAND2_X1 U7939 ( .A1(n6709), .A2(n6798), .ZN(n7059) );
  NAND2_X1 U7940 ( .A1(n7063), .A2(n6799), .ZN(n7057) );
  NAND2_X1 U7941 ( .A1(n6793), .A2(n6708), .ZN(n7062) );
  NAND2_X1 U7942 ( .A1(n6801), .A2(n6709), .ZN(n7060) );
  NAND2_X1 U7943 ( .A1(n8212), .A2(n8211), .ZN(n7063) );
  INV_X1 U7944 ( .A(n8228), .ZN(n7052) );
  INV_X1 U7945 ( .A(n13142), .ZN(n7347) );
  INV_X1 U7946 ( .A(n8247), .ZN(n7038) );
  NAND2_X1 U7947 ( .A1(n7277), .A2(n8839), .ZN(n6945) );
  INV_X1 U7948 ( .A(n7045), .ZN(n7044) );
  INV_X1 U7949 ( .A(n7035), .ZN(n7034) );
  INV_X1 U7950 ( .A(n7159), .ZN(n7158) );
  OAI21_X1 U7951 ( .B1(n7940), .B2(n7160), .A(n7955), .ZN(n7159) );
  INV_X1 U7952 ( .A(n7942), .ZN(n7160) );
  INV_X1 U7953 ( .A(n7497), .ZN(n7496) );
  OAI22_X1 U7954 ( .A1(n14381), .A2(n8744), .B1(n14361), .B2(n14379), .ZN(
        n7497) );
  INV_X1 U7955 ( .A(n14427), .ZN(n7486) );
  INV_X1 U7956 ( .A(n7509), .ZN(n7504) );
  NAND2_X1 U7957 ( .A1(n14249), .A2(n10794), .ZN(n7509) );
  INV_X1 U7958 ( .A(n14462), .ZN(n7477) );
  INV_X1 U7959 ( .A(n8673), .ZN(n7482) );
  AOI21_X1 U7960 ( .B1(n6965), .B2(n8341), .A(n6964), .ZN(n6963) );
  INV_X1 U7961 ( .A(n7596), .ZN(n6964) );
  INV_X1 U7962 ( .A(n6967), .ZN(n6965) );
  INV_X1 U7963 ( .A(n8341), .ZN(n6966) );
  AOI21_X1 U7964 ( .B1(n8477), .B2(n8330), .A(n8490), .ZN(n7559) );
  INV_X1 U7965 ( .A(n8330), .ZN(n7560) );
  OAI21_X1 U7966 ( .B1(n8322), .B2(n7134), .A(n8325), .ZN(n7132) );
  INV_X1 U7967 ( .A(n8465), .ZN(n8325) );
  NOR2_X1 U7968 ( .A1(n7134), .A2(n6942), .ZN(n6941) );
  INV_X1 U7969 ( .A(n8320), .ZN(n6942) );
  NAND2_X1 U7970 ( .A1(n8435), .A2(n8318), .ZN(n8321) );
  INV_X1 U7971 ( .A(n8434), .ZN(n8318) );
  INV_X1 U7972 ( .A(n8313), .ZN(n7515) );
  INV_X1 U7973 ( .A(n7392), .ZN(n7390) );
  AOI21_X1 U7974 ( .B1(n7392), .B2(n7389), .A(n7388), .ZN(n7387) );
  AOI21_X1 U7975 ( .B1(P3_REG1_REG_2__SCAN_IN), .B2(n10115), .A(n10106), .ZN(
        n10041) );
  INV_X1 U7976 ( .A(n8250), .ZN(n7467) );
  INV_X1 U7977 ( .A(n7462), .ZN(n7461) );
  INV_X1 U7978 ( .A(n8249), .ZN(n7457) );
  INV_X1 U7979 ( .A(n7466), .ZN(n12444) );
  OR2_X1 U7980 ( .A1(n12492), .A2(n12203), .ZN(n8237) );
  INV_X1 U7981 ( .A(n8227), .ZN(n7447) );
  INV_X1 U7982 ( .A(n7448), .ZN(n6999) );
  INV_X1 U7983 ( .A(n8226), .ZN(n6998) );
  NOR2_X1 U7984 ( .A1(n12521), .A2(n7452), .ZN(n7451) );
  INV_X1 U7985 ( .A(n8219), .ZN(n7452) );
  AOI21_X1 U7986 ( .B1(n11707), .B2(n7202), .A(n6743), .ZN(n7201) );
  OR2_X1 U7987 ( .A1(n12711), .A2(n12235), .ZN(n8200) );
  AOI21_X1 U7988 ( .B1(n7443), .B2(n8168), .A(n10865), .ZN(n6994) );
  NOR2_X1 U7989 ( .A1(n10722), .A2(n7445), .ZN(n7442) );
  NAND2_X1 U7990 ( .A1(n11077), .A2(n7444), .ZN(n7443) );
  OR2_X1 U7991 ( .A1(n10728), .A2(n7445), .ZN(n7444) );
  AOI21_X1 U7992 ( .B1(n10442), .B2(n7213), .A(n6760), .ZN(n7212) );
  INV_X1 U7993 ( .A(n10438), .ZN(n7213) );
  NAND2_X1 U7994 ( .A1(n6989), .A2(n9157), .ZN(n15350) );
  INV_X1 U7995 ( .A(n7165), .ZN(n7164) );
  OAI21_X1 U7996 ( .B1(n7878), .B2(n7166), .A(n7892), .ZN(n7165) );
  INV_X1 U7997 ( .A(n7880), .ZN(n7166) );
  INV_X1 U7998 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n8305) );
  NAND2_X1 U7999 ( .A1(n9918), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7677) );
  NAND2_X1 U8000 ( .A1(n7321), .A2(n12878), .ZN(n7320) );
  NAND2_X1 U8001 ( .A1(n7322), .A2(n7325), .ZN(n7321) );
  NOR2_X1 U8002 ( .A1(n12960), .A2(n7339), .ZN(n7338) );
  INV_X1 U8003 ( .A(n12827), .ZN(n7339) );
  OR2_X1 U8004 ( .A1(n13980), .A2(n13358), .ZN(n13374) );
  NAND2_X1 U8005 ( .A1(n13884), .A2(n13891), .ZN(n7578) );
  NOR2_X1 U8006 ( .A1(n14030), .A2(n13906), .ZN(n7566) );
  AND2_X1 U8007 ( .A1(n14030), .A2(n13363), .ZN(n7553) );
  OAI22_X1 U8008 ( .A1(n11582), .A2(n11595), .B1(n13264), .B2(n13064), .ZN(
        n11738) );
  NAND2_X1 U8009 ( .A1(n15131), .A2(n13271), .ZN(n7530) );
  AND2_X1 U8010 ( .A1(n10847), .A2(n13013), .ZN(n7531) );
  OR2_X1 U8011 ( .A1(n13013), .A2(n13009), .ZN(n7077) );
  OR2_X1 U8012 ( .A1(n14830), .A2(n13266), .ZN(n6870) );
  NOR2_X1 U8013 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n7342) );
  NOR2_X1 U8014 ( .A1(n7412), .A2(n6881), .ZN(n6880) );
  INV_X1 U8015 ( .A(n6885), .ZN(n6881) );
  OR2_X1 U8016 ( .A1(n12090), .A2(n14163), .ZN(n12095) );
  NOR2_X1 U8017 ( .A1(n12096), .A2(n6907), .ZN(n6906) );
  INV_X1 U8018 ( .A(n12060), .ZN(n6907) );
  OR2_X1 U8019 ( .A1(n14162), .A2(n12090), .ZN(n12096) );
  NAND2_X1 U8020 ( .A1(n14090), .A2(n12017), .ZN(n12023) );
  INV_X1 U8021 ( .A(n14241), .ZN(n11912) );
  NAND2_X1 U8022 ( .A1(n11135), .A2(n10255), .ZN(n8423) );
  NAND2_X1 U8023 ( .A1(n6822), .A2(n6821), .ZN(n8813) );
  INV_X1 U8024 ( .A(n14125), .ZN(n6821) );
  INV_X1 U8025 ( .A(n10246), .ZN(n6822) );
  NAND2_X1 U8026 ( .A1(n11138), .A2(n11137), .ZN(n11136) );
  OAI21_X1 U8027 ( .B1(n8686), .B2(n8376), .A(n8375), .ZN(n8710) );
  NAND2_X1 U8028 ( .A1(n7597), .A2(n7600), .ZN(n8376) );
  NAND2_X1 U8029 ( .A1(n7150), .A2(n8373), .ZN(n8686) );
  NAND2_X1 U8030 ( .A1(n8656), .A2(n8655), .ZN(n7150) );
  AND2_X1 U8031 ( .A1(n8366), .A2(n8365), .ZN(n8631) );
  AND2_X1 U8032 ( .A1(n8360), .A2(n8359), .ZN(n8618) );
  OAI21_X1 U8033 ( .B1(n8568), .B2(n8348), .A(n8347), .ZN(n8596) );
  INV_X1 U8034 ( .A(n8567), .ZN(n8348) );
  OR2_X1 U8035 ( .A1(n8492), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n8507) );
  INV_X1 U8036 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9288) );
  NAND2_X1 U8037 ( .A1(n9305), .A2(n9304), .ZN(n9358) );
  INV_X1 U8038 ( .A(n9219), .ZN(n7386) );
  AND2_X1 U8039 ( .A1(n9228), .A2(n9227), .ZN(n12165) );
  INV_X1 U8040 ( .A(n9224), .ZN(n12166) );
  OR2_X1 U8041 ( .A1(n8020), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8033) );
  XNOR2_X1 U8042 ( .A(n9165), .B(n15200), .ZN(n9168) );
  NAND2_X1 U8043 ( .A1(n15194), .A2(n6742), .ZN(n10484) );
  NOR2_X1 U8044 ( .A1(P3_REG3_REG_25__SCAN_IN), .A2(n8033), .ZN(n8046) );
  NAND2_X1 U8045 ( .A1(n6834), .A2(n7180), .ZN(n6833) );
  XNOR2_X1 U8046 ( .A(n7175), .B(n9145), .ZN(n8145) );
  AND2_X1 U8047 ( .A1(n7177), .A2(n8131), .ZN(n7176) );
  NOR2_X1 U8048 ( .A1(n12408), .A2(n7178), .ZN(n7177) );
  NAND2_X1 U8049 ( .A1(n10059), .A2(n10058), .ZN(n15224) );
  OR2_X1 U8050 ( .A1(n10057), .A2(n10056), .ZN(n10058) );
  INV_X1 U8051 ( .A(n11053), .ZN(n7246) );
  NAND2_X1 U8052 ( .A1(n12318), .A2(n12319), .ZN(n6845) );
  NOR2_X1 U8053 ( .A1(n12304), .A2(n12305), .ZN(n14747) );
  INV_X1 U8054 ( .A(n7248), .ZN(n12302) );
  OR2_X1 U8055 ( .A1(n14747), .A2(n14746), .ZN(n7254) );
  NAND2_X1 U8056 ( .A1(n7997), .A2(n8230), .ZN(n12491) );
  INV_X1 U8057 ( .A(n7451), .ZN(n7450) );
  OR2_X1 U8058 ( .A1(n12508), .A2(n12513), .ZN(n12510) );
  NOR2_X1 U8059 ( .A1(n8217), .A2(n7455), .ZN(n7454) );
  OR2_X1 U8060 ( .A1(n12560), .A2(n12534), .ZN(n8207) );
  AND4_X1 U8061 ( .A1(n7923), .A2(n7922), .A3(n7921), .A4(n7920), .ZN(n12552)
         );
  AND3_X1 U8062 ( .A1(n7954), .A2(n7953), .A3(n7952), .ZN(n12553) );
  NAND2_X1 U8063 ( .A1(n7197), .A2(n7203), .ZN(n7195) );
  AND2_X1 U8064 ( .A1(n8207), .A2(n8213), .ZN(n12550) );
  AOI21_X1 U8065 ( .B1(n7003), .B2(n11568), .A(n6735), .ZN(n7001) );
  INV_X1 U8066 ( .A(n7003), .ZN(n7002) );
  CLKBUF_X1 U8067 ( .A(n11569), .Z(n6847) );
  NAND2_X1 U8068 ( .A1(n15417), .A2(n7827), .ZN(n11353) );
  NAND2_X1 U8069 ( .A1(n10722), .A2(n10728), .ZN(n10721) );
  NAND2_X1 U8070 ( .A1(n15337), .A2(n10438), .ZN(n10443) );
  OR2_X1 U8071 ( .A1(n7674), .A2(n9521), .ZN(n7648) );
  INV_X1 U8072 ( .A(n11952), .ZN(n10542) );
  NAND2_X1 U8073 ( .A1(n7988), .A2(n7987), .ZN(n12387) );
  NAND2_X1 U8074 ( .A1(n9267), .A2(n9260), .ZN(n15351) );
  NAND2_X1 U8075 ( .A1(n9153), .A2(n9152), .ZN(n10453) );
  OAI21_X1 U8076 ( .B1(n8078), .B2(n8077), .A(n8079), .ZN(n8081) );
  NAND2_X1 U8077 ( .A1(n8261), .A2(n7369), .ZN(n8273) );
  NOR2_X1 U8078 ( .A1(P3_IR_REG_23__SCAN_IN), .A2(P3_IR_REG_24__SCAN_IN), .ZN(
        n7369) );
  NOR2_X1 U8079 ( .A1(n7984), .A2(n7186), .ZN(n7185) );
  INV_X1 U8080 ( .A(n7981), .ZN(n7186) );
  AND2_X1 U8081 ( .A1(n8120), .A2(n7402), .ZN(n7403) );
  NOR2_X1 U8082 ( .A1(n8118), .A2(n8267), .ZN(n8119) );
  INV_X1 U8083 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8118) );
  INV_X1 U8084 ( .A(n8146), .ZN(n8123) );
  NAND2_X1 U8085 ( .A1(n7966), .A2(n11293), .ZN(n7969) );
  NAND2_X1 U8086 ( .A1(n7807), .A2(n7806), .ZN(n7815) );
  INV_X1 U8087 ( .A(n7171), .ZN(n7170) );
  OAI21_X1 U8088 ( .B1(n7173), .B2(n7172), .A(n7768), .ZN(n7171) );
  INV_X1 U8089 ( .A(n7765), .ZN(n7172) );
  AND2_X1 U8090 ( .A1(n7731), .A2(n7712), .ZN(n7729) );
  INV_X1 U8091 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7696) );
  AND2_X1 U8092 ( .A1(n7710), .A2(n7692), .ZN(n7708) );
  INV_X1 U8093 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n7693) );
  NAND2_X1 U8094 ( .A1(n9795), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7664) );
  NOR2_X1 U8095 ( .A1(n10572), .A2(n10400), .ZN(n7315) );
  INV_X1 U8096 ( .A(n10571), .ZN(n7318) );
  INV_X1 U8097 ( .A(n12843), .ZN(n7337) );
  INV_X1 U8098 ( .A(n12800), .ZN(n12801) );
  NAND2_X1 U8099 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(n12801), .ZN(n12817) );
  INV_X1 U8100 ( .A(n13875), .ZN(n13207) );
  NAND2_X1 U8101 ( .A1(n11839), .A2(n11840), .ZN(n11866) );
  OR2_X1 U8102 ( .A1(n11546), .A2(n11545), .ZN(n11556) );
  NAND2_X1 U8103 ( .A1(n6728), .A2(n7131), .ZN(n7130) );
  NAND2_X1 U8104 ( .A1(n13246), .A2(n6616), .ZN(n7131) );
  NAND2_X1 U8105 ( .A1(n13234), .A2(n13233), .ZN(n13241) );
  AOI21_X1 U8106 ( .B1(n13227), .B2(n13226), .A(n13225), .ZN(n13243) );
  NAND2_X1 U8107 ( .A1(n13218), .A2(n7126), .ZN(n13247) );
  AND2_X1 U8108 ( .A1(n13217), .A2(n7127), .ZN(n7126) );
  NAND2_X1 U8109 ( .A1(n7128), .A2(n13214), .ZN(n7127) );
  INV_X1 U8110 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6985) );
  BUF_X1 U8111 ( .A(n12775), .Z(n12903) );
  OR2_X1 U8113 ( .A1(n10407), .A2(n9923), .ZN(n9924) );
  NAND2_X1 U8114 ( .A1(n13403), .A2(n6692), .ZN(n13345) );
  INV_X1 U8115 ( .A(n13356), .ZN(n13790) );
  AOI21_X1 U8116 ( .B1(n6975), .B2(n6974), .A(n6764), .ZN(n6973) );
  INV_X1 U8117 ( .A(n6979), .ZN(n6974) );
  NAND2_X1 U8118 ( .A1(n13835), .A2(n6981), .ZN(n6978) );
  NOR2_X1 U8119 ( .A1(n13371), .A2(n6980), .ZN(n6979) );
  INV_X1 U8120 ( .A(n7582), .ZN(n6980) );
  AND2_X1 U8121 ( .A1(n7570), .A2(n7571), .ZN(n7567) );
  NAND2_X1 U8122 ( .A1(n13850), .A2(n13368), .ZN(n7570) );
  OR2_X1 U8123 ( .A1(n13884), .A2(n13365), .ZN(n7583) );
  OR2_X1 U8124 ( .A1(n7070), .A2(n13352), .ZN(n7584) );
  NOR2_X1 U8125 ( .A1(n13878), .A2(n7577), .ZN(n7576) );
  INV_X1 U8126 ( .A(n7584), .ZN(n7577) );
  OR2_X1 U8127 ( .A1(n13916), .A2(n13929), .ZN(n7586) );
  NAND2_X1 U8128 ( .A1(n13894), .A2(n13893), .ZN(n13892) );
  INV_X1 U8129 ( .A(n13351), .ZN(n13893) );
  OR2_X1 U8130 ( .A1(n13349), .A2(n13927), .ZN(n7587) );
  NOR2_X1 U8131 ( .A1(n13940), .A2(n7565), .ZN(n7564) );
  INV_X1 U8132 ( .A(n7587), .ZN(n7565) );
  INV_X1 U8133 ( .A(n13923), .ZN(n13940) );
  NAND2_X1 U8134 ( .A1(n6769), .A2(n13360), .ZN(n7549) );
  INV_X1 U8135 ( .A(n13361), .ZN(n7550) );
  NAND2_X1 U8136 ( .A1(n11754), .A2(n11753), .ZN(n13350) );
  AND2_X1 U8137 ( .A1(n7081), .A2(n13066), .ZN(n6982) );
  OR2_X1 U8138 ( .A1(n7081), .A2(n13265), .ZN(n6861) );
  NOR2_X1 U8139 ( .A1(n10527), .A2(n13009), .ZN(n10692) );
  NAND2_X1 U8140 ( .A1(n10512), .A2(n13191), .ZN(n10688) );
  INV_X1 U8141 ( .A(n10513), .ZN(n10514) );
  NAND2_X1 U8142 ( .A1(n13185), .A2(n10321), .ZN(n10322) );
  OR2_X1 U8143 ( .A1(n9943), .A2(n9786), .ZN(n14784) );
  OR2_X1 U8144 ( .A1(n9750), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n9752) );
  OR2_X1 U8145 ( .A1(n9752), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n10283) );
  NAND2_X1 U8146 ( .A1(n12013), .A2(n7432), .ZN(n14090) );
  NOR2_X1 U8147 ( .A1(n14093), .A2(n7433), .ZN(n7432) );
  INV_X1 U8148 ( .A(n12012), .ZN(n7433) );
  AND2_X1 U8149 ( .A1(n14187), .A2(n12083), .ZN(n14104) );
  AOI21_X1 U8150 ( .B1(n7428), .B2(n7430), .A(n6748), .ZN(n7427) );
  NAND2_X1 U8151 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n8739), .ZN(n8753) );
  AND2_X1 U8152 ( .A1(n10936), .A2(n10935), .ZN(n10946) );
  OR2_X1 U8153 ( .A1(n9430), .A2(n8410), .ZN(n6869) );
  INV_X1 U8154 ( .A(n14200), .ZN(n7437) );
  NOR2_X1 U8155 ( .A1(n14117), .A2(n7440), .ZN(n7439) );
  INV_X1 U8156 ( .A(n12045), .ZN(n7440) );
  NOR2_X1 U8157 ( .A1(n8694), .A2(n14132), .ZN(n8702) );
  NAND2_X1 U8158 ( .A1(n8702), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8719) );
  INV_X1 U8159 ( .A(n10248), .ZN(n10254) );
  NAND2_X1 U8160 ( .A1(n6683), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n8404) );
  OR3_X1 U8161 ( .A1(n8875), .A2(n11515), .A3(n11726), .ZN(n10367) );
  OR2_X1 U8162 ( .A1(n14279), .A2(n14278), .ZN(n7089) );
  NAND2_X1 U8163 ( .A1(n9081), .A2(n9080), .ZN(n14342) );
  NAND2_X1 U8164 ( .A1(n9059), .A2(n9058), .ZN(n14345) );
  OR2_X1 U8165 ( .A1(n14388), .A2(n14389), .ZN(n14386) );
  NAND2_X1 U8166 ( .A1(n8717), .A2(n8716), .ZN(n14423) );
  NAND2_X1 U8167 ( .A1(n6694), .A2(n8838), .ZN(n6952) );
  NOR2_X1 U8168 ( .A1(n6947), .A2(n7277), .ZN(n6951) );
  NOR2_X1 U8169 ( .A1(n14453), .A2(n7278), .ZN(n6947) );
  XNOR2_X1 U8170 ( .A(n6970), .B(n14237), .ZN(n14462) );
  AND2_X1 U8171 ( .A1(n7281), .A2(n7279), .ZN(n14473) );
  NOR2_X1 U8172 ( .A1(n6696), .A2(n6756), .ZN(n7279) );
  OR2_X1 U8173 ( .A1(n14494), .A2(n14495), .ZN(n7483) );
  AND2_X1 U8174 ( .A1(n8992), .A2(n8654), .ZN(n14516) );
  OR2_X1 U8175 ( .A1(n11886), .A2(n11887), .ZN(n11891) );
  AND2_X1 U8176 ( .A1(n8960), .A2(n8972), .ZN(n11821) );
  NOR2_X1 U8177 ( .A1(n11611), .A2(n7298), .ZN(n7297) );
  INV_X1 U8178 ( .A(n8826), .ZN(n7298) );
  NAND2_X1 U8179 ( .A1(n8576), .A2(n8575), .ZN(n11928) );
  OR2_X1 U8180 ( .A1(n14707), .A2(n11912), .ZN(n8566) );
  INV_X1 U8181 ( .A(n9104), .ZN(n11460) );
  NAND2_X1 U8182 ( .A1(n8554), .A2(n8948), .ZN(n14698) );
  OR2_X1 U8183 ( .A1(n11385), .A2(n8953), .ZN(n8554) );
  INV_X1 U8184 ( .A(n7295), .ZN(n7294) );
  NAND2_X1 U8185 ( .A1(n11196), .A2(n8852), .ZN(n14710) );
  AND2_X1 U8186 ( .A1(n9103), .A2(n8523), .ZN(n7501) );
  NAND2_X1 U8187 ( .A1(n8522), .A2(n8521), .ZN(n11112) );
  AOI21_X1 U8188 ( .B1(n10617), .B2(n8814), .A(n7602), .ZN(n10780) );
  NOR2_X1 U8189 ( .A1(n7506), .A2(n10809), .ZN(n7602) );
  INV_X1 U8190 ( .A(n7108), .ZN(n6827) );
  AOI21_X1 U8191 ( .B1(n14561), .B2(n14963), .A(n14560), .ZN(n7108) );
  NAND2_X1 U8192 ( .A1(n8607), .A2(n8606), .ZN(n14634) );
  NAND2_X1 U8193 ( .A1(n9051), .A2(n7117), .ZN(n7119) );
  NAND2_X1 U8194 ( .A1(n7118), .A2(n7112), .ZN(n7111) );
  NOR2_X1 U8195 ( .A1(n7120), .A2(n9042), .ZN(n7112) );
  AND2_X1 U8196 ( .A1(n7122), .A2(n7116), .ZN(n7115) );
  AND2_X1 U8197 ( .A1(n9054), .A2(n6803), .ZN(n7122) );
  NAND2_X1 U8198 ( .A1(n9051), .A2(n7117), .ZN(n7116) );
  NAND2_X1 U8199 ( .A1(n8387), .A2(n6908), .ZN(n8384) );
  NOR2_X1 U8200 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n6908) );
  NAND2_X1 U8201 ( .A1(n7141), .A2(n6710), .ZN(n8775) );
  NAND2_X1 U8202 ( .A1(n8387), .A2(n8288), .ZN(n8389) );
  AOI22_X1 U8203 ( .A1(n7146), .A2(n7144), .B1(n7147), .B2(n7143), .ZN(n7142)
         );
  INV_X1 U8204 ( .A(n8745), .ZN(n7144) );
  INV_X1 U8205 ( .A(n7149), .ZN(n7143) );
  OR2_X1 U8206 ( .A1(n8747), .A2(n7145), .ZN(n7141) );
  NOR2_X1 U8207 ( .A1(n7146), .A2(n7147), .ZN(n7145) );
  AND2_X1 U8208 ( .A1(n8573), .A2(n7240), .ZN(n8859) );
  AND2_X1 U8209 ( .A1(n8797), .A2(n6773), .ZN(n7240) );
  INV_X1 U8210 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n7241) );
  NAND2_X1 U8211 ( .A1(n8369), .A2(n6957), .ZN(n8643) );
  NAND2_X1 U8212 ( .A1(n6962), .A2(n8341), .ZN(n8555) );
  NAND2_X1 U8213 ( .A1(n7151), .A2(n6967), .ZN(n6962) );
  INV_X1 U8214 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n7474) );
  INV_X1 U8215 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n7472) );
  INV_X1 U8216 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7473) );
  XNOR2_X1 U8217 ( .A(n8394), .B(P1_IR_REG_1__SCAN_IN), .ZN(n9458) );
  NOR2_X1 U8218 ( .A1(n9293), .A2(n9292), .ZN(n9342) );
  OAI21_X1 U8219 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n9298), .A(n9297), .ZN(
        n9352) );
  XNOR2_X1 U8220 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(n9301), .ZN(n9322) );
  NOR2_X1 U8221 ( .A1(n9367), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n7267) );
  INV_X1 U8222 ( .A(n9362), .ZN(n7269) );
  AND2_X1 U8223 ( .A1(n14886), .A2(n6933), .ZN(n6932) );
  AND3_X1 U8224 ( .A1(n7756), .A2(n7755), .A3(n7754), .ZN(n11089) );
  NAND2_X1 U8225 ( .A1(n7377), .A2(n9203), .ZN(n11688) );
  OR2_X1 U8226 ( .A1(n11509), .A2(n9204), .ZN(n7377) );
  NOR2_X1 U8227 ( .A1(n7373), .A2(n6702), .ZN(n7370) );
  NAND2_X1 U8228 ( .A1(n15196), .A2(n15195), .ZN(n15194) );
  AND4_X1 U8229 ( .A1(n8038), .A2(n8037), .A3(n8036), .A4(n8035), .ZN(n12448)
         );
  INV_X1 U8230 ( .A(n15193), .ZN(n15207) );
  NOR2_X1 U8231 ( .A1(n12276), .A2(n12275), .ZN(n12304) );
  XNOR2_X1 U8232 ( .A(n12418), .B(n12419), .ZN(n12588) );
  OR2_X1 U8233 ( .A1(n6691), .A2(n12417), .ZN(n12418) );
  NAND2_X1 U8234 ( .A1(n7464), .A2(n8245), .ZN(n12437) );
  OR2_X1 U8235 ( .A1(n11990), .A2(n7674), .ZN(n8084) );
  NOR2_X1 U8236 ( .A1(n6717), .A2(n12585), .ZN(n12655) );
  AOI21_X1 U8237 ( .B1(n12588), .B2(n14775), .A(n12589), .ZN(n12658) );
  NAND2_X1 U8238 ( .A1(n7948), .A2(n7947), .ZN(n12694) );
  NAND2_X1 U8239 ( .A1(n12707), .A2(n14770), .ZN(n12712) );
  INV_X2 U8240 ( .A(n15419), .ZN(n12707) );
  NAND2_X1 U8241 ( .A1(n12858), .A2(n12857), .ZN(n13985) );
  NAND2_X1 U8242 ( .A1(n12762), .A2(n12761), .ZN(n14016) );
  NAND2_X1 U8243 ( .A1(n12798), .A2(n12797), .ZN(n13999) );
  NAND2_X1 U8244 ( .A1(n12768), .A2(n12767), .ZN(n14010) );
  INV_X1 U8245 ( .A(n13263), .ZN(n11751) );
  OR2_X1 U8246 ( .A1(n9943), .A2(n9627), .ZN(n13928) );
  NAND2_X1 U8247 ( .A1(n13179), .A2(n13178), .ZN(n13966) );
  NAND2_X1 U8248 ( .A1(n7521), .A2(n15054), .ZN(n7520) );
  AOI21_X1 U8249 ( .B1(n7535), .B2(n7538), .A(n6767), .ZN(n7533) );
  XNOR2_X1 U8250 ( .A(n13402), .B(n13409), .ZN(n13988) );
  NAND2_X1 U8251 ( .A1(n7539), .A2(n6693), .ZN(n13402) );
  NOR2_X1 U8252 ( .A1(n6703), .A2(n14850), .ZN(n6894) );
  NAND2_X1 U8253 ( .A1(n6897), .A2(n6899), .ZN(n6896) );
  OR2_X1 U8254 ( .A1(n14083), .A2(n7430), .ZN(n6899) );
  AND4_X1 U8255 ( .A1(n8520), .A2(n8519), .A3(n8518), .A4(n8517), .ZN(n11681)
         );
  NAND2_X1 U8256 ( .A1(n8663), .A2(n8662), .ZN(n14616) );
  NAND2_X1 U8257 ( .A1(n14174), .A2(n12060), .ZN(n14102) );
  NAND2_X1 U8258 ( .A1(n8738), .A2(n8737), .ZN(n14578) );
  NAND2_X1 U8259 ( .A1(n8391), .A2(n8390), .ZN(n14585) );
  NAND2_X1 U8260 ( .A1(n11926), .A2(n11925), .ZN(n11931) );
  NAND2_X1 U8261 ( .A1(n6872), .A2(n12038), .ZN(n14199) );
  NAND2_X1 U8262 ( .A1(n14156), .A2(n14157), .ZN(n6872) );
  NAND2_X1 U8263 ( .A1(n8750), .A2(n8749), .ZN(n14572) );
  NAND2_X1 U8264 ( .A1(n12829), .A2(n6617), .ZN(n8750) );
  AND2_X1 U8265 ( .A1(n14844), .A2(n14963), .ZN(n14215) );
  NAND2_X1 U8266 ( .A1(n9875), .A2(n9874), .ZN(n9873) );
  XNOR2_X1 U8267 ( .A(n6937), .B(n11970), .ZN(n14564) );
  NAND2_X1 U8268 ( .A1(n6938), .A2(n6740), .ZN(n6937) );
  AOI21_X1 U8269 ( .B1(n14364), .B2(n8846), .A(n8790), .ZN(n8847) );
  INV_X1 U8270 ( .A(n6938), .ZN(n11964) );
  NAND2_X1 U8271 ( .A1(n8810), .A2(n8809), .ZN(n8811) );
  NAND2_X1 U8272 ( .A1(n14367), .A2(n14366), .ZN(n14566) );
  INV_X1 U8273 ( .A(n14365), .ZN(n14366) );
  NAND2_X1 U8274 ( .A1(n8763), .A2(n8762), .ZN(n14567) );
  NAND2_X1 U8275 ( .A1(n12856), .A2(n6617), .ZN(n8763) );
  NAND2_X1 U8276 ( .A1(n14673), .A2(n9430), .ZN(n14445) );
  AND2_X1 U8277 ( .A1(n6934), .A2(P2_ADDR_REG_1__SCAN_IN), .ZN(n9332) );
  INV_X1 U8278 ( .A(n14691), .ZN(n6921) );
  NAND2_X1 U8279 ( .A1(n6923), .A2(n6721), .ZN(n6922) );
  INV_X1 U8280 ( .A(n6919), .ZN(n6916) );
  AND2_X1 U8281 ( .A1(n6918), .A2(n6917), .ZN(n14694) );
  NOR2_X1 U8282 ( .A1(n14696), .A2(n6919), .ZN(n6917) );
  NAND2_X1 U8283 ( .A1(n14876), .A2(n9362), .ZN(n9366) );
  NAND2_X1 U8284 ( .A1(n14729), .A2(n9376), .ZN(n14677) );
  OR2_X1 U8285 ( .A1(n7361), .A2(n12998), .ZN(n7360) );
  INV_X1 U8286 ( .A(n12997), .ZN(n7361) );
  NAND2_X1 U8287 ( .A1(n8925), .A2(n8927), .ZN(n6867) );
  INV_X1 U8288 ( .A(n13023), .ZN(n7355) );
  NOR2_X1 U8289 ( .A1(n13026), .A2(n13023), .ZN(n7356) );
  NAND2_X1 U8290 ( .A1(n8942), .A2(n8944), .ZN(n7236) );
  NOR2_X1 U8291 ( .A1(n13039), .A2(n13036), .ZN(n7358) );
  INV_X1 U8292 ( .A(n13036), .ZN(n7357) );
  AOI21_X1 U8293 ( .B1(n8971), .B2(n8970), .A(n9082), .ZN(n8976) );
  OAI21_X1 U8294 ( .B1(n8956), .B2(n7231), .A(n7228), .ZN(n8967) );
  NAND2_X1 U8295 ( .A1(n15349), .A2(n7019), .ZN(n7018) );
  NAND2_X1 U8296 ( .A1(n10458), .A2(n8154), .ZN(n7019) );
  NAND2_X1 U8297 ( .A1(n8153), .A2(n9267), .ZN(n7020) );
  NAND2_X1 U8298 ( .A1(n7013), .A2(n7012), .ZN(n8160) );
  OR2_X1 U8299 ( .A1(n8159), .A2(n10458), .ZN(n7012) );
  NAND2_X1 U8300 ( .A1(n7014), .A2(n8157), .ZN(n7013) );
  NOR2_X1 U8301 ( .A1(n10865), .A2(n7068), .ZN(n7067) );
  NOR2_X1 U8302 ( .A1(n8172), .A2(n10458), .ZN(n7068) );
  INV_X1 U8303 ( .A(n8175), .ZN(n7065) );
  OAI22_X1 U8304 ( .A1(n13114), .A2(n7344), .B1(n13115), .B2(n7343), .ZN(
        n13120) );
  INV_X1 U8305 ( .A(n13113), .ZN(n7343) );
  NOR2_X1 U8306 ( .A1(n13116), .A2(n13113), .ZN(n7344) );
  OAI21_X1 U8307 ( .B1(n7069), .B2(n7066), .A(n7064), .ZN(n8181) );
  NOR2_X1 U8308 ( .A1(n7065), .A2(n11092), .ZN(n7064) );
  OAI21_X1 U8309 ( .B1(n8170), .B2(n10458), .A(n7067), .ZN(n7066) );
  AOI21_X1 U8310 ( .B1(n8169), .B2(n8168), .A(n9267), .ZN(n7069) );
  NAND2_X1 U8311 ( .A1(n9029), .A2(n9027), .ZN(n7233) );
  NAND2_X1 U8312 ( .A1(n7364), .A2(n13131), .ZN(n7363) );
  NAND2_X1 U8313 ( .A1(n7063), .A2(n6797), .ZN(n7056) );
  AND2_X1 U8314 ( .A1(n7051), .A2(n8232), .ZN(n7050) );
  NAND2_X1 U8315 ( .A1(n7054), .A2(n7052), .ZN(n7051) );
  AOI21_X1 U8316 ( .B1(n7050), .B2(n12503), .A(n12490), .ZN(n7049) );
  AOI21_X1 U8317 ( .B1(n7046), .B2(n7048), .A(n12478), .ZN(n7045) );
  INV_X1 U8318 ( .A(n7049), .ZN(n7048) );
  NOR2_X1 U8319 ( .A1(n8136), .A2(n7206), .ZN(n8137) );
  NAND2_X1 U8320 ( .A1(n11077), .A2(n7207), .ZN(n7206) );
  INV_X1 U8321 ( .A(n13141), .ZN(n7345) );
  NOR2_X1 U8322 ( .A1(n7347), .A2(n13141), .ZN(n7346) );
  INV_X1 U8323 ( .A(n7397), .ZN(n7389) );
  INV_X1 U8324 ( .A(n9215), .ZN(n7388) );
  AOI21_X1 U8325 ( .B1(n7045), .B2(n7043), .A(n12462), .ZN(n7042) );
  INV_X1 U8326 ( .A(n7046), .ZN(n7043) );
  NAND2_X1 U8327 ( .A1(n12243), .A2(n15343), .ZN(n8157) );
  NOR2_X1 U8328 ( .A1(P3_IR_REG_13__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), .ZN(
        n7607) );
  NAND2_X1 U8329 ( .A1(n13146), .A2(n13147), .ZN(n13145) );
  AND2_X1 U8330 ( .A1(n7139), .A2(n13212), .ZN(n7135) );
  AND2_X1 U8331 ( .A1(n13375), .A2(n13331), .ZN(n7139) );
  XNOR2_X1 U8332 ( .A(n13343), .B(n13377), .ZN(n7140) );
  INV_X1 U8333 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7641) );
  INV_X1 U8334 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7642) );
  INV_X1 U8335 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7639) );
  INV_X1 U8336 ( .A(n10084), .ZN(n10083) );
  NAND2_X1 U8337 ( .A1(n9040), .A2(n9039), .ZN(n9047) );
  OR2_X1 U8338 ( .A1(n14381), .A2(n14389), .ZN(n7498) );
  NOR2_X1 U8339 ( .A1(n6950), .A2(n7278), .ZN(n6949) );
  AOI21_X1 U8340 ( .B1(n6840), .B2(n6948), .A(n6944), .ZN(n6943) );
  NOR2_X1 U8341 ( .A1(n7278), .A2(n6950), .ZN(n6948) );
  NAND2_X1 U8342 ( .A1(n6766), .A2(n6945), .ZN(n6944) );
  INV_X1 U8343 ( .A(n9074), .ZN(n7113) );
  NAND2_X1 U8344 ( .A1(n8383), .A2(n8382), .ZN(n8730) );
  NAND2_X1 U8345 ( .A1(n8632), .A2(n8631), .ZN(n8367) );
  NAND2_X1 U8346 ( .A1(n8342), .A2(n9553), .ZN(n8345) );
  OAI21_X1 U8347 ( .B1(n9794), .B2(n9503), .A(n6830), .ZN(n8323) );
  NAND2_X1 U8348 ( .A1(n9794), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n6830) );
  NOR2_X1 U8349 ( .A1(n12190), .A2(n7398), .ZN(n7397) );
  INV_X1 U8350 ( .A(n12145), .ZN(n7398) );
  OR2_X1 U8351 ( .A1(n11728), .A2(n11727), .ZN(n9207) );
  NAND2_X1 U8352 ( .A1(n12199), .A2(n9218), .ZN(n9220) );
  OR2_X1 U8353 ( .A1(n8248), .A2(n7026), .ZN(n7025) );
  NOR2_X1 U8354 ( .A1(n7024), .A2(n7028), .ZN(n7023) );
  AND2_X1 U8355 ( .A1(n7029), .A2(n7033), .ZN(n7028) );
  NAND2_X1 U8356 ( .A1(n7031), .A2(n7034), .ZN(n7030) );
  NAND2_X1 U8357 ( .A1(n12419), .A2(n7179), .ZN(n7178) );
  AND2_X1 U8358 ( .A1(n8144), .A2(n7040), .ZN(n7179) );
  NAND2_X1 U8359 ( .A1(n15294), .A2(n15295), .ZN(n6842) );
  AOI21_X1 U8360 ( .B1(P3_REG1_REG_10__SCAN_IN), .B2(n11058), .A(n11057), .ZN(
        n11226) );
  NAND2_X1 U8361 ( .A1(n11471), .A2(n6866), .ZN(n12259) );
  OR2_X1 U8362 ( .A1(n11476), .A2(n13689), .ZN(n6866) );
  NAND2_X1 U8363 ( .A1(n12283), .A2(n12277), .ZN(n12316) );
  NAND2_X1 U8364 ( .A1(n6843), .A2(n14736), .ZN(n12321) );
  NAND2_X1 U8365 ( .A1(n6845), .A2(n6844), .ZN(n6843) );
  INV_X1 U8366 ( .A(n14742), .ZN(n6844) );
  NOR2_X1 U8367 ( .A1(n7989), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8009) );
  NOR2_X1 U8368 ( .A1(n12370), .A2(n7198), .ZN(n7197) );
  INV_X1 U8369 ( .A(n7201), .ZN(n7198) );
  OR2_X1 U8370 ( .A1(n12565), .A2(n12574), .ZN(n12370) );
  OR2_X1 U8371 ( .A1(n12574), .A2(n12567), .ZN(n12369) );
  OR2_X1 U8372 ( .A1(n11799), .A2(n11727), .ZN(n8201) );
  NOR2_X1 U8373 ( .A1(n8196), .A2(n7004), .ZN(n7003) );
  INV_X1 U8374 ( .A(n8192), .ZN(n7004) );
  INV_X1 U8375 ( .A(n11287), .ZN(n11325) );
  AND2_X1 U8376 ( .A1(n8161), .A2(n8157), .ZN(n15336) );
  NAND2_X1 U8377 ( .A1(n8017), .A2(n8016), .ZN(n8027) );
  INV_X1 U8378 ( .A(n7608), .ZN(n7469) );
  AOI21_X1 U8379 ( .B1(n7158), .B2(n7160), .A(n6811), .ZN(n7155) );
  INV_X1 U8380 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n8362) );
  NOR2_X2 U8381 ( .A1(n7896), .A2(P3_IR_REG_16__SCAN_IN), .ZN(n8121) );
  INV_X1 U8382 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n8356) );
  INV_X1 U8383 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n7750) );
  NAND2_X1 U8384 ( .A1(n9509), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n7731) );
  NAND2_X1 U8385 ( .A1(n9497), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7710) );
  NAND2_X1 U8386 ( .A1(n9476), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7691) );
  NOR2_X1 U8387 ( .A1(n10766), .A2(n10765), .ZN(n10884) );
  NOR2_X1 U8388 ( .A1(n11161), .A2(n11160), .ZN(n11309) );
  NAND2_X2 U8389 ( .A1(n10171), .A2(n13224), .ZN(n9932) );
  NOR2_X1 U8390 ( .A1(n11556), .A2(n11555), .ZN(n11587) );
  OR2_X1 U8391 ( .A1(n13966), .A2(n13180), .ZN(n13244) );
  INV_X1 U8392 ( .A(n12971), .ZN(n13224) );
  INV_X1 U8393 ( .A(n13219), .ZN(n7128) );
  NAND2_X1 U8394 ( .A1(n13375), .A2(n13374), .ZN(n7526) );
  INV_X1 U8395 ( .A(n13355), .ZN(n7542) );
  NAND2_X1 U8396 ( .A1(n13985), .A2(n13356), .ZN(n7543) );
  NOR2_X1 U8397 ( .A1(n7081), .A2(n13052), .ZN(n7080) );
  NOR2_X1 U8398 ( .A1(n10527), .A2(n7073), .ZN(n7072) );
  NAND2_X1 U8399 ( .A1(n15137), .A2(n7074), .ZN(n7073) );
  INV_X1 U8400 ( .A(n7077), .ZN(n7076) );
  NAND2_X1 U8401 ( .A1(n10508), .A2(n10507), .ZN(n10512) );
  NOR2_X1 U8402 ( .A1(n10133), .A2(n10132), .ZN(n10271) );
  NOR2_X1 U8403 ( .A1(n10476), .A2(n12988), .ZN(n10393) );
  NAND2_X1 U8404 ( .A1(n7071), .A2(n7070), .ZN(n13879) );
  NAND2_X1 U8405 ( .A1(n11414), .A2(n7078), .ZN(n11755) );
  AND2_X1 U8406 ( .A1(n6697), .A2(n7079), .ZN(n7078) );
  NAND2_X1 U8407 ( .A1(n13215), .A2(n10168), .ZN(n9793) );
  INV_X1 U8408 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7341) );
  OR2_X1 U8409 ( .A1(n9554), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n9594) );
  OR2_X1 U8410 ( .A1(n9531), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n9554) );
  NOR2_X1 U8411 ( .A1(n9506), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n9729) );
  NAND2_X1 U8412 ( .A1(n10948), .A2(n10947), .ZN(n7420) );
  NAND2_X1 U8413 ( .A1(n6887), .A2(n6886), .ZN(n6885) );
  INV_X1 U8414 ( .A(n10737), .ZN(n6886) );
  INV_X1 U8415 ( .A(n10736), .ZN(n6887) );
  NAND2_X1 U8416 ( .A1(n11643), .A2(n7092), .ZN(n11645) );
  OR2_X1 U8417 ( .A1(n11644), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7092) );
  NAND2_X1 U8418 ( .A1(n7495), .A2(n14358), .ZN(n7494) );
  INV_X1 U8419 ( .A(n7498), .ZN(n7495) );
  OR2_X1 U8420 ( .A1(n7496), .A2(n8845), .ZN(n7492) );
  NAND2_X1 U8421 ( .A1(n14394), .A2(n7103), .ZN(n7102) );
  NOR2_X1 U8422 ( .A1(n14585), .A2(n14423), .ZN(n7103) );
  AOI21_X1 U8423 ( .B1(n14448), .B2(n8708), .A(n7486), .ZN(n7485) );
  AND2_X1 U8424 ( .A1(n8837), .A2(n7286), .ZN(n7282) );
  INV_X1 U8425 ( .A(n7283), .ZN(n7280) );
  NOR2_X1 U8426 ( .A1(n14516), .A2(n7284), .ZN(n7283) );
  INV_X1 U8427 ( .A(n8982), .ZN(n7284) );
  NAND2_X1 U8428 ( .A1(n8833), .A2(n7286), .ZN(n7285) );
  NAND2_X1 U8429 ( .A1(n9104), .A2(n7490), .ZN(n7489) );
  NAND2_X1 U8430 ( .A1(n14709), .A2(n8566), .ZN(n7490) );
  NOR2_X1 U8431 ( .A1(n7296), .A2(n7293), .ZN(n7292) );
  INV_X1 U8432 ( .A(n8819), .ZN(n7293) );
  NOR2_X1 U8433 ( .A1(n11195), .A2(n14964), .ZN(n11196) );
  NOR2_X1 U8434 ( .A1(n10964), .A2(n14954), .ZN(n7106) );
  AND2_X1 U8435 ( .A1(n8816), .A2(n8476), .ZN(n10777) );
  AOI21_X1 U8436 ( .B1(n7505), .B2(n7504), .A(n6755), .ZN(n7502) );
  INV_X1 U8437 ( .A(n7505), .ZN(n7503) );
  NAND2_X1 U8438 ( .A1(n10939), .A2(n10746), .ZN(n7508) );
  NAND2_X1 U8439 ( .A1(n10621), .A2(n7509), .ZN(n7507) );
  NAND2_X1 U8440 ( .A1(n7100), .A2(n7099), .ZN(n10628) );
  INV_X1 U8441 ( .A(n10825), .ZN(n7100) );
  OAI21_X1 U8442 ( .B1(n14494), .B2(n7479), .A(n7476), .ZN(n14461) );
  AND2_X1 U8443 ( .A1(n8745), .A2(SI_26_), .ZN(n7149) );
  INV_X1 U8444 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8572) );
  NOR2_X1 U8445 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n7408) );
  NOR2_X1 U8446 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n8658) );
  NAND2_X1 U8447 ( .A1(n8367), .A2(n6958), .ZN(n6957) );
  AND2_X1 U8448 ( .A1(n8366), .A2(SI_18_), .ZN(n6958) );
  NAND2_X1 U8449 ( .A1(n8368), .A2(n10002), .ZN(n8369) );
  NAND2_X1 U8450 ( .A1(n8367), .A2(n8366), .ZN(n8368) );
  INV_X1 U8451 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8569) );
  NOR2_X1 U8452 ( .A1(n8336), .A2(n6968), .ZN(n6967) );
  INV_X1 U8453 ( .A(n8334), .ZN(n6968) );
  AOI21_X1 U8454 ( .B1(n8340), .B2(n8539), .A(n8339), .ZN(n8341) );
  NAND2_X1 U8455 ( .A1(n8337), .A2(SI_11_), .ZN(n8539) );
  NAND2_X1 U8456 ( .A1(n7151), .A2(n8334), .ZN(n8536) );
  XNOR2_X1 U8457 ( .A(n8536), .B(SI_10_), .ZN(n8534) );
  XNOR2_X1 U8458 ( .A(n8333), .B(SI_9_), .ZN(n8505) );
  AOI21_X1 U8459 ( .B1(n7559), .B2(n7560), .A(n6757), .ZN(n7556) );
  XNOR2_X1 U8460 ( .A(n8331), .B(SI_8_), .ZN(n8490) );
  OR2_X1 U8461 ( .A1(n8479), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n8492) );
  XNOR2_X1 U8462 ( .A(n8329), .B(SI_7_), .ZN(n8477) );
  OAI21_X1 U8463 ( .B1(n7132), .B2(n6836), .A(n8327), .ZN(n8478) );
  AND2_X1 U8464 ( .A1(n6941), .A2(n8321), .ZN(n6836) );
  NAND2_X1 U8465 ( .A1(n8323), .A2(SI_5_), .ZN(n8324) );
  INV_X1 U8466 ( .A(n8430), .ZN(n8314) );
  XNOR2_X1 U8467 ( .A(n6820), .B(P1_ADDR_REG_1__SCAN_IN), .ZN(n9329) );
  INV_X1 U8468 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n6820) );
  NOR2_X1 U8469 ( .A1(n9287), .A2(n6818), .ZN(n9289) );
  AND2_X1 U8470 ( .A1(n9288), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n6818) );
  NOR2_X1 U8471 ( .A1(n9290), .A2(n6835), .ZN(n9291) );
  AND2_X1 U8472 ( .A1(n14274), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n6835) );
  OR2_X1 U8473 ( .A1(n11507), .A2(n11709), .ZN(n9203) );
  AOI21_X1 U8474 ( .B1(n12220), .B2(n7382), .A(n9230), .ZN(n7381) );
  INV_X1 U8475 ( .A(n12220), .ZN(n7383) );
  INV_X1 U8476 ( .A(n9228), .ZN(n7382) );
  OAI21_X1 U8477 ( .B1(n12190), .B2(n7396), .A(n7400), .ZN(n7395) );
  NOR2_X1 U8478 ( .A1(n12155), .A2(n7395), .ZN(n7392) );
  NAND2_X1 U8479 ( .A1(n6850), .A2(n7397), .ZN(n7393) );
  AND2_X1 U8480 ( .A1(n9207), .A2(n6725), .ZN(n7375) );
  NOR2_X1 U8481 ( .A1(n7376), .A2(n7374), .ZN(n7373) );
  INV_X1 U8482 ( .A(n9207), .ZN(n7374) );
  NAND2_X1 U8483 ( .A1(n7900), .A2(n11857), .ZN(n7918) );
  NAND2_X1 U8484 ( .A1(n9212), .A2(n12233), .ZN(n7396) );
  NOR2_X1 U8486 ( .A1(n7854), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n7872) );
  OR2_X1 U8487 ( .A1(n7836), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7854) );
  NAND2_X1 U8488 ( .A1(n7795), .A2(n7794), .ZN(n7820) );
  NAND2_X1 U8489 ( .A1(n10564), .A2(n10563), .ZN(n7401) );
  OR2_X1 U8490 ( .A1(n7378), .A2(n9206), .ZN(n7376) );
  AOI21_X1 U8491 ( .B1(n9204), .B2(n9203), .A(n7379), .ZN(n7378) );
  INV_X1 U8492 ( .A(n11689), .ZN(n7379) );
  AND2_X1 U8493 ( .A1(n7885), .A2(n12279), .ZN(n7900) );
  AND4_X1 U8494 ( .A1(n8107), .A2(n8088), .A3(n8087), .A4(n8086), .ZN(n12232)
         );
  AND4_X1 U8495 ( .A1(n7651), .A2(n7652), .A3(n7653), .A4(n7650), .ZN(n15354)
         );
  NAND2_X1 U8496 ( .A1(n7666), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n7653) );
  OR2_X1 U8497 ( .A1(n10155), .A2(n10012), .ZN(n10157) );
  AND2_X1 U8498 ( .A1(n10146), .A2(n10039), .ZN(n10107) );
  NAND2_X1 U8499 ( .A1(n10040), .A2(n6741), .ZN(n15247) );
  NAND2_X1 U8500 ( .A1(n7258), .A2(n7257), .ZN(n7256) );
  AND2_X1 U8501 ( .A1(n7259), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7257) );
  NAND2_X1 U8502 ( .A1(n10060), .A2(n7259), .ZN(n7255) );
  NOR2_X1 U8503 ( .A1(n15224), .A2(n10022), .ZN(n15223) );
  OAI21_X1 U8504 ( .B1(n15276), .B2(n7252), .A(n7251), .ZN(n15299) );
  NAND2_X1 U8505 ( .A1(n7253), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7252) );
  NAND2_X1 U8506 ( .A1(n10641), .A2(n7253), .ZN(n7251) );
  INV_X1 U8507 ( .A(n15300), .ZN(n7253) );
  NOR2_X1 U8508 ( .A1(n11062), .A2(n11061), .ZN(n11064) );
  OR2_X1 U8509 ( .A1(n11467), .A2(n11466), .ZN(n11468) );
  XNOR2_X1 U8510 ( .A(n12259), .B(n12249), .ZN(n11472) );
  NOR2_X1 U8511 ( .A1(n12271), .A2(n7250), .ZN(n7249) );
  INV_X1 U8512 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n7250) );
  XOR2_X1 U8513 ( .A(n12316), .B(n12317), .Z(n12278) );
  INV_X1 U8514 ( .A(n7459), .ZN(n7458) );
  AOI21_X1 U8515 ( .B1(n7459), .B2(n7461), .A(n7457), .ZN(n7456) );
  AND2_X1 U8516 ( .A1(n7460), .A2(n7467), .ZN(n7459) );
  NOR2_X1 U8517 ( .A1(n12419), .A2(n7209), .ZN(n7208) );
  INV_X1 U8518 ( .A(n12400), .ZN(n7209) );
  NAND2_X1 U8519 ( .A1(n12480), .A2(n7053), .ZN(n12479) );
  AOI21_X1 U8520 ( .B1(n12513), .B2(n7219), .A(n7218), .ZN(n7217) );
  NOR2_X1 U8521 ( .A1(n12680), .A2(n12488), .ZN(n7218) );
  INV_X1 U8522 ( .A(n7446), .ZN(n7000) );
  AOI21_X1 U8523 ( .B1(n7446), .B2(n6999), .A(n6998), .ZN(n6997) );
  AOI21_X1 U8524 ( .B1(n7448), .B2(n7450), .A(n7447), .ZN(n7446) );
  AND2_X1 U8525 ( .A1(n7950), .A2(n7949), .ZN(n7959) );
  AND3_X1 U8526 ( .A1(n7937), .A2(n7936), .A3(n7935), .ZN(n12534) );
  OR2_X1 U8527 ( .A1(n12363), .A2(n6718), .ZN(n12565) );
  AND2_X1 U8528 ( .A1(n8206), .A2(n8204), .ZN(n11806) );
  NAND2_X1 U8529 ( .A1(n7199), .A2(n7201), .ZN(n12566) );
  NAND2_X1 U8530 ( .A1(n7200), .A2(n11707), .ZN(n7199) );
  NAND2_X1 U8531 ( .A1(n11770), .A2(n11769), .ZN(n11768) );
  OAI21_X1 U8532 ( .B1(n11244), .B2(n11325), .A(n11095), .ZN(n7793) );
  INV_X1 U8533 ( .A(n11329), .ZN(n11095) );
  AND4_X1 U8534 ( .A1(n7741), .A2(n7740), .A3(n7739), .A4(n7738), .ZN(n11094)
         );
  AND4_X1 U8535 ( .A1(n7762), .A2(n7761), .A3(n7760), .A4(n7759), .ZN(n11250)
         );
  NAND2_X1 U8536 ( .A1(n6996), .A2(n8168), .ZN(n10857) );
  OR2_X1 U8537 ( .A1(n7442), .A2(n7443), .ZN(n6996) );
  OR2_X1 U8538 ( .A1(n7721), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7736) );
  NOR2_X1 U8539 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n7702) );
  NAND2_X1 U8540 ( .A1(n7214), .A2(n10430), .ZN(n10429) );
  INV_X1 U8541 ( .A(n15336), .ZN(n15338) );
  AND2_X1 U8542 ( .A1(n10426), .A2(n10457), .ZN(n15373) );
  INV_X1 U8543 ( .A(n15351), .ZN(n15366) );
  AND2_X1 U8544 ( .A1(n9406), .A2(n9405), .ZN(n10540) );
  NAND2_X1 U8545 ( .A1(n8044), .A2(n8043), .ZN(n12398) );
  NAND2_X1 U8546 ( .A1(n8032), .A2(n8031), .ZN(n12396) );
  NAND2_X1 U8547 ( .A1(n8019), .A2(n8018), .ZN(n12392) );
  NAND2_X1 U8548 ( .A1(n7899), .A2(n7898), .ZN(n12365) );
  XNOR2_X1 U8549 ( .A(n8268), .B(P3_IR_REG_26__SCAN_IN), .ZN(n9232) );
  OAI21_X1 U8550 ( .B1(n8273), .B2(P3_IR_REG_25__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8268) );
  OR2_X1 U8551 ( .A1(n8027), .A2(n11448), .ZN(n8028) );
  NAND2_X1 U8552 ( .A1(n8026), .A2(n12136), .ZN(n8029) );
  NAND2_X1 U8553 ( .A1(n8261), .A2(n8260), .ZN(n8269) );
  XNOR2_X1 U8554 ( .A(n8027), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n8026) );
  OAI21_X1 U8555 ( .B1(n7980), .B2(n7184), .A(n7182), .ZN(n8004) );
  AOI21_X1 U8556 ( .B1(n7978), .B2(n7185), .A(n7183), .ZN(n7182) );
  INV_X1 U8557 ( .A(n7185), .ZN(n7184) );
  INV_X1 U8558 ( .A(n7998), .ZN(n7183) );
  NAND2_X1 U8559 ( .A1(n7162), .A2(n7161), .ZN(n7909) );
  AOI21_X1 U8560 ( .B1(n7164), .B2(n7166), .A(n6800), .ZN(n7161) );
  AND2_X1 U8561 ( .A1(n7803), .A2(n7782), .ZN(n7801) );
  OR2_X1 U8562 ( .A1(n7713), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n7715) );
  NOR2_X1 U8563 ( .A1(n7715), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n7751) );
  INV_X1 U8564 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7606) );
  NAND2_X1 U8565 ( .A1(n7645), .A2(n7644), .ZN(n7676) );
  AND2_X1 U8566 ( .A1(n7677), .A2(n7646), .ZN(n7675) );
  INV_X1 U8567 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10409) );
  INV_X1 U8568 ( .A(n11623), .ZN(n7330) );
  INV_X1 U8569 ( .A(n7331), .ZN(n7328) );
  AND2_X1 U8570 ( .A1(n11621), .A2(n11622), .ZN(n7333) );
  AND2_X1 U8571 ( .A1(n12781), .A2(n12780), .ZN(n12782) );
  OR2_X1 U8572 ( .A1(n12730), .A2(n11864), .ZN(n7325) );
  INV_X1 U8573 ( .A(n7323), .ZN(n7322) );
  OAI22_X1 U8574 ( .A1(n12730), .A2(n7324), .B1(n12728), .B2(n12729), .ZN(
        n7323) );
  OR2_X1 U8575 ( .A1(n11840), .A2(n11864), .ZN(n7324) );
  NAND2_X1 U8576 ( .A1(n7316), .A2(n7317), .ZN(n7311) );
  NAND2_X1 U8577 ( .A1(n7313), .A2(n7316), .ZN(n7310) );
  XNOR2_X1 U8578 ( .A(n9932), .B(n12979), .ZN(n7303) );
  OR2_X1 U8579 ( .A1(n10993), .A2(n10992), .ZN(n11161) );
  AND2_X1 U8580 ( .A1(n12929), .A2(n12873), .ZN(n7307) );
  NAND2_X1 U8581 ( .A1(n6828), .A2(n12793), .ZN(n12795) );
  INV_X1 U8582 ( .A(n12794), .ZN(n6828) );
  OR2_X1 U8583 ( .A1(n11871), .A2(n11870), .ZN(n12744) );
  NAND2_X1 U8584 ( .A1(n11307), .A2(n11423), .ZN(n7331) );
  NAND2_X1 U8585 ( .A1(n11299), .A2(n11423), .ZN(n7332) );
  NOR2_X1 U8586 ( .A1(n12771), .A2(n12952), .ZN(n12787) );
  INV_X1 U8587 ( .A(n12817), .ZN(n12815) );
  AND2_X1 U8588 ( .A1(n13244), .A2(n13239), .ZN(n13213) );
  AND4_X1 U8589 ( .A1(n12867), .A2(n12866), .A3(n12865), .A4(n12864), .ZN(
        n13358) );
  OR2_X1 U8590 ( .A1(n12901), .A2(n13796), .ZN(n12838) );
  OR2_X1 U8591 ( .A1(n12901), .A2(n13815), .ZN(n12821) );
  NOR2_X1 U8592 ( .A1(n6704), .A2(n13925), .ZN(n7519) );
  NAND2_X1 U8593 ( .A1(n7522), .A2(n7526), .ZN(n7521) );
  NOR2_X1 U8594 ( .A1(n6614), .A2(n7536), .ZN(n7535) );
  AND2_X1 U8595 ( .A1(n12894), .A2(n12893), .ZN(n13394) );
  NOR2_X1 U8596 ( .A1(n7540), .A2(n7537), .ZN(n7536) );
  INV_X1 U8597 ( .A(n7543), .ZN(n7537) );
  AND2_X1 U8598 ( .A1(n13409), .A2(n7541), .ZN(n7540) );
  NAND2_X1 U8599 ( .A1(n6693), .A2(n7542), .ZN(n7541) );
  NAND2_X1 U8600 ( .A1(n6693), .A2(n7543), .ZN(n7538) );
  OR2_X1 U8601 ( .A1(n13990), .A2(n13354), .ZN(n13355) );
  INV_X1 U8602 ( .A(n13990), .ZN(n13799) );
  OAI22_X1 U8603 ( .A1(n13840), .A2(n13841), .B1(n13850), .B2(n13367), .ZN(
        n13836) );
  AND2_X1 U8604 ( .A1(n13847), .A2(n13827), .ZN(n13829) );
  AND2_X1 U8605 ( .A1(n13861), .A2(n13850), .ZN(n13847) );
  NAND2_X1 U8606 ( .A1(n7575), .A2(n7578), .ZN(n7574) );
  INV_X1 U8607 ( .A(n7576), .ZN(n7575) );
  INV_X1 U8608 ( .A(n7563), .ZN(n7561) );
  AOI21_X1 U8609 ( .B1(n7564), .B2(n13202), .A(n7566), .ZN(n7563) );
  INV_X1 U8610 ( .A(n7545), .ZN(n7544) );
  AOI21_X1 U8611 ( .B1(n13940), .B2(n7548), .A(n7553), .ZN(n7545) );
  NOR2_X1 U8612 ( .A1(n11755), .A2(n14037), .ZN(n13932) );
  NAND2_X1 U8613 ( .A1(n11414), .A2(n6697), .ZN(n11598) );
  AND2_X1 U8614 ( .A1(n11414), .A2(n7080), .ZN(n14809) );
  AND2_X1 U8615 ( .A1(n7517), .A2(n7516), .ZN(n14808) );
  NAND2_X1 U8616 ( .A1(n13052), .A2(n14786), .ZN(n7516) );
  NAND2_X1 U8617 ( .A1(n14808), .A2(n14807), .ZN(n14806) );
  AND2_X1 U8618 ( .A1(n11414), .A2(n14824), .ZN(n14811) );
  INV_X1 U8619 ( .A(n13196), .ZN(n11410) );
  NOR2_X1 U8620 ( .A1(n15142), .A2(n11178), .ZN(n11179) );
  OR2_X1 U8621 ( .A1(n15061), .A2(n11181), .ZN(n15064) );
  NAND2_X1 U8622 ( .A1(n7076), .A2(n7075), .ZN(n10897) );
  NOR2_X1 U8623 ( .A1(n10527), .A2(n13022), .ZN(n7075) );
  OR2_X1 U8624 ( .A1(n13022), .A2(n10922), .ZN(n7528) );
  INV_X1 U8625 ( .A(n13270), .ZN(n10922) );
  INV_X1 U8626 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10579) );
  OR2_X1 U8627 ( .A1(n10580), .A2(n10579), .ZN(n10766) );
  OR2_X1 U8628 ( .A1(n10410), .A2(n10409), .ZN(n10580) );
  INV_X1 U8629 ( .A(n7529), .ZN(n10875) );
  NOR2_X1 U8630 ( .A1(n7077), .A2(n10527), .ZN(n10852) );
  INV_X1 U8631 ( .A(n10512), .ZN(n10511) );
  NAND2_X1 U8632 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n10133) );
  INV_X1 U8633 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10132) );
  CLKBUF_X1 U8634 ( .A(n10516), .Z(n13962) );
  INV_X1 U8635 ( .A(n13185), .ZN(n10473) );
  INV_X1 U8636 ( .A(n14784), .ZN(n13949) );
  OR2_X1 U8637 ( .A1(n9793), .A2(n13226), .ZN(n10164) );
  NOR2_X1 U8638 ( .A1(n10172), .A2(n12976), .ZN(n10173) );
  AND2_X1 U8639 ( .A1(n7572), .A2(n7571), .ZN(n13842) );
  INV_X1 U8640 ( .A(n13064), .ZN(n14048) );
  INV_X1 U8641 ( .A(n7517), .ZN(n14823) );
  INV_X1 U8642 ( .A(n15150), .ZN(n15114) );
  AND2_X1 U8643 ( .A1(n9412), .A2(n6987), .ZN(n6986) );
  NOR2_X1 U8644 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n6987) );
  OR2_X1 U8645 ( .A1(n9594), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n9596) );
  OR2_X1 U8646 ( .A1(n9504), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n9506) );
  INV_X1 U8647 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n9471) );
  INV_X1 U8648 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9795) );
  OAI211_X1 U8649 ( .C1(n6884), .C2(n7414), .A(n6816), .B(n6883), .ZN(n6882)
         );
  NAND2_X1 U8650 ( .A1(n10735), .A2(n6880), .ZN(n6884) );
  NAND2_X1 U8651 ( .A1(n12011), .A2(n12010), .ZN(n12012) );
  INV_X1 U8652 ( .A(n12008), .ZN(n12011) );
  OR2_X1 U8653 ( .A1(n8587), .A2(n11211), .ZN(n8609) );
  NAND2_X1 U8654 ( .A1(n14199), .A2(n14200), .ZN(n7441) );
  OR2_X1 U8655 ( .A1(n8665), .A2(n8298), .ZN(n8677) );
  AOI21_X1 U8656 ( .B1(n6906), .B2(n6904), .A(n6765), .ZN(n6903) );
  INV_X1 U8657 ( .A(n14175), .ZN(n6904) );
  INV_X1 U8658 ( .A(n6906), .ZN(n6905) );
  NAND2_X1 U8659 ( .A1(n12023), .A2(n12022), .ZN(n12024) );
  AOI21_X1 U8660 ( .B1(n12024), .B2(n7410), .A(n14148), .ZN(n7409) );
  INV_X1 U8661 ( .A(n14220), .ZN(n7410) );
  AND2_X1 U8662 ( .A1(n12089), .A2(n12088), .ZN(n14163) );
  OR2_X1 U8663 ( .A1(n12084), .A2(n14104), .ZN(n12089) );
  OR2_X1 U8664 ( .A1(n14103), .A2(n12084), .ZN(n14162) );
  OAI21_X1 U8665 ( .B1(n6607), .B2(n10738), .A(n7434), .ZN(n10085) );
  AOI21_X1 U8666 ( .B1(n12112), .B2(n11130), .A(n7435), .ZN(n7434) );
  NOR2_X1 U8667 ( .A1(n10367), .A2(n8410), .ZN(n7435) );
  NAND2_X1 U8668 ( .A1(n10089), .A2(n10251), .ZN(n10250) );
  OR2_X1 U8669 ( .A1(n12078), .A2(n14185), .ZN(n14187) );
  OR2_X1 U8670 ( .A1(n14102), .A2(n14131), .ZN(n14186) );
  NAND2_X1 U8671 ( .A1(n11899), .A2(n6855), .ZN(n6854) );
  INV_X1 U8672 ( .A(n11901), .ZN(n6855) );
  OR2_X1 U8673 ( .A1(n7418), .A2(n6705), .ZN(n7416) );
  AND2_X1 U8674 ( .A1(n7420), .A2(n10929), .ZN(n7418) );
  AND2_X1 U8675 ( .A1(n7420), .A2(n7417), .ZN(n7415) );
  NAND2_X1 U8676 ( .A1(n10735), .A2(n6885), .ZN(n10740) );
  AOI21_X1 U8677 ( .B1(n6903), .B2(n6905), .A(n6901), .ZN(n6900) );
  INV_X1 U8678 ( .A(n14140), .ZN(n6901) );
  NAND2_X1 U8679 ( .A1(n14219), .A2(n14220), .ZN(n14218) );
  AND4_X1 U8680 ( .A1(n8808), .A2(n8807), .A3(n8806), .A4(n8805), .ZN(n12129)
         );
  INV_X1 U8681 ( .A(n9063), .ZN(n8804) );
  NAND2_X1 U8682 ( .A1(n8445), .A2(n6911), .ZN(n6910) );
  NAND2_X1 U8683 ( .A1(n9063), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6911) );
  NAND2_X1 U8684 ( .A1(n9063), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n8425) );
  NAND2_X1 U8685 ( .A1(n6682), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n8399) );
  AND2_X1 U8686 ( .A1(n9454), .A2(n6772), .ZN(n9455) );
  NOR2_X1 U8687 ( .A1(n9455), .A2(n7098), .ZN(n14262) );
  AND2_X1 U8688 ( .A1(n9458), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7098) );
  INV_X1 U8689 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n14274) );
  NAND2_X1 U8690 ( .A1(n9873), .A2(n7087), .ZN(n9834) );
  OR2_X1 U8691 ( .A1(n9842), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n7087) );
  NOR2_X1 U8692 ( .A1(n10552), .A2(n7091), .ZN(n10556) );
  AND2_X1 U8693 ( .A1(n10553), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7091) );
  NAND2_X1 U8694 ( .A1(n10556), .A2(n10555), .ZN(n10711) );
  NAND2_X1 U8695 ( .A1(n10711), .A2(n7090), .ZN(n10713) );
  NAND2_X1 U8696 ( .A1(n10708), .A2(n10554), .ZN(n7090) );
  NAND2_X1 U8697 ( .A1(n10713), .A2(n10714), .ZN(n11026) );
  NOR2_X1 U8698 ( .A1(n11207), .A2(n7093), .ZN(n11209) );
  AND2_X1 U8699 ( .A1(n11208), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7093) );
  NAND2_X1 U8700 ( .A1(n11209), .A2(n11210), .ZN(n11643) );
  XNOR2_X1 U8701 ( .A(n11645), .B(n11646), .ZN(n14912) );
  AND2_X1 U8702 ( .A1(n14313), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n14320) );
  NAND2_X1 U8703 ( .A1(n12132), .A2(n11965), .ZN(n11966) );
  NAND2_X1 U8704 ( .A1(n9045), .A2(n9044), .ZN(n14561) );
  AND2_X1 U8705 ( .A1(n11978), .A2(n8784), .ZN(n12126) );
  AND2_X1 U8706 ( .A1(n8783), .A2(n8766), .ZN(n14084) );
  NOR2_X1 U8707 ( .A1(n14358), .A2(n7302), .ZN(n7301) );
  INV_X1 U8708 ( .A(n8844), .ZN(n7302) );
  NAND2_X1 U8709 ( .A1(n14380), .A2(n8844), .ZN(n14356) );
  AND2_X1 U8710 ( .A1(n8765), .A2(n8754), .ZN(n14377) );
  NAND2_X1 U8711 ( .A1(n8299), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8300) );
  AND2_X1 U8712 ( .A1(n8718), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8739) );
  NOR2_X1 U8713 ( .A1(n14435), .A2(n7101), .ZN(n14412) );
  INV_X1 U8714 ( .A(n7103), .ZN(n7101) );
  OR2_X1 U8715 ( .A1(n14456), .A2(n14599), .ZN(n14435) );
  OR2_X1 U8716 ( .A1(n14434), .A2(n14448), .ZN(n14432) );
  NOR2_X1 U8717 ( .A1(n14501), .A2(n14609), .ZN(n14481) );
  NAND2_X1 U8718 ( .A1(n14524), .A2(n14507), .ZN(n14501) );
  NAND2_X1 U8719 ( .A1(n7285), .A2(n7283), .ZN(n14490) );
  NAND2_X1 U8720 ( .A1(n7285), .A2(n8982), .ZN(n14513) );
  NAND2_X1 U8721 ( .A1(n8833), .A2(n8832), .ZN(n14535) );
  NAND2_X1 U8722 ( .A1(n11883), .A2(n8853), .ZN(n14534) );
  NOR2_X1 U8723 ( .A1(n8609), .A2(n8608), .ZN(n8626) );
  AND2_X1 U8724 ( .A1(n8626), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8637) );
  NAND2_X1 U8725 ( .A1(n11825), .A2(n14231), .ZN(n11882) );
  NOR2_X1 U8726 ( .A1(n11608), .A2(n14639), .ZN(n11825) );
  NAND2_X1 U8727 ( .A1(n14711), .A2(n14860), .ZN(n11608) );
  NOR2_X1 U8728 ( .A1(n8560), .A2(n8559), .ZN(n8577) );
  OR2_X1 U8729 ( .A1(n8547), .A2(n14845), .ZN(n8560) );
  AOI21_X1 U8730 ( .B1(n7501), .B2(n11109), .A(n6754), .ZN(n7499) );
  INV_X1 U8731 ( .A(n7501), .ZN(n7500) );
  NAND2_X1 U8732 ( .A1(n11192), .A2(n8820), .ZN(n11386) );
  NAND2_X1 U8733 ( .A1(n11107), .A2(n8819), .ZN(n11194) );
  NAND2_X1 U8734 ( .A1(n11194), .A2(n11193), .ZN(n11192) );
  NOR2_X1 U8735 ( .A1(n8513), .A2(n8512), .ZN(n8528) );
  NAND3_X1 U8736 ( .A1(n6698), .A2(n10806), .A3(n14897), .ZN(n11195) );
  INV_X1 U8737 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n8496) );
  OR2_X1 U8738 ( .A1(n8497), .A2(n8496), .ZN(n8513) );
  NAND2_X1 U8739 ( .A1(n10806), .A2(n7106), .ZN(n11007) );
  INV_X1 U8740 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n9866) );
  OR2_X1 U8741 ( .A1(n8484), .A2(n9866), .ZN(n8497) );
  NAND2_X1 U8742 ( .A1(n10806), .A2(n11041), .ZN(n11006) );
  AND2_X1 U8743 ( .A1(n10808), .A2(n14948), .ZN(n10806) );
  NAND2_X1 U8744 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n8458) );
  INV_X1 U8745 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n8457) );
  NOR2_X1 U8746 ( .A1(n8458), .A2(n8457), .ZN(n8470) );
  NAND2_X1 U8747 ( .A1(n7507), .A2(n7508), .ZN(n10812) );
  NOR2_X1 U8748 ( .A1(n10746), .A2(n10628), .ZN(n10808) );
  NAND2_X1 U8749 ( .A1(n9099), .A2(n8898), .ZN(n7288) );
  NAND2_X1 U8750 ( .A1(n8422), .A2(n9099), .ZN(n10235) );
  INV_X1 U8751 ( .A(n9099), .ZN(n10232) );
  NAND2_X1 U8752 ( .A1(n10232), .A2(n10231), .ZN(n10230) );
  NAND2_X1 U8753 ( .A1(n11129), .A2(n10594), .ZN(n10825) );
  AND2_X1 U8754 ( .A1(n8850), .A2(n11277), .ZN(n9822) );
  AND2_X1 U8755 ( .A1(n11823), .A2(n11822), .ZN(n14636) );
  XNOR2_X1 U8756 ( .A(n9078), .B(n9077), .ZN(n14068) );
  INV_X1 U8757 ( .A(n7110), .ZN(n9078) );
  XNOR2_X1 U8758 ( .A(n9052), .B(n9051), .ZN(n13157) );
  NAND2_X1 U8759 ( .A1(n7123), .A2(n9041), .ZN(n9052) );
  NAND2_X1 U8760 ( .A1(n7118), .A2(n7124), .ZN(n7123) );
  AND2_X1 U8761 ( .A1(n8871), .A2(n8870), .ZN(n8874) );
  INV_X1 U8762 ( .A(n8388), .ZN(n8870) );
  CLKBUF_X1 U8763 ( .A(n8387), .Z(n8388) );
  XNOR2_X1 U8764 ( .A(n8760), .B(n8748), .ZN(n12829) );
  CLKBUF_X1 U8765 ( .A(n8866), .Z(n8868) );
  XNOR2_X1 U8766 ( .A(n8733), .B(n8729), .ZN(n12796) );
  INV_X1 U8767 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8877) );
  XNOR2_X1 U8768 ( .A(n8715), .B(n8714), .ZN(n12783) );
  NAND2_X1 U8769 ( .A1(n8712), .A2(n8711), .ZN(n8715) );
  XNOR2_X1 U8770 ( .A(n8798), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9089) );
  INV_X1 U8771 ( .A(n8797), .ZN(n7242) );
  XNOR2_X1 U8772 ( .A(n8691), .B(n8690), .ZN(n12760) );
  NAND2_X1 U8773 ( .A1(n8688), .A2(n8687), .ZN(n8691) );
  INV_X1 U8774 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8791) );
  XNOR2_X1 U8775 ( .A(n8602), .B(n8601), .ZN(n11542) );
  AND2_X1 U8776 ( .A1(n8509), .A2(n8524), .ZN(n10290) );
  XNOR2_X1 U8777 ( .A(n8478), .B(n8477), .ZN(n10574) );
  OAI21_X1 U8778 ( .B1(n8418), .B2(n8417), .A(n8313), .ZN(n8431) );
  INV_X1 U8779 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9331) );
  XNOR2_X1 U8780 ( .A(n9329), .B(n9330), .ZN(n6934) );
  XNOR2_X1 U8781 ( .A(n9289), .B(n15234), .ZN(n9326) );
  XNOR2_X1 U8782 ( .A(n9325), .B(n7274), .ZN(n9333) );
  INV_X1 U8783 ( .A(n9324), .ZN(n7274) );
  NAND2_X1 U8784 ( .A1(n15439), .A2(n9338), .ZN(n9339) );
  OAI22_X1 U8785 ( .A1(n9342), .A2(n9294), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n9340), .ZN(n9345) );
  AND2_X1 U8786 ( .A1(n14691), .A2(n7264), .ZN(n6919) );
  NOR2_X1 U8787 ( .A1(n9303), .A2(n9302), .ZN(n9354) );
  NOR2_X1 U8788 ( .A1(n10649), .A2(n9322), .ZN(n9302) );
  NOR2_X1 U8789 ( .A1(n9310), .A2(n9309), .ZN(n9370) );
  NAND2_X1 U8790 ( .A1(n7385), .A2(n12182), .ZN(n12139) );
  NAND2_X1 U8791 ( .A1(n8007), .A2(n8006), .ZN(n12492) );
  NAND2_X1 U8792 ( .A1(n9195), .A2(n9194), .ZN(n15184) );
  AOI21_X1 U8793 ( .B1(n9498), .B2(n8099), .A(n7811), .ZN(n15189) );
  AND3_X1 U8794 ( .A1(n7682), .A2(n7681), .A3(n7680), .ZN(n15200) );
  CLKBUF_X1 U8795 ( .A(n11046), .Z(n15181) );
  NAND2_X1 U8796 ( .A1(n10210), .A2(n7205), .ZN(n10211) );
  NAND2_X1 U8797 ( .A1(n7393), .A2(n7391), .ZN(n12154) );
  INV_X1 U8798 ( .A(n7395), .ZN(n7391) );
  AND4_X1 U8799 ( .A1(n7825), .A2(n7824), .A3(n7823), .A4(n7822), .ZN(n11526)
         );
  INV_X1 U8800 ( .A(n12465), .ZN(n12489) );
  NAND2_X1 U8801 ( .A1(n7946), .A2(n6991), .ZN(n6990) );
  NAND2_X1 U8802 ( .A1(n6993), .A2(SI_0_), .ZN(n6992) );
  AOI21_X1 U8803 ( .B1(n6850), .B2(n12145), .A(n7394), .ZN(n12191) );
  INV_X1 U8804 ( .A(n7396), .ZN(n7394) );
  NAND2_X1 U8805 ( .A1(n9201), .A2(n11574), .ZN(n6849) );
  AND4_X1 U8806 ( .A1(n7800), .A2(n7799), .A3(n7798), .A4(n7797), .ZN(n11442)
         );
  NAND2_X1 U8807 ( .A1(n7401), .A2(n9175), .ZN(n15208) );
  NAND2_X1 U8808 ( .A1(n12219), .A2(n12220), .ZN(n12218) );
  OR2_X1 U8809 ( .A1(n8059), .A2(n8047), .ZN(n12454) );
  NAND2_X1 U8810 ( .A1(n7372), .A2(n7376), .ZN(n11730) );
  NAND2_X1 U8811 ( .A1(n11509), .A2(n6725), .ZN(n7372) );
  NAND2_X1 U8812 ( .A1(n7022), .A2(n10423), .ZN(n7021) );
  NAND2_X1 U8813 ( .A1(n6833), .A2(n7181), .ZN(n7022) );
  INV_X1 U8814 ( .A(n10635), .ZN(n10427) );
  INV_X1 U8815 ( .A(n11709), .ZN(n12236) );
  INV_X1 U8816 ( .A(n11442), .ZN(n11342) );
  INV_X1 U8817 ( .A(n11094), .ZN(n12240) );
  INV_X1 U8818 ( .A(n10858), .ZN(n12241) );
  INV_X1 U8819 ( .A(n15354), .ZN(n12244) );
  OR2_X1 U8820 ( .A1(n9406), .A2(n12714), .ZN(n12245) );
  INV_X1 U8821 ( .A(n10035), .ZN(n6991) );
  INV_X1 U8822 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n13672) );
  NAND2_X1 U8823 ( .A1(n10157), .A2(n10054), .ZN(n10100) );
  INV_X1 U8824 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n15234) );
  NAND2_X1 U8825 ( .A1(n7256), .A2(n7255), .ZN(n15235) );
  NOR2_X1 U8826 ( .A1(n15276), .A2(n15275), .ZN(n15274) );
  AOI22_X1 U8827 ( .A1(n15283), .A2(n15282), .B1(n10673), .B2(n10672), .ZN(
        n15293) );
  NOR2_X1 U8828 ( .A1(n15311), .A2(n15312), .ZN(n15310) );
  NAND2_X1 U8829 ( .A1(n7246), .A2(n11065), .ZN(n7245) );
  NOR2_X1 U8830 ( .A1(n11223), .A2(n11222), .ZN(n11225) );
  AOI21_X1 U8831 ( .B1(n11054), .B2(n11053), .A(n7247), .ZN(n11223) );
  AOI21_X1 U8832 ( .B1(n12249), .B2(n12248), .A(n12247), .ZN(n12253) );
  INV_X1 U8833 ( .A(n6845), .ZN(n14743) );
  INV_X1 U8834 ( .A(n7254), .ZN(n14748) );
  OAI21_X1 U8835 ( .B1(n14763), .B2(n12311), .A(n12310), .ZN(n12333) );
  XNOR2_X1 U8836 ( .A(n6858), .B(n12346), .ZN(n12347) );
  NAND2_X1 U8837 ( .A1(n6860), .A2(n6859), .ZN(n6858) );
  OR2_X1 U8838 ( .A1(n8071), .A2(n8060), .ZN(n12438) );
  NAND2_X1 U8839 ( .A1(n12510), .A2(n12385), .ZN(n12498) );
  OAI21_X1 U8840 ( .B1(n12545), .B2(n7450), .A(n7448), .ZN(n12514) );
  NAND2_X1 U8841 ( .A1(n12545), .A2(n7454), .ZN(n7453) );
  NAND2_X1 U8842 ( .A1(n12374), .A2(n12373), .ZN(n12549) );
  NAND2_X1 U8843 ( .A1(n7931), .A2(n7930), .ZN(n12560) );
  NAND2_X1 U8844 ( .A1(n7917), .A2(n7916), .ZN(n12636) );
  NAND2_X1 U8845 ( .A1(n6847), .A2(n11568), .ZN(n11708) );
  NAND2_X1 U8846 ( .A1(n7005), .A2(n8192), .ZN(n11576) );
  NAND2_X1 U8847 ( .A1(n11527), .A2(n7202), .ZN(n7005) );
  NAND2_X1 U8848 ( .A1(n10721), .A2(n8163), .ZN(n11075) );
  AND3_X1 U8849 ( .A1(n7720), .A2(n7719), .A3(n7718), .ZN(n10802) );
  NAND2_X1 U8850 ( .A1(n10443), .A2(n10442), .ZN(n10723) );
  NAND2_X1 U8851 ( .A1(n7958), .A2(n7957), .ZN(n12626) );
  AOI21_X1 U8852 ( .B1(n12720), .B2(n8099), .A(n8093), .ZN(n12654) );
  NAND2_X1 U8853 ( .A1(n6824), .A2(n14775), .ZN(n6823) );
  NAND2_X1 U8854 ( .A1(n7971), .A2(n7970), .ZN(n12683) );
  NAND2_X1 U8855 ( .A1(n7869), .A2(n7868), .ZN(n12711) );
  NAND2_X1 U8856 ( .A1(n7853), .A2(n7852), .ZN(n11798) );
  AND3_X1 U8857 ( .A1(n7699), .A2(n7698), .A3(n7697), .ZN(n11274) );
  AOI21_X1 U8858 ( .B1(n11267), .B2(n11266), .A(n11265), .ZN(n15421) );
  INV_X1 U8859 ( .A(n10453), .ZN(n12715) );
  OR2_X1 U8860 ( .A1(n8081), .A2(n8080), .ZN(n8082) );
  NAND2_X1 U8861 ( .A1(n8275), .A2(n8274), .ZN(n9148) );
  OR2_X1 U8862 ( .A1(n8273), .A2(P3_IR_REG_25__SCAN_IN), .ZN(n8274) );
  MUX2_X1 U8863 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8272), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8275) );
  NAND2_X1 U8864 ( .A1(n7187), .A2(n7185), .ZN(n7999) );
  NAND2_X1 U8865 ( .A1(n7187), .A2(n7981), .ZN(n7985) );
  NOR2_X1 U8866 ( .A1(n8123), .A2(n8122), .ZN(n8124) );
  NAND2_X1 U8867 ( .A1(n8128), .A2(n8119), .ZN(n8125) );
  NOR2_X1 U8868 ( .A1(P3_IR_REG_21__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n8122) );
  NAND2_X1 U8869 ( .A1(n7157), .A2(n7942), .ZN(n7956) );
  NAND2_X1 U8870 ( .A1(n7941), .A2(n7940), .ZN(n7157) );
  NAND2_X1 U8871 ( .A1(n7879), .A2(n7878), .ZN(n7163) );
  INV_X1 U8872 ( .A(SI_12_), .ZN(n9553) );
  NAND2_X1 U8873 ( .A1(n7766), .A2(n7765), .ZN(n7769) );
  INV_X1 U8874 ( .A(n10650), .ZN(n15296) );
  NAND2_X1 U8875 ( .A1(n7745), .A2(n7744), .ZN(n7748) );
  INV_X1 U8876 ( .A(n10667), .ZN(n10651) );
  NAND2_X1 U8877 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n7654) );
  NAND2_X1 U8878 ( .A1(n7312), .A2(n7317), .ZN(n10758) );
  NAND2_X1 U8879 ( .A1(n10402), .A2(n7315), .ZN(n7312) );
  OAI21_X1 U8880 ( .B1(n11839), .B2(n7325), .A(n7322), .ZN(n12881) );
  NAND2_X1 U8881 ( .A1(n12735), .A2(n12734), .ZN(n14027) );
  OR2_X1 U8882 ( .A1(n12889), .A2(n7337), .ZN(n7336) );
  INV_X1 U8883 ( .A(n7335), .ZN(n7334) );
  OAI22_X1 U8884 ( .A1(n12889), .A2(n6745), .B1(n12887), .B2(n12888), .ZN(
        n7335) );
  NOR2_X1 U8885 ( .A1(n11301), .A2(n11300), .ZN(n11308) );
  NAND2_X1 U8886 ( .A1(n11304), .A2(n11303), .ZN(n14830) );
  NAND2_X1 U8887 ( .A1(n12813), .A2(n12812), .ZN(n13995) );
  AND3_X1 U8888 ( .A1(n11554), .A2(n11553), .A3(n11552), .ZN(n14785) );
  OAI21_X1 U8889 ( .B1(n11301), .B2(n7332), .A(n7331), .ZN(n11624) );
  NAND2_X1 U8890 ( .A1(n11154), .A2(n11153), .ZN(n13040) );
  NAND2_X1 U8891 ( .A1(n11866), .A2(n11865), .ZN(n12731) );
  NAND2_X1 U8892 ( .A1(n10402), .A2(n10401), .ZN(n10573) );
  NAND2_X1 U8893 ( .A1(n10403), .A2(n10117), .ZN(n10405) );
  NAND2_X1 U8894 ( .A1(n12828), .A2(n12827), .ZN(n12959) );
  AND4_X1 U8895 ( .A1(n11370), .A2(n11369), .A3(n11368), .A4(n11367), .ZN(
        n13066) );
  OAI211_X1 U8896 ( .C1(n7129), .C2(n13247), .A(n13248), .B(n13249), .ZN(n7125) );
  NOR2_X1 U8897 ( .A1(n13245), .A2(n7130), .ZN(n7129) );
  NAND4_X1 U8898 ( .A1(n10278), .A2(n10277), .A3(n10276), .A4(n10275), .ZN(
        n13272) );
  NAND4_X1 U8899 ( .A1(n9940), .A2(n9939), .A3(n9938), .A4(n9937), .ZN(n13948)
         );
  OR2_X1 U8900 ( .A1(n10135), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n9939) );
  OR2_X1 U8901 ( .A1(n10135), .A2(n10478), .ZN(n9926) );
  OR2_X1 U8902 ( .A1(n12775), .A2(n10186), .ZN(n9761) );
  OR2_X1 U8903 ( .A1(n10135), .A2(n9994), .ZN(n9762) );
  INV_X1 U8904 ( .A(n13345), .ZN(n13344) );
  NAND2_X1 U8905 ( .A1(n6972), .A2(n6973), .ZN(n13789) );
  NAND2_X1 U8906 ( .A1(n6977), .A2(n6978), .ZN(n13807) );
  NAND2_X1 U8907 ( .A1(n13369), .A2(n6979), .ZN(n6977) );
  NAND2_X1 U8908 ( .A1(n13369), .A2(n7582), .ZN(n13824) );
  NAND2_X1 U8909 ( .A1(n13874), .A2(n7583), .ZN(n13855) );
  NAND2_X1 U8910 ( .A1(n13892), .A2(n7584), .ZN(n13877) );
  AND2_X1 U8911 ( .A1(n13350), .A2(n7564), .ZN(n13938) );
  NAND2_X1 U8912 ( .A1(n13350), .A2(n7587), .ZN(n13939) );
  NAND2_X1 U8913 ( .A1(n7547), .A2(n7549), .ZN(n13924) );
  NAND2_X1 U8914 ( .A1(n7546), .A2(n6719), .ZN(n7547) );
  AND2_X1 U8915 ( .A1(n7551), .A2(n7554), .ZN(n13362) );
  NAND2_X1 U8916 ( .A1(n7546), .A2(n11737), .ZN(n7551) );
  INV_X1 U8917 ( .A(n13941), .ZN(n15069) );
  AND2_X1 U8918 ( .A1(n7513), .A2(n12970), .ZN(n15086) );
  INV_X1 U8919 ( .A(n10173), .ZN(n7513) );
  INV_X1 U8920 ( .A(n13975), .ZN(n13976) );
  AND2_X1 U8921 ( .A1(n9788), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15082) );
  NAND2_X1 U8922 ( .A1(n9538), .A2(n9539), .ZN(n14069) );
  BUF_X1 U8923 ( .A(n9542), .Z(n11939) );
  NAND2_X1 U8924 ( .A1(n6837), .A2(n10190), .ZN(n10342) );
  INV_X1 U8925 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n13518) );
  AND2_X1 U8926 ( .A1(n9753), .A2(n10283), .ZN(n11359) );
  INV_X1 U8927 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9731) );
  INV_X1 U8928 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10877) );
  INV_X1 U8929 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9556) );
  INV_X1 U8930 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9534) );
  INV_X1 U8931 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9515) );
  INV_X1 U8932 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9509) );
  INV_X1 U8933 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9497) );
  INV_X1 U8934 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9476) );
  INV_X1 U8935 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9918) );
  NAND2_X1 U8936 ( .A1(n12013), .A2(n12012), .ZN(n14092) );
  NAND2_X1 U8937 ( .A1(n7441), .A2(n12045), .ZN(n14116) );
  AND2_X1 U8938 ( .A1(n7431), .A2(n7428), .ZN(n7422) );
  OAI21_X1 U8939 ( .B1(n6737), .B2(n7431), .A(n7424), .ZN(n7423) );
  INV_X1 U8940 ( .A(n7428), .ZN(n7425) );
  NAND2_X1 U8941 ( .A1(n12125), .A2(n7427), .ZN(n7426) );
  NAND2_X1 U8942 ( .A1(n8541), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8396) );
  INV_X1 U8943 ( .A(n11915), .ZN(n11916) );
  NAND2_X1 U8944 ( .A1(n14852), .A2(n11910), .ZN(n11914) );
  AND2_X1 U8945 ( .A1(n6812), .A2(n7419), .ZN(n10949) );
  NAND2_X1 U8946 ( .A1(n10928), .A2(n10929), .ZN(n7419) );
  INV_X1 U8947 ( .A(n11130), .ZN(n10098) );
  INV_X1 U8948 ( .A(n7439), .ZN(n7438) );
  AOI21_X1 U8949 ( .B1(n7439), .B2(n7437), .A(n6795), .ZN(n7436) );
  INV_X1 U8950 ( .A(n14445), .ZN(n14599) );
  NAND2_X1 U8951 ( .A1(n8437), .A2(n14270), .ZN(n7299) );
  NAND2_X1 U8952 ( .A1(n8541), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7300) );
  NAND2_X1 U8953 ( .A1(n8647), .A2(n8646), .ZN(n14620) );
  NAND2_X1 U8954 ( .A1(n8455), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n8401) );
  INV_X1 U8955 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9284) );
  INV_X1 U8956 ( .A(n7089), .ZN(n14277) );
  NAND2_X1 U8957 ( .A1(n14281), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7088) );
  NOR2_X1 U8958 ( .A1(n9857), .A2(n9856), .ZN(n9888) );
  NOR2_X1 U8959 ( .A1(n9854), .A2(n7095), .ZN(n9857) );
  NOR2_X1 U8960 ( .A1(n7097), .A2(n7096), .ZN(n7095) );
  NOR2_X1 U8961 ( .A1(n9888), .A2(n7094), .ZN(n9891) );
  AND2_X1 U8962 ( .A1(n9892), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7094) );
  NAND2_X1 U8963 ( .A1(n9891), .A2(n9890), .ZN(n9954) );
  NOR2_X1 U8964 ( .A1(n14321), .A2(n7086), .ZN(n14313) );
  AND2_X1 U8965 ( .A1(n14311), .A2(n14323), .ZN(n7086) );
  XNOR2_X1 U8966 ( .A(n7085), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n14333) );
  NOR2_X1 U8967 ( .A1(n14320), .A2(n14321), .ZN(n7085) );
  INV_X1 U8968 ( .A(n12132), .ZN(n11998) );
  AND2_X1 U8969 ( .A1(n14386), .A2(n8744), .ZN(n14373) );
  NOR2_X1 U8970 ( .A1(n14397), .A2(n6954), .ZN(n6953) );
  INV_X1 U8971 ( .A(n8842), .ZN(n6954) );
  NAND2_X1 U8972 ( .A1(n7276), .A2(n8842), .ZN(n14398) );
  OAI21_X1 U8973 ( .B1(n6840), .B2(n6694), .A(n8838), .ZN(n14449) );
  NAND2_X1 U8974 ( .A1(n7483), .A2(n8673), .ZN(n14476) );
  NAND2_X1 U8975 ( .A1(n8636), .A2(n8635), .ZN(n14550) );
  NAND2_X1 U8976 ( .A1(n8625), .A2(n8624), .ZN(n14153) );
  NAND2_X1 U8977 ( .A1(n8827), .A2(n8826), .ZN(n11612) );
  OAI21_X1 U8978 ( .B1(n14698), .B2(n14709), .A(n8566), .ZN(n11457) );
  NAND2_X1 U8979 ( .A1(n8558), .A2(n8557), .ZN(n14707) );
  NAND2_X1 U8980 ( .A1(n11112), .A2(n7501), .ZN(n11190) );
  INV_X1 U8981 ( .A(n14506), .ZN(n14706) );
  INV_X1 U8982 ( .A(n14529), .ZN(n14716) );
  OR2_X1 U8983 ( .A1(n10081), .A2(n10369), .ZN(n14498) );
  OR2_X1 U8984 ( .A1(n14526), .A2(n14552), .ZN(n14529) );
  OR2_X1 U8985 ( .A1(n14526), .A2(n14546), .ZN(n14506) );
  NOR2_X1 U8986 ( .A1(n14559), .A2(n6827), .ZN(n6826) );
  OAI21_X1 U8987 ( .B1(n11999), .B2(n14959), .A(n6841), .ZN(n14565) );
  AND2_X1 U8988 ( .A1(n12004), .A2(n8857), .ZN(n6841) );
  NAND2_X1 U8989 ( .A1(n14570), .A2(n7599), .ZN(n14646) );
  AND2_X1 U8990 ( .A1(n14569), .A2(n7591), .ZN(n7599) );
  INV_X1 U8991 ( .A(n14566), .ZN(n14570) );
  AND2_X1 U8992 ( .A1(n6776), .A2(n8288), .ZN(n7510) );
  INV_X1 U8993 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7511) );
  NAND2_X1 U8994 ( .A1(n7111), .A2(n7115), .ZN(n9075) );
  NAND2_X1 U8995 ( .A1(n8389), .A2(n6825), .ZN(n8386) );
  NOR2_X1 U8996 ( .A1(n8289), .A2(n8290), .ZN(n6825) );
  XNOR2_X1 U8997 ( .A(n9043), .B(n9042), .ZN(n12891) );
  OR2_X1 U8998 ( .A1(n8387), .A2(n7290), .ZN(n7289) );
  NAND2_X1 U8999 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n7290) );
  XNOR2_X1 U9000 ( .A(n8772), .B(n8761), .ZN(n12856) );
  NAND2_X1 U9001 ( .A1(n7141), .A2(n7142), .ZN(n8772) );
  INV_X1 U9002 ( .A(n8874), .ZN(n11726) );
  INV_X1 U9003 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n8860) );
  OAI21_X1 U9004 ( .B1(n8876), .B2(P1_IR_REG_23__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8861) );
  XNOR2_X1 U9005 ( .A(n8701), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14673) );
  OR2_X1 U9006 ( .A1(n8859), .A2(n8290), .ZN(n8799) );
  INV_X1 U9007 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9727) );
  INV_X1 U9008 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9733) );
  INV_X1 U9009 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9558) );
  INV_X1 U9010 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9530) );
  INV_X1 U9011 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9517) );
  OR2_X1 U9012 ( .A1(n8452), .A2(n8451), .ZN(n9884) );
  INV_X1 U9013 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9502) );
  INV_X1 U9014 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9488) );
  NAND2_X1 U9015 ( .A1(n8419), .A2(n7474), .ZN(n8428) );
  INV_X1 U9016 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9490) );
  XNOR2_X1 U9017 ( .A(n6934), .B(P2_ADDR_REG_1__SCAN_IN), .ZN(n15452) );
  NAND2_X1 U9018 ( .A1(n6914), .A2(n14681), .ZN(n15448) );
  XNOR2_X1 U9019 ( .A(n7271), .B(n9337), .ZN(n15441) );
  XNOR2_X1 U9020 ( .A(n9339), .B(n7270), .ZN(n14687) );
  AND2_X1 U9021 ( .A1(n7261), .A2(n7260), .ZN(n14873) );
  INV_X1 U9022 ( .A(n14694), .ZN(n7261) );
  OAI21_X1 U9023 ( .B1(n7263), .B2(n7262), .A(P2_ADDR_REG_10__SCAN_IN), .ZN(
        n7260) );
  NAND2_X1 U9024 ( .A1(n7269), .A2(n9365), .ZN(n7268) );
  NAND2_X1 U9025 ( .A1(n14880), .A2(n14879), .ZN(n14878) );
  AOI21_X1 U9026 ( .B1(n6932), .B2(n6931), .A(n9372), .ZN(n6926) );
  NAND2_X1 U9027 ( .A1(n6931), .A2(n6928), .ZN(n6927) );
  NAND2_X1 U9028 ( .A1(n6925), .A2(n6931), .ZN(n6924) );
  INV_X1 U9029 ( .A(n9374), .ZN(n7272) );
  NAND2_X1 U9030 ( .A1(n15194), .A2(n9170), .ZN(n10486) );
  OAI21_X1 U9031 ( .B1(n12655), .B2(n15433), .A(n6831), .ZN(P3_U3488) );
  AOI21_X1 U9032 ( .B1(n12410), .B2(n6853), .A(n6832), .ZN(n6831) );
  NOR2_X1 U9033 ( .A1(n15436), .A2(n12587), .ZN(n6832) );
  OAI21_X1 U9034 ( .B1(n12658), .B2(n15433), .A(n6851), .ZN(P3_U3487) );
  AOI21_X1 U9035 ( .B1(n12426), .B2(n6853), .A(n6852), .ZN(n6851) );
  NOR2_X1 U9036 ( .A1(n15436), .A2(n12590), .ZN(n6852) );
  OR2_X1 U9037 ( .A1(n12707), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n7007) );
  AOI211_X1 U9038 ( .C1(n15068), .C2(n13984), .A(n13416), .B(n13415), .ZN(
        n13417) );
  NAND2_X1 U9039 ( .A1(n6896), .A2(n14904), .ZN(n6895) );
  INV_X1 U9040 ( .A(n6922), .ZN(n14692) );
  NAND2_X1 U9041 ( .A1(n14887), .A2(n14886), .ZN(n14885) );
  OAI21_X1 U9042 ( .B1(n9381), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n14675), .ZN(
        n6819) );
  AND2_X1 U9043 ( .A1(n7464), .A2(n7462), .ZN(n6691) );
  AND3_X1 U9044 ( .A1(n7083), .A2(n13394), .A3(n7082), .ZN(n6692) );
  INV_X1 U9045 ( .A(n11568), .ZN(n7202) );
  OR2_X1 U9046 ( .A1(n13799), .A2(n13373), .ZN(n6693) );
  INV_X1 U9047 ( .A(n14448), .ZN(n7277) );
  NAND2_X1 U9048 ( .A1(n6722), .A2(n7189), .ZN(n7777) );
  OR2_X1 U9049 ( .A1(n14462), .A2(n6969), .ZN(n6694) );
  AOI21_X1 U9050 ( .B1(n7481), .B2(n14495), .A(n6753), .ZN(n7480) );
  INV_X1 U9051 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8289) );
  NOR2_X1 U9052 ( .A1(n8836), .A2(n14495), .ZN(n6696) );
  NAND2_X1 U9053 ( .A1(n11869), .A2(n11868), .ZN(n14030) );
  INV_X1 U9054 ( .A(n12594), .ZN(n6824) );
  AND2_X1 U9055 ( .A1(n7080), .A2(n13064), .ZN(n6697) );
  INV_X1 U9056 ( .A(n12111), .ZN(n7430) );
  INV_X1 U9057 ( .A(n9367), .ZN(n9365) );
  AOI21_X1 U9058 ( .B1(n7040), .B2(n7038), .A(n6750), .ZN(n7037) );
  INV_X1 U9059 ( .A(n7037), .ZN(n7033) );
  AND2_X1 U9060 ( .A1(n7106), .A2(n7105), .ZN(n6698) );
  NAND2_X1 U9061 ( .A1(n11361), .A2(n11360), .ZN(n13052) );
  AND4_X1 U9062 ( .A1(n7605), .A2(n7604), .A3(n7750), .A4(n7696), .ZN(n6699)
         );
  AND2_X1 U9063 ( .A1(n7406), .A2(n7405), .ZN(n8797) );
  NAND2_X1 U9064 ( .A1(n12785), .A2(n12784), .ZN(n14004) );
  INV_X1 U9065 ( .A(n14004), .ZN(n13850) );
  INV_X1 U9066 ( .A(n11673), .ZN(n6890) );
  AND2_X1 U9067 ( .A1(n6892), .A2(n11673), .ZN(n6700) );
  INV_X1 U9068 ( .A(n12503), .ZN(n7054) );
  NOR2_X1 U9069 ( .A1(n6727), .A2(n11010), .ZN(n6701) );
  AND2_X1 U9070 ( .A1(n11728), .A2(n11727), .ZN(n6702) );
  AND2_X1 U9071 ( .A1(n6768), .A2(n6897), .ZN(n6703) );
  INV_X1 U9072 ( .A(n11662), .ZN(n7412) );
  AND2_X1 U9073 ( .A1(n7522), .A2(n6747), .ZN(n6704) );
  AND2_X1 U9074 ( .A1(n7420), .A2(n6729), .ZN(n6705) );
  INV_X1 U9075 ( .A(n8925), .ZN(n7232) );
  OR2_X1 U9076 ( .A1(n11957), .A2(n11673), .ZN(n6706) );
  OR2_X1 U9077 ( .A1(n9289), .A2(n15234), .ZN(n6707) );
  NAND2_X1 U9078 ( .A1(n13159), .A2(n13158), .ZN(n13380) );
  INV_X1 U9079 ( .A(n13380), .ZN(n7083) );
  NAND2_X1 U9080 ( .A1(n6837), .A2(n7342), .ZN(n9613) );
  NAND2_X1 U9081 ( .A1(n8121), .A2(n7914), .ZN(n7943) );
  AND2_X1 U9082 ( .A1(n8204), .A2(n10458), .ZN(n6708) );
  AND2_X1 U9083 ( .A1(n8206), .A2(n9267), .ZN(n6709) );
  AND2_X1 U9084 ( .A1(n7142), .A2(n6809), .ZN(n6710) );
  INV_X1 U9085 ( .A(n11574), .ZN(n12237) );
  AND4_X1 U9086 ( .A1(n7841), .A2(n7840), .A3(n7839), .A4(n7838), .ZN(n11574)
         );
  INV_X1 U9087 ( .A(n12410), .ZN(n12657) );
  NAND2_X1 U9088 ( .A1(n8084), .A2(n8083), .ZN(n12410) );
  AND2_X1 U9089 ( .A1(n11053), .A2(n7247), .ZN(n6711) );
  INV_X1 U9090 ( .A(n9051), .ZN(n7120) );
  INV_X1 U9091 ( .A(n10458), .ZN(n9267) );
  AND2_X1 U9092 ( .A1(n9150), .A2(n9232), .ZN(n6712) );
  AND2_X1 U9093 ( .A1(n7119), .A2(n6803), .ZN(n6713) );
  OR2_X1 U9094 ( .A1(n7115), .A2(n7113), .ZN(n6714) );
  OR2_X1 U9095 ( .A1(n10440), .A2(n10968), .ZN(n6715) );
  INV_X1 U9096 ( .A(n8456), .ZN(n8706) );
  INV_X1 U9097 ( .A(n6970), .ZN(n14460) );
  NAND2_X1 U9098 ( .A1(n8693), .A2(n8692), .ZN(n6970) );
  INV_X1 U9099 ( .A(n8785), .ZN(n8667) );
  XOR2_X1 U9100 ( .A(n12387), .B(n10209), .Z(n6716) );
  INV_X1 U9101 ( .A(n8899), .ZN(n8850) );
  NOR2_X1 U9102 ( .A1(n9111), .A2(n7482), .ZN(n7481) );
  AND2_X1 U9103 ( .A1(n12586), .A2(n14775), .ZN(n6717) );
  NOR2_X1 U9104 ( .A1(n12365), .A2(n12570), .ZN(n6718) );
  INV_X1 U9105 ( .A(n8838), .ZN(n7278) );
  AND2_X1 U9106 ( .A1(n13360), .A2(n11737), .ZN(n6719) );
  AND2_X1 U9107 ( .A1(n10437), .A2(n10436), .ZN(n6720) );
  INV_X1 U9108 ( .A(n11769), .ZN(n8197) );
  AND2_X1 U9109 ( .A1(n8200), .A2(n8202), .ZN(n11769) );
  OR2_X1 U9110 ( .A1(n9350), .A2(n9351), .ZN(n6721) );
  OR2_X1 U9111 ( .A1(n13879), .A2(n14016), .ZN(n6723) );
  OR2_X1 U9112 ( .A1(n11955), .A2(n6891), .ZN(n6724) );
  AND2_X1 U9113 ( .A1(n8168), .A2(n8172), .ZN(n11077) );
  INV_X1 U9114 ( .A(n8253), .ZN(n7180) );
  AND2_X1 U9115 ( .A1(n7380), .A2(n9203), .ZN(n6725) );
  NAND2_X1 U9116 ( .A1(n7453), .A2(n8219), .ZN(n12525) );
  XNOR2_X1 U9117 ( .A(n12132), .B(n14362), .ZN(n9094) );
  AND2_X1 U9118 ( .A1(n12024), .A2(n14218), .ZN(n6726) );
  NAND2_X1 U9119 ( .A1(n14432), .A2(n8708), .ZN(n14419) );
  XNOR2_X1 U9120 ( .A(n10934), .B(n10961), .ZN(n10813) );
  XNOR2_X1 U9121 ( .A(n13999), .B(n13260), .ZN(n13823) );
  XNOR2_X1 U9122 ( .A(n14567), .B(n14234), .ZN(n14358) );
  NOR2_X1 U9123 ( .A1(n14954), .A2(n11657), .ZN(n6727) );
  OR2_X1 U9124 ( .A1(n13239), .A2(n6616), .ZN(n6728) );
  NAND2_X1 U9125 ( .A1(n12743), .A2(n12742), .ZN(n14022) );
  INV_X1 U9126 ( .A(n14022), .ZN(n7070) );
  NAND2_X1 U9127 ( .A1(n10882), .A2(n10881), .ZN(n13027) );
  INV_X1 U9128 ( .A(n13027), .ZN(n7074) );
  AND2_X1 U9129 ( .A1(n10945), .A2(n10946), .ZN(n6729) );
  AND2_X1 U9130 ( .A1(n6699), .A2(n7694), .ZN(n7774) );
  AND2_X1 U9131 ( .A1(n6973), .A2(n6971), .ZN(n6730) );
  AND3_X1 U9132 ( .A1(n13635), .A2(n13636), .A3(n10190), .ZN(n6731) );
  OR2_X1 U9133 ( .A1(n14435), .A2(n7102), .ZN(n6732) );
  NOR2_X1 U9134 ( .A1(n15447), .A2(n6912), .ZN(n6733) );
  INV_X1 U9135 ( .A(n14696), .ZN(n7262) );
  AND2_X1 U9136 ( .A1(n8441), .A2(n8440), .ZN(n10794) );
  AND2_X1 U9137 ( .A1(n8456), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6734) );
  AND2_X1 U9138 ( .A1(n11798), .A2(n12236), .ZN(n6735) );
  AND2_X1 U9139 ( .A1(n13940), .A2(n6719), .ZN(n6736) );
  AND2_X1 U9140 ( .A1(n7427), .A2(n7425), .ZN(n6737) );
  AND2_X1 U9141 ( .A1(n7441), .A2(n7439), .ZN(n6738) );
  NOR2_X1 U9142 ( .A1(n12398), .A2(n12464), .ZN(n6739) );
  AND2_X1 U9143 ( .A1(n11541), .A2(n11540), .ZN(n14816) );
  INV_X1 U9144 ( .A(n14816), .ZN(n7081) );
  NAND2_X1 U9145 ( .A1(n8511), .A2(n8510), .ZN(n11671) );
  XNOR2_X1 U9146 ( .A(n13380), .B(n13259), .ZN(n13375) );
  INV_X1 U9147 ( .A(n8839), .ZN(n6950) );
  NAND2_X1 U9148 ( .A1(n12132), .A2(n14362), .ZN(n6740) );
  INV_X1 U9149 ( .A(n13132), .ZN(n7364) );
  OR2_X1 U9150 ( .A1(n10041), .A2(n15231), .ZN(n6741) );
  INV_X1 U9151 ( .A(n13104), .ZN(n7354) );
  INV_X1 U9152 ( .A(n7104), .ZN(n14422) );
  NOR2_X1 U9153 ( .A1(n14435), .A2(n14423), .ZN(n7104) );
  AND2_X1 U9154 ( .A1(n9171), .A2(n9170), .ZN(n6742) );
  OR2_X1 U9155 ( .A1(n14886), .A2(n6933), .ZN(n6931) );
  AND2_X1 U9156 ( .A1(n11798), .A2(n11709), .ZN(n6743) );
  AND2_X1 U9157 ( .A1(n13892), .A2(n7576), .ZN(n6744) );
  INV_X1 U9158 ( .A(n7317), .ZN(n7314) );
  NAND2_X1 U9159 ( .A1(n10570), .A2(n7318), .ZN(n7317) );
  OR2_X1 U9160 ( .A1(n7338), .A2(n7337), .ZN(n6745) );
  NAND2_X1 U9161 ( .A1(n14567), .A2(n14211), .ZN(n6746) );
  NAND2_X1 U9162 ( .A1(n7598), .A2(n7527), .ZN(n6747) );
  INV_X1 U9163 ( .A(n13353), .ZN(n13811) );
  AND2_X1 U9164 ( .A1(n12118), .A2(n12117), .ZN(n6748) );
  AND2_X1 U9165 ( .A1(n13064), .A2(n14785), .ZN(n6749) );
  NOR3_X1 U9166 ( .A1(n12591), .A2(n12449), .A3(n9267), .ZN(n6750) );
  OR2_X1 U9167 ( .A1(n6705), .A2(n7417), .ZN(n6751) );
  NOR2_X1 U9168 ( .A1(n14209), .A2(n7430), .ZN(n6752) );
  NOR2_X1 U9169 ( .A1(n14609), .A2(n14134), .ZN(n6753) );
  NOR2_X1 U9170 ( .A1(n14964), .A2(n14898), .ZN(n6754) );
  NOR2_X1 U9171 ( .A1(n10961), .A2(n10934), .ZN(n6755) );
  AND2_X1 U9172 ( .A1(n8837), .A2(n7280), .ZN(n6756) );
  INV_X1 U9173 ( .A(n13371), .ZN(n6981) );
  NAND2_X1 U9174 ( .A1(n10755), .A2(n10756), .ZN(n7316) );
  INV_X1 U9175 ( .A(n11707), .ZN(n7203) );
  INV_X1 U9176 ( .A(n6840), .ZN(n14453) );
  NOR2_X1 U9177 ( .A1(n14473), .A2(n14475), .ZN(n6840) );
  INV_X1 U9178 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n13637) );
  INV_X1 U9179 ( .A(n12125), .ZN(n7431) );
  INV_X1 U9180 ( .A(n7084), .ZN(n13382) );
  NOR2_X1 U9181 ( .A1(n13381), .A2(n13380), .ZN(n7084) );
  AND2_X1 U9182 ( .A1(n8331), .A2(SI_8_), .ZN(n6757) );
  AND2_X1 U9183 ( .A1(n12492), .A2(n8233), .ZN(n6758) );
  INV_X1 U9184 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n8290) );
  AND2_X1 U9185 ( .A1(n15151), .A2(n11408), .ZN(n6759) );
  AND2_X1 U9186 ( .A1(n8240), .A2(n8241), .ZN(n12394) );
  INV_X1 U9187 ( .A(n12394), .ZN(n12462) );
  AND2_X1 U9188 ( .A1(n15192), .A2(n11274), .ZN(n6760) );
  INV_X1 U9189 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8266) );
  NOR2_X1 U9190 ( .A1(n12626), .A2(n12535), .ZN(n6761) );
  INV_X1 U9191 ( .A(n8958), .ZN(n7230) );
  INV_X1 U9192 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8288) );
  INV_X1 U9193 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9503) );
  NAND2_X1 U9194 ( .A1(n8955), .A2(n7230), .ZN(n6762) );
  AND2_X1 U9195 ( .A1(n6891), .A2(n6890), .ZN(n6763) );
  NOR2_X1 U9196 ( .A1(n13819), .A2(n13372), .ZN(n6764) );
  NAND2_X1 U9197 ( .A1(n12433), .A2(n7208), .ZN(n7211) );
  NAND2_X1 U9198 ( .A1(n12095), .A2(n12094), .ZN(n6765) );
  NAND2_X1 U9199 ( .A1(n14423), .A2(n14440), .ZN(n6766) );
  NOR2_X1 U9200 ( .A1(n13394), .A2(n13358), .ZN(n6767) );
  INV_X1 U9201 ( .A(n6892), .ZN(n6891) );
  NAND2_X1 U9202 ( .A1(n14083), .A2(n14209), .ZN(n6768) );
  INV_X1 U9203 ( .A(n9013), .ZN(n7226) );
  OR2_X1 U9204 ( .A1(n7550), .A2(n7552), .ZN(n6769) );
  INV_X1 U9205 ( .A(n8959), .ZN(n7227) );
  INV_X1 U9206 ( .A(n12513), .ZN(n12383) );
  AND2_X1 U9207 ( .A1(n8226), .A2(n8227), .ZN(n12513) );
  NAND2_X1 U9208 ( .A1(n13167), .A2(n13166), .ZN(n13343) );
  INV_X1 U9209 ( .A(n13343), .ZN(n7082) );
  AND2_X1 U9210 ( .A1(n9362), .A2(n9367), .ZN(n6770) );
  NOR2_X1 U9211 ( .A1(n10777), .A2(n6727), .ZN(n6771) );
  INV_X1 U9212 ( .A(n8256), .ZN(n7181) );
  INV_X1 U9213 ( .A(n12447), .ZN(n7465) );
  AND2_X1 U9214 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6772) );
  AND2_X1 U9215 ( .A1(n8572), .A2(n7241), .ZN(n6773) );
  AND2_X1 U9216 ( .A1(n9177), .A2(n9175), .ZN(n6774) );
  OR2_X1 U9217 ( .A1(n7354), .A2(n13103), .ZN(n6775) );
  AND2_X1 U9218 ( .A1(n8289), .A2(n7511), .ZN(n6776) );
  NAND2_X1 U9219 ( .A1(n10062), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n6777) );
  AOI21_X1 U9220 ( .B1(n6700), .B2(n11957), .A(n6763), .ZN(n6889) );
  OR2_X1 U9221 ( .A1(n7364), .A2(n13131), .ZN(n6778) );
  OR2_X1 U9222 ( .A1(n13012), .A2(n13010), .ZN(n6779) );
  OR2_X1 U9223 ( .A1(n12999), .A2(n12997), .ZN(n6780) );
  AND2_X1 U9224 ( .A1(n7578), .A2(n13893), .ZN(n6781) );
  AND2_X1 U9225 ( .A1(n11916), .A2(n11910), .ZN(n6782) );
  OR2_X1 U9226 ( .A1(n13049), .A2(n13051), .ZN(n6783) );
  AND2_X1 U9227 ( .A1(n7492), .A2(n6746), .ZN(n6784) );
  OR2_X1 U9228 ( .A1(n7351), .A2(n13050), .ZN(n6785) );
  NAND2_X1 U9229 ( .A1(n13374), .A2(n13181), .ZN(n13357) );
  AND2_X1 U9230 ( .A1(n6721), .A2(n6920), .ZN(n6787) );
  OR2_X1 U9231 ( .A1(n13011), .A2(n7349), .ZN(n6788) );
  INV_X1 U9232 ( .A(n9206), .ZN(n7380) );
  NAND2_X1 U9233 ( .A1(n8926), .A2(n7232), .ZN(n6790) );
  INV_X1 U9234 ( .A(n6976), .ZN(n6975) );
  NAND2_X1 U9235 ( .A1(n13353), .A2(n6978), .ZN(n6976) );
  OR2_X1 U9236 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n6791) );
  NAND2_X1 U9237 ( .A1(n9014), .A2(n7226), .ZN(n6792) );
  NAND2_X1 U9238 ( .A1(n11586), .A2(n11585), .ZN(n14042) );
  INV_X1 U9239 ( .A(n14042), .ZN(n7079) );
  NAND2_X1 U9240 ( .A1(n11838), .A2(n11837), .ZN(n11839) );
  NAND2_X1 U9241 ( .A1(n6837), .A2(n6695), .ZN(n9413) );
  AND4_X1 U9242 ( .A1(n7890), .A2(n7889), .A3(n7888), .A4(n7887), .ZN(n11727)
         );
  AND2_X1 U9243 ( .A1(n11712), .A2(n8200), .ZN(n6793) );
  INV_X1 U9244 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7096) );
  INV_X1 U9245 ( .A(n7071), .ZN(n13910) );
  NOR2_X1 U9246 ( .A1(n13930), .A2(n14027), .ZN(n7071) );
  INV_X1 U9247 ( .A(n12478), .ZN(n7053) );
  OR2_X1 U9248 ( .A1(n14824), .A2(n14786), .ZN(n6794) );
  AND2_X1 U9249 ( .A1(n12052), .A2(n12051), .ZN(n6795) );
  NAND2_X1 U9250 ( .A1(n11900), .A2(n6854), .ZN(n14848) );
  INV_X1 U9251 ( .A(n13906), .ZN(n13363) );
  AND2_X1 U9252 ( .A1(n7393), .A2(n7392), .ZN(n6796) );
  AND4_X1 U9253 ( .A1(n8014), .A2(n8013), .A3(n8012), .A4(n8011), .ZN(n12203)
         );
  OR2_X1 U9254 ( .A1(n12364), .A2(n7058), .ZN(n6797) );
  NAND2_X1 U9255 ( .A1(n8203), .A2(n8204), .ZN(n6798) );
  NAND2_X1 U9256 ( .A1(n7062), .A2(n7060), .ZN(n6799) );
  AND2_X1 U9257 ( .A1(n10348), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n6800) );
  AND2_X1 U9258 ( .A1(n11712), .A2(n8202), .ZN(n6801) );
  NAND2_X1 U9259 ( .A1(n8201), .A2(n8206), .ZN(n6802) );
  INV_X1 U9260 ( .A(n14531), .ZN(n14526) );
  INV_X1 U9261 ( .A(n15072), .ZN(n13944) );
  INV_X1 U9262 ( .A(n11065), .ZN(n7247) );
  INV_X1 U9263 ( .A(n12651), .ZN(n6853) );
  OR2_X1 U9264 ( .A1(n9050), .A2(SI_29_), .ZN(n6803) );
  AND2_X1 U9265 ( .A1(n10806), .A2(n6698), .ZN(n6804) );
  AND2_X1 U9266 ( .A1(n15380), .A2(n10543), .ZN(n12581) );
  INV_X1 U9267 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n7407) );
  INV_X1 U9268 ( .A(n9041), .ZN(n7117) );
  NOR2_X1 U9269 ( .A1(n15274), .A2(n10641), .ZN(n6805) );
  NOR2_X1 U9270 ( .A1(n11283), .A2(n11284), .ZN(n6806) );
  INV_X1 U9271 ( .A(n9042), .ZN(n7124) );
  AND2_X1 U9272 ( .A1(n7505), .A2(n7507), .ZN(n6807) );
  NOR2_X1 U9273 ( .A1(n11308), .A2(n11307), .ZN(n6808) );
  INV_X1 U9274 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7270) );
  NOR2_X1 U9275 ( .A1(n11882), .A2(n14153), .ZN(n11883) );
  OR2_X1 U9276 ( .A1(n8773), .A2(SI_27_), .ZN(n6809) );
  NAND2_X1 U9277 ( .A1(n11112), .A2(n8523), .ZN(n6810) );
  AND2_X1 U9278 ( .A1(n10905), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n6811) );
  AND3_X1 U9279 ( .A1(n9411), .A2(n9614), .A3(n9410), .ZN(n9426) );
  OR2_X1 U9280 ( .A1(n10740), .A2(n10739), .ZN(n6812) );
  AND2_X1 U9281 ( .A1(n6922), .A2(n6921), .ZN(n6813) );
  INV_X1 U9282 ( .A(n7554), .ZN(n7552) );
  NAND2_X1 U9283 ( .A1(n14042), .A2(n11751), .ZN(n7554) );
  OR2_X1 U9284 ( .A1(n7120), .A2(n7114), .ZN(n6814) );
  OR2_X1 U9285 ( .A1(n7120), .A2(n9042), .ZN(n6815) );
  INV_X1 U9286 ( .A(n14850), .ZN(n14904) );
  NAND2_X1 U9287 ( .A1(n8495), .A2(n8494), .ZN(n14956) );
  INV_X1 U9288 ( .A(n14956), .ZN(n7105) );
  NAND2_X1 U9289 ( .A1(n10094), .A2(n10093), .ZN(n14850) );
  NAND2_X1 U9290 ( .A1(n10230), .A2(n8898), .ZN(n10828) );
  INV_X1 U9291 ( .A(n8900), .ZN(n7223) );
  AND2_X1 U9292 ( .A1(n10174), .A2(n13219), .ZN(n13925) );
  NAND2_X1 U9293 ( .A1(n10955), .A2(n10956), .ZN(n6816) );
  INV_X1 U9294 ( .A(n9858), .ZN(n7097) );
  NOR2_X1 U9295 ( .A1(n15223), .A2(n10060), .ZN(n6817) );
  INV_X1 U9296 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n6863) );
  INV_X1 U9297 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n6928) );
  INV_X1 U9298 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7640) );
  INV_X1 U9299 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6913) );
  AOI21_X1 U9300 ( .B1(n8812), .B2(n14701), .A(n8811), .ZN(n12004) );
  INV_X1 U9301 ( .A(n14701), .ZN(n14603) );
  OR2_X2 U9302 ( .A1(n9664), .A2(n10367), .ZN(n14252) );
  NAND2_X1 U9303 ( .A1(n7846), .A2(n7845), .ZN(n7861) );
  NAND2_X1 U9304 ( .A1(n7191), .A2(n7190), .ZN(n12656) );
  OAI21_X1 U9305 ( .B1(n12444), .B2(n7458), .A(n7456), .ZN(n12409) );
  NAND2_X1 U9306 ( .A1(n7462), .A2(n12447), .ZN(n7460) );
  NAND2_X1 U9307 ( .A1(n7711), .A2(n7710), .ZN(n7730) );
  NAND2_X1 U9308 ( .A1(n7154), .A2(n7677), .ZN(n7690) );
  OAI211_X1 U9309 ( .C1(n7022), .C2(n10428), .A(n8257), .B(n7021), .ZN(n7169)
         );
  AND2_X1 U9310 ( .A1(n7035), .A2(n10458), .ZN(n7029) );
  NAND2_X1 U9311 ( .A1(n7192), .A2(n12407), .ZN(n12585) );
  NAND2_X1 U9312 ( .A1(n11344), .A2(n11343), .ZN(n11521) );
  NAND2_X1 U9313 ( .A1(n12655), .A2(n12707), .ZN(n7191) );
  NAND2_X1 U9314 ( .A1(n11327), .A2(n11326), .ZN(n11328) );
  NAND2_X1 U9315 ( .A1(n11079), .A2(n10864), .ZN(n10866) );
  NAND2_X1 U9316 ( .A1(n12380), .A2(n12379), .ZN(n12522) );
  OAI21_X1 U9317 ( .B1(n15337), .B2(n7214), .A(n7212), .ZN(n10727) );
  INV_X1 U9318 ( .A(n7612), .ZN(n7404) );
  OAI211_X1 U9319 ( .C1(n7200), .C2(n7196), .A(n7195), .B(n12369), .ZN(n12371)
         );
  AOI222_X2 U9320 ( .A1(n15369), .A2(n12436), .B1(n12435), .B2(n15366), .C1(
        n12464), .C2(n12406), .ZN(n12593) );
  XNOR2_X1 U9321 ( .A(n6819), .B(n9389), .ZN(SUB_1596_U4) );
  INV_X1 U9322 ( .A(n7273), .ZN(n9325) );
  NAND2_X1 U9323 ( .A1(n6923), .A2(n6787), .ZN(n6918) );
  NAND2_X1 U9324 ( .A1(n14878), .A2(n9368), .ZN(n14882) );
  NOR2_X1 U9325 ( .A1(n14690), .A2(n14689), .ZN(n14688) );
  NOR2_X1 U9326 ( .A1(n14687), .A2(n14686), .ZN(n14685) );
  NOR2_X1 U9327 ( .A1(n14873), .A2(n14874), .ZN(n9356) );
  NAND2_X1 U9328 ( .A1(n15441), .A2(n15440), .ZN(n15439) );
  OAI21_X1 U9329 ( .B1(n9371), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n14881), .ZN(
        n14887) );
  XOR2_X1 U9330 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n9323), .Z(n9336) );
  NAND3_X1 U9331 ( .A1(n7266), .A2(n7268), .A3(n7265), .ZN(n14880) );
  XNOR2_X1 U9332 ( .A(n9344), .B(n15017), .ZN(n15446) );
  NAND2_X1 U9333 ( .A1(n7163), .A2(n7880), .ZN(n7893) );
  NAND2_X1 U9334 ( .A1(n6720), .A2(n15338), .ZN(n15337) );
  NAND2_X2 U9335 ( .A1(n8151), .A2(n9157), .ZN(n7204) );
  NAND2_X2 U9336 ( .A1(n12244), .A2(n10214), .ZN(n8151) );
  NAND2_X1 U9337 ( .A1(n7008), .A2(n7007), .ZN(n12659) );
  NAND2_X1 U9338 ( .A1(n10725), .A2(n10724), .ZN(n10862) );
  NAND3_X1 U9339 ( .A1(n7211), .A2(n15369), .A3(n12421), .ZN(n12425) );
  NAND3_X1 U9340 ( .A1(n12593), .A2(n12592), .A3(n6823), .ZN(n12661) );
  AND3_X1 U9341 ( .A1(n7629), .A2(n7627), .A3(n7628), .ZN(n6848) );
  OAI21_X1 U9342 ( .B1(n8522), .B2(n7500), .A(n7499), .ZN(n11385) );
  AOI21_X1 U9343 ( .B1(n14536), .B2(n14537), .A(n8641), .ZN(n14515) );
  AOI21_X1 U9344 ( .B1(n10779), .B2(n6771), .A(n6701), .ZN(n10977) );
  AOI21_X1 U9345 ( .B1(n8617), .B2(n8970), .A(n7589), .ZN(n11886) );
  NAND2_X1 U9346 ( .A1(n10268), .A2(n10269), .ZN(n10402) );
  NOR2_X1 U9347 ( .A1(n10005), .A2(n10004), .ZN(n10003) );
  AOI21_X2 U9348 ( .B1(n12937), .B2(n12939), .A(n12938), .ZN(n12914) );
  NAND3_X1 U9349 ( .A1(n6984), .A2(n6695), .A3(n9425), .ZN(n9622) );
  AND2_X1 U9350 ( .A1(n9412), .A2(n6985), .ZN(n6984) );
  NAND2_X1 U9351 ( .A1(n10986), .A2(n10985), .ZN(n11150) );
  NOR2_X1 U9352 ( .A1(n7303), .A2(n9916), .ZN(n9987) );
  INV_X1 U9353 ( .A(n7326), .ZN(n14791) );
  NAND2_X1 U9354 ( .A1(n6681), .A2(n9486), .ZN(n9919) );
  AOI22_X1 U9355 ( .A1(n10126), .A2(n10125), .B1(n10124), .B2(n10123), .ZN(
        n10130) );
  NAND2_X1 U9356 ( .A1(n6829), .A2(n7225), .ZN(n9018) );
  NAND3_X1 U9357 ( .A1(n9011), .A2(n9012), .A3(n6792), .ZN(n6829) );
  MUX2_X1 U9358 ( .A(n10255), .B(n14251), .S(n8918), .Z(n8915) );
  NAND2_X1 U9359 ( .A1(n7234), .A2(n7233), .ZN(n9031) );
  INV_X1 U9360 ( .A(n8447), .ZN(n8322) );
  INV_X1 U9361 ( .A(n8954), .ZN(n8955) );
  OR2_X2 U9362 ( .A1(n10648), .A2(n10647), .ZN(n11054) );
  NOR2_X1 U9363 ( .A1(n15310), .A2(n10644), .ZN(n10648) );
  NOR2_X2 U9364 ( .A1(n15256), .A2(n10066), .ZN(n10069) );
  XNOR2_X1 U9365 ( .A(n10643), .B(n10676), .ZN(n15311) );
  NOR2_X1 U9366 ( .A1(n12255), .A2(n12256), .ZN(n12257) );
  NAND2_X2 U9367 ( .A1(n11093), .A2(n11092), .ZN(n11247) );
  NAND2_X2 U9368 ( .A1(n12520), .A2(n12382), .ZN(n12508) );
  NAND2_X1 U9369 ( .A1(n7215), .A2(n10863), .ZN(n11079) );
  INV_X1 U9370 ( .A(n11569), .ZN(n7200) );
  BUF_X4 U9371 ( .A(n7667), .Z(n8103) );
  NAND2_X1 U9372 ( .A1(n7193), .A2(n15369), .ZN(n7192) );
  NAND2_X1 U9373 ( .A1(n11524), .A2(n11523), .ZN(n11569) );
  INV_X2 U9374 ( .A(n15352), .ZN(n12243) );
  NAND2_X1 U9375 ( .A1(n7815), .A2(n7814), .ZN(n7829) );
  NAND2_X1 U9376 ( .A1(n7781), .A2(n7780), .ZN(n7802) );
  NAND2_X1 U9377 ( .A1(n8255), .A2(n8254), .ZN(n6834) );
  XNOR2_X1 U9378 ( .A(n9375), .B(n7272), .ZN(n14731) );
  NAND2_X1 U9379 ( .A1(n6930), .A2(n6929), .ZN(n9373) );
  NAND2_X1 U9380 ( .A1(n14876), .A2(n6770), .ZN(n7266) );
  INV_X1 U9381 ( .A(n9336), .ZN(n7271) );
  NAND2_X1 U9382 ( .A1(n7558), .A2(n8330), .ZN(n8491) );
  AOI21_X2 U9383 ( .B1(n11379), .B2(n11378), .A(n6759), .ZN(n11411) );
  INV_X1 U9384 ( .A(n7197), .ZN(n7196) );
  NAND2_X2 U9385 ( .A1(n7884), .A2(n7883), .ZN(n11799) );
  NAND2_X1 U9386 ( .A1(n12658), .A2(n12707), .ZN(n7008) );
  OAI21_X2 U9387 ( .B1(n7745), .B2(n7172), .A(n7170), .ZN(n7781) );
  OAI21_X1 U9388 ( .B1(n11411), .B2(n11410), .A(n6870), .ZN(n11380) );
  NAND2_X1 U9389 ( .A1(n8317), .A2(n8316), .ZN(n8435) );
  NAND2_X1 U9390 ( .A1(n6865), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n6864) );
  AND2_X1 U9391 ( .A1(n7288), .A2(n10830), .ZN(n6838) );
  NAND2_X1 U9392 ( .A1(n11136), .A2(n8813), .ZN(n10231) );
  NAND2_X1 U9393 ( .A1(n11108), .A2(n11109), .ZN(n11107) );
  NAND2_X1 U9394 ( .A1(n8827), .A2(n7297), .ZN(n11614) );
  NAND2_X1 U9395 ( .A1(n8310), .A2(n8305), .ZN(n6839) );
  NAND2_X1 U9396 ( .A1(n8833), .A2(n7282), .ZN(n7281) );
  NAND2_X1 U9397 ( .A1(n11229), .A2(n11230), .ZN(n11471) );
  NAND2_X1 U9398 ( .A1(n7204), .A2(n15368), .ZN(n10433) );
  CLKBUF_X1 U9399 ( .A(n15354), .Z(n6846) );
  OAI22_X1 U9400 ( .A1(n12475), .A2(n12393), .B1(n12465), .B2(n12392), .ZN(
        n12460) );
  OR2_X2 U9401 ( .A1(n12460), .A2(n12394), .ZN(n12461) );
  XNOR2_X1 U9402 ( .A(n12401), .B(n7194), .ZN(n7193) );
  XNOR2_X2 U9403 ( .A(n7649), .B(n15365), .ZN(n15349) );
  NAND2_X2 U9404 ( .A1(n7626), .A2(n6848), .ZN(n15365) );
  NAND2_X1 U9405 ( .A1(n14791), .A2(n14792), .ZN(n14790) );
  NAND2_X1 U9406 ( .A1(n11781), .A2(n11782), .ZN(n11838) );
  OAI21_X2 U9407 ( .B1(n10402), .B2(n7311), .A(n7310), .ZN(n10762) );
  NAND2_X1 U9408 ( .A1(n12374), .A2(n7221), .ZN(n12547) );
  NAND2_X1 U9409 ( .A1(n7211), .A2(n7210), .ZN(n12401) );
  NAND2_X1 U9410 ( .A1(n7371), .A2(n7370), .ZN(n11852) );
  XNOR2_X1 U9411 ( .A(n12781), .B(n12769), .ZN(n12949) );
  OAI22_X1 U9412 ( .A1(n9919), .A2(n9918), .B1(n6681), .B2(n9917), .ZN(n9922)
         );
  NAND4_X2 U9413 ( .A1(n7613), .A2(n7188), .A3(n6722), .A4(n7469), .ZN(n7635)
         );
  NAND2_X1 U9414 ( .A1(n7643), .A2(n6863), .ZN(n6862) );
  NAND2_X1 U9415 ( .A1(n7557), .A2(n7556), .ZN(n8506) );
  NAND2_X1 U9416 ( .A1(n6868), .A2(n9003), .ZN(n9008) );
  NOR2_X1 U9417 ( .A1(n11056), .A2(n11055), .ZN(n11222) );
  NAND2_X1 U9418 ( .A1(n12957), .A2(n12843), .ZN(n12890) );
  NOR2_X1 U9419 ( .A1(n11469), .A2(n11470), .ZN(n12255) );
  NOR2_X1 U9420 ( .A1(n12257), .A2(n12258), .ZN(n12274) );
  NAND2_X1 U9421 ( .A1(n10762), .A2(n10761), .ZN(n10917) );
  OAI22_X1 U9422 ( .A1(n12914), .A2(n12913), .B1(n12765), .B2(n12764), .ZN(
        n12781) );
  OAI21_X1 U9423 ( .B1(n9990), .B2(n9987), .A(n9988), .ZN(n10005) );
  NAND2_X1 U9424 ( .A1(n6873), .A2(n12031), .ZN(n14156) );
  INV_X1 U9425 ( .A(n8324), .ZN(n7134) );
  NAND2_X1 U9426 ( .A1(n8727), .A2(n8726), .ZN(n14403) );
  NAND2_X1 U9427 ( .A1(n7109), .A2(n7107), .ZN(n14645) );
  NAND2_X2 U9428 ( .A1(n8386), .A2(n8385), .ZN(n12005) );
  NOR2_X4 U9429 ( .A1(n8866), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n8387) );
  OR2_X1 U9430 ( .A1(n10148), .A2(n10149), .ZN(n10150) );
  NAND2_X1 U9431 ( .A1(n12345), .A2(n12344), .ZN(n6859) );
  INV_X1 U9432 ( .A(n12343), .ZN(n6860) );
  NAND2_X1 U9433 ( .A1(n7466), .A2(n7465), .ZN(n7464) );
  NAND2_X1 U9434 ( .A1(n11328), .A2(n11336), .ZN(n11344) );
  NAND2_X1 U9435 ( .A1(n11249), .A2(n11248), .ZN(n11327) );
  NAND2_X1 U9436 ( .A1(n12479), .A2(n8235), .ZN(n12459) );
  AOI21_X1 U9437 ( .B1(n12491), .B2(n8234), .A(n7470), .ZN(n12480) );
  NAND2_X1 U9438 ( .A1(n12433), .A2(n12400), .ZN(n12420) );
  NAND2_X1 U9439 ( .A1(n12502), .A2(n8231), .ZN(n7997) );
  INV_X1 U9440 ( .A(n7006), .ZN(n11770) );
  NAND2_X1 U9441 ( .A1(n7030), .A2(n8252), .ZN(n7024) );
  NAND2_X1 U9442 ( .A1(n7709), .A2(n7708), .ZN(n7711) );
  NAND2_X1 U9443 ( .A1(n7730), .A2(n7729), .ZN(n7732) );
  NAND2_X1 U9444 ( .A1(n7169), .A2(n8263), .ZN(n7168) );
  NAND2_X1 U9445 ( .A1(n7804), .A2(n7803), .ZN(n7807) );
  NAND2_X1 U9446 ( .A1(n7831), .A2(n7830), .ZN(n7844) );
  NAND3_X1 U9447 ( .A1(n7642), .A2(n7641), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n6865) );
  NAND2_X1 U9448 ( .A1(n7555), .A2(n8322), .ZN(n7133) );
  NOR2_X1 U9449 ( .A1(n14014), .A2(n6871), .ZN(n13840) );
  NAND2_X2 U9450 ( .A1(n13810), .A2(n7592), .ZN(n13802) );
  INV_X1 U9451 ( .A(n9004), .ZN(n6868) );
  NAND2_X1 U9452 ( .A1(n9008), .A2(n9007), .ZN(n9010) );
  NAND2_X1 U9453 ( .A1(n15247), .A2(n15246), .ZN(n15245) );
  NAND2_X1 U9454 ( .A1(n15328), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n15327) );
  NAND2_X1 U9455 ( .A1(n11227), .A2(n11228), .ZN(n11229) );
  NAND2_X1 U9456 ( .A1(n11059), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n11227) );
  NAND2_X1 U9457 ( .A1(n6876), .A2(n7406), .ZN(n8864) );
  AOI21_X2 U9458 ( .B1(n8392), .B2(n8393), .A(n8309), .ZN(n8418) );
  AND2_X2 U9459 ( .A1(n13868), .A2(n13867), .ZN(n14014) );
  NAND2_X1 U9460 ( .A1(n10862), .A2(n10861), .ZN(n11078) );
  NOR2_X2 U9463 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n6878) );
  NOR2_X1 U9464 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n6879) );
  NAND2_X1 U9465 ( .A1(n6751), .A2(n7416), .ZN(n7413) );
  NAND3_X1 U9466 ( .A1(n6751), .A2(n7416), .A3(n11662), .ZN(n6883) );
  INV_X1 U9467 ( .A(n6882), .ZN(n14077) );
  NAND2_X1 U9468 ( .A1(n11956), .A2(n6700), .ZN(n6888) );
  OAI211_X1 U9469 ( .C1(n11956), .C2(n6706), .A(n6888), .B(n6889), .ZN(n14895)
         );
  NOR2_X1 U9470 ( .A1(n11956), .A2(n11957), .ZN(n11955) );
  AOI22_X2 U9471 ( .A1(n6724), .A2(n11673), .B1(n14895), .B2(n14894), .ZN(
        n11679) );
  NAND2_X1 U9472 ( .A1(n11668), .A2(n11669), .ZN(n6892) );
  NAND2_X1 U9473 ( .A1(n14208), .A2(n6894), .ZN(n6893) );
  OAI211_X1 U9474 ( .C1(n14208), .C2(n6895), .A(n14089), .B(n6893), .ZN(
        P1_U3214) );
  NAND2_X1 U9475 ( .A1(n14176), .A2(n14175), .ZN(n14174) );
  OAI21_X1 U9476 ( .B1(n14176), .B2(n6905), .A(n6903), .ZN(n14139) );
  NAND2_X1 U9477 ( .A1(n6902), .A2(n6900), .ZN(n12104) );
  NAND2_X1 U9478 ( .A1(n14176), .A2(n6903), .ZN(n6902) );
  NOR2_X1 U9479 ( .A1(n6910), .A2(n6734), .ZN(n6909) );
  AOI21_X1 U9480 ( .B1(n15448), .B2(n15449), .A(n6913), .ZN(n6912) );
  NOR2_X1 U9481 ( .A1(n15448), .A2(n15449), .ZN(n15447) );
  NAND2_X1 U9482 ( .A1(n14682), .A2(n14683), .ZN(n14681) );
  OAI21_X1 U9483 ( .B1(n14682), .B2(n14683), .A(n6915), .ZN(n6914) );
  INV_X1 U9484 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n6915) );
  NAND2_X1 U9485 ( .A1(n14731), .A2(n14730), .ZN(n14729) );
  NAND2_X1 U9486 ( .A1(n14889), .A2(n14891), .ZN(n9375) );
  INV_X1 U9487 ( .A(n14688), .ZN(n6923) );
  INV_X1 U9488 ( .A(n14881), .ZN(n6925) );
  OAI211_X1 U9489 ( .C1(n9371), .C2(n6927), .A(n6926), .B(n6924), .ZN(n14892)
         );
  INV_X1 U9490 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n6933) );
  NAND2_X1 U9491 ( .A1(n14364), .A2(n6935), .ZN(n6938) );
  NAND2_X1 U9492 ( .A1(n7132), .A2(n8327), .ZN(n6940) );
  NAND3_X1 U9493 ( .A1(n6940), .A2(n7559), .A3(n6939), .ZN(n7557) );
  NAND3_X1 U9494 ( .A1(n6941), .A2(n8327), .A3(n8321), .ZN(n6939) );
  NAND2_X1 U9495 ( .A1(n6946), .A2(n6943), .ZN(n8841) );
  NAND2_X1 U9496 ( .A1(n14447), .A2(n8839), .ZN(n14428) );
  NAND2_X1 U9497 ( .A1(n6951), .A2(n6952), .ZN(n14447) );
  NAND2_X1 U9498 ( .A1(n7276), .A2(n6953), .ZN(n14580) );
  NAND2_X1 U9499 ( .A1(n6957), .A2(n6956), .ZN(n6955) );
  NAND2_X1 U9500 ( .A1(n7151), .A2(n6963), .ZN(n6961) );
  NAND3_X1 U9501 ( .A1(n9425), .A2(n6695), .A3(n9412), .ZN(n9535) );
  AOI21_X1 U9502 ( .B1(n13411), .B2(n7598), .A(n13925), .ZN(n6988) );
  NAND2_X1 U9503 ( .A1(n6989), .A2(n9165), .ZN(n9163) );
  NAND2_X1 U9504 ( .A1(n8135), .A2(n8151), .ZN(n6989) );
  INV_X2 U9505 ( .A(n10187), .ZN(n11950) );
  NAND2_X1 U9507 ( .A1(n7442), .A2(n8168), .ZN(n6995) );
  NAND2_X1 U9508 ( .A1(n6995), .A2(n6994), .ZN(n7758) );
  OAI21_X1 U9509 ( .B1(n12545), .B2(n7000), .A(n6997), .ZN(n12502) );
  OAI21_X1 U9510 ( .B1(n11527), .B2(n7002), .A(n7001), .ZN(n7006) );
  AOI21_X2 U9511 ( .B1(n12459), .B2(n12394), .A(n7009), .ZN(n7466) );
  AOI21_X1 U9512 ( .B1(n8155), .B2(n9157), .A(n7018), .ZN(n7017) );
  NAND3_X1 U9513 ( .A1(n7027), .A2(n7025), .A3(n7023), .ZN(n8255) );
  INV_X1 U9514 ( .A(n7029), .ZN(n7026) );
  NAND2_X1 U9515 ( .A1(n8248), .A2(n7031), .ZN(n7027) );
  OR2_X1 U9516 ( .A1(n8229), .A2(n7044), .ZN(n7041) );
  NAND2_X1 U9517 ( .A1(n7041), .A2(n7042), .ZN(n8244) );
  OR2_X1 U9518 ( .A1(n8205), .A2(n7057), .ZN(n7055) );
  NAND2_X1 U9519 ( .A1(n7055), .A2(n7056), .ZN(n8216) );
  NOR2_X2 U9520 ( .A1(n6723), .A2(n14010), .ZN(n13861) );
  NAND2_X1 U9521 ( .A1(n7076), .A2(n7072), .ZN(n11181) );
  MUX2_X1 U9522 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n14974), .S(n9458), .Z(n9454)
         );
  NOR2_X2 U9523 ( .A1(n14710), .A2(n14707), .ZN(n14711) );
  NOR2_X2 U9524 ( .A1(n14534), .A2(n14620), .ZN(n14524) );
  INV_X1 U9525 ( .A(n14939), .ZN(n7099) );
  MUX2_X1 U9526 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n9910), .Z(n8319) );
  INV_X1 U9527 ( .A(n9043), .ZN(n7118) );
  OAI21_X1 U9528 ( .B1(n9043), .B2(n6814), .A(n6714), .ZN(n7110) );
  OAI21_X1 U9529 ( .B1(n9043), .B2(n6815), .A(n6713), .ZN(n7121) );
  NAND2_X1 U9530 ( .A1(n7133), .A2(n8324), .ZN(n8466) );
  NAND4_X1 U9531 ( .A1(n7135), .A2(n13239), .A3(n13244), .A4(n7140), .ZN(n7138) );
  OAI211_X1 U9532 ( .C1(n13213), .C2(n13331), .A(n7138), .B(n7136), .ZN(n13216) );
  NAND2_X1 U9533 ( .A1(n7137), .A2(n13214), .ZN(n7136) );
  NAND3_X1 U9534 ( .A1(n7140), .A2(n13375), .A3(n13212), .ZN(n7137) );
  INV_X1 U9535 ( .A(n13213), .ZN(n13221) );
  OAI21_X1 U9536 ( .B1(n8747), .B2(n8746), .A(n8745), .ZN(n8760) );
  AOI21_X1 U9537 ( .B1(n8746), .B2(n8745), .A(SI_26_), .ZN(n7146) );
  INV_X1 U9538 ( .A(n7664), .ZN(n7152) );
  NAND2_X1 U9539 ( .A1(n7152), .A2(n7656), .ZN(n7645) );
  NAND2_X1 U9540 ( .A1(n7690), .A2(n7689), .ZN(n7153) );
  NAND2_X1 U9541 ( .A1(n7676), .A2(n7675), .ZN(n7154) );
  NAND2_X1 U9542 ( .A1(n7941), .A2(n7158), .ZN(n7156) );
  NAND2_X1 U9543 ( .A1(n7879), .A2(n7164), .ZN(n7162) );
  NAND3_X1 U9544 ( .A1(n7168), .A2(n7167), .A3(n8278), .ZN(P3_U3296) );
  OAI21_X2 U9545 ( .B1(n8053), .B2(n8052), .A(n8054), .ZN(n8066) );
  NAND3_X1 U9546 ( .A1(n7181), .A2(n7180), .A3(n7176), .ZN(n7175) );
  OR2_X1 U9547 ( .A1(n12707), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n7190) );
  OAI21_X1 U9548 ( .B1(n7204), .B2(n8152), .A(n9157), .ZN(n8153) );
  XNOR2_X1 U9549 ( .A(n15368), .B(n7204), .ZN(n15370) );
  AND2_X1 U9550 ( .A1(n10209), .A2(n7204), .ZN(n7205) );
  XNOR2_X1 U9551 ( .A(n8135), .B(n7204), .ZN(n15382) );
  NOR2_X1 U9552 ( .A1(n11092), .A2(n7204), .ZN(n7207) );
  OR2_X2 U9553 ( .A1(n12432), .A2(n7040), .ZN(n12433) );
  INV_X1 U9554 ( .A(n11078), .ZN(n7215) );
  NAND2_X1 U9555 ( .A1(n12508), .A2(n7219), .ZN(n7216) );
  NAND2_X1 U9556 ( .A1(n12547), .A2(n12378), .ZN(n12380) );
  OR2_X1 U9557 ( .A1(n9070), .A2(n7223), .ZN(n7222) );
  NAND2_X1 U9558 ( .A1(n9070), .A2(n9089), .ZN(n7224) );
  XNOR2_X1 U9559 ( .A(n8899), .B(n14334), .ZN(n9070) );
  INV_X1 U9560 ( .A(n9018), .ZN(n9021) );
  NAND2_X1 U9561 ( .A1(n8930), .A2(n8931), .ZN(n8929) );
  INV_X1 U9562 ( .A(n9029), .ZN(n7235) );
  NAND2_X1 U9563 ( .A1(n7237), .A2(n7239), .ZN(n8940) );
  NAND3_X1 U9564 ( .A1(n8935), .A2(n7238), .A3(n8934), .ZN(n7237) );
  OR2_X1 U9565 ( .A1(n8938), .A2(n8936), .ZN(n7238) );
  NAND2_X1 U9566 ( .A1(n8938), .A2(n8936), .ZN(n7239) );
  NAND3_X1 U9567 ( .A1(n7244), .A2(n7243), .A3(n7245), .ZN(n11056) );
  NAND2_X1 U9568 ( .A1(n11054), .A2(n6711), .ZN(n7243) );
  XNOR2_X2 U9569 ( .A(n10640), .B(n10673), .ZN(n15276) );
  XNOR2_X2 U9570 ( .A(n12309), .B(n14753), .ZN(n14761) );
  INV_X1 U9571 ( .A(n15224), .ZN(n7258) );
  NAND3_X1 U9572 ( .A1(n7256), .A2(n7255), .A3(n6777), .ZN(n10065) );
  INV_X1 U9573 ( .A(n15236), .ZN(n7259) );
  NOR2_X2 U9574 ( .A1(n14762), .A2(n14761), .ZN(n14763) );
  AOI21_X1 U9575 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n15296), .A(n15299), .ZN(
        n10643) );
  NAND2_X1 U9576 ( .A1(n10065), .A2(n10064), .ZN(n10063) );
  NAND2_X1 U9577 ( .A1(n11468), .A2(n12260), .ZN(n12254) );
  AOI21_X2 U9578 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n10651), .A(n10639), .ZN(
        n10640) );
  NOR2_X2 U9579 ( .A1(n10069), .A2(n10068), .ZN(n10639) );
  AND2_X4 U9580 ( .A1(n8405), .A2(n9794), .ZN(n8541) );
  NOR2_X4 U9581 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n10052) );
  INV_X1 U9582 ( .A(n15349), .ZN(n10434) );
  NOR2_X1 U9583 ( .A1(n11225), .A2(n11224), .ZN(n11467) );
  NOR2_X1 U9584 ( .A1(n15257), .A2(n15258), .ZN(n15256) );
  AOI21_X1 U9585 ( .B1(n6661), .B2(n9002), .A(n9001), .ZN(n9004) );
  AND2_X4 U9586 ( .A1(n8297), .A2(n8296), .ZN(n8785) );
  NOR2_X2 U9587 ( .A1(n11412), .A2(n14830), .ZN(n11414) );
  NOR2_X1 U9588 ( .A1(n8909), .A2(n8908), .ZN(n8912) );
  NAND2_X1 U9589 ( .A1(n7829), .A2(n7828), .ZN(n7831) );
  NAND2_X1 U9590 ( .A1(n7802), .A2(n7801), .ZN(n7804) );
  NAND2_X1 U9591 ( .A1(n7909), .A2(n7908), .ZN(n7911) );
  NAND2_X1 U9592 ( .A1(n8145), .A2(n9154), .ZN(n8257) );
  XNOR2_X2 U9593 ( .A(n7630), .B(P3_IR_REG_2__SCAN_IN), .ZN(n10050) );
  INV_X1 U9594 ( .A(n7263), .ZN(n14695) );
  INV_X1 U9595 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7264) );
  NAND2_X1 U9596 ( .A1(n14877), .A2(n7267), .ZN(n7265) );
  OAI21_X1 U9597 ( .B1(n9326), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6707), .ZN(
        n7273) );
  INV_X1 U9598 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n7275) );
  NAND2_X1 U9599 ( .A1(n14405), .A2(n14406), .ZN(n7276) );
  NAND2_X1 U9600 ( .A1(n11107), .A2(n7292), .ZN(n7291) );
  NAND2_X1 U9601 ( .A1(n7291), .A2(n7294), .ZN(n8823) );
  NAND2_X1 U9602 ( .A1(n11614), .A2(n8828), .ZN(n11814) );
  NAND2_X2 U9603 ( .A1(n8405), .A2(n9486), .ZN(n9057) );
  NAND2_X1 U9604 ( .A1(n14380), .A2(n7301), .ZN(n14364) );
  NAND2_X1 U9605 ( .A1(n7303), .A2(n9916), .ZN(n9988) );
  NAND2_X1 U9606 ( .A1(n12872), .A2(n7307), .ZN(n7304) );
  INV_X1 U9607 ( .A(n7306), .ZN(n7305) );
  INV_X1 U9608 ( .A(n12929), .ZN(n7308) );
  NAND2_X1 U9609 ( .A1(n7309), .A2(n12795), .ZN(n12930) );
  NAND2_X1 U9610 ( .A1(n12872), .A2(n12873), .ZN(n7309) );
  AOI21_X1 U9611 ( .B1(n11839), .B2(n7322), .A(n7320), .ZN(n7319) );
  INV_X1 U9612 ( .A(n7319), .ZN(n12740) );
  OAI21_X1 U9613 ( .B1(n11301), .B2(n7329), .A(n7327), .ZN(n7326) );
  AOI21_X1 U9614 ( .B1(n7328), .B2(n11623), .A(n7333), .ZN(n7327) );
  OR2_X1 U9615 ( .A1(n7330), .A2(n7332), .ZN(n7329) );
  NAND2_X1 U9616 ( .A1(n12828), .A2(n7338), .ZN(n12957) );
  NAND2_X1 U9617 ( .A1(n13120), .A2(n13119), .ZN(n13118) );
  OAI22_X2 U9618 ( .A1(n13143), .A2(n7346), .B1(n13142), .B2(n7345), .ZN(
        n13146) );
  NAND3_X1 U9619 ( .A1(n13008), .A2(n13007), .A3(n6779), .ZN(n7348) );
  NAND2_X1 U9620 ( .A1(n7348), .A2(n6788), .ZN(n13016) );
  NAND2_X1 U9621 ( .A1(n7350), .A2(n6785), .ZN(n13055) );
  NAND3_X1 U9622 ( .A1(n13048), .A2(n13047), .A3(n6783), .ZN(n7350) );
  NAND2_X1 U9623 ( .A1(n7352), .A2(n7353), .ZN(n13107) );
  NAND3_X1 U9624 ( .A1(n13101), .A2(n13102), .A3(n6775), .ZN(n7352) );
  OAI22_X2 U9625 ( .A1(n13024), .A2(n7356), .B1(n13025), .B2(n7355), .ZN(
        n13030) );
  NAND2_X1 U9626 ( .A1(n13030), .A2(n13031), .ZN(n13029) );
  OAI22_X2 U9627 ( .A1(n13037), .A2(n7358), .B1(n13038), .B2(n7357), .ZN(
        n13043) );
  NAND2_X1 U9628 ( .A1(n13043), .A2(n13044), .ZN(n13042) );
  NAND3_X1 U9629 ( .A1(n12996), .A2(n12995), .A3(n6780), .ZN(n7359) );
  NAND2_X1 U9630 ( .A1(n7359), .A2(n7360), .ZN(n13003) );
  NAND3_X1 U9631 ( .A1(n13130), .A2(n13129), .A3(n6778), .ZN(n7362) );
  NAND2_X1 U9632 ( .A1(n7362), .A2(n7363), .ZN(n13135) );
  NAND3_X1 U9633 ( .A1(n7365), .A2(n12984), .A3(n12983), .ZN(n7367) );
  NAND2_X1 U9634 ( .A1(n7367), .A2(n7366), .ZN(n12991) );
  OR2_X1 U9635 ( .A1(n12986), .A2(n7368), .ZN(n7366) );
  AND2_X2 U9636 ( .A1(n10168), .A2(n13174), .ZN(n12969) );
  AND2_X2 U9637 ( .A1(n9906), .A2(n13214), .ZN(n13174) );
  XNOR2_X2 U9638 ( .A(n9617), .B(n9616), .ZN(n10168) );
  NAND2_X1 U9639 ( .A1(n11509), .A2(n7375), .ZN(n7371) );
  NAND2_X1 U9640 ( .A1(n12164), .A2(n9228), .ZN(n12219) );
  INV_X1 U9641 ( .A(n9390), .ZN(n9393) );
  NAND3_X2 U9642 ( .A1(n7385), .A2(n12203), .A3(n12182), .ZN(n12183) );
  NAND2_X2 U9643 ( .A1(n9220), .A2(n9219), .ZN(n12182) );
  NAND2_X2 U9644 ( .A1(n7384), .A2(n7386), .ZN(n7385) );
  INV_X1 U9645 ( .A(n9220), .ZN(n7384) );
  AOI21_X2 U9646 ( .B1(n12183), .B2(n12182), .A(n12181), .ZN(n12185) );
  OAI21_X1 U9647 ( .B1(n12146), .B2(n7390), .A(n7387), .ZN(n7399) );
  INV_X1 U9648 ( .A(n7399), .ZN(n9216) );
  OR2_X1 U9649 ( .A1(n9213), .A2(n12535), .ZN(n7400) );
  NAND2_X1 U9650 ( .A1(n7401), .A2(n6774), .ZN(n15205) );
  NOR2_X1 U9651 ( .A1(n7612), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n7402) );
  AND2_X2 U9652 ( .A1(n8120), .A2(n7404), .ZN(n7613) );
  NAND4_X1 U9653 ( .A1(n7469), .A2(n7403), .A3(n6699), .A4(n7694), .ZN(n8259)
         );
  NAND3_X1 U9654 ( .A1(n9150), .A2(n9232), .A3(n9151), .ZN(n9153) );
  AND2_X1 U9655 ( .A1(n7408), .A2(n7407), .ZN(n7405) );
  INV_X1 U9656 ( .A(n12024), .ZN(n7411) );
  OAI21_X1 U9657 ( .B1(n7414), .B2(n10740), .A(n7413), .ZN(n11663) );
  NAND2_X1 U9658 ( .A1(n10740), .A2(n10739), .ZN(n10928) );
  INV_X1 U9659 ( .A(n10739), .ZN(n7417) );
  OAI211_X1 U9660 ( .C1(n14208), .C2(n7426), .A(n7423), .B(n7421), .ZN(n12134)
         );
  NAND2_X1 U9661 ( .A1(n14208), .A2(n7422), .ZN(n7421) );
  NAND2_X1 U9662 ( .A1(n7431), .A2(n7427), .ZN(n7424) );
  NAND2_X1 U9663 ( .A1(n14852), .A2(n6782), .ZN(n11926) );
  NAND2_X1 U9664 ( .A1(n7793), .A2(n7792), .ZN(n11337) );
  NAND2_X1 U9665 ( .A1(n12545), .A2(n8207), .ZN(n12537) );
  INV_X1 U9666 ( .A(n8207), .ZN(n7455) );
  NOR2_X2 U9667 ( .A1(n7039), .A2(n7463), .ZN(n7462) );
  XNOR2_X1 U9668 ( .A(n8113), .B(n9145), .ZN(n7468) );
  NOR2_X1 U9669 ( .A1(n7777), .A2(n7608), .ZN(n7866) );
  NAND2_X1 U9670 ( .A1(n15350), .A2(n15349), .ZN(n15348) );
  NAND2_X1 U9671 ( .A1(n7475), .A2(n7480), .ZN(n14463) );
  NAND2_X1 U9672 ( .A1(n14494), .A2(n7481), .ZN(n7475) );
  AOI21_X1 U9673 ( .B1(n7480), .B2(n7478), .A(n7477), .ZN(n7476) );
  INV_X1 U9674 ( .A(n7481), .ZN(n7478) );
  INV_X1 U9675 ( .A(n7480), .ZN(n7479) );
  NAND2_X1 U9676 ( .A1(n7484), .A2(n7485), .ZN(n8725) );
  NAND2_X1 U9677 ( .A1(n14434), .A2(n8708), .ZN(n7484) );
  OAI21_X1 U9678 ( .B1(n14698), .B2(n7489), .A(n7487), .ZN(n11606) );
  INV_X1 U9679 ( .A(n11606), .ZN(n8617) );
  OR2_X1 U9680 ( .A1(n14388), .A2(n7498), .ZN(n7491) );
  AND2_X2 U9681 ( .A1(n7493), .A2(n6784), .ZN(n11967) );
  OAI21_X1 U9682 ( .B1(n10621), .B2(n7503), .A(n7502), .ZN(n10778) );
  AND2_X1 U9683 ( .A1(n7506), .A2(n7508), .ZN(n7505) );
  INV_X1 U9684 ( .A(n10813), .ZN(n7506) );
  NAND2_X1 U9685 ( .A1(n8387), .A2(n7510), .ZN(n7512) );
  OAI211_X1 U9686 ( .C1(n8311), .C2(n7515), .A(n7514), .B(n8314), .ZN(n8317)
         );
  NAND2_X1 U9687 ( .A1(n8418), .A2(n8313), .ZN(n7514) );
  NAND2_X1 U9688 ( .A1(n13411), .A2(n7519), .ZN(n7518) );
  OAI211_X1 U9689 ( .C1(n13411), .C2(n7520), .A(n13379), .B(n7518), .ZN(n13973) );
  INV_X1 U9690 ( .A(n13375), .ZN(n7527) );
  NAND2_X1 U9691 ( .A1(n7532), .A2(n7533), .ZN(n13359) );
  NAND2_X1 U9692 ( .A1(n13802), .A2(n7535), .ZN(n7532) );
  NAND2_X1 U9693 ( .A1(n13802), .A2(n13355), .ZN(n7539) );
  CLKBUF_X1 U9694 ( .A(n11738), .Z(n7546) );
  NAND2_X1 U9695 ( .A1(n8478), .A2(n8328), .ZN(n7558) );
  INV_X1 U9696 ( .A(n11754), .ZN(n7562) );
  INV_X1 U9697 ( .A(n7572), .ZN(n13854) );
  NAND2_X1 U9698 ( .A1(n13894), .A2(n6781), .ZN(n7573) );
  NAND2_X1 U9699 ( .A1(n7573), .A2(n7574), .ZN(n13868) );
  INV_X1 U9700 ( .A(n8405), .ZN(n8437) );
  NAND2_X1 U9701 ( .A1(n14565), .A2(n14973), .ZN(n8897) );
  NAND2_X1 U9702 ( .A1(n13151), .A2(n13150), .ZN(n13154) );
  NOR2_X1 U9703 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n9323), .ZN(n9292) );
  AND2_X4 U9704 ( .A1(n7625), .A2(n7623), .ZN(n8085) );
  XNOR2_X2 U9705 ( .A(n7654), .B(n7655), .ZN(n10162) );
  CLKBUF_X1 U9706 ( .A(n8264), .Z(n12354) );
  OAI21_X1 U9707 ( .B1(n14364), .B2(n14959), .A(n14363), .ZN(n14365) );
  NAND2_X1 U9708 ( .A1(n9430), .A2(n14674), .ZN(n8409) );
  INV_X1 U9709 ( .A(n13199), .ZN(n11378) );
  NAND4_X2 U9710 ( .A1(n8427), .A2(n8426), .A3(n8425), .A4(n8424), .ZN(n14250)
         );
  INV_X1 U9711 ( .A(n8907), .ZN(n8908) );
  OR2_X1 U9712 ( .A1(n11537), .A2(n7674), .ZN(n8070) );
  OR2_X1 U9713 ( .A1(n11964), .A2(n8847), .ZN(n11999) );
  AOI22_X2 U9714 ( .A1(n12175), .A2(n12174), .B1(n9210), .B2(n12372), .ZN(
        n12211) );
  OAI222_X1 U9715 ( .A1(n14668), .A2(n13165), .B1(P1_U3086), .B2(n8295), .C1(
        n11986), .C2(n12137), .ZN(P1_U3325) );
  AND2_X2 U9716 ( .A1(n8295), .A2(n14671), .ZN(n8455) );
  XNOR2_X1 U9717 ( .A(n10746), .B(n10939), .ZN(n10622) );
  OAI22_X2 U9718 ( .A1(n12211), .A2(n12210), .B1(n12534), .B2(n9211), .ZN(
        n12146) );
  AND2_X1 U9719 ( .A1(n9278), .A2(n15193), .ZN(n7580) );
  AND4_X1 U9720 ( .A1(n8658), .A2(n13492), .A3(n13629), .A4(n8657), .ZN(n7581)
         );
  OR2_X1 U9721 ( .A1(n13850), .A2(n13368), .ZN(n7582) );
  AND2_X1 U9722 ( .A1(n8997), .A2(n8989), .ZN(n7585) );
  NOR2_X1 U9723 ( .A1(n8616), .A2(n11817), .ZN(n7589) );
  AND4_X1 U9724 ( .A1(n8260), .A2(n7615), .A3(n8266), .A4(n7614), .ZN(n7590)
         );
  OR2_X1 U9725 ( .A1(n14568), .A2(n14947), .ZN(n7591) );
  OR2_X1 U9726 ( .A1(n13819), .A2(n13791), .ZN(n7592) );
  NOR2_X1 U9727 ( .A1(n13829), .A2(n13828), .ZN(n7593) );
  OR2_X1 U9728 ( .A1(n13827), .A2(n13370), .ZN(n7594) );
  INV_X1 U9729 ( .A(n9094), .ZN(n8790) );
  INV_X1 U9730 ( .A(n10968), .ZN(n8263) );
  INV_X1 U9731 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n7794) );
  NAND4_X1 U9732 ( .A1(n8789), .A2(n8788), .A3(n8787), .A4(n8786), .ZN(n14362)
         );
  INV_X1 U9733 ( .A(n14362), .ZN(n11965) );
  NAND2_X1 U9734 ( .A1(n9267), .A2(n8265), .ZN(n15353) );
  INV_X1 U9735 ( .A(n10932), .ZN(n10252) );
  AND2_X1 U9736 ( .A1(n8345), .A2(n8344), .ZN(n7596) );
  OR2_X1 U9737 ( .A1(n8684), .A2(SI_20_), .ZN(n7597) );
  AND2_X1 U9738 ( .A1(n6614), .A2(n13390), .ZN(n7598) );
  INV_X1 U9739 ( .A(n14358), .ZN(n8845) );
  OR2_X1 U9740 ( .A1(n8689), .A2(SI_21_), .ZN(n7600) );
  INV_X1 U9741 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n8410) );
  INV_X1 U9742 ( .A(n12878), .ZN(n12736) );
  AOI22_X1 U9743 ( .A1(n10246), .A2(n12119), .B1(n12073), .B2(n14125), .ZN(
        n10248) );
  OR2_X1 U9744 ( .A1(n13336), .A2(n13335), .ZN(P2_U3233) );
  INV_X1 U9745 ( .A(n14550), .ZN(n8853) );
  INV_X1 U9746 ( .A(n10246), .ZN(n8910) );
  NAND2_X1 U9747 ( .A1(n6612), .A2(n8910), .ZN(n8911) );
  NAND2_X1 U9748 ( .A1(n12994), .A2(n12993), .ZN(n12995) );
  NAND2_X1 U9749 ( .A1(n13006), .A2(n13005), .ZN(n13007) );
  NAND2_X1 U9750 ( .A1(n8933), .A2(n8932), .ZN(n8934) );
  NAND2_X1 U9751 ( .A1(n13033), .A2(n13032), .ZN(n13034) );
  AND2_X1 U9752 ( .A1(n11611), .A2(n14240), .ZN(n8968) );
  AND2_X1 U9753 ( .A1(n8974), .A2(n14537), .ZN(n8975) );
  NAND2_X1 U9754 ( .A1(n9006), .A2(n9005), .ZN(n9012) );
  INV_X1 U9755 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n7611) );
  INV_X1 U9756 ( .A(n12550), .ZN(n12375) );
  INV_X1 U9757 ( .A(n10728), .ZN(n10724) );
  INV_X1 U9758 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n8279) );
  OR2_X1 U9759 ( .A1(n12566), .A2(n12363), .ZN(n11802) );
  INV_X1 U9760 ( .A(n11077), .ZN(n10863) );
  NAND2_X1 U9761 ( .A1(n10214), .A2(n6846), .ZN(n10432) );
  INV_X1 U9762 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n10765) );
  OR2_X1 U9763 ( .A1(n14027), .A2(n13929), .ZN(n13364) );
  AOI22_X1 U9764 ( .A1(n10246), .A2(n10245), .B1(n12120), .B2(n14125), .ZN(
        n10247) );
  NAND2_X1 U9765 ( .A1(n12015), .A2(n12016), .ZN(n12017) );
  INV_X1 U9766 ( .A(n8719), .ZN(n8299) );
  NAND2_X1 U9767 ( .A1(n8710), .A2(n8379), .ZN(n8383) );
  INV_X1 U9768 ( .A(n8477), .ZN(n8328) );
  INV_X1 U9769 ( .A(n15209), .ZN(n9177) );
  OR2_X1 U9770 ( .A1(n15185), .A2(n15182), .ZN(n9194) );
  INV_X1 U9771 ( .A(n10487), .ZN(n9171) );
  OR2_X1 U9772 ( .A1(n7972), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n7989) );
  NOR2_X1 U9773 ( .A1(n7932), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n7950) );
  AND2_X1 U9774 ( .A1(n8059), .A2(n9398), .ZN(n8071) );
  INV_X1 U9775 ( .A(n15353), .ZN(n12406) );
  INV_X1 U9776 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n7701) );
  NAND2_X1 U9777 ( .A1(n7926), .A2(n7925), .ZN(n7928) );
  NAND2_X1 U9778 ( .A1(n7844), .A2(n7843), .ZN(n7846) );
  INV_X1 U9779 ( .A(n12879), .ZN(n12739) );
  NAND2_X1 U9780 ( .A1(n12815), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n12834) );
  NAND2_X1 U9781 ( .A1(n12752), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n12771) );
  OR2_X1 U9782 ( .A1(n11743), .A2(n11742), .ZN(n11871) );
  AND2_X1 U9783 ( .A1(n13999), .A2(n13370), .ZN(n13371) );
  NAND2_X1 U9784 ( .A1(n10884), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n10993) );
  NAND2_X1 U9785 ( .A1(n10271), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n10410) );
  OR2_X1 U9786 ( .A1(n10135), .A2(n10199), .ZN(n9546) );
  OR2_X1 U9787 ( .A1(n11909), .A2(n11908), .ZN(n11910) );
  AND2_X1 U9788 ( .A1(n9126), .A2(n9131), .ZN(n9121) );
  INV_X1 U9789 ( .A(n8300), .ZN(n8718) );
  NAND2_X2 U9790 ( .A1(n12005), .A2(n14253), .ZN(n8405) );
  INV_X1 U9791 ( .A(n11109), .ZN(n8521) );
  INV_X1 U9792 ( .A(n11196), .ZN(n11396) );
  NAND2_X1 U9793 ( .A1(n8351), .A2(SI_15_), .ZN(n8600) );
  NOR2_X1 U9794 ( .A1(n9363), .A2(n9364), .ZN(n9309) );
  AND2_X1 U9795 ( .A1(n7872), .A2(n7871), .ZN(n7885) );
  NOR2_X1 U9796 ( .A1(n7736), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7786) );
  NOR2_X1 U9797 ( .A1(n11434), .A2(n11435), .ZN(n11451) );
  OR2_X1 U9798 ( .A1(n7918), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n7932) );
  AND2_X1 U9799 ( .A1(n7786), .A2(n7785), .ZN(n7795) );
  NAND2_X1 U9800 ( .A1(n7959), .A2(n12194), .ZN(n7972) );
  OR2_X1 U9801 ( .A1(n7820), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7836) );
  OR2_X1 U9802 ( .A1(n15203), .A2(n15351), .ZN(n12224) );
  AND2_X1 U9803 ( .A1(n8046), .A2(n12223), .ZN(n8059) );
  AOI21_X1 U9804 ( .B1(n12435), .B2(n12406), .A(n12405), .ZN(n12407) );
  INV_X1 U9805 ( .A(n12364), .ZN(n12574) );
  NAND2_X1 U9806 ( .A1(n7702), .A2(n7701), .ZN(n7721) );
  INV_X1 U9807 ( .A(n10428), .ZN(n15376) );
  AND2_X1 U9808 ( .A1(n10440), .A2(n10439), .ZN(n15359) );
  NAND2_X1 U9809 ( .A1(n7860), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7863) );
  AND2_X1 U9810 ( .A1(n7814), .A2(n7805), .ZN(n7806) );
  AND2_X1 U9811 ( .A1(n7691), .A2(n7678), .ZN(n7689) );
  AND2_X1 U9812 ( .A1(n11309), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n11362) );
  INV_X1 U9813 ( .A(n12780), .ZN(n12769) );
  NOR2_X1 U9814 ( .A1(n12744), .A2(n12943), .ZN(n12752) );
  INV_X1 U9815 ( .A(n12903), .ZN(n13168) );
  OR2_X1 U9816 ( .A1(n15019), .A2(n15018), .ZN(n15021) );
  INV_X1 U9817 ( .A(n13995), .ZN(n13819) );
  XNOR2_X1 U9818 ( .A(n13990), .B(n13373), .ZN(n13801) );
  INV_X1 U9819 ( .A(n13052), .ZN(n14824) );
  INV_X1 U9820 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n13635) );
  INV_X1 U9821 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n8512) );
  NAND2_X1 U9822 ( .A1(n11924), .A2(n11923), .ZN(n11925) );
  OR2_X1 U9823 ( .A1(n8677), .A2(n14180), .ZN(n8694) );
  NAND2_X1 U9824 ( .A1(n8637), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8665) );
  INV_X1 U9825 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n14845) );
  OR3_X1 U9826 ( .A1(n11032), .A2(n11031), .A3(n11030), .ZN(n11204) );
  INV_X1 U9827 ( .A(n14404), .ZN(n14210) );
  AND2_X1 U9828 ( .A1(n8899), .A2(n9089), .ZN(n10092) );
  INV_X1 U9829 ( .A(n14540), .ZN(n14466) );
  XNOR2_X1 U9830 ( .A(n8346), .B(n9560), .ZN(n8567) );
  INV_X1 U9831 ( .A(n12230), .ZN(n15213) );
  AND2_X1 U9832 ( .A1(n9253), .A2(n10540), .ZN(n15193) );
  AND4_X1 U9833 ( .A1(n8076), .A2(n8075), .A3(n8074), .A4(n8073), .ZN(n12402)
         );
  AND2_X1 U9834 ( .A1(n7965), .A2(n7964), .ZN(n12535) );
  AND4_X1 U9835 ( .A1(n7859), .A2(n7858), .A3(n7857), .A4(n7856), .ZN(n11709)
         );
  INV_X1 U9836 ( .A(n15320), .ZN(n15266) );
  INV_X1 U9837 ( .A(n15359), .ZN(n15369) );
  AND2_X1 U9838 ( .A1(n10456), .A2(n10455), .ZN(n10538) );
  NAND2_X1 U9839 ( .A1(n15373), .A2(n12595), .ZN(n14775) );
  INV_X1 U9840 ( .A(n10540), .ZN(n11265) );
  INV_X1 U9841 ( .A(n15374), .ZN(n14770) );
  AND2_X1 U9842 ( .A1(n9972), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9405) );
  NAND2_X1 U9843 ( .A1(n11362), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n11546) );
  OR2_X1 U9844 ( .A1(n12901), .A2(n13405), .ZN(n12852) );
  INV_X1 U9845 ( .A(n15026), .ZN(n15045) );
  INV_X1 U9846 ( .A(n13928), .ZN(n14787) );
  INV_X1 U9847 ( .A(n13925), .ZN(n15054) );
  INV_X1 U9848 ( .A(n13937), .ZN(n15068) );
  OR2_X1 U9849 ( .A1(n10164), .A2(n15085), .ZN(n13957) );
  OR2_X1 U9850 ( .A1(n9793), .A2(n13222), .ZN(n15150) );
  INV_X1 U9851 ( .A(n15147), .ZN(n15117) );
  INV_X1 U9852 ( .A(n9729), .ZN(n9531) );
  INV_X1 U9853 ( .A(n11401), .ZN(n9139) );
  INV_X1 U9854 ( .A(n14913), .ZN(n14298) );
  INV_X1 U9855 ( .A(n14386), .ZN(n14387) );
  AND2_X1 U9856 ( .A1(n10092), .A2(n14256), .ZN(n14539) );
  INV_X1 U9857 ( .A(n14705), .ZN(n14531) );
  INV_X1 U9858 ( .A(n14345), .ZN(n14558) );
  INV_X1 U9859 ( .A(n14963), .ZN(n14947) );
  NAND2_X1 U9860 ( .A1(n8849), .A2(n12121), .ZN(n14959) );
  NAND2_X1 U9861 ( .A1(n14546), .A2(n8851), .ZN(n14963) );
  INV_X1 U9862 ( .A(n14959), .ZN(n14965) );
  AND2_X1 U9863 ( .A1(n9984), .A2(n9983), .ZN(n15326) );
  AND2_X1 U9864 ( .A1(n9271), .A2(n9270), .ZN(n15215) );
  INV_X1 U9865 ( .A(n12552), .ZN(n12372) );
  INV_X1 U9866 ( .A(n15326), .ZN(n15308) );
  INV_X1 U9867 ( .A(n15264), .ZN(n15333) );
  NAND2_X1 U9868 ( .A1(n10546), .A2(n12555), .ZN(n15380) );
  INV_X1 U9869 ( .A(n15436), .ZN(n15433) );
  AND3_X2 U9870 ( .A1(n10461), .A2(n10538), .A3(n10460), .ZN(n15436) );
  INV_X1 U9871 ( .A(n15421), .ZN(n15419) );
  INV_X1 U9872 ( .A(SI_13_), .ZN(n9560) );
  INV_X1 U9873 ( .A(n10050), .ZN(n10115) );
  INV_X1 U9874 ( .A(n14796), .ZN(n11848) );
  INV_X1 U9875 ( .A(n14785), .ZN(n13264) );
  OR2_X1 U9876 ( .A1(n9641), .A2(P2_U3088), .ZN(n15035) );
  INV_X1 U9877 ( .A(n13944), .ZN(n15059) );
  AND2_X1 U9878 ( .A1(n13957), .A2(n10195), .ZN(n15072) );
  INV_X1 U9879 ( .A(n15177), .ZN(n15174) );
  INV_X1 U9880 ( .A(n15157), .ZN(n15156) );
  INV_X1 U9881 ( .A(n15078), .ZN(n15079) );
  INV_X1 U9882 ( .A(n15082), .ZN(n15085) );
  INV_X1 U9883 ( .A(n13214), .ZN(n13331) );
  INV_X1 U9884 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n13506) );
  OR2_X1 U9885 ( .A1(n10371), .A2(P1_U3086), .ZN(n14909) );
  INV_X1 U9886 ( .A(n14215), .ZN(n14896) );
  OR2_X1 U9887 ( .A1(n9814), .A2(n14256), .ZN(n14921) );
  OR2_X1 U9888 ( .A1(n14526), .A2(n14959), .ZN(n14511) );
  AND2_X1 U9889 ( .A1(n10226), .A2(n14498), .ZN(n14705) );
  INV_X1 U9890 ( .A(n14982), .ZN(n14980) );
  OR2_X1 U9891 ( .A1(n14614), .A2(n14613), .ZN(n14655) );
  AND3_X1 U9892 ( .A1(n14867), .A2(n14866), .A3(n14865), .ZN(n14871) );
  AND2_X1 U9893 ( .A1(n10366), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9591) );
  OR2_X1 U9894 ( .A1(n8574), .A2(n8659), .ZN(n11205) );
  INV_X1 U9895 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9593) );
  XNOR2_X1 U9896 ( .A(n9388), .B(n9387), .ZN(n9389) );
  INV_X1 U9897 ( .A(n14252), .ZN(P1_U4016) );
  NAND2_X1 U9898 ( .A1(n8897), .A2(n8896), .ZN(P1_U3524) );
  NAND4_X1 U9899 ( .A1(n7607), .A2(n7847), .A3(n13648), .A4(n13643), .ZN(n7608) );
  NAND3_X1 U9900 ( .A1(n13642), .A2(n7894), .A3(n7611), .ZN(n7612) );
  INV_X1 U9901 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7615) );
  INV_X1 U9902 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7614) );
  NOR2_X2 U9903 ( .A1(n7635), .A2(P3_IR_REG_27__SCAN_IN), .ZN(n7631) );
  INV_X1 U9904 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n7616) );
  AND2_X2 U9905 ( .A1(n7631), .A2(n7616), .ZN(n7619) );
  INV_X1 U9906 ( .A(n7619), .ZN(n7633) );
  NAND2_X1 U9907 ( .A1(n7633), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7617) );
  INV_X1 U9909 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7618) );
  NAND2_X1 U9910 ( .A1(n7619), .A2(n7618), .ZN(n7621) );
  NAND2_X2 U9911 ( .A1(n7620), .A2(n7621), .ZN(n7624) );
  XNOR2_X2 U9912 ( .A(n7622), .B(P3_IR_REG_30__SCAN_IN), .ZN(n7625) );
  NAND2_X1 U9913 ( .A1(n8085), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n7629) );
  INV_X1 U9914 ( .A(n7625), .ZN(n12726) );
  NAND2_X1 U9915 ( .A1(n7666), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n7628) );
  AND2_X2 U9916 ( .A1(n7625), .A2(n7624), .ZN(n7667) );
  NAND2_X1 U9917 ( .A1(n7667), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7627) );
  NAND2_X1 U9918 ( .A1(n7595), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7626) );
  OR2_X1 U9919 ( .A1(n7631), .A2(n8267), .ZN(n7632) );
  NAND2_X1 U9920 ( .A1(n7635), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7637) );
  INV_X1 U9921 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7636) );
  NAND3_X1 U9922 ( .A1(n7640), .A2(n7639), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n7643) );
  NAND2_X1 U9923 ( .A1(n8305), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7644) );
  NAND2_X1 U9924 ( .A1(n9490), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7646) );
  XNOR2_X1 U9925 ( .A(n7676), .B(n7675), .ZN(n9521) );
  OR2_X1 U9926 ( .A1(n7672), .A2(SI_2_), .ZN(n7647) );
  OAI211_X1 U9927 ( .C1(n10050), .C2(n9973), .A(n7648), .B(n7647), .ZN(n15360)
         );
  NAND2_X1 U9928 ( .A1(n7667), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n7652) );
  NAND2_X1 U9929 ( .A1(n8085), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n7651) );
  NAND2_X1 U9930 ( .A1(n7595), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7650) );
  INV_X1 U9931 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7655) );
  INV_X1 U9932 ( .A(SI_1_), .ZN(n9512) );
  OR2_X1 U9933 ( .A1(n7672), .A2(n9512), .ZN(n7658) );
  XNOR2_X1 U9934 ( .A(n7656), .B(n7664), .ZN(n9513) );
  OR2_X1 U9935 ( .A1(n7674), .A2(n9513), .ZN(n7657) );
  OAI211_X1 U9936 ( .C1(n9973), .C2(n10162), .A(n7658), .B(n7657), .ZN(n9160)
         );
  NAND2_X1 U9937 ( .A1(n8085), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n7662) );
  NAND2_X1 U9938 ( .A1(n7666), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n7661) );
  NAND2_X1 U9939 ( .A1(n7667), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7660) );
  NAND2_X1 U9940 ( .A1(n7595), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n7659) );
  NAND4_X1 U9941 ( .A1(n7662), .A2(n7661), .A3(n7660), .A4(n7659), .ZN(n15367)
         );
  INV_X1 U9942 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10035) );
  INV_X1 U9943 ( .A(SI_0_), .ZN(n9524) );
  INV_X1 U9944 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8406) );
  NAND2_X1 U9945 ( .A1(n8406), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7663) );
  AND2_X1 U9946 ( .A1(n7664), .A2(n7663), .ZN(n9525) );
  NOR2_X2 U9947 ( .A1(n15367), .A2(n11950), .ZN(n8135) );
  NAND2_X1 U9948 ( .A1(n15354), .A2(n9160), .ZN(n9157) );
  INV_X1 U9949 ( .A(n15365), .ZN(n10435) );
  NAND2_X1 U9950 ( .A1(n10435), .A2(n7649), .ZN(n8156) );
  NAND2_X1 U9951 ( .A1(n15348), .A2(n8156), .ZN(n15335) );
  INV_X1 U9952 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n7665) );
  NAND2_X1 U9953 ( .A1(n7991), .A2(n7665), .ZN(n7671) );
  NAND2_X1 U9954 ( .A1(n7666), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n7670) );
  NAND2_X1 U9955 ( .A1(n7667), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7669) );
  NAND2_X1 U9956 ( .A1(n7684), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7668) );
  AND4_X2 U9957 ( .A1(n7671), .A2(n7670), .A3(n7669), .A4(n7668), .ZN(n15352)
         );
  OR2_X1 U9958 ( .A1(n7672), .A2(SI_3_), .ZN(n7682) );
  NAND2_X1 U9959 ( .A1(n9488), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7678) );
  XNOR2_X1 U9960 ( .A(n7690), .B(n7689), .ZN(n9518) );
  OR2_X1 U9961 ( .A1(n7674), .A2(n9518), .ZN(n7681) );
  OR2_X1 U9962 ( .A1(n7694), .A2(n8267), .ZN(n7679) );
  XNOR2_X1 U9963 ( .A(n7679), .B(n7693), .ZN(n10056) );
  NAND2_X1 U9964 ( .A1(n7946), .A2(n10056), .ZN(n7680) );
  NAND2_X1 U9965 ( .A1(n15352), .A2(n15200), .ZN(n8161) );
  INV_X1 U9966 ( .A(n15200), .ZN(n15343) );
  NAND2_X1 U9967 ( .A1(n15335), .A2(n15336), .ZN(n7683) );
  NAND2_X1 U9968 ( .A1(n7683), .A2(n8161), .ZN(n10430) );
  NAND2_X1 U9969 ( .A1(n7684), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7688) );
  NAND2_X1 U9970 ( .A1(n7870), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n7687) );
  XNOR2_X1 U9971 ( .A(P3_REG3_REG_4__SCAN_IN), .B(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n10547) );
  NAND2_X1 U9972 ( .A1(n8085), .A2(n10547), .ZN(n7686) );
  NAND2_X1 U9973 ( .A1(n8103), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7685) );
  AND4_X2 U9974 ( .A1(n7688), .A2(n7687), .A3(n7686), .A4(n7685), .ZN(n10565)
         );
  OR2_X1 U9975 ( .A1(n7673), .A2(SI_4_), .ZN(n7699) );
  NAND2_X1 U9976 ( .A1(n9502), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n7692) );
  XNOR2_X1 U9977 ( .A(n7709), .B(n7708), .ZN(n9477) );
  OR2_X1 U9978 ( .A1(n7674), .A2(n9477), .ZN(n7698) );
  NAND2_X1 U9979 ( .A1(n7694), .A2(n7693), .ZN(n7713) );
  NAND2_X1 U9980 ( .A1(n7713), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7695) );
  NAND2_X1 U9981 ( .A1(n7946), .A2(n10062), .ZN(n7697) );
  NAND2_X1 U9982 ( .A1(n10565), .A2(n11274), .ZN(n8165) );
  INV_X1 U9983 ( .A(n11274), .ZN(n10490) );
  NAND2_X1 U9984 ( .A1(n15192), .A2(n10490), .ZN(n8162) );
  NAND2_X1 U9985 ( .A1(n8165), .A2(n8162), .ZN(n10442) );
  NAND2_X1 U9986 ( .A1(n10429), .A2(n8165), .ZN(n10722) );
  NAND2_X1 U9987 ( .A1(n7684), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7707) );
  NAND2_X1 U9988 ( .A1(n7870), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n7706) );
  OR2_X1 U9989 ( .A1(n7702), .A2(n7701), .ZN(n7703) );
  NAND2_X1 U9990 ( .A1(n7721), .A2(n7703), .ZN(n10801) );
  NAND2_X1 U9991 ( .A1(n7991), .A2(n10801), .ZN(n7705) );
  NAND2_X1 U9992 ( .A1(n8103), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7704) );
  NAND4_X1 U9993 ( .A1(n7707), .A2(n7706), .A3(n7705), .A4(n7704), .ZN(n12242)
         );
  OR2_X1 U9994 ( .A1(n7673), .A2(SI_5_), .ZN(n7720) );
  NAND2_X1 U9995 ( .A1(n9503), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7712) );
  XNOR2_X1 U9996 ( .A(n7730), .B(n7729), .ZN(n9480) );
  OR2_X1 U9997 ( .A1(n7674), .A2(n9480), .ZN(n7719) );
  NAND2_X1 U9998 ( .A1(n7715), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7714) );
  MUX2_X1 U9999 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7714), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n7717) );
  INV_X1 U10000 ( .A(n7751), .ZN(n7716) );
  NAND2_X1 U10001 ( .A1(n7717), .A2(n7716), .ZN(n10064) );
  NAND2_X1 U10002 ( .A1(n7946), .A2(n10064), .ZN(n7718) );
  XNOR2_X1 U10003 ( .A(n12242), .B(n10802), .ZN(n10728) );
  INV_X1 U10004 ( .A(n12242), .ZN(n10860) );
  NAND2_X1 U10005 ( .A1(n10860), .A2(n10802), .ZN(n8163) );
  NAND2_X1 U10006 ( .A1(n7595), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n7727) );
  NAND2_X1 U10007 ( .A1(n8045), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n7726) );
  NAND2_X1 U10008 ( .A1(n7721), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7722) );
  AND2_X1 U10009 ( .A1(n7736), .A2(n7722), .ZN(n15216) );
  INV_X1 U10010 ( .A(n15216), .ZN(n7723) );
  NAND2_X1 U10011 ( .A1(n7991), .A2(n7723), .ZN(n7725) );
  NAND2_X1 U10012 ( .A1(n8103), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7724) );
  OR2_X1 U10013 ( .A1(n7751), .A2(n8267), .ZN(n7728) );
  XNOR2_X1 U10014 ( .A(n7728), .B(P3_IR_REG_6__SCAN_IN), .ZN(n10667) );
  XNOR2_X1 U10015 ( .A(n9515), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n7733) );
  XNOR2_X1 U10016 ( .A(n7743), .B(n7733), .ZN(n9527) );
  OR2_X1 U10017 ( .A1(n7674), .A2(n9527), .ZN(n7735) );
  INV_X1 U10018 ( .A(SI_6_), .ZN(n9526) );
  OR2_X1 U10019 ( .A1(n7673), .A2(n9526), .ZN(n7734) );
  OAI211_X1 U10020 ( .C1(n9973), .C2(n10651), .A(n7735), .B(n7734), .ZN(n15212) );
  NAND2_X1 U10021 ( .A1(n10858), .A2(n15212), .ZN(n8168) );
  INV_X1 U10022 ( .A(n15212), .ZN(n9176) );
  NAND2_X1 U10023 ( .A1(n12241), .A2(n9176), .ZN(n8172) );
  NAND2_X1 U10024 ( .A1(n7595), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n7741) );
  NAND2_X1 U10025 ( .A1(n7870), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n7740) );
  AND2_X1 U10026 ( .A1(n7736), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7737) );
  OR2_X1 U10027 ( .A1(n7737), .A2(n7786), .ZN(n10870) );
  NAND2_X1 U10028 ( .A1(n8085), .A2(n10870), .ZN(n7739) );
  NAND2_X1 U10029 ( .A1(n8103), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7738) );
  NAND2_X1 U10030 ( .A1(n9517), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7742) );
  NAND2_X1 U10031 ( .A1(n9515), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n7744) );
  NAND2_X1 U10032 ( .A1(n9530), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7765) );
  NAND2_X1 U10033 ( .A1(n9534), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n7746) );
  NAND2_X1 U10034 ( .A1(n7765), .A2(n7746), .ZN(n7747) );
  NAND2_X1 U10035 ( .A1(n7748), .A2(n7747), .ZN(n7749) );
  AND2_X1 U10036 ( .A1(n7766), .A2(n7749), .ZN(n9483) );
  OR2_X1 U10037 ( .A1(n7674), .A2(n9483), .ZN(n7756) );
  OR2_X1 U10038 ( .A1(n7673), .A2(SI_7_), .ZN(n7755) );
  NAND2_X1 U10039 ( .A1(n7751), .A2(n7750), .ZN(n7763) );
  NAND2_X1 U10040 ( .A1(n7763), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7753) );
  INV_X1 U10041 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n7752) );
  XNOR2_X1 U10042 ( .A(n7753), .B(n7752), .ZN(n15279) );
  NAND2_X1 U10043 ( .A1(n7946), .A2(n15279), .ZN(n7754) );
  NAND2_X1 U10044 ( .A1(n11094), .A2(n11089), .ZN(n8173) );
  INV_X1 U10045 ( .A(n11089), .ZN(n7757) );
  NAND2_X1 U10046 ( .A1(n12240), .A2(n7757), .ZN(n8174) );
  NAND2_X1 U10047 ( .A1(n8173), .A2(n8174), .ZN(n10865) );
  INV_X1 U10048 ( .A(n10865), .ZN(n8171) );
  NAND2_X1 U10049 ( .A1(n7758), .A2(n8173), .ZN(n11088) );
  NAND2_X1 U10050 ( .A1(n7684), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7762) );
  NAND2_X1 U10051 ( .A1(n7870), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n7761) );
  INV_X1 U10052 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n13719) );
  XNOR2_X1 U10053 ( .A(n7786), .B(n13719), .ZN(n11101) );
  NAND2_X1 U10054 ( .A1(n7991), .A2(n11101), .ZN(n7760) );
  NAND2_X1 U10055 ( .A1(n8103), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7759) );
  OAI21_X1 U10056 ( .B1(n7763), .B2(P3_IR_REG_7__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7764) );
  XNOR2_X1 U10057 ( .A(n7764), .B(P3_IR_REG_8__SCAN_IN), .ZN(n10650) );
  NAND2_X1 U10058 ( .A1(n9558), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7780) );
  NAND2_X1 U10059 ( .A1(n9556), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n7767) );
  OR2_X1 U10060 ( .A1(n7769), .A2(n7768), .ZN(n7770) );
  NAND2_X1 U10061 ( .A1(n7781), .A2(n7770), .ZN(n9473) );
  OR2_X1 U10062 ( .A1(n7674), .A2(n9473), .ZN(n7772) );
  INV_X1 U10063 ( .A(SI_8_), .ZN(n9474) );
  OR2_X1 U10064 ( .A1(n7673), .A2(n9474), .ZN(n7771) );
  OAI211_X1 U10065 ( .C1(n9973), .C2(n15296), .A(n7772), .B(n7771), .ZN(n11100) );
  NAND2_X1 U10066 ( .A1(n11250), .A2(n11100), .ZN(n8178) );
  INV_X1 U10067 ( .A(n11250), .ZN(n12239) );
  INV_X1 U10068 ( .A(n11100), .ZN(n11245) );
  NAND2_X1 U10069 ( .A1(n12239), .A2(n11245), .ZN(n8177) );
  NAND2_X1 U10070 ( .A1(n8178), .A2(n8177), .ZN(n11092) );
  INV_X1 U10071 ( .A(n11092), .ZN(n8176) );
  NAND2_X1 U10072 ( .A1(n11088), .A2(n8176), .ZN(n7773) );
  NAND2_X1 U10073 ( .A1(n7773), .A2(n8178), .ZN(n11244) );
  NOR2_X1 U10074 ( .A1(n7774), .A2(n8267), .ZN(n7775) );
  MUX2_X1 U10075 ( .A(n8267), .B(n7775), .S(P3_IR_REG_9__SCAN_IN), .Z(n7776)
         );
  INV_X1 U10076 ( .A(n7776), .ZN(n7778) );
  NAND2_X1 U10077 ( .A1(n7778), .A2(n7777), .ZN(n15321) );
  INV_X1 U10078 ( .A(n15321), .ZN(n10676) );
  OAI22_X1 U10079 ( .A1(n7673), .A2(SI_9_), .B1(n10676), .B2(n9973), .ZN(n7779) );
  INV_X1 U10080 ( .A(n7779), .ZN(n7784) );
  NAND2_X1 U10081 ( .A1(n9593), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n7803) );
  NAND2_X1 U10082 ( .A1(n10877), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n7782) );
  XNOR2_X1 U10083 ( .A(n7802), .B(n7801), .ZN(n9529) );
  NAND2_X1 U10084 ( .A1(n9529), .A2(n8099), .ZN(n7783) );
  NAND2_X1 U10085 ( .A1(n7784), .A2(n7783), .ZN(n11287) );
  NAND2_X1 U10086 ( .A1(n7870), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n7791) );
  NAND2_X1 U10087 ( .A1(n8103), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7790) );
  NOR2_X1 U10088 ( .A1(P3_REG3_REG_9__SCAN_IN), .A2(P3_REG3_REG_8__SCAN_IN), 
        .ZN(n7785) );
  INV_X1 U10089 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n15313) );
  AOI21_X1 U10090 ( .B1(n7786), .B2(n13719), .A(n15313), .ZN(n7787) );
  OR2_X1 U10091 ( .A1(n7795), .A2(n7787), .ZN(n11289) );
  NAND2_X1 U10092 ( .A1(n7991), .A2(n11289), .ZN(n7789) );
  NAND2_X1 U10093 ( .A1(n7595), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n7788) );
  NAND4_X1 U10094 ( .A1(n7791), .A2(n7790), .A3(n7789), .A4(n7788), .ZN(n11329) );
  NAND2_X1 U10095 ( .A1(n11244), .A2(n11325), .ZN(n7792) );
  OR2_X1 U10096 ( .A1(n7795), .A2(n7794), .ZN(n7796) );
  AND2_X1 U10097 ( .A1(n7820), .A2(n7796), .ZN(n15191) );
  INV_X1 U10098 ( .A(n15191), .ZN(n11333) );
  NAND2_X1 U10099 ( .A1(n7991), .A2(n11333), .ZN(n7800) );
  NAND2_X1 U10100 ( .A1(n7870), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n7799) );
  NAND2_X1 U10101 ( .A1(n8103), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7798) );
  NAND2_X1 U10102 ( .A1(n8102), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7797) );
  NAND2_X1 U10103 ( .A1(n9733), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n7814) );
  NAND2_X1 U10104 ( .A1(n13506), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n7805) );
  OR2_X1 U10105 ( .A1(n7807), .A2(n7806), .ZN(n7808) );
  NAND2_X1 U10106 ( .A1(n7815), .A2(n7808), .ZN(n9498) );
  NAND2_X1 U10107 ( .A1(n7777), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7809) );
  MUX2_X1 U10108 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7809), .S(
        P3_IR_REG_10__SCAN_IN), .Z(n7810) );
  OR2_X1 U10109 ( .A1(n7777), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n7832) );
  AND2_X1 U10110 ( .A1(n7810), .A2(n7832), .ZN(n10678) );
  OAI22_X1 U10111 ( .A1(n7673), .A2(SI_10_), .B1(n10678), .B2(n9973), .ZN(
        n7811) );
  NAND2_X1 U10112 ( .A1(n11442), .A2(n15189), .ZN(n8187) );
  INV_X1 U10113 ( .A(n15189), .ZN(n7812) );
  NAND2_X1 U10114 ( .A1(n11342), .A2(n7812), .ZN(n11350) );
  NAND2_X1 U10115 ( .A1(n8187), .A2(n11350), .ZN(n11336) );
  INV_X1 U10116 ( .A(n11336), .ZN(n7813) );
  XNOR2_X1 U10117 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n7816) );
  XNOR2_X1 U10118 ( .A(n7829), .B(n7816), .ZN(n9510) );
  NAND2_X1 U10119 ( .A1(n9510), .A2(n8099), .ZN(n7819) );
  INV_X1 U10120 ( .A(SI_11_), .ZN(n9511) );
  NAND2_X1 U10121 ( .A1(n7832), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7817) );
  XNOR2_X1 U10122 ( .A(n7817), .B(n13648), .ZN(n11065) );
  AOI22_X1 U10123 ( .A1(n6993), .A2(n9511), .B1(n7946), .B2(n11065), .ZN(n7818) );
  NAND2_X1 U10124 ( .A1(n7819), .A2(n7818), .ZN(n11522) );
  NAND2_X1 U10125 ( .A1(n7870), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n7825) );
  NAND2_X1 U10126 ( .A1(n8103), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n7824) );
  NAND2_X1 U10127 ( .A1(n7820), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7821) );
  NAND2_X1 U10128 ( .A1(n7836), .A2(n7821), .ZN(n11444) );
  NAND2_X1 U10129 ( .A1(n7991), .A2(n11444), .ZN(n7823) );
  NAND2_X1 U10130 ( .A1(n8102), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n7822) );
  INV_X1 U10131 ( .A(n11526), .ZN(n12238) );
  OR2_X1 U10132 ( .A1(n11522), .A2(n12238), .ZN(n8186) );
  NAND2_X1 U10133 ( .A1(n11522), .A2(n12238), .ZN(n8188) );
  NAND2_X1 U10134 ( .A1(n8186), .A2(n8188), .ZN(n11351) );
  INV_X1 U10135 ( .A(n11350), .ZN(n7826) );
  NOR2_X1 U10136 ( .A1(n11351), .A2(n7826), .ZN(n7827) );
  INV_X1 U10137 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9758) );
  NAND2_X1 U10138 ( .A1(n9758), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n7828) );
  INV_X1 U10139 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9819) );
  NAND2_X1 U10140 ( .A1(n9819), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n7830) );
  XNOR2_X1 U10141 ( .A(n9727), .B(P1_DATAO_REG_12__SCAN_IN), .ZN(n7842) );
  XNOR2_X1 U10142 ( .A(n7844), .B(n7842), .ZN(n9551) );
  NAND2_X1 U10143 ( .A1(n9551), .A2(n8099), .ZN(n7835) );
  NOR2_X1 U10144 ( .A1(n7832), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n7848) );
  OR2_X1 U10145 ( .A1(n7848), .A2(n8267), .ZN(n7833) );
  XNOR2_X1 U10146 ( .A(n7833), .B(P3_IR_REG_12__SCAN_IN), .ZN(n11476) );
  AOI22_X1 U10147 ( .A1(n6993), .A2(SI_12_), .B1(n7946), .B2(n11476), .ZN(
        n7834) );
  NAND2_X1 U10148 ( .A1(n7835), .A2(n7834), .ZN(n11570) );
  NAND2_X1 U10149 ( .A1(n8102), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n7841) );
  NAND2_X1 U10150 ( .A1(n8045), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n7840) );
  NAND2_X1 U10151 ( .A1(n7836), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7837) );
  NAND2_X1 U10152 ( .A1(n7854), .A2(n7837), .ZN(n11528) );
  NAND2_X1 U10153 ( .A1(n8085), .A2(n11528), .ZN(n7839) );
  NAND2_X1 U10154 ( .A1(n8103), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7838) );
  OR2_X1 U10155 ( .A1(n11570), .A2(n11574), .ZN(n8191) );
  NAND2_X1 U10156 ( .A1(n11570), .A2(n11574), .ZN(n8192) );
  NAND2_X1 U10157 ( .A1(n8191), .A2(n8192), .ZN(n11568) );
  INV_X1 U10158 ( .A(n7842), .ZN(n7843) );
  NAND2_X1 U10159 ( .A1(n9727), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n7845) );
  XNOR2_X1 U10160 ( .A(n7860), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n9559) );
  NAND2_X1 U10161 ( .A1(n9559), .A2(n8099), .ZN(n7853) );
  NAND2_X1 U10162 ( .A1(n7848), .A2(n7847), .ZN(n7850) );
  NAND2_X1 U10163 ( .A1(n7850), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7849) );
  MUX2_X1 U10164 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7849), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n7851) );
  OR2_X1 U10165 ( .A1(n7850), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n7864) );
  NAND2_X1 U10166 ( .A1(n7851), .A2(n7864), .ZN(n12260) );
  AOI22_X1 U10167 ( .A1(n6993), .A2(n9560), .B1(n7946), .B2(n12260), .ZN(n7852) );
  NAND2_X1 U10168 ( .A1(n8102), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n7859) );
  NAND2_X1 U10169 ( .A1(n8045), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n7858) );
  AND2_X1 U10170 ( .A1(n7854), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n7855) );
  OR2_X1 U10171 ( .A1(n7855), .A2(n7872), .ZN(n11577) );
  NAND2_X1 U10172 ( .A1(n7991), .A2(n11577), .ZN(n7857) );
  NAND2_X1 U10173 ( .A1(n8103), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n7856) );
  NOR2_X1 U10174 ( .A1(n11798), .A2(n12236), .ZN(n8196) );
  INV_X1 U10175 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n13698) );
  NAND2_X1 U10176 ( .A1(n7861), .A2(n13698), .ZN(n7862) );
  XNOR2_X1 U10177 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n7878) );
  XNOR2_X1 U10178 ( .A(n7879), .B(n7878), .ZN(n9660) );
  NAND2_X1 U10179 ( .A1(n9660), .A2(n8099), .ZN(n7869) );
  INV_X1 U10180 ( .A(SI_14_), .ZN(n9661) );
  NAND2_X1 U10181 ( .A1(n7864), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7865) );
  MUX2_X1 U10182 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7865), .S(
        P3_IR_REG_14__SCAN_IN), .Z(n7867) );
  INV_X1 U10183 ( .A(n7866), .ZN(n7881) );
  NAND2_X1 U10184 ( .A1(n7867), .A2(n7881), .ZN(n12282) );
  AOI22_X1 U10185 ( .A1(n6993), .A2(n9661), .B1(n7946), .B2(n12282), .ZN(n7868) );
  NAND2_X1 U10186 ( .A1(n8102), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n7877) );
  NAND2_X1 U10187 ( .A1(n7870), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n7876) );
  INV_X1 U10188 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n7871) );
  NOR2_X1 U10189 ( .A1(n7872), .A2(n7871), .ZN(n7873) );
  OR2_X1 U10190 ( .A1(n7885), .A2(n7873), .ZN(n11771) );
  NAND2_X1 U10191 ( .A1(n7991), .A2(n11771), .ZN(n7875) );
  NAND2_X1 U10192 ( .A1(n8103), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n7874) );
  NAND4_X1 U10193 ( .A1(n7877), .A2(n7876), .A3(n7875), .A4(n7874), .ZN(n12235) );
  NAND2_X1 U10194 ( .A1(n12711), .A2(n12235), .ZN(n8202) );
  NAND2_X1 U10195 ( .A1(n11768), .A2(n8200), .ZN(n11720) );
  INV_X1 U10196 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10207) );
  NAND2_X1 U10197 ( .A1(n10207), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n7880) );
  INV_X1 U10198 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10348) );
  XNOR2_X1 U10199 ( .A(n10348), .B(P1_DATAO_REG_15__SCAN_IN), .ZN(n7891) );
  XNOR2_X1 U10200 ( .A(n7893), .B(n7891), .ZN(n9725) );
  NAND2_X1 U10201 ( .A1(n9725), .A2(n8099), .ZN(n7884) );
  NAND2_X1 U10202 ( .A1(n7881), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7882) );
  XNOR2_X1 U10203 ( .A(n7882), .B(P3_IR_REG_15__SCAN_IN), .ZN(n12303) );
  AOI22_X1 U10204 ( .A1(n6993), .A2(SI_15_), .B1(n7946), .B2(n12303), .ZN(
        n7883) );
  NAND2_X1 U10205 ( .A1(n8102), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n7890) );
  NAND2_X1 U10206 ( .A1(n8045), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n7889) );
  INV_X1 U10207 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n12279) );
  NOR2_X1 U10208 ( .A1(n7885), .A2(n12279), .ZN(n7886) );
  OR2_X1 U10209 ( .A1(n7900), .A2(n7886), .ZN(n11734) );
  NAND2_X1 U10210 ( .A1(n7991), .A2(n11734), .ZN(n7888) );
  NAND2_X1 U10211 ( .A1(n8103), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7887) );
  NAND2_X1 U10212 ( .A1(n11799), .A2(n11727), .ZN(n8203) );
  NAND2_X1 U10213 ( .A1(n8201), .A2(n8203), .ZN(n11710) );
  NAND2_X1 U10214 ( .A1(n11720), .A2(n11712), .ZN(n11719) );
  NAND2_X1 U10215 ( .A1(n11719), .A2(n8203), .ZN(n11807) );
  INV_X1 U10216 ( .A(n7891), .ZN(n7892) );
  XNOR2_X1 U10217 ( .A(n8356), .B(P1_DATAO_REG_16__SCAN_IN), .ZN(n7907) );
  XNOR2_X1 U10218 ( .A(n7909), .B(n7907), .ZN(n9807) );
  NAND2_X1 U10219 ( .A1(n9807), .A2(n8099), .ZN(n7899) );
  NAND2_X1 U10220 ( .A1(n7866), .A2(n7894), .ZN(n7896) );
  NAND2_X1 U10221 ( .A1(n7896), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7895) );
  MUX2_X1 U10222 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7895), .S(
        P3_IR_REG_16__SCAN_IN), .Z(n7897) );
  INV_X1 U10223 ( .A(n8121), .ZN(n7912) );
  AND2_X1 U10224 ( .A1(n7897), .A2(n7912), .ZN(n12307) );
  AOI22_X1 U10225 ( .A1(n6993), .A2(SI_16_), .B1(n7946), .B2(n12307), .ZN(
        n7898) );
  NAND2_X1 U10226 ( .A1(n8102), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n7905) );
  NAND2_X1 U10227 ( .A1(n8045), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n7904) );
  INV_X1 U10228 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n11857) );
  OR2_X1 U10229 ( .A1(n7900), .A2(n11857), .ZN(n7901) );
  NAND2_X1 U10230 ( .A1(n7918), .A2(n7901), .ZN(n11861) );
  NAND2_X1 U10231 ( .A1(n7991), .A2(n11861), .ZN(n7903) );
  NAND2_X1 U10232 ( .A1(n8103), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n7902) );
  NAND4_X1 U10233 ( .A1(n7905), .A2(n7904), .A3(n7903), .A4(n7902), .ZN(n12570) );
  INV_X1 U10234 ( .A(n12570), .ZN(n7906) );
  OR2_X1 U10235 ( .A1(n12365), .A2(n7906), .ZN(n8206) );
  NAND2_X1 U10236 ( .A1(n12365), .A2(n7906), .ZN(n8204) );
  NAND2_X1 U10237 ( .A1(n11807), .A2(n11806), .ZN(n11805) );
  NAND2_X1 U10238 ( .A1(n11805), .A2(n8204), .ZN(n12575) );
  INV_X1 U10239 ( .A(n7907), .ZN(n7908) );
  NAND2_X1 U10240 ( .A1(n8356), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n7910) );
  XNOR2_X1 U10241 ( .A(n8362), .B(P1_DATAO_REG_17__SCAN_IN), .ZN(n7924) );
  XNOR2_X1 U10242 ( .A(n7926), .B(n7924), .ZN(n9885) );
  NAND2_X1 U10243 ( .A1(n9885), .A2(n8099), .ZN(n7917) );
  NAND2_X1 U10244 ( .A1(n7912), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7913) );
  MUX2_X1 U10245 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7913), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n7915) );
  NAND2_X1 U10246 ( .A1(n7915), .A2(n7943), .ZN(n12320) );
  INV_X1 U10247 ( .A(n12320), .ZN(n14753) );
  AOI22_X1 U10248 ( .A1(n6993), .A2(SI_17_), .B1(n7946), .B2(n14753), .ZN(
        n7916) );
  NAND2_X1 U10249 ( .A1(n7918), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n7919) );
  NAND2_X1 U10250 ( .A1(n7932), .A2(n7919), .ZN(n12576) );
  NAND2_X1 U10251 ( .A1(n12576), .A2(n7991), .ZN(n7923) );
  NAND2_X1 U10252 ( .A1(n8045), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n7922) );
  NAND2_X1 U10253 ( .A1(n8103), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7921) );
  NAND2_X1 U10254 ( .A1(n8102), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n7920) );
  OR2_X1 U10255 ( .A1(n12636), .A2(n12552), .ZN(n8208) );
  NAND2_X1 U10256 ( .A1(n12636), .A2(n12552), .ZN(n12543) );
  NAND2_X1 U10257 ( .A1(n8208), .A2(n12543), .ZN(n12364) );
  NAND2_X1 U10258 ( .A1(n12575), .A2(n12574), .ZN(n12573) );
  INV_X1 U10259 ( .A(n7924), .ZN(n7925) );
  NAND2_X1 U10260 ( .A1(n8362), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n7927) );
  INV_X1 U10261 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10613) );
  XNOR2_X1 U10262 ( .A(n10613), .B(P1_DATAO_REG_18__SCAN_IN), .ZN(n7939) );
  XNOR2_X1 U10263 ( .A(n7941), .B(n7939), .ZN(n10000) );
  NAND2_X1 U10264 ( .A1(n10000), .A2(n8099), .ZN(n7931) );
  NAND2_X1 U10265 ( .A1(n7943), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7929) );
  XNOR2_X1 U10266 ( .A(n7929), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12344) );
  AOI22_X1 U10267 ( .A1(n6993), .A2(SI_18_), .B1(n7946), .B2(n12344), .ZN(
        n7930) );
  INV_X1 U10268 ( .A(n7950), .ZN(n7934) );
  NAND2_X1 U10269 ( .A1(n7932), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n7933) );
  NAND2_X1 U10270 ( .A1(n7934), .A2(n7933), .ZN(n12554) );
  NAND2_X1 U10271 ( .A1(n12554), .A2(n7991), .ZN(n7937) );
  AOI22_X1 U10272 ( .A1(n8045), .A2(P3_REG0_REG_18__SCAN_IN), .B1(n8103), .B2(
        P3_REG2_REG_18__SCAN_IN), .ZN(n7936) );
  NAND2_X1 U10273 ( .A1(n8102), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n7935) );
  NAND2_X1 U10274 ( .A1(n12560), .A2(n12534), .ZN(n8213) );
  INV_X1 U10275 ( .A(n12543), .ZN(n8211) );
  NOR2_X1 U10276 ( .A1(n12375), .A2(n8211), .ZN(n7938) );
  NAND2_X1 U10277 ( .A1(n12573), .A2(n7938), .ZN(n12545) );
  INV_X1 U10278 ( .A(n7939), .ZN(n7940) );
  NAND2_X1 U10279 ( .A1(n10613), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n7942) );
  XNOR2_X1 U10280 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .ZN(n7955) );
  XNOR2_X1 U10281 ( .A(n7956), .B(n7955), .ZN(n11996) );
  NAND2_X1 U10282 ( .A1(n11996), .A2(n8099), .ZN(n7948) );
  INV_X1 U10283 ( .A(SI_19_), .ZN(n11994) );
  NOR2_X2 U10284 ( .A1(n7943), .A2(P3_IR_REG_18__SCAN_IN), .ZN(n8115) );
  INV_X1 U10285 ( .A(n8115), .ZN(n7944) );
  INV_X1 U10286 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8114) );
  AOI22_X1 U10287 ( .A1(n6993), .A2(n11994), .B1(n7946), .B2(n6687), .ZN(n7947) );
  INV_X1 U10288 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n7949) );
  NOR2_X1 U10289 ( .A1(n7950), .A2(n7949), .ZN(n7951) );
  OR2_X1 U10290 ( .A1(n7959), .A2(n7951), .ZN(n12538) );
  NAND2_X1 U10291 ( .A1(n12538), .A2(n7991), .ZN(n7954) );
  AOI22_X1 U10292 ( .A1(n8045), .A2(P3_REG0_REG_19__SCAN_IN), .B1(n8102), .B2(
        P3_REG1_REG_19__SCAN_IN), .ZN(n7953) );
  NAND2_X1 U10293 ( .A1(n8103), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n7952) );
  INV_X1 U10294 ( .A(n12553), .ZN(n12233) );
  AND2_X1 U10295 ( .A1(n12694), .A2(n12233), .ZN(n8217) );
  OR2_X1 U10296 ( .A1(n12694), .A2(n12233), .ZN(n8219) );
  INV_X1 U10297 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10905) );
  INV_X1 U10298 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11203) );
  XNOR2_X1 U10299 ( .A(n7966), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n10503) );
  NAND2_X1 U10300 ( .A1(n10503), .A2(n8099), .ZN(n7958) );
  INV_X1 U10301 ( .A(SI_20_), .ZN(n10505) );
  OR2_X1 U10302 ( .A1(n7673), .A2(n10505), .ZN(n7957) );
  INV_X1 U10303 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n12194) );
  OR2_X1 U10304 ( .A1(n7959), .A2(n12194), .ZN(n7960) );
  NAND2_X1 U10305 ( .A1(n7972), .A2(n7960), .ZN(n12527) );
  NAND2_X1 U10306 ( .A1(n12527), .A2(n7991), .ZN(n7965) );
  INV_X1 U10307 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n12687) );
  NAND2_X1 U10308 ( .A1(n8102), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n7962) );
  NAND2_X1 U10309 ( .A1(n8103), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n7961) );
  OAI211_X1 U10310 ( .C1(n7700), .C2(n12687), .A(n7962), .B(n7961), .ZN(n7963)
         );
  INV_X1 U10311 ( .A(n7963), .ZN(n7964) );
  XNOR2_X1 U10312 ( .A(n12626), .B(n12535), .ZN(n12521) );
  INV_X1 U10313 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11293) );
  NAND2_X1 U10314 ( .A1(n7967), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7968) );
  INV_X1 U10315 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11278) );
  XNOR2_X1 U10316 ( .A(n11278), .B(P1_DATAO_REG_21__SCAN_IN), .ZN(n7978) );
  XNOR2_X1 U10317 ( .A(n7980), .B(n7978), .ZN(n11951) );
  NAND2_X1 U10318 ( .A1(n11951), .A2(n8099), .ZN(n7971) );
  INV_X1 U10319 ( .A(SI_21_), .ZN(n11953) );
  OR2_X1 U10320 ( .A1(n7673), .A2(n11953), .ZN(n7970) );
  NAND2_X1 U10321 ( .A1(n7972), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n7973) );
  NAND2_X1 U10322 ( .A1(n7989), .A2(n7973), .ZN(n12515) );
  INV_X1 U10323 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n7976) );
  NAND2_X1 U10324 ( .A1(n8102), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n7975) );
  NAND2_X1 U10325 ( .A1(n8103), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n7974) );
  OAI211_X1 U10326 ( .C1(n7700), .C2(n7976), .A(n7975), .B(n7974), .ZN(n7977)
         );
  AOI21_X1 U10327 ( .B1(n12515), .B2(n7991), .A(n7977), .ZN(n12202) );
  NAND2_X1 U10328 ( .A1(n12683), .A2(n12202), .ZN(n8227) );
  OR2_X1 U10329 ( .A1(n12683), .A2(n12202), .ZN(n8226) );
  INV_X1 U10330 ( .A(n7978), .ZN(n7979) );
  NAND2_X1 U10331 ( .A1(n11278), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n7981) );
  INV_X1 U10332 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11943) );
  NAND2_X1 U10333 ( .A1(n11943), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n7998) );
  INV_X1 U10334 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7982) );
  NAND2_X1 U10335 ( .A1(n7982), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n7983) );
  NAND2_X1 U10336 ( .A1(n7998), .A2(n7983), .ZN(n7984) );
  NAND2_X1 U10337 ( .A1(n7985), .A2(n7984), .ZN(n7986) );
  NAND2_X1 U10338 ( .A1(n7999), .A2(n7986), .ZN(n10637) );
  NAND2_X1 U10339 ( .A1(n10637), .A2(n8099), .ZN(n7988) );
  INV_X1 U10340 ( .A(SI_22_), .ZN(n8700) );
  OR2_X1 U10341 ( .A1(n7673), .A2(n8700), .ZN(n7987) );
  NAND2_X1 U10342 ( .A1(n7989), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n7990) );
  INV_X1 U10343 ( .A(n8009), .ZN(n8008) );
  NAND2_X1 U10344 ( .A1(n7990), .A2(n8008), .ZN(n12504) );
  NAND2_X1 U10345 ( .A1(n12504), .A2(n7991), .ZN(n7996) );
  INV_X1 U10346 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13711) );
  NAND2_X1 U10347 ( .A1(n8045), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n7993) );
  NAND2_X1 U10348 ( .A1(n8103), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n7992) );
  OAI211_X1 U10349 ( .C1(n6690), .C2(n13711), .A(n7993), .B(n7992), .ZN(n7994)
         );
  INV_X1 U10350 ( .A(n7994), .ZN(n7995) );
  NAND2_X1 U10351 ( .A1(n7996), .A2(n7995), .ZN(n12386) );
  NAND2_X1 U10352 ( .A1(n12387), .A2(n12488), .ZN(n8231) );
  INV_X1 U10353 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8000) );
  NAND2_X1 U10354 ( .A1(n8000), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8016) );
  INV_X1 U10355 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8001) );
  NAND2_X1 U10356 ( .A1(n8001), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8002) );
  AND2_X1 U10357 ( .A1(n8016), .A2(n8002), .ZN(n8003) );
  OR2_X1 U10358 ( .A1(n8004), .A2(n8003), .ZN(n8005) );
  NAND2_X1 U10359 ( .A1(n8017), .A2(n8005), .ZN(n10967) );
  NAND2_X1 U10360 ( .A1(n10967), .A2(n8099), .ZN(n8007) );
  INV_X1 U10361 ( .A(SI_23_), .ZN(n10970) );
  OR2_X1 U10362 ( .A1(n7673), .A2(n10970), .ZN(n8006) );
  NAND2_X1 U10363 ( .A1(n8045), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8014) );
  NAND2_X1 U10364 ( .A1(n8102), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8013) );
  NAND2_X1 U10365 ( .A1(P3_REG3_REG_23__SCAN_IN), .A2(n8008), .ZN(n8010) );
  INV_X1 U10366 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n13725) );
  NAND2_X1 U10367 ( .A1(n13725), .A2(n8009), .ZN(n8020) );
  NAND2_X1 U10368 ( .A1(n8010), .A2(n8020), .ZN(n12493) );
  NAND2_X1 U10369 ( .A1(n7991), .A2(n12493), .ZN(n8012) );
  NAND2_X1 U10370 ( .A1(n8103), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8011) );
  NAND2_X1 U10371 ( .A1(n12492), .A2(n12203), .ZN(n8015) );
  NAND2_X1 U10372 ( .A1(n8237), .A2(n8015), .ZN(n12490) );
  INV_X1 U10373 ( .A(n12490), .ZN(n8234) );
  XNOR2_X1 U10374 ( .A(n8026), .B(P2_DATAO_REG_24__SCAN_IN), .ZN(n11219) );
  NAND2_X1 U10375 ( .A1(n11219), .A2(n8099), .ZN(n8019) );
  INV_X1 U10376 ( .A(SI_24_), .ZN(n11220) );
  OR2_X1 U10377 ( .A1(n7673), .A2(n11220), .ZN(n8018) );
  NAND2_X1 U10378 ( .A1(n8102), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8025) );
  NAND2_X1 U10379 ( .A1(n8045), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8024) );
  NAND2_X1 U10380 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(n8020), .ZN(n8021) );
  NAND2_X1 U10381 ( .A1(n8021), .A2(n8033), .ZN(n12481) );
  NAND2_X1 U10382 ( .A1(n8085), .A2(n12481), .ZN(n8023) );
  NAND2_X1 U10383 ( .A1(n8103), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8022) );
  NAND4_X1 U10384 ( .A1(n8025), .A2(n8024), .A3(n8023), .A4(n8022), .ZN(n12465) );
  OR2_X1 U10385 ( .A1(n12392), .A2(n12489), .ZN(n8236) );
  NAND2_X1 U10386 ( .A1(n12392), .A2(n12489), .ZN(n8235) );
  NAND2_X1 U10387 ( .A1(n8236), .A2(n8235), .ZN(n12478) );
  INV_X1 U10388 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n12136) );
  INV_X1 U10389 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11448) );
  INV_X1 U10390 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n11519) );
  XNOR2_X1 U10391 ( .A(n11519), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n8030) );
  XNOR2_X1 U10392 ( .A(n8040), .B(n8030), .ZN(n11322) );
  NAND2_X1 U10393 ( .A1(n11322), .A2(n8099), .ZN(n8032) );
  INV_X1 U10394 ( .A(SI_25_), .ZN(n11324) );
  OR2_X1 U10395 ( .A1(n7673), .A2(n11324), .ZN(n8031) );
  NAND2_X1 U10396 ( .A1(n8102), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8038) );
  NAND2_X1 U10397 ( .A1(n8045), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8037) );
  AND2_X1 U10398 ( .A1(P3_REG3_REG_25__SCAN_IN), .A2(n8033), .ZN(n8034) );
  OR2_X1 U10399 ( .A1(n8034), .A2(n8046), .ZN(n12469) );
  NAND2_X1 U10400 ( .A1(n8085), .A2(n12469), .ZN(n8036) );
  NAND2_X1 U10401 ( .A1(n8103), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8035) );
  OR2_X1 U10402 ( .A1(n12396), .A2(n12448), .ZN(n8240) );
  NAND2_X1 U10403 ( .A1(n12396), .A2(n12448), .ZN(n8241) );
  INV_X1 U10404 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n11516) );
  AND2_X1 U10405 ( .A1(n11516), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8039) );
  NAND2_X1 U10406 ( .A1(n11519), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8041) );
  INV_X1 U10407 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n11703) );
  INV_X1 U10408 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n13524) );
  AOI22_X1 U10409 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n11703), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n13524), .ZN(n8042) );
  XNOR2_X1 U10410 ( .A(n8053), .B(n8042), .ZN(n11430) );
  NAND2_X1 U10411 ( .A1(n11430), .A2(n8099), .ZN(n8044) );
  INV_X1 U10412 ( .A(SI_26_), .ZN(n11432) );
  OR2_X1 U10413 ( .A1(n7673), .A2(n11432), .ZN(n8043) );
  NAND2_X1 U10414 ( .A1(n8045), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8051) );
  NAND2_X1 U10415 ( .A1(n8103), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8050) );
  INV_X1 U10416 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n12223) );
  NOR2_X1 U10417 ( .A1(n8046), .A2(n12223), .ZN(n8047) );
  NAND2_X1 U10418 ( .A1(n7991), .A2(n12454), .ZN(n8049) );
  NAND2_X1 U10419 ( .A1(n8102), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8048) );
  NAND4_X1 U10420 ( .A1(n8051), .A2(n8050), .A3(n8049), .A4(n8048), .ZN(n12464) );
  NAND2_X1 U10421 ( .A1(n12398), .A2(n9397), .ZN(n8246) );
  NAND2_X1 U10422 ( .A1(n8245), .A2(n8246), .ZN(n12447) );
  NOR2_X1 U10423 ( .A1(n13524), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8052) );
  NAND2_X1 U10424 ( .A1(n13524), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8054) );
  INV_X1 U10425 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n11791) );
  INV_X1 U10426 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n11833) );
  AOI22_X1 U10427 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n11791), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n11833), .ZN(n8055) );
  INV_X1 U10428 ( .A(n8055), .ZN(n8056) );
  XNOR2_X1 U10429 ( .A(n8066), .B(n8056), .ZN(n11533) );
  NAND2_X1 U10430 ( .A1(n11533), .A2(n8099), .ZN(n8058) );
  INV_X1 U10431 ( .A(SI_27_), .ZN(n11534) );
  OR2_X1 U10432 ( .A1(n7673), .A2(n11534), .ZN(n8057) );
  NAND2_X2 U10433 ( .A1(n8058), .A2(n8057), .ZN(n12591) );
  NAND2_X1 U10434 ( .A1(n8045), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8064) );
  NAND2_X1 U10435 ( .A1(n8103), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8063) );
  INV_X1 U10436 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n9398) );
  NOR2_X1 U10437 ( .A1(n8059), .A2(n9398), .ZN(n8060) );
  NAND2_X1 U10438 ( .A1(n7991), .A2(n12438), .ZN(n8062) );
  NAND2_X1 U10439 ( .A1(n8102), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8061) );
  NAND4_X1 U10440 ( .A1(n8064), .A2(n8063), .A3(n8062), .A4(n8061), .ZN(n12422) );
  NOR2_X1 U10441 ( .A1(n11791), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8065) );
  NAND2_X1 U10442 ( .A1(n11791), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8067) );
  INV_X1 U10443 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12007) );
  INV_X1 U10444 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13634) );
  AOI22_X1 U10445 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(
        P2_DATAO_REG_28__SCAN_IN), .B1(n12007), .B2(n13634), .ZN(n8068) );
  XNOR2_X1 U10446 ( .A(n8078), .B(n8068), .ZN(n11537) );
  INV_X1 U10447 ( .A(SI_28_), .ZN(n11536) );
  OR2_X1 U10448 ( .A1(n7673), .A2(n11536), .ZN(n8069) );
  NAND2_X2 U10449 ( .A1(n8070), .A2(n8069), .ZN(n12426) );
  NAND2_X1 U10450 ( .A1(n8045), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8076) );
  NAND2_X1 U10451 ( .A1(n8102), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8075) );
  INV_X1 U10452 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n13684) );
  NAND2_X1 U10453 ( .A1(n8071), .A2(n13684), .ZN(n12358) );
  OR2_X1 U10454 ( .A1(n8071), .A2(n13684), .ZN(n8072) );
  NAND2_X1 U10455 ( .A1(n12358), .A2(n8072), .ZN(n12427) );
  NAND2_X1 U10456 ( .A1(n7991), .A2(n12427), .ZN(n8074) );
  NAND2_X1 U10457 ( .A1(n7667), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8073) );
  NAND2_X1 U10458 ( .A1(n12426), .A2(n12402), .ZN(n8133) );
  NAND2_X1 U10459 ( .A1(n12591), .A2(n12449), .ZN(n12416) );
  NAND2_X1 U10460 ( .A1(n8133), .A2(n12416), .ZN(n8250) );
  INV_X1 U10461 ( .A(n12409), .ZN(n8109) );
  NOR2_X1 U10462 ( .A1(n12007), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8077) );
  NAND2_X1 U10463 ( .A1(n12007), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8079) );
  XNOR2_X1 U10464 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n8080) );
  NAND2_X1 U10465 ( .A1(n8090), .A2(n8082), .ZN(n11990) );
  INV_X1 U10466 ( .A(SI_29_), .ZN(n11993) );
  OR2_X1 U10467 ( .A1(n7673), .A2(n11993), .ZN(n8083) );
  INV_X1 U10468 ( .A(n12358), .ZN(n12411) );
  NAND2_X1 U10469 ( .A1(n8085), .A2(n12411), .ZN(n8107) );
  NAND2_X1 U10470 ( .A1(n8045), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8088) );
  NAND2_X1 U10471 ( .A1(n8103), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8087) );
  NAND2_X1 U10472 ( .A1(n8102), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8086) );
  INV_X1 U10473 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14670) );
  NAND2_X1 U10474 ( .A1(n14670), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8089) );
  NAND2_X1 U10475 ( .A1(n8090), .A2(n8089), .ZN(n8098) );
  INV_X1 U10476 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n11986) );
  XNOR2_X1 U10477 ( .A(n11986), .B(P1_DATAO_REG_30__SCAN_IN), .ZN(n8097) );
  OAI22_X1 U10478 ( .A1(n8098), .A2(n8097), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(n11986), .ZN(n8092) );
  XNOR2_X1 U10479 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n8091) );
  XNOR2_X1 U10480 ( .A(n8092), .B(n8091), .ZN(n12720) );
  NOR2_X1 U10481 ( .A1(n7673), .A2(n13683), .ZN(n8093) );
  NAND2_X1 U10482 ( .A1(n8102), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n8096) );
  NAND2_X1 U10483 ( .A1(n8045), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n8095) );
  NAND2_X1 U10484 ( .A1(n7667), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n8094) );
  NAND4_X1 U10485 ( .A1(n8107), .A2(n8096), .A3(n8095), .A4(n8094), .ZN(n12356) );
  AND2_X1 U10486 ( .A1(n12654), .A2(n12356), .ZN(n8256) );
  XNOR2_X1 U10487 ( .A(n8098), .B(n8097), .ZN(n12722) );
  NAND2_X1 U10488 ( .A1(n12722), .A2(n8099), .ZN(n8101) );
  INV_X1 U10489 ( .A(SI_30_), .ZN(n12724) );
  OR2_X1 U10490 ( .A1(n7673), .A2(n12724), .ZN(n8100) );
  NAND2_X1 U10491 ( .A1(n8101), .A2(n8100), .ZN(n14771) );
  INV_X1 U10492 ( .A(n14771), .ZN(n12362) );
  NAND2_X1 U10493 ( .A1(n8102), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8106) );
  NAND2_X1 U10494 ( .A1(n8045), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8105) );
  NAND2_X1 U10495 ( .A1(n8103), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8104) );
  AND4_X1 U10496 ( .A1(n8107), .A2(n8106), .A3(n8105), .A4(n8104), .ZN(n12404)
         );
  NAND2_X1 U10497 ( .A1(n14771), .A2(n12404), .ZN(n8131) );
  NAND2_X1 U10498 ( .A1(n12410), .A2(n12232), .ZN(n8132) );
  AND2_X1 U10499 ( .A1(n8131), .A2(n8132), .ZN(n8254) );
  OAI21_X1 U10500 ( .B1(n12362), .B2(n12356), .A(n8254), .ZN(n8108) );
  INV_X1 U10501 ( .A(n12404), .ZN(n12231) );
  NAND2_X1 U10502 ( .A1(n12362), .A2(n12231), .ZN(n8130) );
  AOI21_X1 U10503 ( .B1(n12356), .B2(n8130), .A(n12654), .ZN(n8110) );
  NOR2_X1 U10504 ( .A1(n8111), .A2(n8110), .ZN(n8113) );
  NAND2_X1 U10505 ( .A1(n8115), .A2(n8114), .ZN(n8126) );
  INV_X1 U10506 ( .A(n8126), .ZN(n8117) );
  INV_X1 U10507 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8116) );
  NAND2_X1 U10508 ( .A1(n8117), .A2(n8116), .ZN(n8128) );
  NAND2_X1 U10509 ( .A1(n8121), .A2(n8120), .ZN(n8146) );
  NAND2_X1 U10510 ( .A1(n8126), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8127) );
  NAND2_X1 U10511 ( .A1(n10542), .A2(n10448), .ZN(n10440) );
  OAI21_X1 U10512 ( .B1(n12654), .B2(n12356), .A(n8130), .ZN(n8253) );
  NAND2_X1 U10513 ( .A1(n8252), .A2(n8132), .ZN(n12408) );
  AND2_X2 U10514 ( .A1(n8249), .A2(n8133), .ZN(n12419) );
  NAND2_X1 U10515 ( .A1(n8230), .A2(n8231), .ZN(n12503) );
  OR2_X1 U10516 ( .A1(n12694), .A2(n12553), .ZN(n12379) );
  INV_X1 U10517 ( .A(n12379), .ZN(n8134) );
  AND2_X1 U10518 ( .A1(n12694), .A2(n12553), .ZN(n12376) );
  NOR2_X1 U10519 ( .A1(n8134), .A2(n12376), .ZN(n12536) );
  AND2_X1 U10520 ( .A1(n15367), .A2(n11950), .ZN(n8152) );
  NOR2_X1 U10521 ( .A1(n8135), .A2(n8152), .ZN(n10907) );
  NAND4_X1 U10522 ( .A1(n15336), .A2(n7214), .A3(n8171), .A4(n10907), .ZN(
        n8136) );
  NAND3_X1 U10523 ( .A1(n8137), .A2(n10728), .A3(n15349), .ZN(n8138) );
  XNOR2_X1 U10524 ( .A(n11329), .B(n11287), .ZN(n11248) );
  OR4_X1 U10525 ( .A1(n8138), .A2(n11351), .A3(n11336), .A4(n11248), .ZN(n8139) );
  OR2_X1 U10526 ( .A1(n8196), .A2(n6735), .ZN(n11571) );
  NOR4_X1 U10527 ( .A1(n8139), .A2(n8197), .A3(n11568), .A4(n11571), .ZN(n8140) );
  NAND4_X1 U10528 ( .A1(n8140), .A2(n11712), .A3(n11806), .A4(n12574), .ZN(
        n8141) );
  NOR4_X1 U10529 ( .A1(n12503), .A2(n12536), .A3(n12375), .A4(n8141), .ZN(
        n8142) );
  INV_X1 U10530 ( .A(n12521), .ZN(n12526) );
  NAND4_X1 U10531 ( .A1(n8234), .A2(n12513), .A3(n8142), .A4(n12526), .ZN(
        n8143) );
  NOR4_X1 U10532 ( .A1(n12447), .A2(n12462), .A3(n12478), .A4(n8143), .ZN(
        n8144) );
  NAND2_X1 U10533 ( .A1(n10504), .A2(n6687), .ZN(n10449) );
  INV_X1 U10534 ( .A(n10449), .ZN(n10423) );
  NAND2_X1 U10535 ( .A1(n10504), .A2(n9145), .ZN(n10428) );
  NAND2_X1 U10536 ( .A1(n8146), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8147) );
  MUX2_X1 U10537 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8147), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n8148) );
  NAND2_X1 U10538 ( .A1(n8148), .A2(n8259), .ZN(n10635) );
  INV_X1 U10539 ( .A(n8157), .ZN(n8149) );
  AOI21_X1 U10540 ( .B1(n15365), .B2(n15360), .A(n8149), .ZN(n8159) );
  INV_X1 U10541 ( .A(n8152), .ZN(n8150) );
  OAI22_X1 U10542 ( .A1(n8135), .A2(n10542), .B1(n10427), .B2(n8150), .ZN(
        n8155) );
  INV_X1 U10543 ( .A(n8151), .ZN(n8154) );
  AOI21_X1 U10544 ( .B1(n8161), .B2(n8156), .A(n9267), .ZN(n8158) );
  OAI211_X1 U10545 ( .C1(n8161), .C2(n10458), .A(n8160), .B(n7214), .ZN(n8166)
         );
  NAND3_X1 U10546 ( .A1(n8166), .A2(n10728), .A3(n8162), .ZN(n8164) );
  NAND3_X1 U10547 ( .A1(n8164), .A2(n8168), .A3(n8163), .ZN(n8170) );
  NAND3_X1 U10548 ( .A1(n8166), .A2(n10728), .A3(n8165), .ZN(n8167) );
  OAI211_X1 U10549 ( .C1(n10860), .C2(n10802), .A(n8167), .B(n8172), .ZN(n8169) );
  MUX2_X1 U10550 ( .A(n8174), .B(n8173), .S(n9267), .Z(n8175) );
  INV_X1 U10551 ( .A(n11248), .ZN(n8180) );
  MUX2_X1 U10552 ( .A(n8178), .B(n8177), .S(n9267), .Z(n8179) );
  AND3_X1 U10553 ( .A1(n8181), .A2(n8180), .A3(n8179), .ZN(n8185) );
  NOR2_X1 U10554 ( .A1(n11329), .A2(n10458), .ZN(n8183) );
  NOR2_X1 U10555 ( .A1(n11095), .A2(n9267), .ZN(n8182) );
  MUX2_X1 U10556 ( .A(n8183), .B(n8182), .S(n11287), .Z(n8184) );
  NOR4_X1 U10557 ( .A1(n8185), .A2(n8184), .A3(n11351), .A4(n11336), .ZN(n8195) );
  OAI211_X1 U10558 ( .C1(n11351), .C2(n8187), .A(n8192), .B(n8186), .ZN(n8190)
         );
  OAI211_X1 U10559 ( .C1(n11351), .C2(n11350), .A(n8191), .B(n8188), .ZN(n8189) );
  MUX2_X1 U10560 ( .A(n8190), .B(n8189), .S(n9267), .Z(n8194) );
  MUX2_X1 U10561 ( .A(n8192), .B(n8191), .S(n10458), .Z(n8193) );
  OAI21_X1 U10562 ( .B1(n8195), .B2(n8194), .A(n8193), .ZN(n8199) );
  INV_X1 U10563 ( .A(n11571), .ZN(n11575) );
  MUX2_X1 U10564 ( .A(n8196), .B(n6735), .S(n10458), .Z(n8198) );
  AOI211_X1 U10565 ( .C1(n8199), .C2(n11575), .A(n8198), .B(n8197), .ZN(n8205)
         );
  INV_X1 U10566 ( .A(n8213), .ZN(n8209) );
  OAI211_X1 U10567 ( .C1(n8209), .C2(n8208), .A(n9267), .B(n8207), .ZN(n8210)
         );
  OR2_X1 U10568 ( .A1(n8210), .A2(n8217), .ZN(n8212) );
  INV_X1 U10569 ( .A(n8212), .ZN(n8215) );
  AND3_X1 U10570 ( .A1(n8219), .A2(n8213), .A3(n10458), .ZN(n8214) );
  OAI22_X1 U10571 ( .A1(n8216), .A2(n12375), .B1(n8215), .B2(n8214), .ZN(n8221) );
  INV_X1 U10572 ( .A(n8217), .ZN(n8218) );
  MUX2_X1 U10573 ( .A(n8219), .B(n8218), .S(n10458), .Z(n8220) );
  NAND2_X1 U10574 ( .A1(n8221), .A2(n8220), .ZN(n8225) );
  INV_X1 U10575 ( .A(n12535), .ZN(n12381) );
  NAND2_X1 U10576 ( .A1(n12381), .A2(n9267), .ZN(n8223) );
  NAND2_X1 U10577 ( .A1(n12535), .A2(n10458), .ZN(n8222) );
  MUX2_X1 U10578 ( .A(n8223), .B(n8222), .S(n12626), .Z(n8224) );
  OAI211_X1 U10579 ( .C1(n8225), .C2(n12521), .A(n12513), .B(n8224), .ZN(n8229) );
  MUX2_X1 U10580 ( .A(n8227), .B(n8226), .S(n10458), .Z(n8228) );
  MUX2_X1 U10581 ( .A(n8231), .B(n8230), .S(n10458), .Z(n8232) );
  AND2_X1 U10582 ( .A1(n12203), .A2(n9267), .ZN(n8233) );
  INV_X1 U10583 ( .A(n8235), .ZN(n8239) );
  AOI21_X1 U10584 ( .B1(n8237), .B2(n8236), .A(n8239), .ZN(n8238) );
  MUX2_X1 U10585 ( .A(n8239), .B(n8238), .S(n10458), .Z(n8243) );
  MUX2_X1 U10586 ( .A(n8241), .B(n8240), .S(n9267), .Z(n8242) );
  OAI211_X1 U10587 ( .C1(n8244), .C2(n8243), .A(n7465), .B(n8242), .ZN(n8248)
         );
  MUX2_X1 U10588 ( .A(n8246), .B(n8245), .S(n10458), .Z(n8247) );
  OAI21_X1 U10589 ( .B1(n8250), .B2(n10458), .A(n8249), .ZN(n8251) );
  NAND2_X1 U10590 ( .A1(n8259), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8258) );
  MUX2_X1 U10591 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8258), .S(
        P3_IR_REG_23__SCAN_IN), .Z(n8262) );
  INV_X1 U10592 ( .A(n8259), .ZN(n8261) );
  NAND2_X1 U10593 ( .A1(n8262), .A2(n8269), .ZN(n9972) );
  OR2_X1 U10594 ( .A1(n9972), .A2(P3_U3151), .ZN(n10968) );
  INV_X1 U10595 ( .A(n12354), .ZN(n9975) );
  NAND2_X1 U10596 ( .A1(n9975), .A2(n12340), .ZN(n9976) );
  NAND2_X1 U10597 ( .A1(n9976), .A2(n9973), .ZN(n9260) );
  INV_X1 U10598 ( .A(n9260), .ZN(n8265) );
  NAND2_X1 U10599 ( .A1(n8269), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8270) );
  MUX2_X1 U10600 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8270), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8271) );
  NAND2_X1 U10601 ( .A1(n8271), .A2(n8273), .ZN(n9147) );
  INV_X1 U10602 ( .A(n9147), .ZN(n11218) );
  NAND2_X1 U10603 ( .A1(n8273), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8272) );
  INV_X1 U10604 ( .A(n9148), .ZN(n8276) );
  NAND3_X1 U10605 ( .A1(n9232), .A2(n11218), .A3(n8276), .ZN(n9406) );
  NAND4_X1 U10606 ( .A1(n12406), .A2(n10423), .A3(n9975), .A4(n10540), .ZN(
        n8277) );
  OAI211_X1 U10607 ( .C1(n10427), .C2(n10968), .A(n8277), .B(P3_B_REG_SCAN_IN), 
        .ZN(n8278) );
  NAND3_X1 U10608 ( .A1(n8572), .A2(n8569), .A3(n8279), .ZN(n8280) );
  NOR2_X1 U10609 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n8285) );
  NAND4_X1 U10610 ( .A1(n8285), .A2(n8284), .A3(n8283), .A4(n8282), .ZN(n8286)
         );
  NOR2_X2 U10611 ( .A1(n8438), .A2(n8286), .ZN(n8570) );
  NAND2_X1 U10612 ( .A1(n8287), .A2(n8570), .ZN(n8866) );
  INV_X1 U10613 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n8291) );
  NAND2_X1 U10614 ( .A1(n8384), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8293) );
  MUX2_X1 U10615 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8293), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n8294) );
  AND2_X2 U10616 ( .A1(n8295), .A2(n8296), .ZN(n8456) );
  NAND2_X1 U10617 ( .A1(n8781), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8304) );
  BUF_X4 U10618 ( .A(n8460), .Z(n9063) );
  NAND2_X1 U10619 ( .A1(n9063), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8303) );
  INV_X1 U10620 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n14167) );
  NAND2_X1 U10621 ( .A1(n8470), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8484) );
  NAND2_X1 U10622 ( .A1(n8528), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8547) );
  INV_X1 U10623 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n8559) );
  NAND2_X1 U10624 ( .A1(n8577), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8587) );
  INV_X1 U10625 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n11211) );
  INV_X1 U10626 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8608) );
  NAND2_X1 U10627 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n8298) );
  INV_X1 U10628 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n14180) );
  INV_X1 U10629 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n14132) );
  AOI21_X1 U10630 ( .B1(n14167), .B2(n8300), .A(n8739), .ZN(n14414) );
  NAND2_X1 U10631 ( .A1(n8785), .A2(n14414), .ZN(n8302) );
  NAND2_X1 U10632 ( .A1(n9064), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n8301) );
  NAND4_X1 U10633 ( .A1(n8304), .A2(n8303), .A3(n8302), .A4(n8301), .ZN(n14235) );
  INV_X1 U10634 ( .A(n14235), .ZN(n8728) );
  INV_X1 U10635 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9492) );
  AND2_X1 U10636 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8306) );
  NAND2_X1 U10637 ( .A1(n9910), .A2(n8306), .ZN(n8408) );
  AND2_X1 U10638 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8307) );
  NAND2_X1 U10639 ( .A1(n8310), .A2(n8307), .ZN(n9797) );
  NAND2_X1 U10640 ( .A1(n8408), .A2(n9797), .ZN(n8393) );
  NOR2_X1 U10641 ( .A1(n8308), .A2(n9512), .ZN(n8309) );
  MUX2_X1 U10642 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n8310), .Z(n8312) );
  INV_X1 U10643 ( .A(n8417), .ZN(n8311) );
  NAND2_X1 U10644 ( .A1(n8312), .A2(SI_2_), .ZN(n8313) );
  MUX2_X1 U10645 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n8310), .Z(n8315) );
  XNOR2_X1 U10646 ( .A(n8315), .B(SI_3_), .ZN(n8430) );
  NAND2_X1 U10647 ( .A1(n8315), .A2(SI_3_), .ZN(n8316) );
  NAND2_X1 U10648 ( .A1(n8319), .A2(SI_4_), .ZN(n8320) );
  MUX2_X1 U10649 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n9794), .Z(n8326) );
  NAND2_X1 U10650 ( .A1(n8326), .A2(SI_6_), .ZN(n8327) );
  MUX2_X1 U10651 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n9794), .Z(n8329) );
  NAND2_X1 U10652 ( .A1(n8329), .A2(SI_7_), .ZN(n8330) );
  MUX2_X1 U10653 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n9794), .Z(n8331) );
  MUX2_X1 U10654 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n9794), .Z(n8333) );
  NAND2_X1 U10655 ( .A1(n8333), .A2(SI_9_), .ZN(n8334) );
  MUX2_X1 U10656 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n9794), .Z(n8535) );
  INV_X1 U10657 ( .A(n8535), .ZN(n8335) );
  INV_X1 U10658 ( .A(SI_10_), .ZN(n9499) );
  MUX2_X1 U10659 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n9794), .Z(n8337) );
  OAI21_X1 U10660 ( .B1(n8335), .B2(n9499), .A(n8539), .ZN(n8336) );
  NOR2_X1 U10661 ( .A1(n8535), .A2(SI_10_), .ZN(n8340) );
  INV_X1 U10662 ( .A(n8337), .ZN(n8338) );
  NAND2_X1 U10663 ( .A1(n8338), .A2(n9511), .ZN(n8538) );
  INV_X1 U10664 ( .A(n8538), .ZN(n8339) );
  MUX2_X1 U10665 ( .A(n9727), .B(n9731), .S(n9794), .Z(n8342) );
  INV_X1 U10666 ( .A(n8342), .ZN(n8343) );
  NAND2_X1 U10667 ( .A1(n8343), .A2(SI_12_), .ZN(n8344) );
  MUX2_X1 U10668 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n9794), .Z(n8346) );
  NAND2_X1 U10669 ( .A1(n8346), .A2(SI_13_), .ZN(n8347) );
  MUX2_X1 U10670 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n9794), .Z(n8594) );
  INV_X1 U10671 ( .A(n8594), .ZN(n8349) );
  MUX2_X1 U10672 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n9794), .Z(n8351) );
  NOR2_X1 U10673 ( .A1(n8594), .A2(SI_14_), .ZN(n8354) );
  INV_X1 U10674 ( .A(n8351), .ZN(n8352) );
  INV_X1 U10675 ( .A(SI_15_), .ZN(n13779) );
  NAND2_X1 U10676 ( .A1(n8352), .A2(n13779), .ZN(n8599) );
  INV_X1 U10677 ( .A(n8599), .ZN(n8353) );
  MUX2_X1 U10678 ( .A(n8356), .B(n13518), .S(n9794), .Z(n8357) );
  INV_X1 U10679 ( .A(SI_16_), .ZN(n9809) );
  NAND2_X1 U10680 ( .A1(n8357), .A2(n9809), .ZN(n8360) );
  INV_X1 U10681 ( .A(n8357), .ZN(n8358) );
  NAND2_X1 U10682 ( .A1(n8358), .A2(SI_16_), .ZN(n8359) );
  INV_X1 U10683 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10345) );
  MUX2_X1 U10684 ( .A(n8362), .B(n10345), .S(n9794), .Z(n8363) );
  INV_X1 U10685 ( .A(SI_17_), .ZN(n9887) );
  NAND2_X1 U10686 ( .A1(n8363), .A2(n9887), .ZN(n8366) );
  INV_X1 U10687 ( .A(n8363), .ZN(n8364) );
  NAND2_X1 U10688 ( .A1(n8364), .A2(SI_17_), .ZN(n8365) );
  INV_X1 U10689 ( .A(SI_18_), .ZN(n10002) );
  MUX2_X1 U10690 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n9794), .Z(n8642) );
  INV_X1 U10691 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10841) );
  MUX2_X1 U10692 ( .A(n10905), .B(n10841), .S(n9794), .Z(n8370) );
  NAND2_X1 U10693 ( .A1(n8370), .A2(n11994), .ZN(n8373) );
  INV_X1 U10694 ( .A(n8370), .ZN(n8371) );
  NAND2_X1 U10695 ( .A1(n8371), .A2(SI_19_), .ZN(n8372) );
  MUX2_X1 U10696 ( .A(n11293), .B(n11203), .S(n9794), .Z(n8674) );
  MUX2_X1 U10697 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9794), .Z(n8689) );
  NOR2_X1 U10698 ( .A1(n8674), .A2(n10505), .ZN(n8374) );
  AOI22_X1 U10699 ( .A1(n8374), .A2(n7600), .B1(n8689), .B2(SI_21_), .ZN(n8375) );
  MUX2_X1 U10700 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n9794), .Z(n8709) );
  MUX2_X1 U10701 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n9794), .Z(n8713) );
  INV_X1 U10702 ( .A(n8713), .ZN(n8377) );
  NAND2_X1 U10703 ( .A1(n8377), .A2(n10970), .ZN(n8380) );
  OAI21_X1 U10704 ( .B1(SI_22_), .B2(n8709), .A(n8380), .ZN(n8378) );
  INV_X1 U10705 ( .A(n8378), .ZN(n8379) );
  INV_X1 U10706 ( .A(n8709), .ZN(n11940) );
  NOR2_X1 U10707 ( .A1(n11940), .A2(n8700), .ZN(n8381) );
  AOI22_X1 U10708 ( .A1(n8381), .A2(n8380), .B1(n8713), .B2(SI_23_), .ZN(n8382) );
  MUX2_X1 U10709 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n9794), .Z(n8729) );
  NAND2_X1 U10710 ( .A1(n12796), .A2(n6617), .ZN(n8391) );
  NAND2_X1 U10711 ( .A1(n8541), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8390) );
  XNOR2_X1 U10712 ( .A(n8392), .B(n8393), .ZN(n9909) );
  NAND2_X1 U10713 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n8394) );
  NAND2_X1 U10714 ( .A1(n8437), .A2(n9458), .ZN(n8395) );
  OAI211_X2 U10715 ( .C1(n9057), .C2(n9909), .A(n8396), .B(n8395), .ZN(n14125)
         );
  NAND2_X1 U10716 ( .A1(n8456), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8400) );
  NAND2_X1 U10717 ( .A1(n8455), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n8398) );
  NAND2_X1 U10718 ( .A1(n8460), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n8397) );
  NAND2_X1 U10719 ( .A1(n8456), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n8403) );
  NAND2_X1 U10720 ( .A1(n8460), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n8402) );
  OAI21_X1 U10721 ( .B1(n9794), .B2(n9524), .A(n8406), .ZN(n8407) );
  AND2_X1 U10722 ( .A1(n8408), .A2(n8407), .ZN(n14674) );
  OAI21_X1 U10723 ( .B1(n6821), .B2(n10246), .A(n9096), .ZN(n8412) );
  NAND2_X1 U10724 ( .A1(n10246), .A2(n6821), .ZN(n8411) );
  NAND2_X1 U10725 ( .A1(n8412), .A2(n8411), .ZN(n10233) );
  INV_X1 U10726 ( .A(n10233), .ZN(n8422) );
  NAND2_X1 U10727 ( .A1(n8456), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n8416) );
  NAND2_X1 U10728 ( .A1(n8785), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n8415) );
  NAND2_X1 U10729 ( .A1(n8460), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n8414) );
  NAND2_X1 U10730 ( .A1(n8455), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n8413) );
  NAND4_X2 U10731 ( .A1(n8416), .A2(n8415), .A3(n8414), .A4(n8413), .ZN(n14251) );
  XNOR2_X1 U10732 ( .A(n8418), .B(n8417), .ZN(n9920) );
  OR2_X1 U10733 ( .A1(n8419), .A2(n8290), .ZN(n8420) );
  XNOR2_X1 U10734 ( .A(n8420), .B(P1_IR_REG_2__SCAN_IN), .ZN(n14270) );
  NAND2_X1 U10735 ( .A1(n14251), .A2(n10594), .ZN(n8421) );
  AND2_X1 U10736 ( .A1(n8423), .A2(n8421), .ZN(n9099) );
  NAND2_X1 U10737 ( .A1(n10235), .A2(n8423), .ZN(n10821) );
  NAND2_X1 U10738 ( .A1(n8456), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n8427) );
  INV_X1 U10739 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9449) );
  NAND2_X1 U10740 ( .A1(n8785), .A2(n9449), .ZN(n8426) );
  NAND2_X1 U10741 ( .A1(n8455), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n8424) );
  NAND2_X1 U10742 ( .A1(n8428), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8429) );
  XNOR2_X1 U10743 ( .A(n8429), .B(n8281), .ZN(n9836) );
  XNOR2_X1 U10744 ( .A(n8431), .B(n8430), .ZN(n9934) );
  NAND2_X1 U10745 ( .A1(n8436), .A2(n9934), .ZN(n8433) );
  NAND2_X1 U10746 ( .A1(n8541), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8432) );
  OR2_X1 U10747 ( .A1(n14250), .A2(n7099), .ZN(n8920) );
  NAND2_X1 U10748 ( .A1(n14250), .A2(n7099), .ZN(n8919) );
  NAND2_X1 U10749 ( .A1(n8920), .A2(n8919), .ZN(n10830) );
  INV_X1 U10750 ( .A(n10830), .ZN(n10822) );
  NAND2_X1 U10751 ( .A1(n10821), .A2(n10822), .ZN(n10820) );
  NAND2_X1 U10752 ( .A1(n10820), .A2(n8920), .ZN(n10621) );
  XNOR2_X1 U10753 ( .A(n8435), .B(n8434), .ZN(n10118) );
  NAND2_X1 U10754 ( .A1(n10118), .A2(n6617), .ZN(n8441) );
  NAND2_X1 U10755 ( .A1(n8438), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8439) );
  XNOR2_X1 U10756 ( .A(n8439), .B(P1_IR_REG_4__SCAN_IN), .ZN(n14281) );
  AOI22_X1 U10757 ( .A1(n9079), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n8661), .B2(
        n14281), .ZN(n8440) );
  INV_X1 U10758 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n8442) );
  NAND2_X1 U10759 ( .A1(n9449), .A2(n8442), .ZN(n8443) );
  AND2_X1 U10760 ( .A1(n8443), .A2(n8458), .ZN(n10745) );
  NAND2_X1 U10761 ( .A1(n8785), .A2(n10745), .ZN(n8446) );
  INV_X1 U10762 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n8444) );
  OR2_X1 U10763 ( .A1(n8803), .A2(n8444), .ZN(n8445) );
  INV_X1 U10764 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n9837) );
  NAND2_X1 U10765 ( .A1(n10259), .A2(n6617), .ZN(n8454) );
  NOR2_X1 U10766 ( .A1(n8438), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n8450) );
  NOR2_X1 U10767 ( .A1(n8450), .A2(n8290), .ZN(n8448) );
  MUX2_X1 U10768 ( .A(n8290), .B(n8448), .S(P1_IR_REG_5__SCAN_IN), .Z(n8452)
         );
  INV_X1 U10769 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n8449) );
  NAND2_X1 U10770 ( .A1(n8450), .A2(n8449), .ZN(n8479) );
  INV_X1 U10771 ( .A(n8479), .ZN(n8451) );
  INV_X1 U10772 ( .A(n9884), .ZN(n9842) );
  AOI22_X1 U10773 ( .A1(n9079), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n8661), .B2(
        n9842), .ZN(n8453) );
  NAND2_X1 U10774 ( .A1(n8454), .A2(n8453), .ZN(n10934) );
  NAND2_X1 U10775 ( .A1(n8455), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n8464) );
  NAND2_X1 U10776 ( .A1(n8456), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n8463) );
  AND2_X1 U10777 ( .A1(n8458), .A2(n8457), .ZN(n8459) );
  NOR2_X1 U10778 ( .A1(n8470), .A2(n8459), .ZN(n10942) );
  NAND2_X1 U10779 ( .A1(n8785), .A2(n10942), .ZN(n8462) );
  NAND2_X1 U10780 ( .A1(n8460), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n8461) );
  NAND4_X1 U10781 ( .A1(n8464), .A2(n8463), .A3(n8462), .A4(n8461), .ZN(n14248) );
  INV_X1 U10782 ( .A(n10778), .ZN(n10779) );
  XNOR2_X1 U10783 ( .A(n8466), .B(n8465), .ZN(n10403) );
  NAND2_X1 U10784 ( .A1(n10403), .A2(n6617), .ZN(n8469) );
  NAND2_X1 U10785 ( .A1(n8479), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8467) );
  XNOR2_X1 U10786 ( .A(n8467), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9858) );
  AOI22_X1 U10787 ( .A1(n9079), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n8661), .B2(
        n9858), .ZN(n8468) );
  NAND2_X1 U10788 ( .A1(n8469), .A2(n8468), .ZN(n10964) );
  NAND2_X1 U10789 ( .A1(n8781), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n8475) );
  NAND2_X1 U10790 ( .A1(n9064), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n8474) );
  OR2_X1 U10791 ( .A1(n8470), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8471) );
  AND2_X1 U10792 ( .A1(n8484), .A2(n8471), .ZN(n10788) );
  NAND2_X1 U10793 ( .A1(n8785), .A2(n10788), .ZN(n8473) );
  NAND2_X1 U10794 ( .A1(n9063), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n8472) );
  NAND4_X1 U10795 ( .A1(n8475), .A2(n8474), .A3(n8473), .A4(n8472), .ZN(n14247) );
  OR2_X1 U10796 ( .A1(n10964), .A2(n14247), .ZN(n8816) );
  NAND2_X1 U10797 ( .A1(n10964), .A2(n14247), .ZN(n8476) );
  NAND2_X1 U10798 ( .A1(n10574), .A2(n6617), .ZN(n8482) );
  NAND2_X1 U10799 ( .A1(n8492), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8480) );
  XNOR2_X1 U10800 ( .A(n8480), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9892) );
  AOI22_X1 U10801 ( .A1(n9079), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n8661), .B2(
        n9892), .ZN(n8481) );
  INV_X1 U10802 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n8483) );
  OR2_X1 U10803 ( .A1(n8803), .A2(n8483), .ZN(n8489) );
  INV_X2 U10804 ( .A(n8706), .ZN(n8781) );
  NAND2_X1 U10805 ( .A1(n8781), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n8488) );
  NAND2_X1 U10806 ( .A1(n8484), .A2(n9866), .ZN(n8485) );
  AND2_X1 U10807 ( .A1(n8497), .A2(n8485), .ZN(n14078) );
  NAND2_X1 U10808 ( .A1(n8785), .A2(n14078), .ZN(n8487) );
  NAND2_X1 U10809 ( .A1(n9063), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n8486) );
  NAND4_X1 U10810 ( .A1(n8489), .A2(n8488), .A3(n8487), .A4(n8486), .ZN(n14246) );
  INV_X1 U10811 ( .A(n14246), .ZN(n11657) );
  XNOR2_X1 U10812 ( .A(n14954), .B(n14246), .ZN(n11013) );
  INV_X1 U10813 ( .A(n14247), .ZN(n10953) );
  NAND2_X1 U10814 ( .A1(n10964), .A2(n10953), .ZN(n11009) );
  AND2_X1 U10815 ( .A1(n11013), .A2(n11009), .ZN(n11010) );
  XNOR2_X1 U10816 ( .A(n8491), .B(n8490), .ZN(n10750) );
  NAND2_X1 U10817 ( .A1(n10750), .A2(n6617), .ZN(n8495) );
  NAND2_X1 U10818 ( .A1(n8507), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8493) );
  XNOR2_X1 U10819 ( .A(n8493), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9957) );
  AOI22_X1 U10820 ( .A1(n9079), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n8661), .B2(
        n9957), .ZN(n8494) );
  NAND2_X1 U10821 ( .A1(n9064), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n8503) );
  NAND2_X1 U10822 ( .A1(n8781), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n8502) );
  NAND2_X1 U10823 ( .A1(n8497), .A2(n8496), .ZN(n8498) );
  NAND2_X1 U10824 ( .A1(n8513), .A2(n8498), .ZN(n11960) );
  INV_X1 U10825 ( .A(n11960), .ZN(n8499) );
  NAND2_X1 U10826 ( .A1(n8785), .A2(n8499), .ZN(n8501) );
  NAND2_X1 U10827 ( .A1(n9063), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n8500) );
  NAND4_X1 U10828 ( .A1(n8503), .A2(n8502), .A3(n8501), .A4(n8500), .ZN(n14245) );
  XNOR2_X1 U10829 ( .A(n14956), .B(n14245), .ZN(n10976) );
  NAND2_X1 U10830 ( .A1(n10977), .A2(n10976), .ZN(n10975) );
  INV_X1 U10831 ( .A(n14245), .ZN(n14901) );
  OR2_X1 U10832 ( .A1(n14956), .A2(n14901), .ZN(n8504) );
  NAND2_X1 U10833 ( .A1(n10975), .A2(n8504), .ZN(n11110) );
  INV_X1 U10834 ( .A(n11110), .ZN(n8522) );
  XNOR2_X1 U10835 ( .A(n8506), .B(n8505), .ZN(n10876) );
  NAND2_X1 U10836 ( .A1(n10876), .A2(n6617), .ZN(n8511) );
  OAI21_X1 U10837 ( .B1(n8507), .B2(P1_IR_REG_8__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8543) );
  INV_X1 U10838 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8508) );
  OR2_X1 U10839 ( .A1(n8543), .A2(n8508), .ZN(n8509) );
  NAND2_X1 U10840 ( .A1(n8543), .A2(n8508), .ZN(n8524) );
  AOI22_X1 U10841 ( .A1(n9079), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n8661), .B2(
        n10290), .ZN(n8510) );
  NAND2_X1 U10842 ( .A1(n8781), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n8520) );
  INV_X1 U10843 ( .A(n8528), .ZN(n8515) );
  NAND2_X1 U10844 ( .A1(n8513), .A2(n8512), .ZN(n8514) );
  NAND2_X1 U10845 ( .A1(n8515), .A2(n8514), .ZN(n14908) );
  INV_X1 U10846 ( .A(n14908), .ZN(n11116) );
  NAND2_X1 U10847 ( .A1(n8785), .A2(n11116), .ZN(n8519) );
  INV_X1 U10848 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9958) );
  OR2_X1 U10849 ( .A1(n8804), .A2(n9958), .ZN(n8518) );
  INV_X1 U10850 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n8516) );
  OR2_X1 U10851 ( .A1(n8803), .A2(n8516), .ZN(n8517) );
  XNOR2_X1 U10852 ( .A(n11671), .B(n11681), .ZN(n11109) );
  NAND2_X1 U10853 ( .A1(n11671), .A2(n11681), .ZN(n8523) );
  XNOR2_X1 U10854 ( .A(n8534), .B(n8535), .ZN(n10987) );
  NAND2_X1 U10855 ( .A1(n10987), .A2(n6617), .ZN(n8527) );
  NAND2_X1 U10856 ( .A1(n8524), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8525) );
  XNOR2_X1 U10857 ( .A(n8525), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10553) );
  AOI22_X1 U10858 ( .A1(n9079), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n10553), 
        .B2(n8661), .ZN(n8526) );
  NAND2_X1 U10859 ( .A1(n9064), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n8533) );
  NAND2_X1 U10860 ( .A1(n8781), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8532) );
  OR2_X1 U10861 ( .A1(n8528), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8529) );
  AND2_X1 U10862 ( .A1(n8529), .A2(n8547), .ZN(n11684) );
  NAND2_X1 U10863 ( .A1(n8785), .A2(n11684), .ZN(n8531) );
  NAND2_X1 U10864 ( .A1(n9063), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n8530) );
  NAND4_X1 U10865 ( .A1(n8533), .A2(n8532), .A3(n8531), .A4(n8530), .ZN(n14243) );
  XNOR2_X1 U10866 ( .A(n14964), .B(n14243), .ZN(n9103) );
  INV_X1 U10867 ( .A(n14243), .ZN(n14898) );
  INV_X1 U10868 ( .A(n11385), .ZN(n11388) );
  NAND2_X1 U10869 ( .A1(n8536), .A2(SI_10_), .ZN(n8537) );
  NAND2_X1 U10870 ( .A1(n8539), .A2(n8538), .ZN(n8540) );
  NAND2_X1 U10871 ( .A1(n11151), .A2(n6617), .ZN(n8546) );
  OAI21_X1 U10872 ( .B1(P1_IR_REG_9__SCAN_IN), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8542) );
  NAND2_X1 U10873 ( .A1(n8543), .A2(n8542), .ZN(n8544) );
  INV_X1 U10874 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n13708) );
  XNOR2_X1 U10875 ( .A(n8544), .B(n13708), .ZN(n10712) );
  AOI22_X1 U10876 ( .A1(n9079), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n8661), 
        .B2(n10712), .ZN(n8545) );
  NAND2_X1 U10877 ( .A1(n8781), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n8553) );
  INV_X1 U10878 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11395) );
  OR2_X1 U10879 ( .A1(n8804), .A2(n11395), .ZN(n8552) );
  NAND2_X1 U10880 ( .A1(n8547), .A2(n14845), .ZN(n8548) );
  NAND2_X1 U10881 ( .A1(n8560), .A2(n8548), .ZN(n14858) );
  INV_X1 U10882 ( .A(n14858), .ZN(n8549) );
  NAND2_X1 U10883 ( .A1(n8785), .A2(n8549), .ZN(n8551) );
  NAND2_X1 U10884 ( .A1(n9064), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n8550) );
  NAND4_X1 U10885 ( .A1(n8553), .A2(n8552), .A3(n8551), .A4(n8550), .ZN(n14242) );
  INV_X1 U10886 ( .A(n14242), .ZN(n11680) );
  NOR2_X1 U10887 ( .A1(n14843), .A2(n11680), .ZN(n8953) );
  NAND2_X1 U10888 ( .A1(n14843), .A2(n11680), .ZN(n8948) );
  XNOR2_X1 U10889 ( .A(n8555), .B(n7596), .ZN(n11302) );
  NAND2_X1 U10890 ( .A1(n11302), .A2(n6617), .ZN(n8558) );
  OR2_X1 U10891 ( .A1(n8570), .A2(n8290), .ZN(n8556) );
  XNOR2_X1 U10892 ( .A(n8556), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11029) );
  AOI22_X1 U10893 ( .A1(n9079), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n8661), 
        .B2(n11029), .ZN(n8557) );
  NAND2_X1 U10894 ( .A1(n9064), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n8565) );
  NAND2_X1 U10895 ( .A1(n8781), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n8564) );
  AND2_X1 U10896 ( .A1(n8560), .A2(n8559), .ZN(n8561) );
  NOR2_X1 U10897 ( .A1(n8577), .A2(n8561), .ZN(n14704) );
  NAND2_X1 U10898 ( .A1(n8785), .A2(n14704), .ZN(n8563) );
  NAND2_X1 U10899 ( .A1(n9063), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n8562) );
  NAND4_X1 U10900 ( .A1(n8565), .A2(n8564), .A3(n8563), .A4(n8562), .ZN(n14241) );
  XNOR2_X1 U10901 ( .A(n14707), .B(n11912), .ZN(n14709) );
  XNOR2_X1 U10902 ( .A(n8568), .B(n8567), .ZN(n11358) );
  NAND2_X1 U10903 ( .A1(n11358), .A2(n6617), .ZN(n8576) );
  NOR2_X1 U10904 ( .A1(n8573), .A2(n8290), .ZN(n8571) );
  MUX2_X1 U10905 ( .A(n8290), .B(n8571), .S(P1_IR_REG_13__SCAN_IN), .Z(n8574)
         );
  INV_X1 U10906 ( .A(n11205), .ZN(n11208) );
  AOI22_X1 U10907 ( .A1(n9079), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n8661), 
        .B2(n11208), .ZN(n8575) );
  NAND2_X1 U10908 ( .A1(n9064), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n8582) );
  NAND2_X1 U10909 ( .A1(n8781), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8581) );
  OR2_X1 U10910 ( .A1(n8577), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8578) );
  AND2_X1 U10911 ( .A1(n8587), .A2(n8578), .ZN(n11935) );
  NAND2_X1 U10912 ( .A1(n8785), .A2(n11935), .ZN(n8580) );
  NAND2_X1 U10913 ( .A1(n9063), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n8579) );
  NAND4_X1 U10914 ( .A1(n8582), .A2(n8581), .A3(n8580), .A4(n8579), .ZN(n14240) );
  XNOR2_X1 U10915 ( .A(n11928), .B(n14240), .ZN(n9104) );
  INV_X1 U10916 ( .A(n14240), .ZN(n14094) );
  OR2_X1 U10917 ( .A1(n11928), .A2(n14094), .ZN(n8583) );
  XNOR2_X1 U10918 ( .A(n8596), .B(SI_14_), .ZN(n8593) );
  XNOR2_X1 U10919 ( .A(n8593), .B(n8594), .ZN(n11538) );
  NAND2_X1 U10920 ( .A1(n11538), .A2(n6617), .ZN(n8585) );
  NAND2_X1 U10921 ( .A1(n8796), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8604) );
  XNOR2_X1 U10922 ( .A(n8604), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11644) );
  AOI22_X1 U10923 ( .A1(n9079), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n8661), 
        .B2(n11644), .ZN(n8584) );
  NAND2_X1 U10924 ( .A1(n8781), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n8592) );
  INV_X1 U10925 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n8586) );
  OR2_X1 U10926 ( .A1(n8804), .A2(n8586), .ZN(n8591) );
  NAND2_X1 U10927 ( .A1(n8587), .A2(n11211), .ZN(n8588) );
  AND2_X1 U10928 ( .A1(n8609), .A2(n8588), .ZN(n14098) );
  NAND2_X1 U10929 ( .A1(n8785), .A2(n14098), .ZN(n8590) );
  NAND2_X1 U10930 ( .A1(n9064), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n8589) );
  NAND4_X1 U10931 ( .A1(n8592), .A2(n8591), .A3(n8590), .A4(n8589), .ZN(n14239) );
  INV_X1 U10932 ( .A(n14239), .ZN(n14223) );
  NOR2_X1 U10933 ( .A1(n14639), .A2(n14223), .ZN(n11815) );
  INV_X1 U10934 ( .A(n11815), .ZN(n8615) );
  INV_X1 U10935 ( .A(n8593), .ZN(n8595) );
  NAND2_X1 U10936 ( .A1(n8595), .A2(n8594), .ZN(n8598) );
  NAND2_X1 U10937 ( .A1(n8596), .A2(SI_14_), .ZN(n8597) );
  NAND2_X1 U10938 ( .A1(n8598), .A2(n8597), .ZN(n8602) );
  NAND2_X1 U10939 ( .A1(n8600), .A2(n8599), .ZN(n8601) );
  NAND2_X1 U10940 ( .A1(n11542), .A2(n6617), .ZN(n8607) );
  NAND2_X1 U10941 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), 
        .ZN(n8603) );
  NAND2_X1 U10942 ( .A1(n8604), .A2(n8603), .ZN(n8605) );
  XNOR2_X1 U10943 ( .A(n8605), .B(n7407), .ZN(n11646) );
  AOI22_X1 U10944 ( .A1(n8541), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n8661), 
        .B2(n11646), .ZN(n8606) );
  AND2_X1 U10945 ( .A1(n8609), .A2(n8608), .ZN(n8610) );
  OR2_X1 U10946 ( .A1(n8610), .A2(n8626), .ZN(n14222) );
  NAND2_X1 U10947 ( .A1(n9064), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n8612) );
  NAND2_X1 U10948 ( .A1(n8781), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n8611) );
  AND2_X1 U10949 ( .A1(n8612), .A2(n8611), .ZN(n8614) );
  INV_X1 U10950 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n11828) );
  OR2_X1 U10951 ( .A1(n8804), .A2(n11828), .ZN(n8613) );
  OAI211_X1 U10952 ( .C1(n14222), .C2(n8667), .A(n8614), .B(n8613), .ZN(n14238) );
  INV_X1 U10953 ( .A(n14238), .ZN(n14095) );
  AND2_X1 U10954 ( .A1(n8615), .A2(n8960), .ZN(n8970) );
  INV_X1 U10955 ( .A(n8960), .ZN(n8616) );
  NAND2_X1 U10956 ( .A1(n14634), .A2(n14095), .ZN(n8972) );
  NAND2_X1 U10957 ( .A1(n14639), .A2(n14223), .ZN(n11816) );
  AND2_X1 U10958 ( .A1(n11821), .A2(n11816), .ZN(n11817) );
  XNOR2_X1 U10959 ( .A(n8619), .B(n8618), .ZN(n11583) );
  NAND2_X1 U10960 ( .A1(n11583), .A2(n6617), .ZN(n8625) );
  OR3_X1 U10961 ( .A1(n8796), .A2(P1_IR_REG_15__SCAN_IN), .A3(
        P1_IR_REG_14__SCAN_IN), .ZN(n8622) );
  NAND2_X1 U10962 ( .A1(n8622), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8620) );
  MUX2_X1 U10963 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8620), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n8621) );
  INV_X1 U10964 ( .A(n8621), .ZN(n8623) );
  NOR2_X1 U10965 ( .A1(n8622), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n8633) );
  NOR2_X1 U10966 ( .A1(n8623), .A2(n8633), .ZN(n14297) );
  AOI22_X1 U10967 ( .A1(n9079), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n8661), 
        .B2(n14297), .ZN(n8624) );
  NOR2_X1 U10968 ( .A1(n8626), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8627) );
  OR2_X1 U10969 ( .A1(n8637), .A2(n8627), .ZN(n14151) );
  AOI22_X1 U10970 ( .A1(n9064), .A2(P1_REG0_REG_16__SCAN_IN), .B1(n8781), .B2(
        P1_REG1_REG_16__SCAN_IN), .ZN(n8629) );
  NAND2_X1 U10971 ( .A1(n9063), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8628) );
  OAI211_X1 U10972 ( .C1(n14151), .C2(n8667), .A(n8629), .B(n8628), .ZN(n14538) );
  INV_X1 U10973 ( .A(n14538), .ZN(n14224) );
  XNOR2_X1 U10974 ( .A(n14153), .B(n14224), .ZN(n11887) );
  NAND2_X1 U10975 ( .A1(n14153), .A2(n14224), .ZN(n8630) );
  NAND2_X1 U10976 ( .A1(n11891), .A2(n8630), .ZN(n14536) );
  XNOR2_X1 U10977 ( .A(n8632), .B(n8631), .ZN(n11739) );
  NAND2_X1 U10978 ( .A1(n11739), .A2(n6617), .ZN(n8636) );
  INV_X1 U10979 ( .A(n8633), .ZN(n8644) );
  NAND2_X1 U10980 ( .A1(n8644), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8634) );
  XNOR2_X1 U10981 ( .A(n8634), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14310) );
  AOI22_X1 U10982 ( .A1(n9079), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n8661), 
        .B2(n14310), .ZN(n8635) );
  OR2_X1 U10983 ( .A1(n8637), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8638) );
  NAND2_X1 U10984 ( .A1(n8665), .A2(n8638), .ZN(n14547) );
  AOI22_X1 U10985 ( .A1(n9064), .A2(P1_REG0_REG_17__SCAN_IN), .B1(n8781), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n8640) );
  NAND2_X1 U10986 ( .A1(n9063), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8639) );
  OAI211_X1 U10987 ( .C1(n14547), .C2(n8667), .A(n8640), .B(n8639), .ZN(n14517) );
  XNOR2_X1 U10988 ( .A(n14550), .B(n14517), .ZN(n14537) );
  INV_X1 U10989 ( .A(n14517), .ZN(n14203) );
  AND2_X1 U10990 ( .A1(n14550), .A2(n14203), .ZN(n8641) );
  XNOR2_X1 U10991 ( .A(n8643), .B(n8642), .ZN(n11867) );
  NAND2_X1 U10992 ( .A1(n11867), .A2(n6617), .ZN(n8647) );
  OAI21_X1 U10993 ( .B1(n8644), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8645) );
  XNOR2_X1 U10994 ( .A(n8645), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14308) );
  AOI22_X1 U10995 ( .A1(n8541), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n14308), 
        .B2(n8661), .ZN(n8646) );
  XNOR2_X1 U10996 ( .A(n8665), .B(P1_REG3_REG_18__SCAN_IN), .ZN(n14525) );
  NAND2_X1 U10997 ( .A1(n14525), .A2(n8785), .ZN(n8653) );
  INV_X1 U10998 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n8650) );
  NAND2_X1 U10999 ( .A1(n9063), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8649) );
  NAND2_X1 U11000 ( .A1(n8781), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8648) );
  OAI211_X1 U11001 ( .C1(n8803), .C2(n8650), .A(n8649), .B(n8648), .ZN(n8651)
         );
  INV_X1 U11002 ( .A(n8651), .ZN(n8652) );
  NAND2_X1 U11003 ( .A1(n8653), .A2(n8652), .ZN(n14541) );
  INV_X1 U11004 ( .A(n14541), .ZN(n8987) );
  NAND2_X1 U11005 ( .A1(n14620), .A2(n8987), .ZN(n8654) );
  NAND2_X1 U11006 ( .A1(n14515), .A2(n14516), .ZN(n14514) );
  XNOR2_X1 U11007 ( .A(n8656), .B(n8655), .ZN(n12732) );
  NAND2_X1 U11008 ( .A1(n12732), .A2(n6617), .ZN(n8663) );
  INV_X1 U11009 ( .A(n8796), .ZN(n8659) );
  INV_X1 U11010 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n13492) );
  INV_X1 U11011 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n13629) );
  INV_X1 U11012 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n8657) );
  NAND2_X1 U11013 ( .A1(n8659), .A2(n7581), .ZN(n8660) );
  INV_X1 U11014 ( .A(n14334), .ZN(n14552) );
  AOI22_X1 U11015 ( .A1(n8541), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14552), 
        .B2(n8661), .ZN(n8662) );
  INV_X1 U11016 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n14201) );
  INV_X1 U11017 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8664) );
  OAI21_X1 U11018 ( .B1(n8665), .B2(n14201), .A(n8664), .ZN(n8666) );
  NAND2_X1 U11019 ( .A1(n8666), .A2(n8677), .ZN(n14499) );
  OR2_X1 U11020 ( .A1(n14499), .A2(n8667), .ZN(n8672) );
  INV_X1 U11021 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14322) );
  NAND2_X1 U11022 ( .A1(n9064), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8669) );
  NAND2_X1 U11023 ( .A1(n9063), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n8668) );
  OAI211_X1 U11024 ( .C1(n8706), .C2(n14322), .A(n8669), .B(n8668), .ZN(n8670)
         );
  INV_X1 U11025 ( .A(n8670), .ZN(n8671) );
  NAND2_X1 U11026 ( .A1(n8672), .A2(n8671), .ZN(n14518) );
  INV_X1 U11027 ( .A(n14518), .ZN(n14202) );
  XNOR2_X1 U11028 ( .A(n14616), .B(n14202), .ZN(n14495) );
  NAND2_X1 U11029 ( .A1(n14616), .A2(n14202), .ZN(n8673) );
  XNOR2_X1 U11030 ( .A(n8686), .B(SI_20_), .ZN(n8685) );
  XNOR2_X1 U11031 ( .A(n8685), .B(n8674), .ZN(n12741) );
  NAND2_X1 U11032 ( .A1(n12741), .A2(n6617), .ZN(n8676) );
  NAND2_X1 U11033 ( .A1(n9079), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8675) );
  NAND2_X1 U11034 ( .A1(n8677), .A2(n14180), .ZN(n8678) );
  NAND2_X1 U11035 ( .A1(n8694), .A2(n8678), .ZN(n14177) );
  INV_X1 U11036 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n8681) );
  NAND2_X1 U11037 ( .A1(n9063), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8680) );
  NAND2_X1 U11038 ( .A1(n8781), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n8679) );
  OAI211_X1 U11039 ( .C1(n8803), .C2(n8681), .A(n8680), .B(n8679), .ZN(n8682)
         );
  INV_X1 U11040 ( .A(n8682), .ZN(n8683) );
  OAI21_X1 U11041 ( .B1(n14177), .B2(n8667), .A(n8683), .ZN(n14496) );
  INV_X1 U11042 ( .A(n14496), .ZN(n14134) );
  XNOR2_X1 U11043 ( .A(n14609), .B(n14134), .ZN(n9111) );
  NAND2_X1 U11044 ( .A1(n8685), .A2(n8684), .ZN(n8688) );
  OR2_X1 U11045 ( .A1(n8686), .A2(n10505), .ZN(n8687) );
  XNOR2_X1 U11046 ( .A(n8689), .B(SI_21_), .ZN(n8690) );
  NAND2_X1 U11047 ( .A1(n12760), .A2(n6617), .ZN(n8693) );
  NAND2_X1 U11048 ( .A1(n9079), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8692) );
  AND2_X1 U11049 ( .A1(n8694), .A2(n14132), .ZN(n8695) );
  OR2_X1 U11050 ( .A1(n8695), .A2(n8702), .ZN(n14133) );
  INV_X1 U11051 ( .A(n14133), .ZN(n14468) );
  INV_X1 U11052 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n13674) );
  NAND2_X1 U11053 ( .A1(n9063), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8697) );
  NAND2_X1 U11054 ( .A1(n8781), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n8696) );
  OAI211_X1 U11055 ( .C1(n8803), .C2(n13674), .A(n8697), .B(n8696), .ZN(n8698)
         );
  AOI21_X1 U11056 ( .B1(n14468), .B2(n8785), .A(n8698), .ZN(n14439) );
  INV_X1 U11057 ( .A(n14439), .ZN(n14237) );
  NAND2_X1 U11058 ( .A1(n14460), .A2(n14237), .ZN(n8699) );
  NAND2_X1 U11059 ( .A1(n11941), .A2(n9486), .ZN(n8701) );
  OR2_X1 U11060 ( .A1(n8702), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8703) );
  AND2_X1 U11061 ( .A1(n8703), .A2(n8719), .ZN(n14437) );
  INV_X1 U11062 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n13552) );
  NAND2_X1 U11063 ( .A1(n9064), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8705) );
  NAND2_X1 U11064 ( .A1(n9063), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8704) );
  OAI211_X1 U11065 ( .C1(n8706), .C2(n13552), .A(n8705), .B(n8704), .ZN(n8707)
         );
  AOI21_X1 U11066 ( .B1(n14437), .B2(n8785), .A(n8707), .ZN(n14467) );
  INV_X1 U11067 ( .A(n14467), .ZN(n14236) );
  XNOR2_X1 U11068 ( .A(n14445), .B(n14236), .ZN(n14448) );
  OR2_X1 U11069 ( .A1(n14445), .A2(n14236), .ZN(n8708) );
  NAND2_X1 U11070 ( .A1(n11941), .A2(n8709), .ZN(n8712) );
  NAND2_X1 U11071 ( .A1(n8710), .A2(SI_22_), .ZN(n8711) );
  XNOR2_X1 U11072 ( .A(n8713), .B(SI_23_), .ZN(n8714) );
  NAND2_X1 U11073 ( .A1(n12783), .A2(n6617), .ZN(n8717) );
  NAND2_X1 U11074 ( .A1(n8541), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8716) );
  NAND2_X1 U11075 ( .A1(n9064), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8723) );
  NAND2_X1 U11076 ( .A1(n8781), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n8722) );
  INV_X1 U11077 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n14109) );
  AOI21_X1 U11078 ( .B1(n14109), .B2(n8719), .A(n8718), .ZN(n14424) );
  NAND2_X1 U11079 ( .A1(n6683), .A2(n14424), .ZN(n8721) );
  NAND2_X1 U11080 ( .A1(n9063), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n8720) );
  NAND4_X1 U11081 ( .A1(n8723), .A2(n8722), .A3(n8721), .A4(n8720), .ZN(n14440) );
  XNOR2_X1 U11082 ( .A(n14423), .B(n14440), .ZN(n14427) );
  INV_X1 U11083 ( .A(n14440), .ZN(n14169) );
  NAND2_X1 U11084 ( .A1(n14423), .A2(n14169), .ZN(n8724) );
  NAND2_X1 U11085 ( .A1(n8725), .A2(n8724), .ZN(n14401) );
  INV_X1 U11086 ( .A(n14401), .ZN(n8727) );
  INV_X1 U11087 ( .A(n14406), .ZN(n8726) );
  OAI21_X1 U11088 ( .B1(n8728), .B2(n14585), .A(n14403), .ZN(n14388) );
  INV_X1 U11089 ( .A(n8729), .ZN(n8732) );
  NAND2_X1 U11090 ( .A1(n8730), .A2(SI_24_), .ZN(n8731) );
  MUX2_X1 U11091 ( .A(n11516), .B(n11519), .S(n9794), .Z(n8734) );
  NAND2_X1 U11092 ( .A1(n8734), .A2(n11324), .ZN(n8745) );
  INV_X1 U11093 ( .A(n8734), .ZN(n8735) );
  NAND2_X1 U11094 ( .A1(n8735), .A2(SI_25_), .ZN(n8736) );
  NAND2_X1 U11095 ( .A1(n8745), .A2(n8736), .ZN(n8746) );
  XNOR2_X1 U11096 ( .A(n8747), .B(n8746), .ZN(n12811) );
  NAND2_X1 U11097 ( .A1(n12811), .A2(n6617), .ZN(n8738) );
  NAND2_X1 U11098 ( .A1(n9079), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8737) );
  NAND2_X1 U11099 ( .A1(n8781), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8743) );
  NAND2_X1 U11100 ( .A1(n9063), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8742) );
  OAI21_X1 U11101 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n8739), .A(n8753), .ZN(
        n14144) );
  INV_X1 U11102 ( .A(n14144), .ZN(n14391) );
  NAND2_X1 U11103 ( .A1(n8785), .A2(n14391), .ZN(n8741) );
  NAND2_X1 U11104 ( .A1(n9064), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8740) );
  NAND4_X1 U11105 ( .A1(n8743), .A2(n8742), .A3(n8741), .A4(n8740), .ZN(n14404) );
  XNOR2_X1 U11106 ( .A(n14578), .B(n14210), .ZN(n14389) );
  NAND2_X1 U11107 ( .A1(n14578), .A2(n14210), .ZN(n8744) );
  MUX2_X1 U11108 ( .A(n13524), .B(n11703), .S(n9794), .Z(n8759) );
  XNOR2_X1 U11109 ( .A(n8759), .B(SI_26_), .ZN(n8748) );
  NAND2_X1 U11110 ( .A1(n9079), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8749) );
  NAND2_X1 U11111 ( .A1(n9064), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8758) );
  NAND2_X1 U11112 ( .A1(n8781), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8757) );
  INV_X1 U11113 ( .A(n8753), .ZN(n8751) );
  NAND2_X1 U11114 ( .A1(n8751), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8765) );
  INV_X1 U11115 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8752) );
  NAND2_X1 U11116 ( .A1(n8753), .A2(n8752), .ZN(n8754) );
  NAND2_X1 U11117 ( .A1(n6683), .A2(n14377), .ZN(n8756) );
  NAND2_X1 U11118 ( .A1(n9063), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8755) );
  NAND4_X1 U11119 ( .A1(n8758), .A2(n8757), .A3(n8756), .A4(n8755), .ZN(n14361) );
  INV_X1 U11120 ( .A(n14361), .ZN(n14086) );
  INV_X1 U11121 ( .A(n14572), .ZN(n14379) );
  MUX2_X1 U11122 ( .A(n11833), .B(n11791), .S(n9794), .Z(n8771) );
  XNOR2_X1 U11123 ( .A(n8771), .B(SI_27_), .ZN(n8761) );
  NAND2_X1 U11124 ( .A1(n8541), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8762) );
  NAND2_X1 U11125 ( .A1(n9064), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8770) );
  INV_X1 U11126 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n13687) );
  OR2_X1 U11127 ( .A1(n8804), .A2(n13687), .ZN(n8769) );
  NAND2_X1 U11128 ( .A1(n8781), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n8768) );
  INV_X1 U11129 ( .A(n8765), .ZN(n8764) );
  NAND2_X1 U11130 ( .A1(n8764), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8783) );
  INV_X1 U11131 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n14085) );
  NAND2_X1 U11132 ( .A1(n8765), .A2(n14085), .ZN(n8766) );
  NAND2_X1 U11133 ( .A1(n6683), .A2(n14084), .ZN(n8767) );
  NAND4_X1 U11134 ( .A1(n8770), .A2(n8769), .A3(n8768), .A4(n8767), .ZN(n14234) );
  INV_X1 U11135 ( .A(n14234), .ZN(n14211) );
  INV_X1 U11136 ( .A(n8771), .ZN(n8773) );
  NAND2_X1 U11137 ( .A1(n8773), .A2(SI_27_), .ZN(n8774) );
  NAND2_X1 U11138 ( .A1(n8775), .A2(n8774), .ZN(n9043) );
  MUX2_X1 U11139 ( .A(n12007), .B(n13634), .S(n9794), .Z(n8776) );
  NAND2_X1 U11140 ( .A1(n8776), .A2(n11536), .ZN(n9041) );
  INV_X1 U11141 ( .A(n8776), .ZN(n8777) );
  NAND2_X1 U11142 ( .A1(n8777), .A2(SI_28_), .ZN(n8778) );
  NAND2_X1 U11143 ( .A1(n9041), .A2(n8778), .ZN(n9042) );
  NAND2_X1 U11144 ( .A1(n12891), .A2(n6617), .ZN(n8780) );
  NAND2_X1 U11145 ( .A1(n8541), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8779) );
  NAND2_X1 U11146 ( .A1(n9064), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8789) );
  INV_X1 U11147 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n13727) );
  OR2_X1 U11148 ( .A1(n8804), .A2(n13727), .ZN(n8788) );
  NAND2_X1 U11149 ( .A1(n8781), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n8787) );
  INV_X1 U11150 ( .A(n8783), .ZN(n8782) );
  NAND2_X1 U11151 ( .A1(n8782), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n11978) );
  INV_X1 U11152 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n12127) );
  NAND2_X1 U11153 ( .A1(n8783), .A2(n12127), .ZN(n8784) );
  NAND2_X1 U11154 ( .A1(n6683), .A2(n12126), .ZN(n8786) );
  XNOR2_X1 U11155 ( .A(n11967), .B(n8790), .ZN(n8812) );
  NAND2_X1 U11156 ( .A1(n8792), .A2(n8791), .ZN(n8793) );
  INV_X1 U11157 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8794) );
  NAND2_X1 U11158 ( .A1(n8899), .A2(n14552), .ZN(n8800) );
  NAND2_X1 U11159 ( .A1(n8901), .A2(n8800), .ZN(n14701) );
  NAND2_X1 U11160 ( .A1(n8456), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8808) );
  INV_X1 U11161 ( .A(n11978), .ZN(n8801) );
  NAND2_X1 U11162 ( .A1(n8785), .A2(n8801), .ZN(n8807) );
  INV_X1 U11163 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n8802) );
  OR2_X1 U11164 ( .A1(n8803), .A2(n8802), .ZN(n8806) );
  INV_X1 U11165 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n13675) );
  OR2_X1 U11166 ( .A1(n8804), .A2(n13675), .ZN(n8805) );
  INV_X1 U11167 ( .A(n12129), .ZN(n14233) );
  NAND2_X1 U11168 ( .A1(n14233), .A2(n14540), .ZN(n8810) );
  INV_X1 U11169 ( .A(n12005), .ZN(n14256) );
  NAND2_X1 U11170 ( .A1(n14234), .A2(n14539), .ZN(n8809) );
  NAND2_X1 U11171 ( .A1(n10246), .A2(n14125), .ZN(n8907) );
  NAND2_X1 U11172 ( .A1(n6609), .A2(n11130), .ZN(n11137) );
  NAND2_X1 U11173 ( .A1(n11135), .A2(n10594), .ZN(n8898) );
  INV_X1 U11174 ( .A(n14250), .ZN(n10743) );
  NAND2_X1 U11175 ( .A1(n10743), .A2(n7099), .ZN(n10618) );
  NAND2_X1 U11176 ( .A1(n10829), .A2(n10618), .ZN(n10617) );
  AND2_X1 U11177 ( .A1(n10813), .A2(n10622), .ZN(n8814) );
  NAND2_X1 U11178 ( .A1(n10939), .A2(n10794), .ZN(n10809) );
  OR2_X1 U11179 ( .A1(n10934), .A2(n14248), .ZN(n10781) );
  NAND2_X1 U11180 ( .A1(n10780), .A2(n10781), .ZN(n8815) );
  NAND2_X1 U11181 ( .A1(n8815), .A2(n10777), .ZN(n10784) );
  NAND2_X1 U11182 ( .A1(n10784), .A2(n8816), .ZN(n11016) );
  INV_X1 U11183 ( .A(n11013), .ZN(n11017) );
  NAND2_X1 U11184 ( .A1(n11016), .A2(n11017), .ZN(n11015) );
  OR2_X1 U11185 ( .A1(n14954), .A2(n14246), .ZN(n8817) );
  NAND2_X1 U11186 ( .A1(n11015), .A2(n8817), .ZN(n10973) );
  INV_X1 U11187 ( .A(n10976), .ZN(n10972) );
  NAND2_X1 U11188 ( .A1(n10973), .A2(n10972), .ZN(n10971) );
  OR2_X1 U11189 ( .A1(n14956), .A2(n14245), .ZN(n8818) );
  NAND2_X1 U11190 ( .A1(n10971), .A2(n8818), .ZN(n11108) );
  INV_X1 U11191 ( .A(n11681), .ZN(n14244) );
  OR2_X1 U11192 ( .A1(n11671), .A2(n14244), .ZN(n8819) );
  INV_X1 U11193 ( .A(n9103), .ZN(n11193) );
  OR2_X1 U11194 ( .A1(n14964), .A2(n14243), .ZN(n8820) );
  NAND2_X1 U11195 ( .A1(n14843), .A2(n14242), .ZN(n8821) );
  OR2_X1 U11196 ( .A1(n14843), .A2(n14242), .ZN(n8822) );
  NAND2_X1 U11197 ( .A1(n8823), .A2(n8822), .ZN(n14708) );
  NAND2_X1 U11198 ( .A1(n14708), .A2(n14709), .ZN(n8825) );
  OR2_X1 U11199 ( .A1(n14707), .A2(n14241), .ZN(n8824) );
  NAND2_X1 U11200 ( .A1(n8825), .A2(n8824), .ZN(n11461) );
  NAND2_X1 U11201 ( .A1(n11461), .A2(n11460), .ZN(n8827) );
  OR2_X1 U11202 ( .A1(n11928), .A2(n14240), .ZN(n8826) );
  XNOR2_X1 U11203 ( .A(n14639), .B(n14239), .ZN(n11611) );
  NAND2_X1 U11204 ( .A1(n14639), .A2(n14239), .ZN(n8828) );
  INV_X1 U11205 ( .A(n11814), .ZN(n8830) );
  INV_X1 U11206 ( .A(n11821), .ZN(n8829) );
  NAND2_X1 U11207 ( .A1(n8830), .A2(n8829), .ZN(n11812) );
  OR2_X1 U11208 ( .A1(n14634), .A2(n14238), .ZN(n8831) );
  NAND2_X1 U11209 ( .A1(n11812), .A2(n8831), .ZN(n11885) );
  NAND2_X1 U11210 ( .A1(n11885), .A2(n11887), .ZN(n8833) );
  OR2_X1 U11211 ( .A1(n14153), .A2(n14538), .ZN(n8832) );
  NOR2_X1 U11212 ( .A1(n14550), .A2(n14517), .ZN(n8834) );
  NAND2_X1 U11213 ( .A1(n14550), .A2(n14517), .ZN(n8982) );
  OR2_X1 U11214 ( .A1(n14620), .A2(n14541), .ZN(n14489) );
  OR2_X1 U11215 ( .A1(n14616), .A2(n14518), .ZN(n8835) );
  AND2_X1 U11216 ( .A1(n14489), .A2(n8835), .ZN(n8837) );
  INV_X1 U11217 ( .A(n8835), .ZN(n8836) );
  INV_X1 U11218 ( .A(n9111), .ZN(n14475) );
  NAND2_X1 U11219 ( .A1(n14609), .A2(n14496), .ZN(n14454) );
  NAND2_X1 U11220 ( .A1(n14460), .A2(n14439), .ZN(n8838) );
  NAND2_X1 U11221 ( .A1(n14445), .A2(n14467), .ZN(n8839) );
  OR2_X1 U11222 ( .A1(n14423), .A2(n14440), .ZN(n8840) );
  NAND2_X1 U11223 ( .A1(n8841), .A2(n8840), .ZN(n14405) );
  OR2_X1 U11224 ( .A1(n14585), .A2(n14235), .ZN(n8842) );
  INV_X1 U11225 ( .A(n14389), .ZN(n14397) );
  NAND2_X1 U11226 ( .A1(n14578), .A2(n14404), .ZN(n8843) );
  NAND2_X1 U11227 ( .A1(n14572), .A2(n14361), .ZN(n8844) );
  OR2_X1 U11228 ( .A1(n14567), .A2(n14234), .ZN(n8846) );
  NAND2_X1 U11229 ( .A1(n10084), .A2(n8899), .ZN(n8849) );
  NAND2_X1 U11230 ( .A1(n8899), .A2(n14334), .ZN(n8848) );
  NAND2_X1 U11231 ( .A1(n10083), .A2(n8848), .ZN(n10932) );
  NAND2_X1 U11232 ( .A1(n9822), .A2(n7223), .ZN(n14546) );
  NAND2_X1 U11233 ( .A1(n9822), .A2(n14552), .ZN(n8851) );
  INV_X1 U11234 ( .A(n10934), .ZN(n14948) );
  INV_X1 U11235 ( .A(n10964), .ZN(n11041) );
  INV_X1 U11236 ( .A(n11671), .ZN(n14897) );
  INV_X1 U11237 ( .A(n14843), .ZN(n8852) );
  INV_X1 U11238 ( .A(n11928), .ZN(n14860) );
  INV_X1 U11239 ( .A(n14634), .ZN(n14231) );
  INV_X1 U11240 ( .A(n14616), .ZN(n14507) );
  NAND2_X1 U11241 ( .A1(n14481), .A2(n14460), .ZN(n14456) );
  INV_X1 U11242 ( .A(n14578), .ZN(n14394) );
  INV_X1 U11243 ( .A(n8854), .ZN(n14376) );
  NOR2_X2 U11244 ( .A1(n14376), .A2(n14567), .ZN(n14354) );
  INV_X1 U11245 ( .A(n14354), .ZN(n8856) );
  INV_X1 U11246 ( .A(n14712), .ZN(n14503) );
  NAND2_X1 U11247 ( .A1(n11998), .A2(n14354), .ZN(n11972) );
  INV_X1 U11248 ( .A(n11972), .ZN(n8855) );
  AOI211_X1 U11249 ( .C1(n12132), .C2(n8856), .A(n14503), .B(n8855), .ZN(
        n12002) );
  AOI21_X1 U11250 ( .B1(n12132), .B2(n14963), .A(n12002), .ZN(n8857) );
  NAND2_X1 U11251 ( .A1(n8859), .A2(n8858), .ZN(n8876) );
  XNOR2_X1 U11252 ( .A(n8861), .B(n8860), .ZN(n8875) );
  INV_X1 U11253 ( .A(n8875), .ZN(n8863) );
  INV_X1 U11254 ( .A(P1_B_REG_SCAN_IN), .ZN(n8862) );
  NAND2_X1 U11255 ( .A1(n8863), .A2(n8862), .ZN(n8873) );
  OAI21_X1 U11256 ( .B1(n8796), .B2(n8864), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n8865) );
  MUX2_X1 U11257 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8865), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n8867) );
  NAND2_X1 U11258 ( .A1(n8867), .A2(n8868), .ZN(n11515) );
  NAND3_X1 U11259 ( .A1(n8875), .A2(P1_B_REG_SCAN_IN), .A3(n11515), .ZN(n8872)
         );
  NAND2_X1 U11260 ( .A1(n8868), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8869) );
  MUX2_X1 U11261 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8869), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n8871) );
  NAND3_X1 U11262 ( .A1(n8873), .A2(n8872), .A3(n8874), .ZN(n10078) );
  NAND2_X1 U11263 ( .A1(n11515), .A2(n11726), .ZN(n10079) );
  OAI21_X1 U11264 ( .B1(n10078), .B2(P1_D_REG_1__SCAN_IN), .A(n10079), .ZN(
        n8894) );
  NAND2_X1 U11265 ( .A1(n8876), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8878) );
  XNOR2_X1 U11266 ( .A(n8878), .B(n8877), .ZN(n10366) );
  NAND2_X1 U11267 ( .A1(n10367), .A2(n9591), .ZN(n10081) );
  AND2_X1 U11268 ( .A1(n8900), .A2(n14552), .ZN(n10220) );
  NAND2_X1 U11269 ( .A1(n10220), .A2(n9822), .ZN(n10369) );
  NAND2_X1 U11270 ( .A1(n8900), .A2(n14334), .ZN(n8879) );
  NAND2_X1 U11271 ( .A1(n10092), .A2(n8879), .ZN(n10365) );
  NAND2_X1 U11272 ( .A1(n10369), .A2(n10365), .ZN(n8880) );
  NOR2_X1 U11273 ( .A1(n10081), .A2(n8880), .ZN(n8893) );
  NOR4_X1 U11274 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n8884) );
  NOR4_X1 U11275 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n8883) );
  NOR4_X1 U11276 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n8882) );
  NOR4_X1 U11277 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n8881) );
  AND4_X1 U11278 ( .A1(n8884), .A2(n8883), .A3(n8882), .A4(n8881), .ZN(n8890)
         );
  NOR2_X1 U11279 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .ZN(
        n8888) );
  NOR4_X1 U11280 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n8887) );
  NOR4_X1 U11281 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n8886) );
  NOR4_X1 U11282 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n8885) );
  AND4_X1 U11283 ( .A1(n8888), .A2(n8887), .A3(n8886), .A4(n8885), .ZN(n8889)
         );
  NAND2_X1 U11284 ( .A1(n8890), .A2(n8889), .ZN(n10076) );
  INV_X1 U11285 ( .A(n10076), .ZN(n8891) );
  OR2_X1 U11286 ( .A1(n10078), .A2(n8891), .ZN(n8892) );
  AND3_X1 U11287 ( .A1(n8894), .A2(n8893), .A3(n8892), .ZN(n9825) );
  OR2_X1 U11288 ( .A1(n10078), .A2(P1_D_REG_0__SCAN_IN), .ZN(n8895) );
  NAND2_X1 U11289 ( .A1(n8875), .A2(n11726), .ZN(n9663) );
  NAND2_X1 U11290 ( .A1(n8895), .A2(n9663), .ZN(n10364) );
  AND2_X2 U11291 ( .A1(n9825), .A2(n10364), .ZN(n14973) );
  NAND2_X1 U11292 ( .A1(n14971), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8896) );
  INV_X1 U11293 ( .A(n8898), .ZN(n8914) );
  OAI21_X1 U11294 ( .B1(n11130), .B2(n10083), .A(n8903), .ZN(n8902) );
  NAND2_X1 U11295 ( .A1(n6609), .A2(n8902), .ZN(n8906) );
  INV_X1 U11296 ( .A(n8903), .ZN(n8904) );
  NAND2_X1 U11297 ( .A1(n10098), .A2(n8904), .ZN(n8905) );
  NOR2_X1 U11298 ( .A1(n6612), .A2(n14125), .ZN(n8909) );
  NAND2_X1 U11299 ( .A1(n8912), .A2(n8911), .ZN(n8913) );
  OAI21_X1 U11300 ( .B1(n10594), .B2(n11135), .A(n8915), .ZN(n8916) );
  NAND2_X1 U11301 ( .A1(n8917), .A2(n10822), .ZN(n8922) );
  MUX2_X1 U11302 ( .A(n8920), .B(n8919), .S(n9082), .Z(n8921) );
  MUX2_X1 U11303 ( .A(n10939), .B(n10794), .S(n9082), .Z(n8924) );
  MUX2_X1 U11304 ( .A(n14249), .B(n10746), .S(n6612), .Z(n8923) );
  MUX2_X1 U11305 ( .A(n14248), .B(n10934), .S(n6612), .Z(n8926) );
  MUX2_X1 U11306 ( .A(n10934), .B(n14248), .S(n6612), .Z(n8925) );
  INV_X1 U11307 ( .A(n8926), .ZN(n8927) );
  MUX2_X1 U11308 ( .A(n14247), .B(n10964), .S(n9082), .Z(n8931) );
  MUX2_X1 U11309 ( .A(n14247), .B(n10964), .S(n6612), .Z(n8928) );
  NAND2_X1 U11310 ( .A1(n8929), .A2(n8928), .ZN(n8935) );
  INV_X1 U11311 ( .A(n8930), .ZN(n8933) );
  INV_X1 U11312 ( .A(n8931), .ZN(n8932) );
  MUX2_X1 U11313 ( .A(n14246), .B(n14954), .S(n6612), .Z(n8937) );
  MUX2_X1 U11314 ( .A(n14246), .B(n14954), .S(n9082), .Z(n8936) );
  INV_X1 U11315 ( .A(n8937), .ZN(n8938) );
  MUX2_X1 U11316 ( .A(n14245), .B(n14956), .S(n9082), .Z(n8941) );
  MUX2_X1 U11317 ( .A(n14245), .B(n14956), .S(n6612), .Z(n8939) );
  MUX2_X1 U11318 ( .A(n14244), .B(n11671), .S(n6612), .Z(n8943) );
  MUX2_X1 U11319 ( .A(n14244), .B(n11671), .S(n9082), .Z(n8942) );
  INV_X1 U11320 ( .A(n8943), .ZN(n8944) );
  INV_X1 U11321 ( .A(n14964), .ZN(n11687) );
  MUX2_X1 U11322 ( .A(n14898), .B(n11687), .S(n9026), .Z(n8946) );
  MUX2_X1 U11323 ( .A(n14243), .B(n14964), .S(n9082), .Z(n8945) );
  AOI21_X1 U11324 ( .B1(n8947), .B2(n8946), .A(n8945), .ZN(n8951) );
  NOR2_X1 U11325 ( .A1(n8947), .A2(n8946), .ZN(n8950) );
  INV_X1 U11326 ( .A(n8948), .ZN(n8952) );
  OR2_X1 U11327 ( .A1(n8953), .A2(n8952), .ZN(n11389) );
  INV_X1 U11328 ( .A(n11389), .ZN(n8949) );
  MUX2_X1 U11329 ( .A(n8953), .B(n8952), .S(n6612), .Z(n8954) );
  INV_X1 U11330 ( .A(n14707), .ZN(n14721) );
  MUX2_X1 U11331 ( .A(n11912), .B(n14721), .S(n9082), .Z(n8958) );
  MUX2_X1 U11332 ( .A(n14241), .B(n14707), .S(n9026), .Z(n8957) );
  MUX2_X1 U11333 ( .A(n14240), .B(n11928), .S(n9026), .Z(n8959) );
  NAND3_X1 U11334 ( .A1(n8960), .A2(n11611), .A3(n7227), .ZN(n8966) );
  AND4_X1 U11335 ( .A1(n8960), .A2(n11611), .A3(n11928), .A4(n9082), .ZN(n8961) );
  NAND2_X1 U11336 ( .A1(n8969), .A2(n8961), .ZN(n8965) );
  OAI21_X1 U11337 ( .B1(n14238), .B2(n11816), .A(n14231), .ZN(n8963) );
  AOI21_X1 U11338 ( .B1(n11816), .B2(n14238), .A(n9026), .ZN(n8962) );
  NAND2_X1 U11339 ( .A1(n8963), .A2(n8962), .ZN(n8964) );
  OAI211_X1 U11340 ( .C1(n8967), .C2(n8966), .A(n8965), .B(n8964), .ZN(n8977)
         );
  INV_X1 U11341 ( .A(n8972), .ZN(n8973) );
  INV_X1 U11342 ( .A(n14153), .ZN(n14628) );
  MUX2_X1 U11343 ( .A(n14224), .B(n14628), .S(n9082), .Z(n8979) );
  MUX2_X1 U11344 ( .A(n14538), .B(n14153), .S(n9026), .Z(n8978) );
  AOI22_X1 U11345 ( .A1(n8973), .A2(n9026), .B1(n8979), .B2(n8978), .ZN(n8974)
         );
  OAI21_X1 U11346 ( .B1(n8977), .B2(n8976), .A(n8975), .ZN(n8986) );
  INV_X1 U11347 ( .A(n8978), .ZN(n8981) );
  INV_X1 U11348 ( .A(n8979), .ZN(n8980) );
  NAND3_X1 U11349 ( .A1(n14537), .A2(n8981), .A3(n8980), .ZN(n8985) );
  MUX2_X1 U11350 ( .A(n14517), .B(n14550), .S(n9082), .Z(n8983) );
  NAND2_X1 U11351 ( .A1(n8983), .A2(n8982), .ZN(n8984) );
  NAND3_X1 U11352 ( .A1(n8986), .A2(n8985), .A3(n8984), .ZN(n8990) );
  INV_X1 U11353 ( .A(n14495), .ZN(n8997) );
  MUX2_X1 U11354 ( .A(n9082), .B(n14620), .S(n8987), .Z(n8988) );
  NAND2_X1 U11355 ( .A1(n14620), .A2(n9082), .ZN(n8991) );
  NAND2_X1 U11356 ( .A1(n8988), .A2(n8991), .ZN(n8989) );
  OAI22_X1 U11357 ( .A1(n8992), .A2(n9082), .B1(n8991), .B2(n14541), .ZN(n8996) );
  NOR2_X1 U11358 ( .A1(n14616), .A2(n9082), .ZN(n8994) );
  AND2_X1 U11359 ( .A1(n14616), .A2(n9082), .ZN(n8993) );
  MUX2_X1 U11360 ( .A(n8994), .B(n8993), .S(n14202), .Z(n8995) );
  AOI21_X1 U11361 ( .B1(n8997), .B2(n8996), .A(n8995), .ZN(n8998) );
  INV_X1 U11362 ( .A(n14609), .ZN(n14484) );
  MUX2_X1 U11363 ( .A(n14134), .B(n14484), .S(n9026), .Z(n9000) );
  MUX2_X1 U11364 ( .A(n14496), .B(n14609), .S(n9082), .Z(n8999) );
  MUX2_X1 U11365 ( .A(n14237), .B(n6970), .S(n9082), .Z(n9002) );
  MUX2_X1 U11366 ( .A(n14439), .B(n14460), .S(n9026), .Z(n9001) );
  INV_X1 U11367 ( .A(n9008), .ZN(n9006) );
  MUX2_X1 U11368 ( .A(n14236), .B(n14599), .S(n9026), .Z(n9007) );
  INV_X1 U11369 ( .A(n9007), .ZN(n9005) );
  MUX2_X1 U11370 ( .A(n14236), .B(n14599), .S(n9082), .Z(n9009) );
  NAND2_X1 U11371 ( .A1(n9010), .A2(n9009), .ZN(n9011) );
  MUX2_X1 U11372 ( .A(n14440), .B(n14423), .S(n9082), .Z(n9014) );
  MUX2_X1 U11373 ( .A(n14440), .B(n14423), .S(n9026), .Z(n9013) );
  INV_X1 U11374 ( .A(n9014), .ZN(n9015) );
  MUX2_X1 U11375 ( .A(n14235), .B(n14585), .S(n9026), .Z(n9019) );
  NAND2_X1 U11376 ( .A1(n9018), .A2(n9019), .ZN(n9017) );
  MUX2_X1 U11377 ( .A(n14235), .B(n14585), .S(n9082), .Z(n9016) );
  NAND2_X1 U11378 ( .A1(n9017), .A2(n9016), .ZN(n9023) );
  INV_X1 U11379 ( .A(n9019), .ZN(n9020) );
  NAND2_X1 U11380 ( .A1(n9021), .A2(n9020), .ZN(n9022) );
  MUX2_X1 U11381 ( .A(n14404), .B(n14578), .S(n9082), .Z(n9025) );
  MUX2_X1 U11382 ( .A(n14404), .B(n14578), .S(n9026), .Z(n9024) );
  MUX2_X1 U11383 ( .A(n14361), .B(n14572), .S(n9026), .Z(n9028) );
  INV_X1 U11384 ( .A(n9028), .ZN(n9027) );
  MUX2_X1 U11385 ( .A(n14361), .B(n14572), .S(n9082), .Z(n9029) );
  MUX2_X1 U11386 ( .A(n14234), .B(n14567), .S(n9082), .Z(n9032) );
  MUX2_X1 U11387 ( .A(n14234), .B(n14567), .S(n9026), .Z(n9030) );
  MUX2_X1 U11388 ( .A(n14362), .B(n12132), .S(n9026), .Z(n9036) );
  MUX2_X1 U11389 ( .A(n14362), .B(n12132), .S(n9082), .Z(n9033) );
  NAND2_X1 U11390 ( .A1(n9034), .A2(n9033), .ZN(n9040) );
  INV_X1 U11391 ( .A(n9035), .ZN(n9038) );
  INV_X1 U11392 ( .A(n9036), .ZN(n9037) );
  NAND2_X1 U11393 ( .A1(n9038), .A2(n9037), .ZN(n9039) );
  INV_X1 U11394 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n11988) );
  MUX2_X1 U11395 ( .A(n14670), .B(n11988), .S(n9794), .Z(n9049) );
  XNOR2_X1 U11396 ( .A(n9049), .B(SI_29_), .ZN(n9051) );
  NAND2_X1 U11397 ( .A1(n13157), .A2(n6617), .ZN(n9045) );
  NAND2_X1 U11398 ( .A1(n9079), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n9044) );
  MUX2_X1 U11399 ( .A(n14561), .B(n14233), .S(n9026), .Z(n9048) );
  MUX2_X1 U11400 ( .A(n14233), .B(n14561), .S(n9026), .Z(n9046) );
  INV_X1 U11401 ( .A(n9049), .ZN(n9050) );
  MUX2_X1 U11402 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n9794), .Z(n9053) );
  NAND2_X1 U11403 ( .A1(n9053), .A2(SI_30_), .ZN(n9074) );
  OAI21_X1 U11404 ( .B1(n9053), .B2(SI_30_), .A(n9074), .ZN(n9055) );
  INV_X1 U11405 ( .A(n9055), .ZN(n9054) );
  NAND2_X1 U11406 ( .A1(n7121), .A2(n9055), .ZN(n9056) );
  NAND2_X1 U11407 ( .A1(n9075), .A2(n9056), .ZN(n13165) );
  OR2_X1 U11408 ( .A1(n13165), .A2(n9057), .ZN(n9059) );
  NAND2_X1 U11409 ( .A1(n8541), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n9058) );
  NAND2_X1 U11410 ( .A1(n8781), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n9062) );
  NAND2_X1 U11411 ( .A1(n9063), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n9061) );
  NAND2_X1 U11412 ( .A1(n9064), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n9060) );
  NAND3_X1 U11413 ( .A1(n9062), .A2(n9061), .A3(n9060), .ZN(n14341) );
  NAND2_X1 U11414 ( .A1(n8456), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n9067) );
  NAND2_X1 U11415 ( .A1(n9063), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9066) );
  NAND2_X1 U11416 ( .A1(n9064), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n9065) );
  NAND3_X1 U11417 ( .A1(n9067), .A2(n9066), .A3(n9065), .ZN(n14232) );
  OAI21_X1 U11418 ( .B1(n14341), .B2(n8900), .A(n14232), .ZN(n9068) );
  INV_X1 U11419 ( .A(n9068), .ZN(n9069) );
  MUX2_X1 U11420 ( .A(n14345), .B(n9069), .S(n9026), .Z(n9092) );
  NAND2_X1 U11421 ( .A1(n9070), .A2(n11277), .ZN(n9072) );
  NAND2_X1 U11422 ( .A1(n9082), .A2(n14341), .ZN(n9083) );
  INV_X1 U11423 ( .A(n14232), .ZN(n9071) );
  AOI21_X1 U11424 ( .B1(n9072), .B2(n9083), .A(n9071), .ZN(n9073) );
  AOI21_X1 U11425 ( .B1(n14345), .B2(n9026), .A(n9073), .ZN(n9091) );
  NOR2_X1 U11426 ( .A1(n9092), .A2(n9091), .ZN(n9120) );
  MUX2_X1 U11427 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9794), .Z(n9076) );
  XNOR2_X1 U11428 ( .A(n9076), .B(SI_31_), .ZN(n9077) );
  NAND2_X1 U11429 ( .A1(n14068), .A2(n6617), .ZN(n9081) );
  NAND2_X1 U11430 ( .A1(n9079), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n9080) );
  MUX2_X1 U11431 ( .A(n14341), .B(n9082), .S(n14342), .Z(n9084) );
  NAND2_X1 U11432 ( .A1(n9084), .A2(n9083), .ZN(n9129) );
  INV_X1 U11433 ( .A(n10092), .ZN(n9086) );
  NAND2_X1 U11434 ( .A1(n8850), .A2(n8900), .ZN(n9085) );
  NAND2_X1 U11435 ( .A1(n9086), .A2(n9085), .ZN(n9088) );
  NAND2_X1 U11436 ( .A1(n10220), .A2(n9089), .ZN(n9087) );
  NAND2_X1 U11437 ( .A1(n9088), .A2(n9087), .ZN(n9090) );
  OR2_X1 U11438 ( .A1(n8900), .A2(n9089), .ZN(n9119) );
  AND2_X1 U11439 ( .A1(n9090), .A2(n9119), .ZN(n9127) );
  NAND2_X1 U11440 ( .A1(n9129), .A2(n9127), .ZN(n9125) );
  XNOR2_X1 U11441 ( .A(n14342), .B(n14341), .ZN(n9126) );
  INV_X1 U11442 ( .A(n9090), .ZN(n9131) );
  NAND2_X1 U11443 ( .A1(n9092), .A2(n9091), .ZN(n9124) );
  NAND3_X1 U11444 ( .A1(n9093), .A2(n9121), .A3(n9124), .ZN(n9137) );
  INV_X1 U11445 ( .A(n14516), .ZN(n14512) );
  NAND2_X1 U11446 ( .A1(n6609), .A2(n10098), .ZN(n9095) );
  NAND2_X1 U11447 ( .A1(n9096), .A2(n9095), .ZN(n9820) );
  INV_X1 U11448 ( .A(n9820), .ZN(n9098) );
  NAND4_X1 U11449 ( .A1(n9099), .A2(n10822), .A3(n9098), .A4(n9097), .ZN(n9100) );
  NOR2_X1 U11450 ( .A1(n9100), .A2(n10622), .ZN(n9101) );
  INV_X1 U11451 ( .A(n10777), .ZN(n10782) );
  NAND4_X1 U11452 ( .A1(n11013), .A2(n9101), .A3(n10782), .A4(n7506), .ZN(
        n9102) );
  OR3_X1 U11453 ( .A1(n11109), .A2(n10972), .A3(n9102), .ZN(n9106) );
  NAND2_X1 U11454 ( .A1(n9104), .A2(n9103), .ZN(n9105) );
  OR4_X1 U11455 ( .A1(n11389), .A2(n9106), .A3(n14709), .A4(n9105), .ZN(n9107)
         );
  NOR2_X1 U11456 ( .A1(n11887), .A2(n9107), .ZN(n9108) );
  NAND4_X1 U11457 ( .A1(n11821), .A2(n9108), .A3(n14537), .A4(n11611), .ZN(
        n9109) );
  OR3_X1 U11458 ( .A1(n14512), .A2(n14495), .A3(n9109), .ZN(n9110) );
  NOR2_X1 U11459 ( .A1(n9111), .A2(n9110), .ZN(n9112) );
  NAND4_X1 U11460 ( .A1(n14427), .A2(n7277), .A3(n9112), .A4(n14462), .ZN(
        n9113) );
  OR3_X1 U11461 ( .A1(n14389), .A2(n14406), .A3(n9113), .ZN(n9114) );
  NOR4_X1 U11462 ( .A1(n8790), .A2(n8845), .A3(n14381), .A4(n9114), .ZN(n9117)
         );
  INV_X1 U11463 ( .A(n11970), .ZN(n9116) );
  XNOR2_X1 U11464 ( .A(n14345), .B(n14232), .ZN(n9115) );
  NAND4_X1 U11465 ( .A1(n9126), .A2(n9117), .A3(n9116), .A4(n9115), .ZN(n9118)
         );
  XNOR2_X1 U11466 ( .A(n9118), .B(n14552), .ZN(n9135) );
  INV_X1 U11467 ( .A(n9119), .ZN(n9134) );
  INV_X1 U11468 ( .A(n9120), .ZN(n9123) );
  INV_X1 U11469 ( .A(n9121), .ZN(n9122) );
  OAI22_X1 U11470 ( .A1(n9125), .A2(n9124), .B1(n9123), .B2(n9122), .ZN(n9133)
         );
  INV_X1 U11471 ( .A(n9126), .ZN(n9128) );
  AND2_X1 U11472 ( .A1(n9128), .A2(n9127), .ZN(n9130) );
  MUX2_X1 U11473 ( .A(n9131), .B(n9130), .S(n9129), .Z(n9132) );
  AOI211_X1 U11474 ( .C1(n9135), .C2(n9134), .A(n9133), .B(n9132), .ZN(n9136)
         );
  NAND3_X1 U11475 ( .A1(n9138), .A2(n9137), .A3(n9136), .ZN(n9140) );
  OR2_X1 U11476 ( .A1(n10366), .A2(P1_U3086), .ZN(n11401) );
  NAND2_X1 U11477 ( .A1(n9140), .A2(n9139), .ZN(n9144) );
  INV_X1 U11478 ( .A(n14539), .ZN(n14438) );
  INV_X1 U11479 ( .A(n10365), .ZN(n10082) );
  NOR4_X1 U11480 ( .A1(n10081), .A2(n14438), .A3(n10082), .A4(n6684), .ZN(
        n9142) );
  OAI21_X1 U11481 ( .B1(n11401), .B2(n8899), .A(P1_B_REG_SCAN_IN), .ZN(n9141)
         );
  OR2_X1 U11482 ( .A1(n9142), .A2(n9141), .ZN(n9143) );
  NAND2_X1 U11483 ( .A1(n9144), .A2(n9143), .ZN(P1_U3242) );
  NAND2_X1 U11484 ( .A1(n11952), .A2(n9145), .ZN(n9146) );
  NAND2_X1 U11485 ( .A1(n9146), .A2(n10504), .ZN(n9156) );
  XNOR2_X1 U11486 ( .A(n9147), .B(P3_B_REG_SCAN_IN), .ZN(n9149) );
  NAND2_X1 U11487 ( .A1(n9149), .A2(n9148), .ZN(n9150) );
  INV_X1 U11488 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n9151) );
  OR2_X1 U11489 ( .A1(n9232), .A2(n11218), .ZN(n9152) );
  NAND2_X1 U11490 ( .A1(n9154), .A2(n12715), .ZN(n9155) );
  NAND2_X2 U11491 ( .A1(n9155), .A2(n9156), .ZN(n9165) );
  CLKBUF_X3 U11492 ( .A(n9165), .Z(n10209) );
  XNOR2_X1 U11493 ( .A(n11570), .B(n10209), .ZN(n9201) );
  INV_X1 U11494 ( .A(n9165), .ZN(n9161) );
  NAND2_X1 U11495 ( .A1(n10432), .A2(n9161), .ZN(n9159) );
  NAND2_X1 U11496 ( .A1(n9157), .A2(n9165), .ZN(n9158) );
  NAND2_X1 U11497 ( .A1(n9159), .A2(n9158), .ZN(n9164) );
  NAND3_X1 U11498 ( .A1(n12244), .A2(n9161), .A3(n9160), .ZN(n9162) );
  NAND2_X1 U11500 ( .A1(n15367), .A2(n10187), .ZN(n15368) );
  NAND3_X1 U11501 ( .A1(n10212), .A2(n9163), .A3(n15368), .ZN(n10208) );
  NAND2_X1 U11502 ( .A1(n10208), .A2(n9164), .ZN(n10349) );
  XNOR2_X1 U11503 ( .A(n7649), .B(n9165), .ZN(n9166) );
  XNOR2_X1 U11504 ( .A(n9166), .B(n15365), .ZN(n10350) );
  AND2_X1 U11505 ( .A1(n9166), .A2(n10435), .ZN(n9167) );
  XNOR2_X1 U11506 ( .A(n12243), .B(n9168), .ZN(n15195) );
  INV_X1 U11507 ( .A(n9168), .ZN(n9169) );
  NAND2_X1 U11508 ( .A1(n9169), .A2(n12243), .ZN(n9170) );
  XNOR2_X1 U11509 ( .A(n9165), .B(n11274), .ZN(n9172) );
  XNOR2_X1 U11510 ( .A(n9172), .B(n10565), .ZN(n10487) );
  NAND2_X1 U11511 ( .A1(n9172), .A2(n10565), .ZN(n9173) );
  NAND2_X1 U11512 ( .A1(n10484), .A2(n9173), .ZN(n10564) );
  XNOR2_X1 U11513 ( .A(n10209), .B(n10802), .ZN(n9174) );
  XNOR2_X1 U11514 ( .A(n9174), .B(n12242), .ZN(n10563) );
  NAND2_X1 U11515 ( .A1(n9174), .A2(n10860), .ZN(n9175) );
  XNOR2_X1 U11516 ( .A(n10209), .B(n9176), .ZN(n9178) );
  XNOR2_X1 U11517 ( .A(n9178), .B(n12241), .ZN(n15209) );
  NAND2_X1 U11518 ( .A1(n9178), .A2(n12241), .ZN(n9179) );
  NAND2_X1 U11519 ( .A1(n15205), .A2(n9179), .ZN(n10835) );
  XNOR2_X1 U11520 ( .A(n10209), .B(n11089), .ZN(n9180) );
  XNOR2_X1 U11521 ( .A(n9180), .B(n12240), .ZN(n10834) );
  NAND2_X1 U11522 ( .A1(n10835), .A2(n10834), .ZN(n10833) );
  INV_X1 U11523 ( .A(n9180), .ZN(n9181) );
  NAND2_X1 U11524 ( .A1(n9181), .A2(n12240), .ZN(n9182) );
  NAND2_X1 U11525 ( .A1(n10833), .A2(n9182), .ZN(n11046) );
  XNOR2_X1 U11526 ( .A(n10209), .B(n11245), .ZN(n9189) );
  XNOR2_X1 U11527 ( .A(n9189), .B(n11250), .ZN(n11047) );
  XNOR2_X1 U11528 ( .A(n10209), .B(n11325), .ZN(n9190) );
  NAND2_X1 U11529 ( .A1(n9190), .A2(n11095), .ZN(n9188) );
  AND2_X1 U11530 ( .A1(n11047), .A2(n9188), .ZN(n15180) );
  XNOR2_X1 U11531 ( .A(n9255), .B(n15189), .ZN(n9183) );
  NAND2_X1 U11532 ( .A1(n9183), .A2(n11342), .ZN(n9199) );
  INV_X1 U11533 ( .A(n9183), .ZN(n9184) );
  NAND2_X1 U11534 ( .A1(n9184), .A2(n11442), .ZN(n9185) );
  NAND2_X1 U11535 ( .A1(n9199), .A2(n9185), .ZN(n15185) );
  INV_X1 U11536 ( .A(n15185), .ZN(n9186) );
  AND2_X1 U11537 ( .A1(n15180), .A2(n9186), .ZN(n9187) );
  NAND2_X1 U11538 ( .A1(n11046), .A2(n9187), .ZN(n9195) );
  INV_X1 U11539 ( .A(n9188), .ZN(n9193) );
  NAND2_X1 U11540 ( .A1(n9189), .A2(n12239), .ZN(n11281) );
  XNOR2_X1 U11541 ( .A(n9190), .B(n11095), .ZN(n11284) );
  INV_X1 U11542 ( .A(n11284), .ZN(n9191) );
  AND2_X1 U11543 ( .A1(n11281), .A2(n9191), .ZN(n9192) );
  OR2_X1 U11544 ( .A1(n9193), .A2(n9192), .ZN(n15182) );
  INV_X1 U11545 ( .A(n9199), .ZN(n9196) );
  XNOR2_X1 U11546 ( .A(n11522), .B(n10209), .ZN(n9197) );
  NOR3_X2 U11547 ( .A1(n15184), .A2(n9196), .A3(n9197), .ZN(n11438) );
  NOR2_X1 U11548 ( .A1(n11438), .A2(n11526), .ZN(n11434) );
  INV_X1 U11549 ( .A(n15184), .ZN(n9200) );
  INV_X1 U11550 ( .A(n9197), .ZN(n9198) );
  AOI21_X1 U11551 ( .B1(n9200), .B2(n9199), .A(n9198), .ZN(n11435) );
  XNOR2_X1 U11552 ( .A(n9201), .B(n12237), .ZN(n11450) );
  XOR2_X1 U11553 ( .A(n10209), .B(n11798), .Z(n11507) );
  INV_X1 U11554 ( .A(n11507), .ZN(n9202) );
  NOR2_X1 U11555 ( .A1(n9202), .A2(n12236), .ZN(n9204) );
  XNOR2_X1 U11556 ( .A(n12711), .B(n10209), .ZN(n9205) );
  INV_X1 U11557 ( .A(n12235), .ZN(n11711) );
  XNOR2_X1 U11558 ( .A(n9205), .B(n11711), .ZN(n11689) );
  AND2_X1 U11559 ( .A1(n9205), .A2(n12235), .ZN(n9206) );
  XNOR2_X1 U11560 ( .A(n11799), .B(n10209), .ZN(n11728) );
  INV_X1 U11561 ( .A(n11727), .ZN(n12234) );
  XNOR2_X1 U11562 ( .A(n12365), .B(n9255), .ZN(n9208) );
  NAND2_X1 U11563 ( .A1(n9208), .A2(n12570), .ZN(n11854) );
  NOR2_X1 U11564 ( .A1(n9208), .A2(n12570), .ZN(n11853) );
  XNOR2_X1 U11565 ( .A(n12636), .B(n10209), .ZN(n9209) );
  XNOR2_X1 U11566 ( .A(n9209), .B(n12372), .ZN(n12174) );
  INV_X1 U11567 ( .A(n9209), .ZN(n9210) );
  XNOR2_X1 U11568 ( .A(n12560), .B(n10209), .ZN(n9211) );
  XNOR2_X1 U11569 ( .A(n9211), .B(n12534), .ZN(n12210) );
  XNOR2_X1 U11570 ( .A(n12694), .B(n10209), .ZN(n9212) );
  XNOR2_X1 U11571 ( .A(n9212), .B(n12553), .ZN(n12145) );
  XNOR2_X1 U11572 ( .A(n12626), .B(n10209), .ZN(n9213) );
  XNOR2_X1 U11573 ( .A(n9213), .B(n12535), .ZN(n12190) );
  XNOR2_X1 U11574 ( .A(n12683), .B(n10209), .ZN(n9214) );
  NAND2_X1 U11575 ( .A1(n9214), .A2(n12202), .ZN(n9215) );
  OAI21_X1 U11576 ( .B1(n9214), .B2(n12202), .A(n9215), .ZN(n12155) );
  NOR2_X2 U11577 ( .A1(n9216), .A2(n6716), .ZN(n9217) );
  AOI21_X1 U11578 ( .B1(n9216), .B2(n6716), .A(n9217), .ZN(n12200) );
  NAND2_X1 U11579 ( .A1(n12200), .A2(n12488), .ZN(n12199) );
  INV_X1 U11580 ( .A(n9217), .ZN(n9218) );
  XNOR2_X1 U11581 ( .A(n12492), .B(n10209), .ZN(n9219) );
  INV_X1 U11582 ( .A(n12203), .ZN(n12389) );
  XNOR2_X1 U11583 ( .A(n12392), .B(n10209), .ZN(n9221) );
  NAND2_X1 U11584 ( .A1(n9221), .A2(n12489), .ZN(n9224) );
  INV_X1 U11585 ( .A(n9221), .ZN(n9222) );
  NAND2_X1 U11586 ( .A1(n9222), .A2(n12465), .ZN(n9223) );
  NAND2_X1 U11587 ( .A1(n9224), .A2(n9223), .ZN(n12181) );
  XNOR2_X1 U11588 ( .A(n12396), .B(n10209), .ZN(n9225) );
  NAND2_X1 U11589 ( .A1(n9225), .A2(n12448), .ZN(n9228) );
  INV_X1 U11590 ( .A(n9225), .ZN(n9226) );
  INV_X1 U11591 ( .A(n12448), .ZN(n12395) );
  NAND2_X1 U11592 ( .A1(n9226), .A2(n12395), .ZN(n9227) );
  XNOR2_X1 U11593 ( .A(n12398), .B(n9255), .ZN(n9229) );
  NOR2_X1 U11594 ( .A1(n9229), .A2(n12464), .ZN(n9230) );
  AOI21_X1 U11595 ( .B1(n9229), .B2(n12464), .A(n9230), .ZN(n12220) );
  XNOR2_X1 U11596 ( .A(n12591), .B(n9255), .ZN(n9274) );
  NOR2_X1 U11597 ( .A1(n9274), .A2(n12422), .ZN(n9254) );
  AOI21_X1 U11598 ( .B1(n9274), .B2(n12422), .A(n9254), .ZN(n9391) );
  NAND2_X1 U11599 ( .A1(n9390), .A2(n9391), .ZN(n9395) );
  INV_X1 U11600 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n9231) );
  NAND2_X1 U11601 ( .A1(n6712), .A2(n9231), .ZN(n9234) );
  INV_X1 U11602 ( .A(n9232), .ZN(n11433) );
  NAND2_X1 U11603 ( .A1(n11433), .A2(n9148), .ZN(n9233) );
  NAND2_X1 U11604 ( .A1(n9234), .A2(n9233), .ZN(n10535) );
  INV_X1 U11605 ( .A(n10535), .ZN(n12713) );
  NOR2_X1 U11606 ( .A1(P3_D_REG_24__SCAN_IN), .A2(P3_D_REG_27__SCAN_IN), .ZN(
        n9238) );
  NOR4_X1 U11607 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_26__SCAN_IN), .A4(P3_D_REG_17__SCAN_IN), .ZN(n9237) );
  NOR4_X1 U11608 ( .A1(P3_D_REG_18__SCAN_IN), .A2(P3_D_REG_29__SCAN_IN), .A3(
        P3_D_REG_10__SCAN_IN), .A4(P3_D_REG_31__SCAN_IN), .ZN(n9236) );
  NOR4_X1 U11609 ( .A1(P3_D_REG_22__SCAN_IN), .A2(P3_D_REG_25__SCAN_IN), .A3(
        P3_D_REG_20__SCAN_IN), .A4(P3_D_REG_19__SCAN_IN), .ZN(n9235) );
  NAND4_X1 U11610 ( .A1(n9238), .A2(n9237), .A3(n9236), .A4(n9235), .ZN(n9244)
         );
  NOR4_X1 U11611 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n9242) );
  NOR4_X1 U11612 ( .A1(P3_D_REG_12__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_11__SCAN_IN), .ZN(n9241) );
  NOR4_X1 U11613 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n9240) );
  NOR4_X1 U11614 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n9239) );
  NAND4_X1 U11615 ( .A1(n9242), .A2(n9241), .A3(n9240), .A4(n9239), .ZN(n9243)
         );
  OAI21_X1 U11616 ( .B1(n9244), .B2(n9243), .A(n6712), .ZN(n10454) );
  AND3_X1 U11617 ( .A1(n12713), .A2(n12715), .A3(n10454), .ZN(n11261) );
  NAND2_X1 U11618 ( .A1(n11952), .A2(n10504), .ZN(n9245) );
  NAND2_X1 U11619 ( .A1(n9245), .A2(n10635), .ZN(n9249) );
  NAND2_X1 U11620 ( .A1(n10504), .A2(n10427), .ZN(n9246) );
  NAND2_X1 U11621 ( .A1(n9246), .A2(n9145), .ZN(n9247) );
  NAND2_X1 U11622 ( .A1(n9247), .A2(n11952), .ZN(n9248) );
  NAND2_X1 U11623 ( .A1(n9249), .A2(n9248), .ZN(n11263) );
  NAND2_X1 U11624 ( .A1(n11952), .A2(n10635), .ZN(n15374) );
  NAND3_X1 U11625 ( .A1(n11261), .A2(n11263), .A3(n15374), .ZN(n9252) );
  NAND2_X1 U11626 ( .A1(n9145), .A2(n10427), .ZN(n10439) );
  INV_X1 U11627 ( .A(n10439), .ZN(n9250) );
  NAND2_X1 U11628 ( .A1(n9154), .A2(n9250), .ZN(n11259) );
  INV_X1 U11629 ( .A(n11259), .ZN(n9262) );
  AND3_X1 U11630 ( .A1(n10453), .A2(n10535), .A3(n10454), .ZN(n11264) );
  NAND2_X1 U11631 ( .A1(n9262), .A2(n11264), .ZN(n9251) );
  NAND2_X1 U11632 ( .A1(n9252), .A2(n9251), .ZN(n9253) );
  INV_X1 U11633 ( .A(n9254), .ZN(n9256) );
  XNOR2_X1 U11634 ( .A(n12419), .B(n9255), .ZN(n9277) );
  NAND4_X1 U11635 ( .A1(n9395), .A2(n15193), .A3(n9256), .A4(n9277), .ZN(n9282) );
  OR2_X1 U11636 ( .A1(n11261), .A2(n15376), .ZN(n9258) );
  NOR2_X1 U11637 ( .A1(n15374), .A2(n11265), .ZN(n9257) );
  NAND2_X1 U11638 ( .A1(n9258), .A2(n9257), .ZN(n12230) );
  AND2_X1 U11639 ( .A1(n10423), .A2(n10540), .ZN(n9259) );
  NAND2_X1 U11640 ( .A1(n11264), .A2(n9259), .ZN(n15203) );
  INV_X1 U11641 ( .A(n11263), .ZN(n9265) );
  NAND2_X1 U11642 ( .A1(n9267), .A2(n10449), .ZN(n10537) );
  AND2_X1 U11643 ( .A1(n9406), .A2(n9972), .ZN(n9261) );
  AND2_X1 U11644 ( .A1(n10537), .A2(n9261), .ZN(n9264) );
  INV_X1 U11645 ( .A(n11264), .ZN(n9268) );
  NAND2_X1 U11646 ( .A1(n9268), .A2(n9262), .ZN(n9263) );
  OAI211_X1 U11647 ( .C1(n11261), .C2(n9265), .A(n9264), .B(n9263), .ZN(n9266)
         );
  NAND2_X1 U11648 ( .A1(n9266), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9271) );
  NAND2_X1 U11649 ( .A1(n9267), .A2(n10423), .ZN(n11260) );
  INV_X1 U11650 ( .A(n11260), .ZN(n9269) );
  NAND3_X1 U11651 ( .A1(n9269), .A2(n10540), .A3(n9268), .ZN(n9270) );
  INV_X1 U11652 ( .A(n15215), .ZN(n12227) );
  NAND2_X1 U11653 ( .A1(n12227), .A2(n12427), .ZN(n9273) );
  OR2_X1 U11654 ( .A1(n15203), .A2(n15353), .ZN(n12222) );
  INV_X1 U11655 ( .A(n12222), .ZN(n12212) );
  AOI22_X1 U11656 ( .A1(n12212), .A2(n12422), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n9272) );
  OAI211_X1 U11657 ( .C1(n12232), .C2(n12224), .A(n9273), .B(n9272), .ZN(n9276) );
  NOR4_X1 U11658 ( .A1(n9277), .A2(n9274), .A3(n15207), .A4(n12422), .ZN(n9275) );
  AOI211_X1 U11659 ( .C1(n15213), .C2(n12426), .A(n9276), .B(n9275), .ZN(n9281) );
  INV_X1 U11660 ( .A(n9395), .ZN(n9279) );
  INV_X1 U11661 ( .A(n9277), .ZN(n9278) );
  NAND2_X1 U11662 ( .A1(n9279), .A2(n7580), .ZN(n9280) );
  NAND3_X1 U11663 ( .A1(n9282), .A2(n9281), .A3(n9280), .ZN(P3_U3160) );
  INV_X1 U11664 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n13724) );
  INV_X1 U11665 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9316) );
  AND2_X1 U11666 ( .A1(n9316), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n9315) );
  INV_X1 U11667 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n13497) );
  INV_X1 U11668 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n13658) );
  NAND2_X1 U11669 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(n13658), .ZN(n9313) );
  INV_X1 U11670 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n13716) );
  NOR2_X1 U11671 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n13716), .ZN(n9310) );
  INV_X1 U11672 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9307) );
  INV_X1 U11673 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n13542) );
  AOI22_X1 U11674 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(P3_ADDR_REG_12__SCAN_IN), 
        .B1(n13542), .B2(n9307), .ZN(n9357) );
  INV_X1 U11675 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n13539) );
  NAND2_X1 U11676 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(n13539), .ZN(n9305) );
  INV_X1 U11677 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9283) );
  AOI22_X1 U11678 ( .A1(P3_ADDR_REG_11__SCAN_IN), .A2(n9283), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n13539), .ZN(n9355) );
  INV_X1 U11679 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9300) );
  XOR2_X1 U11680 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), .Z(
        n9353) );
  INV_X1 U11681 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9298) );
  INV_X1 U11682 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9296) );
  INV_X1 U11683 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n15291) );
  NAND2_X1 U11684 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n15291), .ZN(n9295) );
  NOR2_X1 U11685 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n13672), .ZN(n9286) );
  NAND2_X1 U11686 ( .A1(P3_ADDR_REG_0__SCAN_IN), .A2(n9331), .ZN(n9330) );
  NOR2_X1 U11687 ( .A1(n9330), .A2(n9329), .ZN(n9285) );
  XNOR2_X1 U11688 ( .A(n9288), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n9327) );
  NOR2_X1 U11689 ( .A1(n9328), .A2(n9327), .ZN(n9287) );
  XNOR2_X1 U11690 ( .A(n14274), .B(P3_ADDR_REG_4__SCAN_IN), .ZN(n9324) );
  NOR2_X1 U11691 ( .A1(n9325), .A2(n9324), .ZN(n9290) );
  INV_X1 U11692 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n15273) );
  NOR2_X1 U11693 ( .A1(n9291), .A2(n15273), .ZN(n9293) );
  INV_X1 U11694 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n9340) );
  AND2_X1 U11695 ( .A1(n9340), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9294) );
  INV_X1 U11696 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n15309) );
  XNOR2_X1 U11697 ( .A(n15309), .B(n9298), .ZN(n9348) );
  NAND2_X1 U11698 ( .A1(n9349), .A2(n9348), .ZN(n9297) );
  NOR2_X1 U11699 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n9301), .ZN(n9303) );
  INV_X1 U11700 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n10649) );
  NAND2_X1 U11701 ( .A1(n9355), .A2(n9354), .ZN(n9304) );
  INV_X1 U11702 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9308) );
  AOI22_X1 U11703 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .B1(n9308), .B2(n13716), .ZN(n9364) );
  INV_X1 U11704 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9311) );
  AOI22_X1 U11705 ( .A1(P3_ADDR_REG_14__SCAN_IN), .A2(n9311), .B1(
        P1_ADDR_REG_14__SCAN_IN), .B2(n13658), .ZN(n9369) );
  NAND2_X1 U11706 ( .A1(n9370), .A2(n9369), .ZN(n9312) );
  NAND2_X1 U11707 ( .A1(n9313), .A2(n9312), .ZN(n9320) );
  INV_X1 U11708 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14927) );
  NAND2_X1 U11709 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n14927), .ZN(n9314) );
  AOI22_X1 U11710 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n13497), .B1(n9320), 
        .B2(n9314), .ZN(n9317) );
  OAI22_X1 U11711 ( .A1(n9315), .A2(n9317), .B1(P3_ADDR_REG_16__SCAN_IN), .B2(
        n9316), .ZN(n9377) );
  XNOR2_X1 U11712 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n9377), .ZN(n9378) );
  XOR2_X1 U11713 ( .A(n13724), .B(n9378), .Z(n9374) );
  XOR2_X1 U11714 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n9316), .Z(n9318) );
  XOR2_X1 U11715 ( .A(n9318), .B(n9317), .Z(n9372) );
  NAND2_X1 U11716 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n13497), .ZN(n9319) );
  OAI21_X1 U11717 ( .B1(n13497), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n9319), .ZN(
        n9321) );
  XOR2_X1 U11718 ( .A(n9321), .B(n9320), .Z(n14886) );
  XOR2_X1 U11719 ( .A(n10649), .B(n9322), .Z(n14696) );
  INV_X1 U11720 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n9334) );
  NAND2_X1 U11721 ( .A1(n9333), .A2(n9334), .ZN(n9335) );
  XOR2_X1 U11722 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n9326), .Z(n15449) );
  XOR2_X1 U11723 ( .A(n9328), .B(n9327), .Z(n14683) );
  OAI21_X1 U11724 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n9331), .A(n9330), .ZN(
        n15442) );
  NAND2_X1 U11725 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15442), .ZN(n15453) );
  NOR2_X1 U11726 ( .A1(n15453), .A2(n15452), .ZN(n15451) );
  NOR2_X1 U11727 ( .A1(n9332), .A2(n15451), .ZN(n14682) );
  XOR2_X1 U11728 ( .A(n9334), .B(n9333), .Z(n15438) );
  NAND2_X1 U11729 ( .A1(n6733), .A2(n15438), .ZN(n15437) );
  NAND2_X1 U11730 ( .A1(n9335), .A2(n15437), .ZN(n9337) );
  NAND2_X1 U11731 ( .A1(n9336), .A2(n9337), .ZN(n9338) );
  INV_X1 U11732 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15440) );
  NOR2_X1 U11733 ( .A1(n9339), .A2(n7270), .ZN(n9343) );
  XNOR2_X1 U11734 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n9340), .ZN(n9341) );
  XOR2_X1 U11735 ( .A(n9342), .B(n9341), .Z(n14686) );
  INV_X1 U11736 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n15017) );
  NOR2_X1 U11737 ( .A1(n9344), .A2(n15017), .ZN(n9347) );
  XOR2_X1 U11738 ( .A(n15291), .B(P1_ADDR_REG_7__SCAN_IN), .Z(n9346) );
  XOR2_X1 U11739 ( .A(n9346), .B(n9345), .Z(n15445) );
  XNOR2_X1 U11740 ( .A(n9349), .B(n9348), .ZN(n9351) );
  INV_X1 U11741 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14690) );
  XNOR2_X1 U11742 ( .A(n9351), .B(n9350), .ZN(n14689) );
  XOR2_X1 U11743 ( .A(n9353), .B(n9352), .Z(n14691) );
  XNOR2_X1 U11744 ( .A(n9355), .B(n9354), .ZN(n14874) );
  NAND2_X1 U11745 ( .A1(n14873), .A2(n14874), .ZN(n14872) );
  XOR2_X1 U11746 ( .A(n9358), .B(n9357), .Z(n9361) );
  INV_X1 U11747 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15036) );
  NAND2_X1 U11748 ( .A1(n9361), .A2(n9360), .ZN(n9362) );
  XOR2_X1 U11749 ( .A(n9364), .B(n9363), .Z(n9367) );
  INV_X1 U11750 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14879) );
  NAND2_X1 U11751 ( .A1(n9367), .A2(n9366), .ZN(n9368) );
  XNOR2_X1 U11752 ( .A(n9370), .B(n9369), .ZN(n14883) );
  NOR2_X1 U11753 ( .A1(n14882), .A2(n14883), .ZN(n9371) );
  NAND2_X1 U11754 ( .A1(n14883), .A2(n14882), .ZN(n14881) );
  INV_X1 U11755 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n14893) );
  NAND2_X1 U11756 ( .A1(n14893), .A2(n14892), .ZN(n14889) );
  NAND2_X1 U11757 ( .A1(n9374), .A2(n9375), .ZN(n9376) );
  INV_X1 U11758 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n14730) );
  INV_X1 U11759 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9385) );
  XOR2_X1 U11760 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(n9385), .Z(n9383) );
  NOR2_X1 U11761 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n9377), .ZN(n9380) );
  NOR2_X1 U11762 ( .A1(n13724), .A2(n9378), .ZN(n9379) );
  NOR2_X1 U11763 ( .A1(n9380), .A2(n9379), .ZN(n9382) );
  XNOR2_X1 U11764 ( .A(n9383), .B(n9382), .ZN(n14676) );
  NOR2_X1 U11765 ( .A1(n14677), .A2(n14676), .ZN(n9381) );
  NAND2_X1 U11766 ( .A1(n14677), .A2(n14676), .ZN(n14675) );
  NAND2_X1 U11767 ( .A1(n9383), .A2(n9382), .ZN(n9384) );
  OAI21_X1 U11768 ( .B1(n9385), .B2(P3_ADDR_REG_18__SCAN_IN), .A(n9384), .ZN(
        n9388) );
  XNOR2_X1 U11769 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n9386) );
  XNOR2_X1 U11770 ( .A(n9386), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n9387) );
  INV_X1 U11771 ( .A(n9391), .ZN(n9392) );
  NAND2_X1 U11772 ( .A1(n9393), .A2(n9392), .ZN(n9394) );
  NAND2_X1 U11773 ( .A1(n9395), .A2(n9394), .ZN(n9396) );
  NAND2_X1 U11774 ( .A1(n9396), .A2(n15193), .ZN(n9404) );
  INV_X1 U11775 ( .A(n12591), .ZN(n12440) );
  NOR2_X1 U11776 ( .A1(n12222), .A2(n9397), .ZN(n9400) );
  OAI22_X1 U11777 ( .A1(n12224), .A2(n12402), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n9398), .ZN(n9399) );
  AOI211_X1 U11778 ( .C1(n12227), .C2(n12438), .A(n9400), .B(n9399), .ZN(n9401) );
  OAI21_X1 U11779 ( .B1(n12440), .B2(n12230), .A(n9401), .ZN(n9402) );
  INV_X1 U11780 ( .A(n9402), .ZN(n9403) );
  NAND2_X1 U11781 ( .A1(n9404), .A2(n9403), .ZN(P3_U3154) );
  INV_X1 U11782 ( .A(n9591), .ZN(n9664) );
  INV_X1 U11783 ( .A(n9405), .ZN(n12714) );
  INV_X2 U11784 ( .A(n12245), .ZN(P3_U3897) );
  NOR2_X1 U11785 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), 
        .ZN(n9411) );
  NOR2_X1 U11786 ( .A1(n9413), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n9417) );
  INV_X1 U11787 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n9414) );
  NAND2_X1 U11788 ( .A1(n9417), .A2(n9414), .ZN(n9419) );
  NAND2_X1 U11789 ( .A1(n9419), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9415) );
  MUX2_X1 U11790 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9415), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n9416) );
  AND2_X1 U11791 ( .A1(n9535), .A2(n9416), .ZN(n9766) );
  INV_X1 U11792 ( .A(n9417), .ZN(n9422) );
  NAND2_X1 U11793 ( .A1(n9422), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9418) );
  MUX2_X1 U11794 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9418), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n9420) );
  NAND2_X1 U11795 ( .A1(n9420), .A2(n9419), .ZN(n11517) );
  NAND2_X1 U11796 ( .A1(n9413), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9421) );
  MUX2_X1 U11797 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9421), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n9423) );
  NAND2_X1 U11798 ( .A1(n9423), .A2(n9422), .ZN(n11447) );
  NOR2_X1 U11799 ( .A1(n11517), .A2(n11447), .ZN(n9424) );
  NAND2_X1 U11800 ( .A1(n9766), .A2(n9424), .ZN(n9779) );
  INV_X1 U11801 ( .A(n9779), .ZN(n9429) );
  INV_X1 U11802 ( .A(n9426), .ZN(n9427) );
  OAI21_X1 U11803 ( .B1(n9613), .B2(n9427), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n9428) );
  XNOR2_X1 U11804 ( .A(n9428), .B(n13635), .ZN(n11403) );
  NAND2_X1 U11805 ( .A1(n9429), .A2(n11403), .ZN(n9625) );
  OR2_X2 U11806 ( .A1(n9625), .A2(P2_U3088), .ZN(n13273) );
  INV_X1 U11807 ( .A(n13273), .ZN(P2_U3947) );
  NAND2_X1 U11808 ( .A1(n10081), .A2(n11401), .ZN(n9448) );
  NAND2_X1 U11809 ( .A1(n10366), .A2(n10092), .ZN(n9431) );
  NAND2_X1 U11810 ( .A1(n9431), .A2(n9430), .ZN(n9447) );
  INV_X1 U11811 ( .A(n9447), .ZN(n9432) );
  NAND2_X1 U11812 ( .A1(n9448), .A2(n9432), .ZN(n9814) );
  OR3_X1 U11813 ( .A1(n9814), .A2(n6684), .A3(n12005), .ZN(n14917) );
  INV_X1 U11814 ( .A(n14917), .ZN(n14332) );
  INV_X1 U11815 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10592) );
  MUX2_X1 U11816 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10592), .S(n14270), .Z(
        n9435) );
  INV_X1 U11817 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9459) );
  MUX2_X1 U11818 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n9459), .S(n9458), .Z(n9433)
         );
  AND2_X1 U11819 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14255) );
  NAND2_X1 U11820 ( .A1(n9433), .A2(n14255), .ZN(n14264) );
  NAND2_X1 U11821 ( .A1(n9458), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n14263) );
  NAND2_X1 U11822 ( .A1(n14264), .A2(n14263), .ZN(n9434) );
  NAND2_X1 U11823 ( .A1(n9435), .A2(n9434), .ZN(n14267) );
  NAND2_X1 U11824 ( .A1(n14270), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9439) );
  NAND2_X1 U11825 ( .A1(n14267), .A2(n9439), .ZN(n9438) );
  INV_X1 U11826 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n9436) );
  MUX2_X1 U11827 ( .A(n9436), .B(P1_REG2_REG_3__SCAN_IN), .S(n9836), .Z(n9437)
         );
  NAND2_X1 U11828 ( .A1(n9438), .A2(n9437), .ZN(n14284) );
  MUX2_X1 U11829 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n9436), .S(n9836), .Z(n9440)
         );
  NAND3_X1 U11830 ( .A1(n14267), .A2(n9440), .A3(n9439), .ZN(n9441) );
  AND3_X1 U11831 ( .A1(n14332), .A2(n14284), .A3(n9441), .ZN(n9453) );
  INV_X1 U11832 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n14974) );
  INV_X1 U11833 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9442) );
  MUX2_X1 U11834 ( .A(n9442), .B(P1_REG1_REG_2__SCAN_IN), .S(n14270), .Z(
        n14261) );
  NOR2_X1 U11835 ( .A1(n14262), .A2(n14261), .ZN(n14260) );
  AOI21_X1 U11836 ( .B1(P1_REG1_REG_2__SCAN_IN), .B2(n14270), .A(n14260), .ZN(
        n9446) );
  INV_X1 U11837 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9443) );
  MUX2_X1 U11838 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9443), .S(n9836), .Z(n9445)
         );
  NOR2_X1 U11839 ( .A1(n9446), .A2(n9445), .ZN(n9830) );
  INV_X1 U11840 ( .A(n9814), .ZN(n9444) );
  AND2_X1 U11841 ( .A1(n9444), .A2(n6684), .ZN(n14913) );
  AOI211_X1 U11842 ( .C1(n9446), .C2(n9445), .A(n9830), .B(n14298), .ZN(n9452)
         );
  NOR2_X1 U11843 ( .A1(n14921), .A2(n9836), .ZN(n9451) );
  NAND2_X1 U11844 ( .A1(n9448), .A2(n9447), .ZN(n14926) );
  OAI22_X1 U11845 ( .A1(n14926), .A2(n7275), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9449), .ZN(n9450) );
  OR4_X1 U11846 ( .A1(n9453), .A2(n9452), .A3(n9451), .A4(n9450), .ZN(P1_U3246) );
  NAND2_X1 U11847 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9457) );
  INV_X1 U11848 ( .A(n9454), .ZN(n9456) );
  AOI211_X1 U11849 ( .C1(n9457), .C2(n9456), .A(n9455), .B(n14298), .ZN(n9467)
         );
  INV_X1 U11850 ( .A(n9458), .ZN(n9491) );
  NOR2_X1 U11851 ( .A1(n14921), .A2(n9491), .ZN(n9466) );
  INV_X1 U11852 ( .A(n14255), .ZN(n9462) );
  MUX2_X1 U11853 ( .A(n9459), .B(P1_REG2_REG_1__SCAN_IN), .S(n9458), .Z(n9461)
         );
  INV_X1 U11854 ( .A(n14264), .ZN(n9460) );
  AOI211_X1 U11855 ( .C1(n9462), .C2(n9461), .A(n9460), .B(n14917), .ZN(n9465)
         );
  INV_X1 U11856 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9463) );
  OAI22_X1 U11857 ( .A1(n14926), .A2(n9284), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9463), .ZN(n9464) );
  OR4_X1 U11858 ( .A1(n9467), .A2(n9466), .A3(n9465), .A4(n9464), .ZN(P1_U3244) );
  AND2_X1 U11859 ( .A1(n9794), .A2(P2_U3088), .ZN(n11849) );
  NOR2_X1 U11860 ( .A1(n9794), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14071) );
  NAND2_X1 U11861 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n9468) );
  XNOR2_X1 U11862 ( .A(n9468), .B(P2_IR_REG_1__SCAN_IN), .ZN(n9911) );
  AOI22_X1 U11863 ( .A1(n14071), .A2(P1_DATAO_REG_1__SCAN_IN), .B1(n9911), 
        .B2(P2_STATE_REG_SCAN_IN), .ZN(n9469) );
  OAI21_X1 U11864 ( .B1(n9909), .B2(n6618), .A(n9469), .ZN(P2_U3326) );
  INV_X2 U11865 ( .A(n14071), .ZN(n11987) );
  OR2_X1 U11866 ( .A1(n9470), .A2(n6642), .ZN(n9472) );
  XNOR2_X1 U11867 ( .A(n9472), .B(n9471), .ZN(n9917) );
  OAI222_X1 U11868 ( .A1(n11987), .A2(n9918), .B1(n6618), .B2(n9920), .C1(
        P2_U3088), .C2(n9917), .ZN(P2_U3325) );
  NAND2_X1 U11869 ( .A1(n9794), .A2(P3_U3151), .ZN(n11995) );
  NOR2_X1 U11870 ( .A1(n9794), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12719) );
  OAI222_X1 U11871 ( .A1(P3_U3151), .A2(n15296), .B1(n11995), .B2(n9474), .C1(
        n11991), .C2(n9473), .ZN(P3_U3287) );
  INV_X1 U11872 ( .A(n9934), .ZN(n9487) );
  OR2_X1 U11873 ( .A1(n9494), .A2(n6642), .ZN(n9475) );
  XNOR2_X1 U11874 ( .A(n9475), .B(P2_IR_REG_3__SCAN_IN), .ZN(n9933) );
  INV_X1 U11875 ( .A(n9933), .ZN(n14993) );
  OAI222_X1 U11876 ( .A1(n11987), .A2(n9476), .B1(n6618), .B2(n9487), .C1(
        P2_U3088), .C2(n14993), .ZN(P2_U3324) );
  CLKBUF_X1 U11877 ( .A(n11995), .Z(n12725) );
  INV_X1 U11878 ( .A(SI_4_), .ZN(n9479) );
  INV_X1 U11879 ( .A(n9477), .ZN(n9478) );
  OAI222_X1 U11880 ( .A1(P3_U3151), .A2(n10062), .B1(n12725), .B2(n9479), .C1(
        n11991), .C2(n9478), .ZN(P3_U3291) );
  INV_X1 U11881 ( .A(SI_5_), .ZN(n9482) );
  INV_X1 U11882 ( .A(n9480), .ZN(n9481) );
  OAI222_X1 U11883 ( .A1(P3_U3151), .A2(n10064), .B1(n12725), .B2(n9482), .C1(
        n11991), .C2(n9481), .ZN(P3_U3290) );
  INV_X1 U11884 ( .A(SI_7_), .ZN(n9485) );
  INV_X1 U11885 ( .A(n9483), .ZN(n9484) );
  OAI222_X1 U11886 ( .A1(P3_U3151), .A2(n15279), .B1(n12725), .B2(n9485), .C1(
        n11991), .C2(n9484), .ZN(P3_U3288) );
  OAI222_X1 U11887 ( .A1(n12137), .A2(n9488), .B1(n14668), .B2(n9487), .C1(
        P1_U3086), .C2(n9836), .ZN(P1_U3352) );
  INV_X1 U11888 ( .A(n14270), .ZN(n9489) );
  OAI222_X1 U11889 ( .A1(n12137), .A2(n9490), .B1(n14668), .B2(n9920), .C1(
        P1_U3086), .C2(n9489), .ZN(P1_U3353) );
  OAI222_X1 U11890 ( .A1(n12137), .A2(n9492), .B1(n14668), .B2(n9909), .C1(
        P1_U3086), .C2(n9491), .ZN(P1_U3354) );
  INV_X1 U11891 ( .A(n10118), .ZN(n9501) );
  NAND2_X1 U11892 ( .A1(n9494), .A2(n9493), .ZN(n9504) );
  NAND2_X1 U11893 ( .A1(n9504), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9495) );
  XNOR2_X1 U11894 ( .A(n9495), .B(P2_IR_REG_4__SCAN_IN), .ZN(n10119) );
  INV_X1 U11895 ( .A(n10119), .ZN(n9496) );
  OAI222_X1 U11896 ( .A1(n11987), .A2(n9497), .B1(n6618), .B2(n9501), .C1(
        P2_U3088), .C2(n9496), .ZN(P2_U3323) );
  INV_X1 U11897 ( .A(n10678), .ZN(n11058) );
  OAI222_X1 U11898 ( .A1(P3_U3151), .A2(n11058), .B1(n12725), .B2(n9499), .C1(
        n11991), .C2(n9498), .ZN(P3_U3285) );
  INV_X1 U11899 ( .A(n14281), .ZN(n9500) );
  OAI222_X1 U11900 ( .A1(n12137), .A2(n9502), .B1(n14668), .B2(n9501), .C1(
        P1_U3086), .C2(n9500), .ZN(P1_U3351) );
  INV_X1 U11901 ( .A(n10259), .ZN(n9508) );
  OAI222_X1 U11902 ( .A1(n12137), .A2(n9503), .B1(n14668), .B2(n9508), .C1(
        P1_U3086), .C2(n9884), .ZN(P1_U3350) );
  NAND2_X1 U11903 ( .A1(n9506), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9505) );
  MUX2_X1 U11904 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9505), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n9507) );
  NAND2_X1 U11905 ( .A1(n9507), .A2(n9531), .ZN(n9708) );
  OAI222_X1 U11906 ( .A1(n11987), .A2(n9509), .B1(n6618), .B2(n9508), .C1(
        P2_U3088), .C2(n9708), .ZN(P2_U3322) );
  OAI222_X1 U11907 ( .A1(P3_U3151), .A2(n11065), .B1(n12725), .B2(n9511), .C1(
        n11991), .C2(n9510), .ZN(P3_U3284) );
  OAI222_X1 U11908 ( .A1(n11991), .A2(n9513), .B1(n12725), .B2(n9512), .C1(
        P3_U3151), .C2(n10162), .ZN(P3_U3294) );
  INV_X1 U11909 ( .A(n10403), .ZN(n9516) );
  NAND2_X1 U11910 ( .A1(n9531), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9514) );
  XNOR2_X1 U11911 ( .A(n9514), .B(P2_IR_REG_6__SCAN_IN), .ZN(n13276) );
  INV_X1 U11912 ( .A(n13276), .ZN(n13283) );
  OAI222_X1 U11913 ( .A1(n11987), .A2(n9515), .B1(n6618), .B2(n9516), .C1(
        P2_U3088), .C2(n13283), .ZN(P2_U3321) );
  OAI222_X1 U11914 ( .A1(n12137), .A2(n9517), .B1(n14668), .B2(n9516), .C1(
        P1_U3086), .C2(n7097), .ZN(P1_U3349) );
  INV_X1 U11915 ( .A(SI_3_), .ZN(n9520) );
  INV_X1 U11916 ( .A(n9518), .ZN(n9519) );
  OAI222_X1 U11917 ( .A1(P3_U3151), .A2(n10056), .B1(n12725), .B2(n9520), .C1(
        n11991), .C2(n9519), .ZN(P3_U3292) );
  INV_X1 U11918 ( .A(SI_2_), .ZN(n9523) );
  INV_X1 U11919 ( .A(n9521), .ZN(n9522) );
  OAI222_X1 U11920 ( .A1(P3_U3151), .A2(n10115), .B1(n12725), .B2(n9523), .C1(
        n11991), .C2(n9522), .ZN(P3_U3293) );
  OAI222_X1 U11921 ( .A1(P3_U3151), .A2(n10035), .B1(n11991), .B2(n9525), .C1(
        n9524), .C2(n12725), .ZN(P3_U3295) );
  OAI222_X1 U11922 ( .A1(n10651), .A2(P3_U3151), .B1(n11991), .B2(n9527), .C1(
        n9526), .C2(n11995), .ZN(P3_U3289) );
  INV_X1 U11923 ( .A(SI_9_), .ZN(n9528) );
  OAI222_X1 U11924 ( .A1(n15321), .A2(P3_U3151), .B1(n11991), .B2(n9529), .C1(
        n9528), .C2(n11995), .ZN(P3_U3286) );
  INV_X1 U11925 ( .A(n10574), .ZN(n9533) );
  INV_X1 U11926 ( .A(n9892), .ZN(n9870) );
  OAI222_X1 U11927 ( .A1(n12137), .A2(n9530), .B1(n14668), .B2(n9533), .C1(
        P1_U3086), .C2(n9870), .ZN(P1_U3348) );
  NAND2_X1 U11928 ( .A1(n9554), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9532) );
  XNOR2_X1 U11929 ( .A(n9532), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10575) );
  INV_X1 U11930 ( .A(n10575), .ZN(n15010) );
  OAI222_X1 U11931 ( .A1(n11987), .A2(n9534), .B1(n6618), .B2(n9533), .C1(
        P2_U3088), .C2(n15010), .ZN(P2_U3320) );
  INV_X1 U11932 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n9539) );
  INV_X1 U11933 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9536) );
  NAND2_X1 U11934 ( .A1(n10406), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n9549) );
  INV_X1 U11935 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9666) );
  OR2_X1 U11936 ( .A1(n10407), .A2(n9666), .ZN(n9548) );
  INV_X1 U11937 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9543) );
  OR2_X1 U11938 ( .A1(n12775), .A2(n9543), .ZN(n9547) );
  INV_X1 U11939 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10199) );
  NAND2_X1 U11940 ( .A1(n10172), .A2(P2_U3947), .ZN(n9550) );
  OAI21_X1 U11941 ( .B1(P2_U3947), .B2(n8406), .A(n9550), .ZN(P2_U3531) );
  INV_X1 U11942 ( .A(n11476), .ZN(n11239) );
  INV_X1 U11943 ( .A(n9551), .ZN(n9552) );
  OAI222_X1 U11944 ( .A1(P3_U3151), .A2(n11239), .B1(n12725), .B2(n9553), .C1(
        n11991), .C2(n9552), .ZN(P3_U3283) );
  INV_X1 U11945 ( .A(n10750), .ZN(n9557) );
  NAND2_X1 U11946 ( .A1(n9594), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9555) );
  XNOR2_X1 U11947 ( .A(n9555), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10751) );
  INV_X1 U11948 ( .A(n10751), .ZN(n9648) );
  OAI222_X1 U11949 ( .A1(n11987), .A2(n9556), .B1(n6618), .B2(n9557), .C1(
        P2_U3088), .C2(n9648), .ZN(P2_U3319) );
  INV_X1 U11950 ( .A(n9957), .ZN(n9902) );
  OAI222_X1 U11951 ( .A1(n12137), .A2(n9558), .B1(n14668), .B2(n9557), .C1(
        P1_U3086), .C2(n9902), .ZN(P1_U3347) );
  OAI222_X1 U11952 ( .A1(P3_U3151), .A2(n12260), .B1(n12725), .B2(n9560), .C1(
        n11991), .C2(n9559), .ZN(P3_U3282) );
  NOR2_X1 U11953 ( .A1(n6712), .A2(n12714), .ZN(n9562) );
  CLKBUF_X1 U11954 ( .A(n9562), .Z(n9589) );
  INV_X1 U11955 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n9561) );
  NOR2_X1 U11956 ( .A1(n9589), .A2(n9561), .ZN(P3_U3253) );
  INV_X1 U11957 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n9563) );
  NOR2_X1 U11958 ( .A1(n9589), .A2(n9563), .ZN(P3_U3240) );
  INV_X1 U11959 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n9564) );
  NOR2_X1 U11960 ( .A1(n9562), .A2(n9564), .ZN(P3_U3244) );
  INV_X1 U11961 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n9565) );
  NOR2_X1 U11962 ( .A1(n9589), .A2(n9565), .ZN(P3_U3248) );
  INV_X1 U11963 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n9566) );
  NOR2_X1 U11964 ( .A1(n9562), .A2(n9566), .ZN(P3_U3242) );
  INV_X1 U11965 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n9567) );
  NOR2_X1 U11966 ( .A1(n9589), .A2(n9567), .ZN(P3_U3249) );
  INV_X1 U11967 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n9568) );
  NOR2_X1 U11968 ( .A1(n9562), .A2(n9568), .ZN(P3_U3260) );
  INV_X1 U11969 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n9569) );
  NOR2_X1 U11970 ( .A1(n9589), .A2(n9569), .ZN(P3_U3259) );
  INV_X1 U11971 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n9570) );
  NOR2_X1 U11972 ( .A1(n9562), .A2(n9570), .ZN(P3_U3258) );
  INV_X1 U11973 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n9571) );
  NOR2_X1 U11974 ( .A1(n9589), .A2(n9571), .ZN(P3_U3263) );
  INV_X1 U11975 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n9572) );
  NOR2_X1 U11976 ( .A1(n9589), .A2(n9572), .ZN(P3_U3256) );
  INV_X1 U11977 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n9573) );
  NOR2_X1 U11978 ( .A1(n9589), .A2(n9573), .ZN(P3_U3255) );
  INV_X1 U11979 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n9574) );
  NOR2_X1 U11980 ( .A1(n9589), .A2(n9574), .ZN(P3_U3254) );
  INV_X1 U11981 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n13607) );
  NOR2_X1 U11982 ( .A1(n9562), .A2(n13607), .ZN(P3_U3238) );
  INV_X1 U11983 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n9575) );
  NOR2_X1 U11984 ( .A1(n9589), .A2(n9575), .ZN(P3_U3252) );
  INV_X1 U11985 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n9576) );
  NOR2_X1 U11986 ( .A1(n9589), .A2(n9576), .ZN(P3_U3257) );
  INV_X1 U11987 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n9577) );
  NOR2_X1 U11988 ( .A1(n9562), .A2(n9577), .ZN(P3_U3245) );
  INV_X1 U11989 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n9578) );
  NOR2_X1 U11990 ( .A1(n9562), .A2(n9578), .ZN(P3_U3234) );
  INV_X1 U11991 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n9579) );
  NOR2_X1 U11992 ( .A1(n9589), .A2(n9579), .ZN(P3_U3247) );
  INV_X1 U11993 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n9580) );
  NOR2_X1 U11994 ( .A1(n9562), .A2(n9580), .ZN(P3_U3262) );
  INV_X1 U11995 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n9581) );
  NOR2_X1 U11996 ( .A1(n9589), .A2(n9581), .ZN(P3_U3246) );
  INV_X1 U11997 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n9582) );
  NOR2_X1 U11998 ( .A1(n9589), .A2(n9582), .ZN(P3_U3250) );
  INV_X1 U11999 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n9583) );
  NOR2_X1 U12000 ( .A1(n9589), .A2(n9583), .ZN(P3_U3261) );
  INV_X1 U12001 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n9584) );
  NOR2_X1 U12002 ( .A1(n9562), .A2(n9584), .ZN(P3_U3243) );
  INV_X1 U12003 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n9585) );
  NOR2_X1 U12004 ( .A1(n9562), .A2(n9585), .ZN(P3_U3236) );
  INV_X1 U12005 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n13491) );
  NOR2_X1 U12006 ( .A1(n9562), .A2(n13491), .ZN(P3_U3241) );
  INV_X1 U12007 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n13728) );
  NOR2_X1 U12008 ( .A1(n9589), .A2(n13728), .ZN(P3_U3239) );
  INV_X1 U12009 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n9586) );
  NOR2_X1 U12010 ( .A1(n9589), .A2(n9586), .ZN(P3_U3237) );
  INV_X1 U12011 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n9587) );
  NOR2_X1 U12012 ( .A1(n9589), .A2(n9587), .ZN(P3_U3235) );
  INV_X1 U12013 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n9588) );
  NOR2_X1 U12014 ( .A1(n9589), .A2(n9588), .ZN(P3_U3251) );
  INV_X1 U12015 ( .A(n10081), .ZN(n10224) );
  NAND2_X1 U12016 ( .A1(n10224), .A2(n10078), .ZN(n14930) );
  INV_X1 U12017 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10075) );
  INV_X1 U12018 ( .A(n10079), .ZN(n9590) );
  AOI22_X1 U12019 ( .A1(n14930), .A2(n10075), .B1(n9591), .B2(n9590), .ZN(
        P1_U3446) );
  INV_X1 U12020 ( .A(n14926), .ZN(n14316) );
  NOR2_X1 U12021 ( .A1(n14316), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U12022 ( .A(P3_DATAO_REG_9__SCAN_IN), .ZN(n13551) );
  NAND2_X1 U12023 ( .A1(n11329), .A2(P3_U3897), .ZN(n9592) );
  OAI21_X1 U12024 ( .B1(P3_U3897), .B2(n13551), .A(n9592), .ZN(P3_U3500) );
  INV_X1 U12025 ( .A(n10876), .ZN(n9600) );
  INV_X1 U12026 ( .A(n10290), .ZN(n9968) );
  OAI222_X1 U12027 ( .A1(n12137), .A2(n9593), .B1(n14668), .B2(n9600), .C1(
        P1_U3086), .C2(n9968), .ZN(P1_U3346) );
  NAND2_X1 U12028 ( .A1(n9596), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9595) );
  MUX2_X1 U12029 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9595), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n9599) );
  INV_X1 U12030 ( .A(n9596), .ZN(n9598) );
  INV_X1 U12031 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n9597) );
  NAND2_X1 U12032 ( .A1(n9598), .A2(n9597), .ZN(n9736) );
  NAND2_X1 U12033 ( .A1(n9599), .A2(n9736), .ZN(n10879) );
  OAI222_X1 U12034 ( .A1(n11987), .A2(n10877), .B1(n6618), .B2(n9600), .C1(
        P2_U3088), .C2(n10879), .ZN(P2_U3318) );
  INV_X1 U12035 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9923) );
  MUX2_X1 U12036 ( .A(n9923), .B(P2_REG2_REG_2__SCAN_IN), .S(n9917), .Z(n9603)
         );
  INV_X1 U12037 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9759) );
  MUX2_X1 U12038 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n9759), .S(n9911), .Z(n9667)
         );
  AND2_X1 U12039 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9601) );
  NAND2_X1 U12040 ( .A1(n9667), .A2(n9601), .ZN(n9684) );
  NAND2_X1 U12041 ( .A1(n9911), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9683) );
  NAND2_X1 U12042 ( .A1(n9684), .A2(n9683), .ZN(n9602) );
  NAND2_X1 U12043 ( .A1(n9603), .A2(n9602), .ZN(n9687) );
  INV_X1 U12044 ( .A(n9917), .ZN(n9682) );
  NAND2_X1 U12045 ( .A1(n9682), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n9604) );
  NAND2_X1 U12046 ( .A1(n9687), .A2(n9604), .ZN(n15000) );
  INV_X1 U12047 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10334) );
  MUX2_X1 U12048 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10334), .S(n9933), .Z(
        n14999) );
  NAND2_X1 U12049 ( .A1(n15000), .A2(n14999), .ZN(n14998) );
  NAND2_X1 U12050 ( .A1(n9933), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9720) );
  NAND2_X1 U12051 ( .A1(n14998), .A2(n9720), .ZN(n9606) );
  INV_X1 U12052 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n13952) );
  MUX2_X1 U12053 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n13952), .S(n10119), .Z(
        n9605) );
  NAND2_X1 U12054 ( .A1(n9606), .A2(n9605), .ZN(n9722) );
  NAND2_X1 U12055 ( .A1(n10119), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9709) );
  NAND2_X1 U12056 ( .A1(n9722), .A2(n9709), .ZN(n9608) );
  INV_X1 U12057 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10392) );
  MUX2_X1 U12058 ( .A(n10392), .B(P2_REG2_REG_5__SCAN_IN), .S(n9708), .Z(n9607) );
  NAND2_X1 U12059 ( .A1(n9608), .A2(n9607), .ZN(n13279) );
  INV_X1 U12060 ( .A(n9708), .ZN(n10260) );
  NAND2_X1 U12061 ( .A1(n10260), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n13278) );
  NAND2_X1 U12062 ( .A1(n13279), .A2(n13278), .ZN(n9610) );
  INV_X1 U12063 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10525) );
  MUX2_X1 U12064 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10525), .S(n13276), .Z(
        n9609) );
  NAND2_X1 U12065 ( .A1(n9610), .A2(n9609), .ZN(n13281) );
  NAND2_X1 U12066 ( .A1(n13276), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n9611) );
  NAND2_X1 U12067 ( .A1(n13281), .A2(n9611), .ZN(n15014) );
  INV_X1 U12068 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10408) );
  MUX2_X1 U12069 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10408), .S(n10575), .Z(
        n15013) );
  NAND2_X1 U12070 ( .A1(n15014), .A2(n15013), .ZN(n15012) );
  OR2_X1 U12071 ( .A1(n15010), .A2(n10408), .ZN(n9630) );
  INV_X1 U12072 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n9612) );
  MUX2_X1 U12073 ( .A(n9612), .B(P2_REG2_REG_8__SCAN_IN), .S(n10751), .Z(n9629) );
  AOI21_X1 U12074 ( .B1(n15012), .B2(n9630), .A(n9629), .ZN(n9651) );
  NAND2_X1 U12075 ( .A1(n9783), .A2(n9614), .ZN(n9780) );
  INV_X1 U12076 ( .A(n9780), .ZN(n9615) );
  INV_X1 U12077 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n9781) );
  NAND2_X1 U12078 ( .A1(n9615), .A2(n9781), .ZN(n9618) );
  INV_X1 U12079 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n9616) );
  INV_X1 U12080 ( .A(n10168), .ZN(n13254) );
  NAND2_X1 U12081 ( .A1(n13254), .A2(n6610), .ZN(n9943) );
  INV_X1 U12082 ( .A(n11403), .ZN(n9624) );
  NAND2_X1 U12083 ( .A1(n9535), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9621) );
  OAI21_X1 U12084 ( .B1(n9943), .B2(n9624), .A(n6681), .ZN(n9626) );
  NAND2_X1 U12085 ( .A1(n9626), .A2(n9625), .ZN(n9641) );
  INV_X1 U12086 ( .A(n13253), .ZN(n13339) );
  NAND2_X1 U12087 ( .A1(n13339), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11789) );
  NOR2_X1 U12088 ( .A1(n11789), .A2(n9627), .ZN(n9628) );
  NAND2_X1 U12089 ( .A1(n9641), .A2(n9628), .ZN(n15026) );
  NAND3_X1 U12090 ( .A1(n15012), .A2(n9630), .A3(n9629), .ZN(n9631) );
  NAND2_X1 U12091 ( .A1(n15045), .A2(n9631), .ZN(n9646) );
  INV_X1 U12092 ( .A(n15035), .ZN(n15043) );
  AND2_X1 U12093 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n10773) );
  AND2_X1 U12094 ( .A1(n9627), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9632) );
  NAND2_X1 U12095 ( .A1(n9641), .A2(n9632), .ZN(n15051) );
  NOR2_X1 U12096 ( .A1(n15051), .A2(n9648), .ZN(n9633) );
  AOI211_X1 U12097 ( .C1(n15043), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n10773), .B(
        n9633), .ZN(n9645) );
  INV_X1 U12098 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n15170) );
  MUX2_X1 U12099 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n15170), .S(n10751), .Z(
        n9643) );
  INV_X1 U12100 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10412) );
  INV_X1 U12101 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n15159) );
  MUX2_X1 U12102 ( .A(n15159), .B(P2_REG1_REG_2__SCAN_IN), .S(n9917), .Z(n9679) );
  INV_X1 U12103 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10186) );
  MUX2_X1 U12104 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n10186), .S(n9911), .Z(n9670) );
  AND2_X1 U12105 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9669) );
  NAND2_X1 U12106 ( .A1(n9670), .A2(n9669), .ZN(n9668) );
  NAND2_X1 U12107 ( .A1(n9911), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9634) );
  NAND2_X1 U12108 ( .A1(n9668), .A2(n9634), .ZN(n9678) );
  NAND2_X1 U12109 ( .A1(n9679), .A2(n9678), .ZN(n9677) );
  NAND2_X1 U12110 ( .A1(n9682), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9635) );
  NAND2_X1 U12111 ( .A1(n9677), .A2(n9635), .ZN(n14991) );
  INV_X1 U12112 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n15161) );
  MUX2_X1 U12113 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n15161), .S(n9933), .Z(
        n14992) );
  NAND2_X1 U12114 ( .A1(n14991), .A2(n14992), .ZN(n14990) );
  NAND2_X1 U12115 ( .A1(n9933), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9636) );
  NAND2_X1 U12116 ( .A1(n14990), .A2(n9636), .ZN(n9715) );
  INV_X1 U12117 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n15163) );
  MUX2_X1 U12118 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n15163), .S(n10119), .Z(
        n9716) );
  NAND2_X1 U12119 ( .A1(n9715), .A2(n9716), .ZN(n9714) );
  NAND2_X1 U12120 ( .A1(n10119), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9637) );
  NAND2_X1 U12121 ( .A1(n9714), .A2(n9637), .ZN(n9704) );
  INV_X1 U12122 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n15165) );
  MUX2_X1 U12123 ( .A(n15165), .B(P2_REG1_REG_5__SCAN_IN), .S(n9708), .Z(n9705) );
  NAND2_X1 U12124 ( .A1(n9704), .A2(n9705), .ZN(n9703) );
  NAND2_X1 U12125 ( .A1(n10260), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9638) );
  NAND2_X1 U12126 ( .A1(n9703), .A2(n9638), .ZN(n13288) );
  INV_X1 U12127 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n15167) );
  MUX2_X1 U12128 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n15167), .S(n13276), .Z(
        n13289) );
  NAND2_X1 U12129 ( .A1(n13288), .A2(n13289), .ZN(n13287) );
  NAND2_X1 U12130 ( .A1(n13276), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9639) );
  NAND2_X1 U12131 ( .A1(n13287), .A2(n9639), .ZN(n15005) );
  MUX2_X1 U12132 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10412), .S(n10575), .Z(
        n15004) );
  NAND2_X1 U12133 ( .A1(n15005), .A2(n15004), .ZN(n15003) );
  OAI21_X1 U12134 ( .B1(n10412), .B2(n15010), .A(n15003), .ZN(n9642) );
  OR2_X1 U12135 ( .A1(n9627), .A2(P2_U3088), .ZN(n11850) );
  NOR2_X1 U12136 ( .A1(n11850), .A2(n13339), .ZN(n9640) );
  NAND2_X1 U12137 ( .A1(n9641), .A2(n9640), .ZN(n15037) );
  INV_X1 U12138 ( .A(n15037), .ZN(n14984) );
  NAND2_X1 U12139 ( .A1(n9642), .A2(n9643), .ZN(n9647) );
  OAI211_X1 U12140 ( .C1(n9643), .C2(n9642), .A(n14984), .B(n9647), .ZN(n9644)
         );
  OAI211_X1 U12141 ( .C1(n9651), .C2(n9646), .A(n9645), .B(n9644), .ZN(
        P2_U3222) );
  INV_X1 U12142 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n11128) );
  MUX2_X1 U12143 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n11128), .S(n10879), .Z(
        n9650) );
  OAI21_X1 U12144 ( .B1(n15170), .B2(n9648), .A(n9647), .ZN(n9649) );
  NOR2_X1 U12145 ( .A1(n9649), .A2(n9650), .ZN(n9698) );
  AOI21_X1 U12146 ( .B1(n9650), .B2(n9649), .A(n9698), .ZN(n9659) );
  AOI21_X1 U12147 ( .B1(n10751), .B2(P2_REG2_REG_8__SCAN_IN), .A(n9651), .ZN(
        n9654) );
  INV_X1 U12148 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n9652) );
  MUX2_X1 U12149 ( .A(n9652), .B(P2_REG2_REG_9__SCAN_IN), .S(n10879), .Z(n9653) );
  NAND2_X1 U12150 ( .A1(n9654), .A2(n9653), .ZN(n9691) );
  OAI21_X1 U12151 ( .B1(n9654), .B2(n9653), .A(n9691), .ZN(n9657) );
  NOR2_X1 U12152 ( .A1(n15035), .A2(n7264), .ZN(n9656) );
  NAND2_X1 U12153 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n10921) );
  OAI21_X1 U12154 ( .B1(n15051), .B2(n10879), .A(n10921), .ZN(n9655) );
  AOI211_X1 U12155 ( .C1(n9657), .C2(n15045), .A(n9656), .B(n9655), .ZN(n9658)
         );
  OAI21_X1 U12156 ( .B1(n9659), .B2(n15037), .A(n9658), .ZN(P2_U3223) );
  OAI222_X1 U12157 ( .A1(P3_U3151), .A2(n12282), .B1(n11995), .B2(n9661), .C1(
        n11991), .C2(n9660), .ZN(P3_U3281) );
  INV_X1 U12158 ( .A(P3_DATAO_REG_10__SCAN_IN), .ZN(n13718) );
  NAND2_X1 U12159 ( .A1(n11342), .A2(P3_U3897), .ZN(n9662) );
  OAI21_X1 U12160 ( .B1(P3_U3897), .B2(n13718), .A(n9662), .ZN(P3_U3501) );
  INV_X1 U12161 ( .A(n14930), .ZN(n14929) );
  OAI22_X1 U12162 ( .A1(n14929), .A2(P1_D_REG_0__SCAN_IN), .B1(n9664), .B2(
        n9663), .ZN(n9665) );
  INV_X1 U12163 ( .A(n9665), .ZN(P1_U3445) );
  INV_X1 U12164 ( .A(n9684), .ZN(n9676) );
  NOR2_X1 U12165 ( .A1(n15026), .A2(n9666), .ZN(n14983) );
  AOI22_X1 U12166 ( .A1(n14983), .A2(P2_IR_REG_0__SCAN_IN), .B1(n15045), .B2(
        n9667), .ZN(n9675) );
  INV_X1 U12167 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9994) );
  INV_X1 U12168 ( .A(n15051), .ZN(n15032) );
  AOI22_X1 U12169 ( .A1(n15043), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(n15032), 
        .B2(n9911), .ZN(n9672) );
  OAI211_X1 U12170 ( .C1(n9670), .C2(n9669), .A(n14984), .B(n9668), .ZN(n9671)
         );
  OAI211_X1 U12171 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n9994), .A(n9672), .B(
        n9671), .ZN(n9673) );
  INV_X1 U12172 ( .A(n9673), .ZN(n9674) );
  OAI21_X1 U12173 ( .B1(n9676), .B2(n9675), .A(n9674), .ZN(P2_U3215) );
  INV_X1 U12174 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10478) );
  OAI211_X1 U12175 ( .C1(n9679), .C2(n9678), .A(n14984), .B(n9677), .ZN(n9680)
         );
  OAI21_X1 U12176 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n10478), .A(n9680), .ZN(
        n9681) );
  AOI21_X1 U12177 ( .B1(n9682), .B2(n15032), .A(n9681), .ZN(n9689) );
  MUX2_X1 U12178 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n9923), .S(n9917), .Z(n9685)
         );
  NAND3_X1 U12179 ( .A1(n9685), .A2(n9684), .A3(n9683), .ZN(n9686) );
  NAND3_X1 U12180 ( .A1(n15045), .A2(n9687), .A3(n9686), .ZN(n9688) );
  OAI211_X1 U12181 ( .C1(n6915), .C2(n15035), .A(n9689), .B(n9688), .ZN(
        P2_U3216) );
  NAND2_X1 U12182 ( .A1(n9736), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9690) );
  XNOR2_X1 U12183 ( .A(n9690), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10988) );
  INV_X1 U12184 ( .A(n10988), .ZN(n9745) );
  NAND2_X1 U12185 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n11001)
         );
  OAI21_X1 U12186 ( .B1(n15051), .B2(n9745), .A(n11001), .ZN(n9697) );
  INV_X1 U12187 ( .A(n10879), .ZN(n9692) );
  OAI21_X1 U12188 ( .B1(n9692), .B2(P2_REG2_REG_9__SCAN_IN), .A(n9691), .ZN(
        n9695) );
  INV_X1 U12189 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n9693) );
  MUX2_X1 U12190 ( .A(n9693), .B(P2_REG2_REG_10__SCAN_IN), .S(n10988), .Z(
        n9694) );
  NOR2_X1 U12191 ( .A1(n9695), .A2(n9694), .ZN(n9735) );
  AOI211_X1 U12192 ( .C1(n9695), .C2(n9694), .A(n15026), .B(n9735), .ZN(n9696)
         );
  AOI211_X1 U12193 ( .C1(n15043), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n9697), .B(
        n9696), .ZN(n9702) );
  AOI21_X1 U12194 ( .B1(n10879), .B2(n11128), .A(n9698), .ZN(n9700) );
  INV_X1 U12195 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n15172) );
  MUX2_X1 U12196 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n15172), .S(n10988), .Z(
        n9699) );
  NAND2_X1 U12197 ( .A1(n9700), .A2(n9699), .ZN(n9744) );
  OAI211_X1 U12198 ( .C1(n9700), .C2(n9699), .A(n9744), .B(n14984), .ZN(n9701)
         );
  NAND2_X1 U12199 ( .A1(n9702), .A2(n9701), .ZN(P2_U3224) );
  AND2_X1 U12200 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n10280) );
  OAI211_X1 U12201 ( .C1(n9705), .C2(n9704), .A(n14984), .B(n9703), .ZN(n9706)
         );
  INV_X1 U12202 ( .A(n9706), .ZN(n9707) );
  AOI211_X1 U12203 ( .C1(n15032), .C2(n10260), .A(n10280), .B(n9707), .ZN(
        n9713) );
  MUX2_X1 U12204 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10392), .S(n9708), .Z(n9710) );
  NAND3_X1 U12205 ( .A1(n9710), .A2(n9722), .A3(n9709), .ZN(n9711) );
  NAND3_X1 U12206 ( .A1(n15045), .A2(n13279), .A3(n9711), .ZN(n9712) );
  OAI211_X1 U12207 ( .C1(n15440), .C2(n15035), .A(n9713), .B(n9712), .ZN(
        P2_U3219) );
  AND2_X1 U12208 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n10142) );
  OAI211_X1 U12209 ( .C1(n9716), .C2(n9715), .A(n14984), .B(n9714), .ZN(n9717)
         );
  INV_X1 U12210 ( .A(n9717), .ZN(n9718) );
  AOI211_X1 U12211 ( .C1(n15032), .C2(n10119), .A(n10142), .B(n9718), .ZN(
        n9724) );
  MUX2_X1 U12212 ( .A(n13952), .B(P2_REG2_REG_4__SCAN_IN), .S(n10119), .Z(
        n9719) );
  NAND3_X1 U12213 ( .A1(n14998), .A2(n9720), .A3(n9719), .ZN(n9721) );
  NAND3_X1 U12214 ( .A1(n15045), .A2(n9722), .A3(n9721), .ZN(n9723) );
  OAI211_X1 U12215 ( .C1(n9334), .C2(n15035), .A(n9724), .B(n9723), .ZN(
        P2_U3218) );
  INV_X1 U12216 ( .A(n12303), .ZN(n12317) );
  INV_X1 U12217 ( .A(n9725), .ZN(n9726) );
  OAI222_X1 U12218 ( .A1(P3_U3151), .A2(n12317), .B1(n11995), .B2(n13779), 
        .C1(n11991), .C2(n9726), .ZN(P3_U3280) );
  INV_X1 U12219 ( .A(n11302), .ZN(n9732) );
  INV_X1 U12220 ( .A(n11029), .ZN(n10716) );
  OAI222_X1 U12221 ( .A1(n12137), .A2(n9727), .B1(n14668), .B2(n9732), .C1(
        n10716), .C2(P1_U3086), .ZN(P1_U3343) );
  NAND2_X1 U12222 ( .A1(n9729), .A2(n9728), .ZN(n9750) );
  NAND2_X1 U12223 ( .A1(n9750), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9730) );
  XNOR2_X1 U12224 ( .A(n9730), .B(P2_IR_REG_12__SCAN_IN), .ZN(n15031) );
  INV_X1 U12225 ( .A(n15031), .ZN(n10303) );
  OAI222_X1 U12226 ( .A1(P2_U3088), .A2(n10303), .B1(n6618), .B2(n9732), .C1(
        n9731), .C2(n11987), .ZN(P2_U3315) );
  INV_X1 U12227 ( .A(n10987), .ZN(n9734) );
  INV_X1 U12228 ( .A(n10553), .ZN(n10296) );
  OAI222_X1 U12229 ( .A1(n12137), .A2(n9733), .B1(n14668), .B2(n9734), .C1(
        P1_U3086), .C2(n10296), .ZN(P1_U3345) );
  OAI222_X1 U12230 ( .A1(n11987), .A2(n13506), .B1(n6618), .B2(n9734), .C1(
        P2_U3088), .C2(n9745), .ZN(P2_U3317) );
  AOI21_X1 U12231 ( .B1(n10988), .B2(P2_REG2_REG_10__SCAN_IN), .A(n9735), .ZN(
        n9739) );
  INV_X1 U12232 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10302) );
  OAI21_X1 U12233 ( .B1(n9736), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9737) );
  XNOR2_X1 U12234 ( .A(n9737), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11152) );
  MUX2_X1 U12235 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n10302), .S(n11152), .Z(
        n9738) );
  NAND2_X1 U12236 ( .A1(n9739), .A2(n9738), .ZN(n15025) );
  OAI21_X1 U12237 ( .B1(n9739), .B2(n9738), .A(n15025), .ZN(n9743) );
  INV_X1 U12238 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n9740) );
  NOR2_X1 U12239 ( .A1(n15035), .A2(n9740), .ZN(n9742) );
  INV_X1 U12240 ( .A(n11152), .ZN(n10309) );
  NAND2_X1 U12241 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n11167)
         );
  OAI21_X1 U12242 ( .B1(n15051), .B2(n10309), .A(n11167), .ZN(n9741) );
  AOI211_X1 U12243 ( .C1(n9743), .C2(n15045), .A(n9742), .B(n9741), .ZN(n9749)
         );
  OAI21_X1 U12244 ( .B1(n15172), .B2(n9745), .A(n9744), .ZN(n9747) );
  INV_X1 U12245 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n15175) );
  MUX2_X1 U12246 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n15175), .S(n11152), .Z(
        n9746) );
  NAND2_X1 U12247 ( .A1(n9747), .A2(n9746), .ZN(n10308) );
  OAI211_X1 U12248 ( .C1(n9747), .C2(n9746), .A(n10308), .B(n14984), .ZN(n9748) );
  NAND2_X1 U12249 ( .A1(n9749), .A2(n9748), .ZN(P2_U3225) );
  NAND2_X1 U12250 ( .A1(n9752), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9751) );
  MUX2_X1 U12251 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9751), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n9753) );
  INV_X1 U12252 ( .A(n11359), .ZN(n9755) );
  INV_X1 U12253 ( .A(n11358), .ZN(n9756) );
  INV_X1 U12254 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9754) );
  OAI222_X1 U12255 ( .A1(P2_U3088), .A2(n9755), .B1(n6618), .B2(n9756), .C1(
        n9754), .C2(n11987), .ZN(P2_U3314) );
  OAI222_X1 U12256 ( .A1(P1_U3086), .A2(n11205), .B1(n14668), .B2(n9756), .C1(
        n13698), .C2(n12137), .ZN(P1_U3342) );
  INV_X1 U12257 ( .A(P3_DATAO_REG_21__SCAN_IN), .ZN(n13612) );
  INV_X1 U12258 ( .A(n12202), .ZN(n12384) );
  NAND2_X1 U12259 ( .A1(n12384), .A2(P3_U3897), .ZN(n9757) );
  OAI21_X1 U12260 ( .B1(P3_U3897), .B2(n13612), .A(n9757), .ZN(P3_U3512) );
  INV_X1 U12261 ( .A(n11151), .ZN(n9818) );
  OAI222_X1 U12262 ( .A1(n11987), .A2(n9758), .B1(n6618), .B2(n9818), .C1(
        P2_U3088), .C2(n10309), .ZN(P2_U3316) );
  OR2_X1 U12263 ( .A1(n10407), .A2(n9759), .ZN(n9763) );
  NAND2_X1 U12264 ( .A1(n10406), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n9760) );
  XNOR2_X1 U12265 ( .A(n11447), .B(P2_B_REG_SCAN_IN), .ZN(n9764) );
  NAND2_X1 U12266 ( .A1(n9764), .A2(n11517), .ZN(n9765) );
  AND2_X1 U12267 ( .A1(n9765), .A2(n9766), .ZN(n15073) );
  INV_X1 U12268 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15084) );
  INV_X1 U12269 ( .A(n9766), .ZN(n11704) );
  AOI22_X1 U12270 ( .A1(n15073), .A2(n15084), .B1(n11704), .B2(n11517), .ZN(
        n10165) );
  NOR4_X1 U12271 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n9775) );
  INV_X1 U12272 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n15076) );
  INV_X1 U12273 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n15074) );
  INV_X1 U12274 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n15075) );
  INV_X1 U12275 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n15077) );
  NAND4_X1 U12276 ( .A1(n15076), .A2(n15074), .A3(n15075), .A4(n15077), .ZN(
        n9772) );
  NOR4_X1 U12277 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n9770) );
  NOR4_X1 U12278 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n9769) );
  NOR4_X1 U12279 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9768) );
  NOR4_X1 U12280 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n9767) );
  NAND4_X1 U12281 ( .A1(n9770), .A2(n9769), .A3(n9768), .A4(n9767), .ZN(n9771)
         );
  NOR4_X1 U12282 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        n9772), .A4(n9771), .ZN(n9774) );
  NOR4_X1 U12283 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n9773) );
  NAND3_X1 U12284 ( .A1(n9775), .A2(n9774), .A3(n9773), .ZN(n9776) );
  NAND2_X1 U12285 ( .A1(n15073), .A2(n9776), .ZN(n10163) );
  AND2_X1 U12286 ( .A1(n10165), .A2(n10163), .ZN(n10194) );
  INV_X1 U12287 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15080) );
  NAND2_X1 U12288 ( .A1(n15073), .A2(n15080), .ZN(n9778) );
  NAND2_X1 U12289 ( .A1(n11704), .A2(n11447), .ZN(n9777) );
  NAND2_X1 U12290 ( .A1(n9778), .A2(n9777), .ZN(n15081) );
  INV_X1 U12291 ( .A(n15081), .ZN(n10182) );
  NAND2_X1 U12292 ( .A1(n10194), .A2(n10182), .ZN(n9787) );
  AND2_X1 U12293 ( .A1(n9779), .A2(n11403), .ZN(n9788) );
  OR2_X1 U12294 ( .A1(n9787), .A2(n15085), .ZN(n9791) );
  NAND2_X1 U12295 ( .A1(n9780), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9782) );
  XNOR2_X1 U12296 ( .A(n9782), .B(n9781), .ZN(n9906) );
  INV_X1 U12297 ( .A(n9783), .ZN(n9784) );
  NAND2_X1 U12298 ( .A1(n9784), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9785) );
  XNOR2_X1 U12299 ( .A(n9785), .B(P2_IR_REG_19__SCAN_IN), .ZN(n13214) );
  NAND2_X1 U12300 ( .A1(n9906), .A2(n13331), .ZN(n13252) );
  NOR2_X2 U12301 ( .A1(n9791), .A2(n13252), .ZN(n14795) );
  INV_X1 U12302 ( .A(n9627), .ZN(n9786) );
  NAND2_X1 U12303 ( .A1(n14795), .A2(n13949), .ZN(n12962) );
  INV_X1 U12304 ( .A(n6610), .ZN(n13215) );
  INV_X1 U12305 ( .A(n13174), .ZN(n13226) );
  NAND2_X1 U12306 ( .A1(n9787), .A2(n10164), .ZN(n9790) );
  INV_X1 U12307 ( .A(n13252), .ZN(n13222) );
  OR2_X1 U12308 ( .A1(n9943), .A2(n13222), .ZN(n10193) );
  AND2_X1 U12309 ( .A1(n10193), .A2(n9788), .ZN(n9789) );
  NAND2_X1 U12310 ( .A1(n9790), .A2(n9789), .ZN(n9941) );
  NOR2_X1 U12311 ( .A1(n9941), .A2(P2_U3088), .ZN(n10006) );
  INV_X1 U12312 ( .A(n10006), .ZN(n9801) );
  INV_X1 U12313 ( .A(n9791), .ZN(n9802) );
  AND2_X1 U12314 ( .A1(n15150), .A2(n9943), .ZN(n9792) );
  NAND2_X1 U12315 ( .A1(n9802), .A2(n9792), .ZN(n12967) );
  INV_X1 U12316 ( .A(n9793), .ZN(n10198) );
  INV_X1 U12317 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9799) );
  NAND2_X1 U12318 ( .A1(n9794), .A2(SI_0_), .ZN(n9796) );
  NAND2_X1 U12319 ( .A1(n9796), .A2(n9795), .ZN(n9798) );
  NAND2_X1 U12320 ( .A1(n9798), .A2(n9797), .ZN(n14073) );
  MUX2_X1 U12321 ( .A(n9799), .B(n14073), .S(n10878), .Z(n12976) );
  NAND2_X1 U12322 ( .A1(n10172), .A2(n12976), .ZN(n12970) );
  NOR3_X1 U12323 ( .A1(n12967), .A2(n11374), .A3(n12970), .ZN(n9800) );
  AOI21_X1 U12324 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n9801), .A(n9800), .ZN(
        n9806) );
  AOI21_X1 U12325 ( .B1(n6611), .B2(n10172), .A(n12967), .ZN(n9804) );
  INV_X1 U12326 ( .A(n9906), .ZN(n13184) );
  AND2_X1 U12327 ( .A1(n10198), .A2(n13184), .ZN(n10337) );
  NAND2_X1 U12328 ( .A1(n9802), .A2(n10337), .ZN(n9803) );
  NAND2_X1 U12329 ( .A1(n9803), .A2(n13957), .ZN(n14796) );
  INV_X1 U12330 ( .A(n12976), .ZN(n12973) );
  OAI21_X1 U12331 ( .B1(n9804), .B2(n14796), .A(n12973), .ZN(n9805) );
  OAI211_X1 U12332 ( .C1(n10324), .C2(n12962), .A(n9806), .B(n9805), .ZN(
        P2_U3204) );
  INV_X1 U12333 ( .A(n12307), .ZN(n14733) );
  INV_X1 U12334 ( .A(n9807), .ZN(n9808) );
  OAI222_X1 U12335 ( .A1(P3_U3151), .A2(n14733), .B1(n11995), .B2(n9809), .C1(
        n11991), .C2(n9808), .ZN(P3_U3279) );
  INV_X1 U12336 ( .A(n6684), .ZN(n11974) );
  NOR2_X1 U12337 ( .A1(n6684), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9810) );
  NOR2_X1 U12338 ( .A1(n12005), .A2(n9810), .ZN(n14259) );
  OAI21_X1 U12339 ( .B1(n11974), .B2(P1_REG1_REG_0__SCAN_IN), .A(n14259), .ZN(
        n9811) );
  MUX2_X1 U12340 ( .A(n9811), .B(n14259), .S(P1_IR_REG_0__SCAN_IN), .Z(n9813)
         );
  INV_X1 U12341 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9812) );
  OAI22_X1 U12342 ( .A1(n9814), .A2(n9813), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9812), .ZN(n9816) );
  NOR3_X1 U12343 ( .A1(n14298), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n8410), .ZN(
        n9815) );
  AOI211_X1 U12344 ( .C1(n14316), .C2(P1_ADDR_REG_0__SCAN_IN), .A(n9816), .B(
        n9815), .ZN(n9817) );
  INV_X1 U12345 ( .A(n9817), .ZN(P1_U3243) );
  INV_X1 U12346 ( .A(n10712), .ZN(n10708) );
  OAI222_X1 U12347 ( .A1(n9819), .A2(n12137), .B1(P1_U3086), .B2(n10708), .C1(
        n14668), .C2(n9818), .ZN(P1_U3344) );
  OAI21_X1 U12348 ( .B1(n14965), .B2(n14701), .A(n9820), .ZN(n9821) );
  OAI21_X1 U12349 ( .B1(n8910), .B2(n14466), .A(n9821), .ZN(n10221) );
  INV_X1 U12350 ( .A(n9822), .ZN(n9823) );
  NOR2_X1 U12351 ( .A1(n10098), .A2(n9823), .ZN(n10223) );
  NOR2_X1 U12352 ( .A1(n10221), .A2(n10223), .ZN(n9829) );
  INV_X1 U12353 ( .A(n10364), .ZN(n9824) );
  AND2_X2 U12354 ( .A1(n9825), .A2(n9824), .ZN(n14982) );
  NAND2_X1 U12355 ( .A1(n14980), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9826) );
  OAI21_X1 U12356 ( .B1(n9829), .B2(n14980), .A(n9826), .ZN(P1_U3528) );
  INV_X1 U12357 ( .A(n14973), .ZN(n14971) );
  INV_X1 U12358 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9827) );
  OR2_X1 U12359 ( .A1(n14973), .A2(n9827), .ZN(n9828) );
  OAI21_X1 U12360 ( .B1(n9829), .B2(n14971), .A(n9828), .ZN(P1_U3459) );
  MUX2_X1 U12361 ( .A(n7096), .B(P1_REG1_REG_6__SCAN_IN), .S(n9858), .Z(n9835)
         );
  INV_X1 U12362 ( .A(n9836), .ZN(n9831) );
  AOI21_X1 U12363 ( .B1(n9831), .B2(P1_REG1_REG_3__SCAN_IN), .A(n9830), .ZN(
        n14279) );
  INV_X1 U12364 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9832) );
  MUX2_X1 U12365 ( .A(n9832), .B(P1_REG1_REG_4__SCAN_IN), .S(n14281), .Z(
        n14278) );
  INV_X1 U12366 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9833) );
  MUX2_X1 U12367 ( .A(n9833), .B(P1_REG1_REG_5__SCAN_IN), .S(n9884), .Z(n9874)
         );
  NOR2_X1 U12368 ( .A1(n9834), .A2(n9835), .ZN(n9854) );
  AOI211_X1 U12369 ( .C1(n9835), .C2(n9834), .A(n14298), .B(n9854), .ZN(n9850)
         );
  INV_X1 U12370 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10817) );
  MUX2_X1 U12371 ( .A(n10817), .B(P1_REG2_REG_5__SCAN_IN), .S(n9884), .Z(n9841) );
  OR2_X1 U12372 ( .A1(n9836), .A2(n9436), .ZN(n14283) );
  NAND2_X1 U12373 ( .A1(n14284), .A2(n14283), .ZN(n9839) );
  MUX2_X1 U12374 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n9837), .S(n14281), .Z(n9838) );
  NAND2_X1 U12375 ( .A1(n9839), .A2(n9838), .ZN(n14286) );
  NAND2_X1 U12376 ( .A1(n14281), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9876) );
  NAND2_X1 U12377 ( .A1(n14286), .A2(n9876), .ZN(n9840) );
  NAND2_X1 U12378 ( .A1(n9841), .A2(n9840), .ZN(n9879) );
  NAND2_X1 U12379 ( .A1(n9842), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9847) );
  NAND2_X1 U12380 ( .A1(n9879), .A2(n9847), .ZN(n9845) );
  INV_X1 U12381 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9843) );
  MUX2_X1 U12382 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n9843), .S(n9858), .Z(n9844)
         );
  NAND2_X1 U12383 ( .A1(n9845), .A2(n9844), .ZN(n9864) );
  MUX2_X1 U12384 ( .A(n9843), .B(P1_REG2_REG_6__SCAN_IN), .S(n9858), .Z(n9846)
         );
  NAND3_X1 U12385 ( .A1(n9879), .A2(n9847), .A3(n9846), .ZN(n9848) );
  AND3_X1 U12386 ( .A1(n14332), .A2(n9864), .A3(n9848), .ZN(n9849) );
  NOR2_X1 U12387 ( .A1(n9850), .A2(n9849), .ZN(n9853) );
  INV_X1 U12388 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n13662) );
  NOR2_X1 U12389 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n13662), .ZN(n9851) );
  AOI21_X1 U12390 ( .B1(n14316), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n9851), .ZN(
        n9852) );
  OAI211_X1 U12391 ( .C1(n7097), .C2(n14921), .A(n9853), .B(n9852), .ZN(
        P1_U3249) );
  INV_X1 U12392 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9855) );
  MUX2_X1 U12393 ( .A(n9855), .B(P1_REG1_REG_7__SCAN_IN), .S(n9892), .Z(n9856)
         );
  AOI211_X1 U12394 ( .C1(n9857), .C2(n9856), .A(n14298), .B(n9888), .ZN(n9872)
         );
  NAND2_X1 U12395 ( .A1(n9858), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9863) );
  NAND2_X1 U12396 ( .A1(n9864), .A2(n9863), .ZN(n9861) );
  INV_X1 U12397 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9859) );
  MUX2_X1 U12398 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n9859), .S(n9892), .Z(n9860)
         );
  NAND2_X1 U12399 ( .A1(n9861), .A2(n9860), .ZN(n9897) );
  MUX2_X1 U12400 ( .A(n9859), .B(P1_REG2_REG_7__SCAN_IN), .S(n9892), .Z(n9862)
         );
  NAND3_X1 U12401 ( .A1(n9864), .A2(n9863), .A3(n9862), .ZN(n9865) );
  NAND3_X1 U12402 ( .A1(n14332), .A2(n9897), .A3(n9865), .ZN(n9869) );
  NOR2_X1 U12403 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9866), .ZN(n9867) );
  AOI21_X1 U12404 ( .B1(n14316), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n9867), .ZN(
        n9868) );
  OAI211_X1 U12405 ( .C1(n14921), .C2(n9870), .A(n9869), .B(n9868), .ZN(n9871)
         );
  OR2_X1 U12406 ( .A1(n9872), .A2(n9871), .ZN(P1_U3250) );
  OAI21_X1 U12407 ( .B1(n9875), .B2(n9874), .A(n9873), .ZN(n9881) );
  MUX2_X1 U12408 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10817), .S(n9884), .Z(n9877) );
  NAND3_X1 U12409 ( .A1(n9877), .A2(n14286), .A3(n9876), .ZN(n9878) );
  AND3_X1 U12410 ( .A1(n14332), .A2(n9879), .A3(n9878), .ZN(n9880) );
  AOI21_X1 U12411 ( .B1(n9881), .B2(n14913), .A(n9880), .ZN(n9883) );
  AND2_X1 U12412 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10941) );
  AOI21_X1 U12413 ( .B1(n14316), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n10941), .ZN(
        n9882) );
  OAI211_X1 U12414 ( .C1(n9884), .C2(n14921), .A(n9883), .B(n9882), .ZN(
        P1_U3248) );
  INV_X1 U12415 ( .A(n9885), .ZN(n9886) );
  OAI222_X1 U12416 ( .A1(P3_U3151), .A2(n12320), .B1(n12725), .B2(n9887), .C1(
        n11991), .C2(n9886), .ZN(P3_U3278) );
  INV_X1 U12417 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9889) );
  MUX2_X1 U12418 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n9889), .S(n9957), .Z(n9890)
         );
  OAI21_X1 U12419 ( .B1(n9891), .B2(n9890), .A(n9954), .ZN(n9904) );
  NAND2_X1 U12420 ( .A1(n9892), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9896) );
  NAND2_X1 U12421 ( .A1(n9897), .A2(n9896), .ZN(n9894) );
  INV_X1 U12422 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10980) );
  MUX2_X1 U12423 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10980), .S(n9957), .Z(n9893) );
  NAND2_X1 U12424 ( .A1(n9894), .A2(n9893), .ZN(n9963) );
  MUX2_X1 U12425 ( .A(n10980), .B(P1_REG2_REG_8__SCAN_IN), .S(n9957), .Z(n9895) );
  NAND3_X1 U12426 ( .A1(n9897), .A2(n9896), .A3(n9895), .ZN(n9898) );
  NAND3_X1 U12427 ( .A1(n14332), .A2(n9963), .A3(n9898), .ZN(n9901) );
  NAND2_X1 U12428 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n11958) );
  INV_X1 U12429 ( .A(n11958), .ZN(n9899) );
  AOI21_X1 U12430 ( .B1(n14316), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n9899), .ZN(
        n9900) );
  OAI211_X1 U12431 ( .C1(n14921), .C2(n9902), .A(n9901), .B(n9900), .ZN(n9903)
         );
  AOI21_X1 U12432 ( .B1(n9904), .B2(n14913), .A(n9903), .ZN(n9905) );
  INV_X1 U12433 ( .A(n9905), .ZN(P1_U3251) );
  XNOR2_X1 U12434 ( .A(n12971), .B(n10168), .ZN(n9908) );
  AND2_X1 U12435 ( .A1(n12973), .A2(n10172), .ZN(n10170) );
  AOI22_X1 U12436 ( .A1(n11155), .A2(n12976), .B1(n10170), .B2(n6611), .ZN(
        n9990) );
  NAND2_X1 U12437 ( .A1(n6613), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n9913) );
  AND3_X2 U12438 ( .A1(n9914), .A2(n9913), .A3(n9912), .ZN(n9993) );
  NOR2_X1 U12439 ( .A1(n9920), .A2(n13164), .ZN(n9921) );
  XNOR2_X1 U12440 ( .A(n9932), .B(n15093), .ZN(n9929) );
  NAND2_X1 U12441 ( .A1(n10406), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n9927) );
  OR2_X1 U12442 ( .A1(n12775), .A2(n15159), .ZN(n9925) );
  NAND2_X1 U12443 ( .A1(n10319), .A2(n6611), .ZN(n9928) );
  NAND2_X1 U12444 ( .A1(n9929), .A2(n9928), .ZN(n9930) );
  OAI21_X1 U12445 ( .B1(n9929), .B2(n9928), .A(n9930), .ZN(n10004) );
  INV_X1 U12446 ( .A(n9930), .ZN(n9931) );
  NOR2_X1 U12447 ( .A1(n10003), .A2(n9931), .ZN(n10126) );
  AOI22_X1 U12448 ( .A1(n6613), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n12733), 
        .B2(n9933), .ZN(n9936) );
  NAND2_X1 U12449 ( .A1(n9934), .A2(n10117), .ZN(n9935) );
  XNOR2_X1 U12450 ( .A(n12895), .B(n12988), .ZN(n10123) );
  NAND2_X1 U12451 ( .A1(n10406), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n9940) );
  OR2_X1 U12452 ( .A1(n12775), .A2(n15161), .ZN(n9938) );
  OR2_X1 U12453 ( .A1(n10407), .A2(n10334), .ZN(n9937) );
  NAND2_X1 U12454 ( .A1(n13948), .A2(n6611), .ZN(n10122) );
  XNOR2_X1 U12455 ( .A(n10123), .B(n10122), .ZN(n10125) );
  XNOR2_X1 U12456 ( .A(n10126), .B(n10125), .ZN(n9952) );
  NAND2_X1 U12457 ( .A1(n9941), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14799) );
  INV_X1 U12458 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9942) );
  OAI22_X1 U12459 ( .A1(n14799), .A2(P2_REG3_REG_3__SCAN_IN), .B1(
        P2_STATE_REG_SCAN_IN), .B2(n9942), .ZN(n9950) );
  INV_X1 U12460 ( .A(n10319), .ZN(n9992) );
  NAND2_X1 U12461 ( .A1(n14795), .A2(n14787), .ZN(n12963) );
  INV_X2 U12462 ( .A(n10407), .ZN(n12900) );
  NAND2_X1 U12463 ( .A1(n12900), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9948) );
  INV_X1 U12464 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9944) );
  OR2_X1 U12465 ( .A1(n12845), .A2(n9944), .ZN(n9947) );
  OAI21_X1 U12466 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n10133), .ZN(n13956) );
  OR2_X1 U12467 ( .A1(n10135), .A2(n13956), .ZN(n9946) );
  OR2_X1 U12468 ( .A1(n12775), .A2(n15163), .ZN(n9945) );
  INV_X1 U12469 ( .A(n13274), .ZN(n10388) );
  OAI22_X1 U12470 ( .A1(n9992), .A2(n12963), .B1(n12962), .B2(n10388), .ZN(
        n9949) );
  AOI211_X1 U12471 ( .C1(n12988), .C2(n14796), .A(n9950), .B(n9949), .ZN(n9951) );
  OAI21_X1 U12472 ( .B1(n9952), .B2(n12967), .A(n9951), .ZN(P2_U3190) );
  INV_X1 U12473 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9953) );
  MUX2_X1 U12474 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n9953), .S(n10290), .Z(n9956) );
  OAI21_X1 U12475 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n9957), .A(n9954), .ZN(
        n9955) );
  NAND2_X1 U12476 ( .A1(n9955), .A2(n9956), .ZN(n10287) );
  OAI21_X1 U12477 ( .B1(n9956), .B2(n9955), .A(n10287), .ZN(n9970) );
  NAND2_X1 U12478 ( .A1(n9957), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9962) );
  NAND2_X1 U12479 ( .A1(n9963), .A2(n9962), .ZN(n9960) );
  MUX2_X1 U12480 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n9958), .S(n10290), .Z(n9959) );
  NAND2_X1 U12481 ( .A1(n9960), .A2(n9959), .ZN(n10295) );
  MUX2_X1 U12482 ( .A(n9958), .B(P1_REG2_REG_9__SCAN_IN), .S(n10290), .Z(n9961) );
  NAND3_X1 U12483 ( .A1(n9963), .A2(n9962), .A3(n9961), .ZN(n9964) );
  NAND3_X1 U12484 ( .A1(n14332), .A2(n10295), .A3(n9964), .ZN(n9967) );
  NAND2_X1 U12485 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n14906) );
  INV_X1 U12486 ( .A(n14906), .ZN(n9965) );
  AOI21_X1 U12487 ( .B1(n14316), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n9965), .ZN(
        n9966) );
  OAI211_X1 U12488 ( .C1(n14921), .C2(n9968), .A(n9967), .B(n9966), .ZN(n9969)
         );
  AOI21_X1 U12489 ( .B1(n9970), .B2(n14913), .A(n9969), .ZN(n9971) );
  INV_X1 U12490 ( .A(n9971), .ZN(P1_U3252) );
  INV_X1 U12491 ( .A(n9972), .ZN(n9974) );
  OAI21_X1 U12492 ( .B1(n10458), .B2(n9974), .A(n9973), .ZN(n9984) );
  NOR2_X1 U12493 ( .A1(n10540), .A2(n8263), .ZN(n9982) );
  OR2_X1 U12494 ( .A1(n9984), .A2(n9982), .ZN(n9977) );
  MUX2_X1 U12495 ( .A(n9977), .B(n12245), .S(n9975), .Z(n15320) );
  NOR2_X1 U12496 ( .A1(n9977), .A2(n9976), .ZN(n15264) );
  NAND2_X1 U12497 ( .A1(P3_U3897), .A2(n12354), .ZN(n15322) );
  NOR2_X2 U12498 ( .A1(n9977), .A2(n12340), .ZN(n15329) );
  INV_X1 U12499 ( .A(n15329), .ZN(n15297) );
  NAND3_X1 U12500 ( .A1(n15333), .A2(n15322), .A3(n15297), .ZN(n9981) );
  INV_X1 U12501 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10051) );
  INV_X1 U12502 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n9978) );
  MUX2_X1 U12503 ( .A(n10051), .B(n9978), .S(n7638), .Z(n9979) );
  NAND2_X1 U12504 ( .A1(n9979), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10149) );
  OAI21_X1 U12505 ( .B1(n6991), .B2(n9979), .A(n10149), .ZN(n9980) );
  NAND2_X1 U12506 ( .A1(n9981), .A2(n9980), .ZN(n9986) );
  INV_X1 U12507 ( .A(n9982), .ZN(n9983) );
  AOI22_X1 U12508 ( .A1(n15326), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n9985) );
  OAI211_X1 U12509 ( .C1(n15320), .C2(n10035), .A(n9986), .B(n9985), .ZN(
        P3_U3182) );
  INV_X1 U12510 ( .A(n9987), .ZN(n9989) );
  NAND2_X1 U12511 ( .A1(n9989), .A2(n9988), .ZN(n9991) );
  XNOR2_X1 U12512 ( .A(n9991), .B(n9990), .ZN(n9999) );
  INV_X1 U12513 ( .A(n12963), .ZN(n9997) );
  NOR2_X1 U12514 ( .A1(n12962), .A2(n9992), .ZN(n9996) );
  OAI22_X1 U12515 ( .A1(n11848), .A2(n9993), .B1(n10006), .B2(n9994), .ZN(
        n9995) );
  AOI211_X1 U12516 ( .C1(n9997), .C2(n10172), .A(n9996), .B(n9995), .ZN(n9998)
         );
  OAI21_X1 U12517 ( .B1(n9999), .B2(n12967), .A(n9998), .ZN(P2_U3194) );
  INV_X1 U12518 ( .A(n12344), .ZN(n12336) );
  INV_X1 U12519 ( .A(n10000), .ZN(n10001) );
  OAI222_X1 U12520 ( .A1(P3_U3151), .A2(n12336), .B1(n12725), .B2(n10002), 
        .C1(n11991), .C2(n10001), .ZN(P3_U3277) );
  AOI21_X1 U12521 ( .B1(n10005), .B2(n10004), .A(n10003), .ZN(n10010) );
  INV_X1 U12522 ( .A(n13948), .ZN(n10140) );
  OAI22_X1 U12523 ( .A1(n10324), .A2(n12963), .B1(n12962), .B2(n10140), .ZN(
        n10008) );
  OAI22_X1 U12524 ( .A1(n11848), .A2(n15093), .B1(n10006), .B2(n10478), .ZN(
        n10007) );
  NOR2_X1 U12525 ( .A1(n10008), .A2(n10007), .ZN(n10009) );
  OAI21_X1 U12526 ( .B1(n10010), .B2(n12967), .A(n10009), .ZN(P2_U3209) );
  INV_X1 U12527 ( .A(n15322), .ZN(n15305) );
  INV_X1 U12528 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10012) );
  INV_X1 U12529 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10011) );
  MUX2_X1 U12530 ( .A(n10012), .B(n10011), .S(n7638), .Z(n10013) );
  INV_X1 U12531 ( .A(n10162), .ZN(n10037) );
  NAND2_X1 U12532 ( .A1(n10013), .A2(n10037), .ZN(n10103) );
  INV_X1 U12533 ( .A(n10013), .ZN(n10014) );
  NAND2_X1 U12534 ( .A1(n10014), .A2(n10162), .ZN(n10015) );
  NAND2_X1 U12535 ( .A1(n10103), .A2(n10015), .ZN(n10148) );
  NAND2_X1 U12536 ( .A1(n10150), .A2(n10103), .ZN(n10021) );
  INV_X1 U12537 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10017) );
  INV_X1 U12538 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10016) );
  MUX2_X1 U12539 ( .A(n10017), .B(n10016), .S(n7638), .Z(n10018) );
  NAND2_X1 U12540 ( .A1(n10018), .A2(n10050), .ZN(n15219) );
  INV_X1 U12541 ( .A(n10018), .ZN(n10019) );
  NAND2_X1 U12542 ( .A1(n10019), .A2(n10115), .ZN(n10020) );
  AND2_X1 U12543 ( .A1(n15219), .A2(n10020), .ZN(n10102) );
  NAND2_X1 U12544 ( .A1(n10021), .A2(n10102), .ZN(n15220) );
  NAND2_X1 U12545 ( .A1(n15220), .A2(n15219), .ZN(n10026) );
  INV_X1 U12546 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10022) );
  INV_X1 U12547 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15225) );
  MUX2_X1 U12548 ( .A(n10022), .B(n15225), .S(n6688), .Z(n10023) );
  INV_X1 U12549 ( .A(n10056), .ZN(n15231) );
  NAND2_X1 U12550 ( .A1(n10023), .A2(n15231), .ZN(n10027) );
  INV_X1 U12551 ( .A(n10023), .ZN(n10024) );
  NAND2_X1 U12552 ( .A1(n10024), .A2(n10056), .ZN(n10025) );
  AND2_X1 U12553 ( .A1(n10027), .A2(n10025), .ZN(n15217) );
  NAND2_X1 U12554 ( .A1(n10026), .A2(n15217), .ZN(n15222) );
  NAND2_X1 U12555 ( .A1(n15222), .A2(n10027), .ZN(n15239) );
  MUX2_X1 U12556 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n14735), .Z(n10028) );
  INV_X1 U12557 ( .A(n10062), .ZN(n15241) );
  XNOR2_X1 U12558 ( .A(n10028), .B(n15241), .ZN(n15238) );
  NAND2_X1 U12559 ( .A1(n15239), .A2(n15238), .ZN(n15237) );
  INV_X1 U12560 ( .A(n10028), .ZN(n10029) );
  NAND2_X1 U12561 ( .A1(n10029), .A2(n15241), .ZN(n10030) );
  NAND2_X1 U12562 ( .A1(n15237), .A2(n10030), .ZN(n15255) );
  MUX2_X1 U12563 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n14735), .Z(n10031) );
  NAND2_X1 U12564 ( .A1(n10031), .A2(n10064), .ZN(n15253) );
  NAND2_X1 U12565 ( .A1(n15255), .A2(n15253), .ZN(n10033) );
  INV_X1 U12566 ( .A(n10031), .ZN(n10032) );
  INV_X1 U12567 ( .A(n10064), .ZN(n15265) );
  NAND2_X1 U12568 ( .A1(n10032), .A2(n15265), .ZN(n15252) );
  NAND2_X1 U12569 ( .A1(n10033), .A2(n15252), .ZN(n10665) );
  MUX2_X1 U12570 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n14735), .Z(n10666) );
  XNOR2_X1 U12571 ( .A(n10666), .B(n10667), .ZN(n10664) );
  XNOR2_X1 U12572 ( .A(n10665), .B(n10664), .ZN(n10073) );
  NAND2_X1 U12573 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n15202) );
  INV_X1 U12574 ( .A(n15202), .ZN(n10034) );
  AOI21_X1 U12575 ( .B1(n15326), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n10034), .ZN(
        n10049) );
  INV_X1 U12576 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15425) );
  AOI22_X1 U12577 ( .A1(n10667), .A2(n15425), .B1(P3_REG1_REG_6__SCAN_IN), 
        .B2(n10651), .ZN(n10046) );
  NAND2_X1 U12578 ( .A1(P3_REG1_REG_4__SCAN_IN), .A2(n10062), .ZN(n10042) );
  INV_X1 U12579 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10462) );
  AOI22_X1 U12580 ( .A1(n15241), .A2(n10462), .B1(P3_REG1_REG_4__SCAN_IN), 
        .B2(n10062), .ZN(n15246) );
  NAND2_X1 U12581 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n10035), .ZN(n10036) );
  NOR3_X1 U12582 ( .A1(n9978), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n10038) );
  AOI21_X1 U12583 ( .B1(n10037), .B2(n10036), .A(n10038), .ZN(n10147) );
  NAND2_X1 U12584 ( .A1(n10147), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n10146) );
  INV_X1 U12585 ( .A(n10038), .ZN(n10039) );
  MUX2_X1 U12586 ( .A(P3_REG1_REG_2__SCAN_IN), .B(n10016), .S(n10050), .Z(
        n10108) );
  XNOR2_X1 U12587 ( .A(n10041), .B(n10056), .ZN(n15226) );
  NAND2_X1 U12588 ( .A1(n15226), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n10040) );
  NAND2_X1 U12589 ( .A1(n10042), .A2(n15245), .ZN(n10043) );
  NAND2_X1 U12590 ( .A1(n10043), .A2(n10064), .ZN(n10044) );
  XNOR2_X1 U12591 ( .A(n10043), .B(n15265), .ZN(n15261) );
  NAND2_X1 U12592 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(n15261), .ZN(n15260) );
  NAND2_X1 U12593 ( .A1(n10044), .A2(n15260), .ZN(n10045) );
  NAND2_X1 U12594 ( .A1(n10046), .A2(n10045), .ZN(n10652) );
  OAI21_X1 U12595 ( .B1(n10046), .B2(n10045), .A(n10652), .ZN(n10047) );
  NAND2_X1 U12596 ( .A1(n15329), .A2(n10047), .ZN(n10048) );
  OAI211_X1 U12597 ( .C1(n15320), .C2(n10651), .A(n10049), .B(n10048), .ZN(
        n10072) );
  XNOR2_X1 U12598 ( .A(n10050), .B(P3_REG2_REG_2__SCAN_IN), .ZN(n10101) );
  NOR2_X1 U12599 ( .A1(n10051), .A2(n6991), .ZN(n10053) );
  NAND2_X1 U12600 ( .A1(n10052), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10054) );
  OAI21_X1 U12601 ( .B1(n10162), .B2(n10053), .A(n10054), .ZN(n10155) );
  NAND2_X1 U12602 ( .A1(n10101), .A2(n10100), .ZN(n10099) );
  NAND2_X1 U12603 ( .A1(n10115), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10055) );
  NAND2_X1 U12604 ( .A1(n10099), .A2(n10055), .ZN(n10057) );
  NAND2_X1 U12605 ( .A1(n10057), .A2(n10056), .ZN(n10059) );
  INV_X1 U12606 ( .A(n10059), .ZN(n10060) );
  NAND2_X1 U12607 ( .A1(P3_REG2_REG_4__SCAN_IN), .A2(n10062), .ZN(n10061) );
  OAI21_X1 U12608 ( .B1(P3_REG2_REG_4__SCAN_IN), .B2(n10062), .A(n10061), .ZN(
        n15236) );
  INV_X1 U12609 ( .A(n10063), .ZN(n10066) );
  INV_X1 U12610 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n15257) );
  OAI21_X1 U12611 ( .B1(n10065), .B2(n10064), .A(n10063), .ZN(n15258) );
  NAND2_X1 U12612 ( .A1(P3_REG2_REG_6__SCAN_IN), .A2(n10651), .ZN(n10067) );
  OAI21_X1 U12613 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n10651), .A(n10067), .ZN(
        n10068) );
  AOI21_X1 U12614 ( .B1(n10069), .B2(n10068), .A(n10639), .ZN(n10070) );
  NOR2_X1 U12615 ( .A1(n15333), .A2(n10070), .ZN(n10071) );
  AOI211_X1 U12616 ( .C1(n15305), .C2(n10073), .A(n10072), .B(n10071), .ZN(
        n10074) );
  INV_X1 U12617 ( .A(n10074), .ZN(P3_U3188) );
  NOR2_X1 U12618 ( .A1(n10076), .A2(n10075), .ZN(n10077) );
  OR2_X1 U12619 ( .A1(n10078), .A2(n10077), .ZN(n10080) );
  NAND2_X1 U12620 ( .A1(n10080), .A2(n10079), .ZN(n10363) );
  OR3_X1 U12621 ( .A1(n10364), .A2(n10363), .A3(n10081), .ZN(n10091) );
  NAND2_X1 U12622 ( .A1(n10091), .A2(n14498), .ZN(n14844) );
  NOR2_X1 U12623 ( .A1(n10091), .A2(n10082), .ZN(n14855) );
  NAND2_X1 U12624 ( .A1(n14855), .A2(n14540), .ZN(n14899) );
  INV_X1 U12625 ( .A(n14899), .ZN(n14193) );
  INV_X1 U12626 ( .A(n10085), .ZN(n10089) );
  NAND2_X1 U12627 ( .A1(n6609), .A2(n12112), .ZN(n10088) );
  INV_X1 U12628 ( .A(n10367), .ZN(n10086) );
  NAND2_X1 U12629 ( .A1(n10086), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10087) );
  OAI211_X1 U12630 ( .C1(n10243), .C2(n10098), .A(n10088), .B(n10087), .ZN(
        n10251) );
  OAI21_X1 U12631 ( .B1(n10089), .B2(n10251), .A(n10250), .ZN(n10090) );
  INV_X1 U12632 ( .A(n10090), .ZN(n14254) );
  INV_X1 U12633 ( .A(n10091), .ZN(n10094) );
  NOR2_X1 U12634 ( .A1(n14963), .A2(n10092), .ZN(n10093) );
  NAND2_X1 U12635 ( .A1(n14844), .A2(n10365), .ZN(n14126) );
  NAND2_X1 U12636 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n14126), .ZN(n10095) );
  OAI21_X1 U12637 ( .B1(n14254), .B2(n14850), .A(n10095), .ZN(n10096) );
  AOI21_X1 U12638 ( .B1(n14193), .B2(n10246), .A(n10096), .ZN(n10097) );
  OAI21_X1 U12639 ( .B1(n10098), .B2(n14896), .A(n10097), .ZN(P1_U3232) );
  OAI21_X1 U12640 ( .B1(n10101), .B2(n10100), .A(n10099), .ZN(n10113) );
  INV_X1 U12641 ( .A(n10102), .ZN(n10104) );
  NAND3_X1 U12642 ( .A1(n10104), .A2(n10103), .A3(n10150), .ZN(n10105) );
  AOI21_X1 U12643 ( .B1(n15220), .B2(n10105), .A(n15322), .ZN(n10112) );
  AOI21_X1 U12644 ( .B1(n10108), .B2(n10107), .A(n10106), .ZN(n10110) );
  AOI22_X1 U12645 ( .A1(n15326), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10109) );
  OAI21_X1 U12646 ( .B1(n15297), .B2(n10110), .A(n10109), .ZN(n10111) );
  AOI211_X1 U12647 ( .C1(n15264), .C2(n10113), .A(n10112), .B(n10111), .ZN(
        n10114) );
  OAI21_X1 U12648 ( .B1(n10115), .B2(n15320), .A(n10114), .ZN(P3_U3184) );
  INV_X1 U12649 ( .A(n11583), .ZN(n10192) );
  INV_X1 U12650 ( .A(n12137), .ZN(n14666) );
  AOI22_X1 U12651 ( .A1(n14297), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n14666), .ZN(n10116) );
  OAI21_X1 U12652 ( .B1(n10192), .B2(n14668), .A(n10116), .ZN(P1_U3339) );
  NAND2_X1 U12653 ( .A1(n10118), .A2(n10117), .ZN(n10121) );
  AOI22_X1 U12654 ( .A1(n6613), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n12733), 
        .B2(n10119), .ZN(n10120) );
  INV_X1 U12655 ( .A(n15106), .ZN(n13958) );
  INV_X1 U12656 ( .A(n10122), .ZN(n10124) );
  AND2_X1 U12657 ( .A1(n13274), .A2(n6611), .ZN(n10128) );
  XNOR2_X1 U12658 ( .A(n12895), .B(n15106), .ZN(n10127) );
  NOR2_X1 U12659 ( .A1(n10127), .A2(n10128), .ZN(n10265) );
  AOI21_X1 U12660 ( .B1(n10128), .B2(n10127), .A(n10265), .ZN(n10129) );
  NAND2_X1 U12661 ( .A1(n10130), .A2(n10129), .ZN(n10267) );
  OAI21_X1 U12662 ( .B1(n10130), .B2(n10129), .A(n10267), .ZN(n10131) );
  INV_X1 U12663 ( .A(n12967), .ZN(n14793) );
  NAND2_X1 U12664 ( .A1(n10131), .A2(n14793), .ZN(n10145) );
  INV_X1 U12665 ( .A(n13956), .ZN(n10143) );
  INV_X1 U12666 ( .A(n14799), .ZN(n11786) );
  NAND2_X1 U12667 ( .A1(n10406), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n10139) );
  OR2_X1 U12668 ( .A1(n10407), .A2(n10392), .ZN(n10138) );
  INV_X1 U12669 ( .A(n10271), .ZN(n10273) );
  NAND2_X1 U12670 ( .A1(n10133), .A2(n10132), .ZN(n10134) );
  NAND2_X1 U12671 ( .A1(n10273), .A2(n10134), .ZN(n10395) );
  OR2_X1 U12672 ( .A1(n10135), .A2(n10395), .ZN(n10137) );
  OR2_X1 U12673 ( .A1(n12775), .A2(n15165), .ZN(n10136) );
  INV_X1 U12674 ( .A(n13950), .ZN(n10519) );
  OAI22_X1 U12675 ( .A1(n10140), .A2(n12963), .B1(n12962), .B2(n10519), .ZN(
        n10141) );
  AOI211_X1 U12676 ( .C1(n10143), .C2(n11786), .A(n10142), .B(n10141), .ZN(
        n10144) );
  OAI211_X1 U12677 ( .C1(n13958), .C2(n11848), .A(n10145), .B(n10144), .ZN(
        P2_U3202) );
  OAI21_X1 U12678 ( .B1(P3_REG1_REG_1__SCAN_IN), .B2(n10147), .A(n10146), .ZN(
        n10160) );
  INV_X1 U12679 ( .A(n10148), .ZN(n10152) );
  INV_X1 U12680 ( .A(n10149), .ZN(n10151) );
  OAI21_X1 U12681 ( .B1(n10152), .B2(n10151), .A(n10150), .ZN(n10153) );
  AOI22_X1 U12682 ( .A1(n15305), .A2(n10153), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(P3_U3151), .ZN(n10154) );
  OAI21_X1 U12683 ( .B1(n15308), .B2(n13672), .A(n10154), .ZN(n10159) );
  NAND2_X1 U12684 ( .A1(n10155), .A2(n10012), .ZN(n10156) );
  AOI21_X1 U12685 ( .B1(n10157), .B2(n10156), .A(n15333), .ZN(n10158) );
  AOI211_X1 U12686 ( .C1(n15329), .C2(n10160), .A(n10159), .B(n10158), .ZN(
        n10161) );
  OAI21_X1 U12687 ( .B1(n10162), .B2(n15320), .A(n10161), .ZN(P3_U3183) );
  AND3_X1 U12688 ( .A1(n10164), .A2(n10193), .A3(n10163), .ZN(n10167) );
  INV_X1 U12689 ( .A(n10165), .ZN(n10166) );
  AND2_X1 U12690 ( .A1(n10166), .A2(n15082), .ZN(n15083) );
  AND2_X1 U12691 ( .A1(n10167), .A2(n15083), .ZN(n10183) );
  AND2_X2 U12692 ( .A1(n10183), .A2(n15081), .ZN(n15157) );
  INV_X1 U12693 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10181) );
  INV_X1 U12694 ( .A(n10471), .ZN(n10169) );
  AOI21_X1 U12695 ( .B1(n10170), .B2(n13183), .A(n10169), .ZN(n10178) );
  INV_X1 U12696 ( .A(n10178), .ZN(n10500) );
  NAND2_X1 U12697 ( .A1(n9993), .A2(n12976), .ZN(n10475) );
  OAI211_X1 U12698 ( .C1(n9993), .C2(n12976), .A(n15065), .B(n10475), .ZN(
        n10495) );
  OAI21_X1 U12699 ( .B1(n9993), .B2(n15150), .A(n10495), .ZN(n10179) );
  AOI22_X1 U12700 ( .A1(n14787), .A2(n10172), .B1(n13949), .B2(n10319), .ZN(
        n10177) );
  OAI21_X1 U12701 ( .B1(n10173), .B2(n13183), .A(n10325), .ZN(n10175) );
  OR2_X1 U12702 ( .A1(n10168), .A2(n13331), .ZN(n10174) );
  NAND2_X1 U12703 ( .A1(n6610), .A2(n13184), .ZN(n13219) );
  NAND2_X1 U12704 ( .A1(n10175), .A2(n15054), .ZN(n10176) );
  OAI211_X1 U12705 ( .C1(n10178), .C2(n10171), .A(n10177), .B(n10176), .ZN(
        n10494) );
  AOI211_X1 U12706 ( .C1(n12969), .C2(n10500), .A(n10179), .B(n10494), .ZN(
        n10184) );
  OR2_X1 U12707 ( .A1(n10184), .A2(n15156), .ZN(n10180) );
  OAI21_X1 U12708 ( .B1(n15157), .B2(n10181), .A(n10180), .ZN(P2_U3433) );
  AND2_X2 U12709 ( .A1(n10183), .A2(n10182), .ZN(n15177) );
  OR2_X1 U12710 ( .A1(n10184), .A2(n15174), .ZN(n10185) );
  OAI21_X1 U12711 ( .B1(n15177), .B2(n10186), .A(n10185), .ZN(P2_U3500) );
  NAND2_X1 U12712 ( .A1(n15215), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10353) );
  NAND2_X1 U12713 ( .A1(n10353), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10189) );
  INV_X1 U12714 ( .A(n12224), .ZN(n12169) );
  AOI22_X1 U12715 ( .A1(n15213), .A2(n10187), .B1(n12169), .B2(n12244), .ZN(
        n10188) );
  OAI211_X1 U12716 ( .C1(n10907), .C2(n15207), .A(n10189), .B(n10188), .ZN(
        P3_U3172) );
  XNOR2_X1 U12717 ( .A(n10191), .B(n10190), .ZN(n15050) );
  OAI222_X1 U12718 ( .A1(P2_U3088), .A2(n15050), .B1(n6618), .B2(n10192), .C1(
        n13518), .C2(n11987), .ZN(P2_U3311) );
  NAND4_X1 U12719 ( .A1(n10194), .A2(n10193), .A3(n15082), .A4(n15081), .ZN(
        n10195) );
  NAND2_X1 U12720 ( .A1(n6610), .A2(n13174), .ZN(n10376) );
  INV_X1 U12721 ( .A(n10376), .ZN(n10196) );
  NAND2_X1 U12722 ( .A1(n13944), .A2(n10196), .ZN(n10900) );
  INV_X1 U12723 ( .A(n10171), .ZN(n15155) );
  NOR2_X1 U12724 ( .A1(n15155), .A2(n15054), .ZN(n10197) );
  OAI22_X1 U12725 ( .A1(n10197), .A2(n15086), .B1(n10324), .B2(n14784), .ZN(
        n15088) );
  NAND2_X1 U12726 ( .A1(n10198), .A2(n12973), .ZN(n15087) );
  OAI22_X1 U12727 ( .A1(n13957), .A2(n10199), .B1(n15087), .B2(n13174), .ZN(
        n10200) );
  OAI21_X1 U12728 ( .B1(n15088), .B2(n10200), .A(n13944), .ZN(n10202) );
  NAND2_X1 U12729 ( .A1(n15059), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n10201) );
  OAI211_X1 U12730 ( .C1(n15086), .C2(n10900), .A(n10202), .B(n10201), .ZN(
        P2_U3265) );
  INV_X1 U12731 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10205) );
  INV_X1 U12732 ( .A(n11538), .ZN(n10206) );
  NAND2_X1 U12733 ( .A1(n10283), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10203) );
  XNOR2_X1 U12734 ( .A(n10203), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11539) );
  INV_X1 U12735 ( .A(n11539), .ZN(n10204) );
  OAI222_X1 U12736 ( .A1(n11987), .A2(n10205), .B1(n6618), .B2(n10206), .C1(
        P2_U3088), .C2(n10204), .ZN(P2_U3313) );
  INV_X1 U12737 ( .A(n11644), .ZN(n11213) );
  OAI222_X1 U12738 ( .A1(n12137), .A2(n10207), .B1(n14668), .B2(n10206), .C1(
        P1_U3086), .C2(n11213), .ZN(P1_U3341) );
  INV_X1 U12739 ( .A(n10353), .ZN(n10219) );
  INV_X1 U12740 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10218) );
  INV_X1 U12741 ( .A(n8135), .ZN(n10210) );
  OAI211_X1 U12742 ( .C1(n10212), .C2(n15368), .A(n10208), .B(n10211), .ZN(
        n10213) );
  NAND2_X1 U12743 ( .A1(n10213), .A2(n15193), .ZN(n10217) );
  OAI22_X1 U12744 ( .A1(n12230), .A2(n10214), .B1(n12224), .B2(n10435), .ZN(
        n10215) );
  AOI21_X1 U12745 ( .B1(n12212), .B2(n15367), .A(n10215), .ZN(n10216) );
  OAI211_X1 U12746 ( .C1(n10219), .C2(n10218), .A(n10217), .B(n10216), .ZN(
        P3_U3162) );
  INV_X1 U12747 ( .A(n10220), .ZN(n10222) );
  AOI21_X1 U12748 ( .B1(n10223), .B2(n10222), .A(n10221), .ZN(n10228) );
  INV_X1 U12749 ( .A(n10363), .ZN(n10225) );
  NAND4_X1 U12750 ( .A1(n10225), .A2(n10224), .A3(n10364), .A4(n10365), .ZN(
        n10226) );
  INV_X1 U12751 ( .A(n14498), .ZN(n14703) );
  AOI22_X1 U12752 ( .A1(n14705), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n14703), .ZN(n10227) );
  OAI21_X1 U12753 ( .B1(n10228), .B2(n14705), .A(n10227), .ZN(P1_U3293) );
  INV_X1 U12754 ( .A(n11739), .ZN(n10346) );
  AOI22_X1 U12755 ( .A1(n14310), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n14666), .ZN(n10229) );
  OAI21_X1 U12756 ( .B1(n10346), .B2(n14668), .A(n10229), .ZN(P1_U3338) );
  OAI21_X1 U12757 ( .B1(n10231), .B2(n10232), .A(n10230), .ZN(n10238) );
  OAI22_X1 U12758 ( .A1(n8910), .A2(n14438), .B1(n10743), .B2(n14466), .ZN(
        n10237) );
  NAND2_X1 U12759 ( .A1(n10233), .A2(n10232), .ZN(n10234) );
  AOI21_X1 U12760 ( .B1(n10235), .B2(n10234), .A(n14603), .ZN(n10236) );
  AOI211_X1 U12761 ( .C1(n14965), .C2(n10238), .A(n10237), .B(n10236), .ZN(
        n10591) );
  OAI211_X1 U12762 ( .C1(n11129), .C2(n10594), .A(n10825), .B(n14712), .ZN(
        n10598) );
  OAI211_X1 U12763 ( .C1(n10594), .C2(n14947), .A(n10591), .B(n10598), .ZN(
        n10240) );
  NAND2_X1 U12764 ( .A1(n10240), .A2(n14982), .ZN(n10239) );
  OAI21_X1 U12765 ( .B1(n14982), .B2(n9442), .A(n10239), .ZN(P1_U3530) );
  INV_X1 U12766 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10242) );
  NAND2_X1 U12767 ( .A1(n10240), .A2(n14973), .ZN(n10241) );
  OAI21_X1 U12768 ( .B1(n14973), .B2(n10242), .A(n10241), .ZN(P1_U3465) );
  AOI22_X1 U12769 ( .A1(n12119), .A2(n14251), .B1(n12073), .B2(n10255), .ZN(
        n10356) );
  AOI22_X1 U12770 ( .A1(n14251), .A2(n12073), .B1(n12120), .B2(n10255), .ZN(
        n10244) );
  XNOR2_X1 U12771 ( .A(n10244), .B(n10932), .ZN(n10357) );
  XOR2_X1 U12772 ( .A(n10356), .B(n10357), .Z(n10358) );
  XNOR2_X1 U12773 ( .A(n10247), .B(n10932), .ZN(n10249) );
  INV_X1 U12774 ( .A(n10249), .ZN(n10253) );
  XNOR2_X1 U12775 ( .A(n10254), .B(n10249), .ZN(n14123) );
  OAI21_X1 U12776 ( .B1(n10252), .B2(n10251), .A(n10250), .ZN(n14122) );
  NAND2_X1 U12777 ( .A1(n14123), .A2(n14122), .ZN(n14121) );
  OAI21_X1 U12778 ( .B1(n10254), .B2(n10253), .A(n14121), .ZN(n10359) );
  XOR2_X1 U12779 ( .A(n10358), .B(n10359), .Z(n10258) );
  NAND2_X1 U12780 ( .A1(n14855), .A2(n14539), .ZN(n14900) );
  INV_X1 U12781 ( .A(n14900), .ZN(n14194) );
  AOI22_X1 U12782 ( .A1(n14194), .A2(n10246), .B1(n14215), .B2(n10255), .ZN(
        n10257) );
  AOI22_X1 U12783 ( .A1(n14193), .A2(n14250), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n14126), .ZN(n10256) );
  OAI211_X1 U12784 ( .C1(n10258), .C2(n14850), .A(n10257), .B(n10256), .ZN(
        P1_U3237) );
  NAND2_X1 U12785 ( .A1(n10259), .A2(n10117), .ZN(n10262) );
  AOI22_X1 U12786 ( .A1(n6613), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n12733), 
        .B2(n10260), .ZN(n10261) );
  NAND2_X2 U12787 ( .A1(n10262), .A2(n10261), .ZN(n15113) );
  INV_X1 U12788 ( .A(n15113), .ZN(n10396) );
  AND2_X1 U12789 ( .A1(n13950), .A2(n12855), .ZN(n10264) );
  XNOR2_X1 U12790 ( .A(n15113), .B(n12895), .ZN(n10263) );
  NOR2_X1 U12791 ( .A1(n10263), .A2(n10264), .ZN(n10400) );
  AOI21_X1 U12792 ( .B1(n10264), .B2(n10263), .A(n10400), .ZN(n10269) );
  INV_X1 U12793 ( .A(n10265), .ZN(n10266) );
  NAND2_X1 U12794 ( .A1(n10267), .A2(n10266), .ZN(n10268) );
  OAI21_X1 U12795 ( .B1(n10269), .B2(n10268), .A(n10402), .ZN(n10270) );
  NAND2_X1 U12796 ( .A1(n10270), .A2(n14793), .ZN(n10282) );
  NAND2_X1 U12797 ( .A1(n10406), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n10278) );
  OR2_X1 U12798 ( .A1(n10407), .A2(n10525), .ZN(n10277) );
  INV_X1 U12799 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10272) );
  NAND2_X1 U12800 ( .A1(n10273), .A2(n10272), .ZN(n10274) );
  NAND2_X1 U12801 ( .A1(n10410), .A2(n10274), .ZN(n10529) );
  OR2_X1 U12802 ( .A1(n10135), .A2(n10529), .ZN(n10276) );
  OR2_X1 U12803 ( .A1(n12775), .A2(n15167), .ZN(n10275) );
  INV_X1 U12804 ( .A(n13272), .ZN(n10586) );
  OAI22_X1 U12805 ( .A1(n10388), .A2(n13928), .B1(n10586), .B2(n14784), .ZN(
        n10390) );
  NOR2_X1 U12806 ( .A1(n14799), .A2(n10395), .ZN(n10279) );
  AOI211_X1 U12807 ( .C1(n14795), .C2(n10390), .A(n10280), .B(n10279), .ZN(
        n10281) );
  OAI211_X1 U12808 ( .C1(n10396), .C2(n11848), .A(n10282), .B(n10281), .ZN(
        P2_U3199) );
  INV_X1 U12809 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10285) );
  INV_X1 U12810 ( .A(n11542), .ZN(n10347) );
  OAI21_X1 U12811 ( .B1(n10283), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n10284) );
  XNOR2_X1 U12812 ( .A(n10284), .B(P2_IR_REG_15__SCAN_IN), .ZN(n13296) );
  INV_X1 U12813 ( .A(n13296), .ZN(n11497) );
  OAI222_X1 U12814 ( .A1(n11987), .A2(n10285), .B1(n6618), .B2(n10347), .C1(
        P2_U3088), .C2(n11497), .ZN(P2_U3312) );
  INV_X1 U12815 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10286) );
  MUX2_X1 U12816 ( .A(n10286), .B(P1_REG1_REG_10__SCAN_IN), .S(n10553), .Z(
        n10289) );
  OAI21_X1 U12817 ( .B1(n10290), .B2(P1_REG1_REG_9__SCAN_IN), .A(n10287), .ZN(
        n10288) );
  NOR2_X1 U12818 ( .A1(n10288), .A2(n10289), .ZN(n10552) );
  AOI211_X1 U12819 ( .C1(n10289), .C2(n10288), .A(n14298), .B(n10552), .ZN(
        n10301) );
  NAND2_X1 U12820 ( .A1(n10290), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10294) );
  INV_X1 U12821 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10291) );
  MUX2_X1 U12822 ( .A(n10291), .B(P1_REG2_REG_10__SCAN_IN), .S(n10553), .Z(
        n10293) );
  NAND3_X1 U12823 ( .A1(n10295), .A2(n10294), .A3(n10293), .ZN(n10292) );
  NAND2_X1 U12824 ( .A1(n14332), .A2(n10292), .ZN(n10299) );
  AOI21_X1 U12825 ( .B1(n10295), .B2(n10294), .A(n10293), .ZN(n10551) );
  AND2_X1 U12826 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n11683) );
  AOI21_X1 U12827 ( .B1(n14316), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n11683), 
        .ZN(n10298) );
  OR2_X1 U12828 ( .A1(n14921), .A2(n10296), .ZN(n10297) );
  OAI211_X1 U12829 ( .C1(n10299), .C2(n10551), .A(n10298), .B(n10297), .ZN(
        n10300) );
  OR2_X1 U12830 ( .A1(n10301), .A2(n10300), .ZN(P1_U3253) );
  NAND2_X1 U12831 ( .A1(n11359), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n10603) );
  OAI21_X1 U12832 ( .B1(n11359), .B2(P2_REG2_REG_13__SCAN_IN), .A(n10603), 
        .ZN(n10599) );
  INV_X1 U12833 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n10304) );
  NAND2_X1 U12834 ( .A1(n10309), .A2(n10302), .ZN(n15023) );
  MUX2_X1 U12835 ( .A(n10304), .B(P2_REG2_REG_12__SCAN_IN), .S(n15031), .Z(
        n15024) );
  AOI21_X1 U12836 ( .B1(n15025), .B2(n15023), .A(n15024), .ZN(n15022) );
  AOI21_X1 U12837 ( .B1(n10304), .B2(n10303), .A(n15022), .ZN(n10601) );
  XOR2_X1 U12838 ( .A(n10599), .B(n10601), .Z(n10315) );
  INV_X1 U12839 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n11310) );
  NOR2_X1 U12840 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11310), .ZN(n10305) );
  AOI21_X1 U12841 ( .B1(n15043), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n10305), 
        .ZN(n10306) );
  INV_X1 U12842 ( .A(n10306), .ZN(n10313) );
  INV_X1 U12843 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n14829) );
  NOR2_X1 U12844 ( .A1(n11359), .A2(n14829), .ZN(n10307) );
  AOI21_X1 U12845 ( .B1(n11359), .B2(n14829), .A(n10307), .ZN(n10311) );
  OAI21_X1 U12846 ( .B1(n15175), .B2(n10309), .A(n10308), .ZN(n15019) );
  INV_X1 U12847 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n14836) );
  MUX2_X1 U12848 ( .A(n14836), .B(P2_REG1_REG_12__SCAN_IN), .S(n15031), .Z(
        n15018) );
  OAI21_X1 U12849 ( .B1(n15031), .B2(P2_REG1_REG_12__SCAN_IN), .A(n15021), 
        .ZN(n10310) );
  NOR2_X1 U12850 ( .A1(n10310), .A2(n10311), .ZN(n10605) );
  AOI211_X1 U12851 ( .C1(n10311), .C2(n10310), .A(n15037), .B(n10605), .ZN(
        n10312) );
  AOI211_X1 U12852 ( .C1(n15032), .C2(n11359), .A(n10313), .B(n10312), .ZN(
        n10314) );
  OAI21_X1 U12853 ( .B1(n15026), .B2(n10315), .A(n10314), .ZN(P2_U3227) );
  OR2_X1 U12854 ( .A1(n13948), .A2(n15100), .ZN(n10386) );
  NAND2_X1 U12855 ( .A1(n13948), .A2(n15100), .ZN(n10316) );
  NAND2_X1 U12856 ( .A1(n10386), .A2(n10316), .ZN(n13186) );
  NAND2_X1 U12857 ( .A1(n10324), .A2(n9993), .ZN(n10470) );
  OR2_X1 U12858 ( .A1(n10319), .A2(n10317), .ZN(n10321) );
  AND2_X1 U12859 ( .A1(n10470), .A2(n10321), .ZN(n10318) );
  NAND2_X1 U12860 ( .A1(n10471), .A2(n10318), .ZN(n10323) );
  OR2_X1 U12861 ( .A1(n10319), .A2(n15093), .ZN(n10329) );
  NAND2_X1 U12862 ( .A1(n10319), .A2(n15093), .ZN(n10320) );
  AND2_X2 U12863 ( .A1(n10329), .A2(n10320), .ZN(n13185) );
  AND2_X1 U12864 ( .A1(n10323), .A2(n10322), .ZN(n10379) );
  XNOR2_X1 U12865 ( .A(n10379), .B(n10327), .ZN(n15098) );
  AOI22_X1 U12866 ( .A1(n14787), .A2(n10319), .B1(n13949), .B2(n13274), .ZN(
        n10333) );
  NAND2_X1 U12867 ( .A1(n10324), .A2(n12979), .ZN(n10465) );
  NAND2_X1 U12868 ( .A1(n10326), .A2(n13185), .ZN(n10328) );
  INV_X1 U12869 ( .A(n10387), .ZN(n10331) );
  AND3_X1 U12870 ( .A1(n13186), .A2(n10329), .A3(n10328), .ZN(n10330) );
  OAI21_X1 U12871 ( .B1(n10331), .B2(n10330), .A(n15054), .ZN(n10332) );
  OAI211_X1 U12872 ( .C1(n15098), .C2(n10171), .A(n10333), .B(n10332), .ZN(
        n15101) );
  INV_X1 U12873 ( .A(n15101), .ZN(n10335) );
  MUX2_X1 U12874 ( .A(n10335), .B(n10334), .S(n15059), .Z(n10341) );
  NAND2_X1 U12875 ( .A1(n13944), .A2(n13331), .ZN(n13937) );
  OR2_X1 U12876 ( .A1(n10475), .A2(n10317), .ZN(n10476) );
  INV_X1 U12877 ( .A(n10476), .ZN(n10336) );
  INV_X1 U12878 ( .A(n10393), .ZN(n13955) );
  OAI211_X1 U12879 ( .C1(n15100), .C2(n10336), .A(n13955), .B(n11374), .ZN(
        n15099) );
  INV_X1 U12880 ( .A(n15099), .ZN(n10339) );
  NAND2_X1 U12881 ( .A1(n13944), .A2(n10337), .ZN(n13959) );
  OAI22_X1 U12882 ( .A1(n13959), .A2(n15100), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n13957), .ZN(n10338) );
  AOI21_X1 U12883 ( .B1(n15068), .B2(n10339), .A(n10338), .ZN(n10340) );
  OAI211_X1 U12884 ( .C1(n15098), .C2(n10900), .A(n10341), .B(n10340), .ZN(
        P2_U3262) );
  NAND2_X1 U12885 ( .A1(n10342), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10343) );
  MUX2_X1 U12886 ( .A(n10343), .B(P2_IR_REG_31__SCAN_IN), .S(n13636), .Z(
        n10344) );
  NAND2_X1 U12887 ( .A1(n10344), .A2(n9613), .ZN(n13310) );
  OAI222_X1 U12888 ( .A1(P2_U3088), .A2(n13310), .B1(n6618), .B2(n10346), .C1(
        n10345), .C2(n11987), .ZN(P2_U3310) );
  INV_X1 U12889 ( .A(n11646), .ZN(n14922) );
  OAI222_X1 U12890 ( .A1(n10348), .A2(n12137), .B1(P1_U3086), .B2(n14922), 
        .C1(n14668), .C2(n10347), .ZN(P1_U3340) );
  XOR2_X1 U12891 ( .A(n10350), .B(n10349), .Z(n10355) );
  AOI22_X1 U12892 ( .A1(n15213), .A2(n7649), .B1(n12169), .B2(n12243), .ZN(
        n10351) );
  OAI21_X1 U12893 ( .B1(n6846), .B2(n12222), .A(n10351), .ZN(n10352) );
  AOI21_X1 U12894 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n10353), .A(n10352), .ZN(
        n10354) );
  OAI21_X1 U12895 ( .B1(n10355), .B2(n15207), .A(n10354), .ZN(P3_U3177) );
  AOI22_X1 U12896 ( .A1(n10359), .A2(n10358), .B1(n10357), .B2(n10356), .ZN(
        n10362) );
  AOI22_X1 U12897 ( .A1(n12119), .A2(n14250), .B1(n12073), .B2(n14939), .ZN(
        n10737) );
  AOI22_X1 U12898 ( .A1(n14250), .A2(n12054), .B1(n12120), .B2(n14939), .ZN(
        n10360) );
  XNOR2_X1 U12899 ( .A(n10360), .B(n10932), .ZN(n10736) );
  XOR2_X1 U12900 ( .A(n10737), .B(n10736), .Z(n10361) );
  NAND2_X1 U12901 ( .A1(n10362), .A2(n10361), .ZN(n10735) );
  OAI211_X1 U12902 ( .C1(n10362), .C2(n10361), .A(n10735), .B(n14904), .ZN(
        n10375) );
  OR2_X1 U12903 ( .A1(n10364), .A2(n10363), .ZN(n10370) );
  NAND3_X1 U12904 ( .A1(n10367), .A2(n10366), .A3(n10365), .ZN(n10368) );
  AOI21_X1 U12905 ( .B1(n10370), .B2(n10369), .A(n10368), .ZN(n10371) );
  INV_X1 U12906 ( .A(n14909), .ZN(n14228) );
  MUX2_X1 U12907 ( .A(n14228), .B(P1_U3086), .S(P1_REG3_REG_3__SCAN_IN), .Z(
        n10373) );
  OAI22_X1 U12908 ( .A1(n14896), .A2(n7099), .B1(n14900), .B2(n11135), .ZN(
        n10372) );
  AOI211_X1 U12909 ( .C1(n14193), .C2(n14249), .A(n10373), .B(n10372), .ZN(
        n10374) );
  NAND2_X1 U12910 ( .A1(n10375), .A2(n10374), .ZN(P1_U3218) );
  NAND2_X1 U12911 ( .A1(n10171), .A2(n10376), .ZN(n10377) );
  NAND2_X1 U12912 ( .A1(n13944), .A2(n10377), .ZN(n13941) );
  NAND2_X1 U12913 ( .A1(n13948), .A2(n12988), .ZN(n10378) );
  NAND2_X1 U12914 ( .A1(n10379), .A2(n10378), .ZN(n10381) );
  OR2_X1 U12915 ( .A1(n13948), .A2(n12988), .ZN(n10380) );
  NAND2_X1 U12916 ( .A1(n10381), .A2(n10380), .ZN(n10516) );
  OR2_X1 U12917 ( .A1(n13962), .A2(n13961), .ZN(n15108) );
  NAND2_X1 U12918 ( .A1(n15106), .A2(n13274), .ZN(n10382) );
  NAND2_X1 U12919 ( .A1(n15108), .A2(n10382), .ZN(n10385) );
  INV_X1 U12920 ( .A(n13190), .ZN(n10384) );
  OR2_X1 U12921 ( .A1(n13961), .A2(n13190), .ZN(n10513) );
  OR2_X1 U12922 ( .A1(n13962), .A2(n10513), .ZN(n10509) );
  AND2_X1 U12923 ( .A1(n10508), .A2(n10509), .ZN(n10383) );
  OAI21_X1 U12924 ( .B1(n10385), .B2(n10384), .A(n10383), .ZN(n15118) );
  NAND2_X1 U12925 ( .A1(n10388), .A2(n15106), .ZN(n10389) );
  XNOR2_X1 U12926 ( .A(n13190), .B(n10522), .ZN(n10391) );
  AOI21_X1 U12927 ( .B1(n10391), .B2(n15054), .A(n10390), .ZN(n15116) );
  MUX2_X1 U12928 ( .A(n10392), .B(n15116), .S(n13944), .Z(n10399) );
  NAND2_X1 U12929 ( .A1(n10393), .A2(n13958), .ZN(n13953) );
  OR2_X1 U12930 ( .A1(n13953), .A2(n15113), .ZN(n10527) );
  INV_X1 U12931 ( .A(n10527), .ZN(n10394) );
  AOI211_X1 U12932 ( .C1(n15113), .C2(n13953), .A(n6611), .B(n10394), .ZN(
        n15112) );
  OAI22_X1 U12933 ( .A1(n13959), .A2(n10396), .B1(n13957), .B2(n10395), .ZN(
        n10397) );
  AOI21_X1 U12934 ( .B1(n15112), .B2(n15068), .A(n10397), .ZN(n10398) );
  OAI211_X1 U12935 ( .C1(n13941), .C2(n15118), .A(n10399), .B(n10398), .ZN(
        P2_U3260) );
  INV_X1 U12936 ( .A(n10400), .ZN(n10401) );
  NAND2_X1 U12937 ( .A1(n13272), .A2(n12855), .ZN(n10571) );
  AOI22_X1 U12938 ( .A1(n6613), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n12733), 
        .B2(n13276), .ZN(n10404) );
  XNOR2_X1 U12939 ( .A(n13009), .B(n12895), .ZN(n10570) );
  XOR2_X1 U12940 ( .A(n10571), .B(n10570), .Z(n10572) );
  XNOR2_X1 U12941 ( .A(n10573), .B(n10572), .ZN(n10422) );
  NAND2_X1 U12942 ( .A1(n14787), .A2(n13950), .ZN(n10418) );
  NAND2_X1 U12943 ( .A1(n13169), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n10416) );
  OR2_X1 U12944 ( .A1(n13172), .A2(n10408), .ZN(n10415) );
  NAND2_X1 U12945 ( .A1(n10410), .A2(n10409), .ZN(n10411) );
  NAND2_X1 U12946 ( .A1(n10580), .A2(n10411), .ZN(n10694) );
  OR2_X1 U12947 ( .A1(n12901), .A2(n10694), .ZN(n10414) );
  OR2_X1 U12948 ( .A1(n12903), .A2(n10412), .ZN(n10413) );
  NAND4_X1 U12949 ( .A1(n10416), .A2(n10415), .A3(n10414), .A4(n10413), .ZN(
        n13271) );
  NAND2_X1 U12950 ( .A1(n13949), .A2(n13271), .ZN(n10417) );
  NAND2_X1 U12951 ( .A1(n10418), .A2(n10417), .ZN(n10523) );
  NAND2_X1 U12952 ( .A1(n14795), .A2(n10523), .ZN(n10419) );
  NAND2_X1 U12953 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n13285) );
  OAI211_X1 U12954 ( .C1(n14799), .C2(n10529), .A(n10419), .B(n13285), .ZN(
        n10420) );
  AOI21_X1 U12955 ( .B1(n13009), .B2(n14796), .A(n10420), .ZN(n10421) );
  OAI21_X1 U12956 ( .B1(n10422), .B2(n12967), .A(n10421), .ZN(P2_U3211) );
  AND2_X1 U12957 ( .A1(n15374), .A2(n10423), .ZN(n10424) );
  NAND2_X1 U12958 ( .A1(n11263), .A2(n10424), .ZN(n10426) );
  NAND2_X1 U12959 ( .A1(n6687), .A2(n10427), .ZN(n10447) );
  INV_X1 U12960 ( .A(n10447), .ZN(n10425) );
  NAND2_X1 U12961 ( .A1(n10448), .A2(n10425), .ZN(n10457) );
  OR2_X1 U12962 ( .A1(n10428), .A2(n10427), .ZN(n12595) );
  INV_X1 U12963 ( .A(n14775), .ZN(n15413) );
  OAI21_X1 U12964 ( .B1(n10430), .B2(n7214), .A(n10429), .ZN(n10431) );
  INV_X1 U12965 ( .A(n10431), .ZN(n10550) );
  NAND2_X1 U12966 ( .A1(n10433), .A2(n10432), .ZN(n15347) );
  NAND2_X1 U12967 ( .A1(n15347), .A2(n10434), .ZN(n10437) );
  NAND2_X1 U12968 ( .A1(n10435), .A2(n15360), .ZN(n10436) );
  NAND2_X1 U12969 ( .A1(n12243), .A2(n15200), .ZN(n10438) );
  INV_X1 U12970 ( .A(n10443), .ZN(n10441) );
  AOI21_X1 U12971 ( .B1(n10441), .B2(n7214), .A(n15359), .ZN(n10446) );
  NAND2_X1 U12972 ( .A1(n15366), .A2(n12242), .ZN(n10445) );
  OR2_X1 U12973 ( .A1(n15352), .A2(n15353), .ZN(n10444) );
  NAND2_X1 U12974 ( .A1(n10445), .A2(n10444), .ZN(n10488) );
  AOI21_X1 U12975 ( .B1(n10446), .B2(n10723), .A(n10488), .ZN(n10544) );
  OAI21_X1 U12976 ( .B1(n15413), .B2(n10550), .A(n10544), .ZN(n11273) );
  OAI21_X1 U12977 ( .B1(n15374), .B2(n10448), .A(n10447), .ZN(n10450) );
  NAND2_X1 U12978 ( .A1(n10450), .A2(n10449), .ZN(n10451) );
  NAND2_X1 U12979 ( .A1(n10451), .A2(n10458), .ZN(n10452) );
  NAND2_X1 U12980 ( .A1(n10452), .A2(n10535), .ZN(n10461) );
  XNOR2_X1 U12981 ( .A(n10453), .B(n12713), .ZN(n10456) );
  AND2_X1 U12982 ( .A1(n10454), .A2(n10540), .ZN(n10455) );
  NAND2_X1 U12983 ( .A1(n10458), .A2(n10457), .ZN(n10536) );
  NAND2_X1 U12984 ( .A1(n10537), .A2(n10536), .ZN(n10459) );
  NAND2_X1 U12985 ( .A1(n10459), .A2(n12713), .ZN(n10460) );
  NAND2_X1 U12986 ( .A1(n15436), .A2(n14770), .ZN(n12651) );
  OAI22_X1 U12987 ( .A1(n12651), .A2(n10490), .B1(n15436), .B2(n10462), .ZN(
        n10463) );
  AOI21_X1 U12988 ( .B1(n11273), .B2(n15436), .A(n10463), .ZN(n10464) );
  INV_X1 U12989 ( .A(n10464), .ZN(P3_U3463) );
  NAND3_X1 U12990 ( .A1(n10325), .A2(n10473), .A3(n10465), .ZN(n10466) );
  NAND2_X1 U12991 ( .A1(n10328), .A2(n10466), .ZN(n10467) );
  NAND2_X1 U12992 ( .A1(n10467), .A2(n15054), .ZN(n10469) );
  AOI22_X1 U12993 ( .A1(n13275), .A2(n14787), .B1(n13949), .B2(n13948), .ZN(
        n10468) );
  NAND2_X1 U12994 ( .A1(n10469), .A2(n10468), .ZN(n15094) );
  INV_X1 U12995 ( .A(n15094), .ZN(n10483) );
  NAND2_X1 U12996 ( .A1(n10471), .A2(n10470), .ZN(n10474) );
  NAND2_X1 U12997 ( .A1(n10474), .A2(n10473), .ZN(n10472) );
  OAI21_X1 U12998 ( .B1(n10474), .B2(n10473), .A(n10472), .ZN(n15096) );
  INV_X1 U12999 ( .A(n10475), .ZN(n10477) );
  OAI211_X1 U13000 ( .C1(n10477), .C2(n15093), .A(n15065), .B(n10476), .ZN(
        n15092) );
  INV_X1 U13001 ( .A(n13959), .ZN(n15060) );
  OAI22_X1 U13002 ( .A1(n13944), .A2(n9923), .B1(n10478), .B2(n13957), .ZN(
        n10479) );
  AOI21_X1 U13003 ( .B1(n15060), .B2(n10317), .A(n10479), .ZN(n10480) );
  OAI21_X1 U13004 ( .B1(n13937), .B2(n15092), .A(n10480), .ZN(n10481) );
  AOI21_X1 U13005 ( .B1(n15069), .B2(n15096), .A(n10481), .ZN(n10482) );
  OAI21_X1 U13006 ( .B1(n15072), .B2(n10483), .A(n10482), .ZN(P2_U3263) );
  INV_X1 U13007 ( .A(n10484), .ZN(n10485) );
  AOI21_X1 U13008 ( .B1(n10487), .B2(n10486), .A(n10485), .ZN(n10493) );
  INV_X1 U13009 ( .A(n15203), .ZN(n12158) );
  AOI22_X1 U13010 ( .A1(n10488), .A2(n12158), .B1(P3_REG3_REG_4__SCAN_IN), 
        .B2(P3_U3151), .ZN(n10489) );
  OAI21_X1 U13011 ( .B1(n10490), .B2(n12230), .A(n10489), .ZN(n10491) );
  AOI21_X1 U13012 ( .B1(n10547), .B2(n12227), .A(n10491), .ZN(n10492) );
  OAI21_X1 U13013 ( .B1(n10493), .B2(n15207), .A(n10492), .ZN(P3_U3170) );
  INV_X1 U13014 ( .A(n10494), .ZN(n10502) );
  INV_X1 U13015 ( .A(n10900), .ZN(n10499) );
  NOR2_X1 U13016 ( .A1(n13937), .A2(n10495), .ZN(n10498) );
  INV_X1 U13017 ( .A(n13957), .ZN(n15058) );
  AOI22_X1 U13018 ( .A1(n15059), .A2(P2_REG2_REG_1__SCAN_IN), .B1(n15058), 
        .B2(P2_REG3_REG_1__SCAN_IN), .ZN(n10496) );
  OAI21_X1 U13019 ( .B1(n13959), .B2(n9993), .A(n10496), .ZN(n10497) );
  AOI211_X1 U13020 ( .C1(n10500), .C2(n10499), .A(n10498), .B(n10497), .ZN(
        n10501) );
  OAI21_X1 U13021 ( .B1(n10502), .B2(n15072), .A(n10501), .ZN(P2_U3264) );
  INV_X1 U13022 ( .A(n10503), .ZN(n10506) );
  OAI222_X1 U13023 ( .A1(n11991), .A2(n10506), .B1(n12725), .B2(n10505), .C1(
        P3_U3151), .C2(n10504), .ZN(P3_U3275) );
  NAND2_X1 U13024 ( .A1(n15113), .A2(n13950), .ZN(n10507) );
  NAND2_X1 U13025 ( .A1(n10509), .A2(n10511), .ZN(n10510) );
  XNOR2_X2 U13026 ( .A(n13009), .B(n10586), .ZN(n13191) );
  OR2_X1 U13027 ( .A1(n10510), .A2(n13191), .ZN(n10518) );
  NAND2_X1 U13028 ( .A1(n10514), .A2(n13191), .ZN(n10515) );
  OR2_X2 U13029 ( .A1(n10516), .A2(n10515), .ZN(n10691) );
  AND2_X1 U13030 ( .A1(n10688), .A2(n10691), .ZN(n10517) );
  AND2_X1 U13031 ( .A1(n10518), .A2(n10517), .ZN(n15124) );
  INV_X1 U13032 ( .A(n15124), .ZN(n10534) );
  OR2_X1 U13033 ( .A1(n15113), .A2(n10519), .ZN(n10521) );
  AND2_X1 U13034 ( .A1(n15113), .A2(n10519), .ZN(n10520) );
  XNOR2_X1 U13035 ( .A(n10698), .B(n13191), .ZN(n10524) );
  AOI21_X1 U13036 ( .B1(n10524), .B2(n15054), .A(n10523), .ZN(n15126) );
  MUX2_X1 U13037 ( .A(n10525), .B(n15126), .S(n13944), .Z(n10533) );
  NAND2_X1 U13038 ( .A1(n10527), .A2(n13009), .ZN(n10526) );
  NAND2_X1 U13039 ( .A1(n10526), .A2(n15065), .ZN(n10528) );
  OR2_X1 U13040 ( .A1(n10528), .A2(n10692), .ZN(n15121) );
  INV_X1 U13041 ( .A(n15121), .ZN(n10531) );
  INV_X1 U13042 ( .A(n13009), .ZN(n15122) );
  OAI22_X1 U13043 ( .A1(n15122), .A2(n13959), .B1(n13957), .B2(n10529), .ZN(
        n10530) );
  AOI21_X1 U13044 ( .B1(n10531), .B2(n15068), .A(n10530), .ZN(n10532) );
  OAI211_X1 U13045 ( .C1(n13941), .C2(n10534), .A(n10533), .B(n10532), .ZN(
        P2_U3259) );
  XNOR2_X1 U13046 ( .A(n10536), .B(n10535), .ZN(n10539) );
  NAND3_X1 U13047 ( .A1(n10539), .A2(n10538), .A3(n10537), .ZN(n10546) );
  AND2_X1 U13048 ( .A1(n15376), .A2(n10540), .ZN(n10541) );
  NAND2_X1 U13049 ( .A1(n10541), .A2(n14770), .ZN(n12555) );
  NAND2_X1 U13050 ( .A1(n10542), .A2(n15376), .ZN(n15377) );
  NAND2_X1 U13051 ( .A1(n15373), .A2(n15377), .ZN(n10543) );
  INV_X1 U13052 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10545) );
  MUX2_X1 U13053 ( .A(n10545), .B(n10544), .S(n15380), .Z(n10549) );
  NOR2_X1 U13054 ( .A1(n10546), .A2(n15376), .ZN(n15344) );
  NAND2_X1 U13055 ( .A1(n15344), .A2(n14770), .ZN(n12578) );
  INV_X1 U13056 ( .A(n12578), .ZN(n12559) );
  INV_X2 U13057 ( .A(n12555), .ZN(n15379) );
  AOI22_X1 U13058 ( .A1(n12559), .A2(n11274), .B1(n15379), .B2(n10547), .ZN(
        n10548) );
  OAI211_X1 U13059 ( .C1(n10550), .C2(n12563), .A(n10549), .B(n10548), .ZN(
        P3_U3229) );
  AOI21_X1 U13060 ( .B1(n10553), .B2(P1_REG2_REG_10__SCAN_IN), .A(n10551), 
        .ZN(n10706) );
  MUX2_X1 U13061 ( .A(n11395), .B(P1_REG2_REG_11__SCAN_IN), .S(n10712), .Z(
        n10705) );
  XNOR2_X1 U13062 ( .A(n10706), .B(n10705), .ZN(n10562) );
  INV_X1 U13063 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10554) );
  MUX2_X1 U13064 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10554), .S(n10712), .Z(
        n10555) );
  OAI21_X1 U13065 ( .B1(n10556), .B2(n10555), .A(n10711), .ZN(n10557) );
  NAND2_X1 U13066 ( .A1(n10557), .A2(n14913), .ZN(n10561) );
  NOR2_X1 U13067 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14845), .ZN(n10559) );
  NOR2_X1 U13068 ( .A1(n14921), .A2(n10708), .ZN(n10558) );
  AOI211_X1 U13069 ( .C1(n14316), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n10559), 
        .B(n10558), .ZN(n10560) );
  OAI211_X1 U13070 ( .C1(n14917), .C2(n10562), .A(n10561), .B(n10560), .ZN(
        P1_U3254) );
  XOR2_X1 U13071 ( .A(n10564), .B(n10563), .Z(n10569) );
  INV_X1 U13072 ( .A(n10802), .ZN(n11269) );
  OAI22_X1 U13073 ( .A1(n10565), .A2(n15353), .B1(n10858), .B2(n15351), .ZN(
        n10729) );
  AOI22_X1 U13074 ( .A1(n10729), .A2(n12158), .B1(P3_REG3_REG_5__SCAN_IN), 
        .B2(P3_U3151), .ZN(n10566) );
  OAI21_X1 U13075 ( .B1(n11269), .B2(n12230), .A(n10566), .ZN(n10567) );
  AOI21_X1 U13076 ( .B1(n10801), .B2(n12227), .A(n10567), .ZN(n10568) );
  OAI21_X1 U13077 ( .B1(n10569), .B2(n15207), .A(n10568), .ZN(P3_U3167) );
  NAND2_X1 U13078 ( .A1(n10574), .A2(n10117), .ZN(n10577) );
  AOI22_X1 U13079 ( .A1(n12892), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n12733), 
        .B2(n10575), .ZN(n10576) );
  NAND2_X1 U13080 ( .A1(n10577), .A2(n10576), .ZN(n13013) );
  XNOR2_X1 U13081 ( .A(n13013), .B(n12895), .ZN(n10755) );
  NAND2_X1 U13082 ( .A1(n13271), .A2(n12855), .ZN(n10754) );
  XNOR2_X1 U13083 ( .A(n10755), .B(n10754), .ZN(n10757) );
  XNOR2_X1 U13084 ( .A(n10758), .B(n10757), .ZN(n10590) );
  NAND2_X1 U13085 ( .A1(n12900), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10585) );
  INV_X1 U13086 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10578) );
  OR2_X1 U13087 ( .A1(n12845), .A2(n10578), .ZN(n10584) );
  NAND2_X1 U13088 ( .A1(n10580), .A2(n10579), .ZN(n10581) );
  NAND2_X1 U13089 ( .A1(n10766), .A2(n10581), .ZN(n10851) );
  OR2_X1 U13090 ( .A1(n12901), .A2(n10851), .ZN(n10583) );
  OR2_X1 U13091 ( .A1(n12775), .A2(n15170), .ZN(n10582) );
  NAND4_X1 U13092 ( .A1(n10585), .A2(n10584), .A3(n10583), .A4(n10582), .ZN(
        n13270) );
  OAI22_X1 U13093 ( .A1(n10586), .A2(n13928), .B1(n10922), .B2(n14784), .ZN(
        n10699) );
  NAND2_X1 U13094 ( .A1(n10699), .A2(n14795), .ZN(n10587) );
  NAND2_X1 U13095 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n15009) );
  OAI211_X1 U13096 ( .C1(n14799), .C2(n10694), .A(n10587), .B(n15009), .ZN(
        n10588) );
  AOI21_X1 U13097 ( .B1(n13013), .B2(n14796), .A(n10588), .ZN(n10589) );
  OAI21_X1 U13098 ( .B1(n10590), .B2(n12967), .A(n10589), .ZN(P2_U3185) );
  MUX2_X1 U13099 ( .A(n10592), .B(n10591), .S(n14531), .Z(n10597) );
  INV_X1 U13100 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10593) );
  OAI22_X1 U13101 ( .A1(n14506), .A2(n10594), .B1(n14498), .B2(n10593), .ZN(
        n10595) );
  INV_X1 U13102 ( .A(n10595), .ZN(n10596) );
  OAI211_X1 U13103 ( .C1(n14529), .C2(n10598), .A(n10597), .B(n10596), .ZN(
        P1_U3291) );
  INV_X1 U13104 ( .A(n10599), .ZN(n10600) );
  NAND2_X1 U13105 ( .A1(n10601), .A2(n10600), .ZN(n10602) );
  NAND2_X1 U13106 ( .A1(n10603), .A2(n10602), .ZN(n11494) );
  XNOR2_X1 U13107 ( .A(n11539), .B(n11494), .ZN(n10604) );
  NOR2_X1 U13108 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n10604), .ZN(n11495) );
  AOI21_X1 U13109 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n10604), .A(n11495), 
        .ZN(n10612) );
  NAND2_X1 U13110 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14797)
         );
  OAI21_X1 U13111 ( .B1(n15035), .B2(n6928), .A(n14797), .ZN(n10610) );
  AOI21_X1 U13112 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n11359), .A(n10605), 
        .ZN(n10608) );
  INV_X1 U13113 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n14821) );
  NOR2_X1 U13114 ( .A1(n11539), .A2(n14821), .ZN(n10606) );
  AOI21_X1 U13115 ( .B1(n11539), .B2(n14821), .A(n10606), .ZN(n10607) );
  NOR2_X1 U13116 ( .A1(n10608), .A2(n10607), .ZN(n11488) );
  AOI211_X1 U13117 ( .C1(n10608), .C2(n10607), .A(n11488), .B(n15037), .ZN(
        n10609) );
  AOI211_X1 U13118 ( .C1(n15032), .C2(n11539), .A(n10610), .B(n10609), .ZN(
        n10611) );
  OAI21_X1 U13119 ( .B1(n10612), .B2(n15026), .A(n10611), .ZN(P2_U3228) );
  INV_X1 U13120 ( .A(n11867), .ZN(n10615) );
  INV_X1 U13121 ( .A(n14308), .ZN(n14323) );
  OAI222_X1 U13122 ( .A1(n12137), .A2(n10613), .B1(n14668), .B2(n10615), .C1(
        n14323), .C2(P1_U3086), .ZN(P1_U3337) );
  INV_X1 U13123 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10616) );
  NAND2_X1 U13124 ( .A1(n9613), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10614) );
  XNOR2_X1 U13125 ( .A(n10614), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13318) );
  INV_X1 U13126 ( .A(n13318), .ZN(n13322) );
  OAI222_X1 U13127 ( .A1(n11987), .A2(n10616), .B1(n6618), .B2(n10615), .C1(
        n13322), .C2(P2_U3088), .ZN(P2_U3309) );
  NAND2_X1 U13128 ( .A1(n10617), .A2(n10622), .ZN(n10810) );
  INV_X1 U13129 ( .A(n10810), .ZN(n10627) );
  OAI22_X1 U13130 ( .A1(n10743), .A2(n14438), .B1(n10961), .B2(n14466), .ZN(
        n10626) );
  NAND3_X1 U13131 ( .A1(n10829), .A2(n14965), .A3(n10618), .ZN(n10620) );
  NAND2_X1 U13132 ( .A1(n10621), .A2(n14701), .ZN(n10619) );
  NAND2_X1 U13133 ( .A1(n10620), .A2(n10619), .ZN(n10624) );
  NOR2_X1 U13134 ( .A1(n10621), .A2(n14603), .ZN(n10623) );
  MUX2_X1 U13135 ( .A(n10624), .B(n10623), .S(n10622), .Z(n10625) );
  AOI211_X1 U13136 ( .C1(n14965), .C2(n10627), .A(n10626), .B(n10625), .ZN(
        n10793) );
  INV_X1 U13137 ( .A(n10628), .ZN(n10824) );
  INV_X1 U13138 ( .A(n10808), .ZN(n10629) );
  OAI211_X1 U13139 ( .C1(n10794), .C2(n10824), .A(n10629), .B(n14712), .ZN(
        n10792) );
  INV_X1 U13140 ( .A(n10792), .ZN(n10632) );
  AOI22_X1 U13141 ( .A1(n14705), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n10745), 
        .B2(n14703), .ZN(n10630) );
  OAI21_X1 U13142 ( .B1(n14506), .B2(n10794), .A(n10630), .ZN(n10631) );
  AOI21_X1 U13143 ( .B1(n14716), .B2(n10632), .A(n10631), .ZN(n10633) );
  OAI21_X1 U13144 ( .B1(n10793), .B2(n14705), .A(n10633), .ZN(P1_U3289) );
  NOR2_X1 U13145 ( .A1(n11995), .A2(SI_22_), .ZN(n10634) );
  AOI21_X1 U13146 ( .B1(n10635), .B2(P3_STATE_REG_SCAN_IN), .A(n10634), .ZN(
        n10636) );
  OAI21_X1 U13147 ( .B1(n10637), .B2(n11991), .A(n10636), .ZN(n10638) );
  INV_X1 U13148 ( .A(n10638), .ZN(P3_U3273) );
  INV_X1 U13149 ( .A(n15279), .ZN(n10673) );
  NOR2_X1 U13150 ( .A1(n10673), .A2(n10640), .ZN(n10641) );
  INV_X1 U13151 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n15275) );
  NAND2_X1 U13152 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n15296), .ZN(n10642) );
  OAI21_X1 U13153 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n15296), .A(n10642), .ZN(
        n15300) );
  NOR2_X1 U13154 ( .A1(n10676), .A2(n10643), .ZN(n10644) );
  INV_X1 U13155 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n15312) );
  NAND2_X1 U13156 ( .A1(n11058), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n11053) );
  INV_X1 U13157 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11335) );
  NAND2_X1 U13158 ( .A1(n10678), .A2(n11335), .ZN(n10645) );
  NAND2_X1 U13159 ( .A1(n11053), .A2(n10645), .ZN(n10647) );
  INV_X1 U13160 ( .A(n11054), .ZN(n10646) );
  AOI21_X1 U13161 ( .B1(n10648), .B2(n10647), .A(n10646), .ZN(n10686) );
  NAND2_X1 U13162 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n15178)
         );
  OAI21_X1 U13163 ( .B1(n15308), .B2(n10649), .A(n15178), .ZN(n10663) );
  INV_X1 U13164 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n15434) );
  MUX2_X1 U13165 ( .A(P3_REG1_REG_10__SCAN_IN), .B(n15434), .S(n10678), .Z(
        n10660) );
  NAND2_X1 U13166 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n15296), .ZN(n10656) );
  INV_X1 U13167 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15429) );
  AOI22_X1 U13168 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n15296), .B1(n10650), 
        .B2(n15429), .ZN(n15295) );
  NAND2_X1 U13169 ( .A1(P3_REG1_REG_6__SCAN_IN), .A2(n10651), .ZN(n10653) );
  NAND2_X1 U13170 ( .A1(n15279), .A2(n10654), .ZN(n10655) );
  NAND2_X1 U13171 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n15278), .ZN(n15277) );
  NAND2_X1 U13172 ( .A1(n10655), .A2(n15277), .ZN(n15294) );
  NAND2_X1 U13173 ( .A1(n15321), .A2(n10657), .ZN(n10658) );
  XNOR2_X1 U13174 ( .A(n10676), .B(n10657), .ZN(n15328) );
  AOI21_X1 U13175 ( .B1(n10660), .B2(n10659), .A(n11057), .ZN(n10661) );
  NOR2_X1 U13176 ( .A1(n10661), .A2(n15297), .ZN(n10662) );
  AOI211_X1 U13177 ( .C1(n15266), .C2(n10678), .A(n10663), .B(n10662), .ZN(
        n10685) );
  NAND2_X1 U13178 ( .A1(n10665), .A2(n10664), .ZN(n10670) );
  INV_X1 U13179 ( .A(n10666), .ZN(n10668) );
  NAND2_X1 U13180 ( .A1(n10668), .A2(n10667), .ZN(n10669) );
  NAND2_X1 U13181 ( .A1(n10670), .A2(n10669), .ZN(n15283) );
  MUX2_X1 U13182 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n14735), .Z(n10671) );
  XNOR2_X1 U13183 ( .A(n10671), .B(n10673), .ZN(n15282) );
  INV_X1 U13184 ( .A(n10671), .ZN(n10672) );
  MUX2_X1 U13185 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n14735), .Z(n10674) );
  XNOR2_X1 U13186 ( .A(n10674), .B(n15296), .ZN(n15292) );
  OAI22_X1 U13187 ( .A1(n15293), .A2(n15292), .B1(n10674), .B2(n15296), .ZN(
        n15315) );
  MUX2_X1 U13188 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n14735), .Z(n10675) );
  NAND2_X1 U13189 ( .A1(n10675), .A2(n15321), .ZN(n15316) );
  NAND2_X1 U13190 ( .A1(n15315), .A2(n15316), .ZN(n15314) );
  INV_X1 U13191 ( .A(n10675), .ZN(n10677) );
  NAND2_X1 U13192 ( .A1(n10677), .A2(n10676), .ZN(n15318) );
  MUX2_X1 U13193 ( .A(n11335), .B(n15434), .S(n14735), .Z(n10679) );
  NAND2_X1 U13194 ( .A1(n10679), .A2(n10678), .ZN(n11060) );
  INV_X1 U13195 ( .A(n10679), .ZN(n10680) );
  NAND2_X1 U13196 ( .A1(n10680), .A2(n11058), .ZN(n10681) );
  NAND2_X1 U13197 ( .A1(n11060), .A2(n10681), .ZN(n10682) );
  AOI21_X1 U13198 ( .B1(n15314), .B2(n15318), .A(n10682), .ZN(n11062) );
  AND3_X1 U13199 ( .A1(n15314), .A2(n15318), .A3(n10682), .ZN(n10683) );
  OAI21_X1 U13200 ( .B1(n11062), .B2(n10683), .A(n15305), .ZN(n10684) );
  OAI211_X1 U13201 ( .C1(n10686), .C2(n15333), .A(n10685), .B(n10684), .ZN(
        P3_U3192) );
  INV_X1 U13202 ( .A(P3_DATAO_REG_27__SCAN_IN), .ZN(n13695) );
  NAND2_X1 U13203 ( .A1(n12422), .A2(P3_U3897), .ZN(n10687) );
  OAI21_X1 U13204 ( .B1(P3_U3897), .B2(n13695), .A(n10687), .ZN(P3_U3518) );
  NAND2_X1 U13205 ( .A1(n13009), .A2(n13272), .ZN(n10689) );
  AND2_X1 U13206 ( .A1(n10689), .A2(n10688), .ZN(n10690) );
  OR2_X1 U13207 ( .A1(n13013), .A2(n13271), .ZN(n10843) );
  NAND2_X1 U13208 ( .A1(n13013), .A2(n13271), .ZN(n10842) );
  NAND2_X1 U13209 ( .A1(n10843), .A2(n10842), .ZN(n13188) );
  XNOR2_X1 U13210 ( .A(n10845), .B(n13188), .ZN(n15133) );
  INV_X1 U13211 ( .A(n13013), .ZN(n15131) );
  OAI21_X1 U13212 ( .B1(n10692), .B2(n15131), .A(n15065), .ZN(n10693) );
  OR2_X1 U13213 ( .A1(n10693), .A2(n10852), .ZN(n15129) );
  INV_X1 U13214 ( .A(n10694), .ZN(n10695) );
  AOI22_X1 U13215 ( .A1(n15059), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n15058), 
        .B2(n10695), .ZN(n10697) );
  NAND2_X1 U13216 ( .A1(n15060), .A2(n13013), .ZN(n10696) );
  OAI211_X1 U13217 ( .C1(n15129), .C2(n13937), .A(n10697), .B(n10696), .ZN(
        n10702) );
  XNOR2_X1 U13218 ( .A(n10846), .B(n13188), .ZN(n10700) );
  AOI21_X1 U13219 ( .B1(n10700), .B2(n15054), .A(n10699), .ZN(n15130) );
  NOR2_X1 U13220 ( .A1(n15130), .A2(n15059), .ZN(n10701) );
  AOI211_X1 U13221 ( .C1(n15069), .C2(n15133), .A(n10702), .B(n10701), .ZN(
        n10703) );
  INV_X1 U13222 ( .A(n10703), .ZN(P2_U3258) );
  INV_X1 U13223 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10704) );
  AOI22_X1 U13224 ( .A1(n11029), .A2(n10704), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n10716), .ZN(n10710) );
  OR2_X1 U13225 ( .A1(n10706), .A2(n10705), .ZN(n10707) );
  OAI21_X1 U13226 ( .B1(n11395), .B2(n10708), .A(n10707), .ZN(n10709) );
  NOR2_X1 U13227 ( .A1(n10710), .A2(n10709), .ZN(n11032) );
  AOI21_X1 U13228 ( .B1(n10710), .B2(n10709), .A(n11032), .ZN(n10720) );
  INV_X1 U13229 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n14727) );
  AOI22_X1 U13230 ( .A1(n11029), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n14727), 
        .B2(n10716), .ZN(n10714) );
  OAI21_X1 U13231 ( .B1(n10714), .B2(n10713), .A(n11026), .ZN(n10718) );
  AOI22_X1 U13232 ( .A1(n14316), .A2(P1_ADDR_REG_12__SCAN_IN), .B1(
        P1_REG3_REG_12__SCAN_IN), .B2(P1_U3086), .ZN(n10715) );
  OAI21_X1 U13233 ( .B1(n10716), .B2(n14921), .A(n10715), .ZN(n10717) );
  AOI21_X1 U13234 ( .B1(n10718), .B2(n14913), .A(n10717), .ZN(n10719) );
  OAI21_X1 U13235 ( .B1(n10720), .B2(n14917), .A(n10719), .ZN(P1_U3255) );
  OAI21_X1 U13236 ( .B1(n10722), .B2(n10728), .A(n10721), .ZN(n10798) );
  INV_X1 U13237 ( .A(n10727), .ZN(n10725) );
  INV_X1 U13238 ( .A(n10862), .ZN(n10726) );
  AOI21_X1 U13239 ( .B1(n10728), .B2(n10727), .A(n10726), .ZN(n10731) );
  INV_X1 U13240 ( .A(n10729), .ZN(n10730) );
  OAI21_X1 U13241 ( .B1(n10731), .B2(n15359), .A(n10730), .ZN(n10799) );
  AOI21_X1 U13242 ( .B1(n14775), .B2(n10798), .A(n10799), .ZN(n11272) );
  INV_X1 U13243 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n10732) );
  OAI22_X1 U13244 ( .A1(n12651), .A2(n11269), .B1(n15436), .B2(n10732), .ZN(
        n10733) );
  INV_X1 U13245 ( .A(n10733), .ZN(n10734) );
  OAI21_X1 U13246 ( .B1(n11272), .B2(n15433), .A(n10734), .ZN(P3_U3464) );
  OAI22_X1 U13247 ( .A1(n10939), .A2(n12062), .B1(n10794), .B2(n12063), .ZN(
        n10739) );
  NAND2_X1 U13248 ( .A1(n6812), .A2(n10928), .ZN(n10742) );
  AOI22_X1 U13249 ( .A1(n12054), .A2(n14249), .B1(n12120), .B2(n10746), .ZN(
        n10741) );
  XNOR2_X1 U13250 ( .A(n10741), .B(n12121), .ZN(n10929) );
  XNOR2_X1 U13251 ( .A(n10742), .B(n10929), .ZN(n10749) );
  AND2_X1 U13252 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n14276) );
  OAI22_X1 U13253 ( .A1(n10743), .A2(n14900), .B1(n14899), .B2(n10961), .ZN(
        n10744) );
  AOI211_X1 U13254 ( .C1(n14228), .C2(n10745), .A(n14276), .B(n10744), .ZN(
        n10748) );
  NAND2_X1 U13255 ( .A1(n14215), .A2(n10746), .ZN(n10747) );
  OAI211_X1 U13256 ( .C1(n10749), .C2(n14850), .A(n10748), .B(n10747), .ZN(
        P1_U3230) );
  NAND2_X1 U13257 ( .A1(n10750), .A2(n10117), .ZN(n10753) );
  AOI22_X1 U13258 ( .A1(n12892), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n12733), 
        .B2(n10751), .ZN(n10752) );
  INV_X1 U13259 ( .A(n13022), .ZN(n15137) );
  INV_X1 U13260 ( .A(n10754), .ZN(n10756) );
  AND2_X1 U13261 ( .A1(n13270), .A2(n12855), .ZN(n10760) );
  XNOR2_X1 U13262 ( .A(n13022), .B(n12895), .ZN(n10759) );
  NOR2_X1 U13263 ( .A1(n10759), .A2(n10760), .ZN(n10915) );
  AOI21_X1 U13264 ( .B1(n10760), .B2(n10759), .A(n10915), .ZN(n10761) );
  OAI21_X1 U13265 ( .B1(n10762), .B2(n10761), .A(n10917), .ZN(n10763) );
  NAND2_X1 U13266 ( .A1(n10763), .A2(n14793), .ZN(n10776) );
  INV_X1 U13267 ( .A(n10851), .ZN(n10774) );
  INV_X1 U13268 ( .A(n13271), .ZN(n10847) );
  NAND2_X1 U13269 ( .A1(n12900), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n10771) );
  INV_X1 U13270 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10764) );
  OR2_X1 U13271 ( .A1(n12845), .A2(n10764), .ZN(n10770) );
  INV_X1 U13272 ( .A(n10884), .ZN(n10886) );
  NAND2_X1 U13273 ( .A1(n10766), .A2(n10765), .ZN(n10767) );
  NAND2_X1 U13274 ( .A1(n10886), .A2(n10767), .ZN(n10898) );
  OR2_X1 U13275 ( .A1(n12901), .A2(n10898), .ZN(n10769) );
  OR2_X1 U13276 ( .A1(n12903), .A2(n11128), .ZN(n10768) );
  NAND4_X1 U13277 ( .A1(n10771), .A2(n10770), .A3(n10769), .A4(n10768), .ZN(
        n13269) );
  INV_X1 U13278 ( .A(n13269), .ZN(n11172) );
  OAI22_X1 U13279 ( .A1(n10847), .A2(n12963), .B1(n12962), .B2(n11172), .ZN(
        n10772) );
  AOI211_X1 U13280 ( .C1(n10774), .C2(n11786), .A(n10773), .B(n10772), .ZN(
        n10775) );
  OAI211_X1 U13281 ( .C1(n15137), .C2(n11848), .A(n10776), .B(n10775), .ZN(
        P2_U3193) );
  OR2_X1 U13282 ( .A1(n10778), .A2(n10777), .ZN(n11011) );
  OAI21_X1 U13283 ( .B1(n10779), .B2(n10782), .A(n11011), .ZN(n10787) );
  OAI22_X1 U13284 ( .A1(n10961), .A2(n14438), .B1(n11657), .B2(n14466), .ZN(
        n10786) );
  NAND3_X1 U13285 ( .A1(n10780), .A2(n10782), .A3(n10781), .ZN(n10783) );
  AOI21_X1 U13286 ( .B1(n10784), .B2(n10783), .A(n14959), .ZN(n10785) );
  AOI211_X1 U13287 ( .C1(n14701), .C2(n10787), .A(n10786), .B(n10785), .ZN(
        n11040) );
  INV_X1 U13288 ( .A(n10788), .ZN(n10960) );
  OAI22_X1 U13289 ( .A1(n14531), .A2(n9843), .B1(n10960), .B2(n14498), .ZN(
        n10790) );
  OAI211_X1 U13290 ( .C1(n10806), .C2(n11041), .A(n14712), .B(n11006), .ZN(
        n11039) );
  NOR2_X1 U13291 ( .A1(n11039), .A2(n14529), .ZN(n10789) );
  AOI211_X1 U13292 ( .C1(n14706), .C2(n10964), .A(n10790), .B(n10789), .ZN(
        n10791) );
  OAI21_X1 U13293 ( .B1(n11040), .B2(n14705), .A(n10791), .ZN(P1_U3287) );
  OAI211_X1 U13294 ( .C1(n10794), .C2(n14947), .A(n10793), .B(n10792), .ZN(
        n10796) );
  NAND2_X1 U13295 ( .A1(n10796), .A2(n14982), .ZN(n10795) );
  OAI21_X1 U13296 ( .B1(n14982), .B2(n9832), .A(n10795), .ZN(P1_U3532) );
  NAND2_X1 U13297 ( .A1(n10796), .A2(n14973), .ZN(n10797) );
  OAI21_X1 U13298 ( .B1(n14973), .B2(n8444), .A(n10797), .ZN(P1_U3471) );
  INV_X1 U13299 ( .A(n10798), .ZN(n10805) );
  INV_X1 U13300 ( .A(n12581), .ZN(n12563) );
  INV_X1 U13301 ( .A(n10799), .ZN(n10800) );
  MUX2_X1 U13302 ( .A(n15257), .B(n10800), .S(n15380), .Z(n10804) );
  AOI22_X1 U13303 ( .A1(n12559), .A2(n10802), .B1(n15379), .B2(n10801), .ZN(
        n10803) );
  OAI211_X1 U13304 ( .C1(n10805), .C2(n12563), .A(n10804), .B(n10803), .ZN(
        P3_U3228) );
  INV_X1 U13305 ( .A(n10806), .ZN(n10807) );
  OAI211_X1 U13306 ( .C1(n14948), .C2(n10808), .A(n10807), .B(n14712), .ZN(
        n14945) );
  NAND2_X1 U13307 ( .A1(n10810), .A2(n10809), .ZN(n10811) );
  OAI21_X1 U13308 ( .B1(n10813), .B2(n10811), .A(n10780), .ZN(n10816) );
  OAI22_X1 U13309 ( .A1(n10953), .A2(n14466), .B1(n10939), .B2(n14438), .ZN(
        n10815) );
  AOI211_X1 U13310 ( .C1(n10813), .C2(n10812), .A(n14603), .B(n6807), .ZN(
        n10814) );
  AOI211_X1 U13311 ( .C1(n14965), .C2(n10816), .A(n10815), .B(n10814), .ZN(
        n14946) );
  MUX2_X1 U13312 ( .A(n10817), .B(n14946), .S(n14531), .Z(n10819) );
  AOI22_X1 U13313 ( .A1(n14706), .A2(n10934), .B1(n14703), .B2(n10942), .ZN(
        n10818) );
  OAI211_X1 U13314 ( .C1(n14529), .C2(n14945), .A(n10819), .B(n10818), .ZN(
        P1_U3288) );
  OAI21_X1 U13315 ( .B1(n10822), .B2(n10821), .A(n10820), .ZN(n10823) );
  AOI222_X1 U13316 ( .A1(n14701), .A2(n10823), .B1(n14249), .B2(n14540), .C1(
        n14251), .C2(n14539), .ZN(n14936) );
  AOI211_X1 U13317 ( .C1(n14939), .C2(n10825), .A(n14503), .B(n10824), .ZN(
        n14938) );
  NOR2_X1 U13318 ( .A1(n14506), .A2(n7099), .ZN(n10827) );
  OAI22_X1 U13319 ( .A1(n14531), .A2(n9436), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n14498), .ZN(n10826) );
  AOI211_X1 U13320 ( .C1(n14938), .C2(n14716), .A(n10827), .B(n10826), .ZN(
        n10832) );
  OAI21_X1 U13321 ( .B1(n10828), .B2(n10830), .A(n10829), .ZN(n14937) );
  INV_X1 U13322 ( .A(n14511), .ZN(n14717) );
  NAND2_X1 U13323 ( .A1(n14937), .A2(n14717), .ZN(n10831) );
  OAI211_X1 U13324 ( .C1(n14936), .C2(n14705), .A(n10832), .B(n10831), .ZN(
        P1_U3290) );
  INV_X1 U13325 ( .A(n10870), .ZN(n10840) );
  OAI211_X1 U13326 ( .C1(n10835), .C2(n10834), .A(n10833), .B(n15193), .ZN(
        n10839) );
  NAND2_X1 U13327 ( .A1(P3_REG3_REG_7__SCAN_IN), .A2(P3_U3151), .ZN(n15289) );
  INV_X1 U13328 ( .A(n15289), .ZN(n10837) );
  OAI22_X1 U13329 ( .A1(n10858), .A2(n12222), .B1(n12224), .B2(n11250), .ZN(
        n10836) );
  AOI211_X1 U13330 ( .C1(n11089), .C2(n15213), .A(n10837), .B(n10836), .ZN(
        n10838) );
  OAI211_X1 U13331 ( .C1(n10840), .C2(n15215), .A(n10839), .B(n10838), .ZN(
        P3_U3153) );
  INV_X1 U13332 ( .A(n12732), .ZN(n10904) );
  OAI222_X1 U13333 ( .A1(n11987), .A2(n10841), .B1(n6618), .B2(n10904), .C1(
        n13331), .C2(P2_U3088), .ZN(P2_U3308) );
  INV_X1 U13334 ( .A(n10842), .ZN(n10844) );
  XNOR2_X1 U13335 ( .A(n13022), .B(n10922), .ZN(n13192) );
  INV_X1 U13336 ( .A(n13192), .ZN(n10892) );
  XNOR2_X1 U13337 ( .A(n10893), .B(n10892), .ZN(n15135) );
  XNOR2_X1 U13338 ( .A(n10875), .B(n10892), .ZN(n10849) );
  OAI22_X1 U13339 ( .A1(n10847), .A2(n13928), .B1(n11172), .B2(n14784), .ZN(
        n10848) );
  AOI21_X1 U13340 ( .B1(n10849), .B2(n15054), .A(n10848), .ZN(n10850) );
  OAI21_X1 U13341 ( .B1(n10171), .B2(n15135), .A(n10850), .ZN(n15138) );
  NAND2_X1 U13342 ( .A1(n15138), .A2(n13944), .ZN(n10856) );
  OAI22_X1 U13343 ( .A1(n13944), .A2(n9612), .B1(n10851), .B2(n13957), .ZN(
        n10854) );
  OAI211_X1 U13344 ( .C1(n10852), .C2(n15137), .A(n15065), .B(n10897), .ZN(
        n15136) );
  NOR2_X1 U13345 ( .A1(n15136), .A2(n13937), .ZN(n10853) );
  AOI211_X1 U13346 ( .C1(n15060), .C2(n13022), .A(n10854), .B(n10853), .ZN(
        n10855) );
  OAI211_X1 U13347 ( .C1(n15135), .C2(n10900), .A(n10856), .B(n10855), .ZN(
        P2_U3257) );
  XNOR2_X1 U13348 ( .A(n10857), .B(n10865), .ZN(n10869) );
  OAI22_X1 U13349 ( .A1(n10858), .A2(n15353), .B1(n11250), .B2(n15351), .ZN(
        n10859) );
  INV_X1 U13350 ( .A(n10859), .ZN(n10868) );
  NAND2_X1 U13351 ( .A1(n10860), .A2(n11269), .ZN(n10861) );
  NAND2_X1 U13352 ( .A1(n12241), .A2(n15212), .ZN(n10864) );
  NAND2_X1 U13353 ( .A1(n10866), .A2(n10865), .ZN(n11091) );
  OAI211_X1 U13354 ( .C1(n10866), .C2(n10865), .A(n11091), .B(n15369), .ZN(
        n10867) );
  OAI211_X1 U13355 ( .C1(n10869), .C2(n15373), .A(n10868), .B(n10867), .ZN(
        n15400) );
  INV_X1 U13356 ( .A(n15400), .ZN(n10874) );
  INV_X2 U13357 ( .A(n15380), .ZN(n12443) );
  INV_X1 U13358 ( .A(n10869), .ZN(n15402) );
  INV_X1 U13359 ( .A(n15377), .ZN(n15342) );
  AND2_X1 U13360 ( .A1(n15380), .A2(n15342), .ZN(n12472) );
  AND2_X1 U13361 ( .A1(n14770), .A2(n11089), .ZN(n15401) );
  AOI22_X1 U13362 ( .A1(n15344), .A2(n15401), .B1(n15379), .B2(n10870), .ZN(
        n10871) );
  OAI21_X1 U13363 ( .B1(n15275), .B2(n15380), .A(n10871), .ZN(n10872) );
  AOI21_X1 U13364 ( .B1(n15402), .B2(n12472), .A(n10872), .ZN(n10873) );
  OAI21_X1 U13365 ( .B1(n10874), .B2(n12443), .A(n10873), .ZN(P3_U3226) );
  NAND2_X1 U13366 ( .A1(n10876), .A2(n10117), .ZN(n10882) );
  OAI22_X1 U13367 ( .A1(n10879), .A2(n10878), .B1(n9919), .B2(n10877), .ZN(
        n10880) );
  INV_X1 U13368 ( .A(n10880), .ZN(n10881) );
  XNOR2_X1 U13369 ( .A(n13027), .B(n11172), .ZN(n13194) );
  XNOR2_X1 U13370 ( .A(n11174), .B(n13194), .ZN(n10896) );
  NAND2_X1 U13371 ( .A1(n13168), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10891) );
  OR2_X1 U13372 ( .A1(n13172), .A2(n9693), .ZN(n10890) );
  INV_X1 U13373 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10883) );
  OR2_X1 U13374 ( .A1(n12845), .A2(n10883), .ZN(n10889) );
  INV_X1 U13375 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10885) );
  NAND2_X1 U13376 ( .A1(n10886), .A2(n10885), .ZN(n10887) );
  NAND2_X1 U13377 ( .A1(n10993), .A2(n10887), .ZN(n15056) );
  OR2_X1 U13378 ( .A1(n12901), .A2(n15056), .ZN(n10888) );
  NAND4_X1 U13379 ( .A1(n10891), .A2(n10890), .A3(n10889), .A4(n10888), .ZN(
        n13268) );
  INV_X1 U13380 ( .A(n13268), .ZN(n11178) );
  OAI22_X1 U13381 ( .A1(n10922), .A2(n13928), .B1(n11178), .B2(n14784), .ZN(
        n10895) );
  XNOR2_X1 U13382 ( .A(n11177), .B(n13194), .ZN(n11124) );
  NOR2_X1 U13383 ( .A1(n11124), .A2(n10171), .ZN(n10894) );
  AOI211_X1 U13384 ( .C1(n10896), .C2(n15054), .A(n10895), .B(n10894), .ZN(
        n11123) );
  INV_X1 U13385 ( .A(n11181), .ZN(n15066) );
  AOI211_X1 U13386 ( .C1(n13027), .C2(n10897), .A(n6611), .B(n15066), .ZN(
        n11121) );
  INV_X1 U13387 ( .A(n10898), .ZN(n10925) );
  AOI22_X1 U13388 ( .A1(n15059), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n15058), 
        .B2(n10925), .ZN(n10899) );
  OAI21_X1 U13389 ( .B1(n7074), .B2(n13959), .A(n10899), .ZN(n10902) );
  NOR2_X1 U13390 ( .A1(n11124), .A2(n10900), .ZN(n10901) );
  AOI211_X1 U13391 ( .C1(n11121), .C2(n15068), .A(n10902), .B(n10901), .ZN(
        n10903) );
  OAI21_X1 U13392 ( .B1(n11123), .B2(n15072), .A(n10903), .ZN(P2_U3256) );
  OAI222_X1 U13393 ( .A1(n12137), .A2(n10905), .B1(P1_U3086), .B2(n14334), 
        .C1(n14668), .C2(n10904), .ZN(P1_U3336) );
  NAND2_X1 U13394 ( .A1(n11260), .A2(n15374), .ZN(n10906) );
  OR2_X1 U13395 ( .A1(n10907), .A2(n10906), .ZN(n10909) );
  OR2_X1 U13396 ( .A1(n6846), .A2(n15351), .ZN(n10908) );
  NAND2_X1 U13397 ( .A1(n10909), .A2(n10908), .ZN(n11948) );
  MUX2_X1 U13398 ( .A(n11948), .B(P3_REG2_REG_0__SCAN_IN), .S(n12443), .Z(
        n10912) );
  INV_X1 U13399 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10910) );
  OAI22_X1 U13400 ( .A1(n12578), .A2(n11950), .B1(n12555), .B2(n10910), .ZN(
        n10911) );
  OR2_X1 U13401 ( .A1(n10912), .A2(n10911), .ZN(P3_U3233) );
  AND2_X1 U13402 ( .A1(n13269), .A2(n12855), .ZN(n10914) );
  XNOR2_X1 U13403 ( .A(n13027), .B(n12895), .ZN(n10913) );
  NOR2_X1 U13404 ( .A1(n10913), .A2(n10914), .ZN(n10984) );
  AOI21_X1 U13405 ( .B1(n10914), .B2(n10913), .A(n10984), .ZN(n10919) );
  INV_X1 U13406 ( .A(n10915), .ZN(n10916) );
  NAND2_X1 U13407 ( .A1(n10917), .A2(n10916), .ZN(n10918) );
  NAND2_X1 U13408 ( .A1(n10918), .A2(n10919), .ZN(n10986) );
  OAI21_X1 U13409 ( .B1(n10919), .B2(n10918), .A(n10986), .ZN(n10920) );
  NAND2_X1 U13410 ( .A1(n10920), .A2(n14793), .ZN(n10927) );
  INV_X1 U13411 ( .A(n10921), .ZN(n10924) );
  OAI22_X1 U13412 ( .A1(n10922), .A2(n12963), .B1(n12962), .B2(n11178), .ZN(
        n10923) );
  AOI211_X1 U13413 ( .C1(n10925), .C2(n11786), .A(n10924), .B(n10923), .ZN(
        n10926) );
  OAI211_X1 U13414 ( .C1(n7074), .C2(n11848), .A(n10927), .B(n10926), .ZN(
        P2_U3203) );
  NAND2_X1 U13415 ( .A1(n10934), .A2(n12120), .ZN(n10931) );
  NAND2_X1 U13416 ( .A1(n14248), .A2(n12054), .ZN(n10930) );
  NAND2_X1 U13417 ( .A1(n10931), .A2(n10930), .ZN(n10933) );
  XNOR2_X1 U13418 ( .A(n10933), .B(n10252), .ZN(n10945) );
  NAND2_X1 U13419 ( .A1(n12119), .A2(n14248), .ZN(n10936) );
  NAND2_X1 U13420 ( .A1(n10934), .A2(n12073), .ZN(n10935) );
  XNOR2_X1 U13421 ( .A(n10945), .B(n10946), .ZN(n10937) );
  XNOR2_X1 U13422 ( .A(n10949), .B(n10937), .ZN(n10938) );
  NAND2_X1 U13423 ( .A1(n10938), .A2(n14904), .ZN(n10944) );
  OAI22_X1 U13424 ( .A1(n10939), .A2(n14900), .B1(n14899), .B2(n10953), .ZN(
        n10940) );
  AOI211_X1 U13425 ( .C1(n14228), .C2(n10942), .A(n10941), .B(n10940), .ZN(
        n10943) );
  OAI211_X1 U13426 ( .C1(n14948), .C2(n14896), .A(n10944), .B(n10943), .ZN(
        P1_U3227) );
  INV_X1 U13427 ( .A(n10945), .ZN(n10948) );
  INV_X1 U13428 ( .A(n10946), .ZN(n10947) );
  NAND2_X1 U13429 ( .A1(n10964), .A2(n12120), .ZN(n10951) );
  NAND2_X1 U13430 ( .A1(n14247), .A2(n12112), .ZN(n10950) );
  NAND2_X1 U13431 ( .A1(n10951), .A2(n10950), .ZN(n10952) );
  XNOR2_X1 U13432 ( .A(n10952), .B(n10252), .ZN(n10955) );
  NOR2_X1 U13433 ( .A1(n10953), .A2(n12062), .ZN(n10954) );
  AOI21_X1 U13434 ( .B1(n10964), .B2(n12054), .A(n10954), .ZN(n10956) );
  INV_X1 U13435 ( .A(n10955), .ZN(n10958) );
  INV_X1 U13436 ( .A(n10956), .ZN(n10957) );
  NAND2_X1 U13437 ( .A1(n10958), .A2(n10957), .ZN(n11662) );
  NAND2_X1 U13438 ( .A1(n6816), .A2(n11662), .ZN(n10959) );
  XNOR2_X1 U13439 ( .A(n11663), .B(n10959), .ZN(n10966) );
  OAI22_X1 U13440 ( .A1(n14909), .A2(n10960), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13662), .ZN(n10963) );
  OAI22_X1 U13441 ( .A1(n10961), .A2(n14900), .B1(n14899), .B2(n11657), .ZN(
        n10962) );
  AOI211_X1 U13442 ( .C1(n14215), .C2(n10964), .A(n10963), .B(n10962), .ZN(
        n10965) );
  OAI21_X1 U13443 ( .B1(n10966), .B2(n14850), .A(n10965), .ZN(P1_U3239) );
  NAND2_X1 U13444 ( .A1(n10967), .A2(n12719), .ZN(n10969) );
  OAI211_X1 U13445 ( .C1(n10970), .C2(n12725), .A(n10969), .B(n10968), .ZN(
        P3_U3272) );
  OAI21_X1 U13446 ( .B1(n10973), .B2(n10972), .A(n10971), .ZN(n10974) );
  INV_X1 U13447 ( .A(n10974), .ZN(n14960) );
  OAI211_X1 U13448 ( .C1(n10977), .C2(n10976), .A(n10975), .B(n14701), .ZN(
        n10979) );
  AOI22_X1 U13449 ( .A1(n14244), .A2(n14540), .B1(n14539), .B2(n14246), .ZN(
        n10978) );
  AND2_X1 U13450 ( .A1(n10979), .A2(n10978), .ZN(n14958) );
  MUX2_X1 U13451 ( .A(n14958), .B(n10980), .S(n14526), .Z(n10983) );
  AOI211_X1 U13452 ( .C1(n14956), .C2(n11007), .A(n14503), .B(n6804), .ZN(
        n14955) );
  OAI22_X1 U13453 ( .A1(n7105), .A2(n14506), .B1(n11960), .B2(n14498), .ZN(
        n10981) );
  AOI21_X1 U13454 ( .B1(n14955), .B2(n14716), .A(n10981), .ZN(n10982) );
  OAI211_X1 U13455 ( .C1(n14960), .C2(n14511), .A(n10983), .B(n10982), .ZN(
        P1_U3285) );
  INV_X1 U13456 ( .A(n10984), .ZN(n10985) );
  NAND2_X1 U13457 ( .A1(n13268), .A2(n12855), .ZN(n11147) );
  NAND2_X1 U13458 ( .A1(n10987), .A2(n10117), .ZN(n10990) );
  AOI22_X1 U13459 ( .A1(n10988), .A2(n12733), .B1(n12892), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n10989) );
  XNOR2_X1 U13460 ( .A(n15061), .B(n12895), .ZN(n11146) );
  XOR2_X1 U13461 ( .A(n11147), .B(n11146), .Z(n11149) );
  XNOR2_X1 U13462 ( .A(n11150), .B(n11149), .ZN(n11005) );
  NAND2_X1 U13463 ( .A1(n14787), .A2(n13269), .ZN(n11000) );
  NAND2_X1 U13464 ( .A1(n12900), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n10998) );
  INV_X1 U13465 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10991) );
  OR2_X1 U13466 ( .A1(n12845), .A2(n10991), .ZN(n10997) );
  INV_X1 U13467 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10992) );
  NAND2_X1 U13468 ( .A1(n10993), .A2(n10992), .ZN(n10994) );
  NAND2_X1 U13469 ( .A1(n11161), .A2(n10994), .ZN(n11183) );
  OR2_X1 U13470 ( .A1(n12901), .A2(n11183), .ZN(n10996) );
  OR2_X1 U13471 ( .A1(n12775), .A2(n15175), .ZN(n10995) );
  NAND4_X1 U13472 ( .A1(n10998), .A2(n10997), .A3(n10996), .A4(n10995), .ZN(
        n13267) );
  NAND2_X1 U13473 ( .A1(n13949), .A2(n13267), .ZN(n10999) );
  NAND2_X1 U13474 ( .A1(n11000), .A2(n10999), .ZN(n15053) );
  NAND2_X1 U13475 ( .A1(n14795), .A2(n15053), .ZN(n11002) );
  OAI211_X1 U13476 ( .C1(n14799), .C2(n15056), .A(n11002), .B(n11001), .ZN(
        n11003) );
  AOI21_X1 U13477 ( .B1(n15061), .B2(n14796), .A(n11003), .ZN(n11004) );
  OAI21_X1 U13478 ( .B1(n11005), .B2(n12967), .A(n11004), .ZN(P2_U3189) );
  AOI21_X1 U13479 ( .B1(n11006), .B2(n14954), .A(n14503), .ZN(n11008) );
  NAND2_X1 U13480 ( .A1(n11008), .A2(n11007), .ZN(n14951) );
  AND2_X1 U13481 ( .A1(n11011), .A2(n11009), .ZN(n11014) );
  NAND2_X1 U13482 ( .A1(n11011), .A2(n11010), .ZN(n11012) );
  OAI211_X1 U13483 ( .C1(n11014), .C2(n11013), .A(n11012), .B(n14701), .ZN(
        n11021) );
  AOI22_X1 U13484 ( .A1(n14539), .A2(n14247), .B1(n14245), .B2(n14540), .ZN(
        n11020) );
  OAI21_X1 U13485 ( .B1(n11017), .B2(n11016), .A(n11015), .ZN(n11018) );
  NAND2_X1 U13486 ( .A1(n11018), .A2(n14965), .ZN(n11019) );
  NAND3_X1 U13487 ( .A1(n11021), .A2(n11020), .A3(n11019), .ZN(n14952) );
  MUX2_X1 U13488 ( .A(n14952), .B(P1_REG2_REG_7__SCAN_IN), .S(n14526), .Z(
        n11022) );
  INV_X1 U13489 ( .A(n11022), .ZN(n11024) );
  AOI22_X1 U13490 ( .A1(n14706), .A2(n14954), .B1(n14078), .B2(n14703), .ZN(
        n11023) );
  OAI211_X1 U13491 ( .C1(n14529), .C2(n14951), .A(n11024), .B(n11023), .ZN(
        P1_U3286) );
  INV_X1 U13492 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11025) );
  MUX2_X1 U13493 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n11025), .S(n11205), .Z(
        n11028) );
  OAI21_X1 U13494 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n11029), .A(n11026), 
        .ZN(n11027) );
  NOR2_X1 U13495 ( .A1(n11027), .A2(n11028), .ZN(n11207) );
  AOI211_X1 U13496 ( .C1(n11028), .C2(n11027), .A(n14298), .B(n11207), .ZN(
        n11038) );
  NOR2_X1 U13497 ( .A1(n11029), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n11031) );
  INV_X1 U13498 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11206) );
  MUX2_X1 U13499 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n11206), .S(n11205), .Z(
        n11030) );
  OAI21_X1 U13500 ( .B1(n11032), .B2(n11031), .A(n11030), .ZN(n11033) );
  NAND3_X1 U13501 ( .A1(n11204), .A2(n14332), .A3(n11033), .ZN(n11036) );
  NAND2_X1 U13502 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n11932)
         );
  INV_X1 U13503 ( .A(n11932), .ZN(n11034) );
  AOI21_X1 U13504 ( .B1(n14316), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n11034), 
        .ZN(n11035) );
  OAI211_X1 U13505 ( .C1(n14921), .C2(n11205), .A(n11036), .B(n11035), .ZN(
        n11037) );
  OR2_X1 U13506 ( .A1(n11038), .A2(n11037), .ZN(P1_U3256) );
  INV_X1 U13507 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n11043) );
  OAI211_X1 U13508 ( .C1(n11041), .C2(n14947), .A(n11040), .B(n11039), .ZN(
        n11044) );
  NAND2_X1 U13509 ( .A1(n11044), .A2(n14973), .ZN(n11042) );
  OAI21_X1 U13510 ( .B1(n14973), .B2(n11043), .A(n11042), .ZN(P1_U3477) );
  NAND2_X1 U13511 ( .A1(n11044), .A2(n14982), .ZN(n11045) );
  OAI21_X1 U13512 ( .B1(n14982), .B2(n7096), .A(n11045), .ZN(P1_U3534) );
  INV_X1 U13513 ( .A(n11101), .ZN(n11052) );
  NAND2_X1 U13514 ( .A1(n15181), .A2(n11047), .ZN(n11282) );
  OAI211_X1 U13515 ( .C1(n15181), .C2(n11047), .A(n11282), .B(n15193), .ZN(
        n11051) );
  NAND2_X1 U13516 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_U3151), .ZN(n15306) );
  INV_X1 U13517 ( .A(n15306), .ZN(n11049) );
  OAI22_X1 U13518 ( .A1(n11094), .A2(n12222), .B1(n12224), .B2(n11095), .ZN(
        n11048) );
  AOI211_X1 U13519 ( .C1(n15213), .C2(n11100), .A(n11049), .B(n11048), .ZN(
        n11050) );
  OAI211_X1 U13520 ( .C1(n15215), .C2(n11052), .A(n11051), .B(n11050), .ZN(
        P3_U3161) );
  INV_X1 U13521 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11055) );
  AOI21_X1 U13522 ( .B1(n11056), .B2(n11055), .A(n11222), .ZN(n11074) );
  XNOR2_X1 U13523 ( .A(n11226), .B(n11065), .ZN(n11059) );
  OAI21_X1 U13524 ( .B1(n11059), .B2(P3_REG1_REG_11__SCAN_IN), .A(n11227), 
        .ZN(n11072) );
  INV_X1 U13525 ( .A(n11060), .ZN(n11061) );
  MUX2_X1 U13526 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n14735), .Z(n11231) );
  XNOR2_X1 U13527 ( .A(n11231), .B(n11065), .ZN(n11063) );
  NOR2_X1 U13528 ( .A1(n11064), .A2(n11063), .ZN(n11232) );
  AOI21_X1 U13529 ( .B1(n11064), .B2(n11063), .A(n11232), .ZN(n11070) );
  INV_X1 U13530 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11066) );
  NOR2_X1 U13531 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11066), .ZN(n11068) );
  NOR2_X1 U13532 ( .A1(n15308), .A2(n13539), .ZN(n11067) );
  AOI211_X1 U13533 ( .C1(n15266), .C2(n7247), .A(n11068), .B(n11067), .ZN(
        n11069) );
  OAI21_X1 U13534 ( .B1(n11070), .B2(n15322), .A(n11069), .ZN(n11071) );
  AOI21_X1 U13535 ( .B1(n11072), .B2(n15329), .A(n11071), .ZN(n11073) );
  OAI21_X1 U13536 ( .B1(n11074), .B2(n15333), .A(n11073), .ZN(P3_U3193) );
  XNOR2_X1 U13537 ( .A(n11075), .B(n11077), .ZN(n15398) );
  INV_X1 U13538 ( .A(n15344), .ZN(n11076) );
  NAND2_X1 U13539 ( .A1(n14770), .A2(n15212), .ZN(n15395) );
  OAI22_X1 U13540 ( .A1(n11076), .A2(n15395), .B1(n15216), .B2(n12555), .ZN(
        n11086) );
  AOI21_X1 U13541 ( .B1(n11078), .B2(n11077), .A(n15359), .ZN(n11080) );
  NAND2_X1 U13542 ( .A1(n11080), .A2(n11079), .ZN(n11084) );
  INV_X1 U13543 ( .A(n15373), .ZN(n15356) );
  NAND2_X1 U13544 ( .A1(n15398), .A2(n15356), .ZN(n11083) );
  OR2_X1 U13545 ( .A1(n11094), .A2(n15351), .ZN(n11082) );
  NAND2_X1 U13546 ( .A1(n12406), .A2(n12242), .ZN(n11081) );
  AND2_X1 U13547 ( .A1(n11082), .A2(n11081), .ZN(n15204) );
  NAND3_X1 U13548 ( .A1(n11084), .A2(n11083), .A3(n15204), .ZN(n15396) );
  MUX2_X1 U13549 ( .A(n15396), .B(P3_REG2_REG_6__SCAN_IN), .S(n12443), .Z(
        n11085) );
  AOI211_X1 U13550 ( .C1(n15398), .C2(n12472), .A(n11086), .B(n11085), .ZN(
        n11087) );
  INV_X1 U13551 ( .A(n11087), .ZN(P3_U3227) );
  XNOR2_X1 U13552 ( .A(n11088), .B(n11092), .ZN(n11099) );
  NAND2_X1 U13553 ( .A1(n12240), .A2(n11089), .ZN(n11090) );
  AND2_X2 U13554 ( .A1(n11091), .A2(n11090), .ZN(n11093) );
  OAI21_X1 U13555 ( .B1(n11093), .B2(n11092), .A(n11247), .ZN(n11097) );
  OAI22_X1 U13556 ( .A1(n11095), .A2(n15351), .B1(n11094), .B2(n15353), .ZN(
        n11096) );
  AOI21_X1 U13557 ( .B1(n11097), .B2(n15369), .A(n11096), .ZN(n11098) );
  OAI21_X1 U13558 ( .B1(n15373), .B2(n11099), .A(n11098), .ZN(n15404) );
  INV_X1 U13559 ( .A(n15404), .ZN(n11106) );
  INV_X1 U13560 ( .A(n11099), .ZN(n15406) );
  INV_X1 U13561 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11103) );
  AND2_X1 U13562 ( .A1(n14770), .A2(n11100), .ZN(n15405) );
  AOI22_X1 U13563 ( .A1(n15344), .A2(n15405), .B1(n11101), .B2(n15379), .ZN(
        n11102) );
  OAI21_X1 U13564 ( .B1(n11103), .B2(n15380), .A(n11102), .ZN(n11104) );
  AOI21_X1 U13565 ( .B1(n15406), .B2(n12472), .A(n11104), .ZN(n11105) );
  OAI21_X1 U13566 ( .B1(n11106), .B2(n12443), .A(n11105), .ZN(P3_U3225) );
  OAI21_X1 U13567 ( .B1(n11109), .B2(n11108), .A(n11107), .ZN(n11115) );
  OAI22_X1 U13568 ( .A1(n14901), .A2(n14438), .B1(n14898), .B2(n14466), .ZN(
        n11114) );
  NAND2_X1 U13569 ( .A1(n11110), .A2(n11109), .ZN(n11111) );
  AOI21_X1 U13570 ( .B1(n11112), .B2(n11111), .A(n14603), .ZN(n11113) );
  AOI211_X1 U13571 ( .C1(n14965), .C2(n11115), .A(n11114), .B(n11113), .ZN(
        n11295) );
  OAI211_X1 U13572 ( .C1(n6804), .C2(n14897), .A(n11195), .B(n14712), .ZN(
        n11294) );
  AOI22_X1 U13573 ( .A1(n14705), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n11116), 
        .B2(n14703), .ZN(n11118) );
  NAND2_X1 U13574 ( .A1(n11671), .A2(n14706), .ZN(n11117) );
  OAI211_X1 U13575 ( .C1(n11294), .C2(n14529), .A(n11118), .B(n11117), .ZN(
        n11119) );
  INV_X1 U13576 ( .A(n11119), .ZN(n11120) );
  OAI21_X1 U13577 ( .B1(n11295), .B2(n14705), .A(n11120), .ZN(P1_U3284) );
  INV_X1 U13578 ( .A(n12969), .ZN(n13971) );
  AOI21_X1 U13579 ( .B1(n15114), .B2(n13027), .A(n11121), .ZN(n11122) );
  OAI211_X1 U13580 ( .C1(n11124), .C2(n13971), .A(n11123), .B(n11122), .ZN(
        n11126) );
  NAND2_X1 U13581 ( .A1(n11126), .A2(n15157), .ZN(n11125) );
  OAI21_X1 U13582 ( .B1(n15157), .B2(n10764), .A(n11125), .ZN(P2_U3457) );
  NAND2_X1 U13583 ( .A1(n11126), .A2(n15177), .ZN(n11127) );
  OAI21_X1 U13584 ( .B1(n15177), .B2(n11128), .A(n11127), .ZN(P2_U3508) );
  INV_X1 U13585 ( .A(n11129), .ZN(n11132) );
  NAND2_X1 U13586 ( .A1(n14125), .A2(n11130), .ZN(n11131) );
  NAND2_X1 U13587 ( .A1(n11132), .A2(n11131), .ZN(n11139) );
  XNOR2_X1 U13588 ( .A(n11139), .B(n8910), .ZN(n11133) );
  MUX2_X1 U13589 ( .A(n11133), .B(n9097), .S(n6609), .Z(n11134) );
  OAI222_X1 U13590 ( .A1(n14438), .A2(n6607), .B1(n14466), .B2(n11135), .C1(
        n14603), .C2(n11134), .ZN(n14932) );
  OAI21_X1 U13591 ( .B1(n11138), .B2(n11137), .A(n11136), .ZN(n14934) );
  INV_X1 U13592 ( .A(n11139), .ZN(n11140) );
  NAND2_X1 U13593 ( .A1(n11140), .A2(n14712), .ZN(n14931) );
  INV_X1 U13594 ( .A(n14931), .ZN(n11141) );
  AOI22_X1 U13595 ( .A1(n14717), .A2(n14934), .B1(n14716), .B2(n11141), .ZN(
        n11143) );
  AOI22_X1 U13596 ( .A1(n14705), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n14703), .ZN(n11142) );
  OAI211_X1 U13597 ( .C1(n6821), .C2(n14506), .A(n11143), .B(n11142), .ZN(
        n11144) );
  AOI21_X1 U13598 ( .B1(n14531), .B2(n14932), .A(n11144), .ZN(n11145) );
  INV_X1 U13599 ( .A(n11145), .ZN(P1_U3292) );
  INV_X1 U13600 ( .A(n11146), .ZN(n11148) );
  NAND2_X1 U13601 ( .A1(n11151), .A2(n10117), .ZN(n11154) );
  AOI22_X1 U13602 ( .A1(n11152), .A2(n12733), .B1(n12892), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n11153) );
  XNOR2_X1 U13603 ( .A(n13040), .B(n11155), .ZN(n11157) );
  NAND2_X1 U13604 ( .A1(n13267), .A2(n12855), .ZN(n11156) );
  NAND2_X1 U13605 ( .A1(n11157), .A2(n11156), .ZN(n11299) );
  OAI21_X1 U13606 ( .B1(n11157), .B2(n11156), .A(n11299), .ZN(n11158) );
  AOI21_X1 U13607 ( .B1(n11159), .B2(n11158), .A(n11301), .ZN(n11171) );
  NOR2_X1 U13608 ( .A1(n14799), .A2(n11183), .ZN(n11169) );
  INV_X1 U13609 ( .A(n14795), .ZN(n12951) );
  NAND2_X1 U13610 ( .A1(n13169), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n11166) );
  OR2_X1 U13611 ( .A1(n13172), .A2(n10304), .ZN(n11165) );
  INV_X1 U13612 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n11160) );
  INV_X1 U13613 ( .A(n11309), .ZN(n11311) );
  NAND2_X1 U13614 ( .A1(n11161), .A2(n11160), .ZN(n11162) );
  NAND2_X1 U13615 ( .A1(n11311), .A2(n11162), .ZN(n11416) );
  OR2_X1 U13616 ( .A1(n12901), .A2(n11416), .ZN(n11164) );
  OR2_X1 U13617 ( .A1(n12903), .A2(n14836), .ZN(n11163) );
  NAND4_X1 U13618 ( .A1(n11166), .A2(n11165), .A3(n11164), .A4(n11163), .ZN(
        n13266) );
  AOI22_X1 U13619 ( .A1(n14787), .A2(n13268), .B1(n13949), .B2(n13266), .ZN(
        n11175) );
  OAI21_X1 U13620 ( .B1(n12951), .B2(n11175), .A(n11167), .ZN(n11168) );
  AOI211_X1 U13621 ( .C1(n13040), .C2(n14796), .A(n11169), .B(n11168), .ZN(
        n11170) );
  OAI21_X1 U13622 ( .B1(n11171), .B2(n12967), .A(n11170), .ZN(P2_U3208) );
  NOR2_X1 U13623 ( .A1(n13027), .A2(n11172), .ZN(n11173) );
  XNOR2_X1 U13624 ( .A(n15061), .B(n13268), .ZN(n15062) );
  XNOR2_X1 U13625 ( .A(n13040), .B(n13267), .ZN(n13199) );
  XNOR2_X1 U13626 ( .A(n11357), .B(n13199), .ZN(n11176) );
  OAI21_X1 U13627 ( .B1(n11176), .B2(n13925), .A(n11175), .ZN(n15152) );
  INV_X1 U13628 ( .A(n15152), .ZN(n11189) );
  INV_X1 U13629 ( .A(n15061), .ZN(n15142) );
  XNOR2_X1 U13630 ( .A(n11379), .B(n11378), .ZN(n15154) );
  NAND2_X1 U13631 ( .A1(n13040), .A2(n15064), .ZN(n11182) );
  NAND3_X1 U13632 ( .A1(n11412), .A2(n15065), .A3(n11182), .ZN(n15148) );
  INV_X1 U13633 ( .A(n11183), .ZN(n11184) );
  AOI22_X1 U13634 ( .A1(n15072), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n15058), 
        .B2(n11184), .ZN(n11186) );
  NAND2_X1 U13635 ( .A1(n13040), .A2(n15060), .ZN(n11185) );
  OAI211_X1 U13636 ( .C1(n15148), .C2(n13937), .A(n11186), .B(n11185), .ZN(
        n11187) );
  AOI21_X1 U13637 ( .B1(n15154), .B2(n15069), .A(n11187), .ZN(n11188) );
  OAI21_X1 U13638 ( .B1(n11189), .B2(n15072), .A(n11188), .ZN(P2_U3254) );
  AOI21_X1 U13639 ( .B1(n6810), .B2(n11193), .A(n14603), .ZN(n11191) );
  AOI22_X1 U13640 ( .A1(n11191), .A2(n11190), .B1(n14539), .B2(n14244), .ZN(
        n14968) );
  OAI21_X1 U13641 ( .B1(n11194), .B2(n11193), .A(n11192), .ZN(n14966) );
  INV_X1 U13642 ( .A(n11195), .ZN(n11197) );
  OAI211_X1 U13643 ( .C1(n11687), .C2(n11197), .A(n14712), .B(n11396), .ZN(
        n11198) );
  OAI21_X1 U13644 ( .B1(n11680), .B2(n14466), .A(n11198), .ZN(n14970) );
  NAND2_X1 U13645 ( .A1(n14970), .A2(n14716), .ZN(n11200) );
  AOI22_X1 U13646 ( .A1(n14705), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n11684), 
        .B2(n14703), .ZN(n11199) );
  OAI211_X1 U13647 ( .C1(n11687), .C2(n14506), .A(n11200), .B(n11199), .ZN(
        n11201) );
  AOI21_X1 U13648 ( .B1(n14966), .B2(n14717), .A(n11201), .ZN(n11202) );
  OAI21_X1 U13649 ( .B1(n14968), .B2(n14705), .A(n11202), .ZN(P1_U3283) );
  INV_X1 U13650 ( .A(n12741), .ZN(n11292) );
  OAI222_X1 U13651 ( .A1(n11987), .A2(n11203), .B1(n6618), .B2(n11292), .C1(
        n9906), .C2(P2_U3088), .ZN(P2_U3307) );
  OAI21_X1 U13652 ( .B1(n11206), .B2(n11205), .A(n11204), .ZN(n11638) );
  MUX2_X1 U13653 ( .A(n8586), .B(P1_REG2_REG_14__SCAN_IN), .S(n11644), .Z(
        n11636) );
  XOR2_X1 U13654 ( .A(n11638), .B(n11636), .Z(n11217) );
  XOR2_X1 U13655 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n11644), .Z(n11210) );
  OAI21_X1 U13656 ( .B1(n11210), .B2(n11209), .A(n11643), .ZN(n11215) );
  NOR2_X1 U13657 ( .A1(n11211), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14097) );
  AOI21_X1 U13658 ( .B1(n14316), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n14097), 
        .ZN(n11212) );
  OAI21_X1 U13659 ( .B1(n11213), .B2(n14921), .A(n11212), .ZN(n11214) );
  AOI21_X1 U13660 ( .B1(n11215), .B2(n14913), .A(n11214), .ZN(n11216) );
  OAI21_X1 U13661 ( .B1(n14917), .B2(n11217), .A(n11216), .ZN(P1_U3257) );
  INV_X1 U13662 ( .A(n11219), .ZN(n11221) );
  OAI222_X1 U13663 ( .A1(n9147), .A2(P3_U3151), .B1(n11991), .B2(n11221), .C1(
        n11220), .C2(n11995), .ZN(P3_U3271) );
  INV_X1 U13664 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n13677) );
  AOI22_X1 U13665 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n11476), .B1(n11239), 
        .B2(n13677), .ZN(n11224) );
  AOI21_X1 U13666 ( .B1(n11225), .B2(n11224), .A(n11467), .ZN(n11243) );
  INV_X1 U13667 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n13689) );
  AOI22_X1 U13668 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n11239), .B1(n11476), 
        .B2(n13689), .ZN(n11230) );
  OR2_X1 U13669 ( .A1(n11226), .A2(n7247), .ZN(n11228) );
  OAI21_X1 U13670 ( .B1(n11230), .B2(n11229), .A(n11471), .ZN(n11241) );
  INV_X1 U13671 ( .A(n11231), .ZN(n11233) );
  AOI21_X1 U13672 ( .B1(n7247), .B2(n11233), .A(n11232), .ZN(n11235) );
  MUX2_X1 U13673 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n14735), .Z(n11473) );
  XNOR2_X1 U13674 ( .A(n11473), .B(n11476), .ZN(n11234) );
  NAND2_X1 U13675 ( .A1(n11235), .A2(n11234), .ZN(n11474) );
  OAI211_X1 U13676 ( .C1(n11235), .C2(n11234), .A(n11474), .B(n15305), .ZN(
        n11238) );
  AND2_X1 U13677 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n11236) );
  AOI21_X1 U13678 ( .B1(n15326), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n11236), 
        .ZN(n11237) );
  OAI211_X1 U13679 ( .C1(n15320), .C2(n11239), .A(n11238), .B(n11237), .ZN(
        n11240) );
  AOI21_X1 U13680 ( .B1(n15329), .B2(n11241), .A(n11240), .ZN(n11242) );
  OAI21_X1 U13681 ( .B1(n11243), .B2(n15333), .A(n11242), .ZN(P3_U3194) );
  XNOR2_X1 U13682 ( .A(n11244), .B(n11248), .ZN(n11254) );
  NAND2_X1 U13683 ( .A1(n11250), .A2(n11245), .ZN(n11246) );
  AND2_X2 U13684 ( .A1(n11247), .A2(n11246), .ZN(n11249) );
  OAI211_X1 U13685 ( .C1(n11249), .C2(n11248), .A(n11327), .B(n15369), .ZN(
        n11253) );
  OAI22_X1 U13686 ( .A1(n11442), .A2(n15351), .B1(n11250), .B2(n15353), .ZN(
        n11251) );
  INV_X1 U13687 ( .A(n11251), .ZN(n11252) );
  OAI211_X1 U13688 ( .C1(n15373), .C2(n11254), .A(n11253), .B(n11252), .ZN(
        n15408) );
  INV_X1 U13689 ( .A(n15408), .ZN(n11258) );
  INV_X1 U13690 ( .A(n11254), .ZN(n15411) );
  NOR2_X1 U13691 ( .A1(n11287), .A2(n15374), .ZN(n15409) );
  AOI22_X1 U13692 ( .A1(n15344), .A2(n15409), .B1(n15379), .B2(n11289), .ZN(
        n11255) );
  OAI21_X1 U13693 ( .B1(n15312), .B2(n15380), .A(n11255), .ZN(n11256) );
  AOI21_X1 U13694 ( .B1(n15411), .B2(n12472), .A(n11256), .ZN(n11257) );
  OAI21_X1 U13695 ( .B1(n11258), .B2(n12443), .A(n11257), .ZN(P3_U3224) );
  NAND2_X1 U13696 ( .A1(n11260), .A2(n11259), .ZN(n11262) );
  NAND2_X1 U13697 ( .A1(n11262), .A2(n11261), .ZN(n11267) );
  NAND2_X1 U13698 ( .A1(n11264), .A2(n11263), .ZN(n11266) );
  INV_X1 U13699 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n11268) );
  OAI22_X1 U13700 ( .A1(n12712), .A2(n11269), .B1(n12707), .B2(n11268), .ZN(
        n11270) );
  INV_X1 U13701 ( .A(n11270), .ZN(n11271) );
  OAI21_X1 U13702 ( .B1(n11272), .B2(n15419), .A(n11271), .ZN(P3_U3405) );
  INV_X1 U13703 ( .A(n11273), .ZN(n11276) );
  INV_X1 U13704 ( .A(n12712), .ZN(n12684) );
  AOI22_X1 U13705 ( .A1(n12684), .A2(n11274), .B1(n15419), .B2(
        P3_REG0_REG_4__SCAN_IN), .ZN(n11275) );
  OAI21_X1 U13706 ( .B1(n11276), .B2(n15419), .A(n11275), .ZN(P3_U3402) );
  INV_X1 U13707 ( .A(n12760), .ZN(n11279) );
  OAI222_X1 U13708 ( .A1(n12137), .A2(n11278), .B1(n14668), .B2(n11279), .C1(
        n11277), .C2(P1_U3086), .ZN(P1_U3334) );
  INV_X1 U13709 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11280) );
  OAI222_X1 U13710 ( .A1(n11987), .A2(n11280), .B1(n6618), .B2(n11279), .C1(
        P2_U3088), .C2(n13215), .ZN(P2_U3306) );
  NAND2_X1 U13711 ( .A1(n11282), .A2(n11281), .ZN(n11283) );
  AOI21_X1 U13712 ( .B1(n11284), .B2(n11283), .A(n6806), .ZN(n11291) );
  OAI22_X1 U13713 ( .A1(n12224), .A2(n11442), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15313), .ZN(n11285) );
  AOI21_X1 U13714 ( .B1(n12212), .B2(n12239), .A(n11285), .ZN(n11286) );
  OAI21_X1 U13715 ( .B1(n11287), .B2(n12230), .A(n11286), .ZN(n11288) );
  AOI21_X1 U13716 ( .B1(n11289), .B2(n12227), .A(n11288), .ZN(n11290) );
  OAI21_X1 U13717 ( .B1(n11291), .B2(n15207), .A(n11290), .ZN(P3_U3171) );
  OAI222_X1 U13718 ( .A1(n12137), .A2(n11293), .B1(P1_U3086), .B2(n8900), .C1(
        n14668), .C2(n11292), .ZN(P1_U3335) );
  OAI211_X1 U13719 ( .C1(n14897), .C2(n14947), .A(n11295), .B(n11294), .ZN(
        n11297) );
  NAND2_X1 U13720 ( .A1(n11297), .A2(n14982), .ZN(n11296) );
  OAI21_X1 U13721 ( .B1(n14982), .B2(n9953), .A(n11296), .ZN(P1_U3537) );
  NAND2_X1 U13722 ( .A1(n11297), .A2(n14973), .ZN(n11298) );
  OAI21_X1 U13723 ( .B1(n14973), .B2(n8516), .A(n11298), .ZN(P1_U3486) );
  INV_X1 U13724 ( .A(n11299), .ZN(n11300) );
  NAND2_X1 U13725 ( .A1(n11302), .A2(n10117), .ZN(n11304) );
  AOI22_X1 U13726 ( .A1(n12892), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n12733), 
        .B2(n15031), .ZN(n11303) );
  XNOR2_X1 U13727 ( .A(n14830), .B(n11155), .ZN(n11306) );
  NAND2_X1 U13728 ( .A1(n13266), .A2(n12855), .ZN(n11305) );
  NAND2_X1 U13729 ( .A1(n11306), .A2(n11305), .ZN(n11423) );
  OAI21_X1 U13730 ( .B1(n11306), .B2(n11305), .A(n11423), .ZN(n11307) );
  AOI21_X1 U13731 ( .B1(n11308), .B2(n11307), .A(n6808), .ZN(n11321) );
  NAND2_X1 U13732 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n15033)
         );
  OAI21_X1 U13733 ( .B1(n14799), .B2(n11416), .A(n15033), .ZN(n11319) );
  INV_X1 U13734 ( .A(n13267), .ZN(n11408) );
  NAND2_X1 U13735 ( .A1(n13169), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n11317) );
  INV_X1 U13736 ( .A(n11362), .ZN(n11364) );
  NAND2_X1 U13737 ( .A1(n11311), .A2(n11310), .ZN(n11312) );
  NAND2_X1 U13738 ( .A1(n11364), .A2(n11312), .ZN(n11426) );
  OR2_X1 U13739 ( .A1(n12901), .A2(n11426), .ZN(n11316) );
  OR2_X1 U13740 ( .A1(n12775), .A2(n14829), .ZN(n11315) );
  INV_X1 U13741 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11313) );
  OR2_X1 U13742 ( .A1(n13172), .A2(n11313), .ZN(n11314) );
  NAND4_X1 U13743 ( .A1(n11317), .A2(n11316), .A3(n11315), .A4(n11314), .ZN(
        n14786) );
  INV_X1 U13744 ( .A(n14786), .ZN(n11409) );
  OAI22_X1 U13745 ( .A1(n11408), .A2(n12963), .B1(n12962), .B2(n11409), .ZN(
        n11318) );
  AOI211_X1 U13746 ( .C1(n14830), .C2(n14796), .A(n11319), .B(n11318), .ZN(
        n11320) );
  OAI21_X1 U13747 ( .B1(n11321), .B2(n12967), .A(n11320), .ZN(P2_U3196) );
  INV_X1 U13748 ( .A(n11322), .ZN(n11323) );
  OAI222_X1 U13749 ( .A1(P3_U3151), .A2(n9148), .B1(n12725), .B2(n11324), .C1(
        n11991), .C2(n11323), .ZN(P3_U3270) );
  NAND2_X1 U13750 ( .A1(n11329), .A2(n11325), .ZN(n11326) );
  OAI211_X1 U13751 ( .C1(n11328), .C2(n11336), .A(n11344), .B(n15369), .ZN(
        n11332) );
  OR2_X1 U13752 ( .A1(n11526), .A2(n15351), .ZN(n11331) );
  NAND2_X1 U13753 ( .A1(n12406), .A2(n11329), .ZN(n11330) );
  AND2_X1 U13754 ( .A1(n11331), .A2(n11330), .ZN(n15179) );
  NAND2_X1 U13755 ( .A1(n11332), .A2(n15179), .ZN(n15415) );
  AND2_X1 U13756 ( .A1(n15189), .A2(n14770), .ZN(n15416) );
  AOI22_X1 U13757 ( .A1(n15344), .A2(n15416), .B1(n15379), .B2(n11333), .ZN(
        n11334) );
  OAI21_X1 U13758 ( .B1(n11335), .B2(n15380), .A(n11334), .ZN(n11340) );
  INV_X1 U13759 ( .A(n15417), .ZN(n11338) );
  AND2_X1 U13760 ( .A1(n11337), .A2(n11336), .ZN(n15414) );
  NOR3_X1 U13761 ( .A1(n11338), .A2(n15414), .A3(n12563), .ZN(n11339) );
  AOI211_X1 U13762 ( .C1(n15380), .C2(n15415), .A(n11340), .B(n11339), .ZN(
        n11341) );
  INV_X1 U13763 ( .A(n11341), .ZN(P3_U3223) );
  NAND2_X1 U13764 ( .A1(n15189), .A2(n11342), .ZN(n11343) );
  INV_X1 U13765 ( .A(n11351), .ZN(n11345) );
  XNOR2_X1 U13766 ( .A(n11521), .B(n11345), .ZN(n11347) );
  OAI22_X1 U13767 ( .A1(n11442), .A2(n15353), .B1(n11574), .B2(n15351), .ZN(
        n11346) );
  AOI21_X1 U13768 ( .B1(n11347), .B2(n15369), .A(n11346), .ZN(n14778) );
  NOR2_X1 U13769 ( .A1(n11522), .A2(n15374), .ZN(n14774) );
  INV_X1 U13770 ( .A(n11444), .ZN(n11348) );
  OAI22_X1 U13771 ( .A1(n15380), .A2(n11055), .B1(n11348), .B2(n12555), .ZN(
        n11349) );
  AOI21_X1 U13772 ( .B1(n15344), .B2(n14774), .A(n11349), .ZN(n11356) );
  NAND2_X1 U13773 ( .A1(n15417), .A2(n11350), .ZN(n11352) );
  NAND2_X1 U13774 ( .A1(n11352), .A2(n11351), .ZN(n11354) );
  NAND2_X1 U13775 ( .A1(n11354), .A2(n11353), .ZN(n14776) );
  NAND2_X1 U13776 ( .A1(n14776), .A2(n12581), .ZN(n11355) );
  OAI211_X1 U13777 ( .C1(n14778), .C2(n12443), .A(n11356), .B(n11355), .ZN(
        P3_U3222) );
  INV_X1 U13778 ( .A(n13040), .ZN(n15151) );
  INV_X1 U13779 ( .A(n13266), .ZN(n11371) );
  XNOR2_X1 U13780 ( .A(n14830), .B(n11371), .ZN(n13196) );
  NAND2_X1 U13781 ( .A1(n11358), .A2(n10117), .ZN(n11361) );
  AOI22_X1 U13782 ( .A1(n12892), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n12733), 
        .B2(n11359), .ZN(n11360) );
  XNOR2_X1 U13783 ( .A(n13052), .B(n14786), .ZN(n13197) );
  XNOR2_X1 U13784 ( .A(n11561), .B(n13197), .ZN(n11373) );
  NAND2_X1 U13785 ( .A1(n13169), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n11370) );
  INV_X1 U13786 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n11363) );
  NAND2_X1 U13787 ( .A1(n11364), .A2(n11363), .ZN(n11365) );
  NAND2_X1 U13788 ( .A1(n11546), .A2(n11365), .ZN(n14804) );
  OR2_X1 U13789 ( .A1(n14804), .A2(n12901), .ZN(n11369) );
  OR2_X1 U13790 ( .A1(n12903), .A2(n14821), .ZN(n11368) );
  INV_X1 U13791 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n11366) );
  OR2_X1 U13792 ( .A1(n13172), .A2(n11366), .ZN(n11367) );
  OAI22_X1 U13793 ( .A1(n11371), .A2(n13928), .B1(n13066), .B2(n14784), .ZN(
        n11424) );
  INV_X1 U13794 ( .A(n11424), .ZN(n11372) );
  OAI21_X1 U13795 ( .B1(n11373), .B2(n13925), .A(n11372), .ZN(n14828) );
  INV_X1 U13796 ( .A(n14828), .ZN(n11384) );
  OAI21_X1 U13797 ( .B1(n11414), .B2(n14824), .A(n11374), .ZN(n11375) );
  NOR2_X1 U13798 ( .A1(n11375), .A2(n14811), .ZN(n14826) );
  INV_X1 U13799 ( .A(n11426), .ZN(n11376) );
  AOI22_X1 U13800 ( .A1(n15072), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n15058), 
        .B2(n11376), .ZN(n11377) );
  OAI21_X1 U13801 ( .B1(n14824), .B2(n13959), .A(n11377), .ZN(n11382) );
  AND2_X1 U13802 ( .A1(n11380), .A2(n13197), .ZN(n14822) );
  NOR3_X1 U13803 ( .A1(n14823), .A2(n14822), .A3(n13941), .ZN(n11381) );
  AOI211_X1 U13804 ( .C1(n15068), .C2(n14826), .A(n11382), .B(n11381), .ZN(
        n11383) );
  OAI21_X1 U13805 ( .B1(n11384), .B2(n15072), .A(n11383), .ZN(P2_U3252) );
  OAI22_X1 U13806 ( .A1(n11385), .A2(n14603), .B1(n11386), .B2(n14959), .ZN(
        n11391) );
  INV_X1 U13807 ( .A(n11386), .ZN(n11387) );
  OAI22_X1 U13808 ( .A1(n11388), .A2(n14603), .B1(n11387), .B2(n14959), .ZN(
        n11390) );
  MUX2_X1 U13809 ( .A(n11391), .B(n11390), .S(n11389), .Z(n11394) );
  NAND2_X1 U13810 ( .A1(n14243), .A2(n14539), .ZN(n11393) );
  NAND2_X1 U13811 ( .A1(n14241), .A2(n14540), .ZN(n11392) );
  NAND2_X1 U13812 ( .A1(n11393), .A2(n11392), .ZN(n14854) );
  NOR2_X1 U13813 ( .A1(n11394), .A2(n14854), .ZN(n14867) );
  OAI22_X1 U13814 ( .A1(n14531), .A2(n11395), .B1(n14858), .B2(n14498), .ZN(
        n11399) );
  NAND2_X1 U13815 ( .A1(n14843), .A2(n11396), .ZN(n11397) );
  NAND3_X1 U13816 ( .A1(n14710), .A2(n14712), .A3(n11397), .ZN(n14866) );
  NOR2_X1 U13817 ( .A1(n14866), .A2(n14529), .ZN(n11398) );
  AOI211_X1 U13818 ( .C1(n14706), .C2(n14843), .A(n11399), .B(n11398), .ZN(
        n11400) );
  OAI21_X1 U13819 ( .B1(n14867), .B2(n14705), .A(n11400), .ZN(P1_U3282) );
  INV_X1 U13820 ( .A(n12783), .ZN(n11405) );
  NAND2_X1 U13821 ( .A1(n14666), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n11402) );
  OAI211_X1 U13822 ( .C1(n11405), .C2(n14668), .A(n11402), .B(n11401), .ZN(
        P1_U3332) );
  NAND2_X1 U13823 ( .A1(n14071), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n11404) );
  OR2_X1 U13824 ( .A1(n11403), .A2(P2_U3088), .ZN(n13257) );
  OAI211_X1 U13825 ( .C1(n11405), .C2(n6618), .A(n11404), .B(n13257), .ZN(
        P2_U3304) );
  XNOR2_X1 U13826 ( .A(n11406), .B(n13196), .ZN(n11407) );
  OAI222_X1 U13827 ( .A1(n14784), .A2(n11409), .B1(n13928), .B2(n11408), .C1(
        n13925), .C2(n11407), .ZN(n14833) );
  INV_X1 U13828 ( .A(n14833), .ZN(n11422) );
  XNOR2_X1 U13829 ( .A(n11411), .B(n11410), .ZN(n14835) );
  NAND2_X1 U13830 ( .A1(n11412), .A2(n14830), .ZN(n11413) );
  NAND2_X1 U13831 ( .A1(n11413), .A2(n11374), .ZN(n11415) );
  OR2_X1 U13832 ( .A1(n11415), .A2(n11414), .ZN(n14831) );
  INV_X1 U13833 ( .A(n11416), .ZN(n11417) );
  AOI22_X1 U13834 ( .A1(n15072), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n15058), 
        .B2(n11417), .ZN(n11419) );
  NAND2_X1 U13835 ( .A1(n14830), .A2(n15060), .ZN(n11418) );
  OAI211_X1 U13836 ( .C1(n14831), .C2(n13937), .A(n11419), .B(n11418), .ZN(
        n11420) );
  AOI21_X1 U13837 ( .B1(n14835), .B2(n15069), .A(n11420), .ZN(n11421) );
  OAI21_X1 U13838 ( .B1(n11422), .B2(n15072), .A(n11421), .ZN(P2_U3253) );
  XNOR2_X1 U13839 ( .A(n13052), .B(n12895), .ZN(n11621) );
  NAND2_X1 U13840 ( .A1(n14786), .A2(n6611), .ZN(n11620) );
  XNOR2_X1 U13841 ( .A(n11621), .B(n11620), .ZN(n11623) );
  XNOR2_X1 U13842 ( .A(n11624), .B(n11623), .ZN(n11429) );
  AOI22_X1 U13843 ( .A1(n11424), .A2(n14795), .B1(P2_REG3_REG_13__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11425) );
  OAI21_X1 U13844 ( .B1(n11426), .B2(n14799), .A(n11425), .ZN(n11427) );
  AOI21_X1 U13845 ( .B1(n13052), .B2(n14796), .A(n11427), .ZN(n11428) );
  OAI21_X1 U13846 ( .B1(n11429), .B2(n12967), .A(n11428), .ZN(P2_U3206) );
  INV_X1 U13847 ( .A(n11430), .ZN(n11431) );
  OAI222_X1 U13848 ( .A1(P3_U3151), .A2(n11433), .B1(n12725), .B2(n11432), 
        .C1(n11991), .C2(n11431), .ZN(P3_U3269) );
  INV_X1 U13849 ( .A(n11451), .ZN(n11439) );
  INV_X1 U13850 ( .A(n11434), .ZN(n11436) );
  OAI21_X1 U13851 ( .B1(n11436), .B2(n11435), .A(n12238), .ZN(n11437) );
  OAI21_X1 U13852 ( .B1(n11439), .B2(n11438), .A(n11437), .ZN(n11440) );
  NAND2_X1 U13853 ( .A1(n11440), .A2(n15193), .ZN(n11446) );
  AOI22_X1 U13854 ( .A1(n12169), .A2(n12237), .B1(P3_REG3_REG_11__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11441) );
  OAI21_X1 U13855 ( .B1(n11442), .B2(n12222), .A(n11441), .ZN(n11443) );
  AOI21_X1 U13856 ( .B1(n11444), .B2(n12227), .A(n11443), .ZN(n11445) );
  OAI211_X1 U13857 ( .C1(n12230), .C2(n11522), .A(n11446), .B(n11445), .ZN(
        P3_U3176) );
  INV_X1 U13858 ( .A(n12796), .ZN(n12135) );
  OAI222_X1 U13859 ( .A1(n11987), .A2(n11448), .B1(n6618), .B2(n12135), .C1(
        n11447), .C2(P2_U3088), .ZN(P2_U3303) );
  INV_X1 U13860 ( .A(n11570), .ZN(n11702) );
  OAI21_X1 U13861 ( .B1(n11451), .B2(n11450), .A(n11449), .ZN(n11452) );
  NAND2_X1 U13862 ( .A1(n11452), .A2(n15193), .ZN(n11456) );
  AOI22_X1 U13863 ( .A1(n12169), .A2(n12236), .B1(P3_REG3_REG_12__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11453) );
  OAI21_X1 U13864 ( .B1(n11526), .B2(n12222), .A(n11453), .ZN(n11454) );
  AOI21_X1 U13865 ( .B1(n11528), .B2(n12227), .A(n11454), .ZN(n11455) );
  OAI211_X1 U13866 ( .C1(n11702), .C2(n12230), .A(n11456), .B(n11455), .ZN(
        P3_U3164) );
  XNOR2_X1 U13867 ( .A(n11457), .B(n11460), .ZN(n11459) );
  AOI22_X1 U13868 ( .A1(n14539), .A2(n14241), .B1(n14239), .B2(n14540), .ZN(
        n11933) );
  INV_X1 U13869 ( .A(n11933), .ZN(n11458) );
  AOI21_X1 U13870 ( .B1(n11459), .B2(n14701), .A(n11458), .ZN(n14861) );
  XNOR2_X1 U13871 ( .A(n11461), .B(n11460), .ZN(n14864) );
  OAI211_X1 U13872 ( .C1(n14711), .C2(n14860), .A(n11608), .B(n14712), .ZN(
        n14859) );
  AOI22_X1 U13873 ( .A1(n14705), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n11935), 
        .B2(n14703), .ZN(n11463) );
  NAND2_X1 U13874 ( .A1(n11928), .A2(n14706), .ZN(n11462) );
  OAI211_X1 U13875 ( .C1(n14859), .C2(n14529), .A(n11463), .B(n11462), .ZN(
        n11464) );
  AOI21_X1 U13876 ( .B1(n14864), .B2(n14717), .A(n11464), .ZN(n11465) );
  OAI21_X1 U13877 ( .B1(n14861), .B2(n14705), .A(n11465), .ZN(P1_U3280) );
  NOR2_X1 U13878 ( .A1(n11476), .A2(n13677), .ZN(n11466) );
  OAI21_X1 U13879 ( .B1(n11468), .B2(n12260), .A(n12254), .ZN(n11470) );
  INV_X1 U13880 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n11469) );
  AOI21_X1 U13881 ( .B1(n11470), .B2(n11469), .A(n12255), .ZN(n11487) );
  INV_X1 U13882 ( .A(n12260), .ZN(n12249) );
  NAND2_X1 U13883 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n11472), .ZN(n12261) );
  OAI21_X1 U13884 ( .B1(n11472), .B2(P3_REG1_REG_13__SCAN_IN), .A(n12261), 
        .ZN(n11485) );
  MUX2_X1 U13885 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n14735), .Z(n12246) );
  XNOR2_X1 U13886 ( .A(n12246), .B(n12260), .ZN(n11478) );
  INV_X1 U13887 ( .A(n11473), .ZN(n11475) );
  OAI21_X1 U13888 ( .B1(n11476), .B2(n11475), .A(n11474), .ZN(n11477) );
  NOR2_X1 U13889 ( .A1(n11477), .A2(n11478), .ZN(n12247) );
  AOI21_X1 U13890 ( .B1(n11478), .B2(n11477), .A(n12247), .ZN(n11483) );
  INV_X1 U13891 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n11479) );
  NOR2_X1 U13892 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11479), .ZN(n11481) );
  NOR2_X1 U13893 ( .A1(n15308), .A2(n13716), .ZN(n11480) );
  AOI211_X1 U13894 ( .C1(n15266), .C2(n12249), .A(n11481), .B(n11480), .ZN(
        n11482) );
  OAI21_X1 U13895 ( .B1(n11483), .B2(n15322), .A(n11482), .ZN(n11484) );
  AOI21_X1 U13896 ( .B1(n15329), .B2(n11485), .A(n11484), .ZN(n11486) );
  OAI21_X1 U13897 ( .B1(n11487), .B2(n15333), .A(n11486), .ZN(P3_U3195) );
  INV_X1 U13898 ( .A(n13310), .ZN(n13305) );
  AND2_X1 U13899 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n11843) );
  INV_X1 U13900 ( .A(n15050), .ZN(n11584) );
  AOI21_X1 U13901 ( .B1(n11539), .B2(P2_REG1_REG_14__SCAN_IN), .A(n11488), 
        .ZN(n11489) );
  NOR2_X1 U13902 ( .A1(n11489), .A2(n11497), .ZN(n11490) );
  INV_X1 U13903 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n13298) );
  XNOR2_X1 U13904 ( .A(n11497), .B(n11489), .ZN(n13299) );
  NOR2_X1 U13905 ( .A1(n13298), .A2(n13299), .ZN(n13297) );
  NOR2_X1 U13906 ( .A1(n11490), .A2(n13297), .ZN(n15040) );
  XNOR2_X1 U13907 ( .A(n11584), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n15039) );
  NOR2_X1 U13908 ( .A1(n15040), .A2(n15039), .ZN(n15038) );
  AOI21_X1 U13909 ( .B1(n11584), .B2(P2_REG1_REG_16__SCAN_IN), .A(n15038), 
        .ZN(n11492) );
  XNOR2_X1 U13910 ( .A(n13305), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n11491) );
  NOR2_X1 U13911 ( .A1(n11491), .A2(n11492), .ZN(n13304) );
  AOI211_X1 U13912 ( .C1(n11492), .C2(n11491), .A(n13304), .B(n15037), .ZN(
        n11493) );
  AOI211_X1 U13913 ( .C1(n13305), .C2(n15032), .A(n11843), .B(n11493), .ZN(
        n11506) );
  INV_X1 U13914 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13505) );
  XNOR2_X1 U13915 ( .A(n15050), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n15046) );
  NOR2_X1 U13916 ( .A1(n11539), .A2(n11494), .ZN(n11496) );
  NOR2_X1 U13917 ( .A1(n11496), .A2(n11495), .ZN(n11498) );
  NAND2_X1 U13918 ( .A1(n13296), .A2(n11498), .ZN(n11499) );
  XNOR2_X1 U13919 ( .A(n11498), .B(n11497), .ZN(n13294) );
  NAND2_X1 U13920 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n13294), .ZN(n13293) );
  NAND2_X1 U13921 ( .A1(n11499), .A2(n13293), .ZN(n15047) );
  NAND2_X1 U13922 ( .A1(n15046), .A2(n15047), .ZN(n15044) );
  OAI21_X1 U13923 ( .B1(n15050), .B2(n13505), .A(n15044), .ZN(n11504) );
  NAND2_X1 U13924 ( .A1(n13310), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n11500) );
  OAI21_X1 U13925 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n13310), .A(n11500), 
        .ZN(n11503) );
  INV_X1 U13926 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n11502) );
  NAND2_X1 U13927 ( .A1(n13310), .A2(n11502), .ZN(n11501) );
  OAI211_X1 U13928 ( .C1(n13310), .C2(n11502), .A(n11504), .B(n11501), .ZN(
        n13309) );
  OAI211_X1 U13929 ( .C1(n11504), .C2(n11503), .A(n15045), .B(n13309), .ZN(
        n11505) );
  OAI211_X1 U13930 ( .C1(n14730), .C2(n15035), .A(n11506), .B(n11505), .ZN(
        P2_U3231) );
  XNOR2_X1 U13931 ( .A(n11507), .B(n11709), .ZN(n11508) );
  XNOR2_X1 U13932 ( .A(n11509), .B(n11508), .ZN(n11514) );
  AOI22_X1 U13933 ( .A1(n12212), .A2(n12237), .B1(P3_REG3_REG_13__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11510) );
  OAI21_X1 U13934 ( .B1(n11711), .B2(n12224), .A(n11510), .ZN(n11512) );
  NOR2_X1 U13935 ( .A1(n11798), .A2(n12230), .ZN(n11511) );
  AOI211_X1 U13936 ( .C1(n11577), .C2(n12227), .A(n11512), .B(n11511), .ZN(
        n11513) );
  OAI21_X1 U13937 ( .B1(n11514), .B2(n15207), .A(n11513), .ZN(P3_U3174) );
  INV_X1 U13938 ( .A(n12811), .ZN(n11518) );
  OAI222_X1 U13939 ( .A1(n12137), .A2(n11516), .B1(n14668), .B2(n11518), .C1(
        n11515), .C2(P1_U3086), .ZN(P1_U3330) );
  OAI222_X1 U13940 ( .A1(n11987), .A2(n11519), .B1(n6618), .B2(n11518), .C1(
        n11517), .C2(P2_U3088), .ZN(P2_U3302) );
  NAND2_X1 U13941 ( .A1(n11522), .A2(n11526), .ZN(n11520) );
  NAND2_X1 U13942 ( .A1(n11521), .A2(n11520), .ZN(n11524) );
  OR2_X1 U13943 ( .A1(n11522), .A2(n11526), .ZN(n11523) );
  XNOR2_X1 U13944 ( .A(n6847), .B(n11568), .ZN(n11525) );
  OAI222_X1 U13945 ( .A1(n15351), .A2(n11709), .B1(n15353), .B2(n11526), .C1(
        n11525), .C2(n15359), .ZN(n11697) );
  INV_X1 U13946 ( .A(n11697), .ZN(n11532) );
  XNOR2_X1 U13947 ( .A(n11527), .B(n7202), .ZN(n11698) );
  AOI22_X1 U13948 ( .A1(n12443), .A2(P3_REG2_REG_12__SCAN_IN), .B1(n15379), 
        .B2(n11528), .ZN(n11529) );
  OAI21_X1 U13949 ( .B1(n12578), .B2(n11702), .A(n11529), .ZN(n11530) );
  AOI21_X1 U13950 ( .B1(n11698), .B2(n12581), .A(n11530), .ZN(n11531) );
  OAI21_X1 U13951 ( .B1(n11532), .B2(n12443), .A(n11531), .ZN(P3_U3221) );
  INV_X1 U13952 ( .A(n11533), .ZN(n11535) );
  OAI222_X1 U13953 ( .A1(P3_U3151), .A2(n14735), .B1(n11991), .B2(n11535), 
        .C1(n11534), .C2(n11995), .ZN(P3_U3268) );
  OAI222_X1 U13954 ( .A1(P3_U3151), .A2(n12354), .B1(n11991), .B2(n11537), 
        .C1(n11536), .C2(n12725), .ZN(P3_U3267) );
  INV_X1 U13955 ( .A(n13066), .ZN(n13265) );
  NAND2_X1 U13956 ( .A1(n11538), .A2(n10117), .ZN(n11541) );
  AOI22_X1 U13957 ( .A1(n12892), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n11539), 
        .B2(n12733), .ZN(n11540) );
  XNOR2_X1 U13958 ( .A(n7081), .B(n13265), .ZN(n14800) );
  INV_X1 U13959 ( .A(n14800), .ZN(n14807) );
  NAND2_X1 U13960 ( .A1(n11542), .A2(n10117), .ZN(n11544) );
  AOI22_X1 U13961 ( .A1(n13296), .A2(n12733), .B1(n12892), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n11543) );
  INV_X1 U13962 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n11545) );
  NAND2_X1 U13963 ( .A1(n11546), .A2(n11545), .ZN(n11547) );
  AND2_X1 U13964 ( .A1(n11556), .A2(n11547), .ZN(n11633) );
  INV_X1 U13965 ( .A(n12901), .ZN(n12754) );
  NAND2_X1 U13966 ( .A1(n11633), .A2(n12754), .ZN(n11554) );
  INV_X1 U13967 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n11548) );
  OR2_X1 U13968 ( .A1(n13172), .A2(n11548), .ZN(n11551) );
  INV_X1 U13969 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n11549) );
  OR2_X1 U13970 ( .A1(n12845), .A2(n11549), .ZN(n11550) );
  AND2_X1 U13971 ( .A1(n11551), .A2(n11550), .ZN(n11553) );
  OR2_X1 U13972 ( .A1(n12775), .A2(n13298), .ZN(n11552) );
  XNOR2_X1 U13973 ( .A(n14048), .B(n13264), .ZN(n13204) );
  XNOR2_X1 U13974 ( .A(n11596), .B(n13204), .ZN(n14050) );
  INV_X1 U13975 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n11560) );
  INV_X1 U13976 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n11555) );
  INV_X1 U13977 ( .A(n11587), .ZN(n11589) );
  NAND2_X1 U13978 ( .A1(n11556), .A2(n11555), .ZN(n11557) );
  NAND2_X1 U13979 ( .A1(n11589), .A2(n11557), .ZN(n11600) );
  OR2_X1 U13980 ( .A1(n11600), .A2(n12901), .ZN(n11559) );
  AOI22_X1 U13981 ( .A1(n12900), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n13169), 
        .B2(P2_REG0_REG_16__SCAN_IN), .ZN(n11558) );
  OAI211_X1 U13982 ( .C1(n12903), .C2(n11560), .A(n11559), .B(n11558), .ZN(
        n13263) );
  XNOR2_X1 U13983 ( .A(n11582), .B(n13204), .ZN(n11562) );
  OAI222_X1 U13984 ( .A1(n14784), .A2(n11751), .B1(n13928), .B2(n13066), .C1(
        n13925), .C2(n11562), .ZN(n14046) );
  NAND2_X1 U13985 ( .A1(n14046), .A2(n13944), .ZN(n11567) );
  OR2_X1 U13986 ( .A1(n14809), .A2(n13064), .ZN(n11563) );
  AND3_X1 U13987 ( .A1(n11598), .A2(n11563), .A3(n11374), .ZN(n14047) );
  AOI22_X1 U13988 ( .A1(n15072), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n15058), 
        .B2(n11633), .ZN(n11564) );
  OAI21_X1 U13989 ( .B1(n13064), .B2(n13959), .A(n11564), .ZN(n11565) );
  AOI21_X1 U13990 ( .B1(n14047), .B2(n15068), .A(n11565), .ZN(n11566) );
  OAI211_X1 U13991 ( .C1(n13941), .C2(n14050), .A(n11567), .B(n11566), .ZN(
        P2_U3250) );
  NAND2_X1 U13992 ( .A1(n11570), .A2(n12237), .ZN(n11705) );
  NAND2_X1 U13993 ( .A1(n11708), .A2(n11705), .ZN(n11572) );
  XNOR2_X1 U13994 ( .A(n11572), .B(n11571), .ZN(n11573) );
  OAI222_X1 U13995 ( .A1(n15351), .A2(n11711), .B1(n15353), .B2(n11574), .C1(
        n11573), .C2(n15359), .ZN(n11792) );
  INV_X1 U13996 ( .A(n11792), .ZN(n11581) );
  XNOR2_X1 U13997 ( .A(n11576), .B(n11575), .ZN(n11793) );
  AOI22_X1 U13998 ( .A1(n12443), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n15379), 
        .B2(n11577), .ZN(n11578) );
  OAI21_X1 U13999 ( .B1(n11798), .B2(n12578), .A(n11578), .ZN(n11579) );
  AOI21_X1 U14000 ( .B1(n11793), .B2(n12581), .A(n11579), .ZN(n11580) );
  OAI21_X1 U14001 ( .B1(n11581), .B2(n12443), .A(n11580), .ZN(P3_U3220) );
  INV_X1 U14002 ( .A(n13204), .ZN(n11595) );
  NAND2_X1 U14003 ( .A1(n11583), .A2(n10117), .ZN(n11586) );
  AOI22_X1 U14004 ( .A1(n12892), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n12733), 
        .B2(n11584), .ZN(n11585) );
  XNOR2_X1 U14005 ( .A(n14042), .B(n11751), .ZN(n13201) );
  INV_X1 U14006 ( .A(n13201), .ZN(n11737) );
  XNOR2_X1 U14007 ( .A(n7546), .B(n11737), .ZN(n11594) );
  INV_X1 U14008 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n11593) );
  NAND2_X1 U14009 ( .A1(n11587), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n11743) );
  INV_X1 U14010 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n11588) );
  NAND2_X1 U14011 ( .A1(n11589), .A2(n11588), .ZN(n11590) );
  NAND2_X1 U14012 ( .A1(n11743), .A2(n11590), .ZN(n11842) );
  OR2_X1 U14013 ( .A1(n11842), .A2(n12901), .ZN(n11592) );
  AOI22_X1 U14014 ( .A1(n12900), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13169), 
        .B2(P2_REG0_REG_17__SCAN_IN), .ZN(n11591) );
  OAI211_X1 U14015 ( .C1(n12903), .C2(n11593), .A(n11592), .B(n11591), .ZN(
        n13262) );
  AOI222_X1 U14016 ( .A1(n15054), .A2(n11594), .B1(n13262), .B2(n13949), .C1(
        n13264), .C2(n14787), .ZN(n14044) );
  NAND2_X1 U14017 ( .A1(n11597), .A2(n13201), .ZN(n11752) );
  OAI21_X1 U14018 ( .B1(n11597), .B2(n13201), .A(n11752), .ZN(n14045) );
  INV_X1 U14019 ( .A(n14045), .ZN(n11604) );
  AOI21_X1 U14020 ( .B1(n11598), .B2(n14042), .A(n6611), .ZN(n11599) );
  AND2_X1 U14021 ( .A1(n11599), .A2(n11755), .ZN(n14041) );
  NAND2_X1 U14022 ( .A1(n14041), .A2(n15068), .ZN(n11602) );
  INV_X1 U14023 ( .A(n11600), .ZN(n11785) );
  AOI22_X1 U14024 ( .A1(n15072), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n15058), 
        .B2(n11785), .ZN(n11601) );
  OAI211_X1 U14025 ( .C1(n7079), .C2(n13959), .A(n11602), .B(n11601), .ZN(
        n11603) );
  AOI21_X1 U14026 ( .B1(n11604), .B2(n15069), .A(n11603), .ZN(n11605) );
  OAI21_X1 U14027 ( .B1(n14044), .B2(n15072), .A(n11605), .ZN(P2_U3249) );
  XOR2_X1 U14028 ( .A(n11606), .B(n11611), .Z(n11607) );
  AOI222_X1 U14029 ( .A1(n14701), .A2(n11607), .B1(n14240), .B2(n14539), .C1(
        n14238), .C2(n14540), .ZN(n14641) );
  AOI211_X1 U14030 ( .C1(n14639), .C2(n11608), .A(n14503), .B(n11825), .ZN(
        n14638) );
  INV_X1 U14031 ( .A(n14639), .ZN(n11610) );
  AOI22_X1 U14032 ( .A1(n14705), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n14098), 
        .B2(n14703), .ZN(n11609) );
  OAI21_X1 U14033 ( .B1(n11610), .B2(n14506), .A(n11609), .ZN(n11616) );
  NAND2_X1 U14034 ( .A1(n11612), .A2(n11611), .ZN(n11613) );
  NAND2_X1 U14035 ( .A1(n11614), .A2(n11613), .ZN(n14642) );
  NOR2_X1 U14036 ( .A1(n14642), .A2(n14511), .ZN(n11615) );
  AOI211_X1 U14037 ( .C1(n14638), .C2(n14716), .A(n11616), .B(n11615), .ZN(
        n11617) );
  OAI21_X1 U14038 ( .B1(n14641), .B2(n14705), .A(n11617), .ZN(P1_U3279) );
  NOR2_X1 U14039 ( .A1(n14785), .A2(n15065), .ZN(n11619) );
  XNOR2_X1 U14040 ( .A(n13064), .B(n11155), .ZN(n11618) );
  NOR2_X1 U14041 ( .A1(n11618), .A2(n11619), .ZN(n11778) );
  AOI21_X1 U14042 ( .B1(n11619), .B2(n11618), .A(n11778), .ZN(n11630) );
  INV_X1 U14043 ( .A(n11620), .ZN(n11622) );
  NOR2_X1 U14044 ( .A1(n13066), .A2(n15065), .ZN(n11626) );
  XNOR2_X1 U14045 ( .A(n14816), .B(n11155), .ZN(n11625) );
  NOR2_X1 U14046 ( .A1(n11625), .A2(n11626), .ZN(n11627) );
  AOI21_X1 U14047 ( .B1(n11626), .B2(n11625), .A(n11627), .ZN(n14792) );
  INV_X1 U14048 ( .A(n11627), .ZN(n11628) );
  NAND2_X1 U14049 ( .A1(n14790), .A2(n11628), .ZN(n11629) );
  NAND2_X1 U14050 ( .A1(n11629), .A2(n11630), .ZN(n11780) );
  OAI21_X1 U14051 ( .B1(n11630), .B2(n11629), .A(n11780), .ZN(n11631) );
  NAND2_X1 U14052 ( .A1(n11631), .A2(n14793), .ZN(n11635) );
  AND2_X1 U14053 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3088), .ZN(n13295) );
  OAI22_X1 U14054 ( .A1(n13066), .A2(n12963), .B1(n12962), .B2(n11751), .ZN(
        n11632) );
  AOI211_X1 U14055 ( .C1(n11633), .C2(n11786), .A(n13295), .B(n11632), .ZN(
        n11634) );
  OAI211_X1 U14056 ( .C1(n13064), .C2(n11848), .A(n11635), .B(n11634), .ZN(
        P2_U3213) );
  NAND2_X1 U14057 ( .A1(n11644), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11640) );
  INV_X1 U14058 ( .A(n11636), .ZN(n11637) );
  NAND2_X1 U14059 ( .A1(n11638), .A2(n11637), .ZN(n11639) );
  NAND2_X1 U14060 ( .A1(n11640), .A2(n11639), .ZN(n11641) );
  NOR2_X1 U14061 ( .A1(n11646), .A2(n11641), .ZN(n11642) );
  XOR2_X1 U14062 ( .A(n11641), .B(n14922), .Z(n14916) );
  NOR2_X1 U14063 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14916), .ZN(n14915) );
  NOR2_X1 U14064 ( .A1(n11642), .A2(n14915), .ZN(n14292) );
  INV_X1 U14065 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11895) );
  XNOR2_X1 U14066 ( .A(n14297), .B(n11895), .ZN(n14291) );
  XNOR2_X1 U14067 ( .A(n14292), .B(n14291), .ZN(n11653) );
  INV_X1 U14068 ( .A(n14921), .ZN(n14303) );
  NAND2_X1 U14069 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14149)
         );
  OAI21_X1 U14070 ( .B1(n14926), .B2(n9316), .A(n14149), .ZN(n11651) );
  NAND2_X1 U14071 ( .A1(n14922), .A2(n11645), .ZN(n11647) );
  INV_X1 U14072 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14911) );
  NAND2_X1 U14073 ( .A1(n14912), .A2(n14911), .ZN(n14910) );
  NAND2_X1 U14074 ( .A1(n11647), .A2(n14910), .ZN(n11649) );
  XNOR2_X1 U14075 ( .A(n14297), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n11648) );
  AOI211_X1 U14076 ( .C1(n11649), .C2(n11648), .A(n14298), .B(n14296), .ZN(
        n11650) );
  AOI211_X1 U14077 ( .C1(n14303), .C2(n14297), .A(n11651), .B(n11650), .ZN(
        n11652) );
  OAI21_X1 U14078 ( .B1(n14917), .B2(n11653), .A(n11652), .ZN(P1_U3259) );
  AOI22_X1 U14079 ( .A1(n14956), .A2(n12073), .B1(n12119), .B2(n14245), .ZN(
        n11669) );
  NAND2_X1 U14080 ( .A1(n14956), .A2(n12120), .ZN(n11655) );
  NAND2_X1 U14081 ( .A1(n14245), .A2(n12112), .ZN(n11654) );
  NAND2_X1 U14082 ( .A1(n11655), .A2(n11654), .ZN(n11656) );
  XNOR2_X1 U14083 ( .A(n11656), .B(n12121), .ZN(n11667) );
  INV_X1 U14084 ( .A(n11667), .ZN(n11668) );
  NOR2_X1 U14085 ( .A1(n11657), .A2(n12062), .ZN(n11658) );
  AOI21_X1 U14086 ( .B1(n14954), .B2(n12073), .A(n11658), .ZN(n11666) );
  NAND2_X1 U14087 ( .A1(n14954), .A2(n12120), .ZN(n11660) );
  NAND2_X1 U14088 ( .A1(n14246), .A2(n12112), .ZN(n11659) );
  NAND2_X1 U14089 ( .A1(n11660), .A2(n11659), .ZN(n11661) );
  XNOR2_X1 U14090 ( .A(n11661), .B(n12121), .ZN(n11664) );
  INV_X1 U14091 ( .A(n11664), .ZN(n11665) );
  XNOR2_X1 U14092 ( .A(n11664), .B(n11666), .ZN(n14076) );
  XOR2_X1 U14093 ( .A(n11669), .B(n11667), .Z(n11957) );
  NOR2_X1 U14094 ( .A1(n11681), .A2(n12062), .ZN(n11670) );
  AOI21_X1 U14095 ( .B1(n11671), .B2(n12054), .A(n11670), .ZN(n11673) );
  AOI22_X1 U14096 ( .A1(n11671), .A2(n12120), .B1(n12073), .B2(n14244), .ZN(
        n11672) );
  XNOR2_X1 U14097 ( .A(n11672), .B(n12121), .ZN(n14894) );
  NAND2_X1 U14098 ( .A1(n14964), .A2(n12120), .ZN(n11675) );
  NAND2_X1 U14099 ( .A1(n14243), .A2(n12112), .ZN(n11674) );
  NAND2_X1 U14100 ( .A1(n11675), .A2(n11674), .ZN(n11676) );
  XNOR2_X1 U14101 ( .A(n11676), .B(n12121), .ZN(n11899) );
  NOR2_X1 U14102 ( .A1(n14898), .A2(n12062), .ZN(n11677) );
  AOI21_X1 U14103 ( .B1(n14964), .B2(n12073), .A(n11677), .ZN(n11901) );
  XNOR2_X1 U14104 ( .A(n11899), .B(n11901), .ZN(n11678) );
  NAND2_X1 U14105 ( .A1(n11679), .A2(n11678), .ZN(n11900) );
  OAI211_X1 U14106 ( .C1(n11679), .C2(n11678), .A(n11900), .B(n14904), .ZN(
        n11686) );
  OAI22_X1 U14107 ( .A1(n11681), .A2(n14900), .B1(n14899), .B2(n11680), .ZN(
        n11682) );
  AOI211_X1 U14108 ( .C1(n11684), .C2(n14228), .A(n11683), .B(n11682), .ZN(
        n11685) );
  OAI211_X1 U14109 ( .C1(n11687), .C2(n14896), .A(n11686), .B(n11685), .ZN(
        P1_U3217) );
  XOR2_X1 U14110 ( .A(n11689), .B(n11688), .Z(n11690) );
  NAND2_X1 U14111 ( .A1(n11690), .A2(n15193), .ZN(n11696) );
  OR2_X1 U14112 ( .A1(n11709), .A2(n15353), .ZN(n11692) );
  OR2_X1 U14113 ( .A1(n11727), .A2(n15351), .ZN(n11691) );
  NAND2_X1 U14114 ( .A1(n11692), .A2(n11691), .ZN(n11766) );
  NAND2_X1 U14115 ( .A1(n11766), .A2(n12158), .ZN(n11693) );
  OAI21_X1 U14116 ( .B1(P3_STATE_REG_SCAN_IN), .B2(n7871), .A(n11693), .ZN(
        n11694) );
  AOI21_X1 U14117 ( .B1(n12227), .B2(n11771), .A(n11694), .ZN(n11695) );
  OAI211_X1 U14118 ( .C1(n12230), .C2(n12711), .A(n11696), .B(n11695), .ZN(
        P3_U3155) );
  AOI21_X1 U14119 ( .B1(n11698), .B2(n14775), .A(n11697), .ZN(n11700) );
  MUX2_X1 U14120 ( .A(n13689), .B(n11700), .S(n15436), .Z(n11699) );
  OAI21_X1 U14121 ( .B1(n11702), .B2(n12651), .A(n11699), .ZN(P3_U3471) );
  INV_X1 U14122 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n13706) );
  MUX2_X1 U14123 ( .A(n13706), .B(n11700), .S(n12707), .Z(n11701) );
  OAI21_X1 U14124 ( .B1(n11702), .B2(n12712), .A(n11701), .ZN(P3_U3426) );
  INV_X1 U14125 ( .A(n12829), .ZN(n11725) );
  OAI222_X1 U14126 ( .A1(n11704), .A2(P2_U3088), .B1(n6618), .B2(n11725), .C1(
        n11703), .C2(n11987), .ZN(P2_U3301) );
  OR2_X1 U14127 ( .A1(n11798), .A2(n11709), .ZN(n11706) );
  AND2_X1 U14128 ( .A1(n11706), .A2(n11705), .ZN(n11707) );
  INV_X1 U14129 ( .A(n11710), .ZN(n11712) );
  OR2_X1 U14130 ( .A1(n11769), .A2(n11712), .ZN(n12363) );
  OR2_X1 U14131 ( .A1(n12711), .A2(n11711), .ZN(n11713) );
  OR2_X1 U14132 ( .A1(n11712), .A2(n11713), .ZN(n11800) );
  AND2_X1 U14133 ( .A1(n11802), .A2(n11800), .ZN(n11715) );
  OR2_X1 U14134 ( .A1(n12566), .A2(n11769), .ZN(n11764) );
  NAND3_X1 U14135 ( .A1(n11764), .A2(n11712), .A3(n11713), .ZN(n11714) );
  NAND3_X1 U14136 ( .A1(n11715), .A2(n15369), .A3(n11714), .ZN(n11718) );
  NAND2_X1 U14137 ( .A1(n12406), .A2(n12235), .ZN(n11717) );
  NAND2_X1 U14138 ( .A1(n15366), .A2(n12570), .ZN(n11716) );
  AND2_X1 U14139 ( .A1(n11717), .A2(n11716), .ZN(n11731) );
  NAND2_X1 U14140 ( .A1(n11718), .A2(n11731), .ZN(n12643) );
  INV_X1 U14141 ( .A(n12643), .ZN(n11724) );
  OAI21_X1 U14142 ( .B1(n11720), .B2(n11712), .A(n11719), .ZN(n12644) );
  INV_X1 U14143 ( .A(n11799), .ZN(n12706) );
  AOI22_X1 U14144 ( .A1(n12443), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15379), 
        .B2(n11734), .ZN(n11721) );
  OAI21_X1 U14145 ( .B1(n12706), .B2(n12578), .A(n11721), .ZN(n11722) );
  AOI21_X1 U14146 ( .B1(n12644), .B2(n12581), .A(n11722), .ZN(n11723) );
  OAI21_X1 U14147 ( .B1(n11724), .B2(n12443), .A(n11723), .ZN(P3_U3218) );
  OAI222_X1 U14148 ( .A1(n12137), .A2(n13524), .B1(P1_U3086), .B2(n11726), 
        .C1(n14668), .C2(n11725), .ZN(P1_U3329) );
  XNOR2_X1 U14149 ( .A(n11728), .B(n11727), .ZN(n11729) );
  XNOR2_X1 U14150 ( .A(n11730), .B(n11729), .ZN(n11736) );
  OAI22_X1 U14151 ( .A1(n11731), .A2(n15203), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12279), .ZN(n11733) );
  NOR2_X1 U14152 ( .A1(n12706), .A2(n12230), .ZN(n11732) );
  AOI211_X1 U14153 ( .C1(n11734), .C2(n12227), .A(n11733), .B(n11732), .ZN(
        n11735) );
  OAI21_X1 U14154 ( .B1(n11736), .B2(n15207), .A(n11735), .ZN(P3_U3181) );
  NAND2_X1 U14155 ( .A1(n11739), .A2(n10117), .ZN(n11741) );
  AOI22_X1 U14156 ( .A1(n12892), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n12733), 
        .B2(n13305), .ZN(n11740) );
  XNOR2_X1 U14157 ( .A(n14037), .B(n13262), .ZN(n13202) );
  INV_X1 U14158 ( .A(n13202), .ZN(n11753) );
  XNOR2_X1 U14159 ( .A(n13362), .B(n11753), .ZN(n11750) );
  INV_X1 U14160 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n11742) );
  NAND2_X1 U14161 ( .A1(n11743), .A2(n11742), .ZN(n11744) );
  NAND2_X1 U14162 ( .A1(n11871), .A2(n11744), .ZN(n13933) );
  OR2_X1 U14163 ( .A1(n13933), .A2(n12901), .ZN(n11749) );
  INV_X1 U14164 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n13306) );
  NAND2_X1 U14165 ( .A1(n12900), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n11746) );
  NAND2_X1 U14166 ( .A1(n13169), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n11745) );
  OAI211_X1 U14167 ( .C1(n13306), .C2(n12903), .A(n11746), .B(n11745), .ZN(
        n11747) );
  INV_X1 U14168 ( .A(n11747), .ZN(n11748) );
  NAND2_X1 U14169 ( .A1(n11749), .A2(n11748), .ZN(n13906) );
  OAI22_X1 U14170 ( .A1(n13363), .A2(n14784), .B1(n11751), .B2(n13928), .ZN(
        n11845) );
  AOI21_X1 U14171 ( .B1(n11750), .B2(n15054), .A(n11845), .ZN(n14039) );
  OAI21_X1 U14172 ( .B1(n11754), .B2(n11753), .A(n13350), .ZN(n14040) );
  INV_X1 U14173 ( .A(n14040), .ZN(n11762) );
  INV_X1 U14174 ( .A(n14037), .ZN(n13349) );
  NAND2_X1 U14175 ( .A1(n11755), .A2(n14037), .ZN(n11756) );
  NAND2_X1 U14176 ( .A1(n11756), .A2(n11374), .ZN(n11757) );
  NOR2_X1 U14177 ( .A1(n13932), .A2(n11757), .ZN(n14036) );
  NAND2_X1 U14178 ( .A1(n14036), .A2(n15068), .ZN(n11760) );
  INV_X1 U14179 ( .A(n11842), .ZN(n11758) );
  AOI22_X1 U14180 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n15059), .B1(n11758), 
        .B2(n15058), .ZN(n11759) );
  OAI211_X1 U14181 ( .C1(n13349), .C2(n13959), .A(n11760), .B(n11759), .ZN(
        n11761) );
  AOI21_X1 U14182 ( .B1(n11762), .B2(n15069), .A(n11761), .ZN(n11763) );
  OAI21_X1 U14183 ( .B1(n14039), .B2(n15072), .A(n11763), .ZN(P2_U3248) );
  INV_X1 U14184 ( .A(n11764), .ZN(n11765) );
  AOI211_X1 U14185 ( .C1(n11769), .C2(n12566), .A(n15359), .B(n11765), .ZN(
        n11767) );
  OR2_X1 U14186 ( .A1(n11767), .A2(n11766), .ZN(n12647) );
  INV_X1 U14187 ( .A(n12647), .ZN(n11775) );
  OAI21_X1 U14188 ( .B1(n11770), .B2(n11769), .A(n11768), .ZN(n12648) );
  AOI22_X1 U14189 ( .A1(n12443), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n15379), 
        .B2(n11771), .ZN(n11772) );
  OAI21_X1 U14190 ( .B1(n12711), .B2(n12578), .A(n11772), .ZN(n11773) );
  AOI21_X1 U14191 ( .B1(n12648), .B2(n12581), .A(n11773), .ZN(n11774) );
  OAI21_X1 U14192 ( .B1(n11775), .B2(n12443), .A(n11774), .ZN(P3_U3219) );
  AND2_X1 U14193 ( .A1(n13263), .A2(n6611), .ZN(n11777) );
  XNOR2_X1 U14194 ( .A(n14042), .B(n12895), .ZN(n11776) );
  NOR2_X1 U14195 ( .A1(n11776), .A2(n11777), .ZN(n11836) );
  AOI21_X1 U14196 ( .B1(n11777), .B2(n11776), .A(n11836), .ZN(n11782) );
  INV_X1 U14197 ( .A(n11778), .ZN(n11779) );
  NAND2_X1 U14198 ( .A1(n11780), .A2(n11779), .ZN(n11781) );
  OAI21_X1 U14199 ( .B1(n11782), .B2(n11781), .A(n11838), .ZN(n11783) );
  NAND2_X1 U14200 ( .A1(n11783), .A2(n14793), .ZN(n11788) );
  AND2_X1 U14201 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n15042) );
  INV_X1 U14202 ( .A(n13262), .ZN(n13927) );
  OAI22_X1 U14203 ( .A1(n14785), .A2(n12963), .B1(n12962), .B2(n13927), .ZN(
        n11784) );
  AOI211_X1 U14204 ( .C1(n11786), .C2(n11785), .A(n15042), .B(n11784), .ZN(
        n11787) );
  OAI211_X1 U14205 ( .C1(n7079), .C2(n11848), .A(n11788), .B(n11787), .ZN(
        P2_U3198) );
  NAND2_X1 U14206 ( .A1(n12856), .A2(n11849), .ZN(n11790) );
  OAI211_X1 U14207 ( .C1(n11987), .C2(n11791), .A(n11790), .B(n11789), .ZN(
        P2_U3300) );
  INV_X1 U14208 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n13541) );
  AOI21_X1 U14209 ( .B1(n11793), .B2(n14775), .A(n11792), .ZN(n11795) );
  MUX2_X1 U14210 ( .A(n13541), .B(n11795), .S(n15436), .Z(n11794) );
  OAI21_X1 U14211 ( .B1(n12651), .B2(n11798), .A(n11794), .ZN(P3_U3472) );
  INV_X1 U14212 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n11796) );
  MUX2_X1 U14213 ( .A(n11796), .B(n11795), .S(n12707), .Z(n11797) );
  OAI21_X1 U14214 ( .B1(n12712), .B2(n11798), .A(n11797), .ZN(P3_U3429) );
  NAND2_X1 U14215 ( .A1(n11799), .A2(n12234), .ZN(n11801) );
  AND2_X1 U14216 ( .A1(n11801), .A2(n11800), .ZN(n12367) );
  NAND2_X1 U14217 ( .A1(n11802), .A2(n12367), .ZN(n11803) );
  XOR2_X1 U14218 ( .A(n11806), .B(n11803), .Z(n11804) );
  AOI22_X1 U14219 ( .A1(n15366), .A2(n12372), .B1(n12234), .B2(n12406), .ZN(
        n11858) );
  OAI21_X1 U14220 ( .B1(n11804), .B2(n15359), .A(n11858), .ZN(n12640) );
  INV_X1 U14221 ( .A(n12640), .ZN(n11811) );
  OAI21_X1 U14222 ( .B1(n11807), .B2(n11806), .A(n11805), .ZN(n12641) );
  INV_X1 U14223 ( .A(n12365), .ZN(n12702) );
  AOI22_X1 U14224 ( .A1(n12443), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15379), 
        .B2(n11861), .ZN(n11808) );
  OAI21_X1 U14225 ( .B1(n12702), .B2(n12578), .A(n11808), .ZN(n11809) );
  AOI21_X1 U14226 ( .B1(n12641), .B2(n12581), .A(n11809), .ZN(n11810) );
  OAI21_X1 U14227 ( .B1(n11811), .B2(n12443), .A(n11810), .ZN(P3_U3217) );
  INV_X1 U14228 ( .A(n11812), .ZN(n11813) );
  AOI21_X1 U14229 ( .B1(n11821), .B2(n11814), .A(n11813), .ZN(n14637) );
  OR2_X1 U14230 ( .A1(n11606), .A2(n11815), .ZN(n11818) );
  AND2_X1 U14231 ( .A1(n11818), .A2(n11816), .ZN(n11820) );
  NAND2_X1 U14232 ( .A1(n11818), .A2(n11817), .ZN(n11819) );
  OAI211_X1 U14233 ( .C1(n11821), .C2(n11820), .A(n11819), .B(n14701), .ZN(
        n11823) );
  AOI22_X1 U14234 ( .A1(n14538), .A2(n14540), .B1(n14539), .B2(n14239), .ZN(
        n11822) );
  OAI21_X1 U14235 ( .B1(n14222), .B2(n14498), .A(n14636), .ZN(n11824) );
  NAND2_X1 U14236 ( .A1(n11824), .A2(n14531), .ZN(n11831) );
  INV_X1 U14237 ( .A(n11825), .ZN(n11827) );
  INV_X1 U14238 ( .A(n11882), .ZN(n11826) );
  AOI211_X1 U14239 ( .C1(n14634), .C2(n11827), .A(n14503), .B(n11826), .ZN(
        n14633) );
  OAI22_X1 U14240 ( .A1(n14231), .A2(n14506), .B1(n14531), .B2(n11828), .ZN(
        n11829) );
  AOI21_X1 U14241 ( .B1(n14633), .B2(n14716), .A(n11829), .ZN(n11830) );
  OAI211_X1 U14242 ( .C1(n14637), .C2(n14511), .A(n11831), .B(n11830), .ZN(
        P1_U3278) );
  INV_X1 U14243 ( .A(n12856), .ZN(n11832) );
  OAI222_X1 U14244 ( .A1(n12137), .A2(n11833), .B1(P1_U3086), .B2(n6684), .C1(
        n14668), .C2(n11832), .ZN(P1_U3328) );
  AND2_X1 U14245 ( .A1(n13262), .A2(n6611), .ZN(n11835) );
  XNOR2_X1 U14246 ( .A(n14037), .B(n12895), .ZN(n11834) );
  NOR2_X1 U14247 ( .A1(n11834), .A2(n11835), .ZN(n11864) );
  AOI21_X1 U14248 ( .B1(n11835), .B2(n11834), .A(n11864), .ZN(n11840) );
  INV_X1 U14249 ( .A(n11836), .ZN(n11837) );
  OAI21_X1 U14250 ( .B1(n11840), .B2(n11839), .A(n11866), .ZN(n11841) );
  NAND2_X1 U14251 ( .A1(n11841), .A2(n14793), .ZN(n11847) );
  NOR2_X1 U14252 ( .A1(n14799), .A2(n11842), .ZN(n11844) );
  AOI211_X1 U14253 ( .C1(n11845), .C2(n14795), .A(n11844), .B(n11843), .ZN(
        n11846) );
  OAI211_X1 U14254 ( .C1(n13349), .C2(n11848), .A(n11847), .B(n11846), .ZN(
        P2_U3200) );
  NAND2_X1 U14255 ( .A1(n12891), .A2(n11849), .ZN(n11851) );
  OAI211_X1 U14256 ( .C1(n11987), .C2(n13634), .A(n11851), .B(n11850), .ZN(
        P2_U3299) );
  INV_X1 U14257 ( .A(n11853), .ZN(n11855) );
  NAND2_X1 U14258 ( .A1(n11855), .A2(n11854), .ZN(n11856) );
  XNOR2_X1 U14259 ( .A(n11852), .B(n11856), .ZN(n11863) );
  OAI22_X1 U14260 ( .A1(n11858), .A2(n15203), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11857), .ZN(n11860) );
  NOR2_X1 U14261 ( .A1(n12702), .A2(n12230), .ZN(n11859) );
  AOI211_X1 U14262 ( .C1(n11861), .C2(n12227), .A(n11860), .B(n11859), .ZN(
        n11862) );
  OAI21_X1 U14263 ( .B1(n11863), .B2(n15207), .A(n11862), .ZN(P3_U3166) );
  INV_X1 U14264 ( .A(n11864), .ZN(n11865) );
  NAND2_X1 U14265 ( .A1(n13906), .A2(n6611), .ZN(n12728) );
  NAND2_X1 U14266 ( .A1(n11867), .A2(n10117), .ZN(n11869) );
  AOI22_X1 U14267 ( .A1(n12892), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n12733), 
        .B2(n13318), .ZN(n11868) );
  XNOR2_X1 U14268 ( .A(n14030), .B(n12895), .ZN(n12727) );
  XOR2_X1 U14269 ( .A(n12728), .B(n12727), .Z(n12730) );
  XNOR2_X1 U14270 ( .A(n12731), .B(n12730), .ZN(n11881) );
  NAND2_X1 U14271 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13308)
         );
  OAI21_X1 U14272 ( .B1(n14799), .B2(n13933), .A(n13308), .ZN(n11879) );
  INV_X1 U14273 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n11870) );
  NAND2_X1 U14274 ( .A1(n11871), .A2(n11870), .ZN(n11872) );
  NAND2_X1 U14275 ( .A1(n12744), .A2(n11872), .ZN(n13912) );
  INV_X1 U14276 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n11875) );
  NAND2_X1 U14277 ( .A1(n13168), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n11874) );
  NAND2_X1 U14278 ( .A1(n13169), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n11873) );
  OAI211_X1 U14279 ( .C1(n13172), .C2(n11875), .A(n11874), .B(n11873), .ZN(
        n11876) );
  INV_X1 U14280 ( .A(n11876), .ZN(n11877) );
  OAI21_X1 U14281 ( .B1(n13912), .B2(n12901), .A(n11877), .ZN(n13261) );
  INV_X1 U14282 ( .A(n13261), .ZN(n13929) );
  OAI22_X1 U14283 ( .A1(n13929), .A2(n12962), .B1(n13927), .B2(n12963), .ZN(
        n11878) );
  AOI211_X1 U14284 ( .C1(n14030), .C2(n14796), .A(n11879), .B(n11878), .ZN(
        n11880) );
  OAI21_X1 U14285 ( .B1(n11881), .B2(n12967), .A(n11880), .ZN(P2_U3210) );
  AOI21_X1 U14286 ( .B1(n11882), .B2(n14153), .A(n14503), .ZN(n11884) );
  INV_X1 U14287 ( .A(n11883), .ZN(n14533) );
  NAND2_X1 U14288 ( .A1(n11884), .A2(n14533), .ZN(n14627) );
  OR2_X1 U14289 ( .A1(n11885), .A2(n14959), .ZN(n11889) );
  AOI22_X1 U14290 ( .A1(n11886), .A2(n14701), .B1(n14965), .B2(n11885), .ZN(
        n11888) );
  MUX2_X1 U14291 ( .A(n11889), .B(n11888), .S(n11887), .Z(n11894) );
  AOI22_X1 U14292 ( .A1(n14517), .A2(n14540), .B1(n14539), .B2(n14238), .ZN(
        n11890) );
  OAI21_X1 U14293 ( .B1(n11891), .B2(n14603), .A(n11890), .ZN(n11892) );
  INV_X1 U14294 ( .A(n11892), .ZN(n11893) );
  NAND2_X1 U14295 ( .A1(n11894), .A2(n11893), .ZN(n14630) );
  NAND2_X1 U14296 ( .A1(n14630), .A2(n14531), .ZN(n11898) );
  OAI22_X1 U14297 ( .A1(n14531), .A2(n11895), .B1(n14151), .B2(n14498), .ZN(
        n11896) );
  AOI21_X1 U14298 ( .B1(n14153), .B2(n14706), .A(n11896), .ZN(n11897) );
  OAI211_X1 U14299 ( .C1(n14627), .C2(n14529), .A(n11898), .B(n11897), .ZN(
        P1_U3277) );
  AOI22_X1 U14300 ( .A1(n14843), .A2(n12073), .B1(n12119), .B2(n14242), .ZN(
        n11907) );
  NAND2_X1 U14301 ( .A1(n14843), .A2(n12120), .ZN(n11903) );
  NAND2_X1 U14302 ( .A1(n14242), .A2(n12054), .ZN(n11902) );
  NAND2_X1 U14303 ( .A1(n11903), .A2(n11902), .ZN(n11904) );
  XNOR2_X1 U14304 ( .A(n11904), .B(n12121), .ZN(n11909) );
  XOR2_X1 U14305 ( .A(n11907), .B(n11909), .Z(n14849) );
  INV_X1 U14306 ( .A(n14849), .ZN(n11905) );
  INV_X1 U14307 ( .A(n11907), .ZN(n11908) );
  AOI22_X1 U14308 ( .A1(n14707), .A2(n12120), .B1(n12054), .B2(n14241), .ZN(
        n11911) );
  XNOR2_X1 U14309 ( .A(n11911), .B(n12121), .ZN(n11921) );
  NOR2_X1 U14310 ( .A1(n11912), .A2(n12062), .ZN(n11913) );
  AOI21_X1 U14311 ( .B1(n14707), .B2(n12054), .A(n11913), .ZN(n11922) );
  XNOR2_X1 U14312 ( .A(n11921), .B(n11922), .ZN(n11915) );
  AOI21_X1 U14313 ( .B1(n11914), .B2(n11915), .A(n14850), .ZN(n11917) );
  NAND2_X1 U14314 ( .A1(n11917), .A2(n11926), .ZN(n11920) );
  INV_X1 U14315 ( .A(n14855), .ZN(n14181) );
  AOI22_X1 U14316 ( .A1(n14539), .A2(n14242), .B1(n14240), .B2(n14540), .ZN(
        n14699) );
  OAI22_X1 U14317 ( .A1(n14181), .A2(n14699), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8559), .ZN(n11918) );
  AOI21_X1 U14318 ( .B1(n14704), .B2(n14228), .A(n11918), .ZN(n11919) );
  OAI211_X1 U14319 ( .C1(n14721), .C2(n14896), .A(n11920), .B(n11919), .ZN(
        P1_U3224) );
  INV_X1 U14320 ( .A(n11921), .ZN(n11924) );
  INV_X1 U14321 ( .A(n11922), .ZN(n11923) );
  NOR2_X1 U14322 ( .A1(n14094), .A2(n12062), .ZN(n11927) );
  AOI21_X1 U14323 ( .B1(n11928), .B2(n12054), .A(n11927), .ZN(n12009) );
  AOI22_X1 U14324 ( .A1(n11928), .A2(n12120), .B1(n12054), .B2(n14240), .ZN(
        n11929) );
  XNOR2_X1 U14325 ( .A(n11929), .B(n12121), .ZN(n12008) );
  XOR2_X1 U14326 ( .A(n12009), .B(n12008), .Z(n11930) );
  OAI211_X1 U14327 ( .C1(n11931), .C2(n11930), .A(n12013), .B(n14904), .ZN(
        n11937) );
  OAI21_X1 U14328 ( .B1(n14181), .B2(n11933), .A(n11932), .ZN(n11934) );
  AOI21_X1 U14329 ( .B1(n11935), .B2(n14228), .A(n11934), .ZN(n11936) );
  OAI211_X1 U14330 ( .C1(n14860), .C2(n14896), .A(n11937), .B(n11936), .ZN(
        P1_U3234) );
  INV_X1 U14331 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n11938) );
  OAI222_X1 U14332 ( .A1(n6618), .A2(n13165), .B1(P2_U3088), .B2(n11939), .C1(
        n11938), .C2(n11987), .ZN(P2_U3297) );
  XNOR2_X1 U14333 ( .A(n11941), .B(n11940), .ZN(n12766) );
  INV_X1 U14334 ( .A(n12766), .ZN(n11942) );
  OAI222_X1 U14335 ( .A1(n11987), .A2(n11943), .B1(n6618), .B2(n11942), .C1(
        n10168), .C2(P2_U3088), .ZN(P2_U3305) );
  INV_X1 U14336 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n11944) );
  NOR2_X1 U14337 ( .A1(n12707), .A2(n11944), .ZN(n11945) );
  AOI21_X1 U14338 ( .B1(n12707), .B2(n11948), .A(n11945), .ZN(n11946) );
  OAI21_X1 U14339 ( .B1(n11950), .B2(n12712), .A(n11946), .ZN(P3_U3390) );
  NOR2_X1 U14340 ( .A1(n15436), .A2(n9978), .ZN(n11947) );
  AOI21_X1 U14341 ( .B1(n15436), .B2(n11948), .A(n11947), .ZN(n11949) );
  OAI21_X1 U14342 ( .B1(n11950), .B2(n12651), .A(n11949), .ZN(P3_U3459) );
  INV_X1 U14343 ( .A(n11951), .ZN(n11954) );
  OAI222_X1 U14344 ( .A1(n11991), .A2(n11954), .B1(n11995), .B2(n11953), .C1(
        P3_U3151), .C2(n11952), .ZN(P3_U3274) );
  AOI21_X1 U14345 ( .B1(n11957), .B2(n11956), .A(n11955), .ZN(n11963) );
  AOI22_X1 U14346 ( .A1(n14194), .A2(n14246), .B1(n14193), .B2(n14244), .ZN(
        n11959) );
  OAI211_X1 U14347 ( .C1(n11960), .C2(n14909), .A(n11959), .B(n11958), .ZN(
        n11961) );
  AOI21_X1 U14348 ( .B1(n14215), .B2(n14956), .A(n11961), .ZN(n11962) );
  OAI21_X1 U14349 ( .B1(n11963), .B2(n14850), .A(n11962), .ZN(P1_U3221) );
  NAND2_X1 U14350 ( .A1(n11967), .A2(n11966), .ZN(n11969) );
  NAND2_X1 U14351 ( .A1(n11998), .A2(n14362), .ZN(n11968) );
  NAND2_X1 U14352 ( .A1(n11969), .A2(n11968), .ZN(n11971) );
  XNOR2_X1 U14353 ( .A(n11971), .B(n11970), .ZN(n14562) );
  NOR2_X1 U14354 ( .A1(n14705), .A2(n14603), .ZN(n14390) );
  NAND2_X1 U14355 ( .A1(n14562), .A2(n14390), .ZN(n11985) );
  AOI21_X1 U14356 ( .B1(n11972), .B2(n14561), .A(n14503), .ZN(n11973) );
  NAND2_X1 U14357 ( .A1(n14561), .A2(n14706), .ZN(n11982) );
  NAND2_X1 U14358 ( .A1(n14362), .A2(n14539), .ZN(n11977) );
  NAND2_X1 U14359 ( .A1(n11974), .A2(P1_B_REG_SCAN_IN), .ZN(n11975) );
  AND2_X1 U14360 ( .A1(n14540), .A2(n11975), .ZN(n14340) );
  NAND2_X1 U14361 ( .A1(n14232), .A2(n14340), .ZN(n11976) );
  NAND2_X1 U14362 ( .A1(n11977), .A2(n11976), .ZN(n14560) );
  INV_X1 U14363 ( .A(n14560), .ZN(n11979) );
  OAI22_X1 U14364 ( .A1(n14526), .A2(n11979), .B1(n11978), .B2(n14498), .ZN(
        n11980) );
  INV_X1 U14365 ( .A(n11980), .ZN(n11981) );
  OAI211_X1 U14366 ( .C1(n14531), .C2(n13675), .A(n11982), .B(n11981), .ZN(
        n11983) );
  AOI21_X1 U14367 ( .B1(n14559), .B2(n14716), .A(n11983), .ZN(n11984) );
  OAI211_X1 U14368 ( .C1(n14564), .C2(n14511), .A(n11985), .B(n11984), .ZN(
        P1_U3356) );
  INV_X1 U14369 ( .A(n13157), .ZN(n14672) );
  OAI222_X1 U14370 ( .A1(n6618), .A2(n14672), .B1(P2_U3088), .B2(n11989), .C1(
        n11988), .C2(n11987), .ZN(P2_U3298) );
  OAI222_X1 U14371 ( .A1(n11995), .A2(n11993), .B1(P3_U3151), .B2(n7624), .C1(
        n11991), .C2(n11990), .ZN(P3_U3266) );
  OAI222_X1 U14372 ( .A1(n11991), .A2(n11996), .B1(n11995), .B2(n11994), .C1(
        P3_U3151), .C2(n6687), .ZN(P3_U3276) );
  AOI22_X1 U14373 ( .A1(n14526), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n12126), 
        .B2(n14703), .ZN(n11997) );
  OAI21_X1 U14374 ( .B1(n11998), .B2(n14506), .A(n11997), .ZN(n12001) );
  NOR2_X1 U14375 ( .A1(n11999), .A2(n14511), .ZN(n12000) );
  OAI21_X1 U14376 ( .B1(n12004), .B2(n14705), .A(n12003), .ZN(P1_U3265) );
  INV_X1 U14377 ( .A(n12891), .ZN(n12006) );
  OAI222_X1 U14378 ( .A1(n12137), .A2(n12007), .B1(n14668), .B2(n12006), .C1(
        n12005), .C2(P1_U3086), .ZN(P1_U3327) );
  INV_X1 U14379 ( .A(n12009), .ZN(n12010) );
  AOI22_X1 U14380 ( .A1(n14639), .A2(n12120), .B1(n12073), .B2(n14239), .ZN(
        n12014) );
  XNOR2_X1 U14381 ( .A(n12014), .B(n12121), .ZN(n12015) );
  AOI22_X1 U14382 ( .A1(n14639), .A2(n12073), .B1(n12119), .B2(n14239), .ZN(
        n12016) );
  XNOR2_X1 U14383 ( .A(n12015), .B(n12016), .ZN(n14093) );
  NAND2_X1 U14384 ( .A1(n14634), .A2(n12120), .ZN(n12019) );
  NAND2_X1 U14385 ( .A1(n14238), .A2(n12054), .ZN(n12018) );
  NAND2_X1 U14386 ( .A1(n12019), .A2(n12018), .ZN(n12020) );
  XNOR2_X1 U14387 ( .A(n12020), .B(n12121), .ZN(n12021) );
  AOI22_X1 U14388 ( .A1(n14634), .A2(n12073), .B1(n12119), .B2(n14238), .ZN(
        n14220) );
  INV_X1 U14389 ( .A(n12021), .ZN(n12022) );
  AOI22_X1 U14390 ( .A1(n14153), .A2(n12073), .B1(n12119), .B2(n14538), .ZN(
        n12028) );
  NAND2_X1 U14391 ( .A1(n14153), .A2(n12120), .ZN(n12026) );
  NAND2_X1 U14392 ( .A1(n14538), .A2(n12073), .ZN(n12025) );
  NAND2_X1 U14393 ( .A1(n12026), .A2(n12025), .ZN(n12027) );
  XNOR2_X1 U14394 ( .A(n12027), .B(n12121), .ZN(n12030) );
  XOR2_X1 U14395 ( .A(n12028), .B(n12030), .Z(n14148) );
  INV_X1 U14396 ( .A(n12028), .ZN(n12029) );
  NAND2_X1 U14397 ( .A1(n14550), .A2(n12120), .ZN(n12033) );
  NAND2_X1 U14398 ( .A1(n14517), .A2(n12073), .ZN(n12032) );
  NAND2_X1 U14399 ( .A1(n12033), .A2(n12032), .ZN(n12034) );
  XNOR2_X1 U14400 ( .A(n12034), .B(n12121), .ZN(n12035) );
  AOI22_X1 U14401 ( .A1(n14550), .A2(n12073), .B1(n12119), .B2(n14517), .ZN(
        n12036) );
  XNOR2_X1 U14402 ( .A(n12035), .B(n12036), .ZN(n14157) );
  INV_X1 U14403 ( .A(n12035), .ZN(n12037) );
  NAND2_X1 U14404 ( .A1(n12037), .A2(n12036), .ZN(n12038) );
  NAND2_X1 U14405 ( .A1(n14620), .A2(n12120), .ZN(n12040) );
  NAND2_X1 U14406 ( .A1(n14541), .A2(n12073), .ZN(n12039) );
  NAND2_X1 U14407 ( .A1(n12040), .A2(n12039), .ZN(n12041) );
  XNOR2_X1 U14408 ( .A(n12041), .B(n12121), .ZN(n12042) );
  AOI22_X1 U14409 ( .A1(n14620), .A2(n12073), .B1(n12119), .B2(n14541), .ZN(
        n12043) );
  XNOR2_X1 U14410 ( .A(n12042), .B(n12043), .ZN(n14200) );
  INV_X1 U14411 ( .A(n12042), .ZN(n12044) );
  NAND2_X1 U14412 ( .A1(n12044), .A2(n12043), .ZN(n12045) );
  AND2_X1 U14413 ( .A1(n14518), .A2(n12119), .ZN(n12046) );
  AOI21_X1 U14414 ( .B1(n14616), .B2(n12054), .A(n12046), .ZN(n12050) );
  NAND2_X1 U14415 ( .A1(n14616), .A2(n12120), .ZN(n12048) );
  NAND2_X1 U14416 ( .A1(n14518), .A2(n12073), .ZN(n12047) );
  NAND2_X1 U14417 ( .A1(n12048), .A2(n12047), .ZN(n12049) );
  XNOR2_X1 U14418 ( .A(n12049), .B(n12121), .ZN(n12052) );
  XOR2_X1 U14419 ( .A(n12050), .B(n12052), .Z(n14117) );
  INV_X1 U14420 ( .A(n12050), .ZN(n12051) );
  AND2_X1 U14421 ( .A1(n14496), .A2(n12119), .ZN(n12053) );
  AOI21_X1 U14422 ( .B1(n14609), .B2(n12054), .A(n12053), .ZN(n12057) );
  AOI22_X1 U14423 ( .A1(n14609), .A2(n12120), .B1(n12054), .B2(n14496), .ZN(
        n12055) );
  XNOR2_X1 U14424 ( .A(n12055), .B(n12121), .ZN(n12056) );
  XOR2_X1 U14425 ( .A(n12057), .B(n12056), .Z(n14175) );
  INV_X1 U14426 ( .A(n12056), .ZN(n12059) );
  INV_X1 U14427 ( .A(n12057), .ZN(n12058) );
  NAND2_X1 U14428 ( .A1(n12059), .A2(n12058), .ZN(n12060) );
  OAI22_X1 U14429 ( .A1(n14460), .A2(n10243), .B1(n14439), .B2(n12063), .ZN(
        n12061) );
  XNOR2_X1 U14430 ( .A(n12061), .B(n12121), .ZN(n12074) );
  OAI22_X1 U14431 ( .A1(n14460), .A2(n12063), .B1(n14439), .B2(n12062), .ZN(
        n12075) );
  XNOR2_X1 U14432 ( .A(n12074), .B(n12075), .ZN(n14131) );
  OR2_X1 U14433 ( .A1(n14445), .A2(n12063), .ZN(n12065) );
  NAND2_X1 U14434 ( .A1(n14236), .A2(n12119), .ZN(n12064) );
  NAND2_X1 U14435 ( .A1(n12065), .A2(n12064), .ZN(n12080) );
  OAI22_X1 U14436 ( .A1(n14445), .A2(n10243), .B1(n14467), .B2(n12063), .ZN(
        n12066) );
  XNOR2_X1 U14437 ( .A(n12066), .B(n12121), .ZN(n12079) );
  XOR2_X1 U14438 ( .A(n12080), .B(n12079), .Z(n14191) );
  INV_X1 U14439 ( .A(n14191), .ZN(n12078) );
  OR2_X1 U14440 ( .A1(n14131), .A2(n12078), .ZN(n14103) );
  NAND2_X1 U14441 ( .A1(n14423), .A2(n12120), .ZN(n12068) );
  NAND2_X1 U14442 ( .A1(n14440), .A2(n12054), .ZN(n12067) );
  NAND2_X1 U14443 ( .A1(n12068), .A2(n12067), .ZN(n12069) );
  XNOR2_X1 U14444 ( .A(n12069), .B(n12121), .ZN(n12085) );
  AOI22_X1 U14445 ( .A1(n14423), .A2(n12073), .B1(n12119), .B2(n14440), .ZN(
        n12086) );
  XNOR2_X1 U14446 ( .A(n12085), .B(n12086), .ZN(n14106) );
  INV_X1 U14447 ( .A(n14106), .ZN(n12084) );
  NAND2_X1 U14448 ( .A1(n14585), .A2(n12120), .ZN(n12071) );
  NAND2_X1 U14449 ( .A1(n14235), .A2(n12112), .ZN(n12070) );
  NAND2_X1 U14450 ( .A1(n12071), .A2(n12070), .ZN(n12072) );
  XNOR2_X1 U14451 ( .A(n12072), .B(n12121), .ZN(n12091) );
  AOI22_X1 U14452 ( .A1(n14585), .A2(n12073), .B1(n12119), .B2(n14235), .ZN(
        n12092) );
  XNOR2_X1 U14453 ( .A(n12091), .B(n12092), .ZN(n14166) );
  INV_X1 U14454 ( .A(n14166), .ZN(n12090) );
  INV_X1 U14455 ( .A(n12074), .ZN(n12077) );
  INV_X1 U14456 ( .A(n12075), .ZN(n12076) );
  NAND2_X1 U14457 ( .A1(n12077), .A2(n12076), .ZN(n14185) );
  INV_X1 U14458 ( .A(n12079), .ZN(n12082) );
  INV_X1 U14459 ( .A(n12080), .ZN(n12081) );
  NAND2_X1 U14460 ( .A1(n12082), .A2(n12081), .ZN(n12083) );
  INV_X1 U14461 ( .A(n12085), .ZN(n12087) );
  NAND2_X1 U14462 ( .A1(n12087), .A2(n12086), .ZN(n12088) );
  INV_X1 U14463 ( .A(n12091), .ZN(n12093) );
  NAND2_X1 U14464 ( .A1(n12093), .A2(n12092), .ZN(n12094) );
  NAND2_X1 U14465 ( .A1(n14578), .A2(n12120), .ZN(n12098) );
  NAND2_X1 U14466 ( .A1(n14404), .A2(n12112), .ZN(n12097) );
  NAND2_X1 U14467 ( .A1(n12098), .A2(n12097), .ZN(n12099) );
  XNOR2_X1 U14468 ( .A(n12099), .B(n12121), .ZN(n12100) );
  AOI22_X1 U14469 ( .A1(n14578), .A2(n12073), .B1(n12119), .B2(n14404), .ZN(
        n12101) );
  XNOR2_X1 U14470 ( .A(n12100), .B(n12101), .ZN(n14140) );
  INV_X1 U14471 ( .A(n12100), .ZN(n12102) );
  NAND2_X1 U14472 ( .A1(n12102), .A2(n12101), .ZN(n12103) );
  NAND2_X1 U14473 ( .A1(n12104), .A2(n12103), .ZN(n14208) );
  NAND2_X1 U14474 ( .A1(n14572), .A2(n12120), .ZN(n12106) );
  NAND2_X1 U14475 ( .A1(n14361), .A2(n12112), .ZN(n12105) );
  NAND2_X1 U14476 ( .A1(n12106), .A2(n12105), .ZN(n12107) );
  XNOR2_X1 U14477 ( .A(n12107), .B(n12121), .ZN(n12108) );
  AOI22_X1 U14478 ( .A1(n14572), .A2(n12073), .B1(n12119), .B2(n14361), .ZN(
        n12109) );
  XNOR2_X1 U14479 ( .A(n12108), .B(n12109), .ZN(n14209) );
  INV_X1 U14480 ( .A(n12108), .ZN(n12110) );
  NAND2_X1 U14481 ( .A1(n12110), .A2(n12109), .ZN(n12111) );
  NAND2_X1 U14482 ( .A1(n14567), .A2(n12120), .ZN(n12114) );
  NAND2_X1 U14483 ( .A1(n14234), .A2(n12112), .ZN(n12113) );
  NAND2_X1 U14484 ( .A1(n12114), .A2(n12113), .ZN(n12115) );
  XNOR2_X1 U14485 ( .A(n12115), .B(n12121), .ZN(n12116) );
  AOI22_X1 U14486 ( .A1(n14567), .A2(n12054), .B1(n12119), .B2(n14234), .ZN(
        n12117) );
  XNOR2_X1 U14487 ( .A(n12116), .B(n12117), .ZN(n14083) );
  INV_X1 U14488 ( .A(n12116), .ZN(n12118) );
  AOI22_X1 U14489 ( .A1(n12132), .A2(n12073), .B1(n12119), .B2(n14362), .ZN(
        n12124) );
  AOI22_X1 U14490 ( .A1(n12132), .A2(n12120), .B1(n12073), .B2(n14362), .ZN(
        n12122) );
  XNOR2_X1 U14491 ( .A(n12122), .B(n12121), .ZN(n12123) );
  XOR2_X1 U14492 ( .A(n12124), .B(n12123), .Z(n12125) );
  INV_X1 U14493 ( .A(n12126), .ZN(n12128) );
  OAI22_X1 U14494 ( .A1(n14909), .A2(n12128), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12127), .ZN(n12131) );
  OAI22_X1 U14495 ( .A1(n12129), .A2(n14899), .B1(n14900), .B2(n14211), .ZN(
        n12130) );
  AOI211_X1 U14496 ( .C1(n12132), .C2(n14215), .A(n12131), .B(n12130), .ZN(
        n12133) );
  OAI21_X1 U14497 ( .B1(n12134), .B2(n14850), .A(n12133), .ZN(P1_U3220) );
  OAI222_X1 U14498 ( .A1(n12137), .A2(n12136), .B1(n14668), .B2(n12135), .C1(
        n8875), .C2(P1_U3086), .ZN(P1_U3331) );
  INV_X1 U14499 ( .A(n12183), .ZN(n12138) );
  AOI21_X1 U14500 ( .B1(n12389), .B2(n12139), .A(n12138), .ZN(n12144) );
  OAI22_X1 U14501 ( .A1(n12224), .A2(n12489), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13725), .ZN(n12141) );
  NOR2_X1 U14502 ( .A1(n12488), .A2(n12222), .ZN(n12140) );
  AOI211_X1 U14503 ( .C1(n12493), .C2(n12227), .A(n12141), .B(n12140), .ZN(
        n12143) );
  NAND2_X1 U14504 ( .A1(n12492), .A2(n15213), .ZN(n12142) );
  OAI211_X1 U14505 ( .C1(n12144), .C2(n15207), .A(n12143), .B(n12142), .ZN(
        P3_U3156) );
  XOR2_X1 U14506 ( .A(n6850), .B(n12145), .Z(n12147) );
  NAND2_X1 U14507 ( .A1(n12147), .A2(n15193), .ZN(n12153) );
  INV_X1 U14508 ( .A(n12538), .ZN(n12148) );
  NOR2_X1 U14509 ( .A1(n15215), .A2(n12148), .ZN(n12151) );
  INV_X1 U14510 ( .A(n12534), .ZN(n12571) );
  NAND2_X1 U14511 ( .A1(n12571), .A2(n12212), .ZN(n12149) );
  NAND2_X1 U14512 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12339)
         );
  OAI211_X1 U14513 ( .C1(n12535), .C2(n12224), .A(n12149), .B(n12339), .ZN(
        n12150) );
  NOR2_X1 U14514 ( .A1(n12151), .A2(n12150), .ZN(n12152) );
  OAI211_X1 U14515 ( .C1(n12230), .C2(n12694), .A(n12153), .B(n12152), .ZN(
        P3_U3159) );
  AOI21_X1 U14516 ( .B1(n12155), .B2(n12154), .A(n6796), .ZN(n12163) );
  INV_X1 U14517 ( .A(n12515), .ZN(n12160) );
  NAND2_X1 U14518 ( .A1(n12386), .A2(n15366), .ZN(n12157) );
  NAND2_X1 U14519 ( .A1(n12381), .A2(n12406), .ZN(n12156) );
  NAND2_X1 U14520 ( .A1(n12157), .A2(n12156), .ZN(n12511) );
  AOI22_X1 U14521 ( .A1(n12511), .A2(n12158), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12159) );
  OAI21_X1 U14522 ( .B1(n12160), .B2(n15215), .A(n12159), .ZN(n12161) );
  AOI21_X1 U14523 ( .B1(n12683), .B2(n15213), .A(n12161), .ZN(n12162) );
  OAI21_X1 U14524 ( .B1(n12163), .B2(n15207), .A(n12162), .ZN(P3_U3163) );
  INV_X1 U14525 ( .A(n12396), .ZN(n12668) );
  INV_X1 U14526 ( .A(n12164), .ZN(n12168) );
  NOR3_X1 U14527 ( .A1(n12185), .A2(n12166), .A3(n12165), .ZN(n12167) );
  OAI21_X1 U14528 ( .B1(n12168), .B2(n12167), .A(n15193), .ZN(n12173) );
  AOI22_X1 U14529 ( .A1(n12169), .A2(n12464), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12170) );
  OAI21_X1 U14530 ( .B1(n12489), .B2(n12222), .A(n12170), .ZN(n12171) );
  AOI21_X1 U14531 ( .B1(n12469), .B2(n12227), .A(n12171), .ZN(n12172) );
  OAI211_X1 U14532 ( .C1(n12668), .C2(n12230), .A(n12173), .B(n12172), .ZN(
        P3_U3165) );
  XNOR2_X1 U14533 ( .A(n12175), .B(n12174), .ZN(n12180) );
  NAND2_X1 U14534 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n14765)
         );
  NAND2_X1 U14535 ( .A1(n12212), .A2(n12570), .ZN(n12176) );
  OAI211_X1 U14536 ( .C1(n12534), .C2(n12224), .A(n14765), .B(n12176), .ZN(
        n12177) );
  AOI21_X1 U14537 ( .B1(n12227), .B2(n12576), .A(n12177), .ZN(n12179) );
  NAND2_X1 U14538 ( .A1(n12636), .A2(n15213), .ZN(n12178) );
  OAI211_X1 U14539 ( .C1(n12180), .C2(n15207), .A(n12179), .B(n12178), .ZN(
        P3_U3168) );
  INV_X1 U14540 ( .A(n12392), .ZN(n12672) );
  AND3_X1 U14541 ( .A1(n12183), .A2(n12182), .A3(n12181), .ZN(n12184) );
  OAI21_X1 U14542 ( .B1(n12185), .B2(n12184), .A(n15193), .ZN(n12189) );
  AOI22_X1 U14543 ( .A1(n12406), .A2(n12389), .B1(n12395), .B2(n15366), .ZN(
        n12476) );
  INV_X1 U14544 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n12186) );
  OAI22_X1 U14545 ( .A1(n12476), .A2(n15203), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12186), .ZN(n12187) );
  AOI21_X1 U14546 ( .B1(n12481), .B2(n12227), .A(n12187), .ZN(n12188) );
  OAI211_X1 U14547 ( .C1(n12672), .C2(n12230), .A(n12189), .B(n12188), .ZN(
        P3_U3169) );
  XNOR2_X1 U14548 ( .A(n12191), .B(n12190), .ZN(n12198) );
  OR2_X1 U14549 ( .A1(n12202), .A2(n15351), .ZN(n12193) );
  NAND2_X1 U14550 ( .A1(n12233), .A2(n12406), .ZN(n12192) );
  AND2_X1 U14551 ( .A1(n12193), .A2(n12192), .ZN(n12523) );
  OAI22_X1 U14552 ( .A1(n12523), .A2(n15203), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12194), .ZN(n12196) );
  INV_X1 U14553 ( .A(n12626), .ZN(n12690) );
  NOR2_X1 U14554 ( .A1(n12690), .A2(n12230), .ZN(n12195) );
  AOI211_X1 U14555 ( .C1(n12527), .C2(n12227), .A(n12196), .B(n12195), .ZN(
        n12197) );
  OAI21_X1 U14556 ( .B1(n12198), .B2(n15207), .A(n12197), .ZN(P3_U3173) );
  INV_X1 U14557 ( .A(n12387), .ZN(n12680) );
  OAI21_X1 U14558 ( .B1(n12488), .B2(n12200), .A(n12199), .ZN(n12201) );
  NAND2_X1 U14559 ( .A1(n12201), .A2(n15193), .ZN(n12209) );
  OR2_X1 U14560 ( .A1(n12202), .A2(n15353), .ZN(n12205) );
  OR2_X1 U14561 ( .A1(n12203), .A2(n15351), .ZN(n12204) );
  AND2_X1 U14562 ( .A1(n12205), .A2(n12204), .ZN(n12499) );
  INV_X1 U14563 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n12206) );
  OAI22_X1 U14564 ( .A1(n12499), .A2(n15203), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12206), .ZN(n12207) );
  AOI21_X1 U14565 ( .B1(n12504), .B2(n12227), .A(n12207), .ZN(n12208) );
  OAI211_X1 U14566 ( .C1(n12680), .C2(n12230), .A(n12209), .B(n12208), .ZN(
        P3_U3175) );
  XNOR2_X1 U14567 ( .A(n12211), .B(n12210), .ZN(n12217) );
  NAND2_X1 U14568 ( .A1(n12212), .A2(n12372), .ZN(n12213) );
  NAND2_X1 U14569 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12314)
         );
  OAI211_X1 U14570 ( .C1(n12553), .C2(n12224), .A(n12213), .B(n12314), .ZN(
        n12215) );
  INV_X1 U14571 ( .A(n12560), .ZN(n12697) );
  NOR2_X1 U14572 ( .A1(n12697), .A2(n12230), .ZN(n12214) );
  AOI211_X1 U14573 ( .C1(n12554), .C2(n12227), .A(n12215), .B(n12214), .ZN(
        n12216) );
  OAI21_X1 U14574 ( .B1(n12217), .B2(n15207), .A(n12216), .ZN(P3_U3178) );
  INV_X1 U14575 ( .A(n12398), .ZN(n12664) );
  OAI21_X1 U14576 ( .B1(n12220), .B2(n12219), .A(n12218), .ZN(n12221) );
  NAND2_X1 U14577 ( .A1(n12221), .A2(n15193), .ZN(n12229) );
  NOR2_X1 U14578 ( .A1(n12222), .A2(n12448), .ZN(n12226) );
  OAI22_X1 U14579 ( .A1(n12224), .A2(n12449), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12223), .ZN(n12225) );
  AOI211_X1 U14580 ( .C1(n12227), .C2(n12454), .A(n12226), .B(n12225), .ZN(
        n12228) );
  OAI211_X1 U14581 ( .C1(n12664), .C2(n12230), .A(n12229), .B(n12228), .ZN(
        P3_U3180) );
  MUX2_X1 U14582 ( .A(n12356), .B(P3_DATAO_REG_31__SCAN_IN), .S(n12245), .Z(
        P3_U3522) );
  MUX2_X1 U14583 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(n12231), .S(P3_U3897), .Z(
        P3_U3521) );
  INV_X1 U14584 ( .A(n12232), .ZN(n12423) );
  MUX2_X1 U14585 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(n12423), .S(P3_U3897), .Z(
        P3_U3520) );
  INV_X1 U14586 ( .A(n12402), .ZN(n12435) );
  MUX2_X1 U14587 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12435), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14588 ( .A(n12464), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12245), .Z(
        P3_U3517) );
  MUX2_X1 U14589 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12395), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14590 ( .A(n12465), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12245), .Z(
        P3_U3515) );
  MUX2_X1 U14591 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n12389), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U14592 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12386), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14593 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12381), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14594 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n12233), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U14595 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12571), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14596 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12372), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14597 ( .A(n12570), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12245), .Z(
        P3_U3507) );
  MUX2_X1 U14598 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12234), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U14599 ( .A(n12235), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12245), .Z(
        P3_U3505) );
  MUX2_X1 U14600 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n12236), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14601 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12237), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14602 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n12238), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U14603 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12239), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14604 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12240), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14605 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12241), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14606 ( .A(n12242), .B(P3_DATAO_REG_5__SCAN_IN), .S(n12245), .Z(
        P3_U3496) );
  MUX2_X1 U14607 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n15192), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14608 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12243), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14609 ( .A(n15365), .B(P3_DATAO_REG_2__SCAN_IN), .S(n12245), .Z(
        P3_U3493) );
  MUX2_X1 U14610 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n12244), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U14611 ( .A(n15367), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12245), .Z(
        P3_U3491) );
  INV_X1 U14612 ( .A(n12246), .ZN(n12248) );
  INV_X1 U14613 ( .A(n12282), .ZN(n12271) );
  INV_X1 U14614 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12649) );
  NAND2_X1 U14615 ( .A1(n12271), .A2(n12649), .ZN(n12250) );
  NAND2_X1 U14616 ( .A1(n12282), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12283) );
  AND2_X1 U14617 ( .A1(n12250), .A2(n12283), .ZN(n12264) );
  XNOR2_X1 U14618 ( .A(n12282), .B(P3_REG2_REG_14__SCAN_IN), .ZN(n12258) );
  INV_X1 U14619 ( .A(n12258), .ZN(n12251) );
  MUX2_X1 U14620 ( .A(n12264), .B(n12251), .S(n12340), .Z(n12252) );
  OAI211_X1 U14621 ( .C1(n12253), .C2(n12252), .A(n12286), .B(n15305), .ZN(
        n12273) );
  INV_X1 U14622 ( .A(n12254), .ZN(n12256) );
  AOI21_X1 U14623 ( .B1(n12258), .B2(n12257), .A(n12274), .ZN(n12269) );
  NAND2_X1 U14624 ( .A1(n12260), .A2(n12259), .ZN(n12262) );
  NAND2_X1 U14625 ( .A1(n12262), .A2(n12261), .ZN(n12263) );
  NAND2_X1 U14626 ( .A1(n12264), .A2(n12263), .ZN(n12277) );
  OAI21_X1 U14627 ( .B1(n12264), .B2(n12263), .A(n12277), .ZN(n12267) );
  NOR2_X1 U14628 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n7871), .ZN(n12266) );
  NOR2_X1 U14629 ( .A1(n15308), .A2(n13658), .ZN(n12265) );
  AOI211_X1 U14630 ( .C1(n15329), .C2(n12267), .A(n12266), .B(n12265), .ZN(
        n12268) );
  OAI21_X1 U14631 ( .B1(n12269), .B2(n15333), .A(n12268), .ZN(n12270) );
  AOI21_X1 U14632 ( .B1(n12271), .B2(n15266), .A(n12270), .ZN(n12272) );
  NAND2_X1 U14633 ( .A1(n12273), .A2(n12272), .ZN(P3_U3196) );
  INV_X1 U14634 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12276) );
  AOI21_X1 U14635 ( .B1(n12276), .B2(n12275), .A(n12304), .ZN(n12294) );
  NAND2_X1 U14636 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n12278), .ZN(n12318) );
  OAI21_X1 U14637 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n12278), .A(n12318), 
        .ZN(n12292) );
  NOR2_X1 U14638 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12279), .ZN(n12280) );
  AOI21_X1 U14639 ( .B1(n15326), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n12280), 
        .ZN(n12281) );
  OAI21_X1 U14640 ( .B1(n15320), .B2(n12317), .A(n12281), .ZN(n12291) );
  NAND2_X1 U14641 ( .A1(n12282), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12284) );
  MUX2_X1 U14642 ( .A(n12284), .B(n12283), .S(n14735), .Z(n12285) );
  NAND2_X1 U14643 ( .A1(n12286), .A2(n12285), .ZN(n12296) );
  XNOR2_X1 U14644 ( .A(n12296), .B(n12317), .ZN(n12288) );
  MUX2_X1 U14645 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n14735), .Z(n12287) );
  NAND2_X1 U14646 ( .A1(n12288), .A2(n12287), .ZN(n12289) );
  AOI21_X1 U14647 ( .B1(n12295), .B2(n12289), .A(n15322), .ZN(n12290) );
  AOI211_X1 U14648 ( .C1(n12292), .C2(n15329), .A(n12291), .B(n12290), .ZN(
        n12293) );
  OAI21_X1 U14649 ( .B1(n12294), .B2(n15333), .A(n12293), .ZN(P3_U3197) );
  MUX2_X1 U14650 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n14735), .Z(n12301) );
  MUX2_X1 U14651 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n14735), .Z(n12299) );
  INV_X1 U14652 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12306) );
  INV_X1 U14653 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13686) );
  MUX2_X1 U14654 ( .A(n12306), .B(n13686), .S(n14735), .Z(n12297) );
  OAI21_X1 U14655 ( .B1(n12296), .B2(n12317), .A(n12295), .ZN(n14740) );
  OAI21_X1 U14656 ( .B1(n12307), .B2(n12297), .A(n14740), .ZN(n12298) );
  NAND2_X1 U14657 ( .A1(n12297), .A2(n12307), .ZN(n14739) );
  NAND2_X1 U14658 ( .A1(n12298), .A2(n14739), .ZN(n14757) );
  XNOR2_X1 U14659 ( .A(n12299), .B(n12320), .ZN(n14758) );
  NOR2_X1 U14660 ( .A1(n14757), .A2(n14758), .ZN(n14756) );
  AOI21_X1 U14661 ( .B1(n12299), .B2(n12320), .A(n14756), .ZN(n12345) );
  XNOR2_X1 U14662 ( .A(n12345), .B(n12344), .ZN(n12300) );
  NOR2_X1 U14663 ( .A1(n12300), .A2(n12301), .ZN(n12343) );
  AOI21_X1 U14664 ( .B1(n12301), .B2(n12300), .A(n12343), .ZN(n12330) );
  INV_X1 U14665 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14762) );
  NOR2_X1 U14666 ( .A1(n12303), .A2(n12302), .ZN(n12305) );
  NAND2_X1 U14667 ( .A1(n14733), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n14737) );
  NAND2_X1 U14668 ( .A1(n12307), .A2(n12306), .ZN(n12308) );
  NAND2_X1 U14669 ( .A1(n14737), .A2(n12308), .ZN(n14746) );
  NOR2_X1 U14670 ( .A1(n12309), .A2(n14753), .ZN(n12311) );
  INV_X1 U14671 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12557) );
  NOR2_X1 U14672 ( .A1(n12344), .A2(n12557), .ZN(n12331) );
  AOI21_X1 U14673 ( .B1(n12344), .B2(n12557), .A(n12331), .ZN(n12310) );
  INV_X1 U14674 ( .A(n12333), .ZN(n12313) );
  NOR3_X1 U14675 ( .A1(n14763), .A2(n12311), .A3(n12310), .ZN(n12312) );
  OAI21_X1 U14676 ( .B1(n12313), .B2(n12312), .A(n15264), .ZN(n12329) );
  INV_X1 U14677 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n12315) );
  OAI21_X1 U14678 ( .B1(n15308), .B2(n12315), .A(n12314), .ZN(n12327) );
  NAND2_X1 U14679 ( .A1(n12317), .A2(n12316), .ZN(n12319) );
  XNOR2_X1 U14680 ( .A(n14733), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n14742) );
  NAND2_X1 U14681 ( .A1(n14733), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n14736) );
  XNOR2_X1 U14682 ( .A(n14753), .B(n12321), .ZN(n14755) );
  NAND2_X1 U14683 ( .A1(P3_REG1_REG_17__SCAN_IN), .A2(n14755), .ZN(n14754) );
  NAND2_X1 U14684 ( .A1(n12321), .A2(n12320), .ZN(n12322) );
  INV_X1 U14685 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12634) );
  XNOR2_X1 U14686 ( .A(n12344), .B(n12634), .ZN(n12323) );
  INV_X1 U14687 ( .A(n12335), .ZN(n12325) );
  NAND3_X1 U14688 ( .A1(n14754), .A2(n12323), .A3(n12322), .ZN(n12324) );
  AOI21_X1 U14689 ( .B1(n12325), .B2(n12324), .A(n15297), .ZN(n12326) );
  AOI211_X1 U14690 ( .C1(n15266), .C2(n12344), .A(n12327), .B(n12326), .ZN(
        n12328) );
  OAI211_X1 U14691 ( .C1(n12330), .C2(n15322), .A(n12329), .B(n12328), .ZN(
        P3_U3200) );
  INV_X1 U14692 ( .A(n12331), .ZN(n12332) );
  NAND2_X1 U14693 ( .A1(n12333), .A2(n12332), .ZN(n12334) );
  XNOR2_X1 U14694 ( .A(n6687), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12341) );
  XNOR2_X1 U14695 ( .A(n12334), .B(n12341), .ZN(n12352) );
  AOI21_X1 U14696 ( .B1(P3_REG1_REG_18__SCAN_IN), .B2(n12336), .A(n12335), 
        .ZN(n12337) );
  XNOR2_X1 U14697 ( .A(n6687), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12342) );
  XNOR2_X1 U14698 ( .A(n12337), .B(n12342), .ZN(n12350) );
  NAND2_X1 U14699 ( .A1(n15326), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12338) );
  OAI211_X1 U14700 ( .C1(n15320), .C2(n6687), .A(n12339), .B(n12338), .ZN(
        n12349) );
  MUX2_X1 U14701 ( .A(n12342), .B(n12341), .S(n12340), .Z(n12346) );
  NOR2_X1 U14702 ( .A1(n12347), .A2(n15322), .ZN(n12348) );
  OAI21_X1 U14703 ( .B1(n12352), .B2(n15333), .A(n12351), .ZN(P3_U3201) );
  INV_X1 U14704 ( .A(P3_B_REG_SCAN_IN), .ZN(n12353) );
  NOR2_X1 U14705 ( .A1(n12354), .A2(n12353), .ZN(n12355) );
  OR2_X1 U14706 ( .A1(n15351), .A2(n12355), .ZN(n12403) );
  INV_X1 U14707 ( .A(n12403), .ZN(n12357) );
  NAND2_X1 U14708 ( .A1(n12357), .A2(n12356), .ZN(n14768) );
  OAI22_X1 U14709 ( .A1(n12443), .A2(n14768), .B1(n12358), .B2(n12555), .ZN(
        n12360) );
  AOI21_X1 U14710 ( .B1(n12443), .B2(P3_REG2_REG_31__SCAN_IN), .A(n12360), 
        .ZN(n12359) );
  OAI21_X1 U14711 ( .B1(n12654), .B2(n12578), .A(n12359), .ZN(P3_U3202) );
  AOI21_X1 U14712 ( .B1(n12443), .B2(P3_REG2_REG_30__SCAN_IN), .A(n12360), 
        .ZN(n12361) );
  OAI21_X1 U14713 ( .B1(n12362), .B2(n12578), .A(n12361), .ZN(P3_U3203) );
  NAND2_X1 U14714 ( .A1(n12365), .A2(n12570), .ZN(n12366) );
  AND2_X1 U14715 ( .A1(n12367), .A2(n12366), .ZN(n12368) );
  INV_X1 U14716 ( .A(n12371), .ZN(n12374) );
  NAND2_X1 U14717 ( .A1(n12636), .A2(n12372), .ZN(n12373) );
  OR2_X1 U14718 ( .A1(n12560), .A2(n12571), .ZN(n12531) );
  INV_X1 U14719 ( .A(n12376), .ZN(n12377) );
  AND2_X1 U14720 ( .A1(n12531), .A2(n12377), .ZN(n12378) );
  NAND2_X1 U14721 ( .A1(n12522), .A2(n12521), .ZN(n12520) );
  NAND2_X1 U14722 ( .A1(n12626), .A2(n12381), .ZN(n12382) );
  OR2_X1 U14723 ( .A1(n12683), .A2(n12384), .ZN(n12385) );
  NOR2_X1 U14724 ( .A1(n12387), .A2(n12386), .ZN(n12388) );
  NAND2_X1 U14725 ( .A1(n12486), .A2(n12490), .ZN(n12391) );
  NAND2_X1 U14726 ( .A1(n12492), .A2(n12389), .ZN(n12390) );
  AND2_X1 U14727 ( .A1(n12392), .A2(n12465), .ZN(n12393) );
  NAND2_X1 U14728 ( .A1(n12396), .A2(n12395), .ZN(n12445) );
  NAND2_X1 U14729 ( .A1(n12398), .A2(n12464), .ZN(n12397) );
  AND2_X1 U14730 ( .A1(n12445), .A2(n12397), .ZN(n12399) );
  OR2_X1 U14731 ( .A1(n12591), .A2(n12422), .ZN(n12400) );
  NOR2_X1 U14732 ( .A1(n12404), .A2(n12403), .ZN(n12405) );
  INV_X1 U14733 ( .A(n12585), .ZN(n12415) );
  XNOR2_X1 U14734 ( .A(n12409), .B(n12408), .ZN(n12586) );
  AOI22_X1 U14735 ( .A1(n12443), .A2(P3_REG2_REG_29__SCAN_IN), .B1(n12411), 
        .B2(n15379), .ZN(n12412) );
  OAI21_X1 U14736 ( .B1(n12657), .B2(n12578), .A(n12412), .ZN(n12413) );
  AOI21_X1 U14737 ( .B1(n12586), .B2(n12581), .A(n12413), .ZN(n12414) );
  OAI21_X1 U14738 ( .B1(n12415), .B2(n12443), .A(n12414), .ZN(P3_U3204) );
  INV_X1 U14739 ( .A(n12416), .ZN(n12417) );
  INV_X1 U14740 ( .A(n12588), .ZN(n12431) );
  NAND2_X1 U14741 ( .A1(n12420), .A2(n12419), .ZN(n12421) );
  AOI22_X1 U14742 ( .A1(n12423), .A2(n15366), .B1(n12406), .B2(n12422), .ZN(
        n12424) );
  NAND2_X1 U14743 ( .A1(n12425), .A2(n12424), .ZN(n12589) );
  INV_X1 U14744 ( .A(n12426), .ZN(n12660) );
  AOI22_X1 U14745 ( .A1(n12443), .A2(P3_REG2_REG_28__SCAN_IN), .B1(n15379), 
        .B2(n12427), .ZN(n12428) );
  OAI21_X1 U14746 ( .B1(n12660), .B2(n12578), .A(n12428), .ZN(n12429) );
  AOI21_X1 U14747 ( .B1(n12589), .B2(n15380), .A(n12429), .ZN(n12430) );
  OAI21_X1 U14748 ( .B1(n12431), .B2(n12563), .A(n12430), .ZN(P3_U3205) );
  INV_X1 U14749 ( .A(n12432), .ZN(n12434) );
  OAI21_X1 U14750 ( .B1(n12434), .B2(n7039), .A(n12433), .ZN(n12436) );
  AOI21_X1 U14751 ( .B1(n7039), .B2(n12437), .A(n6691), .ZN(n12594) );
  AOI22_X1 U14752 ( .A1(n12443), .A2(P3_REG2_REG_27__SCAN_IN), .B1(n15379), 
        .B2(n12438), .ZN(n12439) );
  OAI21_X1 U14753 ( .B1(n12440), .B2(n12578), .A(n12439), .ZN(n12441) );
  AOI21_X1 U14754 ( .B1(n6824), .B2(n12581), .A(n12441), .ZN(n12442) );
  OAI21_X1 U14755 ( .B1(n12593), .B2(n12443), .A(n12442), .ZN(P3_U3206) );
  XNOR2_X1 U14756 ( .A(n12444), .B(n12447), .ZN(n12453) );
  NAND2_X1 U14757 ( .A1(n12461), .A2(n12445), .ZN(n12446) );
  XOR2_X1 U14758 ( .A(n12447), .B(n12446), .Z(n12451) );
  OAI22_X1 U14759 ( .A1(n12449), .A2(n15351), .B1(n12448), .B2(n15353), .ZN(
        n12450) );
  AOI21_X1 U14760 ( .B1(n12451), .B2(n15369), .A(n12450), .ZN(n12452) );
  OAI21_X1 U14761 ( .B1(n15373), .B2(n12453), .A(n12452), .ZN(n12596) );
  INV_X1 U14762 ( .A(n12596), .ZN(n12458) );
  INV_X1 U14763 ( .A(n12453), .ZN(n12597) );
  AOI22_X1 U14764 ( .A1(n12443), .A2(P3_REG2_REG_26__SCAN_IN), .B1(n15379), 
        .B2(n12454), .ZN(n12455) );
  OAI21_X1 U14765 ( .B1(n12664), .B2(n12578), .A(n12455), .ZN(n12456) );
  AOI21_X1 U14766 ( .B1(n12597), .B2(n12472), .A(n12456), .ZN(n12457) );
  OAI21_X1 U14767 ( .B1(n12458), .B2(n12443), .A(n12457), .ZN(P3_U3207) );
  XNOR2_X1 U14768 ( .A(n12459), .B(n12462), .ZN(n12468) );
  INV_X1 U14769 ( .A(n12460), .ZN(n12463) );
  OAI211_X1 U14770 ( .C1(n12463), .C2(n12462), .A(n15369), .B(n12461), .ZN(
        n12467) );
  AOI22_X1 U14771 ( .A1(n12406), .A2(n12465), .B1(n15366), .B2(n12464), .ZN(
        n12466) );
  OAI211_X1 U14772 ( .C1(n15373), .C2(n12468), .A(n12467), .B(n12466), .ZN(
        n12600) );
  INV_X1 U14773 ( .A(n12600), .ZN(n12474) );
  INV_X1 U14774 ( .A(n12468), .ZN(n12601) );
  AOI22_X1 U14775 ( .A1(n12443), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n15379), 
        .B2(n12469), .ZN(n12470) );
  OAI21_X1 U14776 ( .B1(n12668), .B2(n12578), .A(n12470), .ZN(n12471) );
  AOI21_X1 U14777 ( .B1(n12601), .B2(n12472), .A(n12471), .ZN(n12473) );
  OAI21_X1 U14778 ( .B1(n12474), .B2(n12443), .A(n12473), .ZN(P3_U3208) );
  XNOR2_X1 U14779 ( .A(n12475), .B(n12478), .ZN(n12477) );
  OAI21_X1 U14780 ( .B1(n12477), .B2(n15359), .A(n12476), .ZN(n12604) );
  INV_X1 U14781 ( .A(n12604), .ZN(n12485) );
  OAI21_X1 U14782 ( .B1(n12480), .B2(n7053), .A(n12479), .ZN(n12605) );
  AOI22_X1 U14783 ( .A1(n12443), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n15379), 
        .B2(n12481), .ZN(n12482) );
  OAI21_X1 U14784 ( .B1(n12672), .B2(n12578), .A(n12482), .ZN(n12483) );
  AOI21_X1 U14785 ( .B1(n12605), .B2(n12581), .A(n12483), .ZN(n12484) );
  OAI21_X1 U14786 ( .B1(n12485), .B2(n12443), .A(n12484), .ZN(P3_U3209) );
  XNOR2_X1 U14787 ( .A(n12486), .B(n12490), .ZN(n12487) );
  OAI222_X1 U14788 ( .A1(n15351), .A2(n12489), .B1(n15353), .B2(n12488), .C1(
        n12487), .C2(n15359), .ZN(n12608) );
  INV_X1 U14789 ( .A(n12608), .ZN(n12497) );
  XNOR2_X1 U14790 ( .A(n12491), .B(n12490), .ZN(n12609) );
  INV_X1 U14791 ( .A(n12492), .ZN(n12676) );
  AOI22_X1 U14792 ( .A1(n12443), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n15379), 
        .B2(n12493), .ZN(n12494) );
  OAI21_X1 U14793 ( .B1(n12676), .B2(n12578), .A(n12494), .ZN(n12495) );
  AOI21_X1 U14794 ( .B1(n12609), .B2(n12581), .A(n12495), .ZN(n12496) );
  OAI21_X1 U14795 ( .B1(n12497), .B2(n12443), .A(n12496), .ZN(P3_U3210) );
  XNOR2_X1 U14796 ( .A(n12498), .B(n12503), .ZN(n12501) );
  INV_X1 U14797 ( .A(n12499), .ZN(n12500) );
  AOI21_X1 U14798 ( .B1(n12501), .B2(n15369), .A(n12500), .ZN(n12614) );
  XNOR2_X1 U14799 ( .A(n12502), .B(n12503), .ZN(n12612) );
  AOI22_X1 U14800 ( .A1(n12443), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n15379), 
        .B2(n12504), .ZN(n12505) );
  OAI21_X1 U14801 ( .B1(n12680), .B2(n12578), .A(n12505), .ZN(n12506) );
  AOI21_X1 U14802 ( .B1(n12612), .B2(n12581), .A(n12506), .ZN(n12507) );
  OAI21_X1 U14803 ( .B1(n12614), .B2(n12443), .A(n12507), .ZN(P3_U3211) );
  NAND2_X1 U14804 ( .A1(n12508), .A2(n12513), .ZN(n12509) );
  NAND2_X1 U14805 ( .A1(n12510), .A2(n12509), .ZN(n12512) );
  AOI21_X1 U14806 ( .B1(n12512), .B2(n15369), .A(n12511), .ZN(n12619) );
  XNOR2_X1 U14807 ( .A(n12514), .B(n12383), .ZN(n12617) );
  INV_X1 U14808 ( .A(n12683), .ZN(n12517) );
  AOI22_X1 U14809 ( .A1(n12443), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15379), 
        .B2(n12515), .ZN(n12516) );
  OAI21_X1 U14810 ( .B1(n12517), .B2(n12578), .A(n12516), .ZN(n12518) );
  AOI21_X1 U14811 ( .B1(n12617), .B2(n12581), .A(n12518), .ZN(n12519) );
  OAI21_X1 U14812 ( .B1(n12619), .B2(n12443), .A(n12519), .ZN(P3_U3212) );
  OAI211_X1 U14813 ( .C1(n12522), .C2(n12521), .A(n12520), .B(n15369), .ZN(
        n12524) );
  AND2_X1 U14814 ( .A1(n12524), .A2(n12523), .ZN(n12624) );
  XNOR2_X1 U14815 ( .A(n12525), .B(n12526), .ZN(n12622) );
  AOI22_X1 U14816 ( .A1(n12443), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15379), 
        .B2(n12527), .ZN(n12528) );
  OAI21_X1 U14817 ( .B1(n12690), .B2(n12578), .A(n12528), .ZN(n12529) );
  AOI21_X1 U14818 ( .B1(n12622), .B2(n12581), .A(n12529), .ZN(n12530) );
  OAI21_X1 U14819 ( .B1(n12624), .B2(n12443), .A(n12530), .ZN(P3_U3213) );
  NAND2_X1 U14820 ( .A1(n12547), .A2(n12531), .ZN(n12532) );
  XOR2_X1 U14821 ( .A(n12536), .B(n12532), .Z(n12533) );
  OAI222_X1 U14822 ( .A1(n15351), .A2(n12535), .B1(n15353), .B2(n12534), .C1(
        n12533), .C2(n15359), .ZN(n12628) );
  INV_X1 U14823 ( .A(n12628), .ZN(n12542) );
  XNOR2_X1 U14824 ( .A(n12537), .B(n12536), .ZN(n12629) );
  AOI22_X1 U14825 ( .A1(n12443), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15379), 
        .B2(n12538), .ZN(n12539) );
  OAI21_X1 U14826 ( .B1(n12694), .B2(n12578), .A(n12539), .ZN(n12540) );
  AOI21_X1 U14827 ( .B1(n12629), .B2(n12581), .A(n12540), .ZN(n12541) );
  OAI21_X1 U14828 ( .B1(n12542), .B2(n12443), .A(n12541), .ZN(P3_U3214) );
  NAND2_X1 U14829 ( .A1(n12573), .A2(n12543), .ZN(n12544) );
  NAND2_X1 U14830 ( .A1(n12544), .A2(n12375), .ZN(n12546) );
  AND2_X1 U14831 ( .A1(n12546), .A2(n12545), .ZN(n12633) );
  INV_X1 U14832 ( .A(n12633), .ZN(n12564) );
  INV_X1 U14833 ( .A(n12547), .ZN(n12548) );
  AOI21_X1 U14834 ( .B1(n12550), .B2(n12549), .A(n12548), .ZN(n12551) );
  OAI222_X1 U14835 ( .A1(n15351), .A2(n12553), .B1(n15353), .B2(n12552), .C1(
        n15359), .C2(n12551), .ZN(n12632) );
  NAND2_X1 U14836 ( .A1(n12632), .A2(n15380), .ZN(n12562) );
  INV_X1 U14837 ( .A(n12554), .ZN(n12556) );
  OAI22_X1 U14838 ( .A1(n15380), .A2(n12557), .B1(n12556), .B2(n12555), .ZN(
        n12558) );
  AOI21_X1 U14839 ( .B1(n12560), .B2(n12559), .A(n12558), .ZN(n12561) );
  OAI211_X1 U14840 ( .C1(n12564), .C2(n12563), .A(n12562), .B(n12561), .ZN(
        P3_U3215) );
  OR2_X1 U14841 ( .A1(n12566), .A2(n12565), .ZN(n12568) );
  NAND2_X1 U14842 ( .A1(n12568), .A2(n12567), .ZN(n12569) );
  XNOR2_X1 U14843 ( .A(n12569), .B(n12574), .ZN(n12572) );
  AOI222_X1 U14844 ( .A1(n15369), .A2(n12572), .B1(n12571), .B2(n15366), .C1(
        n12570), .C2(n12406), .ZN(n12639) );
  OAI21_X1 U14845 ( .B1(n12575), .B2(n12574), .A(n12573), .ZN(n12637) );
  INV_X1 U14846 ( .A(n12636), .ZN(n12579) );
  AOI22_X1 U14847 ( .A1(n12443), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15379), 
        .B2(n12576), .ZN(n12577) );
  OAI21_X1 U14848 ( .B1(n12579), .B2(n12578), .A(n12577), .ZN(n12580) );
  AOI21_X1 U14849 ( .B1(n12637), .B2(n12581), .A(n12580), .ZN(n12582) );
  OAI21_X1 U14850 ( .B1(n12639), .B2(n12443), .A(n12582), .ZN(P3_U3216) );
  INV_X1 U14851 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n12583) );
  MUX2_X1 U14852 ( .A(n12583), .B(n14768), .S(n15436), .Z(n12584) );
  OAI21_X1 U14853 ( .B1(n12654), .B2(n12651), .A(n12584), .ZN(P3_U3490) );
  INV_X1 U14854 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n12587) );
  INV_X1 U14855 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n12590) );
  NAND2_X1 U14856 ( .A1(n12591), .A2(n14770), .ZN(n12592) );
  MUX2_X1 U14857 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n12661), .S(n15436), .Z(
        P3_U3486) );
  INV_X1 U14858 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12598) );
  INV_X1 U14859 ( .A(n12595), .ZN(n15410) );
  AOI21_X1 U14860 ( .B1(n15410), .B2(n12597), .A(n12596), .ZN(n12662) );
  MUX2_X1 U14861 ( .A(n12598), .B(n12662), .S(n15436), .Z(n12599) );
  OAI21_X1 U14862 ( .B1(n12664), .B2(n12651), .A(n12599), .ZN(P3_U3485) );
  INV_X1 U14863 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n12602) );
  AOI21_X1 U14864 ( .B1(n15410), .B2(n12601), .A(n12600), .ZN(n12665) );
  MUX2_X1 U14865 ( .A(n12602), .B(n12665), .S(n15436), .Z(n12603) );
  OAI21_X1 U14866 ( .B1(n12668), .B2(n12651), .A(n12603), .ZN(P3_U3484) );
  INV_X1 U14867 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12606) );
  AOI21_X1 U14868 ( .B1(n14775), .B2(n12605), .A(n12604), .ZN(n12669) );
  MUX2_X1 U14869 ( .A(n12606), .B(n12669), .S(n15436), .Z(n12607) );
  OAI21_X1 U14870 ( .B1(n12672), .B2(n12651), .A(n12607), .ZN(P3_U3483) );
  INV_X1 U14871 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12610) );
  AOI21_X1 U14872 ( .B1(n14775), .B2(n12609), .A(n12608), .ZN(n12673) );
  MUX2_X1 U14873 ( .A(n12610), .B(n12673), .S(n15436), .Z(n12611) );
  OAI21_X1 U14874 ( .B1(n12676), .B2(n12651), .A(n12611), .ZN(P3_U3482) );
  NAND2_X1 U14875 ( .A1(n12612), .A2(n14775), .ZN(n12613) );
  NAND2_X1 U14876 ( .A1(n12614), .A2(n12613), .ZN(n12677) );
  MUX2_X1 U14877 ( .A(P3_REG1_REG_22__SCAN_IN), .B(n12677), .S(n15436), .Z(
        n12615) );
  INV_X1 U14878 ( .A(n12615), .ZN(n12616) );
  OAI21_X1 U14879 ( .B1(n12680), .B2(n12651), .A(n12616), .ZN(P3_U3481) );
  NAND2_X1 U14880 ( .A1(n12617), .A2(n14775), .ZN(n12618) );
  NAND2_X1 U14881 ( .A1(n12619), .A2(n12618), .ZN(n12681) );
  MUX2_X1 U14882 ( .A(n12681), .B(P3_REG1_REG_21__SCAN_IN), .S(n15433), .Z(
        n12620) );
  AOI21_X1 U14883 ( .B1(n6853), .B2(n12683), .A(n12620), .ZN(n12621) );
  INV_X1 U14884 ( .A(n12621), .ZN(P3_U3480) );
  NAND2_X1 U14885 ( .A1(n12622), .A2(n14775), .ZN(n12623) );
  NAND2_X1 U14886 ( .A1(n12624), .A2(n12623), .ZN(n12686) );
  MUX2_X1 U14887 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n12686), .S(n15436), .Z(
        n12625) );
  AOI21_X1 U14888 ( .B1(n6853), .B2(n12626), .A(n12625), .ZN(n12627) );
  INV_X1 U14889 ( .A(n12627), .ZN(P3_U3479) );
  INV_X1 U14890 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12630) );
  AOI21_X1 U14891 ( .B1(n12629), .B2(n14775), .A(n12628), .ZN(n12691) );
  MUX2_X1 U14892 ( .A(n12630), .B(n12691), .S(n15436), .Z(n12631) );
  OAI21_X1 U14893 ( .B1(n12651), .B2(n12694), .A(n12631), .ZN(P3_U3478) );
  AOI21_X1 U14894 ( .B1(n12633), .B2(n14775), .A(n12632), .ZN(n12695) );
  MUX2_X1 U14895 ( .A(n12634), .B(n12695), .S(n15436), .Z(n12635) );
  OAI21_X1 U14896 ( .B1(n12697), .B2(n12651), .A(n12635), .ZN(P3_U3477) );
  AOI22_X1 U14897 ( .A1(n12637), .A2(n14775), .B1(n14770), .B2(n12636), .ZN(
        n12638) );
  NAND2_X1 U14898 ( .A1(n12639), .A2(n12638), .ZN(n12698) );
  MUX2_X1 U14899 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n12698), .S(n15436), .Z(
        P3_U3476) );
  AOI21_X1 U14900 ( .B1(n14775), .B2(n12641), .A(n12640), .ZN(n12699) );
  MUX2_X1 U14901 ( .A(n13686), .B(n12699), .S(n15436), .Z(n12642) );
  OAI21_X1 U14902 ( .B1(n12702), .B2(n12651), .A(n12642), .ZN(P3_U3475) );
  INV_X1 U14903 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12645) );
  AOI21_X1 U14904 ( .B1(n14775), .B2(n12644), .A(n12643), .ZN(n12703) );
  MUX2_X1 U14905 ( .A(n12645), .B(n12703), .S(n15436), .Z(n12646) );
  OAI21_X1 U14906 ( .B1(n12706), .B2(n12651), .A(n12646), .ZN(P3_U3474) );
  AOI21_X1 U14907 ( .B1(n14775), .B2(n12648), .A(n12647), .ZN(n12708) );
  MUX2_X1 U14908 ( .A(n12649), .B(n12708), .S(n15436), .Z(n12650) );
  OAI21_X1 U14909 ( .B1(n12651), .B2(n12711), .A(n12650), .ZN(P3_U3473) );
  INV_X1 U14910 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n12652) );
  MUX2_X1 U14911 ( .A(n12652), .B(n14768), .S(n12707), .Z(n12653) );
  OAI21_X1 U14912 ( .B1(n12654), .B2(n12712), .A(n12653), .ZN(P3_U3458) );
  OAI21_X1 U14913 ( .B1(n12657), .B2(n12712), .A(n12656), .ZN(P3_U3456) );
  OAI21_X1 U14914 ( .B1(n12660), .B2(n12712), .A(n12659), .ZN(P3_U3455) );
  MUX2_X1 U14915 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n12661), .S(n12707), .Z(
        P3_U3454) );
  INV_X1 U14916 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13574) );
  MUX2_X1 U14917 ( .A(n13574), .B(n12662), .S(n12707), .Z(n12663) );
  OAI21_X1 U14918 ( .B1(n12664), .B2(n12712), .A(n12663), .ZN(P3_U3453) );
  INV_X1 U14919 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n12666) );
  MUX2_X1 U14920 ( .A(n12666), .B(n12665), .S(n12707), .Z(n12667) );
  OAI21_X1 U14921 ( .B1(n12668), .B2(n12712), .A(n12667), .ZN(P3_U3452) );
  INV_X1 U14922 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n12670) );
  MUX2_X1 U14923 ( .A(n12670), .B(n12669), .S(n12707), .Z(n12671) );
  OAI21_X1 U14924 ( .B1(n12672), .B2(n12712), .A(n12671), .ZN(P3_U3451) );
  INV_X1 U14925 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n12674) );
  MUX2_X1 U14926 ( .A(n12674), .B(n12673), .S(n12707), .Z(n12675) );
  OAI21_X1 U14927 ( .B1(n12676), .B2(n12712), .A(n12675), .ZN(P3_U3450) );
  MUX2_X1 U14928 ( .A(P3_REG0_REG_22__SCAN_IN), .B(n12677), .S(n12707), .Z(
        n12678) );
  INV_X1 U14929 ( .A(n12678), .ZN(n12679) );
  OAI21_X1 U14930 ( .B1(n12680), .B2(n12712), .A(n12679), .ZN(P3_U3449) );
  MUX2_X1 U14931 ( .A(n12681), .B(P3_REG0_REG_21__SCAN_IN), .S(n15419), .Z(
        n12682) );
  AOI21_X1 U14932 ( .B1(n12684), .B2(n12683), .A(n12682), .ZN(n12685) );
  INV_X1 U14933 ( .A(n12685), .ZN(P3_U3448) );
  INV_X1 U14934 ( .A(n12686), .ZN(n12688) );
  MUX2_X1 U14935 ( .A(n12688), .B(n12687), .S(n15419), .Z(n12689) );
  OAI21_X1 U14936 ( .B1(n12690), .B2(n12712), .A(n12689), .ZN(P3_U3447) );
  INV_X1 U14937 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n12692) );
  MUX2_X1 U14938 ( .A(n12692), .B(n12691), .S(n12707), .Z(n12693) );
  OAI21_X1 U14939 ( .B1(n12712), .B2(n12694), .A(n12693), .ZN(P3_U3446) );
  INV_X1 U14940 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13710) );
  MUX2_X1 U14941 ( .A(n13710), .B(n12695), .S(n12707), .Z(n12696) );
  OAI21_X1 U14942 ( .B1(n12697), .B2(n12712), .A(n12696), .ZN(P3_U3444) );
  MUX2_X1 U14943 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n12698), .S(n12707), .Z(
        P3_U3441) );
  INV_X1 U14944 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n12700) );
  MUX2_X1 U14945 ( .A(n12700), .B(n12699), .S(n12707), .Z(n12701) );
  OAI21_X1 U14946 ( .B1(n12702), .B2(n12712), .A(n12701), .ZN(P3_U3438) );
  INV_X1 U14947 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n12704) );
  MUX2_X1 U14948 ( .A(n12704), .B(n12703), .S(n12707), .Z(n12705) );
  OAI21_X1 U14949 ( .B1(n12706), .B2(n12712), .A(n12705), .ZN(P3_U3435) );
  INV_X1 U14950 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n12709) );
  MUX2_X1 U14951 ( .A(n12709), .B(n12708), .S(n12707), .Z(n12710) );
  OAI21_X1 U14952 ( .B1(n12712), .B2(n12711), .A(n12710), .ZN(P3_U3432) );
  MUX2_X1 U14953 ( .A(n12713), .B(P3_D_REG_1__SCAN_IN), .S(n12714), .Z(
        P3_U3377) );
  MUX2_X1 U14954 ( .A(n12715), .B(P3_D_REG_0__SCAN_IN), .S(n12714), .Z(
        P3_U3376) );
  INV_X1 U14955 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n12716) );
  NAND3_X1 U14956 ( .A1(n12716), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n12717) );
  OAI22_X1 U14957 ( .A1(n7621), .A2(n12717), .B1(n13683), .B2(n12725), .ZN(
        n12718) );
  AOI21_X1 U14958 ( .B1(n12720), .B2(n12719), .A(n12718), .ZN(n12721) );
  INV_X1 U14959 ( .A(n12721), .ZN(P3_U3264) );
  INV_X1 U14960 ( .A(n12722), .ZN(n12723) );
  OAI222_X1 U14961 ( .A1(n12726), .A2(P3_U3151), .B1(n12725), .B2(n12724), 
        .C1(n11991), .C2(n12723), .ZN(P3_U3265) );
  INV_X1 U14962 ( .A(n12727), .ZN(n12729) );
  NAND2_X1 U14963 ( .A1(n12732), .A2(n10117), .ZN(n12735) );
  AOI22_X1 U14964 ( .A1(n12892), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n12733), 
        .B2(n13214), .ZN(n12734) );
  XNOR2_X1 U14965 ( .A(n14027), .B(n11155), .ZN(n12738) );
  NAND2_X1 U14966 ( .A1(n13261), .A2(n6611), .ZN(n12737) );
  NAND2_X1 U14967 ( .A1(n12738), .A2(n12737), .ZN(n12878) );
  NOR2_X1 U14968 ( .A1(n12738), .A2(n12737), .ZN(n12879) );
  NAND2_X1 U14969 ( .A1(n12740), .A2(n12739), .ZN(n12937) );
  NAND2_X1 U14970 ( .A1(n12741), .A2(n10117), .ZN(n12743) );
  NAND2_X1 U14971 ( .A1(n12892), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n12742) );
  XNOR2_X1 U14972 ( .A(n14022), .B(n11155), .ZN(n12751) );
  INV_X1 U14973 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n12943) );
  AND2_X1 U14974 ( .A1(n12744), .A2(n12943), .ZN(n12745) );
  OR2_X1 U14975 ( .A1(n12745), .A2(n12752), .ZN(n13896) );
  INV_X1 U14976 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n13895) );
  NAND2_X1 U14977 ( .A1(n13169), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n12747) );
  NAND2_X1 U14978 ( .A1(n13168), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n12746) );
  OAI211_X1 U14979 ( .C1(n13895), .C2(n13172), .A(n12747), .B(n12746), .ZN(
        n12748) );
  INV_X1 U14980 ( .A(n12748), .ZN(n12749) );
  OAI21_X1 U14981 ( .B1(n13896), .B2(n12901), .A(n12749), .ZN(n13907) );
  NAND2_X1 U14982 ( .A1(n13907), .A2(n6611), .ZN(n12750) );
  NAND2_X1 U14983 ( .A1(n12751), .A2(n12750), .ZN(n12939) );
  NOR2_X1 U14984 ( .A1(n12751), .A2(n12750), .ZN(n12938) );
  OR2_X1 U14985 ( .A1(n12752), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n12753) );
  AND2_X1 U14986 ( .A1(n12753), .A2(n12771), .ZN(n13881) );
  NAND2_X1 U14987 ( .A1(n13881), .A2(n12754), .ZN(n12759) );
  INV_X1 U14988 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n13659) );
  NAND2_X1 U14989 ( .A1(n12900), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n12756) );
  NAND2_X1 U14990 ( .A1(n13168), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n12755) );
  OAI211_X1 U14991 ( .C1(n12845), .C2(n13659), .A(n12756), .B(n12755), .ZN(
        n12757) );
  INV_X1 U14992 ( .A(n12757), .ZN(n12758) );
  NAND2_X1 U14993 ( .A1(n12759), .A2(n12758), .ZN(n13365) );
  NAND2_X1 U14994 ( .A1(n13365), .A2(n12855), .ZN(n12764) );
  NAND2_X1 U14995 ( .A1(n12760), .A2(n10117), .ZN(n12762) );
  NAND2_X1 U14996 ( .A1(n12892), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n12761) );
  XNOR2_X1 U14997 ( .A(n14016), .B(n12895), .ZN(n12763) );
  XOR2_X1 U14998 ( .A(n12764), .B(n12763), .Z(n12913) );
  INV_X1 U14999 ( .A(n12763), .ZN(n12765) );
  NAND2_X1 U15000 ( .A1(n12766), .A2(n10117), .ZN(n12768) );
  NAND2_X1 U15001 ( .A1(n12892), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n12767) );
  XNOR2_X1 U15002 ( .A(n14010), .B(n12895), .ZN(n12780) );
  NAND2_X1 U15003 ( .A1(n12900), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n12779) );
  INV_X1 U15004 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n12770) );
  OR2_X1 U15005 ( .A1(n12845), .A2(n12770), .ZN(n12778) );
  INV_X1 U15006 ( .A(n12771), .ZN(n12773) );
  INV_X1 U15007 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n12952) );
  INV_X1 U15008 ( .A(n12787), .ZN(n12772) );
  OAI21_X1 U15009 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(n12773), .A(n12772), 
        .ZN(n13862) );
  OR2_X1 U15010 ( .A1(n12901), .A2(n13862), .ZN(n12777) );
  INV_X1 U15011 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n12774) );
  OR2_X1 U15012 ( .A1(n12775), .A2(n12774), .ZN(n12776) );
  NAND4_X1 U15013 ( .A1(n12779), .A2(n12778), .A3(n12777), .A4(n12776), .ZN(
        n13875) );
  NOR2_X1 U15014 ( .A1(n13207), .A2(n15065), .ZN(n12948) );
  AOI21_X2 U15015 ( .B1(n12949), .B2(n12948), .A(n12782), .ZN(n12794) );
  NAND2_X1 U15016 ( .A1(n12783), .A2(n10117), .ZN(n12785) );
  NAND2_X1 U15017 ( .A1(n12892), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n12784) );
  XNOR2_X1 U15018 ( .A(n14004), .B(n12895), .ZN(n12793) );
  NAND2_X1 U15019 ( .A1(n12900), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n12792) );
  INV_X1 U15020 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n12786) );
  OR2_X1 U15021 ( .A1(n12845), .A2(n12786), .ZN(n12791) );
  NAND2_X1 U15022 ( .A1(n12787), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n12800) );
  OAI21_X1 U15023 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(n12787), .A(n12800), 
        .ZN(n13845) );
  OR2_X1 U15024 ( .A1(n12901), .A2(n13845), .ZN(n12790) );
  INV_X1 U15025 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n12788) );
  OR2_X1 U15026 ( .A1(n12903), .A2(n12788), .ZN(n12789) );
  NAND4_X1 U15027 ( .A1(n12792), .A2(n12791), .A3(n12790), .A4(n12789), .ZN(
        n13368) );
  INV_X1 U15028 ( .A(n13368), .ZN(n13367) );
  NOR2_X1 U15029 ( .A1(n13367), .A2(n11374), .ZN(n12873) );
  NAND2_X1 U15030 ( .A1(n12796), .A2(n10117), .ZN(n12798) );
  NAND2_X1 U15031 ( .A1(n12892), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n12797) );
  XNOR2_X1 U15032 ( .A(n13999), .B(n12895), .ZN(n12809) );
  NAND2_X1 U15033 ( .A1(n13169), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n12806) );
  INV_X1 U15034 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n12799) );
  OR2_X1 U15035 ( .A1(n13172), .A2(n12799), .ZN(n12805) );
  OAI21_X1 U15036 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(n12801), .A(n12817), 
        .ZN(n13830) );
  OR2_X1 U15037 ( .A1(n12901), .A2(n13830), .ZN(n12804) );
  INV_X1 U15038 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n12802) );
  OR2_X1 U15039 ( .A1(n12903), .A2(n12802), .ZN(n12803) );
  NAND4_X1 U15040 ( .A1(n12806), .A2(n12805), .A3(n12804), .A4(n12803), .ZN(
        n13260) );
  NAND2_X1 U15041 ( .A1(n13260), .A2(n12855), .ZN(n12807) );
  XNOR2_X1 U15042 ( .A(n12809), .B(n12807), .ZN(n12929) );
  INV_X1 U15043 ( .A(n12807), .ZN(n12808) );
  NAND2_X1 U15044 ( .A1(n12809), .A2(n12808), .ZN(n12810) );
  NAND2_X1 U15045 ( .A1(n12811), .A2(n10117), .ZN(n12813) );
  NAND2_X1 U15046 ( .A1(n12892), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n12812) );
  XNOR2_X1 U15047 ( .A(n13995), .B(n12895), .ZN(n12826) );
  NAND2_X1 U15048 ( .A1(n12900), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n12823) );
  INV_X1 U15049 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n12814) );
  OR2_X1 U15050 ( .A1(n12845), .A2(n12814), .ZN(n12822) );
  INV_X1 U15051 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n12816) );
  NAND2_X1 U15052 ( .A1(n12817), .A2(n12816), .ZN(n12818) );
  NAND2_X1 U15053 ( .A1(n12834), .A2(n12818), .ZN(n13815) );
  INV_X1 U15054 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n12819) );
  OR2_X1 U15055 ( .A1(n12903), .A2(n12819), .ZN(n12820) );
  NAND4_X1 U15056 ( .A1(n12823), .A2(n12822), .A3(n12821), .A4(n12820), .ZN(
        n13372) );
  NAND2_X1 U15057 ( .A1(n13372), .A2(n6611), .ZN(n12824) );
  XNOR2_X1 U15058 ( .A(n12826), .B(n12824), .ZN(n12921) );
  INV_X1 U15059 ( .A(n12824), .ZN(n12825) );
  NAND2_X1 U15060 ( .A1(n12826), .A2(n12825), .ZN(n12827) );
  NAND2_X1 U15061 ( .A1(n12829), .A2(n10117), .ZN(n12831) );
  NAND2_X1 U15062 ( .A1(n12892), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n12830) );
  XNOR2_X1 U15063 ( .A(n13990), .B(n11155), .ZN(n12842) );
  NAND2_X1 U15064 ( .A1(n12900), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n12840) );
  INV_X1 U15065 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n12832) );
  OR2_X1 U15066 ( .A1(n12845), .A2(n12832), .ZN(n12839) );
  INV_X1 U15067 ( .A(n12834), .ZN(n12833) );
  NAND2_X1 U15068 ( .A1(n12833), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n12848) );
  INV_X1 U15069 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n12961) );
  NAND2_X1 U15070 ( .A1(n12834), .A2(n12961), .ZN(n12835) );
  NAND2_X1 U15071 ( .A1(n12848), .A2(n12835), .ZN(n13796) );
  INV_X1 U15072 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n12836) );
  OR2_X1 U15073 ( .A1(n12903), .A2(n12836), .ZN(n12837) );
  NAND4_X1 U15074 ( .A1(n12840), .A2(n12839), .A3(n12838), .A4(n12837), .ZN(
        n13354) );
  NAND2_X1 U15075 ( .A1(n13354), .A2(n12855), .ZN(n12841) );
  NAND2_X1 U15076 ( .A1(n12842), .A2(n12841), .ZN(n12843) );
  OAI21_X1 U15077 ( .B1(n12842), .B2(n12841), .A(n12843), .ZN(n12960) );
  NAND2_X1 U15078 ( .A1(n12900), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n12854) );
  INV_X1 U15079 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n12844) );
  OR2_X1 U15080 ( .A1(n12845), .A2(n12844), .ZN(n12853) );
  INV_X1 U15081 ( .A(n12848), .ZN(n12846) );
  NAND2_X1 U15082 ( .A1(n12846), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n12861) );
  INV_X1 U15083 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n12847) );
  NAND2_X1 U15084 ( .A1(n12848), .A2(n12847), .ZN(n12849) );
  NAND2_X1 U15085 ( .A1(n12861), .A2(n12849), .ZN(n13405) );
  INV_X1 U15086 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n12850) );
  OR2_X1 U15087 ( .A1(n12903), .A2(n12850), .ZN(n12851) );
  NAND4_X1 U15088 ( .A1(n12854), .A2(n12853), .A3(n12852), .A4(n12851), .ZN(
        n13356) );
  NAND2_X1 U15089 ( .A1(n13356), .A2(n12855), .ZN(n12887) );
  NAND2_X1 U15090 ( .A1(n12856), .A2(n10117), .ZN(n12858) );
  NAND2_X1 U15091 ( .A1(n12892), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n12857) );
  XNOR2_X1 U15092 ( .A(n13985), .B(n12895), .ZN(n12886) );
  XOR2_X1 U15093 ( .A(n12887), .B(n12886), .Z(n12889) );
  XNOR2_X1 U15094 ( .A(n12890), .B(n12889), .ZN(n12871) );
  NAND2_X1 U15095 ( .A1(n13169), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n12867) );
  INV_X1 U15096 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13396) );
  OR2_X1 U15097 ( .A1(n13172), .A2(n13396), .ZN(n12866) );
  INV_X1 U15098 ( .A(n12861), .ZN(n12859) );
  NAND2_X1 U15099 ( .A1(n12859), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n13383) );
  INV_X1 U15100 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n12860) );
  NAND2_X1 U15101 ( .A1(n12861), .A2(n12860), .ZN(n12862) );
  NAND2_X1 U15102 ( .A1(n13383), .A2(n12862), .ZN(n13395) );
  OR2_X1 U15103 ( .A1(n12901), .A2(n13395), .ZN(n12865) );
  INV_X1 U15104 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n12863) );
  OR2_X1 U15105 ( .A1(n12903), .A2(n12863), .ZN(n12864) );
  OAI22_X1 U15106 ( .A1(n13373), .A2(n13928), .B1(n13358), .B2(n14784), .ZN(
        n13413) );
  AOI22_X1 U15107 ( .A1(n13413), .A2(n14795), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12868) );
  OAI21_X1 U15108 ( .B1(n13405), .B2(n14799), .A(n12868), .ZN(n12869) );
  AOI21_X1 U15109 ( .B1(n13985), .B2(n14796), .A(n12869), .ZN(n12870) );
  OAI21_X1 U15110 ( .B1(n12871), .B2(n12967), .A(n12870), .ZN(P2_U3186) );
  XNOR2_X1 U15111 ( .A(n12872), .B(n12873), .ZN(n12877) );
  INV_X1 U15112 ( .A(n13260), .ZN(n13370) );
  OAI22_X1 U15113 ( .A1(n13207), .A2(n13928), .B1(n13370), .B2(n14784), .ZN(
        n13843) );
  AOI22_X1 U15114 ( .A1(n13843), .A2(n14795), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12874) );
  OAI21_X1 U15115 ( .B1(n13845), .B2(n14799), .A(n12874), .ZN(n12875) );
  AOI21_X1 U15116 ( .B1(n14004), .B2(n14796), .A(n12875), .ZN(n12876) );
  OAI21_X1 U15117 ( .B1(n12877), .B2(n12967), .A(n12876), .ZN(P2_U3188) );
  NOR2_X1 U15118 ( .A1(n12879), .A2(n12736), .ZN(n12880) );
  XNOR2_X1 U15119 ( .A(n12881), .B(n12880), .ZN(n12885) );
  NAND2_X1 U15120 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13334)
         );
  OAI21_X1 U15121 ( .B1(n13912), .B2(n14799), .A(n13334), .ZN(n12883) );
  INV_X1 U15122 ( .A(n13907), .ZN(n13352) );
  OAI22_X1 U15123 ( .A1(n13352), .A2(n12962), .B1(n13363), .B2(n12963), .ZN(
        n12882) );
  AOI211_X1 U15124 ( .C1(n14027), .C2(n14796), .A(n12883), .B(n12882), .ZN(
        n12884) );
  OAI21_X1 U15125 ( .B1(n12885), .B2(n12967), .A(n12884), .ZN(P2_U3191) );
  INV_X1 U15126 ( .A(n12886), .ZN(n12888) );
  NAND2_X1 U15127 ( .A1(n12891), .A2(n10117), .ZN(n12894) );
  NAND2_X1 U15128 ( .A1(n12892), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n12893) );
  NOR2_X1 U15129 ( .A1(n13358), .A2(n15065), .ZN(n12896) );
  XNOR2_X1 U15130 ( .A(n12896), .B(n12895), .ZN(n12897) );
  XNOR2_X1 U15131 ( .A(n13394), .B(n12897), .ZN(n12898) );
  XNOR2_X1 U15132 ( .A(n12899), .B(n12898), .ZN(n12912) );
  NAND2_X1 U15133 ( .A1(n12900), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n12907) );
  NAND2_X1 U15134 ( .A1(n13169), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n12906) );
  OR2_X1 U15135 ( .A1(n12901), .A2(n13383), .ZN(n12905) );
  INV_X1 U15136 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n12902) );
  OR2_X1 U15137 ( .A1(n12903), .A2(n12902), .ZN(n12904) );
  NAND4_X1 U15138 ( .A1(n12907), .A2(n12906), .A3(n12905), .A4(n12904), .ZN(
        n13259) );
  INV_X1 U15139 ( .A(n13259), .ZN(n12908) );
  OAI22_X1 U15140 ( .A1(n12908), .A2(n14784), .B1(n13790), .B2(n13928), .ZN(
        n13391) );
  AOI22_X1 U15141 ( .A1(n13391), .A2(n14795), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12909) );
  OAI21_X1 U15142 ( .B1(n13395), .B2(n14799), .A(n12909), .ZN(n12910) );
  AOI21_X1 U15143 ( .B1(n13980), .B2(n14796), .A(n12910), .ZN(n12911) );
  OAI21_X1 U15144 ( .B1(n12912), .B2(n12967), .A(n12911), .ZN(P2_U3192) );
  XNOR2_X1 U15145 ( .A(n12914), .B(n12913), .ZN(n12920) );
  INV_X1 U15146 ( .A(n13881), .ZN(n12916) );
  INV_X1 U15147 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n12915) );
  OAI22_X1 U15148 ( .A1(n12916), .A2(n14799), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12915), .ZN(n12918) );
  OAI22_X1 U15149 ( .A1(n13352), .A2(n12963), .B1(n13207), .B2(n12962), .ZN(
        n12917) );
  AOI211_X1 U15150 ( .C1(n14016), .C2(n14796), .A(n12918), .B(n12917), .ZN(
        n12919) );
  OAI21_X1 U15151 ( .B1(n12920), .B2(n12967), .A(n12919), .ZN(P2_U3195) );
  XNOR2_X1 U15152 ( .A(n12922), .B(n12921), .ZN(n12928) );
  NAND2_X1 U15153 ( .A1(n14787), .A2(n13260), .ZN(n12924) );
  NAND2_X1 U15154 ( .A1(n13949), .A2(n13354), .ZN(n12923) );
  NAND2_X1 U15155 ( .A1(n12924), .A2(n12923), .ZN(n13808) );
  AOI22_X1 U15156 ( .A1(n14795), .A2(n13808), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12925) );
  OAI21_X1 U15157 ( .B1(n13815), .B2(n14799), .A(n12925), .ZN(n12926) );
  AOI21_X1 U15158 ( .B1(n13995), .B2(n14796), .A(n12926), .ZN(n12927) );
  OAI21_X1 U15159 ( .B1(n12928), .B2(n12967), .A(n12927), .ZN(P2_U3197) );
  XNOR2_X1 U15160 ( .A(n12930), .B(n12929), .ZN(n12936) );
  NAND2_X1 U15161 ( .A1(n14787), .A2(n13368), .ZN(n12932) );
  NAND2_X1 U15162 ( .A1(n13949), .A2(n13372), .ZN(n12931) );
  NAND2_X1 U15163 ( .A1(n12932), .A2(n12931), .ZN(n13825) );
  AOI22_X1 U15164 ( .A1(n14795), .A2(n13825), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12933) );
  OAI21_X1 U15165 ( .B1(n13830), .B2(n14799), .A(n12933), .ZN(n12934) );
  AOI21_X1 U15166 ( .B1(n13999), .B2(n14796), .A(n12934), .ZN(n12935) );
  OAI21_X1 U15167 ( .B1(n12936), .B2(n12967), .A(n12935), .ZN(P2_U3201) );
  INV_X1 U15168 ( .A(n12937), .ZN(n12942) );
  INV_X1 U15169 ( .A(n12938), .ZN(n12940) );
  NAND2_X1 U15170 ( .A1(n12940), .A2(n12939), .ZN(n12941) );
  XNOR2_X1 U15171 ( .A(n12942), .B(n12941), .ZN(n12947) );
  OAI22_X1 U15172 ( .A1(n13896), .A2(n14799), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12943), .ZN(n12945) );
  INV_X1 U15173 ( .A(n13365), .ZN(n13891) );
  OAI22_X1 U15174 ( .A1(n13891), .A2(n12962), .B1(n13929), .B2(n12963), .ZN(
        n12944) );
  AOI211_X1 U15175 ( .C1(n14022), .C2(n14796), .A(n12945), .B(n12944), .ZN(
        n12946) );
  OAI21_X1 U15176 ( .B1(n12947), .B2(n12967), .A(n12946), .ZN(P2_U3205) );
  XNOR2_X1 U15177 ( .A(n12949), .B(n12948), .ZN(n12956) );
  AND2_X1 U15178 ( .A1(n13949), .A2(n13368), .ZN(n12950) );
  AOI21_X1 U15179 ( .B1(n13365), .B2(n14787), .A(n12950), .ZN(n13856) );
  NOR2_X1 U15180 ( .A1(n13856), .A2(n12951), .ZN(n12954) );
  OAI22_X1 U15181 ( .A1(n14799), .A2(n13862), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12952), .ZN(n12953) );
  AOI211_X1 U15182 ( .C1(n14010), .C2(n14796), .A(n12954), .B(n12953), .ZN(
        n12955) );
  OAI21_X1 U15183 ( .B1(n12956), .B2(n12967), .A(n12955), .ZN(P2_U3207) );
  INV_X1 U15184 ( .A(n12957), .ZN(n12958) );
  AOI21_X1 U15185 ( .B1(n12960), .B2(n12959), .A(n12958), .ZN(n12968) );
  OAI22_X1 U15186 ( .A1(n14799), .A2(n13796), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12961), .ZN(n12965) );
  INV_X1 U15187 ( .A(n13372), .ZN(n13791) );
  OAI22_X1 U15188 ( .A1(n13791), .A2(n12963), .B1(n12962), .B2(n13790), .ZN(
        n12964) );
  AOI211_X1 U15189 ( .C1(n13990), .C2(n14796), .A(n12965), .B(n12964), .ZN(
        n12966) );
  OAI21_X1 U15190 ( .B1(n12968), .B2(n12967), .A(n12966), .ZN(P2_U3212) );
  NAND2_X1 U15191 ( .A1(n12970), .A2(n13000), .ZN(n12972) );
  NAND2_X1 U15192 ( .A1(n12972), .A2(n12971), .ZN(n12975) );
  INV_X2 U15193 ( .A(n13000), .ZN(n13228) );
  NAND2_X1 U15194 ( .A1(n13173), .A2(n12973), .ZN(n12974) );
  NAND2_X1 U15195 ( .A1(n12975), .A2(n12974), .ZN(n12978) );
  OAI211_X1 U15196 ( .C1(n12976), .C2(n13224), .A(n10172), .B(n13228), .ZN(
        n12977) );
  NAND2_X1 U15197 ( .A1(n12978), .A2(n12977), .ZN(n12982) );
  MUX2_X1 U15198 ( .A(n10324), .B(n9993), .S(n6685), .Z(n12981) );
  MUX2_X1 U15199 ( .A(n12979), .B(n13275), .S(n13228), .Z(n12980) );
  NAND2_X1 U15200 ( .A1(n12982), .A2(n12981), .ZN(n12983) );
  MUX2_X1 U15201 ( .A(n10317), .B(n10319), .S(n6685), .Z(n12986) );
  MUX2_X1 U15202 ( .A(n10319), .B(n10317), .S(n13173), .Z(n12985) );
  INV_X1 U15203 ( .A(n12986), .ZN(n12987) );
  MUX2_X1 U15204 ( .A(n13948), .B(n12988), .S(n13228), .Z(n12992) );
  NAND2_X1 U15205 ( .A1(n12991), .A2(n12992), .ZN(n12990) );
  MUX2_X1 U15206 ( .A(n12988), .B(n13948), .S(n13228), .Z(n12989) );
  NAND2_X1 U15207 ( .A1(n12990), .A2(n12989), .ZN(n12996) );
  INV_X1 U15208 ( .A(n12991), .ZN(n12994) );
  INV_X1 U15209 ( .A(n12992), .ZN(n12993) );
  MUX2_X1 U15210 ( .A(n15106), .B(n13274), .S(n13228), .Z(n12998) );
  MUX2_X1 U15211 ( .A(n13274), .B(n15106), .S(n13228), .Z(n12997) );
  INV_X1 U15212 ( .A(n12998), .ZN(n12999) );
  MUX2_X1 U15213 ( .A(n13950), .B(n15113), .S(n13228), .Z(n13004) );
  NAND2_X1 U15214 ( .A1(n13003), .A2(n13004), .ZN(n13002) );
  MUX2_X1 U15215 ( .A(n13950), .B(n15113), .S(n6616), .Z(n13001) );
  NAND2_X1 U15216 ( .A1(n13002), .A2(n13001), .ZN(n13008) );
  INV_X1 U15217 ( .A(n13003), .ZN(n13006) );
  INV_X1 U15218 ( .A(n13004), .ZN(n13005) );
  MUX2_X1 U15219 ( .A(n13272), .B(n13009), .S(n6616), .Z(n13011) );
  MUX2_X1 U15220 ( .A(n13272), .B(n13009), .S(n13228), .Z(n13010) );
  INV_X1 U15221 ( .A(n13011), .ZN(n13012) );
  MUX2_X1 U15222 ( .A(n13271), .B(n13013), .S(n13173), .Z(n13017) );
  NAND2_X1 U15223 ( .A1(n13016), .A2(n13017), .ZN(n13015) );
  MUX2_X1 U15224 ( .A(n13271), .B(n13013), .S(n6616), .Z(n13014) );
  NAND2_X1 U15225 ( .A1(n13015), .A2(n13014), .ZN(n13021) );
  INV_X1 U15226 ( .A(n13016), .ZN(n13019) );
  INV_X1 U15227 ( .A(n13017), .ZN(n13018) );
  NAND2_X1 U15228 ( .A1(n13019), .A2(n13018), .ZN(n13020) );
  NAND2_X1 U15229 ( .A1(n13021), .A2(n13020), .ZN(n13024) );
  MUX2_X1 U15230 ( .A(n13270), .B(n13022), .S(n6616), .Z(n13025) );
  MUX2_X1 U15231 ( .A(n13270), .B(n13022), .S(n13228), .Z(n13023) );
  INV_X1 U15232 ( .A(n13025), .ZN(n13026) );
  MUX2_X1 U15233 ( .A(n13269), .B(n13027), .S(n13228), .Z(n13031) );
  MUX2_X1 U15234 ( .A(n13269), .B(n13027), .S(n6616), .Z(n13028) );
  NAND2_X1 U15235 ( .A1(n13029), .A2(n13028), .ZN(n13035) );
  INV_X1 U15236 ( .A(n13030), .ZN(n13033) );
  INV_X1 U15237 ( .A(n13031), .ZN(n13032) );
  NAND2_X1 U15238 ( .A1(n13035), .A2(n13034), .ZN(n13037) );
  MUX2_X1 U15239 ( .A(n13268), .B(n15061), .S(n6616), .Z(n13038) );
  MUX2_X1 U15240 ( .A(n13268), .B(n15061), .S(n13228), .Z(n13036) );
  INV_X1 U15241 ( .A(n13038), .ZN(n13039) );
  MUX2_X1 U15242 ( .A(n13267), .B(n13040), .S(n13173), .Z(n13044) );
  MUX2_X1 U15243 ( .A(n13267), .B(n13040), .S(n6616), .Z(n13041) );
  NAND2_X1 U15244 ( .A1(n13042), .A2(n13041), .ZN(n13048) );
  INV_X1 U15245 ( .A(n13043), .ZN(n13046) );
  INV_X1 U15246 ( .A(n13044), .ZN(n13045) );
  NAND2_X1 U15247 ( .A1(n13046), .A2(n13045), .ZN(n13047) );
  MUX2_X1 U15248 ( .A(n13266), .B(n14830), .S(n6616), .Z(n13050) );
  MUX2_X1 U15249 ( .A(n13266), .B(n14830), .S(n13228), .Z(n13049) );
  INV_X1 U15250 ( .A(n13050), .ZN(n13051) );
  MUX2_X1 U15251 ( .A(n14786), .B(n13052), .S(n13228), .Z(n13056) );
  NAND2_X1 U15252 ( .A1(n13055), .A2(n13056), .ZN(n13054) );
  MUX2_X1 U15253 ( .A(n14786), .B(n13052), .S(n6616), .Z(n13053) );
  NAND2_X1 U15254 ( .A1(n13054), .A2(n13053), .ZN(n13060) );
  INV_X1 U15255 ( .A(n13055), .ZN(n13058) );
  INV_X1 U15256 ( .A(n13056), .ZN(n13057) );
  NAND2_X1 U15257 ( .A1(n13058), .A2(n13057), .ZN(n13059) );
  NAND2_X1 U15258 ( .A1(n13060), .A2(n13059), .ZN(n13096) );
  MUX2_X1 U15259 ( .A(n13263), .B(n14042), .S(n6616), .Z(n13074) );
  NAND2_X1 U15260 ( .A1(n13202), .A2(n13074), .ZN(n13063) );
  OR2_X1 U15261 ( .A1(n14037), .A2(n13927), .ZN(n13360) );
  NAND2_X1 U15262 ( .A1(n14037), .A2(n13927), .ZN(n13361) );
  AND2_X1 U15263 ( .A1(n13263), .A2(n6616), .ZN(n13061) );
  AOI21_X1 U15264 ( .B1(n14042), .B2(n13228), .A(n13061), .ZN(n13062) );
  NAND3_X1 U15265 ( .A1(n13360), .A2(n13361), .A3(n13062), .ZN(n13079) );
  NAND2_X1 U15266 ( .A1(n13063), .A2(n13079), .ZN(n13085) );
  MUX2_X1 U15267 ( .A(n14785), .B(n13064), .S(n6616), .Z(n13082) );
  MUX2_X1 U15268 ( .A(n13264), .B(n14048), .S(n13173), .Z(n13081) );
  NAND2_X1 U15269 ( .A1(n13082), .A2(n13081), .ZN(n13065) );
  NAND2_X1 U15270 ( .A1(n13085), .A2(n13065), .ZN(n13089) );
  MUX2_X1 U15271 ( .A(n13066), .B(n14816), .S(n6616), .Z(n13071) );
  MUX2_X1 U15272 ( .A(n13265), .B(n7081), .S(n13228), .Z(n13070) );
  AND2_X1 U15273 ( .A1(n13071), .A2(n13070), .ZN(n13067) );
  NOR2_X1 U15274 ( .A1(n13089), .A2(n13067), .ZN(n13095) );
  MUX2_X1 U15275 ( .A(n13906), .B(n14030), .S(n6616), .Z(n13069) );
  AND2_X1 U15276 ( .A1(n13095), .A2(n13069), .ZN(n13068) );
  NAND2_X1 U15277 ( .A1(n13096), .A2(n13068), .ZN(n13094) );
  INV_X1 U15278 ( .A(n13069), .ZN(n13098) );
  INV_X1 U15279 ( .A(n13070), .ZN(n13073) );
  INV_X1 U15280 ( .A(n13071), .ZN(n13072) );
  NAND2_X1 U15281 ( .A1(n13073), .A2(n13072), .ZN(n13088) );
  INV_X1 U15282 ( .A(n13074), .ZN(n13078) );
  AND2_X1 U15283 ( .A1(n13262), .A2(n13173), .ZN(n13076) );
  OAI21_X1 U15284 ( .B1(n13262), .B2(n6685), .A(n14037), .ZN(n13075) );
  OAI21_X1 U15285 ( .B1(n13076), .B2(n14037), .A(n13075), .ZN(n13077) );
  OAI21_X1 U15286 ( .B1(n13079), .B2(n13078), .A(n13077), .ZN(n13080) );
  INV_X1 U15287 ( .A(n13080), .ZN(n13087) );
  INV_X1 U15288 ( .A(n13081), .ZN(n13084) );
  INV_X1 U15289 ( .A(n13082), .ZN(n13083) );
  NAND3_X1 U15290 ( .A1(n13085), .A2(n13084), .A3(n13083), .ZN(n13086) );
  OAI211_X1 U15291 ( .C1(n13089), .C2(n13088), .A(n13087), .B(n13086), .ZN(
        n13090) );
  INV_X1 U15292 ( .A(n13090), .ZN(n13097) );
  OR2_X1 U15293 ( .A1(n13098), .A2(n13097), .ZN(n13092) );
  MUX2_X1 U15294 ( .A(n13906), .B(n14030), .S(n13173), .Z(n13091) );
  AND2_X1 U15295 ( .A1(n13092), .A2(n13091), .ZN(n13093) );
  NAND2_X1 U15296 ( .A1(n13094), .A2(n13093), .ZN(n13102) );
  NAND2_X1 U15297 ( .A1(n13096), .A2(n13095), .ZN(n13100) );
  AND2_X1 U15298 ( .A1(n13098), .A2(n13097), .ZN(n13099) );
  NAND2_X1 U15299 ( .A1(n13100), .A2(n13099), .ZN(n13101) );
  MUX2_X1 U15300 ( .A(n13261), .B(n14027), .S(n6685), .Z(n13104) );
  MUX2_X1 U15301 ( .A(n13261), .B(n14027), .S(n6616), .Z(n13103) );
  MUX2_X1 U15302 ( .A(n13907), .B(n14022), .S(n6616), .Z(n13108) );
  NAND2_X1 U15303 ( .A1(n13107), .A2(n13108), .ZN(n13106) );
  MUX2_X1 U15304 ( .A(n13907), .B(n14022), .S(n13173), .Z(n13105) );
  NAND2_X1 U15305 ( .A1(n13106), .A2(n13105), .ZN(n13112) );
  INV_X1 U15306 ( .A(n13107), .ZN(n13110) );
  INV_X1 U15307 ( .A(n13108), .ZN(n13109) );
  NAND2_X1 U15308 ( .A1(n13110), .A2(n13109), .ZN(n13111) );
  NAND2_X1 U15309 ( .A1(n13112), .A2(n13111), .ZN(n13114) );
  MUX2_X1 U15310 ( .A(n13365), .B(n14016), .S(n13228), .Z(n13115) );
  MUX2_X1 U15311 ( .A(n13365), .B(n14016), .S(n6616), .Z(n13113) );
  INV_X1 U15312 ( .A(n13115), .ZN(n13116) );
  MUX2_X1 U15313 ( .A(n13875), .B(n14010), .S(n6616), .Z(n13119) );
  MUX2_X1 U15314 ( .A(n13875), .B(n14010), .S(n13228), .Z(n13117) );
  NAND2_X1 U15315 ( .A1(n13118), .A2(n13117), .ZN(n13125) );
  OR2_X2 U15316 ( .A1(n13120), .A2(n13119), .ZN(n13124) );
  NAND2_X1 U15317 ( .A1(n13125), .A2(n13124), .ZN(n13121) );
  MUX2_X1 U15318 ( .A(n13368), .B(n14004), .S(n13228), .Z(n13126) );
  NAND2_X1 U15319 ( .A1(n13121), .A2(n13126), .ZN(n13123) );
  MUX2_X1 U15320 ( .A(n13368), .B(n14004), .S(n6616), .Z(n13122) );
  NAND2_X1 U15321 ( .A1(n13123), .A2(n13122), .ZN(n13130) );
  AND2_X1 U15322 ( .A1(n13125), .A2(n13124), .ZN(n13128) );
  INV_X1 U15323 ( .A(n13126), .ZN(n13127) );
  NAND2_X1 U15324 ( .A1(n13128), .A2(n13127), .ZN(n13129) );
  MUX2_X1 U15325 ( .A(n13260), .B(n13999), .S(n6616), .Z(n13132) );
  MUX2_X1 U15326 ( .A(n13260), .B(n13999), .S(n6685), .Z(n13131) );
  MUX2_X1 U15327 ( .A(n13372), .B(n13995), .S(n6685), .Z(n13136) );
  NAND2_X1 U15328 ( .A1(n13135), .A2(n13136), .ZN(n13134) );
  MUX2_X1 U15329 ( .A(n13372), .B(n13995), .S(n6616), .Z(n13133) );
  NAND2_X1 U15330 ( .A1(n13134), .A2(n13133), .ZN(n13140) );
  INV_X1 U15331 ( .A(n13135), .ZN(n13138) );
  INV_X1 U15332 ( .A(n13136), .ZN(n13137) );
  NAND2_X1 U15333 ( .A1(n13138), .A2(n13137), .ZN(n13139) );
  NAND2_X1 U15334 ( .A1(n13140), .A2(n13139), .ZN(n13143) );
  MUX2_X1 U15335 ( .A(n13354), .B(n13990), .S(n6616), .Z(n13142) );
  MUX2_X1 U15336 ( .A(n13354), .B(n13990), .S(n13173), .Z(n13141) );
  MUX2_X1 U15337 ( .A(n13356), .B(n13985), .S(n13228), .Z(n13147) );
  MUX2_X1 U15338 ( .A(n13356), .B(n13985), .S(n6616), .Z(n13144) );
  NAND2_X1 U15339 ( .A1(n13145), .A2(n13144), .ZN(n13151) );
  INV_X1 U15340 ( .A(n13146), .ZN(n13149) );
  INV_X1 U15341 ( .A(n13147), .ZN(n13148) );
  NAND2_X1 U15342 ( .A1(n13149), .A2(n13148), .ZN(n13150) );
  MUX2_X1 U15343 ( .A(n13358), .B(n13394), .S(n6616), .Z(n13155) );
  INV_X1 U15344 ( .A(n13155), .ZN(n13153) );
  MUX2_X1 U15345 ( .A(n13358), .B(n13394), .S(n13173), .Z(n13152) );
  INV_X1 U15346 ( .A(n13236), .ZN(n13220) );
  INV_X1 U15347 ( .A(n13154), .ZN(n13156) );
  NAND2_X1 U15348 ( .A1(n13156), .A2(n13155), .ZN(n13238) );
  NAND2_X1 U15349 ( .A1(n13157), .A2(n10117), .ZN(n13159) );
  NAND2_X1 U15350 ( .A1(n12892), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13158) );
  MUX2_X1 U15351 ( .A(n13259), .B(n13380), .S(n6616), .Z(n13160) );
  INV_X1 U15352 ( .A(n13160), .ZN(n13230) );
  MUX2_X1 U15353 ( .A(n13380), .B(n13259), .S(n6616), .Z(n13229) );
  INV_X1 U15354 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n13538) );
  NAND2_X1 U15355 ( .A1(n13168), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n13163) );
  NAND2_X1 U15356 ( .A1(n13169), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n13162) );
  OAI211_X1 U15357 ( .C1(n13172), .C2(n13538), .A(n13163), .B(n13162), .ZN(
        n13377) );
  NAND2_X1 U15358 ( .A1(n12892), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13166) );
  MUX2_X1 U15359 ( .A(n13377), .B(n13343), .S(n13173), .Z(n13232) );
  INV_X1 U15360 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n13338) );
  NAND2_X1 U15361 ( .A1(n13168), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n13171) );
  NAND2_X1 U15362 ( .A1(n13169), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n13170) );
  OAI211_X1 U15363 ( .C1(n13172), .C2(n13338), .A(n13171), .B(n13170), .ZN(
        n13340) );
  NAND2_X1 U15364 ( .A1(n13340), .A2(n13228), .ZN(n13175) );
  NAND2_X1 U15365 ( .A1(n13254), .A2(n13174), .ZN(n13217) );
  NAND4_X1 U15366 ( .A1(n6610), .A2(n13175), .A3(n13252), .A4(n13217), .ZN(
        n13176) );
  AND2_X1 U15367 ( .A1(n13176), .A2(n13377), .ZN(n13177) );
  AOI21_X1 U15368 ( .B1(n13343), .B2(n6616), .A(n13177), .ZN(n13231) );
  AND2_X1 U15369 ( .A1(n13232), .A2(n13231), .ZN(n13240) );
  NAND2_X1 U15370 ( .A1(n14068), .A2(n10117), .ZN(n13179) );
  NAND2_X1 U15371 ( .A1(n12892), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n13178) );
  INV_X1 U15372 ( .A(n13340), .ZN(n13180) );
  NAND2_X1 U15373 ( .A1(n13966), .A2(n13180), .ZN(n13239) );
  AOI211_X1 U15374 ( .C1(n13230), .C2(n13229), .A(n13240), .B(n13221), .ZN(
        n13237) );
  NAND2_X1 U15375 ( .A1(n13980), .A2(n13358), .ZN(n13181) );
  NAND2_X1 U15376 ( .A1(n13985), .A2(n13790), .ZN(n13390) );
  XNOR2_X1 U15377 ( .A(n13995), .B(n13372), .ZN(n13353) );
  XNOR2_X1 U15378 ( .A(n14016), .B(n13365), .ZN(n13878) );
  XNOR2_X1 U15379 ( .A(n14030), .B(n13363), .ZN(n13923) );
  NAND4_X1 U15380 ( .A1(n13185), .A2(n15086), .A3(n13184), .A4(n13183), .ZN(
        n13187) );
  NOR2_X1 U15381 ( .A1(n13187), .A2(n13186), .ZN(n13189) );
  NAND4_X1 U15382 ( .A1(n13190), .A2(n13189), .A3(n13188), .A4(n13961), .ZN(
        n13193) );
  OR4_X1 U15383 ( .A1(n13194), .A2(n13193), .A3(n13192), .A4(n13191), .ZN(
        n13195) );
  NOR2_X1 U15384 ( .A1(n13196), .A2(n13195), .ZN(n13198) );
  NAND4_X1 U15385 ( .A1(n13199), .A2(n13198), .A3(n13197), .A4(n15062), .ZN(
        n13200) );
  NOR2_X1 U15386 ( .A1(n13201), .A2(n13200), .ZN(n13203) );
  NAND4_X1 U15387 ( .A1(n13204), .A2(n13203), .A3(n13202), .A4(n14800), .ZN(
        n13205) );
  NOR2_X1 U15388 ( .A1(n13923), .A2(n13205), .ZN(n13206) );
  XNOR2_X1 U15389 ( .A(n14022), .B(n13907), .ZN(n13351) );
  XNOR2_X1 U15390 ( .A(n14027), .B(n13261), .ZN(n13904) );
  NAND4_X1 U15391 ( .A1(n13878), .A2(n13206), .A3(n13351), .A4(n13904), .ZN(
        n13208) );
  NOR2_X1 U15392 ( .A1(n13208), .A2(n13867), .ZN(n13209) );
  XNOR2_X1 U15393 ( .A(n14004), .B(n13368), .ZN(n13841) );
  NAND4_X1 U15394 ( .A1(n13353), .A2(n13209), .A3(n13823), .A4(n13841), .ZN(
        n13210) );
  OR3_X1 U15395 ( .A1(n13409), .A2(n13801), .A3(n13210), .ZN(n13211) );
  NOR2_X1 U15396 ( .A1(n13357), .A2(n13211), .ZN(n13212) );
  AND2_X1 U15397 ( .A1(n13216), .A2(n13215), .ZN(n13227) );
  INV_X1 U15398 ( .A(n13227), .ZN(n13218) );
  NAND4_X1 U15399 ( .A1(n13220), .A2(n13238), .A3(n13237), .A4(n13247), .ZN(
        n13251) );
  AOI21_X1 U15400 ( .B1(n6610), .B2(n13331), .A(n13222), .ZN(n13223) );
  OAI21_X1 U15401 ( .B1(n13254), .B2(n13224), .A(n13223), .ZN(n13225) );
  INV_X1 U15402 ( .A(n13243), .ZN(n13235) );
  MUX2_X1 U15403 ( .A(n13239), .B(n13244), .S(n6685), .Z(n13234) );
  OAI22_X1 U15404 ( .A1(n13232), .A2(n13231), .B1(n13230), .B2(n13229), .ZN(
        n13233) );
  NAND4_X1 U15405 ( .A1(n13236), .A2(n13213), .A3(n13235), .A4(n13241), .ZN(
        n13250) );
  NAND3_X1 U15406 ( .A1(n13238), .A2(n13237), .A3(n13241), .ZN(n13249) );
  NOR2_X1 U15407 ( .A1(n13241), .A2(n13240), .ZN(n13245) );
  INV_X1 U15408 ( .A(n13245), .ZN(n13242) );
  NAND3_X1 U15409 ( .A1(n13243), .A2(n6728), .A3(n13242), .ZN(n13248) );
  INV_X1 U15410 ( .A(n13244), .ZN(n13246) );
  NOR4_X1 U15411 ( .A1(n13928), .A2(n15085), .A3(n13253), .A4(n13252), .ZN(
        n13256) );
  OAI21_X1 U15412 ( .B1(n13254), .B2(n13257), .A(P2_B_REG_SCAN_IN), .ZN(n13255) );
  OAI22_X1 U15413 ( .A1(n13258), .A2(n13257), .B1(n13256), .B2(n13255), .ZN(
        P2_U3328) );
  MUX2_X1 U15414 ( .A(n13340), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13273), .Z(
        P2_U3562) );
  MUX2_X1 U15415 ( .A(n13377), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13273), .Z(
        P2_U3561) );
  MUX2_X1 U15416 ( .A(n13259), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13273), .Z(
        P2_U3560) );
  INV_X1 U15417 ( .A(n13358), .ZN(n13376) );
  MUX2_X1 U15418 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13376), .S(P2_U3947), .Z(
        P2_U3559) );
  MUX2_X1 U15419 ( .A(n13356), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13273), .Z(
        P2_U3558) );
  MUX2_X1 U15420 ( .A(n13354), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13273), .Z(
        P2_U3557) );
  MUX2_X1 U15421 ( .A(n13372), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13273), .Z(
        P2_U3556) );
  MUX2_X1 U15422 ( .A(n13260), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13273), .Z(
        P2_U3555) );
  MUX2_X1 U15423 ( .A(n13368), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13273), .Z(
        P2_U3554) );
  MUX2_X1 U15424 ( .A(n13875), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13273), .Z(
        P2_U3553) );
  MUX2_X1 U15425 ( .A(n13365), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13273), .Z(
        P2_U3552) );
  MUX2_X1 U15426 ( .A(n13907), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13273), .Z(
        P2_U3551) );
  MUX2_X1 U15427 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13261), .S(P2_U3947), .Z(
        P2_U3550) );
  MUX2_X1 U15428 ( .A(n13906), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13273), .Z(
        P2_U3549) );
  MUX2_X1 U15429 ( .A(n13262), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13273), .Z(
        P2_U3548) );
  MUX2_X1 U15430 ( .A(n13263), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13273), .Z(
        P2_U3547) );
  MUX2_X1 U15431 ( .A(n13264), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13273), .Z(
        P2_U3546) );
  MUX2_X1 U15432 ( .A(n13265), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13273), .Z(
        P2_U3545) );
  MUX2_X1 U15433 ( .A(n14786), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13273), .Z(
        P2_U3544) );
  MUX2_X1 U15434 ( .A(n13266), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13273), .Z(
        P2_U3543) );
  MUX2_X1 U15435 ( .A(n13267), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13273), .Z(
        P2_U3542) );
  MUX2_X1 U15436 ( .A(n13268), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13273), .Z(
        P2_U3541) );
  MUX2_X1 U15437 ( .A(n13269), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13273), .Z(
        P2_U3540) );
  MUX2_X1 U15438 ( .A(n13270), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13273), .Z(
        P2_U3539) );
  MUX2_X1 U15439 ( .A(n13271), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13273), .Z(
        P2_U3538) );
  MUX2_X1 U15440 ( .A(n13272), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13273), .Z(
        P2_U3537) );
  MUX2_X1 U15441 ( .A(n13950), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13273), .Z(
        P2_U3536) );
  MUX2_X1 U15442 ( .A(n13274), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13273), .Z(
        P2_U3535) );
  MUX2_X1 U15443 ( .A(n13948), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13273), .Z(
        P2_U3534) );
  MUX2_X1 U15444 ( .A(n10319), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13273), .Z(
        P2_U3533) );
  MUX2_X1 U15445 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n13275), .S(P2_U3947), .Z(
        P2_U3532) );
  MUX2_X1 U15446 ( .A(n10525), .B(P2_REG2_REG_6__SCAN_IN), .S(n13276), .Z(
        n13277) );
  NAND3_X1 U15447 ( .A1(n13279), .A2(n13278), .A3(n13277), .ZN(n13280) );
  NAND2_X1 U15448 ( .A1(n13281), .A2(n13280), .ZN(n13282) );
  OAI22_X1 U15449 ( .A1(n13283), .A2(n15051), .B1(n15026), .B2(n13282), .ZN(
        n13284) );
  INV_X1 U15450 ( .A(n13284), .ZN(n13292) );
  INV_X1 U15451 ( .A(n13285), .ZN(n13286) );
  AOI21_X1 U15452 ( .B1(n15043), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n13286), .ZN(
        n13291) );
  OAI211_X1 U15453 ( .C1(n13289), .C2(n13288), .A(n14984), .B(n13287), .ZN(
        n13290) );
  NAND3_X1 U15454 ( .A1(n13292), .A2(n13291), .A3(n13290), .ZN(P2_U3220) );
  OAI211_X1 U15455 ( .C1(n13294), .C2(P2_REG2_REG_15__SCAN_IN), .A(n15045), 
        .B(n13293), .ZN(n13303) );
  AOI21_X1 U15456 ( .B1(n15032), .B2(n13296), .A(n13295), .ZN(n13302) );
  AOI211_X1 U15457 ( .C1(n13299), .C2(n13298), .A(n13297), .B(n15037), .ZN(
        n13300) );
  AOI21_X1 U15458 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(n15043), .A(n13300), 
        .ZN(n13301) );
  NAND3_X1 U15459 ( .A1(n13303), .A2(n13302), .A3(n13301), .ZN(P2_U3229) );
  AOI21_X1 U15460 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n13305), .A(n13304), 
        .ZN(n13323) );
  XNOR2_X1 U15461 ( .A(n13323), .B(n13322), .ZN(n13307) );
  NOR2_X1 U15462 ( .A1(n13306), .A2(n13307), .ZN(n13325) );
  AOI211_X1 U15463 ( .C1(n13307), .C2(n13306), .A(n13325), .B(n15037), .ZN(
        n13316) );
  OAI21_X1 U15464 ( .B1(n15051), .B2(n13322), .A(n13308), .ZN(n13315) );
  INV_X1 U15465 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n13313) );
  OAI21_X1 U15466 ( .B1(n11502), .B2(n13310), .A(n13309), .ZN(n13317) );
  XNOR2_X1 U15467 ( .A(n13317), .B(n13318), .ZN(n13311) );
  NOR2_X1 U15468 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n13311), .ZN(n13320) );
  AOI21_X1 U15469 ( .B1(n13311), .B2(P2_REG2_REG_18__SCAN_IN), .A(n13320), 
        .ZN(n13312) );
  OAI22_X1 U15470 ( .A1(n15035), .A2(n13313), .B1(n15026), .B2(n13312), .ZN(
        n13314) );
  OR3_X1 U15471 ( .A1(n13316), .A2(n13315), .A3(n13314), .ZN(P2_U3232) );
  NOR2_X1 U15472 ( .A1(n13318), .A2(n13317), .ZN(n13319) );
  NOR2_X1 U15473 ( .A1(n13320), .A2(n13319), .ZN(n13321) );
  XOR2_X1 U15474 ( .A(n13321), .B(n11875), .Z(n13329) );
  AOI21_X1 U15475 ( .B1(n13329), .B2(n15045), .A(n15032), .ZN(n13328) );
  NOR2_X1 U15476 ( .A1(n13323), .A2(n13322), .ZN(n13324) );
  NOR2_X1 U15477 ( .A1(n13325), .A2(n13324), .ZN(n13326) );
  XOR2_X1 U15478 ( .A(n13326), .B(P2_REG1_REG_19__SCAN_IN), .Z(n13330) );
  NAND2_X1 U15479 ( .A1(n13330), .A2(n14984), .ZN(n13327) );
  NAND2_X1 U15480 ( .A1(n13328), .A2(n13327), .ZN(n13333) );
  OAI22_X1 U15481 ( .A1(n13330), .A2(n15037), .B1(n13329), .B2(n15026), .ZN(
        n13332) );
  MUX2_X1 U15482 ( .A(n13333), .B(n13332), .S(n13331), .Z(n13336) );
  OAI21_X1 U15483 ( .B1(n15035), .B2(n7640), .A(n13334), .ZN(n13335) );
  INV_X1 U15484 ( .A(n14030), .ZN(n13931) );
  NAND2_X1 U15485 ( .A1(n13932), .A2(n13931), .ZN(n13930) );
  INV_X1 U15486 ( .A(n13999), .ZN(n13827) );
  NAND2_X1 U15487 ( .A1(n13829), .A2(n13819), .ZN(n13814) );
  NOR2_X2 U15488 ( .A1(n13794), .A2(n13985), .ZN(n13403) );
  XNOR2_X1 U15489 ( .A(n13966), .B(n13344), .ZN(n13337) );
  NAND2_X1 U15490 ( .A1(n13337), .A2(n11374), .ZN(n13967) );
  NOR2_X1 U15491 ( .A1(n13944), .A2(n13338), .ZN(n13341) );
  AOI21_X1 U15492 ( .B1(n13339), .B2(P2_B_REG_SCAN_IN), .A(n14784), .ZN(n13378) );
  NAND2_X1 U15493 ( .A1(n13378), .A2(n13340), .ZN(n13969) );
  NOR2_X1 U15494 ( .A1(n13969), .A2(n15059), .ZN(n13347) );
  AOI211_X1 U15495 ( .C1(n13966), .C2(n15060), .A(n13341), .B(n13347), .ZN(
        n13342) );
  OAI21_X1 U15496 ( .B1(n13967), .B2(n13937), .A(n13342), .ZN(P2_U3234) );
  OAI211_X1 U15497 ( .C1(n7084), .C2(n7082), .A(n13345), .B(n15065), .ZN(
        n13970) );
  NOR2_X1 U15498 ( .A1(n7082), .A2(n13959), .ZN(n13346) );
  AOI211_X1 U15499 ( .C1(n15059), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13347), 
        .B(n13346), .ZN(n13348) );
  OAI21_X1 U15500 ( .B1(n13937), .B2(n13970), .A(n13348), .ZN(P2_U3235) );
  INV_X1 U15501 ( .A(n14016), .ZN(n13884) );
  INV_X1 U15502 ( .A(n13904), .ZN(n13918) );
  INV_X1 U15503 ( .A(n14027), .ZN(n13916) );
  INV_X1 U15504 ( .A(n13823), .ZN(n13835) );
  NAND2_X1 U15505 ( .A1(n13836), .A2(n13835), .ZN(n13834) );
  NAND2_X1 U15506 ( .A1(n13834), .A2(n7594), .ZN(n13812) );
  NAND2_X1 U15507 ( .A1(n13812), .A2(n13811), .ZN(n13810) );
  XNOR2_X1 U15508 ( .A(n13359), .B(n13375), .ZN(n13972) );
  INV_X1 U15509 ( .A(n13972), .ZN(n13389) );
  INV_X1 U15510 ( .A(n14010), .ZN(n13366) );
  NOR2_X1 U15511 ( .A1(n7070), .A2(n13907), .ZN(n13872) );
  NOR2_X1 U15512 ( .A1(n13990), .A2(n13373), .ZN(n13410) );
  OR3_X2 U15513 ( .A1(n13788), .A2(n13410), .A3(n13409), .ZN(n13411) );
  AOI22_X1 U15514 ( .A1(n13378), .A2(n13377), .B1(n13376), .B2(n14787), .ZN(
        n13379) );
  INV_X1 U15515 ( .A(n13381), .ZN(n13392) );
  OAI211_X1 U15516 ( .C1(n7083), .C2(n13392), .A(n11374), .B(n13382), .ZN(
        n13974) );
  NOR2_X1 U15517 ( .A1(n13974), .A2(n13937), .ZN(n13387) );
  INV_X1 U15518 ( .A(n13383), .ZN(n13384) );
  AOI22_X1 U15519 ( .A1(n15059), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n15058), 
        .B2(n13384), .ZN(n13385) );
  OAI21_X1 U15520 ( .B1(n7083), .B2(n13959), .A(n13385), .ZN(n13386) );
  AOI211_X1 U15521 ( .C1(n13973), .C2(n13944), .A(n13387), .B(n13386), .ZN(
        n13388) );
  OAI21_X1 U15522 ( .B1(n13389), .B2(n13941), .A(n13388), .ZN(P2_U3236) );
  INV_X1 U15523 ( .A(n13403), .ZN(n13393) );
  AOI211_X1 U15524 ( .C1(n13980), .C2(n13393), .A(n6611), .B(n13392), .ZN(
        n13979) );
  NOR2_X1 U15525 ( .A1(n13394), .A2(n13959), .ZN(n13398) );
  OAI22_X1 U15526 ( .A1(n13944), .A2(n13396), .B1(n13395), .B2(n13957), .ZN(
        n13397) );
  AOI211_X1 U15527 ( .C1(n13979), .C2(n15068), .A(n13398), .B(n13397), .ZN(
        n13401) );
  XNOR2_X1 U15528 ( .A(n13399), .B(n6614), .ZN(n13983) );
  OR2_X1 U15529 ( .A1(n13983), .A2(n13941), .ZN(n13400) );
  OAI211_X1 U15530 ( .C1(n13982), .C2(n15059), .A(n13401), .B(n13400), .ZN(
        P2_U3237) );
  AOI211_X1 U15531 ( .C1(n13985), .C2(n13794), .A(n6611), .B(n13403), .ZN(
        n13984) );
  INV_X1 U15532 ( .A(n13985), .ZN(n13408) );
  INV_X1 U15533 ( .A(n13405), .ZN(n13406) );
  AOI22_X1 U15534 ( .A1(n15059), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n15058), 
        .B2(n13406), .ZN(n13407) );
  OAI21_X1 U15535 ( .B1(n13408), .B2(n13959), .A(n13407), .ZN(n13416) );
  OAI21_X1 U15536 ( .B1(n13788), .B2(n13410), .A(n13409), .ZN(n13412) );
  AOI21_X1 U15537 ( .B1(n13412), .B2(n13411), .A(n13925), .ZN(n13414) );
  NOR2_X1 U15538 ( .A1(n13987), .A2(n15059), .ZN(n13415) );
  OAI21_X1 U15539 ( .B1(n13988), .B2(n13941), .A(n13417), .ZN(P2_U3238) );
  AOI22_X1 U15540 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(keyinput225), .B1(
        P3_IR_REG_16__SCAN_IN), .B2(keyinput154), .ZN(n13418) );
  OAI221_X1 U15541 ( .B1(P1_DATAO_REG_2__SCAN_IN), .B2(keyinput225), .C1(
        P3_IR_REG_16__SCAN_IN), .C2(keyinput154), .A(n13418), .ZN(n13425) );
  AOI22_X1 U15542 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(keyinput146), .B1(
        P2_REG2_REG_19__SCAN_IN), .B2(keyinput202), .ZN(n13419) );
  OAI221_X1 U15543 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(keyinput146), .C1(
        P2_REG2_REG_19__SCAN_IN), .C2(keyinput202), .A(n13419), .ZN(n13424) );
  AOI22_X1 U15544 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(keyinput210), .B1(
        P3_REG3_REG_8__SCAN_IN), .B2(keyinput221), .ZN(n13420) );
  OAI221_X1 U15545 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(keyinput210), .C1(
        P3_REG3_REG_8__SCAN_IN), .C2(keyinput221), .A(n13420), .ZN(n13423) );
  AOI22_X1 U15546 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(keyinput165), .B1(
        P3_REG3_REG_23__SCAN_IN), .B2(keyinput242), .ZN(n13421) );
  OAI221_X1 U15547 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(keyinput165), .C1(
        P3_REG3_REG_23__SCAN_IN), .C2(keyinput242), .A(n13421), .ZN(n13422) );
  NOR4_X1 U15548 ( .A1(n13425), .A2(n13424), .A3(n13423), .A4(n13422), .ZN(
        n13453) );
  AOI22_X1 U15549 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(keyinput247), .B1(
        P1_REG3_REG_6__SCAN_IN), .B2(keyinput243), .ZN(n13426) );
  OAI221_X1 U15550 ( .B1(P3_ADDR_REG_1__SCAN_IN), .B2(keyinput247), .C1(
        P1_REG3_REG_6__SCAN_IN), .C2(keyinput243), .A(n13426), .ZN(n13433) );
  AOI22_X1 U15551 ( .A1(P2_REG2_REG_28__SCAN_IN), .A2(keyinput159), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(keyinput183), .ZN(n13427) );
  OAI221_X1 U15552 ( .B1(P2_REG2_REG_28__SCAN_IN), .B2(keyinput159), .C1(
        P2_DATAO_REG_4__SCAN_IN), .C2(keyinput183), .A(n13427), .ZN(n13432) );
  AOI22_X1 U15553 ( .A1(P2_REG1_REG_23__SCAN_IN), .A2(keyinput238), .B1(
        P3_IR_REG_13__SCAN_IN), .B2(keyinput192), .ZN(n13428) );
  OAI221_X1 U15554 ( .B1(P2_REG1_REG_23__SCAN_IN), .B2(keyinput238), .C1(
        P3_IR_REG_13__SCAN_IN), .C2(keyinput192), .A(n13428), .ZN(n13431) );
  AOI22_X1 U15555 ( .A1(P3_WR_REG_SCAN_IN), .A2(keyinput204), .B1(
        P3_REG3_REG_16__SCAN_IN), .B2(keyinput180), .ZN(n13429) );
  OAI221_X1 U15556 ( .B1(P3_WR_REG_SCAN_IN), .B2(keyinput204), .C1(
        P3_REG3_REG_16__SCAN_IN), .C2(keyinput180), .A(n13429), .ZN(n13430) );
  NOR4_X1 U15557 ( .A1(n13433), .A2(n13432), .A3(n13431), .A4(n13430), .ZN(
        n13452) );
  AOI22_X1 U15558 ( .A1(P1_REG2_REG_3__SCAN_IN), .A2(keyinput235), .B1(SI_28_), 
        .B2(keyinput237), .ZN(n13434) );
  OAI221_X1 U15559 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(keyinput235), .C1(SI_28_), .C2(keyinput237), .A(n13434), .ZN(n13441) );
  AOI22_X1 U15560 ( .A1(P1_REG0_REG_21__SCAN_IN), .A2(keyinput236), .B1(
        P2_REG0_REG_10__SCAN_IN), .B2(keyinput254), .ZN(n13435) );
  OAI221_X1 U15561 ( .B1(P1_REG0_REG_21__SCAN_IN), .B2(keyinput236), .C1(
        P2_REG0_REG_10__SCAN_IN), .C2(keyinput254), .A(n13435), .ZN(n13440) );
  AOI22_X1 U15562 ( .A1(P1_REG0_REG_7__SCAN_IN), .A2(keyinput147), .B1(
        P1_IR_REG_18__SCAN_IN), .B2(keyinput174), .ZN(n13436) );
  OAI221_X1 U15563 ( .B1(P1_REG0_REG_7__SCAN_IN), .B2(keyinput147), .C1(
        P1_IR_REG_18__SCAN_IN), .C2(keyinput174), .A(n13436), .ZN(n13439) );
  AOI22_X1 U15564 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(keyinput188), .B1(
        P3_REG1_REG_29__SCAN_IN), .B2(keyinput246), .ZN(n13437) );
  OAI221_X1 U15565 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(keyinput188), .C1(
        P3_REG1_REG_29__SCAN_IN), .C2(keyinput246), .A(n13437), .ZN(n13438) );
  NOR4_X1 U15566 ( .A1(n13441), .A2(n13440), .A3(n13439), .A4(n13438), .ZN(
        n13451) );
  AOI22_X1 U15567 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(keyinput157), .B1(
        P2_IR_REG_17__SCAN_IN), .B2(keyinput207), .ZN(n13442) );
  OAI221_X1 U15568 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(keyinput157), .C1(
        P2_IR_REG_17__SCAN_IN), .C2(keyinput207), .A(n13442), .ZN(n13449) );
  AOI22_X1 U15569 ( .A1(SI_31_), .A2(keyinput137), .B1(P1_REG1_REG_5__SCAN_IN), 
        .B2(keyinput233), .ZN(n13443) );
  OAI221_X1 U15570 ( .B1(SI_31_), .B2(keyinput137), .C1(P1_REG1_REG_5__SCAN_IN), .C2(keyinput233), .A(n13443), .ZN(n13448) );
  AOI22_X1 U15571 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(keyinput158), .B1(
        P3_REG1_REG_19__SCAN_IN), .B2(keyinput178), .ZN(n13444) );
  OAI221_X1 U15572 ( .B1(P1_DATAO_REG_30__SCAN_IN), .B2(keyinput158), .C1(
        P3_REG1_REG_19__SCAN_IN), .C2(keyinput178), .A(n13444), .ZN(n13447) );
  AOI22_X1 U15573 ( .A1(P3_REG0_REG_23__SCAN_IN), .A2(keyinput255), .B1(
        P1_ADDR_REG_19__SCAN_IN), .B2(keyinput148), .ZN(n13445) );
  OAI221_X1 U15574 ( .B1(P3_REG0_REG_23__SCAN_IN), .B2(keyinput255), .C1(
        P1_ADDR_REG_19__SCAN_IN), .C2(keyinput148), .A(n13445), .ZN(n13446) );
  NOR4_X1 U15575 ( .A1(n13449), .A2(n13448), .A3(n13447), .A4(n13446), .ZN(
        n13450) );
  NAND4_X1 U15576 ( .A1(n13453), .A2(n13452), .A3(n13451), .A4(n13450), .ZN(
        n13589) );
  AOI22_X1 U15577 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(keyinput156), .B1(
        P3_REG1_REG_9__SCAN_IN), .B2(keyinput234), .ZN(n13454) );
  OAI221_X1 U15578 ( .B1(P2_IR_REG_18__SCAN_IN), .B2(keyinput156), .C1(
        P3_REG1_REG_9__SCAN_IN), .C2(keyinput234), .A(n13454), .ZN(n13461) );
  AOI22_X1 U15579 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(keyinput155), .B1(
        P1_D_REG_10__SCAN_IN), .B2(keyinput252), .ZN(n13455) );
  OAI221_X1 U15580 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(keyinput155), .C1(
        P1_D_REG_10__SCAN_IN), .C2(keyinput252), .A(n13455), .ZN(n13460) );
  AOI22_X1 U15581 ( .A1(P1_REG0_REG_29__SCAN_IN), .A2(keyinput196), .B1(SI_4_), 
        .B2(keyinput150), .ZN(n13456) );
  OAI221_X1 U15582 ( .B1(P1_REG0_REG_29__SCAN_IN), .B2(keyinput196), .C1(SI_4_), .C2(keyinput150), .A(n13456), .ZN(n13459) );
  AOI22_X1 U15583 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(keyinput223), .B1(
        P3_REG1_REG_12__SCAN_IN), .B2(keyinput203), .ZN(n13457) );
  OAI221_X1 U15584 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(keyinput223), .C1(
        P3_REG1_REG_12__SCAN_IN), .C2(keyinput203), .A(n13457), .ZN(n13458) );
  NOR4_X1 U15585 ( .A1(n13461), .A2(n13460), .A3(n13459), .A4(n13458), .ZN(
        n13489) );
  AOI22_X1 U15586 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(keyinput142), .B1(
        P1_REG2_REG_29__SCAN_IN), .B2(keyinput170), .ZN(n13462) );
  OAI221_X1 U15587 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(keyinput142), .C1(
        P1_REG2_REG_29__SCAN_IN), .C2(keyinput170), .A(n13462), .ZN(n13469) );
  AOI22_X1 U15588 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(keyinput177), .B1(
        P1_D_REG_15__SCAN_IN), .B2(keyinput138), .ZN(n13463) );
  OAI221_X1 U15589 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(keyinput177), .C1(
        P1_D_REG_15__SCAN_IN), .C2(keyinput138), .A(n13463), .ZN(n13468) );
  AOI22_X1 U15590 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(keyinput149), .B1(
        P3_D_REG_27__SCAN_IN), .B2(keyinput200), .ZN(n13464) );
  OAI221_X1 U15591 ( .B1(P2_DATAO_REG_19__SCAN_IN), .B2(keyinput149), .C1(
        P3_D_REG_27__SCAN_IN), .C2(keyinput200), .A(n13464), .ZN(n13467) );
  AOI22_X1 U15592 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(keyinput164), .B1(
        P3_REG0_REG_2__SCAN_IN), .B2(keyinput151), .ZN(n13465) );
  OAI221_X1 U15593 ( .B1(P2_ADDR_REG_1__SCAN_IN), .B2(keyinput164), .C1(
        P3_REG0_REG_2__SCAN_IN), .C2(keyinput151), .A(n13465), .ZN(n13466) );
  NOR4_X1 U15594 ( .A1(n13469), .A2(n13468), .A3(n13467), .A4(n13466), .ZN(
        n13488) );
  AOI22_X1 U15595 ( .A1(P3_REG3_REG_20__SCAN_IN), .A2(keyinput198), .B1(
        P3_IR_REG_23__SCAN_IN), .B2(keyinput224), .ZN(n13470) );
  OAI221_X1 U15596 ( .B1(P3_REG3_REG_20__SCAN_IN), .B2(keyinput198), .C1(
        P3_IR_REG_23__SCAN_IN), .C2(keyinput224), .A(n13470), .ZN(n13477) );
  AOI22_X1 U15597 ( .A1(P2_REG0_REG_21__SCAN_IN), .A2(keyinput191), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(keyinput143), .ZN(n13471) );
  OAI221_X1 U15598 ( .B1(P2_REG0_REG_21__SCAN_IN), .B2(keyinput191), .C1(
        P2_DATAO_REG_16__SCAN_IN), .C2(keyinput143), .A(n13471), .ZN(n13476)
         );
  AOI22_X1 U15599 ( .A1(P3_REG0_REG_12__SCAN_IN), .A2(keyinput128), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(keyinput244), .ZN(n13472) );
  OAI221_X1 U15600 ( .B1(P3_REG0_REG_12__SCAN_IN), .B2(keyinput128), .C1(
        P1_DATAO_REG_13__SCAN_IN), .C2(keyinput244), .A(n13472), .ZN(n13475)
         );
  AOI22_X1 U15601 ( .A1(P2_REG2_REG_1__SCAN_IN), .A2(keyinput229), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(keyinput218), .ZN(n13473) );
  OAI221_X1 U15602 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(keyinput229), .C1(
        P2_DATAO_REG_29__SCAN_IN), .C2(keyinput218), .A(n13473), .ZN(n13474)
         );
  NOR4_X1 U15603 ( .A1(n13477), .A2(n13476), .A3(n13475), .A4(n13474), .ZN(
        n13487) );
  AOI22_X1 U15604 ( .A1(P1_REG1_REG_19__SCAN_IN), .A2(keyinput130), .B1(
        P3_IR_REG_21__SCAN_IN), .B2(keyinput140), .ZN(n13478) );
  OAI221_X1 U15605 ( .B1(P1_REG1_REG_19__SCAN_IN), .B2(keyinput130), .C1(
        P3_IR_REG_21__SCAN_IN), .C2(keyinput140), .A(n13478), .ZN(n13485) );
  AOI22_X1 U15606 ( .A1(P3_DATAO_REG_21__SCAN_IN), .A2(keyinput190), .B1(
        SI_16_), .B2(keyinput153), .ZN(n13479) );
  OAI221_X1 U15607 ( .B1(P3_DATAO_REG_21__SCAN_IN), .B2(keyinput190), .C1(
        SI_16_), .C2(keyinput153), .A(n13479), .ZN(n13484) );
  AOI22_X1 U15608 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(keyinput206), .B1(
        P3_D_REG_26__SCAN_IN), .B2(keyinput166), .ZN(n13480) );
  OAI221_X1 U15609 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(keyinput206), .C1(
        P3_D_REG_26__SCAN_IN), .C2(keyinput166), .A(n13480), .ZN(n13483) );
  AOI22_X1 U15610 ( .A1(P3_DATAO_REG_27__SCAN_IN), .A2(keyinput139), .B1(
        P2_D_REG_12__SCAN_IN), .B2(keyinput182), .ZN(n13481) );
  OAI221_X1 U15611 ( .B1(P3_DATAO_REG_27__SCAN_IN), .B2(keyinput139), .C1(
        P2_D_REG_12__SCAN_IN), .C2(keyinput182), .A(n13481), .ZN(n13482) );
  NOR4_X1 U15612 ( .A1(n13485), .A2(n13484), .A3(n13483), .A4(n13482), .ZN(
        n13486) );
  NAND4_X1 U15613 ( .A1(n13489), .A2(n13488), .A3(n13487), .A4(n13486), .ZN(
        n13588) );
  AOI22_X1 U15614 ( .A1(n9942), .A2(keyinput173), .B1(n13491), .B2(keyinput172), .ZN(n13490) );
  OAI221_X1 U15615 ( .B1(n9942), .B2(keyinput173), .C1(n13491), .C2(
        keyinput172), .A(n13490), .ZN(n13495) );
  XNOR2_X1 U15616 ( .A(n13492), .B(keyinput217), .ZN(n13494) );
  XNOR2_X1 U15617 ( .A(n15077), .B(keyinput152), .ZN(n13493) );
  OR3_X1 U15618 ( .A1(n13495), .A2(n13494), .A3(n13493), .ZN(n13501) );
  AOI22_X1 U15619 ( .A1(n13497), .A2(keyinput187), .B1(n15076), .B2(
        keyinput160), .ZN(n13496) );
  OAI221_X1 U15620 ( .B1(n13497), .B2(keyinput187), .C1(n15076), .C2(
        keyinput160), .A(n13496), .ZN(n13500) );
  AOI22_X1 U15621 ( .A1(n13687), .A2(keyinput197), .B1(n15075), .B2(
        keyinput216), .ZN(n13498) );
  OAI221_X1 U15622 ( .B1(n13687), .B2(keyinput197), .C1(n15075), .C2(
        keyinput216), .A(n13498), .ZN(n13499) );
  NOR3_X1 U15623 ( .A1(n13501), .A2(n13500), .A3(n13499), .ZN(n13536) );
  INV_X1 U15624 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n13503) );
  AOI22_X1 U15625 ( .A1(n13658), .A2(keyinput133), .B1(n13503), .B2(
        keyinput195), .ZN(n13502) );
  OAI221_X1 U15626 ( .B1(n13658), .B2(keyinput133), .C1(n13503), .C2(
        keyinput195), .A(n13502), .ZN(n13513) );
  AOI22_X1 U15627 ( .A1(n13506), .A2(keyinput214), .B1(keyinput205), .B2(
        n13505), .ZN(n13504) );
  OAI221_X1 U15628 ( .B1(n13506), .B2(keyinput214), .C1(n13505), .C2(
        keyinput205), .A(n13504), .ZN(n13512) );
  XNOR2_X1 U15629 ( .A(P2_IR_REG_23__SCAN_IN), .B(keyinput163), .ZN(n13510) );
  XNOR2_X1 U15630 ( .A(P3_IR_REG_31__SCAN_IN), .B(keyinput212), .ZN(n13509) );
  XNOR2_X1 U15631 ( .A(P3_REG2_REG_25__SCAN_IN), .B(keyinput213), .ZN(n13508)
         );
  XNOR2_X1 U15632 ( .A(keyinput141), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n13507)
         );
  NAND4_X1 U15633 ( .A1(n13510), .A2(n13509), .A3(n13508), .A4(n13507), .ZN(
        n13511) );
  NOR3_X1 U15634 ( .A1(n13513), .A2(n13512), .A3(n13511), .ZN(n13535) );
  AOI22_X1 U15635 ( .A1(n7794), .A2(keyinput181), .B1(keyinput134), .B2(n13698), .ZN(n13514) );
  OAI221_X1 U15636 ( .B1(n7794), .B2(keyinput181), .C1(n13698), .C2(
        keyinput134), .A(n13514), .ZN(n13522) );
  AOI22_X1 U15637 ( .A1(n14180), .A2(keyinput168), .B1(keyinput131), .B2(n7275), .ZN(n13515) );
  OAI221_X1 U15638 ( .B1(n14180), .B2(keyinput168), .C1(n7275), .C2(
        keyinput131), .A(n13515), .ZN(n13521) );
  INV_X1 U15639 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n14935) );
  INV_X1 U15640 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n13610) );
  AOI22_X1 U15641 ( .A1(n14935), .A2(keyinput249), .B1(n13610), .B2(
        keyinput161), .ZN(n13516) );
  OAI221_X1 U15642 ( .B1(n14935), .B2(keyinput249), .C1(n13610), .C2(
        keyinput161), .A(n13516), .ZN(n13520) );
  AOI22_X1 U15643 ( .A1(n13634), .A2(keyinput136), .B1(keyinput208), .B2(
        n13518), .ZN(n13517) );
  OAI221_X1 U15644 ( .B1(n13634), .B2(keyinput136), .C1(n13518), .C2(
        keyinput208), .A(n13517), .ZN(n13519) );
  NOR4_X1 U15645 ( .A1(n13522), .A2(n13521), .A3(n13520), .A4(n13519), .ZN(
        n13534) );
  INV_X1 U15646 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n13694) );
  AOI22_X1 U15647 ( .A1(n13694), .A2(keyinput186), .B1(keyinput241), .B2(
        n13724), .ZN(n13523) );
  OAI221_X1 U15648 ( .B1(n13694), .B2(keyinput186), .C1(n13724), .C2(
        keyinput241), .A(n13523), .ZN(n13532) );
  XNOR2_X1 U15649 ( .A(n13524), .B(keyinput189), .ZN(n13531) );
  XNOR2_X1 U15650 ( .A(keyinput194), .B(n13952), .ZN(n13530) );
  XNOR2_X1 U15651 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput250), .ZN(n13528) );
  XNOR2_X1 U15652 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput185), .ZN(n13527) );
  XNOR2_X1 U15653 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput167), .ZN(n13526) );
  XNOR2_X1 U15654 ( .A(P3_IR_REG_25__SCAN_IN), .B(keyinput184), .ZN(n13525) );
  NAND4_X1 U15655 ( .A1(n13528), .A2(n13527), .A3(n13526), .A4(n13525), .ZN(
        n13529) );
  NOR4_X1 U15656 ( .A1(n13532), .A2(n13531), .A3(n13530), .A4(n13529), .ZN(
        n13533) );
  NAND4_X1 U15657 ( .A1(n13536), .A2(n13535), .A3(n13534), .A4(n13533), .ZN(
        n13587) );
  AOI22_X1 U15658 ( .A1(n13539), .A2(keyinput240), .B1(n13538), .B2(
        keyinput215), .ZN(n13537) );
  OAI221_X1 U15659 ( .B1(n13539), .B2(keyinput240), .C1(n13538), .C2(
        keyinput215), .A(n13537), .ZN(n13549) );
  AOI22_X1 U15660 ( .A1(n13541), .A2(keyinput162), .B1(keyinput211), .B2(
        n14911), .ZN(n13540) );
  OAI221_X1 U15661 ( .B1(n13541), .B2(keyinput162), .C1(n14911), .C2(
        keyinput211), .A(n13540), .ZN(n13548) );
  XNOR2_X1 U15662 ( .A(n13542), .B(keyinput179), .ZN(n13547) );
  XNOR2_X1 U15663 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(keyinput171), .ZN(n13545)
         );
  XNOR2_X1 U15664 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput232), .ZN(n13544) );
  XNOR2_X1 U15665 ( .A(P3_REG0_REG_18__SCAN_IN), .B(keyinput248), .ZN(n13543)
         );
  NAND3_X1 U15666 ( .A1(n13545), .A2(n13544), .A3(n13543), .ZN(n13546) );
  NOR4_X1 U15667 ( .A1(n13549), .A2(n13548), .A3(n13547), .A4(n13546), .ZN(
        n13585) );
  AOI22_X1 U15668 ( .A1(n13552), .A2(keyinput228), .B1(keyinput132), .B2(
        n13551), .ZN(n13550) );
  OAI221_X1 U15669 ( .B1(n13552), .B2(keyinput228), .C1(n13551), .C2(
        keyinput132), .A(n13550), .ZN(n13560) );
  AOI22_X1 U15670 ( .A1(n15074), .A2(keyinput227), .B1(n13779), .B2(
        keyinput145), .ZN(n13553) );
  OAI221_X1 U15671 ( .B1(n15074), .B2(keyinput227), .C1(n13779), .C2(
        keyinput145), .A(n13553), .ZN(n13559) );
  XNOR2_X1 U15672 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput245), .ZN(n13557) );
  XNOR2_X1 U15673 ( .A(P2_IR_REG_28__SCAN_IN), .B(keyinput201), .ZN(n13556) );
  XNOR2_X1 U15674 ( .A(P3_IR_REG_11__SCAN_IN), .B(keyinput230), .ZN(n13555) );
  XNOR2_X1 U15675 ( .A(P3_REG3_REG_28__SCAN_IN), .B(keyinput175), .ZN(n13554)
         );
  NAND4_X1 U15676 ( .A1(n13557), .A2(n13556), .A3(n13555), .A4(n13554), .ZN(
        n13558) );
  NOR3_X1 U15677 ( .A1(n13560), .A2(n13559), .A3(n13558), .ZN(n13584) );
  AOI22_X1 U15678 ( .A1(n13711), .A2(keyinput135), .B1(keyinput193), .B2(
        n13716), .ZN(n13561) );
  OAI221_X1 U15679 ( .B1(n13711), .B2(keyinput135), .C1(n13716), .C2(
        keyinput193), .A(n13561), .ZN(n13571) );
  INV_X1 U15680 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n13564) );
  INV_X1 U15681 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n13563) );
  AOI22_X1 U15682 ( .A1(n13564), .A2(keyinput199), .B1(keyinput129), .B2(
        n13563), .ZN(n13562) );
  OAI221_X1 U15683 ( .B1(n13564), .B2(keyinput199), .C1(n13563), .C2(
        keyinput129), .A(n13562), .ZN(n13570) );
  XNOR2_X1 U15684 ( .A(P3_IR_REG_5__SCAN_IN), .B(keyinput220), .ZN(n13567) );
  XNOR2_X1 U15685 ( .A(P3_IR_REG_10__SCAN_IN), .B(keyinput222), .ZN(n13566) );
  XNOR2_X1 U15686 ( .A(P3_REG1_REG_28__SCAN_IN), .B(keyinput239), .ZN(n13565)
         );
  NAND3_X1 U15687 ( .A1(n13567), .A2(n13566), .A3(n13565), .ZN(n13569) );
  XNOR2_X1 U15688 ( .A(n13718), .B(keyinput209), .ZN(n13568) );
  NOR4_X1 U15689 ( .A1(n13571), .A2(n13570), .A3(n13569), .A4(n13568), .ZN(
        n13583) );
  AOI22_X1 U15690 ( .A1(n9978), .A2(keyinput169), .B1(n13686), .B2(keyinput144), .ZN(n13572) );
  OAI221_X1 U15691 ( .B1(n9978), .B2(keyinput169), .C1(n13686), .C2(
        keyinput144), .A(n13572), .ZN(n13581) );
  AOI22_X1 U15692 ( .A1(n13727), .A2(keyinput251), .B1(n13574), .B2(
        keyinput219), .ZN(n13573) );
  OAI221_X1 U15693 ( .B1(n13727), .B2(keyinput251), .C1(n13574), .C2(
        keyinput219), .A(n13573), .ZN(n13580) );
  INV_X1 U15694 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n13661) );
  XOR2_X1 U15695 ( .A(n13661), .B(keyinput253), .Z(n13578) );
  XNOR2_X1 U15696 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput226), .ZN(n13577) );
  XNOR2_X1 U15697 ( .A(P2_REG3_REG_5__SCAN_IN), .B(keyinput176), .ZN(n13576)
         );
  XNOR2_X1 U15698 ( .A(P3_IR_REG_30__SCAN_IN), .B(keyinput231), .ZN(n13575) );
  NAND4_X1 U15699 ( .A1(n13578), .A2(n13577), .A3(n13576), .A4(n13575), .ZN(
        n13579) );
  NOR3_X1 U15700 ( .A1(n13581), .A2(n13580), .A3(n13579), .ZN(n13582) );
  NAND4_X1 U15701 ( .A1(n13585), .A2(n13584), .A3(n13583), .A4(n13582), .ZN(
        n13586) );
  NOR4_X1 U15702 ( .A1(n13589), .A2(n13588), .A3(n13587), .A4(n13586), .ZN(
        n13787) );
  AOI22_X1 U15703 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput45), .B1(
        P3_REG3_REG_18__SCAN_IN), .B2(keyinput71), .ZN(n13590) );
  OAI221_X1 U15704 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput45), .C1(
        P3_REG3_REG_18__SCAN_IN), .C2(keyinput71), .A(n13590), .ZN(n13597) );
  AOI22_X1 U15705 ( .A1(P2_REG2_REG_2__SCAN_IN), .A2(keyinput13), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(keyinput55), .ZN(n13591) );
  OAI221_X1 U15706 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(keyinput13), .C1(
        P2_DATAO_REG_4__SCAN_IN), .C2(keyinput55), .A(n13591), .ZN(n13596) );
  AOI22_X1 U15707 ( .A1(P3_ADDR_REG_12__SCAN_IN), .A2(keyinput51), .B1(
        P2_IR_REG_18__SCAN_IN), .B2(keyinput28), .ZN(n13592) );
  OAI221_X1 U15708 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(keyinput51), .C1(
        P2_IR_REG_18__SCAN_IN), .C2(keyinput28), .A(n13592), .ZN(n13595) );
  AOI22_X1 U15709 ( .A1(P3_ADDR_REG_11__SCAN_IN), .A2(keyinput112), .B1(
        P2_REG1_REG_15__SCAN_IN), .B2(keyinput78), .ZN(n13593) );
  OAI221_X1 U15710 ( .B1(P3_ADDR_REG_11__SCAN_IN), .B2(keyinput112), .C1(
        P2_REG1_REG_15__SCAN_IN), .C2(keyinput78), .A(n13593), .ZN(n13594) );
  NOR4_X1 U15711 ( .A1(n13597), .A2(n13596), .A3(n13595), .A4(n13594), .ZN(
        n13628) );
  AOI22_X1 U15712 ( .A1(P3_DATAO_REG_9__SCAN_IN), .A2(keyinput4), .B1(
        P2_ADDR_REG_9__SCAN_IN), .B2(keyinput60), .ZN(n13598) );
  OAI221_X1 U15713 ( .B1(P3_DATAO_REG_9__SCAN_IN), .B2(keyinput4), .C1(
        P2_ADDR_REG_9__SCAN_IN), .C2(keyinput60), .A(n13598), .ZN(n13605) );
  AOI22_X1 U15714 ( .A1(P3_REG0_REG_26__SCAN_IN), .A2(keyinput91), .B1(
        P3_REG1_REG_29__SCAN_IN), .B2(keyinput118), .ZN(n13599) );
  OAI221_X1 U15715 ( .B1(P3_REG0_REG_26__SCAN_IN), .B2(keyinput91), .C1(
        P3_REG1_REG_29__SCAN_IN), .C2(keyinput118), .A(n13599), .ZN(n13604) );
  AOI22_X1 U15716 ( .A1(P3_REG0_REG_4__SCAN_IN), .A2(keyinput1), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(keyinput21), .ZN(n13600) );
  OAI221_X1 U15717 ( .B1(P3_REG0_REG_4__SCAN_IN), .B2(keyinput1), .C1(
        P2_DATAO_REG_19__SCAN_IN), .C2(keyinput21), .A(n13600), .ZN(n13603) );
  AOI22_X1 U15718 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(keyinput18), .B1(
        P2_REG2_REG_16__SCAN_IN), .B2(keyinput77), .ZN(n13601) );
  OAI221_X1 U15719 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(keyinput18), .C1(
        P2_REG2_REG_16__SCAN_IN), .C2(keyinput77), .A(n13601), .ZN(n13602) );
  NOR4_X1 U15720 ( .A1(n13605), .A2(n13604), .A3(n13603), .A4(n13602), .ZN(
        n13627) );
  AOI22_X1 U15721 ( .A1(n13607), .A2(keyinput72), .B1(keyinput66), .B2(n13952), 
        .ZN(n13606) );
  OAI221_X1 U15722 ( .B1(n13607), .B2(keyinput72), .C1(n13952), .C2(keyinput66), .A(n13606), .ZN(n13616) );
  AOI22_X1 U15723 ( .A1(P1_REG1_REG_19__SCAN_IN), .A2(keyinput2), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(keyinput80), .ZN(n13608) );
  OAI221_X1 U15724 ( .B1(P1_REG1_REG_19__SCAN_IN), .B2(keyinput2), .C1(
        P1_DATAO_REG_16__SCAN_IN), .C2(keyinput80), .A(n13608), .ZN(n13615) );
  AOI22_X1 U15725 ( .A1(n13610), .A2(keyinput33), .B1(n9978), .B2(keyinput41), 
        .ZN(n13609) );
  OAI221_X1 U15726 ( .B1(n13610), .B2(keyinput33), .C1(n9978), .C2(keyinput41), 
        .A(n13609), .ZN(n13614) );
  INV_X1 U15727 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15390) );
  AOI22_X1 U15728 ( .A1(n15390), .A2(keyinput23), .B1(keyinput62), .B2(n13612), 
        .ZN(n13611) );
  OAI221_X1 U15729 ( .B1(n15390), .B2(keyinput23), .C1(n13612), .C2(keyinput62), .A(n13611), .ZN(n13613) );
  NOR4_X1 U15730 ( .A1(n13616), .A2(n13615), .A3(n13614), .A4(n13613), .ZN(
        n13626) );
  AOI22_X1 U15731 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(keyinput59), .B1(
        P3_REG2_REG_25__SCAN_IN), .B2(keyinput85), .ZN(n13617) );
  OAI221_X1 U15732 ( .B1(P3_ADDR_REG_15__SCAN_IN), .B2(keyinput59), .C1(
        P3_REG2_REG_25__SCAN_IN), .C2(keyinput85), .A(n13617), .ZN(n13624) );
  AOI22_X1 U15733 ( .A1(P2_REG2_REG_28__SCAN_IN), .A2(keyinput31), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(keyinput61), .ZN(n13618) );
  OAI221_X1 U15734 ( .B1(P2_REG2_REG_28__SCAN_IN), .B2(keyinput31), .C1(
        P2_DATAO_REG_26__SCAN_IN), .C2(keyinput61), .A(n13618), .ZN(n13623) );
  AOI22_X1 U15735 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(keyinput52), .B1(
        P3_IR_REG_31__SCAN_IN), .B2(keyinput84), .ZN(n13619) );
  OAI221_X1 U15736 ( .B1(P3_REG3_REG_16__SCAN_IN), .B2(keyinput52), .C1(
        P3_IR_REG_31__SCAN_IN), .C2(keyinput84), .A(n13619), .ZN(n13622) );
  AOI22_X1 U15737 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(keyinput36), .B1(
        P2_REG2_REG_1__SCAN_IN), .B2(keyinput101), .ZN(n13620) );
  OAI221_X1 U15738 ( .B1(P2_ADDR_REG_1__SCAN_IN), .B2(keyinput36), .C1(
        P2_REG2_REG_1__SCAN_IN), .C2(keyinput101), .A(n13620), .ZN(n13621) );
  NOR4_X1 U15739 ( .A1(n13624), .A2(n13623), .A3(n13622), .A4(n13621), .ZN(
        n13625) );
  NAND4_X1 U15740 ( .A1(n13628), .A2(n13627), .A3(n13626), .A4(n13625), .ZN(
        n13786) );
  XOR2_X1 U15741 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput117), .Z(n13633) );
  XOR2_X1 U15742 ( .A(P1_REG2_REG_0__SCAN_IN), .B(keyinput82), .Z(n13632) );
  XOR2_X1 U15743 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput39), .Z(n13631) );
  XNOR2_X1 U15744 ( .A(n13629), .B(keyinput46), .ZN(n13630) );
  NOR4_X1 U15745 ( .A1(n13633), .A2(n13632), .A3(n13631), .A4(n13630), .ZN(
        n13656) );
  XNOR2_X1 U15746 ( .A(n13634), .B(keyinput8), .ZN(n13641) );
  XNOR2_X1 U15747 ( .A(n13635), .B(keyinput35), .ZN(n13640) );
  XNOR2_X1 U15748 ( .A(n13636), .B(keyinput79), .ZN(n13639) );
  XNOR2_X1 U15749 ( .A(n13637), .B(keyinput73), .ZN(n13638) );
  NOR4_X1 U15750 ( .A1(n13641), .A2(n13640), .A3(n13639), .A4(n13638), .ZN(
        n13655) );
  XOR2_X1 U15751 ( .A(P3_IR_REG_5__SCAN_IN), .B(keyinput92), .Z(n13647) );
  XOR2_X1 U15752 ( .A(P2_REG2_REG_30__SCAN_IN), .B(keyinput87), .Z(n13646) );
  XNOR2_X1 U15753 ( .A(n13642), .B(keyinput26), .ZN(n13645) );
  XNOR2_X1 U15754 ( .A(n13643), .B(keyinput94), .ZN(n13644) );
  NOR4_X1 U15755 ( .A1(n13647), .A2(n13646), .A3(n13645), .A4(n13644), .ZN(
        n13654) );
  XOR2_X1 U15756 ( .A(P3_IR_REG_21__SCAN_IN), .B(keyinput12), .Z(n13652) );
  XOR2_X1 U15757 ( .A(P3_IR_REG_30__SCAN_IN), .B(keyinput103), .Z(n13651) );
  XNOR2_X1 U15758 ( .A(n8260), .B(keyinput96), .ZN(n13650) );
  XNOR2_X1 U15759 ( .A(n13648), .B(keyinput102), .ZN(n13649) );
  NOR4_X1 U15760 ( .A1(n13652), .A2(n13651), .A3(n13650), .A4(n13649), .ZN(
        n13653) );
  NAND4_X1 U15761 ( .A1(n13656), .A2(n13655), .A3(n13654), .A4(n13653), .ZN(
        n13670) );
  AOI22_X1 U15762 ( .A1(n13659), .A2(keyinput63), .B1(keyinput5), .B2(n13658), 
        .ZN(n13657) );
  OAI221_X1 U15763 ( .B1(n13659), .B2(keyinput63), .C1(n13658), .C2(keyinput5), 
        .A(n13657), .ZN(n13669) );
  INV_X1 U15764 ( .A(P3_WR_REG_SCAN_IN), .ZN(n13660) );
  XNOR2_X1 U15765 ( .A(n13660), .B(keyinput76), .ZN(n13668) );
  XOR2_X1 U15766 ( .A(keyinput125), .B(n13661), .Z(n13666) );
  XOR2_X1 U15767 ( .A(keyinput115), .B(n13662), .Z(n13665) );
  XOR2_X1 U15768 ( .A(keyinput29), .B(n11502), .Z(n13664) );
  XOR2_X1 U15769 ( .A(keyinput3), .B(n7275), .Z(n13663) );
  NAND4_X1 U15770 ( .A1(n13666), .A2(n13665), .A3(n13664), .A4(n13663), .ZN(
        n13667) );
  NOR4_X1 U15771 ( .A1(n13670), .A2(n13669), .A3(n13668), .A4(n13667), .ZN(
        n13704) );
  AOI22_X1 U15772 ( .A1(n13672), .A2(keyinput119), .B1(n8483), .B2(keyinput19), 
        .ZN(n13671) );
  OAI221_X1 U15773 ( .B1(n13672), .B2(keyinput119), .C1(n8483), .C2(keyinput19), .A(n13671), .ZN(n13681) );
  AOI22_X1 U15774 ( .A1(n13675), .A2(keyinput42), .B1(n13674), .B2(keyinput108), .ZN(n13673) );
  OAI221_X1 U15775 ( .B1(n13675), .B2(keyinput42), .C1(n13674), .C2(
        keyinput108), .A(n13673), .ZN(n13680) );
  AOI22_X1 U15776 ( .A1(n14180), .A2(keyinput40), .B1(n13677), .B2(keyinput95), 
        .ZN(n13676) );
  OAI221_X1 U15777 ( .B1(n14180), .B2(keyinput40), .C1(n13677), .C2(keyinput95), .A(n13676), .ZN(n13679) );
  INV_X1 U15778 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n14928) );
  XNOR2_X1 U15779 ( .A(n14928), .B(keyinput10), .ZN(n13678) );
  NOR4_X1 U15780 ( .A1(n13681), .A2(n13680), .A3(n13679), .A4(n13678), .ZN(
        n13703) );
  INV_X1 U15781 ( .A(SI_31_), .ZN(n13683) );
  AOI22_X1 U15782 ( .A1(n13684), .A2(keyinput47), .B1(keyinput9), .B2(n13683), 
        .ZN(n13682) );
  OAI221_X1 U15783 ( .B1(n13684), .B2(keyinput47), .C1(n13683), .C2(keyinput9), 
        .A(n13682), .ZN(n13692) );
  AOI22_X1 U15784 ( .A1(n13687), .A2(keyinput69), .B1(n13686), .B2(keyinput16), 
        .ZN(n13685) );
  OAI221_X1 U15785 ( .B1(n13687), .B2(keyinput69), .C1(n13686), .C2(keyinput16), .A(n13685), .ZN(n13691) );
  AOI22_X1 U15786 ( .A1(n13689), .A2(keyinput75), .B1(n14670), .B2(keyinput90), 
        .ZN(n13688) );
  OAI221_X1 U15787 ( .B1(n13689), .B2(keyinput75), .C1(n14670), .C2(keyinput90), .A(n13688), .ZN(n13690) );
  NOR3_X1 U15788 ( .A1(n13692), .A2(n13691), .A3(n13690), .ZN(n13702) );
  AOI22_X1 U15789 ( .A1(n13695), .A2(keyinput11), .B1(n13694), .B2(keyinput58), 
        .ZN(n13693) );
  OAI221_X1 U15790 ( .B1(n13695), .B2(keyinput11), .C1(n13694), .C2(keyinput58), .A(n13693), .ZN(n13700) );
  INV_X1 U15791 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n13697) );
  AOI22_X1 U15792 ( .A1(n13698), .A2(keyinput6), .B1(keyinput37), .B2(n13697), 
        .ZN(n13696) );
  OAI221_X1 U15793 ( .B1(n13698), .B2(keyinput6), .C1(n13697), .C2(keyinput37), 
        .A(n13696), .ZN(n13699) );
  NOR2_X1 U15794 ( .A1(n13700), .A2(n13699), .ZN(n13701) );
  NAND4_X1 U15795 ( .A1(n13704), .A2(n13703), .A3(n13702), .A4(n13701), .ZN(
        n13785) );
  AOI22_X1 U15796 ( .A1(n13706), .A2(keyinput0), .B1(keyinput105), .B2(n9833), 
        .ZN(n13705) );
  OAI221_X1 U15797 ( .B1(n13706), .B2(keyinput0), .C1(n9833), .C2(keyinput105), 
        .A(n13705), .ZN(n13714) );
  AOI22_X1 U15798 ( .A1(n13708), .A2(keyinput122), .B1(keyinput83), .B2(n14911), .ZN(n13707) );
  OAI221_X1 U15799 ( .B1(n13708), .B2(keyinput122), .C1(n14911), .C2(
        keyinput83), .A(n13707), .ZN(n13713) );
  AOI22_X1 U15800 ( .A1(n13711), .A2(keyinput7), .B1(n13710), .B2(keyinput120), 
        .ZN(n13709) );
  OAI221_X1 U15801 ( .B1(n13711), .B2(keyinput7), .C1(n13710), .C2(keyinput120), .A(n13709), .ZN(n13712) );
  OR3_X1 U15802 ( .A1(n13714), .A2(n13713), .A3(n13712), .ZN(n13722) );
  AOI22_X1 U15803 ( .A1(n13716), .A2(keyinput65), .B1(n14935), .B2(keyinput121), .ZN(n13715) );
  OAI221_X1 U15804 ( .B1(n13716), .B2(keyinput65), .C1(n14935), .C2(
        keyinput121), .A(n13715), .ZN(n13721) );
  AOI22_X1 U15805 ( .A1(n13719), .A2(keyinput93), .B1(keyinput81), .B2(n13718), 
        .ZN(n13717) );
  OAI221_X1 U15806 ( .B1(n13719), .B2(keyinput93), .C1(n13718), .C2(keyinput81), .A(n13717), .ZN(n13720) );
  NOR3_X1 U15807 ( .A1(n13722), .A2(n13721), .A3(n13720), .ZN(n13739) );
  XOR2_X1 U15808 ( .A(n15074), .B(keyinput99), .Z(n13738) );
  XOR2_X1 U15809 ( .A(n15076), .B(keyinput32), .Z(n13737) );
  AOI22_X1 U15810 ( .A1(n13725), .A2(keyinput114), .B1(keyinput113), .B2(
        n13724), .ZN(n13723) );
  OAI221_X1 U15811 ( .B1(n13725), .B2(keyinput114), .C1(n13724), .C2(
        keyinput113), .A(n13723), .ZN(n13735) );
  AOI22_X1 U15812 ( .A1(n13728), .A2(keyinput38), .B1(keyinput123), .B2(n13727), .ZN(n13726) );
  OAI221_X1 U15813 ( .B1(n13728), .B2(keyinput38), .C1(n13727), .C2(
        keyinput123), .A(n13726), .ZN(n13734) );
  XNOR2_X1 U15814 ( .A(SI_4_), .B(keyinput22), .ZN(n13732) );
  XNOR2_X1 U15815 ( .A(SI_16_), .B(keyinput25), .ZN(n13731) );
  XNOR2_X1 U15816 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput57), .ZN(n13730) );
  XNOR2_X1 U15817 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput89), .ZN(n13729) );
  NAND4_X1 U15818 ( .A1(n13732), .A2(n13731), .A3(n13730), .A4(n13729), .ZN(
        n13733) );
  NOR3_X1 U15819 ( .A1(n13735), .A2(n13734), .A3(n13733), .ZN(n13736) );
  NAND4_X1 U15820 ( .A1(n13739), .A2(n13738), .A3(n13737), .A4(n13736), .ZN(
        n13777) );
  AOI22_X1 U15821 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(keyinput27), .B1(
        P1_ADDR_REG_19__SCAN_IN), .B2(keyinput20), .ZN(n13740) );
  OAI221_X1 U15822 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(keyinput27), .C1(
        P1_ADDR_REG_19__SCAN_IN), .C2(keyinput20), .A(n13740), .ZN(n13747) );
  AOI22_X1 U15823 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(keyinput67), .B1(
        P2_D_REG_8__SCAN_IN), .B2(keyinput24), .ZN(n13741) );
  OAI221_X1 U15824 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(keyinput67), .C1(
        P2_D_REG_8__SCAN_IN), .C2(keyinput24), .A(n13741), .ZN(n13746) );
  AOI22_X1 U15825 ( .A1(P2_REG0_REG_10__SCAN_IN), .A2(keyinput126), .B1(
        P3_IR_REG_25__SCAN_IN), .B2(keyinput56), .ZN(n13742) );
  OAI221_X1 U15826 ( .B1(P2_REG0_REG_10__SCAN_IN), .B2(keyinput126), .C1(
        P3_IR_REG_25__SCAN_IN), .C2(keyinput56), .A(n13742), .ZN(n13745) );
  AOI22_X1 U15827 ( .A1(P2_D_REG_19__SCAN_IN), .A2(keyinput88), .B1(
        P3_IR_REG_13__SCAN_IN), .B2(keyinput64), .ZN(n13743) );
  OAI221_X1 U15828 ( .B1(P2_D_REG_19__SCAN_IN), .B2(keyinput88), .C1(
        P3_IR_REG_13__SCAN_IN), .C2(keyinput64), .A(n13743), .ZN(n13744) );
  NOR4_X1 U15829 ( .A1(n13747), .A2(n13746), .A3(n13745), .A4(n13744), .ZN(
        n13775) );
  AOI22_X1 U15830 ( .A1(P1_REG0_REG_29__SCAN_IN), .A2(keyinput68), .B1(
        P3_REG1_REG_28__SCAN_IN), .B2(keyinput111), .ZN(n13748) );
  OAI221_X1 U15831 ( .B1(P1_REG0_REG_29__SCAN_IN), .B2(keyinput68), .C1(
        P3_REG1_REG_28__SCAN_IN), .C2(keyinput111), .A(n13748), .ZN(n13755) );
  AOI22_X1 U15832 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(keyinput30), .B1(
        P2_D_REG_12__SCAN_IN), .B2(keyinput54), .ZN(n13749) );
  OAI221_X1 U15833 ( .B1(P1_DATAO_REG_30__SCAN_IN), .B2(keyinput30), .C1(
        P2_D_REG_12__SCAN_IN), .C2(keyinput54), .A(n13749), .ZN(n13754) );
  AOI22_X1 U15834 ( .A1(P1_D_REG_10__SCAN_IN), .A2(keyinput124), .B1(
        P2_REG3_REG_5__SCAN_IN), .B2(keyinput48), .ZN(n13750) );
  OAI221_X1 U15835 ( .B1(P1_D_REG_10__SCAN_IN), .B2(keyinput124), .C1(
        P2_REG3_REG_5__SCAN_IN), .C2(keyinput48), .A(n13750), .ZN(n13753) );
  AOI22_X1 U15836 ( .A1(P2_REG1_REG_23__SCAN_IN), .A2(keyinput110), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(keyinput43), .ZN(n13751) );
  OAI221_X1 U15837 ( .B1(P2_REG1_REG_23__SCAN_IN), .B2(keyinput110), .C1(
        P2_DATAO_REG_5__SCAN_IN), .C2(keyinput43), .A(n13751), .ZN(n13752) );
  NOR4_X1 U15838 ( .A1(n13755), .A2(n13754), .A3(n13753), .A4(n13752), .ZN(
        n13774) );
  AOI22_X1 U15839 ( .A1(P1_REG1_REG_22__SCAN_IN), .A2(keyinput100), .B1(
        P3_REG1_REG_9__SCAN_IN), .B2(keyinput106), .ZN(n13756) );
  OAI221_X1 U15840 ( .B1(P1_REG1_REG_22__SCAN_IN), .B2(keyinput100), .C1(
        P3_REG1_REG_9__SCAN_IN), .C2(keyinput106), .A(n13756), .ZN(n13763) );
  AOI22_X1 U15841 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(keyinput49), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(keyinput97), .ZN(n13757) );
  OAI221_X1 U15842 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(keyinput49), .C1(
        P1_DATAO_REG_2__SCAN_IN), .C2(keyinput97), .A(n13757), .ZN(n13762) );
  AOI22_X1 U15843 ( .A1(P3_REG1_REG_19__SCAN_IN), .A2(keyinput50), .B1(SI_28_), 
        .B2(keyinput109), .ZN(n13758) );
  OAI221_X1 U15844 ( .B1(P3_REG1_REG_19__SCAN_IN), .B2(keyinput50), .C1(SI_28_), .C2(keyinput109), .A(n13758), .ZN(n13761) );
  AOI22_X1 U15845 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(keyinput98), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(keyinput86), .ZN(n13759) );
  OAI221_X1 U15846 ( .B1(P1_IR_REG_13__SCAN_IN), .B2(keyinput98), .C1(
        P1_DATAO_REG_10__SCAN_IN), .C2(keyinput86), .A(n13759), .ZN(n13760) );
  NOR4_X1 U15847 ( .A1(n13763), .A2(n13762), .A3(n13761), .A4(n13760), .ZN(
        n13773) );
  AOI22_X1 U15848 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(keyinput104), .B1(
        P3_REG3_REG_20__SCAN_IN), .B2(keyinput70), .ZN(n13764) );
  OAI221_X1 U15849 ( .B1(P1_IR_REG_6__SCAN_IN), .B2(keyinput104), .C1(
        P3_REG3_REG_20__SCAN_IN), .C2(keyinput70), .A(n13764), .ZN(n13771) );
  AOI22_X1 U15850 ( .A1(P3_REG0_REG_23__SCAN_IN), .A2(keyinput127), .B1(
        P3_D_REG_24__SCAN_IN), .B2(keyinput44), .ZN(n13765) );
  OAI221_X1 U15851 ( .B1(P3_REG0_REG_23__SCAN_IN), .B2(keyinput127), .C1(
        P3_D_REG_24__SCAN_IN), .C2(keyinput44), .A(n13765), .ZN(n13770) );
  AOI22_X1 U15852 ( .A1(P1_REG2_REG_3__SCAN_IN), .A2(keyinput107), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(keyinput116), .ZN(n13766) );
  OAI221_X1 U15853 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(keyinput107), .C1(
        P1_DATAO_REG_13__SCAN_IN), .C2(keyinput116), .A(n13766), .ZN(n13769)
         );
  AOI22_X1 U15854 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(keyinput34), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(keyinput15), .ZN(n13767) );
  OAI221_X1 U15855 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(keyinput34), .C1(
        P2_DATAO_REG_16__SCAN_IN), .C2(keyinput15), .A(n13767), .ZN(n13768) );
  NOR4_X1 U15856 ( .A1(n13771), .A2(n13770), .A3(n13769), .A4(n13768), .ZN(
        n13772) );
  NAND4_X1 U15857 ( .A1(n13775), .A2(n13774), .A3(n13773), .A4(n13772), .ZN(
        n13776) );
  NOR2_X1 U15858 ( .A1(n13777), .A2(n13776), .ZN(n13783) );
  OAI22_X1 U15859 ( .A1(n13779), .A2(keyinput17), .B1(n15036), .B2(keyinput14), 
        .ZN(n13778) );
  AOI221_X1 U15860 ( .B1(n13779), .B2(keyinput17), .C1(keyinput14), .C2(n15036), .A(n13778), .ZN(n13782) );
  OAI22_X1 U15861 ( .A1(n7794), .A2(keyinput53), .B1(n11875), .B2(keyinput74), 
        .ZN(n13780) );
  AOI221_X1 U15862 ( .B1(n7794), .B2(keyinput53), .C1(keyinput74), .C2(n11875), 
        .A(n13780), .ZN(n13781) );
  NAND3_X1 U15863 ( .A1(n13783), .A2(n13782), .A3(n13781), .ZN(n13784) );
  NOR4_X1 U15864 ( .A1(n13787), .A2(n13786), .A3(n13785), .A4(n13784), .ZN(
        n13806) );
  AOI211_X1 U15865 ( .C1(n13801), .C2(n13789), .A(n13925), .B(n13788), .ZN(
        n13793) );
  OAI22_X1 U15866 ( .A1(n13791), .A2(n13928), .B1(n13790), .B2(n14784), .ZN(
        n13792) );
  NOR2_X1 U15867 ( .A1(n13793), .A2(n13792), .ZN(n13992) );
  INV_X1 U15868 ( .A(n13794), .ZN(n13795) );
  AOI211_X1 U15869 ( .C1(n13990), .C2(n13814), .A(n6611), .B(n13795), .ZN(
        n13989) );
  INV_X1 U15870 ( .A(n13796), .ZN(n13797) );
  AOI22_X1 U15871 ( .A1(n15059), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n15058), 
        .B2(n13797), .ZN(n13798) );
  OAI21_X1 U15872 ( .B1(n13799), .B2(n13959), .A(n13798), .ZN(n13800) );
  AOI21_X1 U15873 ( .B1(n13989), .B2(n15068), .A(n13800), .ZN(n13804) );
  XNOR2_X1 U15874 ( .A(n13802), .B(n13801), .ZN(n13993) );
  OAI211_X1 U15875 ( .C1(n13992), .C2(n15072), .A(n13804), .B(n13803), .ZN(
        n13805) );
  XOR2_X1 U15876 ( .A(n13806), .B(n13805), .Z(P2_U3239) );
  XNOR2_X1 U15877 ( .A(n13807), .B(n13811), .ZN(n13809) );
  AOI21_X1 U15878 ( .B1(n13809), .B2(n15054), .A(n13808), .ZN(n13997) );
  OAI21_X1 U15879 ( .B1(n13812), .B2(n13811), .A(n13810), .ZN(n13998) );
  INV_X1 U15880 ( .A(n13998), .ZN(n13821) );
  OR2_X1 U15881 ( .A1(n13829), .A2(n13819), .ZN(n13813) );
  AND3_X1 U15882 ( .A1(n13814), .A2(n13813), .A3(n11374), .ZN(n13994) );
  NAND2_X1 U15883 ( .A1(n13994), .A2(n15068), .ZN(n13818) );
  INV_X1 U15884 ( .A(n13815), .ZN(n13816) );
  AOI22_X1 U15885 ( .A1(n15072), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n15058), 
        .B2(n13816), .ZN(n13817) );
  OAI211_X1 U15886 ( .C1(n13819), .C2(n13959), .A(n13818), .B(n13817), .ZN(
        n13820) );
  AOI21_X1 U15887 ( .B1(n13821), .B2(n15069), .A(n13820), .ZN(n13822) );
  OAI21_X1 U15888 ( .B1(n15059), .B2(n13997), .A(n13822), .ZN(P2_U3240) );
  XNOR2_X1 U15889 ( .A(n13824), .B(n13823), .ZN(n13826) );
  AOI21_X1 U15890 ( .B1(n13826), .B2(n15054), .A(n13825), .ZN(n14001) );
  OAI21_X1 U15891 ( .B1(n13847), .B2(n13827), .A(n11374), .ZN(n13828) );
  NAND2_X1 U15892 ( .A1(n13999), .A2(n15060), .ZN(n13833) );
  INV_X1 U15893 ( .A(n13830), .ZN(n13831) );
  AOI22_X1 U15894 ( .A1(n15072), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n15058), 
        .B2(n13831), .ZN(n13832) );
  NAND2_X1 U15895 ( .A1(n13833), .A2(n13832), .ZN(n13838) );
  OAI21_X1 U15896 ( .B1(n13836), .B2(n13835), .A(n13834), .ZN(n14002) );
  NOR2_X1 U15897 ( .A1(n14002), .A2(n13941), .ZN(n13837) );
  AOI211_X1 U15898 ( .C1(n7593), .C2(n15068), .A(n13838), .B(n13837), .ZN(
        n13839) );
  OAI21_X1 U15899 ( .B1(n15059), .B2(n14001), .A(n13839), .ZN(P2_U3241) );
  XNOR2_X1 U15900 ( .A(n13840), .B(n13841), .ZN(n14007) );
  XNOR2_X1 U15901 ( .A(n13842), .B(n13841), .ZN(n13844) );
  AOI21_X1 U15902 ( .B1(n13844), .B2(n15054), .A(n13843), .ZN(n14006) );
  OAI21_X1 U15903 ( .B1(n13845), .B2(n13957), .A(n14006), .ZN(n13846) );
  NAND2_X1 U15904 ( .A1(n13846), .A2(n13944), .ZN(n13853) );
  INV_X1 U15905 ( .A(n13861), .ZN(n13848) );
  AOI211_X1 U15906 ( .C1(n14004), .C2(n13848), .A(n6611), .B(n13847), .ZN(
        n14003) );
  INV_X1 U15907 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n13849) );
  OAI22_X1 U15908 ( .A1(n13850), .A2(n13959), .B1(n13944), .B2(n13849), .ZN(
        n13851) );
  AOI21_X1 U15909 ( .B1(n14003), .B2(n15068), .A(n13851), .ZN(n13852) );
  OAI211_X1 U15910 ( .C1(n14007), .C2(n13941), .A(n13853), .B(n13852), .ZN(
        P2_U3242) );
  AOI211_X1 U15911 ( .C1(n13867), .C2(n13855), .A(n13925), .B(n13854), .ZN(
        n13858) );
  INV_X1 U15912 ( .A(n13856), .ZN(n13857) );
  NOR2_X1 U15913 ( .A1(n13858), .A2(n13857), .ZN(n14012) );
  NAND2_X1 U15914 ( .A1(n6723), .A2(n14010), .ZN(n13859) );
  NAND2_X1 U15915 ( .A1(n13859), .A2(n15065), .ZN(n13860) );
  NOR2_X1 U15916 ( .A1(n13861), .A2(n13860), .ZN(n14009) );
  NAND2_X1 U15917 ( .A1(n14010), .A2(n15060), .ZN(n13865) );
  INV_X1 U15918 ( .A(n13862), .ZN(n13863) );
  AOI22_X1 U15919 ( .A1(n15072), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n15058), 
        .B2(n13863), .ZN(n13864) );
  NAND2_X1 U15920 ( .A1(n13865), .A2(n13864), .ZN(n13866) );
  AOI21_X1 U15921 ( .B1(n14009), .B2(n15068), .A(n13866), .ZN(n13871) );
  INV_X1 U15922 ( .A(n14014), .ZN(n13869) );
  OR2_X1 U15923 ( .A1(n13868), .A2(n13867), .ZN(n14008) );
  NAND3_X1 U15924 ( .A1(n13869), .A2(n15069), .A3(n14008), .ZN(n13870) );
  OAI211_X1 U15925 ( .C1(n14012), .C2(n15059), .A(n13871), .B(n13870), .ZN(
        P2_U3243) );
  OR3_X1 U15926 ( .A1(n13888), .A2(n13872), .A3(n13878), .ZN(n13873) );
  NAND2_X1 U15927 ( .A1(n13874), .A2(n13873), .ZN(n13876) );
  AOI222_X1 U15928 ( .A1(n15054), .A2(n13876), .B1(n13907), .B2(n14787), .C1(
        n13875), .C2(n13949), .ZN(n14018) );
  AOI21_X1 U15929 ( .B1(n13878), .B2(n13877), .A(n6744), .ZN(n14019) );
  INV_X1 U15930 ( .A(n14019), .ZN(n13886) );
  AOI21_X1 U15931 ( .B1(n14016), .B2(n13879), .A(n6611), .ZN(n13880) );
  AND2_X1 U15932 ( .A1(n13880), .A2(n6723), .ZN(n14015) );
  NAND2_X1 U15933 ( .A1(n14015), .A2(n15068), .ZN(n13883) );
  AOI22_X1 U15934 ( .A1(n13881), .A2(n15058), .B1(P2_REG2_REG_21__SCAN_IN), 
        .B2(n15059), .ZN(n13882) );
  OAI211_X1 U15935 ( .C1(n13884), .C2(n13959), .A(n13883), .B(n13882), .ZN(
        n13885) );
  AOI21_X1 U15936 ( .B1(n13886), .B2(n15069), .A(n13885), .ZN(n13887) );
  OAI21_X1 U15937 ( .B1(n14018), .B2(n15059), .A(n13887), .ZN(P2_U3244) );
  AOI21_X1 U15938 ( .B1(n13893), .B2(n13889), .A(n13888), .ZN(n13890) );
  OAI222_X1 U15939 ( .A1(n14784), .A2(n13891), .B1(n13928), .B2(n13929), .C1(
        n13925), .C2(n13890), .ZN(n14020) );
  OAI21_X1 U15940 ( .B1(n13894), .B2(n13893), .A(n13892), .ZN(n14024) );
  OAI22_X1 U15941 ( .A1(n13896), .A2(n13957), .B1(n13895), .B2(n13944), .ZN(
        n13897) );
  AOI21_X1 U15942 ( .B1(n14022), .B2(n15060), .A(n13897), .ZN(n13900) );
  XNOR2_X1 U15943 ( .A(n14022), .B(n7071), .ZN(n13898) );
  AND2_X1 U15944 ( .A1(n13898), .A2(n11374), .ZN(n14021) );
  NAND2_X1 U15945 ( .A1(n14021), .A2(n15068), .ZN(n13899) );
  OAI211_X1 U15946 ( .C1(n14024), .C2(n13941), .A(n13900), .B(n13899), .ZN(
        n13901) );
  AOI21_X1 U15947 ( .B1(n14020), .B2(n13944), .A(n13901), .ZN(n13902) );
  INV_X1 U15948 ( .A(n13902), .ZN(P2_U3245) );
  OAI211_X1 U15949 ( .C1(n13905), .C2(n13904), .A(n13903), .B(n15054), .ZN(
        n13909) );
  AOI22_X1 U15950 ( .A1(n13907), .A2(n13949), .B1(n14787), .B2(n13906), .ZN(
        n13908) );
  NAND2_X1 U15951 ( .A1(n13909), .A2(n13908), .ZN(n14025) );
  AOI21_X1 U15952 ( .B1(n13930), .B2(n14027), .A(n6611), .ZN(n13911) );
  AND2_X1 U15953 ( .A1(n13911), .A2(n13910), .ZN(n14026) );
  NAND2_X1 U15954 ( .A1(n14026), .A2(n15068), .ZN(n13915) );
  INV_X1 U15955 ( .A(n13912), .ZN(n13913) );
  AOI22_X1 U15956 ( .A1(n13913), .A2(n15058), .B1(P2_REG2_REG_19__SCAN_IN), 
        .B2(n15059), .ZN(n13914) );
  OAI211_X1 U15957 ( .C1(n13916), .C2(n13959), .A(n13915), .B(n13914), .ZN(
        n13921) );
  OAI21_X1 U15958 ( .B1(n13919), .B2(n13918), .A(n13917), .ZN(n14029) );
  NOR2_X1 U15959 ( .A1(n14029), .A2(n13941), .ZN(n13920) );
  AOI211_X1 U15960 ( .C1(n13944), .C2(n14025), .A(n13921), .B(n13920), .ZN(
        n13922) );
  INV_X1 U15961 ( .A(n13922), .ZN(P2_U3246) );
  XNOR2_X1 U15962 ( .A(n13924), .B(n13923), .ZN(n13926) );
  OAI222_X1 U15963 ( .A1(n14784), .A2(n13929), .B1(n13928), .B2(n13927), .C1(
        n13926), .C2(n13925), .ZN(n14035) );
  OAI211_X1 U15964 ( .C1(n13932), .C2(n13931), .A(n15065), .B(n13930), .ZN(
        n14031) );
  INV_X1 U15965 ( .A(n13933), .ZN(n13934) );
  AOI22_X1 U15966 ( .A1(n13934), .A2(n15058), .B1(n15059), .B2(
        P2_REG2_REG_18__SCAN_IN), .ZN(n13936) );
  NAND2_X1 U15967 ( .A1(n14030), .A2(n15060), .ZN(n13935) );
  OAI211_X1 U15968 ( .C1(n14031), .C2(n13937), .A(n13936), .B(n13935), .ZN(
        n13943) );
  AOI21_X1 U15969 ( .B1(n13940), .B2(n13939), .A(n13938), .ZN(n14033) );
  NOR2_X1 U15970 ( .A1(n14033), .A2(n13941), .ZN(n13942) );
  AOI211_X1 U15971 ( .C1(n13944), .C2(n14035), .A(n13943), .B(n13942), .ZN(
        n13945) );
  INV_X1 U15972 ( .A(n13945), .ZN(P2_U3247) );
  OAI21_X1 U15973 ( .B1(n13947), .B2(n13961), .A(n13946), .ZN(n13951) );
  AOI222_X1 U15974 ( .A1(n15054), .A2(n13951), .B1(n13950), .B2(n13949), .C1(
        n13948), .C2(n14787), .ZN(n15111) );
  MUX2_X1 U15975 ( .A(n13952), .B(n15111), .S(n13944), .Z(n13965) );
  INV_X1 U15976 ( .A(n13953), .ZN(n13954) );
  AOI211_X1 U15977 ( .C1(n15106), .C2(n13955), .A(n6611), .B(n13954), .ZN(
        n15105) );
  OAI22_X1 U15978 ( .A1(n13959), .A2(n13958), .B1(n13957), .B2(n13956), .ZN(
        n13960) );
  AOI21_X1 U15979 ( .B1(n15105), .B2(n15068), .A(n13960), .ZN(n13964) );
  NAND2_X1 U15980 ( .A1(n13962), .A2(n13961), .ZN(n15107) );
  NAND3_X1 U15981 ( .A1(n15108), .A2(n15069), .A3(n15107), .ZN(n13963) );
  NAND3_X1 U15982 ( .A1(n13965), .A2(n13964), .A3(n13963), .ZN(P2_U3261) );
  INV_X1 U15983 ( .A(n13966), .ZN(n13968) );
  OAI211_X1 U15984 ( .C1(n13968), .C2(n15150), .A(n13967), .B(n13969), .ZN(
        n14051) );
  MUX2_X1 U15985 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n14051), .S(n15177), .Z(
        P2_U3530) );
  OAI211_X1 U15986 ( .C1(n7082), .C2(n15150), .A(n13970), .B(n13969), .ZN(
        n14052) );
  MUX2_X1 U15987 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n14052), .S(n15177), .Z(
        P2_U3529) );
  NAND2_X1 U15988 ( .A1(n10171), .A2(n13971), .ZN(n15147) );
  NAND2_X1 U15989 ( .A1(n13972), .A2(n15147), .ZN(n13978) );
  INV_X1 U15990 ( .A(n13973), .ZN(n13977) );
  OAI21_X1 U15991 ( .B1(n7083), .B2(n15150), .A(n13974), .ZN(n13975) );
  NAND3_X1 U15992 ( .A1(n13978), .A2(n13977), .A3(n13976), .ZN(n14053) );
  MUX2_X1 U15993 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n14053), .S(n15177), .Z(
        P2_U3528) );
  AOI21_X1 U15994 ( .B1(n15114), .B2(n13980), .A(n13979), .ZN(n13981) );
  MUX2_X1 U15995 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n14054), .S(n15177), .Z(
        P2_U3527) );
  AOI21_X1 U15996 ( .B1(n15114), .B2(n13985), .A(n13984), .ZN(n13986) );
  OAI211_X1 U15997 ( .C1(n13988), .C2(n15117), .A(n13987), .B(n13986), .ZN(
        n14055) );
  MUX2_X1 U15998 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n14055), .S(n15177), .Z(
        P2_U3526) );
  AOI21_X1 U15999 ( .B1(n15114), .B2(n13990), .A(n13989), .ZN(n13991) );
  OAI211_X1 U16000 ( .C1(n15117), .C2(n13993), .A(n13992), .B(n13991), .ZN(
        n14056) );
  MUX2_X1 U16001 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14056), .S(n15177), .Z(
        P2_U3525) );
  AOI21_X1 U16002 ( .B1(n15114), .B2(n13995), .A(n13994), .ZN(n13996) );
  OAI211_X1 U16003 ( .C1(n13998), .C2(n15117), .A(n13997), .B(n13996), .ZN(
        n14057) );
  MUX2_X1 U16004 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n14057), .S(n15177), .Z(
        P2_U3524) );
  AOI21_X1 U16005 ( .B1(n15114), .B2(n13999), .A(n7593), .ZN(n14000) );
  OAI211_X1 U16006 ( .C1(n14002), .C2(n15117), .A(n14001), .B(n14000), .ZN(
        n14058) );
  MUX2_X1 U16007 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14058), .S(n15177), .Z(
        P2_U3523) );
  AOI21_X1 U16008 ( .B1(n15114), .B2(n14004), .A(n14003), .ZN(n14005) );
  OAI211_X1 U16009 ( .C1(n14007), .C2(n15117), .A(n14006), .B(n14005), .ZN(
        n14059) );
  MUX2_X1 U16010 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14059), .S(n15177), .Z(
        P2_U3522) );
  NAND2_X1 U16011 ( .A1(n14008), .A2(n15147), .ZN(n14013) );
  AOI21_X1 U16012 ( .B1(n15114), .B2(n14010), .A(n14009), .ZN(n14011) );
  OAI211_X1 U16013 ( .C1(n14014), .C2(n14013), .A(n14012), .B(n14011), .ZN(
        n14060) );
  MUX2_X1 U16014 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n14060), .S(n15177), .Z(
        P2_U3521) );
  AOI21_X1 U16015 ( .B1(n15114), .B2(n14016), .A(n14015), .ZN(n14017) );
  OAI211_X1 U16016 ( .C1(n15117), .C2(n14019), .A(n14018), .B(n14017), .ZN(
        n14061) );
  MUX2_X1 U16017 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n14061), .S(n15177), .Z(
        P2_U3520) );
  AOI211_X1 U16018 ( .C1(n15114), .C2(n14022), .A(n14021), .B(n14020), .ZN(
        n14023) );
  OAI21_X1 U16019 ( .B1(n15117), .B2(n14024), .A(n14023), .ZN(n14062) );
  MUX2_X1 U16020 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14062), .S(n15177), .Z(
        P2_U3519) );
  AOI211_X1 U16021 ( .C1(n15114), .C2(n14027), .A(n14026), .B(n14025), .ZN(
        n14028) );
  OAI21_X1 U16022 ( .B1(n15117), .B2(n14029), .A(n14028), .ZN(n14063) );
  MUX2_X1 U16023 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n14063), .S(n15177), .Z(
        P2_U3518) );
  NAND2_X1 U16024 ( .A1(n14030), .A2(n15114), .ZN(n14032) );
  OAI211_X1 U16025 ( .C1(n14033), .C2(n15117), .A(n14032), .B(n14031), .ZN(
        n14034) );
  OR2_X1 U16026 ( .A1(n14035), .A2(n14034), .ZN(n14064) );
  MUX2_X1 U16027 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14064), .S(n15177), .Z(
        P2_U3517) );
  AOI21_X1 U16028 ( .B1(n15114), .B2(n14037), .A(n14036), .ZN(n14038) );
  OAI211_X1 U16029 ( .C1(n15117), .C2(n14040), .A(n14039), .B(n14038), .ZN(
        n14065) );
  MUX2_X1 U16030 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n14065), .S(n15177), .Z(
        P2_U3516) );
  AOI21_X1 U16031 ( .B1(n15114), .B2(n14042), .A(n14041), .ZN(n14043) );
  OAI211_X1 U16032 ( .C1(n15117), .C2(n14045), .A(n14044), .B(n14043), .ZN(
        n14066) );
  MUX2_X1 U16033 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14066), .S(n15177), .Z(
        P2_U3515) );
  AOI211_X1 U16034 ( .C1(n15114), .C2(n14048), .A(n14047), .B(n14046), .ZN(
        n14049) );
  OAI21_X1 U16035 ( .B1(n15117), .B2(n14050), .A(n14049), .ZN(n14067) );
  MUX2_X1 U16036 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n14067), .S(n15177), .Z(
        P2_U3514) );
  MUX2_X1 U16037 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n14051), .S(n15157), .Z(
        P2_U3498) );
  MUX2_X1 U16038 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n14052), .S(n15157), .Z(
        P2_U3497) );
  MUX2_X1 U16039 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n14053), .S(n15157), .Z(
        P2_U3496) );
  MUX2_X1 U16040 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n14054), .S(n15157), .Z(
        P2_U3495) );
  MUX2_X1 U16041 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n14055), .S(n15157), .Z(
        P2_U3494) );
  MUX2_X1 U16042 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14056), .S(n15157), .Z(
        P2_U3493) );
  MUX2_X1 U16043 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n14057), .S(n15157), .Z(
        P2_U3492) );
  MUX2_X1 U16044 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14058), .S(n15157), .Z(
        P2_U3491) );
  MUX2_X1 U16045 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14059), .S(n15157), .Z(
        P2_U3490) );
  MUX2_X1 U16046 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n14060), .S(n15157), .Z(
        P2_U3489) );
  MUX2_X1 U16047 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n14061), .S(n15157), .Z(
        P2_U3488) );
  MUX2_X1 U16048 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14062), .S(n15157), .Z(
        P2_U3487) );
  MUX2_X1 U16049 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n14063), .S(n15157), .Z(
        P2_U3486) );
  MUX2_X1 U16050 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14064), .S(n15157), .Z(
        P2_U3484) );
  MUX2_X1 U16051 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n14065), .S(n15157), .Z(
        P2_U3481) );
  MUX2_X1 U16052 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n14066), .S(n15157), .Z(
        P2_U3478) );
  MUX2_X1 U16053 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n14067), .S(n15157), .Z(
        P2_U3475) );
  INV_X1 U16054 ( .A(n14068), .ZN(n14669) );
  NOR4_X1 U16055 ( .A1(n14069), .A2(P2_IR_REG_30__SCAN_IN), .A3(n6642), .A4(
        P2_U3088), .ZN(n14070) );
  AOI21_X1 U16056 ( .B1(n14071), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n14070), 
        .ZN(n14072) );
  OAI21_X1 U16057 ( .B1(n14669), .B2(n6618), .A(n14072), .ZN(P2_U3296) );
  INV_X1 U16058 ( .A(n14073), .ZN(n14074) );
  MUX2_X1 U16059 ( .A(n14074), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  OAI211_X1 U16060 ( .C1(n14077), .C2(n14076), .A(n14075), .B(n14904), .ZN(
        n14082) );
  AOI22_X1 U16061 ( .A1(n14228), .A2(n14078), .B1(P1_REG3_REG_7__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14081) );
  AOI22_X1 U16062 ( .A1(n14194), .A2(n14247), .B1(n14193), .B2(n14245), .ZN(
        n14080) );
  NAND2_X1 U16063 ( .A1(n14215), .A2(n14954), .ZN(n14079) );
  NAND4_X1 U16064 ( .A1(n14082), .A2(n14081), .A3(n14080), .A4(n14079), .ZN(
        P1_U3213) );
  INV_X1 U16065 ( .A(n14084), .ZN(n14369) );
  OAI22_X1 U16066 ( .A1(n14909), .A2(n14369), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14085), .ZN(n14088) );
  OAI22_X1 U16067 ( .A1(n11965), .A2(n14899), .B1(n14900), .B2(n14086), .ZN(
        n14087) );
  AOI211_X1 U16068 ( .C1(n14567), .C2(n14215), .A(n14088), .B(n14087), .ZN(
        n14089) );
  INV_X1 U16069 ( .A(n14090), .ZN(n14091) );
  AOI21_X1 U16070 ( .B1(n14093), .B2(n14092), .A(n14091), .ZN(n14101) );
  OAI22_X1 U16071 ( .A1(n14095), .A2(n14899), .B1(n14900), .B2(n14094), .ZN(
        n14096) );
  AOI211_X1 U16072 ( .C1(n14228), .C2(n14098), .A(n14097), .B(n14096), .ZN(
        n14100) );
  NAND2_X1 U16073 ( .A1(n14639), .A2(n14215), .ZN(n14099) );
  OAI211_X1 U16074 ( .C1(n14101), .C2(n14850), .A(n14100), .B(n14099), .ZN(
        P1_U3215) );
  NAND2_X1 U16075 ( .A1(n14188), .A2(n14104), .ZN(n14105) );
  XOR2_X1 U16076 ( .A(n14106), .B(n14105), .Z(n14114) );
  OR2_X1 U16077 ( .A1(n14467), .A2(n14438), .ZN(n14108) );
  NAND2_X1 U16078 ( .A1(n14235), .A2(n14540), .ZN(n14107) );
  NAND2_X1 U16079 ( .A1(n14108), .A2(n14107), .ZN(n14420) );
  INV_X1 U16080 ( .A(n14424), .ZN(n14110) );
  OAI22_X1 U16081 ( .A1(n14909), .A2(n14110), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14109), .ZN(n14111) );
  AOI21_X1 U16082 ( .B1(n14420), .B2(n14855), .A(n14111), .ZN(n14113) );
  INV_X1 U16083 ( .A(n14423), .ZN(n14426) );
  NOR2_X1 U16084 ( .A1(n14426), .A2(n14947), .ZN(n14592) );
  NAND2_X1 U16085 ( .A1(n14592), .A2(n14844), .ZN(n14112) );
  OAI211_X1 U16086 ( .C1(n14114), .C2(n14850), .A(n14113), .B(n14112), .ZN(
        P1_U3216) );
  AOI22_X1 U16087 ( .A1(n14194), .A2(n14541), .B1(n14193), .B2(n14496), .ZN(
        n14115) );
  NAND2_X1 U16088 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14337)
         );
  OAI211_X1 U16089 ( .C1(n14909), .C2(n14499), .A(n14115), .B(n14337), .ZN(
        n14119) );
  AOI211_X1 U16090 ( .C1(n14117), .C2(n14116), .A(n14850), .B(n6738), .ZN(
        n14118) );
  AOI211_X1 U16091 ( .C1(n14215), .C2(n14616), .A(n14119), .B(n14118), .ZN(
        n14120) );
  INV_X1 U16092 ( .A(n14120), .ZN(P1_U3219) );
  OAI21_X1 U16093 ( .B1(n14123), .B2(n14122), .A(n14121), .ZN(n14124) );
  NAND2_X1 U16094 ( .A1(n14124), .A2(n14904), .ZN(n14129) );
  AOI22_X1 U16095 ( .A1(n14194), .A2(n6609), .B1(n14215), .B2(n14125), .ZN(
        n14128) );
  AOI22_X1 U16096 ( .A1(n14193), .A2(n14251), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n14126), .ZN(n14127) );
  NAND3_X1 U16097 ( .A1(n14129), .A2(n14128), .A3(n14127), .ZN(P1_U3222) );
  INV_X1 U16098 ( .A(n14186), .ZN(n14130) );
  AOI21_X1 U16099 ( .B1(n14131), .B2(n14102), .A(n14130), .ZN(n14138) );
  OAI22_X1 U16100 ( .A1(n14133), .A2(n14909), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14132), .ZN(n14136) );
  OAI22_X1 U16101 ( .A1(n14467), .A2(n14899), .B1(n14134), .B2(n14900), .ZN(
        n14135) );
  AOI211_X1 U16102 ( .C1(n6970), .C2(n14215), .A(n14136), .B(n14135), .ZN(
        n14137) );
  OAI21_X1 U16103 ( .B1(n14138), .B2(n14850), .A(n14137), .ZN(P1_U3223) );
  XOR2_X1 U16104 ( .A(n14140), .B(n14139), .Z(n14147) );
  NAND2_X1 U16105 ( .A1(n14235), .A2(n14539), .ZN(n14142) );
  NAND2_X1 U16106 ( .A1(n14361), .A2(n14540), .ZN(n14141) );
  NAND2_X1 U16107 ( .A1(n14142), .A2(n14141), .ZN(n14577) );
  AOI22_X1 U16108 ( .A1(n14855), .A2(n14577), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14143) );
  OAI21_X1 U16109 ( .B1(n14144), .B2(n14909), .A(n14143), .ZN(n14145) );
  AOI21_X1 U16110 ( .B1(n14578), .B2(n14215), .A(n14145), .ZN(n14146) );
  OAI21_X1 U16111 ( .B1(n14147), .B2(n14850), .A(n14146), .ZN(P1_U3225) );
  XOR2_X1 U16112 ( .A(n14148), .B(n6726), .Z(n14155) );
  AOI22_X1 U16113 ( .A1(n14193), .A2(n14517), .B1(n14194), .B2(n14238), .ZN(
        n14150) );
  OAI211_X1 U16114 ( .C1(n14909), .C2(n14151), .A(n14150), .B(n14149), .ZN(
        n14152) );
  AOI21_X1 U16115 ( .B1(n14153), .B2(n14215), .A(n14152), .ZN(n14154) );
  OAI21_X1 U16116 ( .B1(n14155), .B2(n14850), .A(n14154), .ZN(P1_U3226) );
  XOR2_X1 U16117 ( .A(n14157), .B(n14156), .Z(n14161) );
  AOI22_X1 U16118 ( .A1(n14193), .A2(n14541), .B1(n14194), .B2(n14538), .ZN(
        n14158) );
  NAND2_X1 U16119 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14294)
         );
  OAI211_X1 U16120 ( .C1(n14909), .C2(n14547), .A(n14158), .B(n14294), .ZN(
        n14159) );
  AOI21_X1 U16121 ( .B1(n14550), .B2(n14215), .A(n14159), .ZN(n14160) );
  OAI21_X1 U16122 ( .B1(n14161), .B2(n14850), .A(n14160), .ZN(P1_U3228) );
  OR2_X1 U16123 ( .A1(n14102), .A2(n14162), .ZN(n14164) );
  NAND2_X1 U16124 ( .A1(n14164), .A2(n14163), .ZN(n14165) );
  XOR2_X1 U16125 ( .A(n14166), .B(n14165), .Z(n14173) );
  INV_X1 U16126 ( .A(n14414), .ZN(n14168) );
  OAI22_X1 U16127 ( .A1(n14909), .A2(n14168), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14167), .ZN(n14171) );
  OAI22_X1 U16128 ( .A1(n14210), .A2(n14899), .B1(n14900), .B2(n14169), .ZN(
        n14170) );
  AOI211_X1 U16129 ( .C1(n14585), .C2(n14215), .A(n14171), .B(n14170), .ZN(
        n14172) );
  OAI21_X1 U16130 ( .B1(n14173), .B2(n14850), .A(n14172), .ZN(P1_U3229) );
  OAI211_X1 U16131 ( .C1(n14176), .C2(n14175), .A(n14174), .B(n14904), .ZN(
        n14184) );
  INV_X1 U16132 ( .A(n14177), .ZN(n14482) );
  OR2_X1 U16133 ( .A1(n14439), .A2(n14466), .ZN(n14179) );
  NAND2_X1 U16134 ( .A1(n14518), .A2(n14539), .ZN(n14178) );
  AND2_X1 U16135 ( .A1(n14179), .A2(n14178), .ZN(n14478) );
  OAI22_X1 U16136 ( .A1(n14478), .A2(n14181), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14180), .ZN(n14182) );
  AOI21_X1 U16137 ( .B1(n14482), .B2(n14228), .A(n14182), .ZN(n14183) );
  OAI211_X1 U16138 ( .C1(n14484), .C2(n14896), .A(n14184), .B(n14183), .ZN(
        P1_U3233) );
  NAND2_X1 U16139 ( .A1(n14186), .A2(n14185), .ZN(n14190) );
  AND2_X1 U16140 ( .A1(n14188), .A2(n14187), .ZN(n14189) );
  OAI21_X1 U16141 ( .B1(n14191), .B2(n14190), .A(n14189), .ZN(n14192) );
  NAND2_X1 U16142 ( .A1(n14192), .A2(n14904), .ZN(n14198) );
  AOI22_X1 U16143 ( .A1(n14437), .A2(n14228), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14197) );
  AOI22_X1 U16144 ( .A1(n14237), .A2(n14194), .B1(n14193), .B2(n14440), .ZN(
        n14196) );
  NAND2_X1 U16145 ( .A1(n14599), .A2(n14215), .ZN(n14195) );
  NAND4_X1 U16146 ( .A1(n14198), .A2(n14197), .A3(n14196), .A4(n14195), .ZN(
        P1_U3235) );
  XOR2_X1 U16147 ( .A(n14200), .B(n14199), .Z(n14207) );
  NOR2_X1 U16148 ( .A1(n14201), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14315) );
  OAI22_X1 U16149 ( .A1(n14203), .A2(n14900), .B1(n14899), .B2(n14202), .ZN(
        n14204) );
  AOI211_X1 U16150 ( .C1(n14228), .C2(n14525), .A(n14315), .B(n14204), .ZN(
        n14206) );
  NAND2_X1 U16151 ( .A1(n14620), .A2(n14215), .ZN(n14205) );
  OAI211_X1 U16152 ( .C1(n14207), .C2(n14850), .A(n14206), .B(n14205), .ZN(
        P1_U3238) );
  XOR2_X1 U16153 ( .A(n14209), .B(n14208), .Z(n14217) );
  INV_X1 U16154 ( .A(n14377), .ZN(n14213) );
  OAI22_X1 U16155 ( .A1(n14211), .A2(n14466), .B1(n14210), .B2(n14438), .ZN(
        n14374) );
  AOI22_X1 U16156 ( .A1(n14855), .A2(n14374), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14212) );
  OAI21_X1 U16157 ( .B1(n14213), .B2(n14909), .A(n14212), .ZN(n14214) );
  AOI21_X1 U16158 ( .B1(n14572), .B2(n14215), .A(n14214), .ZN(n14216) );
  OAI21_X1 U16159 ( .B1(n14217), .B2(n14850), .A(n14216), .ZN(P1_U3240) );
  OAI21_X1 U16160 ( .B1(n14220), .B2(n14219), .A(n14218), .ZN(n14221) );
  NAND2_X1 U16161 ( .A1(n14221), .A2(n14904), .ZN(n14230) );
  INV_X1 U16162 ( .A(n14222), .ZN(n14227) );
  NAND2_X1 U16163 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14924)
         );
  INV_X1 U16164 ( .A(n14924), .ZN(n14226) );
  OAI22_X1 U16165 ( .A1(n14224), .A2(n14899), .B1(n14900), .B2(n14223), .ZN(
        n14225) );
  AOI211_X1 U16166 ( .C1(n14228), .C2(n14227), .A(n14226), .B(n14225), .ZN(
        n14229) );
  OAI211_X1 U16167 ( .C1(n14231), .C2(n14896), .A(n14230), .B(n14229), .ZN(
        P1_U3241) );
  MUX2_X1 U16168 ( .A(n14341), .B(P1_DATAO_REG_31__SCAN_IN), .S(n14252), .Z(
        P1_U3591) );
  MUX2_X1 U16169 ( .A(n14232), .B(P1_DATAO_REG_30__SCAN_IN), .S(n14252), .Z(
        P1_U3590) );
  MUX2_X1 U16170 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14233), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16171 ( .A(n14362), .B(P1_DATAO_REG_28__SCAN_IN), .S(n14252), .Z(
        P1_U3588) );
  MUX2_X1 U16172 ( .A(n14234), .B(P1_DATAO_REG_27__SCAN_IN), .S(n14252), .Z(
        P1_U3587) );
  MUX2_X1 U16173 ( .A(n14361), .B(P1_DATAO_REG_26__SCAN_IN), .S(n14252), .Z(
        P1_U3586) );
  MUX2_X1 U16174 ( .A(n14404), .B(P1_DATAO_REG_25__SCAN_IN), .S(n14252), .Z(
        P1_U3585) );
  MUX2_X1 U16175 ( .A(n14235), .B(P1_DATAO_REG_24__SCAN_IN), .S(n14252), .Z(
        P1_U3584) );
  MUX2_X1 U16176 ( .A(n14440), .B(P1_DATAO_REG_23__SCAN_IN), .S(n14252), .Z(
        P1_U3583) );
  MUX2_X1 U16177 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14236), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16178 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14237), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16179 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14496), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16180 ( .A(n14518), .B(P1_DATAO_REG_19__SCAN_IN), .S(n14252), .Z(
        P1_U3579) );
  MUX2_X1 U16181 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14541), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16182 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14517), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16183 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14538), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U16184 ( .A(n14238), .B(P1_DATAO_REG_15__SCAN_IN), .S(n14252), .Z(
        P1_U3575) );
  MUX2_X1 U16185 ( .A(n14239), .B(P1_DATAO_REG_14__SCAN_IN), .S(n14252), .Z(
        P1_U3574) );
  MUX2_X1 U16186 ( .A(n14240), .B(P1_DATAO_REG_13__SCAN_IN), .S(n14252), .Z(
        P1_U3573) );
  MUX2_X1 U16187 ( .A(n14241), .B(P1_DATAO_REG_12__SCAN_IN), .S(n14252), .Z(
        P1_U3572) );
  MUX2_X1 U16188 ( .A(n14242), .B(P1_DATAO_REG_11__SCAN_IN), .S(n14252), .Z(
        P1_U3571) );
  MUX2_X1 U16189 ( .A(n14243), .B(P1_DATAO_REG_10__SCAN_IN), .S(n14252), .Z(
        P1_U3570) );
  MUX2_X1 U16190 ( .A(n14244), .B(P1_DATAO_REG_9__SCAN_IN), .S(n14252), .Z(
        P1_U3569) );
  MUX2_X1 U16191 ( .A(n14245), .B(P1_DATAO_REG_8__SCAN_IN), .S(n14252), .Z(
        P1_U3568) );
  MUX2_X1 U16192 ( .A(n14246), .B(P1_DATAO_REG_7__SCAN_IN), .S(n14252), .Z(
        P1_U3567) );
  MUX2_X1 U16193 ( .A(n14247), .B(P1_DATAO_REG_6__SCAN_IN), .S(n14252), .Z(
        P1_U3566) );
  MUX2_X1 U16194 ( .A(n14248), .B(P1_DATAO_REG_5__SCAN_IN), .S(n14252), .Z(
        P1_U3565) );
  MUX2_X1 U16195 ( .A(n14249), .B(P1_DATAO_REG_4__SCAN_IN), .S(n14252), .Z(
        P1_U3564) );
  MUX2_X1 U16196 ( .A(n14250), .B(P1_DATAO_REG_3__SCAN_IN), .S(n14252), .Z(
        P1_U3563) );
  MUX2_X1 U16197 ( .A(n14251), .B(P1_DATAO_REG_2__SCAN_IN), .S(n14252), .Z(
        P1_U3562) );
  MUX2_X1 U16198 ( .A(n10246), .B(P1_DATAO_REG_1__SCAN_IN), .S(n14252), .Z(
        P1_U3561) );
  MUX2_X1 U16199 ( .A(n6609), .B(P1_DATAO_REG_0__SCAN_IN), .S(n14252), .Z(
        P1_U3560) );
  MUX2_X1 U16200 ( .A(n14255), .B(n14254), .S(n6684), .Z(n14257) );
  NAND2_X1 U16201 ( .A1(n14257), .A2(n14256), .ZN(n14258) );
  OAI211_X1 U16202 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n14259), .A(n14258), .B(
        P1_U4016), .ZN(n14290) );
  AOI22_X1 U16203 ( .A1(n14316), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n14273) );
  AOI211_X1 U16204 ( .C1(n14262), .C2(n14261), .A(n14260), .B(n14298), .ZN(
        n14269) );
  MUX2_X1 U16205 ( .A(n10592), .B(P1_REG2_REG_2__SCAN_IN), .S(n14270), .Z(
        n14265) );
  NAND3_X1 U16206 ( .A1(n14265), .A2(n14264), .A3(n14263), .ZN(n14266) );
  AND3_X1 U16207 ( .A1(n14332), .A2(n14267), .A3(n14266), .ZN(n14268) );
  NOR2_X1 U16208 ( .A1(n14269), .A2(n14268), .ZN(n14272) );
  NAND2_X1 U16209 ( .A1(n14303), .A2(n14270), .ZN(n14271) );
  NAND4_X1 U16210 ( .A1(n14290), .A2(n14273), .A3(n14272), .A4(n14271), .ZN(
        P1_U3245) );
  NOR2_X1 U16211 ( .A1(n14926), .A2(n14274), .ZN(n14275) );
  AOI211_X1 U16212 ( .C1(n14303), .C2(n14281), .A(n14276), .B(n14275), .ZN(
        n14289) );
  AOI211_X1 U16213 ( .C1(n14279), .C2(n14278), .A(n14277), .B(n14298), .ZN(
        n14280) );
  INV_X1 U16214 ( .A(n14280), .ZN(n14288) );
  MUX2_X1 U16215 ( .A(n9837), .B(P1_REG2_REG_4__SCAN_IN), .S(n14281), .Z(
        n14282) );
  NAND3_X1 U16216 ( .A1(n14284), .A2(n14283), .A3(n14282), .ZN(n14285) );
  NAND3_X1 U16217 ( .A1(n14332), .A2(n14286), .A3(n14285), .ZN(n14287) );
  NAND4_X1 U16218 ( .A1(n14290), .A2(n14289), .A3(n14288), .A4(n14287), .ZN(
        P1_U3247) );
  AOI22_X1 U16219 ( .A1(n14292), .A2(n14291), .B1(P1_REG2_REG_16__SCAN_IN), 
        .B2(n14297), .ZN(n14293) );
  INV_X1 U16220 ( .A(n14293), .ZN(n14307) );
  XOR2_X1 U16221 ( .A(P1_REG2_REG_17__SCAN_IN), .B(n14310), .Z(n14306) );
  XNOR2_X1 U16222 ( .A(n14307), .B(n14306), .ZN(n14305) );
  INV_X1 U16223 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n14295) );
  OAI21_X1 U16224 ( .B1(n14926), .B2(n14295), .A(n14294), .ZN(n14302) );
  AOI21_X1 U16225 ( .B1(n14297), .B2(P1_REG1_REG_16__SCAN_IN), .A(n14296), 
        .ZN(n14300) );
  XNOR2_X1 U16226 ( .A(n14310), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n14299) );
  NOR2_X1 U16227 ( .A1(n14300), .A2(n14299), .ZN(n14309) );
  AOI211_X1 U16228 ( .C1(n14300), .C2(n14299), .A(n14298), .B(n14309), .ZN(
        n14301) );
  AOI211_X1 U16229 ( .C1(n14303), .C2(n14310), .A(n14302), .B(n14301), .ZN(
        n14304) );
  OAI21_X1 U16230 ( .B1(n14305), .B2(n14917), .A(n14304), .ZN(P1_U3260) );
  AOI22_X1 U16231 ( .A1(n14307), .A2(n14306), .B1(P1_REG2_REG_17__SCAN_IN), 
        .B2(n14310), .ZN(n14324) );
  XNOR2_X1 U16232 ( .A(n14324), .B(n14308), .ZN(n14325) );
  XNOR2_X1 U16233 ( .A(n14325), .B(P1_REG2_REG_18__SCAN_IN), .ZN(n14319) );
  AOI21_X1 U16234 ( .B1(n14310), .B2(P1_REG1_REG_17__SCAN_IN), .A(n14309), 
        .ZN(n14311) );
  NOR2_X1 U16235 ( .A1(n14311), .A2(n14323), .ZN(n14321) );
  INV_X1 U16236 ( .A(n14320), .ZN(n14312) );
  OAI211_X1 U16237 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n14313), .A(n14312), 
        .B(n14913), .ZN(n14318) );
  NOR2_X1 U16238 ( .A1(n14921), .A2(n14323), .ZN(n14314) );
  AOI211_X1 U16239 ( .C1(n14316), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n14315), 
        .B(n14314), .ZN(n14317) );
  OAI211_X1 U16240 ( .C1(n14319), .C2(n14917), .A(n14318), .B(n14317), .ZN(
        P1_U3261) );
  INV_X1 U16241 ( .A(n14333), .ZN(n14330) );
  OR2_X1 U16242 ( .A1(n14324), .A2(n14323), .ZN(n14327) );
  NAND2_X1 U16243 ( .A1(n14325), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n14326) );
  NAND2_X1 U16244 ( .A1(n14327), .A2(n14326), .ZN(n14328) );
  XOR2_X1 U16245 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n14328), .Z(n14331) );
  OAI21_X1 U16246 ( .B1(n14331), .B2(n14917), .A(n14921), .ZN(n14329) );
  AOI21_X1 U16247 ( .B1(n14330), .B2(n14913), .A(n14329), .ZN(n14336) );
  AOI22_X1 U16248 ( .A1(n14333), .A2(n14913), .B1(n14332), .B2(n14331), .ZN(
        n14335) );
  MUX2_X1 U16249 ( .A(n14336), .B(n14335), .S(n14334), .Z(n14338) );
  OAI211_X1 U16250 ( .C1(n6863), .C2(n14926), .A(n14338), .B(n14337), .ZN(
        P1_U3262) );
  NOR2_X1 U16251 ( .A1(n14345), .A2(n7601), .ZN(n14346) );
  XNOR2_X1 U16252 ( .A(n14346), .B(n14342), .ZN(n14339) );
  NAND2_X1 U16253 ( .A1(n14339), .A2(n14712), .ZN(n14554) );
  NAND2_X1 U16254 ( .A1(n14341), .A2(n14340), .ZN(n14556) );
  NOR2_X1 U16255 ( .A1(n14705), .A2(n14556), .ZN(n14350) );
  INV_X1 U16256 ( .A(n14342), .ZN(n14555) );
  NOR2_X1 U16257 ( .A1(n14555), .A2(n14506), .ZN(n14343) );
  AOI211_X1 U16258 ( .C1(n14526), .C2(P1_REG2_REG_31__SCAN_IN), .A(n14350), 
        .B(n14343), .ZN(n14344) );
  OAI21_X1 U16259 ( .B1(n14529), .B2(n14554), .A(n14344), .ZN(P1_U3263) );
  INV_X1 U16260 ( .A(n7601), .ZN(n14348) );
  INV_X1 U16261 ( .A(n14346), .ZN(n14347) );
  OAI211_X1 U16262 ( .C1(n14348), .C2(n14558), .A(n14347), .B(n14712), .ZN(
        n14557) );
  NOR2_X1 U16263 ( .A1(n14558), .A2(n14506), .ZN(n14349) );
  AOI211_X1 U16264 ( .C1(n14526), .C2(P1_REG2_REG_30__SCAN_IN), .A(n14350), 
        .B(n14349), .ZN(n14351) );
  OAI21_X1 U16265 ( .B1(n14529), .B2(n14557), .A(n14351), .ZN(P1_U3264) );
  NAND2_X1 U16266 ( .A1(n14376), .A2(n14567), .ZN(n14352) );
  NAND2_X1 U16267 ( .A1(n14352), .A2(n14712), .ZN(n14353) );
  INV_X1 U16268 ( .A(n14357), .ZN(n14355) );
  NAND2_X1 U16269 ( .A1(n14355), .A2(n14701), .ZN(n14360) );
  AOI22_X1 U16270 ( .A1(n14357), .A2(n14701), .B1(n14965), .B2(n14356), .ZN(
        n14359) );
  MUX2_X1 U16271 ( .A(n14360), .B(n14359), .S(n14358), .Z(n14367) );
  AOI22_X1 U16272 ( .A1(n14540), .A2(n14362), .B1(n14361), .B2(n14539), .ZN(
        n14363) );
  NAND2_X1 U16273 ( .A1(n14566), .A2(n14531), .ZN(n14372) );
  NAND2_X1 U16274 ( .A1(n14526), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n14368) );
  OAI21_X1 U16275 ( .B1(n14498), .B2(n14369), .A(n14368), .ZN(n14370) );
  AOI21_X1 U16276 ( .B1(n14567), .B2(n14706), .A(n14370), .ZN(n14371) );
  OAI211_X1 U16277 ( .C1(n14529), .C2(n14569), .A(n14372), .B(n14371), .ZN(
        P1_U3266) );
  XNOR2_X1 U16278 ( .A(n14373), .B(n14381), .ZN(n14375) );
  AOI21_X1 U16279 ( .B1(n14375), .B2(n14701), .A(n14374), .ZN(n14574) );
  AOI211_X1 U16280 ( .C1(n14572), .C2(n6732), .A(n14503), .B(n8854), .ZN(
        n14571) );
  AOI22_X1 U16281 ( .A1(n14526), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n14377), 
        .B2(n14703), .ZN(n14378) );
  OAI21_X1 U16282 ( .B1(n14379), .B2(n14506), .A(n14378), .ZN(n14384) );
  OAI21_X1 U16283 ( .B1(n14382), .B2(n14381), .A(n14380), .ZN(n14575) );
  NOR2_X1 U16284 ( .A1(n14575), .A2(n14511), .ZN(n14383) );
  AOI211_X1 U16285 ( .C1(n14571), .C2(n14716), .A(n14384), .B(n14383), .ZN(
        n14385) );
  OAI21_X1 U16286 ( .B1(n14574), .B2(n14526), .A(n14385), .ZN(P1_U3267) );
  AOI21_X1 U16287 ( .B1(n14389), .B2(n14388), .A(n14387), .ZN(n14576) );
  INV_X1 U16288 ( .A(n14390), .ZN(n14452) );
  OAI211_X1 U16289 ( .C1(n14412), .C2(n14394), .A(n6732), .B(n14712), .ZN(
        n14581) );
  INV_X1 U16290 ( .A(n14581), .ZN(n14396) );
  AOI22_X1 U16291 ( .A1(n14531), .A2(n14577), .B1(n14391), .B2(n14703), .ZN(
        n14393) );
  NAND2_X1 U16292 ( .A1(n14526), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n14392) );
  OAI211_X1 U16293 ( .C1(n14394), .C2(n14506), .A(n14393), .B(n14392), .ZN(
        n14395) );
  AOI21_X1 U16294 ( .B1(n14396), .B2(n14716), .A(n14395), .ZN(n14400) );
  NAND2_X1 U16295 ( .A1(n14398), .A2(n14397), .ZN(n14579) );
  NAND3_X1 U16296 ( .A1(n14580), .A2(n14579), .A3(n14717), .ZN(n14399) );
  OAI211_X1 U16297 ( .C1(n14576), .C2(n14452), .A(n14400), .B(n14399), .ZN(
        P1_U3268) );
  NAND2_X1 U16298 ( .A1(n14401), .A2(n14406), .ZN(n14402) );
  NAND3_X1 U16299 ( .A1(n14403), .A2(n14701), .A3(n14402), .ZN(n14410) );
  AOI22_X1 U16300 ( .A1(n14540), .A2(n14404), .B1(n14440), .B2(n14539), .ZN(
        n14409) );
  XNOR2_X1 U16301 ( .A(n14405), .B(n14406), .ZN(n14407) );
  NAND2_X1 U16302 ( .A1(n14407), .A2(n14965), .ZN(n14408) );
  NAND3_X1 U16303 ( .A1(n14410), .A2(n14409), .A3(n14408), .ZN(n14589) );
  NAND2_X1 U16304 ( .A1(n14422), .A2(n14585), .ZN(n14411) );
  NAND2_X1 U16305 ( .A1(n14411), .A2(n14712), .ZN(n14413) );
  OR2_X1 U16306 ( .A1(n14413), .A2(n14412), .ZN(n14586) );
  AOI22_X1 U16307 ( .A1(n14526), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n14414), 
        .B2(n14703), .ZN(n14416) );
  NAND2_X1 U16308 ( .A1(n14585), .A2(n14706), .ZN(n14415) );
  OAI211_X1 U16309 ( .C1(n14586), .C2(n14529), .A(n14416), .B(n14415), .ZN(
        n14417) );
  AOI21_X1 U16310 ( .B1(n14589), .B2(n14531), .A(n14417), .ZN(n14418) );
  INV_X1 U16311 ( .A(n14418), .ZN(P1_U3269) );
  XNOR2_X1 U16312 ( .A(n14419), .B(n14427), .ZN(n14421) );
  AOI21_X1 U16313 ( .B1(n14421), .B2(n14701), .A(n14420), .ZN(n14595) );
  AOI211_X1 U16314 ( .C1(n14423), .C2(n14435), .A(n14503), .B(n7104), .ZN(
        n14593) );
  AOI22_X1 U16315 ( .A1(n14526), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n14424), 
        .B2(n14703), .ZN(n14425) );
  OAI21_X1 U16316 ( .B1(n14426), .B2(n14506), .A(n14425), .ZN(n14430) );
  XNOR2_X1 U16317 ( .A(n14428), .B(n14427), .ZN(n14596) );
  NOR2_X1 U16318 ( .A1(n14596), .A2(n14511), .ZN(n14429) );
  AOI211_X1 U16319 ( .C1(n14593), .C2(n14716), .A(n14430), .B(n14429), .ZN(
        n14431) );
  OAI21_X1 U16320 ( .B1(n14595), .B2(n14526), .A(n14431), .ZN(P1_U3270) );
  INV_X1 U16321 ( .A(n14432), .ZN(n14433) );
  AOI21_X1 U16322 ( .B1(n14448), .B2(n14434), .A(n14433), .ZN(n14604) );
  AOI21_X1 U16323 ( .B1(n14456), .B2(n14599), .A(n14503), .ZN(n14436) );
  AND2_X1 U16324 ( .A1(n14436), .A2(n14435), .ZN(n14597) );
  AOI22_X1 U16325 ( .A1(n14437), .A2(n14703), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n14526), .ZN(n14444) );
  OR2_X1 U16326 ( .A1(n14439), .A2(n14438), .ZN(n14442) );
  NAND2_X1 U16327 ( .A1(n14440), .A2(n14540), .ZN(n14441) );
  NAND2_X1 U16328 ( .A1(n14442), .A2(n14441), .ZN(n14598) );
  NAND2_X1 U16329 ( .A1(n14598), .A2(n14531), .ZN(n14443) );
  OAI211_X1 U16330 ( .C1(n14445), .C2(n14506), .A(n14444), .B(n14443), .ZN(
        n14446) );
  AOI21_X1 U16331 ( .B1(n14597), .B2(n14716), .A(n14446), .ZN(n14451) );
  OAI21_X1 U16332 ( .B1(n14449), .B2(n14448), .A(n14447), .ZN(n14600) );
  NAND2_X1 U16333 ( .A1(n14600), .A2(n14717), .ZN(n14450) );
  OAI211_X1 U16334 ( .C1(n14604), .C2(n14452), .A(n14451), .B(n14450), .ZN(
        P1_U3271) );
  NAND2_X1 U16335 ( .A1(n14453), .A2(n14454), .ZN(n14455) );
  XOR2_X1 U16336 ( .A(n14462), .B(n14455), .Z(n14608) );
  INV_X1 U16337 ( .A(n14481), .ZN(n14458) );
  INV_X1 U16338 ( .A(n14456), .ZN(n14457) );
  AOI211_X1 U16339 ( .C1(n6970), .C2(n14458), .A(n14503), .B(n14457), .ZN(
        n14606) );
  INV_X1 U16340 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n14459) );
  OAI22_X1 U16341 ( .A1(n14460), .A2(n14506), .B1(n14531), .B2(n14459), .ZN(
        n14471) );
  OAI211_X1 U16342 ( .C1(n14463), .C2(n14462), .A(n14461), .B(n14701), .ZN(
        n14465) );
  NAND2_X1 U16343 ( .A1(n14496), .A2(n14539), .ZN(n14464) );
  OAI211_X1 U16344 ( .C1(n14467), .C2(n14466), .A(n14465), .B(n14464), .ZN(
        n14605) );
  AOI21_X1 U16345 ( .B1(n14468), .B2(n14703), .A(n14605), .ZN(n14469) );
  NOR2_X1 U16346 ( .A1(n14469), .A2(n14705), .ZN(n14470) );
  AOI211_X1 U16347 ( .C1(n14606), .C2(n14716), .A(n14471), .B(n14470), .ZN(
        n14472) );
  OAI21_X1 U16348 ( .B1(n14608), .B2(n14511), .A(n14472), .ZN(P1_U3272) );
  NAND2_X1 U16349 ( .A1(n14473), .A2(n14475), .ZN(n14474) );
  NAND2_X1 U16350 ( .A1(n14453), .A2(n14474), .ZN(n14612) );
  XNOR2_X1 U16351 ( .A(n14476), .B(n14475), .ZN(n14477) );
  NAND2_X1 U16352 ( .A1(n14477), .A2(n14701), .ZN(n14479) );
  NAND2_X1 U16353 ( .A1(n14479), .A2(n14478), .ZN(n14614) );
  NAND2_X1 U16354 ( .A1(n14614), .A2(n14531), .ZN(n14488) );
  AND2_X1 U16355 ( .A1(n14609), .A2(n14501), .ZN(n14480) );
  OR3_X1 U16356 ( .A1(n14481), .A2(n14480), .A3(n14503), .ZN(n14610) );
  INV_X1 U16357 ( .A(n14610), .ZN(n14486) );
  AOI22_X1 U16358 ( .A1(n14705), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n14482), 
        .B2(n14703), .ZN(n14483) );
  OAI21_X1 U16359 ( .B1(n14484), .B2(n14506), .A(n14483), .ZN(n14485) );
  AOI21_X1 U16360 ( .B1(n14486), .B2(n14716), .A(n14485), .ZN(n14487) );
  OAI211_X1 U16361 ( .C1(n14612), .C2(n14511), .A(n14488), .B(n14487), .ZN(
        P1_U3273) );
  NAND2_X1 U16362 ( .A1(n14490), .A2(n14489), .ZN(n14492) );
  NAND2_X1 U16363 ( .A1(n14492), .A2(n14495), .ZN(n14491) );
  OAI21_X1 U16364 ( .B1(n14492), .B2(n14495), .A(n14491), .ZN(n14493) );
  INV_X1 U16365 ( .A(n14493), .ZN(n14619) );
  XNOR2_X1 U16366 ( .A(n14494), .B(n14495), .ZN(n14497) );
  AOI222_X1 U16367 ( .A1(n14701), .A2(n14497), .B1(n14496), .B2(n14540), .C1(
        n14541), .C2(n14539), .ZN(n14618) );
  OAI21_X1 U16368 ( .B1(n14499), .B2(n14498), .A(n14618), .ZN(n14500) );
  NAND2_X1 U16369 ( .A1(n14500), .A2(n14531), .ZN(n14510) );
  INV_X1 U16370 ( .A(n14524), .ZN(n14504) );
  INV_X1 U16371 ( .A(n14501), .ZN(n14502) );
  AOI211_X1 U16372 ( .C1(n14616), .C2(n14504), .A(n14503), .B(n14502), .ZN(
        n14615) );
  INV_X1 U16373 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n14505) );
  OAI22_X1 U16374 ( .A1(n14507), .A2(n14506), .B1(n14505), .B2(n14531), .ZN(
        n14508) );
  AOI21_X1 U16375 ( .B1(n14615), .B2(n14716), .A(n14508), .ZN(n14509) );
  OAI211_X1 U16376 ( .C1(n14619), .C2(n14511), .A(n14510), .B(n14509), .ZN(
        P1_U3274) );
  XNOR2_X1 U16377 ( .A(n14513), .B(n14512), .ZN(n14521) );
  OAI211_X1 U16378 ( .C1(n14516), .C2(n14515), .A(n14514), .B(n14701), .ZN(
        n14520) );
  AOI22_X1 U16379 ( .A1(n14518), .A2(n14540), .B1(n14539), .B2(n14517), .ZN(
        n14519) );
  OAI211_X1 U16380 ( .C1(n14521), .C2(n14959), .A(n14520), .B(n14519), .ZN(
        n14621) );
  NAND2_X1 U16381 ( .A1(n14534), .A2(n14620), .ZN(n14522) );
  NAND2_X1 U16382 ( .A1(n14522), .A2(n14712), .ZN(n14523) );
  OR2_X1 U16383 ( .A1(n14524), .A2(n14523), .ZN(n14622) );
  AOI22_X1 U16384 ( .A1(n14526), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14525), 
        .B2(n14703), .ZN(n14528) );
  NAND2_X1 U16385 ( .A1(n14620), .A2(n14706), .ZN(n14527) );
  OAI211_X1 U16386 ( .C1(n14622), .C2(n14529), .A(n14528), .B(n14527), .ZN(
        n14530) );
  AOI21_X1 U16387 ( .B1(n14621), .B2(n14531), .A(n14530), .ZN(n14532) );
  INV_X1 U16388 ( .A(n14532), .ZN(P1_U3275) );
  OAI211_X1 U16389 ( .C1(n11883), .C2(n8853), .A(n14712), .B(n14534), .ZN(
        n14625) );
  XOR2_X1 U16390 ( .A(n14537), .B(n14535), .Z(n14545) );
  XOR2_X1 U16391 ( .A(n14536), .B(n14537), .Z(n14543) );
  AOI22_X1 U16392 ( .A1(n14541), .A2(n14540), .B1(n14539), .B2(n14538), .ZN(
        n14542) );
  OAI21_X1 U16393 ( .B1(n14543), .B2(n14603), .A(n14542), .ZN(n14544) );
  AOI21_X1 U16394 ( .B1(n14965), .B2(n14545), .A(n14544), .ZN(n14626) );
  INV_X1 U16395 ( .A(n14546), .ZN(n14549) );
  INV_X1 U16396 ( .A(n14547), .ZN(n14548) );
  AOI22_X1 U16397 ( .A1(n14550), .A2(n14549), .B1(n14548), .B2(n14703), .ZN(
        n14551) );
  OAI211_X1 U16398 ( .C1(n14552), .C2(n14625), .A(n14626), .B(n14551), .ZN(
        n14553) );
  MUX2_X1 U16399 ( .A(P1_REG2_REG_17__SCAN_IN), .B(n14553), .S(n14531), .Z(
        P1_U3276) );
  OAI211_X1 U16400 ( .C1(n14947), .C2(n14555), .A(n14554), .B(n14556), .ZN(
        n14643) );
  MUX2_X1 U16401 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14643), .S(n14982), .Z(
        P1_U3559) );
  OAI211_X1 U16402 ( .C1(n14947), .C2(n14558), .A(n14557), .B(n14556), .ZN(
        n14644) );
  MUX2_X1 U16403 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14644), .S(n14982), .Z(
        P1_U3558) );
  NAND2_X1 U16404 ( .A1(n14562), .A2(n14701), .ZN(n14563) );
  MUX2_X1 U16405 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14645), .S(n14982), .Z(
        P1_U3557) );
  MUX2_X1 U16406 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14565), .S(n14982), .Z(
        P1_U3556) );
  INV_X1 U16407 ( .A(n14567), .ZN(n14568) );
  MUX2_X1 U16408 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14646), .S(n14982), .Z(
        P1_U3555) );
  AOI21_X1 U16409 ( .B1(n14572), .B2(n14963), .A(n14571), .ZN(n14573) );
  OAI211_X1 U16410 ( .C1(n14959), .C2(n14575), .A(n14574), .B(n14573), .ZN(
        n14647) );
  MUX2_X1 U16411 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14647), .S(n14982), .Z(
        P1_U3554) );
  OR2_X1 U16412 ( .A1(n14576), .A2(n14603), .ZN(n14584) );
  AOI21_X1 U16413 ( .B1(n14578), .B2(n14963), .A(n14577), .ZN(n14583) );
  NAND3_X1 U16414 ( .A1(n14580), .A2(n14965), .A3(n14579), .ZN(n14582) );
  NAND4_X1 U16415 ( .A1(n14584), .A2(n14583), .A3(n14582), .A4(n14581), .ZN(
        n14648) );
  MUX2_X1 U16416 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14648), .S(n14982), .Z(
        P1_U3553) );
  INV_X1 U16417 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n14590) );
  INV_X1 U16418 ( .A(n14585), .ZN(n14587) );
  OAI21_X1 U16419 ( .B1(n14587), .B2(n14947), .A(n14586), .ZN(n14588) );
  NOR2_X1 U16420 ( .A1(n14589), .A2(n14588), .ZN(n14649) );
  MUX2_X1 U16421 ( .A(n14590), .B(n14649), .S(n14982), .Z(n14591) );
  INV_X1 U16422 ( .A(n14591), .ZN(P1_U3552) );
  NOR2_X1 U16423 ( .A1(n14593), .A2(n14592), .ZN(n14594) );
  OAI211_X1 U16424 ( .C1(n14959), .C2(n14596), .A(n14595), .B(n14594), .ZN(
        n14652) );
  MUX2_X1 U16425 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14652), .S(n14982), .Z(
        P1_U3551) );
  AOI211_X1 U16426 ( .C1(n14599), .C2(n14963), .A(n14598), .B(n14597), .ZN(
        n14602) );
  NAND2_X1 U16427 ( .A1(n14600), .A2(n14965), .ZN(n14601) );
  OAI211_X1 U16428 ( .C1(n14604), .C2(n14603), .A(n14602), .B(n14601), .ZN(
        n14653) );
  MUX2_X1 U16429 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14653), .S(n14982), .Z(
        P1_U3550) );
  AOI211_X1 U16430 ( .C1(n6970), .C2(n14963), .A(n14606), .B(n14605), .ZN(
        n14607) );
  OAI21_X1 U16431 ( .B1(n14608), .B2(n14959), .A(n14607), .ZN(n14654) );
  MUX2_X1 U16432 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14654), .S(n14982), .Z(
        P1_U3549) );
  NAND2_X1 U16433 ( .A1(n14609), .A2(n14963), .ZN(n14611) );
  OAI211_X1 U16434 ( .C1(n14612), .C2(n14959), .A(n14611), .B(n14610), .ZN(
        n14613) );
  MUX2_X1 U16435 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14655), .S(n14982), .Z(
        P1_U3548) );
  AOI21_X1 U16436 ( .B1(n14616), .B2(n14963), .A(n14615), .ZN(n14617) );
  OAI211_X1 U16437 ( .C1(n14619), .C2(n14959), .A(n14618), .B(n14617), .ZN(
        n14656) );
  MUX2_X1 U16438 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14656), .S(n14982), .Z(
        P1_U3547) );
  INV_X1 U16439 ( .A(n14620), .ZN(n14624) );
  INV_X1 U16440 ( .A(n14621), .ZN(n14623) );
  OAI211_X1 U16441 ( .C1(n14624), .C2(n14947), .A(n14623), .B(n14622), .ZN(
        n14657) );
  MUX2_X1 U16442 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14657), .S(n14982), .Z(
        P1_U3546) );
  OAI211_X1 U16443 ( .C1(n8853), .C2(n14947), .A(n14626), .B(n14625), .ZN(
        n14658) );
  MUX2_X1 U16444 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14658), .S(n14982), .Z(
        P1_U3545) );
  INV_X1 U16445 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n14631) );
  OAI21_X1 U16446 ( .B1(n14628), .B2(n14947), .A(n14627), .ZN(n14629) );
  NOR2_X1 U16447 ( .A1(n14630), .A2(n14629), .ZN(n14659) );
  MUX2_X1 U16448 ( .A(n14631), .B(n14659), .S(n14982), .Z(n14632) );
  INV_X1 U16449 ( .A(n14632), .ZN(P1_U3544) );
  AOI21_X1 U16450 ( .B1(n14634), .B2(n14963), .A(n14633), .ZN(n14635) );
  OAI211_X1 U16451 ( .C1(n14637), .C2(n14959), .A(n14636), .B(n14635), .ZN(
        n14662) );
  MUX2_X1 U16452 ( .A(n14662), .B(P1_REG1_REG_15__SCAN_IN), .S(n14980), .Z(
        P1_U3543) );
  AOI21_X1 U16453 ( .B1(n14639), .B2(n14963), .A(n14638), .ZN(n14640) );
  OAI211_X1 U16454 ( .C1(n14959), .C2(n14642), .A(n14641), .B(n14640), .ZN(
        n14663) );
  MUX2_X1 U16455 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n14663), .S(n14982), .Z(
        P1_U3542) );
  MUX2_X1 U16456 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14643), .S(n14973), .Z(
        P1_U3527) );
  MUX2_X1 U16457 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14644), .S(n14973), .Z(
        P1_U3526) );
  MUX2_X1 U16458 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14645), .S(n14973), .Z(
        P1_U3525) );
  MUX2_X1 U16459 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14646), .S(n14973), .Z(
        P1_U3523) );
  MUX2_X1 U16460 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14647), .S(n14973), .Z(
        P1_U3522) );
  MUX2_X1 U16461 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14648), .S(n14973), .Z(
        P1_U3521) );
  INV_X1 U16462 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n14650) );
  MUX2_X1 U16463 ( .A(n14650), .B(n14649), .S(n14973), .Z(n14651) );
  INV_X1 U16464 ( .A(n14651), .ZN(P1_U3520) );
  MUX2_X1 U16465 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14652), .S(n14973), .Z(
        P1_U3519) );
  MUX2_X1 U16466 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14653), .S(n14973), .Z(
        P1_U3518) );
  MUX2_X1 U16467 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14654), .S(n14973), .Z(
        P1_U3517) );
  MUX2_X1 U16468 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14655), .S(n14973), .Z(
        P1_U3516) );
  MUX2_X1 U16469 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14656), .S(n14973), .Z(
        P1_U3515) );
  MUX2_X1 U16470 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14657), .S(n14973), .Z(
        P1_U3513) );
  MUX2_X1 U16471 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14658), .S(n14973), .Z(
        P1_U3510) );
  INV_X1 U16472 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n14660) );
  MUX2_X1 U16473 ( .A(n14660), .B(n14659), .S(n14973), .Z(n14661) );
  INV_X1 U16474 ( .A(n14661), .ZN(P1_U3507) );
  MUX2_X1 U16475 ( .A(n14662), .B(P1_REG0_REG_15__SCAN_IN), .S(n14971), .Z(
        P1_U3504) );
  MUX2_X1 U16476 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n14663), .S(n14973), .Z(
        P1_U3501) );
  NOR4_X1 U16477 ( .A1(n7512), .A2(P1_IR_REG_30__SCAN_IN), .A3(n8290), .A4(
        P1_U3086), .ZN(n14665) );
  AOI21_X1 U16478 ( .B1(n14666), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n14665), 
        .ZN(n14667) );
  OAI21_X1 U16479 ( .B1(n14669), .B2(n14668), .A(n14667), .ZN(P1_U3324) );
  OAI222_X1 U16480 ( .A1(n14668), .A2(n14672), .B1(P1_U3086), .B2(n14671), 
        .C1(n14670), .C2(n12137), .ZN(P1_U3326) );
  MUX2_X1 U16481 ( .A(n14673), .B(n8899), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  MUX2_X1 U16482 ( .A(n14674), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  OAI21_X1 U16483 ( .B1(n14677), .B2(n14676), .A(n14675), .ZN(n14678) );
  XNOR2_X1 U16484 ( .A(n14678), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16485 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14679) );
  OAI21_X1 U16486 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14679), 
        .ZN(U28) );
  AOI21_X1 U16487 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14680) );
  OAI21_X1 U16488 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14680), 
        .ZN(U29) );
  OAI21_X1 U16489 ( .B1(n14683), .B2(n14682), .A(n14681), .ZN(n14684) );
  XNOR2_X1 U16490 ( .A(n14684), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  AOI21_X1 U16491 ( .B1(n14687), .B2(n14686), .A(n14685), .ZN(SUB_1596_U57) );
  AOI21_X1 U16492 ( .B1(n14690), .B2(n14689), .A(n14688), .ZN(SUB_1596_U55) );
  AOI21_X1 U16493 ( .B1(n14692), .B2(n14691), .A(n6813), .ZN(n14693) );
  XOR2_X1 U16494 ( .A(n14693), .B(P2_ADDR_REG_9__SCAN_IN), .Z(SUB_1596_U54) );
  AOI21_X1 U16495 ( .B1(n14696), .B2(n14695), .A(n14694), .ZN(n14697) );
  XOR2_X1 U16496 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n14697), .Z(SUB_1596_U70)
         );
  XOR2_X1 U16497 ( .A(n14709), .B(n14698), .Z(n14702) );
  INV_X1 U16498 ( .A(n14699), .ZN(n14700) );
  AOI21_X1 U16499 ( .B1(n14702), .B2(n14701), .A(n14700), .ZN(n14722) );
  AOI222_X1 U16500 ( .A1(n14707), .A2(n14706), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n14705), .C1(n14704), .C2(n14703), .ZN(n14719) );
  XNOR2_X1 U16501 ( .A(n14708), .B(n14709), .ZN(n14725) );
  INV_X1 U16502 ( .A(n14710), .ZN(n14714) );
  INV_X1 U16503 ( .A(n14711), .ZN(n14713) );
  OAI211_X1 U16504 ( .C1(n14721), .C2(n14714), .A(n14713), .B(n14712), .ZN(
        n14720) );
  INV_X1 U16505 ( .A(n14720), .ZN(n14715) );
  AOI22_X1 U16506 ( .A1(n14725), .A2(n14717), .B1(n14716), .B2(n14715), .ZN(
        n14718) );
  OAI211_X1 U16507 ( .C1(n14526), .C2(n14722), .A(n14719), .B(n14718), .ZN(
        P1_U3281) );
  OAI21_X1 U16508 ( .B1(n14721), .B2(n14947), .A(n14720), .ZN(n14724) );
  INV_X1 U16509 ( .A(n14722), .ZN(n14723) );
  AOI211_X1 U16510 ( .C1(n14965), .C2(n14725), .A(n14724), .B(n14723), .ZN(
        n14728) );
  INV_X1 U16511 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14726) );
  AOI22_X1 U16512 ( .A1(n14973), .A2(n14728), .B1(n14726), .B2(n14971), .ZN(
        P1_U3495) );
  AOI22_X1 U16513 ( .A1(n14982), .A2(n14728), .B1(n14727), .B2(n14980), .ZN(
        P1_U3540) );
  OAI21_X1 U16514 ( .B1(n14731), .B2(n14730), .A(n14729), .ZN(SUB_1596_U63) );
  INV_X1 U16515 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14732) );
  OAI22_X1 U16516 ( .A1(n15320), .A2(n14733), .B1(n15308), .B2(n14732), .ZN(
        n14734) );
  INV_X1 U16517 ( .A(n14734), .ZN(n14752) );
  MUX2_X1 U16518 ( .A(n14737), .B(n14736), .S(n14735), .Z(n14738) );
  NAND2_X1 U16519 ( .A1(n14739), .A2(n14738), .ZN(n14741) );
  XOR2_X1 U16520 ( .A(n14741), .B(n14740), .Z(n14745) );
  XNOR2_X1 U16521 ( .A(n14743), .B(n14742), .ZN(n14744) );
  AOI22_X1 U16522 ( .A1(n14745), .A2(n15305), .B1(n15329), .B2(n14744), .ZN(
        n14751) );
  NAND2_X1 U16523 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(P3_U3151), .ZN(n14750)
         );
  OAI221_X1 U16524 ( .B1(n14748), .B2(n14747), .C1(n14748), .C2(n14746), .A(
        n15264), .ZN(n14749) );
  NAND4_X1 U16525 ( .A1(n14752), .A2(n14751), .A3(n14750), .A4(n14749), .ZN(
        P3_U3198) );
  AOI22_X1 U16526 ( .A1(n15266), .A2(n14753), .B1(n15326), .B2(
        P3_ADDR_REG_17__SCAN_IN), .ZN(n14767) );
  OAI21_X1 U16527 ( .B1(P3_REG1_REG_17__SCAN_IN), .B2(n14755), .A(n14754), 
        .ZN(n14760) );
  AOI211_X1 U16528 ( .C1(n14758), .C2(n14757), .A(n15322), .B(n14756), .ZN(
        n14759) );
  AOI21_X1 U16529 ( .B1(n15329), .B2(n14760), .A(n14759), .ZN(n14766) );
  OAI221_X1 U16530 ( .B1(n14763), .B2(n14762), .C1(n14763), .C2(n14761), .A(
        n15264), .ZN(n14764) );
  NAND4_X1 U16531 ( .A1(n14767), .A2(n14766), .A3(n14765), .A4(n14764), .ZN(
        P3_U3199) );
  INV_X1 U16532 ( .A(n14768), .ZN(n14769) );
  AOI21_X1 U16533 ( .B1(n14771), .B2(n14770), .A(n14769), .ZN(n14781) );
  INV_X1 U16534 ( .A(n14781), .ZN(n14772) );
  OAI22_X1 U16535 ( .A1(n15433), .A2(n14772), .B1(P3_REG1_REG_30__SCAN_IN), 
        .B2(n15436), .ZN(n14773) );
  INV_X1 U16536 ( .A(n14773), .ZN(P3_U3489) );
  AOI21_X1 U16537 ( .B1(n14776), .B2(n14775), .A(n14774), .ZN(n14777) );
  AND2_X1 U16538 ( .A1(n14778), .A2(n14777), .ZN(n14783) );
  INV_X1 U16539 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14779) );
  AOI22_X1 U16540 ( .A1(n15436), .A2(n14783), .B1(n14779), .B2(n15433), .ZN(
        P3_U3470) );
  INV_X1 U16541 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n14780) );
  AOI22_X1 U16542 ( .A1(n15421), .A2(n14781), .B1(n14780), .B2(n15419), .ZN(
        P3_U3457) );
  INV_X1 U16543 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14782) );
  AOI22_X1 U16544 ( .A1(n15421), .A2(n14783), .B1(n14782), .B2(n15419), .ZN(
        P3_U3423) );
  OR2_X1 U16545 ( .A1(n14785), .A2(n14784), .ZN(n14789) );
  NAND2_X1 U16546 ( .A1(n14787), .A2(n14786), .ZN(n14788) );
  NAND2_X1 U16547 ( .A1(n14789), .A2(n14788), .ZN(n14802) );
  OAI21_X1 U16548 ( .B1(n14792), .B2(n14791), .A(n14790), .ZN(n14794) );
  AOI222_X1 U16549 ( .A1(n14796), .A2(n7081), .B1(n14802), .B2(n14795), .C1(
        n14794), .C2(n14793), .ZN(n14798) );
  OAI211_X1 U16550 ( .C1(n14799), .C2(n14804), .A(n14798), .B(n14797), .ZN(
        P2_U3187) );
  XNOR2_X1 U16551 ( .A(n14801), .B(n14800), .ZN(n14803) );
  AOI21_X1 U16552 ( .B1(n14803), .B2(n15054), .A(n14802), .ZN(n14817) );
  INV_X1 U16553 ( .A(n14804), .ZN(n14805) );
  AOI222_X1 U16554 ( .A1(n7081), .A2(n15060), .B1(P2_REG2_REG_14__SCAN_IN), 
        .B2(n15059), .C1(n15058), .C2(n14805), .ZN(n14814) );
  OAI21_X1 U16555 ( .B1(n14808), .B2(n14807), .A(n14806), .ZN(n14820) );
  INV_X1 U16556 ( .A(n14809), .ZN(n14810) );
  OAI211_X1 U16557 ( .C1(n14816), .C2(n14811), .A(n14810), .B(n15065), .ZN(
        n14815) );
  INV_X1 U16558 ( .A(n14815), .ZN(n14812) );
  AOI22_X1 U16559 ( .A1(n14820), .A2(n15069), .B1(n15068), .B2(n14812), .ZN(
        n14813) );
  OAI211_X1 U16560 ( .C1(n15059), .C2(n14817), .A(n14814), .B(n14813), .ZN(
        P2_U3251) );
  OAI21_X1 U16561 ( .B1(n14816), .B2(n15150), .A(n14815), .ZN(n14819) );
  INV_X1 U16562 ( .A(n14817), .ZN(n14818) );
  AOI211_X1 U16563 ( .C1(n15147), .C2(n14820), .A(n14819), .B(n14818), .ZN(
        n14838) );
  AOI22_X1 U16564 ( .A1(n15177), .A2(n14838), .B1(n14821), .B2(n15174), .ZN(
        P2_U3513) );
  NOR3_X1 U16565 ( .A1(n14823), .A2(n14822), .A3(n15117), .ZN(n14827) );
  NOR2_X1 U16566 ( .A1(n14824), .A2(n15150), .ZN(n14825) );
  NOR4_X1 U16567 ( .A1(n14828), .A2(n14827), .A3(n14826), .A4(n14825), .ZN(
        n14840) );
  AOI22_X1 U16568 ( .A1(n15177), .A2(n14840), .B1(n14829), .B2(n15174), .ZN(
        P2_U3512) );
  INV_X1 U16569 ( .A(n14830), .ZN(n14832) );
  OAI21_X1 U16570 ( .B1(n14832), .B2(n15150), .A(n14831), .ZN(n14834) );
  AOI211_X1 U16571 ( .C1(n14835), .C2(n15147), .A(n14834), .B(n14833), .ZN(
        n14842) );
  AOI22_X1 U16572 ( .A1(n15177), .A2(n14842), .B1(n14836), .B2(n15174), .ZN(
        P2_U3511) );
  INV_X1 U16573 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n14837) );
  AOI22_X1 U16574 ( .A1(n15157), .A2(n14838), .B1(n14837), .B2(n15156), .ZN(
        P2_U3472) );
  INV_X1 U16575 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n14839) );
  AOI22_X1 U16576 ( .A1(n15157), .A2(n14840), .B1(n14839), .B2(n15156), .ZN(
        P2_U3469) );
  INV_X1 U16577 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14841) );
  AOI22_X1 U16578 ( .A1(n15157), .A2(n14842), .B1(n14841), .B2(n15156), .ZN(
        P2_U3466) );
  NAND2_X1 U16579 ( .A1(n14843), .A2(n14963), .ZN(n14865) );
  INV_X1 U16580 ( .A(n14844), .ZN(n14846) );
  OAI22_X1 U16581 ( .A1(n14865), .A2(n14846), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14845), .ZN(n14847) );
  INV_X1 U16582 ( .A(n14847), .ZN(n14857) );
  NAND2_X1 U16583 ( .A1(n14848), .A2(n14849), .ZN(n14851) );
  AOI21_X1 U16584 ( .B1(n14852), .B2(n14851), .A(n14850), .ZN(n14853) );
  AOI21_X1 U16585 ( .B1(n14855), .B2(n14854), .A(n14853), .ZN(n14856) );
  OAI211_X1 U16586 ( .C1(n14858), .C2(n14909), .A(n14857), .B(n14856), .ZN(
        P1_U3236) );
  OAI21_X1 U16587 ( .B1(n14860), .B2(n14947), .A(n14859), .ZN(n14863) );
  INV_X1 U16588 ( .A(n14861), .ZN(n14862) );
  AOI211_X1 U16589 ( .C1(n14965), .C2(n14864), .A(n14863), .B(n14862), .ZN(
        n14869) );
  AOI22_X1 U16590 ( .A1(n14982), .A2(n14869), .B1(n11025), .B2(n14980), .ZN(
        P1_U3541) );
  AOI22_X1 U16591 ( .A1(n14982), .A2(n14871), .B1(n10554), .B2(n14980), .ZN(
        P1_U3539) );
  INV_X1 U16592 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14868) );
  AOI22_X1 U16593 ( .A1(n14973), .A2(n14869), .B1(n14868), .B2(n14971), .ZN(
        P1_U3498) );
  INV_X1 U16594 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14870) );
  AOI22_X1 U16595 ( .A1(n14973), .A2(n14871), .B1(n14870), .B2(n14971), .ZN(
        P1_U3492) );
  OAI21_X1 U16596 ( .B1(n14874), .B2(n14873), .A(n14872), .ZN(n14875) );
  XNOR2_X1 U16597 ( .A(n14875), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  OAI21_X1 U16598 ( .B1(n14877), .B2(n15036), .A(n14876), .ZN(SUB_1596_U68) );
  OAI21_X1 U16599 ( .B1(n14880), .B2(n14879), .A(n14878), .ZN(SUB_1596_U67) );
  OAI21_X1 U16600 ( .B1(n14883), .B2(n14882), .A(n14881), .ZN(n14884) );
  XNOR2_X1 U16601 ( .A(n14884), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  OAI21_X1 U16602 ( .B1(n14887), .B2(n14886), .A(n14885), .ZN(n14888) );
  XNOR2_X1 U16603 ( .A(n14888), .B(P2_ADDR_REG_15__SCAN_IN), .ZN(SUB_1596_U65)
         );
  INV_X1 U16604 ( .A(n14891), .ZN(n14890) );
  OAI222_X1 U16605 ( .A1(n14893), .A2(n14892), .B1(n14893), .B2(n14891), .C1(
        n14890), .C2(n14889), .ZN(SUB_1596_U64) );
  XNOR2_X1 U16606 ( .A(n14895), .B(n14894), .ZN(n14905) );
  NOR2_X1 U16607 ( .A1(n14897), .A2(n14896), .ZN(n14903) );
  OAI22_X1 U16608 ( .A1(n14901), .A2(n14900), .B1(n14899), .B2(n14898), .ZN(
        n14902) );
  AOI211_X1 U16609 ( .C1(n14905), .C2(n14904), .A(n14903), .B(n14902), .ZN(
        n14907) );
  OAI211_X1 U16610 ( .C1(n14909), .C2(n14908), .A(n14907), .B(n14906), .ZN(
        P1_U3231) );
  OAI21_X1 U16611 ( .B1(n14912), .B2(n14911), .A(n14910), .ZN(n14914) );
  NAND2_X1 U16612 ( .A1(n14914), .A2(n14913), .ZN(n14920) );
  AOI21_X1 U16613 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14916), .A(n14915), 
        .ZN(n14918) );
  OR2_X1 U16614 ( .A1(n14918), .A2(n14917), .ZN(n14919) );
  OAI211_X1 U16615 ( .C1(n14922), .C2(n14921), .A(n14920), .B(n14919), .ZN(
        n14923) );
  INV_X1 U16616 ( .A(n14923), .ZN(n14925) );
  OAI211_X1 U16617 ( .C1(n14927), .C2(n14926), .A(n14925), .B(n14924), .ZN(
        P1_U3258) );
  AND2_X1 U16618 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14930), .ZN(P1_U3294) );
  AND2_X1 U16619 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14930), .ZN(P1_U3295) );
  AND2_X1 U16620 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14930), .ZN(P1_U3296) );
  AND2_X1 U16621 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14930), .ZN(P1_U3297) );
  AND2_X1 U16622 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14930), .ZN(P1_U3298) );
  AND2_X1 U16623 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14930), .ZN(P1_U3299) );
  AND2_X1 U16624 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14930), .ZN(P1_U3300) );
  AND2_X1 U16625 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14930), .ZN(P1_U3301) );
  AND2_X1 U16626 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14930), .ZN(P1_U3302) );
  AND2_X1 U16627 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14930), .ZN(P1_U3303) );
  AND2_X1 U16628 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14930), .ZN(P1_U3304) );
  AND2_X1 U16629 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14930), .ZN(P1_U3305) );
  AND2_X1 U16630 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14930), .ZN(P1_U3306) );
  AND2_X1 U16631 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14930), .ZN(P1_U3307) );
  AND2_X1 U16632 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14930), .ZN(P1_U3308) );
  AND2_X1 U16633 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14930), .ZN(P1_U3309) );
  NOR2_X1 U16634 ( .A1(n14929), .A2(n14928), .ZN(P1_U3310) );
  AND2_X1 U16635 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14930), .ZN(P1_U3311) );
  AND2_X1 U16636 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14930), .ZN(P1_U3312) );
  AND2_X1 U16637 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14930), .ZN(P1_U3313) );
  AND2_X1 U16638 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14930), .ZN(P1_U3314) );
  AND2_X1 U16639 ( .A1(n14930), .A2(P1_D_REG_10__SCAN_IN), .ZN(P1_U3315) );
  AND2_X1 U16640 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14930), .ZN(P1_U3316) );
  AND2_X1 U16641 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14930), .ZN(P1_U3317) );
  AND2_X1 U16642 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14930), .ZN(P1_U3318) );
  AND2_X1 U16643 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14930), .ZN(P1_U3319) );
  AND2_X1 U16644 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14930), .ZN(P1_U3320) );
  AND2_X1 U16645 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14930), .ZN(P1_U3321) );
  AND2_X1 U16646 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14930), .ZN(P1_U3322) );
  AND2_X1 U16647 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14930), .ZN(P1_U3323) );
  OAI21_X1 U16648 ( .B1(n6821), .B2(n14947), .A(n14931), .ZN(n14933) );
  AOI211_X1 U16649 ( .C1(n14965), .C2(n14934), .A(n14933), .B(n14932), .ZN(
        n14975) );
  AOI22_X1 U16650 ( .A1(n14973), .A2(n14975), .B1(n14935), .B2(n14971), .ZN(
        P1_U3462) );
  INV_X1 U16651 ( .A(n14936), .ZN(n14943) );
  INV_X1 U16652 ( .A(n14937), .ZN(n14941) );
  AOI21_X1 U16653 ( .B1(n14939), .B2(n14963), .A(n14938), .ZN(n14940) );
  OAI21_X1 U16654 ( .B1(n14941), .B2(n14959), .A(n14940), .ZN(n14942) );
  NOR2_X1 U16655 ( .A1(n14943), .A2(n14942), .ZN(n14976) );
  INV_X1 U16656 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n14944) );
  AOI22_X1 U16657 ( .A1(n14973), .A2(n14976), .B1(n14944), .B2(n14971), .ZN(
        P1_U3468) );
  OAI211_X1 U16658 ( .C1(n14948), .C2(n14947), .A(n14946), .B(n14945), .ZN(
        n14949) );
  INV_X1 U16659 ( .A(n14949), .ZN(n14977) );
  INV_X1 U16660 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n14950) );
  AOI22_X1 U16661 ( .A1(n14973), .A2(n14977), .B1(n14950), .B2(n14971), .ZN(
        P1_U3474) );
  INV_X1 U16662 ( .A(n14951), .ZN(n14953) );
  AOI211_X1 U16663 ( .C1(n14954), .C2(n14963), .A(n14953), .B(n14952), .ZN(
        n14978) );
  AOI22_X1 U16664 ( .A1(n14973), .A2(n14978), .B1(n8483), .B2(n14971), .ZN(
        P1_U3480) );
  AOI21_X1 U16665 ( .B1(n14956), .B2(n14963), .A(n14955), .ZN(n14957) );
  OAI211_X1 U16666 ( .C1(n14960), .C2(n14959), .A(n14958), .B(n14957), .ZN(
        n14961) );
  INV_X1 U16667 ( .A(n14961), .ZN(n14979) );
  INV_X1 U16668 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14962) );
  AOI22_X1 U16669 ( .A1(n14973), .A2(n14979), .B1(n14962), .B2(n14971), .ZN(
        P1_U3483) );
  AOI22_X1 U16670 ( .A1(n14966), .A2(n14965), .B1(n14964), .B2(n14963), .ZN(
        n14967) );
  NAND2_X1 U16671 ( .A1(n14968), .A2(n14967), .ZN(n14969) );
  NOR2_X1 U16672 ( .A1(n14970), .A2(n14969), .ZN(n14981) );
  INV_X1 U16673 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14972) );
  AOI22_X1 U16674 ( .A1(n14973), .A2(n14981), .B1(n14972), .B2(n14971), .ZN(
        P1_U3489) );
  AOI22_X1 U16675 ( .A1(n14982), .A2(n14975), .B1(n14974), .B2(n14980), .ZN(
        P1_U3529) );
  AOI22_X1 U16676 ( .A1(n14982), .A2(n14976), .B1(n9443), .B2(n14980), .ZN(
        P1_U3531) );
  AOI22_X1 U16677 ( .A1(n14982), .A2(n14977), .B1(n9833), .B2(n14980), .ZN(
        P1_U3533) );
  AOI22_X1 U16678 ( .A1(n14982), .A2(n14978), .B1(n9855), .B2(n14980), .ZN(
        P1_U3535) );
  AOI22_X1 U16679 ( .A1(n14982), .A2(n14979), .B1(n9889), .B2(n14980), .ZN(
        P1_U3536) );
  AOI22_X1 U16680 ( .A1(n14982), .A2(n14981), .B1(n10286), .B2(n14980), .ZN(
        P1_U3538) );
  NOR2_X1 U16681 ( .A1(n15043), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI21_X1 U16682 ( .B1(n14984), .B2(P2_REG1_REG_0__SCAN_IN), .A(n14983), .ZN(
        n14989) );
  AOI22_X1 U16683 ( .A1(n15043), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n14988) );
  OAI22_X1 U16684 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n15026), .B1(n15037), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n14986) );
  OAI21_X1 U16685 ( .B1(n15032), .B2(n14986), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n14987) );
  OAI211_X1 U16686 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n14989), .A(n14988), .B(
        n14987), .ZN(P2_U3214) );
  OAI21_X1 U16687 ( .B1(n14992), .B2(n14991), .A(n14990), .ZN(n14996) );
  OR2_X1 U16688 ( .A1(n15051), .A2(n14993), .ZN(n14995) );
  OR2_X1 U16689 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9942), .ZN(n14994) );
  OAI211_X1 U16690 ( .C1(n15037), .C2(n14996), .A(n14995), .B(n14994), .ZN(
        n14997) );
  INV_X1 U16691 ( .A(n14997), .ZN(n15002) );
  OAI211_X1 U16692 ( .C1(n15000), .C2(n14999), .A(n15045), .B(n14998), .ZN(
        n15001) );
  OAI211_X1 U16693 ( .C1(n15035), .C2(n6913), .A(n15002), .B(n15001), .ZN(
        P2_U3217) );
  INV_X1 U16694 ( .A(n15003), .ZN(n15007) );
  NOR2_X1 U16695 ( .A1(n15005), .A2(n15004), .ZN(n15006) );
  OR3_X1 U16696 ( .A1(n15037), .A2(n15007), .A3(n15006), .ZN(n15008) );
  OAI211_X1 U16697 ( .C1(n15051), .C2(n15010), .A(n15009), .B(n15008), .ZN(
        n15011) );
  INV_X1 U16698 ( .A(n15011), .ZN(n15016) );
  OAI211_X1 U16699 ( .C1(n15014), .C2(n15013), .A(n15045), .B(n15012), .ZN(
        n15015) );
  OAI211_X1 U16700 ( .C1(n15035), .C2(n15017), .A(n15016), .B(n15015), .ZN(
        P2_U3221) );
  NAND2_X1 U16701 ( .A1(n15019), .A2(n15018), .ZN(n15020) );
  AOI21_X1 U16702 ( .B1(n15021), .B2(n15020), .A(n15037), .ZN(n15030) );
  INV_X1 U16703 ( .A(n15022), .ZN(n15028) );
  NAND3_X1 U16704 ( .A1(n15025), .A2(n15024), .A3(n15023), .ZN(n15027) );
  AOI21_X1 U16705 ( .B1(n15028), .B2(n15027), .A(n15026), .ZN(n15029) );
  AOI211_X1 U16706 ( .C1(n15032), .C2(n15031), .A(n15030), .B(n15029), .ZN(
        n15034) );
  OAI211_X1 U16707 ( .C1(n15036), .C2(n15035), .A(n15034), .B(n15033), .ZN(
        P2_U3226) );
  AOI211_X1 U16708 ( .C1(n15040), .C2(n15039), .A(n15038), .B(n15037), .ZN(
        n15041) );
  AOI211_X1 U16709 ( .C1(P2_ADDR_REG_16__SCAN_IN), .C2(n15043), .A(n15042), 
        .B(n15041), .ZN(n15049) );
  OAI211_X1 U16710 ( .C1(n15047), .C2(n15046), .A(n15045), .B(n15044), .ZN(
        n15048) );
  OAI211_X1 U16711 ( .C1(n15051), .C2(n15050), .A(n15049), .B(n15048), .ZN(
        P2_U3230) );
  XNOR2_X1 U16712 ( .A(n15052), .B(n15062), .ZN(n15055) );
  AOI21_X1 U16713 ( .B1(n15055), .B2(n15054), .A(n15053), .ZN(n15143) );
  INV_X1 U16714 ( .A(n15056), .ZN(n15057) );
  AOI222_X1 U16715 ( .A1(n15061), .A2(n15060), .B1(P2_REG2_REG_10__SCAN_IN), 
        .B2(n15059), .C1(n15058), .C2(n15057), .ZN(n15071) );
  XOR2_X1 U16716 ( .A(n15063), .B(n15062), .Z(n15146) );
  OAI211_X1 U16717 ( .C1(n15142), .C2(n15066), .A(n15065), .B(n15064), .ZN(
        n15141) );
  INV_X1 U16718 ( .A(n15141), .ZN(n15067) );
  AOI22_X1 U16719 ( .A1(n15146), .A2(n15069), .B1(n15068), .B2(n15067), .ZN(
        n15070) );
  OAI211_X1 U16720 ( .C1(n15072), .C2(n15143), .A(n15071), .B(n15070), .ZN(
        P2_U3255) );
  NOR2_X1 U16721 ( .A1(n15085), .A2(n15073), .ZN(n15078) );
  AND2_X1 U16722 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15079), .ZN(P2_U3266) );
  NOR2_X1 U16723 ( .A1(n15078), .A2(n15074), .ZN(P2_U3267) );
  AND2_X1 U16724 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15079), .ZN(P2_U3268) );
  AND2_X1 U16725 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15079), .ZN(P2_U3269) );
  AND2_X1 U16726 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15079), .ZN(P2_U3270) );
  AND2_X1 U16727 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15079), .ZN(P2_U3271) );
  AND2_X1 U16728 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15079), .ZN(P2_U3272) );
  AND2_X1 U16729 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15079), .ZN(P2_U3273) );
  AND2_X1 U16730 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15079), .ZN(P2_U3274) );
  AND2_X1 U16731 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15079), .ZN(P2_U3275) );
  AND2_X1 U16732 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15079), .ZN(P2_U3276) );
  AND2_X1 U16733 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15079), .ZN(P2_U3277) );
  NOR2_X1 U16734 ( .A1(n15078), .A2(n15075), .ZN(P2_U3278) );
  AND2_X1 U16735 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15079), .ZN(P2_U3279) );
  AND2_X1 U16736 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15079), .ZN(P2_U3280) );
  AND2_X1 U16737 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15079), .ZN(P2_U3281) );
  NOR2_X1 U16738 ( .A1(n15078), .A2(n15076), .ZN(P2_U3282) );
  AND2_X1 U16739 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15079), .ZN(P2_U3283) );
  AND2_X1 U16740 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15079), .ZN(P2_U3284) );
  AND2_X1 U16741 ( .A1(n15079), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3285) );
  AND2_X1 U16742 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15079), .ZN(P2_U3286) );
  AND2_X1 U16743 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15079), .ZN(P2_U3287) );
  AND2_X1 U16744 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15079), .ZN(P2_U3288) );
  NOR2_X1 U16745 ( .A1(n15078), .A2(n15077), .ZN(P2_U3289) );
  AND2_X1 U16746 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15079), .ZN(P2_U3290) );
  AND2_X1 U16747 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15079), .ZN(P2_U3291) );
  AND2_X1 U16748 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15079), .ZN(P2_U3292) );
  AND2_X1 U16749 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15079), .ZN(P2_U3293) );
  AND2_X1 U16750 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15079), .ZN(P2_U3294) );
  AND2_X1 U16751 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15079), .ZN(P2_U3295) );
  AOI22_X1 U16752 ( .A1(n15082), .A2(n15081), .B1(n15080), .B2(n15085), .ZN(
        P2_U3416) );
  AOI21_X1 U16753 ( .B1(n15085), .B2(n15084), .A(n15083), .ZN(P2_U3417) );
  INV_X1 U16754 ( .A(n15086), .ZN(n15090) );
  INV_X1 U16755 ( .A(n15087), .ZN(n15089) );
  AOI211_X1 U16756 ( .C1(n12969), .C2(n15090), .A(n15089), .B(n15088), .ZN(
        n15158) );
  INV_X1 U16757 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n15091) );
  AOI22_X1 U16758 ( .A1(n15157), .A2(n15158), .B1(n15091), .B2(n15156), .ZN(
        P2_U3430) );
  OAI21_X1 U16759 ( .B1(n15093), .B2(n15150), .A(n15092), .ZN(n15095) );
  AOI211_X1 U16760 ( .C1(n15147), .C2(n15096), .A(n15095), .B(n15094), .ZN(
        n15160) );
  INV_X1 U16761 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n15097) );
  AOI22_X1 U16762 ( .A1(n15157), .A2(n15160), .B1(n15097), .B2(n15156), .ZN(
        P2_U3436) );
  INV_X1 U16763 ( .A(n15098), .ZN(n15103) );
  OAI21_X1 U16764 ( .B1(n15100), .B2(n15150), .A(n15099), .ZN(n15102) );
  AOI211_X1 U16765 ( .C1(n12969), .C2(n15103), .A(n15102), .B(n15101), .ZN(
        n15162) );
  INV_X1 U16766 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n15104) );
  AOI22_X1 U16767 ( .A1(n15157), .A2(n15162), .B1(n15104), .B2(n15156), .ZN(
        P2_U3439) );
  AOI21_X1 U16768 ( .B1(n15114), .B2(n15106), .A(n15105), .ZN(n15110) );
  NAND3_X1 U16769 ( .A1(n15108), .A2(n15107), .A3(n15147), .ZN(n15109) );
  AND3_X1 U16770 ( .A1(n15111), .A2(n15110), .A3(n15109), .ZN(n15164) );
  AOI22_X1 U16771 ( .A1(n15157), .A2(n15164), .B1(n9944), .B2(n15156), .ZN(
        P2_U3442) );
  AOI21_X1 U16772 ( .B1(n15114), .B2(n15113), .A(n15112), .ZN(n15115) );
  OAI211_X1 U16773 ( .C1(n15118), .C2(n15117), .A(n15116), .B(n15115), .ZN(
        n15119) );
  INV_X1 U16774 ( .A(n15119), .ZN(n15166) );
  INV_X1 U16775 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n15120) );
  AOI22_X1 U16776 ( .A1(n15157), .A2(n15166), .B1(n15120), .B2(n15156), .ZN(
        P2_U3445) );
  OAI21_X1 U16777 ( .B1(n15122), .B2(n15150), .A(n15121), .ZN(n15123) );
  AOI21_X1 U16778 ( .B1(n15124), .B2(n12969), .A(n15123), .ZN(n15127) );
  NAND2_X1 U16779 ( .A1(n15124), .A2(n15155), .ZN(n15125) );
  AND3_X1 U16780 ( .A1(n15127), .A2(n15126), .A3(n15125), .ZN(n15168) );
  INV_X1 U16781 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n15128) );
  AOI22_X1 U16782 ( .A1(n15157), .A2(n15168), .B1(n15128), .B2(n15156), .ZN(
        P2_U3448) );
  OAI211_X1 U16783 ( .C1(n15131), .C2(n15150), .A(n15130), .B(n15129), .ZN(
        n15132) );
  AOI21_X1 U16784 ( .B1(n15147), .B2(n15133), .A(n15132), .ZN(n15169) );
  INV_X1 U16785 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n15134) );
  AOI22_X1 U16786 ( .A1(n15157), .A2(n15169), .B1(n15134), .B2(n15156), .ZN(
        P2_U3451) );
  INV_X1 U16787 ( .A(n15135), .ZN(n15140) );
  OAI21_X1 U16788 ( .B1(n15137), .B2(n15150), .A(n15136), .ZN(n15139) );
  AOI211_X1 U16789 ( .C1(n12969), .C2(n15140), .A(n15139), .B(n15138), .ZN(
        n15171) );
  AOI22_X1 U16790 ( .A1(n15157), .A2(n15171), .B1(n10578), .B2(n15156), .ZN(
        P2_U3454) );
  OAI21_X1 U16791 ( .B1(n15142), .B2(n15150), .A(n15141), .ZN(n15145) );
  INV_X1 U16792 ( .A(n15143), .ZN(n15144) );
  AOI211_X1 U16793 ( .C1(n15147), .C2(n15146), .A(n15145), .B(n15144), .ZN(
        n15173) );
  AOI22_X1 U16794 ( .A1(n15157), .A2(n15173), .B1(n10883), .B2(n15156), .ZN(
        P2_U3460) );
  NAND2_X1 U16795 ( .A1(n15154), .A2(n12969), .ZN(n15149) );
  OAI211_X1 U16796 ( .C1(n15151), .C2(n15150), .A(n15149), .B(n15148), .ZN(
        n15153) );
  AOI211_X1 U16797 ( .C1(n15155), .C2(n15154), .A(n15153), .B(n15152), .ZN(
        n15176) );
  AOI22_X1 U16798 ( .A1(n15157), .A2(n15176), .B1(n10991), .B2(n15156), .ZN(
        P2_U3463) );
  AOI22_X1 U16799 ( .A1(n15177), .A2(n15158), .B1(n9543), .B2(n15174), .ZN(
        P2_U3499) );
  AOI22_X1 U16800 ( .A1(n15177), .A2(n15160), .B1(n15159), .B2(n15174), .ZN(
        P2_U3501) );
  AOI22_X1 U16801 ( .A1(n15177), .A2(n15162), .B1(n15161), .B2(n15174), .ZN(
        P2_U3502) );
  AOI22_X1 U16802 ( .A1(n15177), .A2(n15164), .B1(n15163), .B2(n15174), .ZN(
        P2_U3503) );
  AOI22_X1 U16803 ( .A1(n15177), .A2(n15166), .B1(n15165), .B2(n15174), .ZN(
        P2_U3504) );
  AOI22_X1 U16804 ( .A1(n15177), .A2(n15168), .B1(n15167), .B2(n15174), .ZN(
        P2_U3505) );
  AOI22_X1 U16805 ( .A1(n15177), .A2(n15169), .B1(n10412), .B2(n15174), .ZN(
        P2_U3506) );
  AOI22_X1 U16806 ( .A1(n15177), .A2(n15171), .B1(n15170), .B2(n15174), .ZN(
        P2_U3507) );
  AOI22_X1 U16807 ( .A1(n15177), .A2(n15173), .B1(n15172), .B2(n15174), .ZN(
        P2_U3509) );
  AOI22_X1 U16808 ( .A1(n15177), .A2(n15176), .B1(n15175), .B2(n15174), .ZN(
        P2_U3510) );
  NOR2_X1 U16809 ( .A1(P3_U3897), .A2(n15326), .ZN(P3_U3150) );
  OAI21_X1 U16810 ( .B1(n15179), .B2(n15203), .A(n15178), .ZN(n15188) );
  NAND2_X1 U16811 ( .A1(n15181), .A2(n15180), .ZN(n15183) );
  AND2_X1 U16812 ( .A1(n15183), .A2(n15182), .ZN(n15186) );
  AOI211_X1 U16813 ( .C1(n15186), .C2(n15185), .A(n15207), .B(n15184), .ZN(
        n15187) );
  AOI211_X1 U16814 ( .C1(n15213), .C2(n15189), .A(n15188), .B(n15187), .ZN(
        n15190) );
  OAI21_X1 U16815 ( .B1(n15191), .B2(n15215), .A(n15190), .ZN(P3_U3157) );
  AOI22_X1 U16816 ( .A1(n15192), .A2(n15366), .B1(n12406), .B2(n15365), .ZN(
        n15340) );
  OAI22_X1 U16817 ( .A1(n15340), .A2(n15203), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n7665), .ZN(n15199) );
  OAI211_X1 U16818 ( .C1(n15196), .C2(n15195), .A(n15194), .B(n15193), .ZN(
        n15197) );
  INV_X1 U16819 ( .A(n15197), .ZN(n15198) );
  AOI211_X1 U16820 ( .C1(n15213), .C2(n15200), .A(n15199), .B(n15198), .ZN(
        n15201) );
  OAI21_X1 U16821 ( .B1(P3_REG3_REG_3__SCAN_IN), .B2(n15215), .A(n15201), .ZN(
        P3_U3158) );
  OAI21_X1 U16822 ( .B1(n15204), .B2(n15203), .A(n15202), .ZN(n15211) );
  INV_X1 U16823 ( .A(n15205), .ZN(n15206) );
  AOI211_X1 U16824 ( .C1(n15209), .C2(n15208), .A(n15207), .B(n15206), .ZN(
        n15210) );
  AOI211_X1 U16825 ( .C1(n15213), .C2(n15212), .A(n15211), .B(n15210), .ZN(
        n15214) );
  OAI21_X1 U16826 ( .B1(n15216), .B2(n15215), .A(n15214), .ZN(P3_U3179) );
  INV_X1 U16827 ( .A(n15217), .ZN(n15218) );
  NAND3_X1 U16828 ( .A1(n15220), .A2(n15219), .A3(n15218), .ZN(n15221) );
  AOI21_X1 U16829 ( .B1(n15222), .B2(n15221), .A(n15322), .ZN(n15230) );
  AOI21_X1 U16830 ( .B1(n10022), .B2(n15224), .A(n15223), .ZN(n15228) );
  XNOR2_X1 U16831 ( .A(n15226), .B(n15225), .ZN(n15227) );
  OAI22_X1 U16832 ( .A1(n15333), .A2(n15228), .B1(n15297), .B2(n15227), .ZN(
        n15229) );
  AOI211_X1 U16833 ( .C1(n15266), .C2(n15231), .A(n15230), .B(n15229), .ZN(
        n15233) );
  NAND2_X1 U16834 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_U3151), .ZN(n15232) );
  OAI211_X1 U16835 ( .C1(n15234), .C2(n15308), .A(n15233), .B(n15232), .ZN(
        P3_U3185) );
  AOI21_X1 U16836 ( .B1(n6817), .B2(n15236), .A(n15235), .ZN(n15251) );
  AND2_X1 U16837 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n15244) );
  OAI21_X1 U16838 ( .B1(n15239), .B2(n15238), .A(n15237), .ZN(n15240) );
  AOI22_X1 U16839 ( .A1(n15266), .A2(n15241), .B1(n15305), .B2(n15240), .ZN(
        n15242) );
  INV_X1 U16840 ( .A(n15242), .ZN(n15243) );
  AOI211_X1 U16841 ( .C1(P3_ADDR_REG_4__SCAN_IN), .C2(n15326), .A(n15244), .B(
        n15243), .ZN(n15250) );
  OAI21_X1 U16842 ( .B1(n15247), .B2(n15246), .A(n15245), .ZN(n15248) );
  NAND2_X1 U16843 ( .A1(n15329), .A2(n15248), .ZN(n15249) );
  OAI211_X1 U16844 ( .C1(n15251), .C2(n15333), .A(n15250), .B(n15249), .ZN(
        P3_U3186) );
  NAND2_X1 U16845 ( .A1(n15253), .A2(n15252), .ZN(n15254) );
  XNOR2_X1 U16846 ( .A(n15255), .B(n15254), .ZN(n15269) );
  AOI21_X1 U16847 ( .B1(n15258), .B2(n15257), .A(n15256), .ZN(n15259) );
  INV_X1 U16848 ( .A(n15259), .ZN(n15263) );
  OAI21_X1 U16849 ( .B1(n15261), .B2(P3_REG1_REG_5__SCAN_IN), .A(n15260), .ZN(
        n15262) );
  AOI22_X1 U16850 ( .A1(n15264), .A2(n15263), .B1(n15329), .B2(n15262), .ZN(
        n15268) );
  NAND2_X1 U16851 ( .A1(n15266), .A2(n15265), .ZN(n15267) );
  OAI211_X1 U16852 ( .C1(n15269), .C2(n15322), .A(n15268), .B(n15267), .ZN(
        n15270) );
  INV_X1 U16853 ( .A(n15270), .ZN(n15272) );
  NAND2_X1 U16854 ( .A1(P3_REG3_REG_5__SCAN_IN), .A2(P3_U3151), .ZN(n15271) );
  OAI211_X1 U16855 ( .C1(n15273), .C2(n15308), .A(n15272), .B(n15271), .ZN(
        P3_U3187) );
  AOI21_X1 U16856 ( .B1(n15276), .B2(n15275), .A(n15274), .ZN(n15287) );
  OAI21_X1 U16857 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n15278), .A(n15277), .ZN(
        n15281) );
  NOR2_X1 U16858 ( .A1(n15320), .A2(n15279), .ZN(n15280) );
  AOI21_X1 U16859 ( .B1(n15281), .B2(n15329), .A(n15280), .ZN(n15286) );
  XNOR2_X1 U16860 ( .A(n15283), .B(n15282), .ZN(n15284) );
  NAND2_X1 U16861 ( .A1(n15284), .A2(n15305), .ZN(n15285) );
  OAI211_X1 U16862 ( .C1(n15287), .C2(n15333), .A(n15286), .B(n15285), .ZN(
        n15288) );
  INV_X1 U16863 ( .A(n15288), .ZN(n15290) );
  OAI211_X1 U16864 ( .C1(n15291), .C2(n15308), .A(n15290), .B(n15289), .ZN(
        P3_U3189) );
  XNOR2_X1 U16865 ( .A(n15293), .B(n15292), .ZN(n15304) );
  XOR2_X1 U16866 ( .A(n15295), .B(n15294), .Z(n15298) );
  OAI22_X1 U16867 ( .A1(n15298), .A2(n15297), .B1(n15296), .B2(n15320), .ZN(
        n15303) );
  AOI21_X1 U16868 ( .B1(n6805), .B2(n15300), .A(n15299), .ZN(n15301) );
  NOR2_X1 U16869 ( .A1(n15301), .A2(n15333), .ZN(n15302) );
  AOI211_X1 U16870 ( .C1(n15305), .C2(n15304), .A(n15303), .B(n15302), .ZN(
        n15307) );
  OAI211_X1 U16871 ( .C1(n15309), .C2(n15308), .A(n15307), .B(n15306), .ZN(
        P3_U3190) );
  AOI21_X1 U16872 ( .B1(n15312), .B2(n15311), .A(n15310), .ZN(n15334) );
  NOR2_X1 U16873 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15313), .ZN(n15325) );
  INV_X1 U16874 ( .A(n15314), .ZN(n15319) );
  AOI21_X1 U16875 ( .B1(n15316), .B2(n15318), .A(n15315), .ZN(n15317) );
  AOI21_X1 U16876 ( .B1(n15319), .B2(n15318), .A(n15317), .ZN(n15323) );
  OAI22_X1 U16877 ( .A1(n15323), .A2(n15322), .B1(n15321), .B2(n15320), .ZN(
        n15324) );
  AOI211_X1 U16878 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n15326), .A(n15325), .B(
        n15324), .ZN(n15332) );
  OAI21_X1 U16879 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n15328), .A(n15327), .ZN(
        n15330) );
  NAND2_X1 U16880 ( .A1(n15330), .A2(n15329), .ZN(n15331) );
  OAI211_X1 U16881 ( .C1(n15334), .C2(n15333), .A(n15332), .B(n15331), .ZN(
        P3_U3191) );
  XOR2_X1 U16882 ( .A(n15336), .B(n15335), .Z(n15341) );
  INV_X1 U16883 ( .A(n15341), .ZN(n15393) );
  OAI211_X1 U16884 ( .C1(n6720), .C2(n15338), .A(n15369), .B(n15337), .ZN(
        n15339) );
  OAI211_X1 U16885 ( .C1(n15341), .C2(n15373), .A(n15340), .B(n15339), .ZN(
        n15391) );
  AOI21_X1 U16886 ( .B1(n15342), .B2(n15393), .A(n15391), .ZN(n15346) );
  NOR2_X1 U16887 ( .A1(n15343), .A2(n15374), .ZN(n15392) );
  AOI22_X1 U16888 ( .A1(n15344), .A2(n15392), .B1(n15379), .B2(n7665), .ZN(
        n15345) );
  OAI221_X1 U16889 ( .B1(n12443), .B2(n15346), .C1(n15380), .C2(n10022), .A(
        n15345), .ZN(P3_U3230) );
  XNOR2_X1 U16890 ( .A(n15347), .B(n15349), .ZN(n15358) );
  OAI21_X1 U16891 ( .B1(n15350), .B2(n15349), .A(n15348), .ZN(n15389) );
  OAI22_X1 U16892 ( .A1(n6846), .A2(n15353), .B1(n15352), .B2(n15351), .ZN(
        n15355) );
  AOI21_X1 U16893 ( .B1(n15389), .B2(n15356), .A(n15355), .ZN(n15357) );
  OAI21_X1 U16894 ( .B1(n15359), .B2(n15358), .A(n15357), .ZN(n15387) );
  INV_X1 U16895 ( .A(n15389), .ZN(n15362) );
  NOR2_X1 U16896 ( .A1(n15374), .A2(n15360), .ZN(n15388) );
  INV_X1 U16897 ( .A(n15388), .ZN(n15361) );
  OAI22_X1 U16898 ( .A1(n15362), .A2(n15377), .B1(n15376), .B2(n15361), .ZN(
        n15363) );
  AOI211_X1 U16899 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n15379), .A(n15387), .B(
        n15363), .ZN(n15364) );
  AOI22_X1 U16900 ( .A1(n12443), .A2(n10017), .B1(n15364), .B2(n15380), .ZN(
        P3_U3231) );
  AOI22_X1 U16901 ( .A1(n12406), .A2(n15367), .B1(n15366), .B2(n15365), .ZN(
        n15372) );
  NAND2_X1 U16902 ( .A1(n15370), .A2(n15369), .ZN(n15371) );
  OAI211_X1 U16903 ( .C1(n15382), .C2(n15373), .A(n15372), .B(n15371), .ZN(
        n15383) );
  NOR2_X1 U16904 ( .A1(n10214), .A2(n15374), .ZN(n15384) );
  INV_X1 U16905 ( .A(n15384), .ZN(n15375) );
  OAI22_X1 U16906 ( .A1(n15382), .A2(n15377), .B1(n15376), .B2(n15375), .ZN(
        n15378) );
  AOI211_X1 U16907 ( .C1(P3_REG3_REG_1__SCAN_IN), .C2(n15379), .A(n15383), .B(
        n15378), .ZN(n15381) );
  AOI22_X1 U16908 ( .A1(n12443), .A2(n10012), .B1(n15381), .B2(n15380), .ZN(
        P3_U3232) );
  INV_X1 U16909 ( .A(n15382), .ZN(n15385) );
  AOI211_X1 U16910 ( .C1(n15410), .C2(n15385), .A(n15384), .B(n15383), .ZN(
        n15422) );
  INV_X1 U16911 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15386) );
  AOI22_X1 U16912 ( .A1(n15421), .A2(n15422), .B1(n15386), .B2(n15419), .ZN(
        P3_U3393) );
  AOI211_X1 U16913 ( .C1(n15410), .C2(n15389), .A(n15388), .B(n15387), .ZN(
        n15423) );
  AOI22_X1 U16914 ( .A1(n15421), .A2(n15423), .B1(n15390), .B2(n15419), .ZN(
        P3_U3396) );
  AOI211_X1 U16915 ( .C1(n15393), .C2(n15410), .A(n15392), .B(n15391), .ZN(
        n15424) );
  INV_X1 U16916 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15394) );
  AOI22_X1 U16917 ( .A1(n15421), .A2(n15424), .B1(n15394), .B2(n15419), .ZN(
        P3_U3399) );
  INV_X1 U16918 ( .A(n15395), .ZN(n15397) );
  AOI211_X1 U16919 ( .C1(n15398), .C2(n15410), .A(n15397), .B(n15396), .ZN(
        n15426) );
  INV_X1 U16920 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15399) );
  AOI22_X1 U16921 ( .A1(n15421), .A2(n15426), .B1(n15399), .B2(n15419), .ZN(
        P3_U3408) );
  AOI211_X1 U16922 ( .C1(n15402), .C2(n15410), .A(n15401), .B(n15400), .ZN(
        n15428) );
  INV_X1 U16923 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15403) );
  AOI22_X1 U16924 ( .A1(n15421), .A2(n15428), .B1(n15403), .B2(n15419), .ZN(
        P3_U3411) );
  AOI211_X1 U16925 ( .C1(n15406), .C2(n15410), .A(n15405), .B(n15404), .ZN(
        n15430) );
  INV_X1 U16926 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15407) );
  AOI22_X1 U16927 ( .A1(n15421), .A2(n15430), .B1(n15407), .B2(n15419), .ZN(
        P3_U3414) );
  AOI211_X1 U16928 ( .C1(n15411), .C2(n15410), .A(n15409), .B(n15408), .ZN(
        n15432) );
  INV_X1 U16929 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15412) );
  AOI22_X1 U16930 ( .A1(n15421), .A2(n15432), .B1(n15412), .B2(n15419), .ZN(
        P3_U3417) );
  NOR2_X1 U16931 ( .A1(n15414), .A2(n15413), .ZN(n15418) );
  AOI211_X1 U16932 ( .C1(n15418), .C2(n15417), .A(n15416), .B(n15415), .ZN(
        n15435) );
  INV_X1 U16933 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15420) );
  AOI22_X1 U16934 ( .A1(n15421), .A2(n15435), .B1(n15420), .B2(n15419), .ZN(
        P3_U3420) );
  AOI22_X1 U16935 ( .A1(n15436), .A2(n15422), .B1(n10011), .B2(n15433), .ZN(
        P3_U3460) );
  AOI22_X1 U16936 ( .A1(n15436), .A2(n15423), .B1(n10016), .B2(n15433), .ZN(
        P3_U3461) );
  AOI22_X1 U16937 ( .A1(n15436), .A2(n15424), .B1(n15225), .B2(n15433), .ZN(
        P3_U3462) );
  AOI22_X1 U16938 ( .A1(n15436), .A2(n15426), .B1(n15425), .B2(n15433), .ZN(
        P3_U3465) );
  INV_X1 U16939 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15427) );
  AOI22_X1 U16940 ( .A1(n15436), .A2(n15428), .B1(n15427), .B2(n15433), .ZN(
        P3_U3466) );
  AOI22_X1 U16941 ( .A1(n15436), .A2(n15430), .B1(n15429), .B2(n15433), .ZN(
        P3_U3467) );
  INV_X1 U16942 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15431) );
  AOI22_X1 U16943 ( .A1(n15436), .A2(n15432), .B1(n15431), .B2(n15433), .ZN(
        P3_U3468) );
  AOI22_X1 U16944 ( .A1(n15436), .A2(n15435), .B1(n15434), .B2(n15433), .ZN(
        P3_U3469) );
  OAI21_X1 U16945 ( .B1(n6733), .B2(n15438), .A(n15437), .ZN(SUB_1596_U59) );
  OAI21_X1 U16946 ( .B1(n15441), .B2(n15440), .A(n15439), .ZN(SUB_1596_U58) );
  OAI21_X1 U16947 ( .B1(n15442), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n15453), .ZN(
        n15443) );
  INV_X1 U16948 ( .A(n15443), .ZN(SUB_1596_U53) );
  AOI21_X1 U16949 ( .B1(n15446), .B2(n15445), .A(n15444), .ZN(SUB_1596_U56) );
  AOI21_X1 U16950 ( .B1(n15449), .B2(n15448), .A(n15447), .ZN(n15450) );
  XOR2_X1 U16951 ( .A(n15450), .B(P2_ADDR_REG_3__SCAN_IN), .Z(SUB_1596_U60) );
  AOI21_X1 U16952 ( .B1(n15453), .B2(n15452), .A(n15451), .ZN(SUB_1596_U5) );
  MUX2_X1 U9908 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7617), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n7620) );
  CLKBUF_X2 U7367 ( .A(n8918), .Z(n9082) );
  NOR2_X1 U7375 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n6877) );
  CLKBUF_X2 U7393 ( .A(n13000), .Z(n6616) );
  AND4_X1 U7399 ( .A1(n6879), .A2(n6878), .A3(n6877), .A4(n8858), .ZN(n6876)
         );
  INV_X1 U7400 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8260) );
  AND2_X1 U7408 ( .A1(n8570), .A2(n8569), .ZN(n8573) );
  AND2_X1 U7409 ( .A1(n9164), .A2(n9162), .ZN(n10212) );
  CLKBUF_X1 U7483 ( .A(n12146), .Z(n6850) );
  NAND2_X1 U7487 ( .A1(n6608), .A2(n9486), .ZN(n7674) );
  CLKBUF_X1 U7503 ( .A(n6613), .Z(n12892) );
  CLKBUF_X1 U7788 ( .A(n10406), .Z(n13169) );
  NOR2_X2 U7802 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n9470) );
  CLKBUF_X1 U8112 ( .A(n8455), .Z(n9064) );
  CLKBUF_X1 U8485 ( .A(n8405), .Z(n9430) );
  CLKBUF_X1 U9461 ( .A(n10135), .Z(n12901) );
  CLKBUF_X1 U9462 ( .A(n9915), .Z(n11374) );
endmodule

